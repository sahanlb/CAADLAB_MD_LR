localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTZ_CHK = {
  {32'h44aee22e, 32'h45056a4a} /* (31, 31, 31) {real, imag} */,
  {32'hc469bb38, 32'hc42a540c} /* (31, 31, 30) {real, imag} */,
  {32'hc1ed377c, 32'hc2abf697} /* (31, 31, 29) {real, imag} */,
  {32'h43bf05ba, 32'h434c6156} /* (31, 31, 28) {real, imag} */,
  {32'hc383d7eb, 32'hc3a9eb88} /* (31, 31, 27) {real, imag} */,
  {32'hc2e27e31, 32'hc3852b92} /* (31, 31, 26) {real, imag} */,
  {32'hc19b0e8c, 32'h430f2998} /* (31, 31, 25) {real, imag} */,
  {32'hc36d59fe, 32'hc08f7240} /* (31, 31, 24) {real, imag} */,
  {32'hc0dca0d0, 32'hc212975a} /* (31, 31, 23) {real, imag} */,
  {32'hc30df27a, 32'hc2698c9c} /* (31, 31, 22) {real, imag} */,
  {32'hc333a85d, 32'h41bec440} /* (31, 31, 21) {real, imag} */,
  {32'hc2bbb80c, 32'hc1e11e30} /* (31, 31, 20) {real, imag} */,
  {32'h418cbd54, 32'hc17487d4} /* (31, 31, 19) {real, imag} */,
  {32'hc29746a2, 32'h422a8e30} /* (31, 31, 18) {real, imag} */,
  {32'h42725e30, 32'h40f12d80} /* (31, 31, 17) {real, imag} */,
  {32'hc175dfc0, 32'h412871c0} /* (31, 31, 16) {real, imag} */,
  {32'h410de2c0, 32'h41040140} /* (31, 31, 15) {real, imag} */,
  {32'h42262744, 32'hc183d560} /* (31, 31, 14) {real, imag} */,
  {32'hc18890bc, 32'h412dc4a4} /* (31, 31, 13) {real, imag} */,
  {32'hbfa17720, 32'hc1c6a150} /* (31, 31, 12) {real, imag} */,
  {32'h433427e7, 32'hc304a240} /* (31, 31, 11) {real, imag} */,
  {32'hc1fd246c, 32'h42a463c6} /* (31, 31, 10) {real, imag} */,
  {32'h4296f753, 32'hc26da69e} /* (31, 31, 9) {real, imag} */,
  {32'h4346baa2, 32'hc3468e96} /* (31, 31, 8) {real, imag} */,
  {32'hc26cf686, 32'h4363589e} /* (31, 31, 7) {real, imag} */,
  {32'hc2b3a163, 32'h40039b40} /* (31, 31, 6) {real, imag} */,
  {32'hc308860c, 32'hc40afaa0} /* (31, 31, 5) {real, imag} */,
  {32'h436ae8c0, 32'h43851d1b} /* (31, 31, 4) {real, imag} */,
  {32'h42f61791, 32'h428da4a9} /* (31, 31, 3) {real, imag} */,
  {32'hc30214a0, 32'hc42518a0} /* (31, 31, 2) {real, imag} */,
  {32'hc35bce04, 32'h44c5580c} /* (31, 31, 1) {real, imag} */,
  {32'h439a3b04, 32'h44a3775c} /* (31, 31, 0) {real, imag} */,
  {32'hc1d02f30, 32'hc49b2789} /* (31, 30, 31) {real, imag} */,
  {32'h411c0840, 32'h4449d71d} /* (31, 30, 30) {real, imag} */,
  {32'hc210f13c, 32'h41d90f62} /* (31, 30, 29) {real, imag} */,
  {32'hc34240cb, 32'hc414b23e} /* (31, 30, 28) {real, imag} */,
  {32'h43edc3cf, 32'h43dee1c2} /* (31, 30, 27) {real, imag} */,
  {32'h41c73c40, 32'h42c7d336} /* (31, 30, 26) {real, imag} */,
  {32'hc23677b0, 32'hc2f1213e} /* (31, 30, 25) {real, imag} */,
  {32'hc27be38e, 32'hc10059bc} /* (31, 30, 24) {real, imag} */,
  {32'h42cc6eb0, 32'h40174080} /* (31, 30, 23) {real, imag} */,
  {32'h41a03630, 32'hc20fc229} /* (31, 30, 22) {real, imag} */,
  {32'h43318582, 32'hc1307034} /* (31, 30, 21) {real, imag} */,
  {32'h421e5de8, 32'h4226ef4a} /* (31, 30, 20) {real, imag} */,
  {32'h40c5b580, 32'h4189ad22} /* (31, 30, 19) {real, imag} */,
  {32'h4172ce8c, 32'h42086b14} /* (31, 30, 18) {real, imag} */,
  {32'hc0990a28, 32'hc153fd70} /* (31, 30, 17) {real, imag} */,
  {32'hc175f6b0, 32'h41f09bf0} /* (31, 30, 16) {real, imag} */,
  {32'h42892af6, 32'hc1c209c8} /* (31, 30, 15) {real, imag} */,
  {32'hc2ab9846, 32'h3e3bec00} /* (31, 30, 14) {real, imag} */,
  {32'h416ff148, 32'h4298cee6} /* (31, 30, 13) {real, imag} */,
  {32'hc1828b0f, 32'hc224341a} /* (31, 30, 12) {real, imag} */,
  {32'hc284c849, 32'h41f5daea} /* (31, 30, 11) {real, imag} */,
  {32'h42774102, 32'h429a4e1c} /* (31, 30, 10) {real, imag} */,
  {32'h42b2c984, 32'hc28368db} /* (31, 30, 9) {real, imag} */,
  {32'hc232dd96, 32'h41b4ccfe} /* (31, 30, 8) {real, imag} */,
  {32'hc2de213c, 32'hc314395d} /* (31, 30, 7) {real, imag} */,
  {32'hc2b34a95, 32'h4218d265} /* (31, 30, 6) {real, imag} */,
  {32'hc2cc0464, 32'h4339e87d} /* (31, 30, 5) {real, imag} */,
  {32'h435ee2b1, 32'hc3462bb4} /* (31, 30, 4) {real, imag} */,
  {32'h42962399, 32'hc149e4b4} /* (31, 30, 3) {real, imag} */,
  {32'hc332d4f8, 32'h44ad535e} /* (31, 30, 2) {real, imag} */,
  {32'hc38e423c, 32'hc500541e} /* (31, 30, 1) {real, imag} */,
  {32'hc38e1240, 32'hc457ec80} /* (31, 30, 0) {real, imag} */,
  {32'h438588fd, 32'h434b8050} /* (31, 29, 31) {real, imag} */,
  {32'hc3b8a910, 32'hc210c644} /* (31, 29, 30) {real, imag} */,
  {32'hc2385564, 32'hc2c25bec} /* (31, 29, 29) {real, imag} */,
  {32'h42a992db, 32'hc3775e66} /* (31, 29, 28) {real, imag} */,
  {32'h420ef24f, 32'h42995e08} /* (31, 29, 27) {real, imag} */,
  {32'hc34d37b4, 32'h4328f63e} /* (31, 29, 26) {real, imag} */,
  {32'hc2735708, 32'hc227e5d6} /* (31, 29, 25) {real, imag} */,
  {32'h41ae92b6, 32'hc097a5f8} /* (31, 29, 24) {real, imag} */,
  {32'h42e3e133, 32'hc23543c8} /* (31, 29, 23) {real, imag} */,
  {32'hc1e70750, 32'h42821767} /* (31, 29, 22) {real, imag} */,
  {32'hc23cfe2f, 32'h426e8187} /* (31, 29, 21) {real, imag} */,
  {32'h423508b9, 32'h4147e3d1} /* (31, 29, 20) {real, imag} */,
  {32'hc0abf5ac, 32'h41dea6e4} /* (31, 29, 19) {real, imag} */,
  {32'hc223f5a6, 32'h4117cc58} /* (31, 29, 18) {real, imag} */,
  {32'h41db9841, 32'h411f6164} /* (31, 29, 17) {real, imag} */,
  {32'hc217f6e5, 32'h40124100} /* (31, 29, 16) {real, imag} */,
  {32'h422fe27c, 32'h428786c8} /* (31, 29, 15) {real, imag} */,
  {32'hc238809a, 32'hc1aee85c} /* (31, 29, 14) {real, imag} */,
  {32'h41569752, 32'hc1700ae8} /* (31, 29, 13) {real, imag} */,
  {32'h411fe324, 32'hc13b623f} /* (31, 29, 12) {real, imag} */,
  {32'hc25e01ad, 32'h4198a956} /* (31, 29, 11) {real, imag} */,
  {32'h42bf6f56, 32'hc2a86f87} /* (31, 29, 10) {real, imag} */,
  {32'h41ed2aec, 32'h41e426f9} /* (31, 29, 9) {real, imag} */,
  {32'hc30e3355, 32'hc27fac37} /* (31, 29, 8) {real, imag} */,
  {32'h42b39b60, 32'h41fb35bb} /* (31, 29, 7) {real, imag} */,
  {32'h424e7562, 32'hc2a529d5} /* (31, 29, 6) {real, imag} */,
  {32'h42bd5bb6, 32'hc2e55d56} /* (31, 29, 5) {real, imag} */,
  {32'h430edb2e, 32'h43427ad2} /* (31, 29, 4) {real, imag} */,
  {32'h42a69bc6, 32'h40ba0920} /* (31, 29, 3) {real, imag} */,
  {32'hc3e80cb8, 32'h43b69bec} /* (31, 29, 2) {real, imag} */,
  {32'h431a3c92, 32'hc3cc4450} /* (31, 29, 1) {real, imag} */,
  {32'h417f378c, 32'hc2c1a6eb} /* (31, 29, 0) {real, imag} */,
  {32'h4252a020, 32'h43bba6dd} /* (31, 28, 31) {real, imag} */,
  {32'hc3af3ab7, 32'hc3c64541} /* (31, 28, 30) {real, imag} */,
  {32'h438aaee5, 32'hc33f032c} /* (31, 28, 29) {real, imag} */,
  {32'h438ccde8, 32'hc2bb54da} /* (31, 28, 28) {real, imag} */,
  {32'hc2b1f275, 32'h4204f2d3} /* (31, 28, 27) {real, imag} */,
  {32'h4296bfda, 32'h431a8b65} /* (31, 28, 26) {real, imag} */,
  {32'hc0943368, 32'hc0a8d3c0} /* (31, 28, 25) {real, imag} */,
  {32'hc3143de2, 32'hc31a4b6b} /* (31, 28, 24) {real, imag} */,
  {32'h41a356b6, 32'h420a0e34} /* (31, 28, 23) {real, imag} */,
  {32'hc2310815, 32'hc12dfee8} /* (31, 28, 22) {real, imag} */,
  {32'hc2d3f798, 32'hc2028f55} /* (31, 28, 21) {real, imag} */,
  {32'h42f26024, 32'h4214f70f} /* (31, 28, 20) {real, imag} */,
  {32'h41c9e494, 32'h41151cac} /* (31, 28, 19) {real, imag} */,
  {32'hc295448e, 32'hc18dd086} /* (31, 28, 18) {real, imag} */,
  {32'hc0d0e3e0, 32'hc183e9ac} /* (31, 28, 17) {real, imag} */,
  {32'h418e5828, 32'h42127f1e} /* (31, 28, 16) {real, imag} */,
  {32'h41f4daa8, 32'h418e50ac} /* (31, 28, 15) {real, imag} */,
  {32'hc1f773ea, 32'hc216cc85} /* (31, 28, 14) {real, imag} */,
  {32'hc128ec28, 32'hc2651cc5} /* (31, 28, 13) {real, imag} */,
  {32'h423856bf, 32'hc08cce48} /* (31, 28, 12) {real, imag} */,
  {32'h41dfbdf8, 32'h42837e7a} /* (31, 28, 11) {real, imag} */,
  {32'hc1ef79a6, 32'h4061de20} /* (31, 28, 10) {real, imag} */,
  {32'hc2908586, 32'h4248c4fc} /* (31, 28, 9) {real, imag} */,
  {32'hc37b328c, 32'hc2fd723a} /* (31, 28, 8) {real, imag} */,
  {32'hc21a62c9, 32'h432f2772} /* (31, 28, 7) {real, imag} */,
  {32'h42e63a0a, 32'hc1cec228} /* (31, 28, 6) {real, imag} */,
  {32'hc18b7804, 32'hc30ba94b} /* (31, 28, 5) {real, imag} */,
  {32'h433b008e, 32'h43873a94} /* (31, 28, 4) {real, imag} */,
  {32'hc24883e8, 32'hc2c7edbc} /* (31, 28, 3) {real, imag} */,
  {32'hc3cb132d, 32'hc3f8aba3} /* (31, 28, 2) {real, imag} */,
  {32'h43af03ac, 32'hc24b0d08} /* (31, 28, 1) {real, imag} */,
  {32'h431b5d25, 32'h4317dda6} /* (31, 28, 0) {real, imag} */,
  {32'hc3c41de1, 32'hc2fb26d4} /* (31, 27, 31) {real, imag} */,
  {32'h43f16f63, 32'h428d178c} /* (31, 27, 30) {real, imag} */,
  {32'h421c567c, 32'h4121ca1f} /* (31, 27, 29) {real, imag} */,
  {32'hc3766d3a, 32'hc19f2f96} /* (31, 27, 28) {real, imag} */,
  {32'h4268e23e, 32'h43252edb} /* (31, 27, 27) {real, imag} */,
  {32'h421c768c, 32'hc20bf6c1} /* (31, 27, 26) {real, imag} */,
  {32'hc2e774a8, 32'hc2d82774} /* (31, 27, 25) {real, imag} */,
  {32'hc1b978c0, 32'h420a04f9} /* (31, 27, 24) {real, imag} */,
  {32'h425bff98, 32'hc2196fa2} /* (31, 27, 23) {real, imag} */,
  {32'h42b05481, 32'hc10500dc} /* (31, 27, 22) {real, imag} */,
  {32'h3f283fc0, 32'h42435bf4} /* (31, 27, 21) {real, imag} */,
  {32'hc207e6a6, 32'hc1215029} /* (31, 27, 20) {real, imag} */,
  {32'h41bacf55, 32'h4164d740} /* (31, 27, 19) {real, imag} */,
  {32'h423c43d4, 32'h4145f258} /* (31, 27, 18) {real, imag} */,
  {32'hc2248974, 32'h42016b10} /* (31, 27, 17) {real, imag} */,
  {32'hc12086c0, 32'h419ef260} /* (31, 27, 16) {real, imag} */,
  {32'hc1ec1130, 32'h40af7d80} /* (31, 27, 15) {real, imag} */,
  {32'hc292856e, 32'hc249e69a} /* (31, 27, 14) {real, imag} */,
  {32'h41eca6d7, 32'hc1cb9320} /* (31, 27, 13) {real, imag} */,
  {32'h407d94a0, 32'hc216a33a} /* (31, 27, 12) {real, imag} */,
  {32'hc23ccccc, 32'h41345c00} /* (31, 27, 11) {real, imag} */,
  {32'hc1fa4c93, 32'hbe408b00} /* (31, 27, 10) {real, imag} */,
  {32'h3e563080, 32'h41e1bb00} /* (31, 27, 9) {real, imag} */,
  {32'hc2d12114, 32'hc21f2cbf} /* (31, 27, 8) {real, imag} */,
  {32'h42473b88, 32'hc25e5bb1} /* (31, 27, 7) {real, imag} */,
  {32'h42ae2ef2, 32'h4283e432} /* (31, 27, 6) {real, imag} */,
  {32'h42ae1ec9, 32'h431b092d} /* (31, 27, 5) {real, imag} */,
  {32'h4291afbc, 32'h41f57c7a} /* (31, 27, 4) {real, imag} */,
  {32'hc22170b8, 32'h4190c4b0} /* (31, 27, 3) {real, imag} */,
  {32'h42969914, 32'h43901265} /* (31, 27, 2) {real, imag} */,
  {32'hc1db0990, 32'hc3cd3627} /* (31, 27, 1) {real, imag} */,
  {32'hc34884ca, 32'hc3144cbc} /* (31, 27, 0) {real, imag} */,
  {32'hc29325b3, 32'h4220501c} /* (31, 26, 31) {real, imag} */,
  {32'hc31d2b10, 32'hc2642998} /* (31, 26, 30) {real, imag} */,
  {32'h4242d701, 32'hc2eee06b} /* (31, 26, 29) {real, imag} */,
  {32'h427c825d, 32'h4256fd6c} /* (31, 26, 28) {real, imag} */,
  {32'hc0417d60, 32'hc2927f71} /* (31, 26, 27) {real, imag} */,
  {32'h403041ec, 32'hc2bfce51} /* (31, 26, 26) {real, imag} */,
  {32'h42b04220, 32'h421e5eca} /* (31, 26, 25) {real, imag} */,
  {32'h3fc764b0, 32'h417e7220} /* (31, 26, 24) {real, imag} */,
  {32'h42cefd75, 32'hc2d18e23} /* (31, 26, 23) {real, imag} */,
  {32'h41a0f210, 32'h429a249f} /* (31, 26, 22) {real, imag} */,
  {32'h411eb18f, 32'h4289e550} /* (31, 26, 21) {real, imag} */,
  {32'hc22c3a64, 32'hbf412dc0} /* (31, 26, 20) {real, imag} */,
  {32'h3f9495a0, 32'hc19b36b3} /* (31, 26, 19) {real, imag} */,
  {32'hc1c8ed14, 32'hc083940e} /* (31, 26, 18) {real, imag} */,
  {32'hc21f8e86, 32'h414688c4} /* (31, 26, 17) {real, imag} */,
  {32'h41c35420, 32'hc12074de} /* (31, 26, 16) {real, imag} */,
  {32'hc202a836, 32'hc1c9b2e8} /* (31, 26, 15) {real, imag} */,
  {32'h410e0ce8, 32'hc18ad092} /* (31, 26, 14) {real, imag} */,
  {32'h422b4863, 32'h424b79b2} /* (31, 26, 13) {real, imag} */,
  {32'hc0510cb0, 32'hc2603589} /* (31, 26, 12) {real, imag} */,
  {32'hc18f8bba, 32'h428a7da2} /* (31, 26, 11) {real, imag} */,
  {32'hc017d62c, 32'h41633ee6} /* (31, 26, 10) {real, imag} */,
  {32'hc24381a6, 32'h42c9d879} /* (31, 26, 9) {real, imag} */,
  {32'h4275a856, 32'hc2c2d044} /* (31, 26, 8) {real, imag} */,
  {32'h4201c5d7, 32'hc20a9d40} /* (31, 26, 7) {real, imag} */,
  {32'h41b60438, 32'h4294a5b1} /* (31, 26, 6) {real, imag} */,
  {32'h42a4f2cd, 32'h42c56e33} /* (31, 26, 5) {real, imag} */,
  {32'hc2bd807f, 32'hc14ee570} /* (31, 26, 4) {real, imag} */,
  {32'h42b6e28a, 32'h41bd9dfc} /* (31, 26, 3) {real, imag} */,
  {32'hc307a412, 32'h4000b6f8} /* (31, 26, 2) {real, imag} */,
  {32'hc2960809, 32'hc29c3448} /* (31, 26, 1) {real, imag} */,
  {32'h431c801d, 32'h428cc446} /* (31, 26, 0) {real, imag} */,
  {32'h4389e06f, 32'h42b026b4} /* (31, 25, 31) {real, imag} */,
  {32'hc3330734, 32'hc2bf21fe} /* (31, 25, 30) {real, imag} */,
  {32'hc2020058, 32'hc291487e} /* (31, 25, 29) {real, imag} */,
  {32'h427019fc, 32'h4045f1e8} /* (31, 25, 28) {real, imag} */,
  {32'h42d65881, 32'h41e549c5} /* (31, 25, 27) {real, imag} */,
  {32'hc2392445, 32'hc247d89d} /* (31, 25, 26) {real, imag} */,
  {32'h427dbfb6, 32'h42443134} /* (31, 25, 25) {real, imag} */,
  {32'h41c22c35, 32'hc228dfb0} /* (31, 25, 24) {real, imag} */,
  {32'h430e6762, 32'hc1fa55ec} /* (31, 25, 23) {real, imag} */,
  {32'h42320cdd, 32'h42b160b4} /* (31, 25, 22) {real, imag} */,
  {32'hc1a8bec0, 32'h425b007c} /* (31, 25, 21) {real, imag} */,
  {32'hc22c496e, 32'hc11b638e} /* (31, 25, 20) {real, imag} */,
  {32'hc08822a4, 32'hc26aba3e} /* (31, 25, 19) {real, imag} */,
  {32'hc1223dd9, 32'h41ded4e0} /* (31, 25, 18) {real, imag} */,
  {32'h406a60c0, 32'hc000f2c2} /* (31, 25, 17) {real, imag} */,
  {32'h41cb9550, 32'hc123cc70} /* (31, 25, 16) {real, imag} */,
  {32'h416d6560, 32'hc12cb390} /* (31, 25, 15) {real, imag} */,
  {32'hc19df544, 32'h41a2f7f8} /* (31, 25, 14) {real, imag} */,
  {32'h418f3ebb, 32'h40d23174} /* (31, 25, 13) {real, imag} */,
  {32'hc1a4d03c, 32'h41c5a7b1} /* (31, 25, 12) {real, imag} */,
  {32'h4134756c, 32'hc1a73cf8} /* (31, 25, 11) {real, imag} */,
  {32'h42053ccb, 32'h4228d0c5} /* (31, 25, 10) {real, imag} */,
  {32'hc28f01cd, 32'hc3083f10} /* (31, 25, 9) {real, imag} */,
  {32'hc1b7bfe5, 32'hc1ea80b8} /* (31, 25, 8) {real, imag} */,
  {32'hc1eda525, 32'h41de9bd9} /* (31, 25, 7) {real, imag} */,
  {32'h42497c81, 32'hc130da7c} /* (31, 25, 6) {real, imag} */,
  {32'h41180928, 32'h4142b73e} /* (31, 25, 5) {real, imag} */,
  {32'hc2a6bcdc, 32'hc1b1b8eb} /* (31, 25, 4) {real, imag} */,
  {32'h41e47f5c, 32'hc2bf1342} /* (31, 25, 3) {real, imag} */,
  {32'hc31c3aa2, 32'hc31d68a2} /* (31, 25, 2) {real, imag} */,
  {32'h41a3916c, 32'h42f64628} /* (31, 25, 1) {real, imag} */,
  {32'h434464ac, 32'h427057d4} /* (31, 25, 0) {real, imag} */,
  {32'hc31045fa, 32'hc3087120} /* (31, 24, 31) {real, imag} */,
  {32'h429bee5f, 32'h4360a0c1} /* (31, 24, 30) {real, imag} */,
  {32'hc14025ca, 32'hc0f4f228} /* (31, 24, 29) {real, imag} */,
  {32'hc307f4ef, 32'hc33296ab} /* (31, 24, 28) {real, imag} */,
  {32'h42c3dd96, 32'h41fa3858} /* (31, 24, 27) {real, imag} */,
  {32'hc2e57110, 32'hc22cbbb5} /* (31, 24, 26) {real, imag} */,
  {32'h429efa44, 32'hc219b3fe} /* (31, 24, 25) {real, imag} */,
  {32'h42ac586f, 32'h429f9ebb} /* (31, 24, 24) {real, imag} */,
  {32'h42355328, 32'hc1f9132d} /* (31, 24, 23) {real, imag} */,
  {32'h41a7b7a6, 32'h421e1118} /* (31, 24, 22) {real, imag} */,
  {32'hc208a511, 32'hc1f810ba} /* (31, 24, 21) {real, imag} */,
  {32'hc14460a4, 32'h41ef9dc4} /* (31, 24, 20) {real, imag} */,
  {32'h4227db64, 32'hc1637ecd} /* (31, 24, 19) {real, imag} */,
  {32'hc08badd3, 32'hbfb8a840} /* (31, 24, 18) {real, imag} */,
  {32'h4192a7f4, 32'hc1cbb3c5} /* (31, 24, 17) {real, imag} */,
  {32'h41a432fc, 32'h41cf8da0} /* (31, 24, 16) {real, imag} */,
  {32'h41645777, 32'hc20c1152} /* (31, 24, 15) {real, imag} */,
  {32'hbfb6a734, 32'h4244c38a} /* (31, 24, 14) {real, imag} */,
  {32'h408cad2c, 32'hc165c9d3} /* (31, 24, 13) {real, imag} */,
  {32'h40341030, 32'h41de7a08} /* (31, 24, 12) {real, imag} */,
  {32'h41d5578e, 32'h4117bd44} /* (31, 24, 11) {real, imag} */,
  {32'h420785ed, 32'h421e6c16} /* (31, 24, 10) {real, imag} */,
  {32'hc154f35a, 32'h420b6ace} /* (31, 24, 9) {real, imag} */,
  {32'hc15d1198, 32'hc2a72a15} /* (31, 24, 8) {real, imag} */,
  {32'h427440bb, 32'hc290e3a9} /* (31, 24, 7) {real, imag} */,
  {32'h428718a4, 32'h41fd1de6} /* (31, 24, 6) {real, imag} */,
  {32'hc27133ec, 32'h438fe8f2} /* (31, 24, 5) {real, imag} */,
  {32'h422d8761, 32'h422c64a4} /* (31, 24, 4) {real, imag} */,
  {32'h41ee5f69, 32'hc22e453f} /* (31, 24, 3) {real, imag} */,
  {32'h42319f12, 32'h43140f39} /* (31, 24, 2) {real, imag} */,
  {32'hc341e188, 32'hc388f062} /* (31, 24, 1) {real, imag} */,
  {32'hc2eba7dd, 32'hc2ee221e} /* (31, 24, 0) {real, imag} */,
  {32'h4300b88f, 32'h426ee25d} /* (31, 23, 31) {real, imag} */,
  {32'hc28ee069, 32'h42f40aae} /* (31, 23, 30) {real, imag} */,
  {32'h4120e8bc, 32'h41e28043} /* (31, 23, 29) {real, imag} */,
  {32'h42a46d48, 32'hc1ca7db0} /* (31, 23, 28) {real, imag} */,
  {32'hc2c14421, 32'hc2a77ef0} /* (31, 23, 27) {real, imag} */,
  {32'h40ce164c, 32'hc2c697a3} /* (31, 23, 26) {real, imag} */,
  {32'h4296ab8e, 32'h41b04e34} /* (31, 23, 25) {real, imag} */,
  {32'h41e0365c, 32'hc0115278} /* (31, 23, 24) {real, imag} */,
  {32'h410f0604, 32'hc121119e} /* (31, 23, 23) {real, imag} */,
  {32'hc17de771, 32'h41b44600} /* (31, 23, 22) {real, imag} */,
  {32'hc21df98b, 32'h412b5e18} /* (31, 23, 21) {real, imag} */,
  {32'h410e7bae, 32'hc18a5c59} /* (31, 23, 20) {real, imag} */,
  {32'hbe16b380, 32'h4179b3bc} /* (31, 23, 19) {real, imag} */,
  {32'hc200eb3a, 32'hc16faa3e} /* (31, 23, 18) {real, imag} */,
  {32'hc0deee40, 32'hc22bcfd4} /* (31, 23, 17) {real, imag} */,
  {32'h42414cfe, 32'h40736ee0} /* (31, 23, 16) {real, imag} */,
  {32'h42123726, 32'h419c849b} /* (31, 23, 15) {real, imag} */,
  {32'hc082d1c8, 32'hc1b76ea5} /* (31, 23, 14) {real, imag} */,
  {32'hc21200f2, 32'hc1a13c92} /* (31, 23, 13) {real, imag} */,
  {32'h41da9b23, 32'h413a7cca} /* (31, 23, 12) {real, imag} */,
  {32'h407e1b50, 32'h41b3e658} /* (31, 23, 11) {real, imag} */,
  {32'hc1a002a6, 32'h41885af4} /* (31, 23, 10) {real, imag} */,
  {32'hc1d50526, 32'h424145b0} /* (31, 23, 9) {real, imag} */,
  {32'hc223bda6, 32'h4208c2cc} /* (31, 23, 8) {real, imag} */,
  {32'hc1448d64, 32'hc0a78bea} /* (31, 23, 7) {real, imag} */,
  {32'hc1f09665, 32'h42ddc9cd} /* (31, 23, 6) {real, imag} */,
  {32'h4207a0fe, 32'hc2c3eb28} /* (31, 23, 5) {real, imag} */,
  {32'hc188c80a, 32'h41e37712} /* (31, 23, 4) {real, imag} */,
  {32'hc2b00d74, 32'h40937d34} /* (31, 23, 3) {real, imag} */,
  {32'hc1c3468d, 32'h406de730} /* (31, 23, 2) {real, imag} */,
  {32'h424e4433, 32'hc2bb9f4a} /* (31, 23, 1) {real, imag} */,
  {32'hc3452506, 32'hc29a2a7b} /* (31, 23, 0) {real, imag} */,
  {32'h425a6777, 32'h42ba254a} /* (31, 22, 31) {real, imag} */,
  {32'hc2f2b96d, 32'h41817f56} /* (31, 22, 30) {real, imag} */,
  {32'h42487475, 32'hbe834500} /* (31, 22, 29) {real, imag} */,
  {32'h42a85f56, 32'hc1dd0c14} /* (31, 22, 28) {real, imag} */,
  {32'hc2c22bee, 32'h42b42088} /* (31, 22, 27) {real, imag} */,
  {32'h42303f0c, 32'h41f29432} /* (31, 22, 26) {real, imag} */,
  {32'h4267590b, 32'hbfafa060} /* (31, 22, 25) {real, imag} */,
  {32'h4085ca34, 32'h423ae7aa} /* (31, 22, 24) {real, imag} */,
  {32'h4186dca2, 32'hbd11a400} /* (31, 22, 23) {real, imag} */,
  {32'hc1be5216, 32'hc21a2037} /* (31, 22, 22) {real, imag} */,
  {32'hc1eba776, 32'h422074ae} /* (31, 22, 21) {real, imag} */,
  {32'h3fddf8a0, 32'h41da2302} /* (31, 22, 20) {real, imag} */,
  {32'h4024b0e0, 32'hc0c474de} /* (31, 22, 19) {real, imag} */,
  {32'h40a3a82a, 32'hc0e9046c} /* (31, 22, 18) {real, imag} */,
  {32'h41fa5521, 32'h4102a849} /* (31, 22, 17) {real, imag} */,
  {32'h41467746, 32'hc117d14d} /* (31, 22, 16) {real, imag} */,
  {32'hc15f9ed6, 32'h419e2d30} /* (31, 22, 15) {real, imag} */,
  {32'hc10128bd, 32'hc0cd123c} /* (31, 22, 14) {real, imag} */,
  {32'h420de142, 32'hc182fa3a} /* (31, 22, 13) {real, imag} */,
  {32'hc0d28038, 32'hc23d0f89} /* (31, 22, 12) {real, imag} */,
  {32'hc24215eb, 32'h41fa71e7} /* (31, 22, 11) {real, imag} */,
  {32'h42000927, 32'hc08d4248} /* (31, 22, 10) {real, imag} */,
  {32'hc2402403, 32'h4221be2d} /* (31, 22, 9) {real, imag} */,
  {32'h412f56e4, 32'h419eabdd} /* (31, 22, 8) {real, imag} */,
  {32'h41af071e, 32'h4131bc86} /* (31, 22, 7) {real, imag} */,
  {32'h424c6d40, 32'h42862900} /* (31, 22, 6) {real, imag} */,
  {32'h42d69fea, 32'h413b80d4} /* (31, 22, 5) {real, imag} */,
  {32'h42636854, 32'h428ee754} /* (31, 22, 4) {real, imag} */,
  {32'h421f50ab, 32'hc2a0e393} /* (31, 22, 3) {real, imag} */,
  {32'hc2d87b5b, 32'hc2d562ca} /* (31, 22, 2) {real, imag} */,
  {32'h42a1f924, 32'h4255dd35} /* (31, 22, 1) {real, imag} */,
  {32'h41ef7455, 32'h41d97a7e} /* (31, 22, 0) {real, imag} */,
  {32'hc304efa7, 32'hc24b3317} /* (31, 21, 31) {real, imag} */,
  {32'h42a43401, 32'hc277ad3b} /* (31, 21, 30) {real, imag} */,
  {32'h41ee98a9, 32'hc1d9adca} /* (31, 21, 29) {real, imag} */,
  {32'hc253304d, 32'h41d2de78} /* (31, 21, 28) {real, imag} */,
  {32'h42074e18, 32'hc19d220e} /* (31, 21, 27) {real, imag} */,
  {32'hc1cd4165, 32'h422fc008} /* (31, 21, 26) {real, imag} */,
  {32'hbfd48870, 32'h41966c2a} /* (31, 21, 25) {real, imag} */,
  {32'h409ed5d3, 32'h42019452} /* (31, 21, 24) {real, imag} */,
  {32'hc19de350, 32'h413a3f43} /* (31, 21, 23) {real, imag} */,
  {32'hc1a1b892, 32'hc236bc46} /* (31, 21, 22) {real, imag} */,
  {32'hc124eefe, 32'hc207eb66} /* (31, 21, 21) {real, imag} */,
  {32'hbfafb5a0, 32'h3f9ba914} /* (31, 21, 20) {real, imag} */,
  {32'hc190e9f7, 32'h408ecd62} /* (31, 21, 19) {real, imag} */,
  {32'h410ed309, 32'h40bc9cf2} /* (31, 21, 18) {real, imag} */,
  {32'hc108b458, 32'h4173777c} /* (31, 21, 17) {real, imag} */,
  {32'h413e3f90, 32'h3ec713f0} /* (31, 21, 16) {real, imag} */,
  {32'h40a82e30, 32'h41231d44} /* (31, 21, 15) {real, imag} */,
  {32'hc0c4ac32, 32'h3eac0020} /* (31, 21, 14) {real, imag} */,
  {32'hc0ff13e3, 32'hc0441dd4} /* (31, 21, 13) {real, imag} */,
  {32'h41441d6a, 32'h41278238} /* (31, 21, 12) {real, imag} */,
  {32'h41644246, 32'h41df5f68} /* (31, 21, 11) {real, imag} */,
  {32'hc213e61b, 32'hc18f1fbd} /* (31, 21, 10) {real, imag} */,
  {32'hc04a0130, 32'hc210e139} /* (31, 21, 9) {real, imag} */,
  {32'hc0ecbdb3, 32'h40d71a68} /* (31, 21, 8) {real, imag} */,
  {32'hc14b00fa, 32'hc2a9f242} /* (31, 21, 7) {real, imag} */,
  {32'h41ae376f, 32'hc0e97dac} /* (31, 21, 6) {real, imag} */,
  {32'hc0881754, 32'h42a7b84e} /* (31, 21, 5) {real, imag} */,
  {32'h41ba1ae2, 32'h4110126f} /* (31, 21, 4) {real, imag} */,
  {32'h40b354fc, 32'hc2862c54} /* (31, 21, 3) {real, imag} */,
  {32'h42cdcf1d, 32'h42c3f802} /* (31, 21, 2) {real, imag} */,
  {32'hc19646e0, 32'hc30e093a} /* (31, 21, 1) {real, imag} */,
  {32'hc2e00824, 32'hc0e2f4ef} /* (31, 21, 0) {real, imag} */,
  {32'hc28b8a2c, 32'h422640cb} /* (31, 20, 31) {real, imag} */,
  {32'h41b3c308, 32'h41e31ed0} /* (31, 20, 30) {real, imag} */,
  {32'h410590aa, 32'hc27ffcb9} /* (31, 20, 29) {real, imag} */,
  {32'hc1b2b2a8, 32'hc1007c9c} /* (31, 20, 28) {real, imag} */,
  {32'hbfade358, 32'h426175e6} /* (31, 20, 27) {real, imag} */,
  {32'h41bda31c, 32'hbf4dac10} /* (31, 20, 26) {real, imag} */,
  {32'hc181c80f, 32'hc20d510a} /* (31, 20, 25) {real, imag} */,
  {32'hc22db9e7, 32'hbf23fbc8} /* (31, 20, 24) {real, imag} */,
  {32'h421adf06, 32'h4287c9b9} /* (31, 20, 23) {real, imag} */,
  {32'hc0a6bbfc, 32'h4231d5a4} /* (31, 20, 22) {real, imag} */,
  {32'hc1da9f96, 32'h4181605a} /* (31, 20, 21) {real, imag} */,
  {32'hc0c375b8, 32'hc0e12750} /* (31, 20, 20) {real, imag} */,
  {32'hbfe47798, 32'hc186fce6} /* (31, 20, 19) {real, imag} */,
  {32'h3ff0b960, 32'hc0a3a71b} /* (31, 20, 18) {real, imag} */,
  {32'hc0b7f6b4, 32'hc1511771} /* (31, 20, 17) {real, imag} */,
  {32'hc0dabad4, 32'h3e913760} /* (31, 20, 16) {real, imag} */,
  {32'hc1146eda, 32'hc17824b7} /* (31, 20, 15) {real, imag} */,
  {32'h40ceaeca, 32'h41147098} /* (31, 20, 14) {real, imag} */,
  {32'hc0958a32, 32'hc0d23f3a} /* (31, 20, 13) {real, imag} */,
  {32'hc18b05e8, 32'hc0de5688} /* (31, 20, 12) {real, imag} */,
  {32'h41a0b3a0, 32'hc05c677e} /* (31, 20, 11) {real, imag} */,
  {32'h41ec31d7, 32'h4085ee4c} /* (31, 20, 10) {real, imag} */,
  {32'h412d854e, 32'hc23afbce} /* (31, 20, 9) {real, imag} */,
  {32'hc2433869, 32'h41851ece} /* (31, 20, 8) {real, imag} */,
  {32'hc2698472, 32'h4270a582} /* (31, 20, 7) {real, imag} */,
  {32'hc180bab6, 32'hc016d16c} /* (31, 20, 6) {real, imag} */,
  {32'h41f6b204, 32'hc20a5836} /* (31, 20, 5) {real, imag} */,
  {32'h4028b070, 32'hc1bb93f0} /* (31, 20, 4) {real, imag} */,
  {32'h411cdab6, 32'h4255f2c5} /* (31, 20, 3) {real, imag} */,
  {32'hc0293c60, 32'hc145c6c3} /* (31, 20, 2) {real, imag} */,
  {32'h428eb778, 32'h42b68df2} /* (31, 20, 1) {real, imag} */,
  {32'h4241e4cc, 32'hc1870442} /* (31, 20, 0) {real, imag} */,
  {32'h42d60461, 32'h4252522a} /* (31, 19, 31) {real, imag} */,
  {32'hc12ea184, 32'h42550303} /* (31, 19, 30) {real, imag} */,
  {32'h41c0eedd, 32'hc21ef386} /* (31, 19, 29) {real, imag} */,
  {32'hc0dec014, 32'hc0132782} /* (31, 19, 28) {real, imag} */,
  {32'hc0593d80, 32'hc0e18578} /* (31, 19, 27) {real, imag} */,
  {32'hc26c52d4, 32'h422c5876} /* (31, 19, 26) {real, imag} */,
  {32'hc0c9928a, 32'hc20ac519} /* (31, 19, 25) {real, imag} */,
  {32'hc253a692, 32'hc20a8ef8} /* (31, 19, 24) {real, imag} */,
  {32'hc196b422, 32'hc00df850} /* (31, 19, 23) {real, imag} */,
  {32'hc145d67b, 32'hc0fad942} /* (31, 19, 22) {real, imag} */,
  {32'h40c4dd14, 32'hc09b92cc} /* (31, 19, 21) {real, imag} */,
  {32'h4098f4c6, 32'hc0fd4136} /* (31, 19, 20) {real, imag} */,
  {32'h41aef196, 32'h415c3bc0} /* (31, 19, 19) {real, imag} */,
  {32'h4190b7a2, 32'hc1859dce} /* (31, 19, 18) {real, imag} */,
  {32'hc14b414b, 32'h4156573c} /* (31, 19, 17) {real, imag} */,
  {32'h3eeac6c0, 32'hc15afd30} /* (31, 19, 16) {real, imag} */,
  {32'hc0694eec, 32'h40de5447} /* (31, 19, 15) {real, imag} */,
  {32'h4035b89c, 32'hbfbcf35c} /* (31, 19, 14) {real, imag} */,
  {32'hc11338a5, 32'h40ff35d8} /* (31, 19, 13) {real, imag} */,
  {32'hc18f2c7c, 32'hc1ce15c2} /* (31, 19, 12) {real, imag} */,
  {32'hc189d3ba, 32'hc07505e8} /* (31, 19, 11) {real, imag} */,
  {32'hc181a8d4, 32'h41a3fbee} /* (31, 19, 10) {real, imag} */,
  {32'hc0ed28a6, 32'hc24aa31b} /* (31, 19, 9) {real, imag} */,
  {32'h41311b70, 32'h3f967930} /* (31, 19, 8) {real, imag} */,
  {32'hc2024fe1, 32'h413d6834} /* (31, 19, 7) {real, imag} */,
  {32'h4279b68c, 32'h41bd6c24} /* (31, 19, 6) {real, imag} */,
  {32'hc1ddfae1, 32'hc28794a8} /* (31, 19, 5) {real, imag} */,
  {32'h422cca1a, 32'h414da4ee} /* (31, 19, 4) {real, imag} */,
  {32'h42111167, 32'hc0a708ac} /* (31, 19, 3) {real, imag} */,
  {32'h42b4bc7c, 32'h426cfcd7} /* (31, 19, 2) {real, imag} */,
  {32'hc2f2207f, 32'h424b6ed2} /* (31, 19, 1) {real, imag} */,
  {32'h422de2fc, 32'hc1c37504} /* (31, 19, 0) {real, imag} */,
  {32'hc2c7efb7, 32'h424420fa} /* (31, 18, 31) {real, imag} */,
  {32'h41b11154, 32'h4121aa1c} /* (31, 18, 30) {real, imag} */,
  {32'hc15d4d72, 32'hc2480060} /* (31, 18, 29) {real, imag} */,
  {32'hc215f331, 32'hc18eeaca} /* (31, 18, 28) {real, imag} */,
  {32'h42919716, 32'h4017a030} /* (31, 18, 27) {real, imag} */,
  {32'h423ad4d2, 32'hc241957e} /* (31, 18, 26) {real, imag} */,
  {32'hc22b065c, 32'hc17748c3} /* (31, 18, 25) {real, imag} */,
  {32'hc13eee4a, 32'hc089bd9a} /* (31, 18, 24) {real, imag} */,
  {32'h40047168, 32'hc11eeba1} /* (31, 18, 23) {real, imag} */,
  {32'hc1b21411, 32'hc0b1dafb} /* (31, 18, 22) {real, imag} */,
  {32'h4075da64, 32'hc16f9b2e} /* (31, 18, 21) {real, imag} */,
  {32'h4028de50, 32'hc0fe8608} /* (31, 18, 20) {real, imag} */,
  {32'hc12c196a, 32'hc0421708} /* (31, 18, 19) {real, imag} */,
  {32'h4189f15c, 32'h3fd02bd0} /* (31, 18, 18) {real, imag} */,
  {32'h411f791a, 32'h3efa0a10} /* (31, 18, 17) {real, imag} */,
  {32'h409253cc, 32'hbff2faa0} /* (31, 18, 16) {real, imag} */,
  {32'hbff8dd14, 32'hc0581d42} /* (31, 18, 15) {real, imag} */,
  {32'hc0c5e6be, 32'hc117935e} /* (31, 18, 14) {real, imag} */,
  {32'hc0f6bfec, 32'h410d1a0e} /* (31, 18, 13) {real, imag} */,
  {32'hbf31d620, 32'h41a909c6} /* (31, 18, 12) {real, imag} */,
  {32'h4114668f, 32'h418b524b} /* (31, 18, 11) {real, imag} */,
  {32'h401771b8, 32'hc06be576} /* (31, 18, 10) {real, imag} */,
  {32'hc1ba4c99, 32'hc181545c} /* (31, 18, 9) {real, imag} */,
  {32'h3f35d060, 32'h4139117d} /* (31, 18, 8) {real, imag} */,
  {32'hc187d04d, 32'hc016baec} /* (31, 18, 7) {real, imag} */,
  {32'hc0ed7900, 32'h419ec8eb} /* (31, 18, 6) {real, imag} */,
  {32'h41b26e32, 32'hc202c892} /* (31, 18, 5) {real, imag} */,
  {32'h4178b0cd, 32'hc209a0ef} /* (31, 18, 4) {real, imag} */,
  {32'h4191496b, 32'h40dd68fc} /* (31, 18, 3) {real, imag} */,
  {32'h3ff2d938, 32'h42019d40} /* (31, 18, 2) {real, imag} */,
  {32'hc2e2a071, 32'h420fd614} /* (31, 18, 1) {real, imag} */,
  {32'hc28496a8, 32'h429175da} /* (31, 18, 0) {real, imag} */,
  {32'h4277127e, 32'hc0c93f96} /* (31, 17, 31) {real, imag} */,
  {32'hc22ac71a, 32'hc1f4a56f} /* (31, 17, 30) {real, imag} */,
  {32'hc1a72d96, 32'h42513974} /* (31, 17, 29) {real, imag} */,
  {32'h41b4da1a, 32'hc131fb9c} /* (31, 17, 28) {real, imag} */,
  {32'hc160c559, 32'hc187aa36} /* (31, 17, 27) {real, imag} */,
  {32'h41705ed8, 32'hc12f18a6} /* (31, 17, 26) {real, imag} */,
  {32'h41249155, 32'hc190ee16} /* (31, 17, 25) {real, imag} */,
  {32'hc1d3c668, 32'h41a6f96a} /* (31, 17, 24) {real, imag} */,
  {32'hc19fd84e, 32'h4133413f} /* (31, 17, 23) {real, imag} */,
  {32'hbe4e1c40, 32'h4166a1c7} /* (31, 17, 22) {real, imag} */,
  {32'h3f17f270, 32'h404637c0} /* (31, 17, 21) {real, imag} */,
  {32'hbf4194c4, 32'h4098517f} /* (31, 17, 20) {real, imag} */,
  {32'hc151767d, 32'h4118cc7a} /* (31, 17, 19) {real, imag} */,
  {32'hc0204738, 32'hc062f9c0} /* (31, 17, 18) {real, imag} */,
  {32'hbf4dd690, 32'hc0d946c6} /* (31, 17, 17) {real, imag} */,
  {32'h413d7e54, 32'h40c15354} /* (31, 17, 16) {real, imag} */,
  {32'hc037f29c, 32'hbf8786e8} /* (31, 17, 15) {real, imag} */,
  {32'h3fca4330, 32'h40833d12} /* (31, 17, 14) {real, imag} */,
  {32'hc1103ca9, 32'h411e5e0a} /* (31, 17, 13) {real, imag} */,
  {32'h4095aa5c, 32'hc18e2483} /* (31, 17, 12) {real, imag} */,
  {32'h41e5df86, 32'hc1f12692} /* (31, 17, 11) {real, imag} */,
  {32'hc1a64b0a, 32'hc221c772} /* (31, 17, 10) {real, imag} */,
  {32'hbfd2a920, 32'hc0ba87d2} /* (31, 17, 9) {real, imag} */,
  {32'hc03f78c0, 32'hbfed7940} /* (31, 17, 8) {real, imag} */,
  {32'h3fccbed8, 32'hc2248f7b} /* (31, 17, 7) {real, imag} */,
  {32'h41ea49fc, 32'h40303fe0} /* (31, 17, 6) {real, imag} */,
  {32'h4208a31f, 32'h4235e92c} /* (31, 17, 5) {real, imag} */,
  {32'h417b565d, 32'h42405243} /* (31, 17, 4) {real, imag} */,
  {32'hc0d2cf34, 32'h420a933c} /* (31, 17, 3) {real, imag} */,
  {32'hc19b260b, 32'h4013c058} /* (31, 17, 2) {real, imag} */,
  {32'h40a44d70, 32'h41b6d400} /* (31, 17, 1) {real, imag} */,
  {32'h4176f21c, 32'h41db9551} /* (31, 17, 0) {real, imag} */,
  {32'h42098b9d, 32'hc149784c} /* (31, 16, 31) {real, imag} */,
  {32'hc1a3d771, 32'h418770ee} /* (31, 16, 30) {real, imag} */,
  {32'hc1d39fab, 32'hc120bec3} /* (31, 16, 29) {real, imag} */,
  {32'hc17a58c8, 32'hc19d1d48} /* (31, 16, 28) {real, imag} */,
  {32'hc1aa7b26, 32'h41219f2c} /* (31, 16, 27) {real, imag} */,
  {32'hc1c22903, 32'h4022d85c} /* (31, 16, 26) {real, imag} */,
  {32'hc0820f8e, 32'h415cd2b7} /* (31, 16, 25) {real, imag} */,
  {32'h41c1283c, 32'h41a2f2af} /* (31, 16, 24) {real, imag} */,
  {32'h41cd6721, 32'hbfd34a70} /* (31, 16, 23) {real, imag} */,
  {32'hbe825a38, 32'hc0d1df1e} /* (31, 16, 22) {real, imag} */,
  {32'h418bbbb5, 32'h412e4bb9} /* (31, 16, 21) {real, imag} */,
  {32'hc0b9e43b, 32'h414e9974} /* (31, 16, 20) {real, imag} */,
  {32'h41235176, 32'h40fdea08} /* (31, 16, 19) {real, imag} */,
  {32'h410c3e05, 32'hc01f78e0} /* (31, 16, 18) {real, imag} */,
  {32'hc184b0e6, 32'h416d9278} /* (31, 16, 17) {real, imag} */,
  {32'h40973015, 32'h405d47f2} /* (31, 16, 16) {real, imag} */,
  {32'hbf04c250, 32'h410960a8} /* (31, 16, 15) {real, imag} */,
  {32'hc0eea78e, 32'hc16f3338} /* (31, 16, 14) {real, imag} */,
  {32'hc14e43da, 32'h40e1be20} /* (31, 16, 13) {real, imag} */,
  {32'h41590dac, 32'hbeb331f0} /* (31, 16, 12) {real, imag} */,
  {32'hc169687d, 32'hc12d999b} /* (31, 16, 11) {real, imag} */,
  {32'h3d3c3e40, 32'h4190d0fa} /* (31, 16, 10) {real, imag} */,
  {32'hc1ae8e87, 32'hbfa570a0} /* (31, 16, 9) {real, imag} */,
  {32'hc069e614, 32'hc208feb1} /* (31, 16, 8) {real, imag} */,
  {32'hc1597bb1, 32'h41cc31ac} /* (31, 16, 7) {real, imag} */,
  {32'h4219db56, 32'hc1b547ba} /* (31, 16, 6) {real, imag} */,
  {32'h407b8358, 32'h40e9cee5} /* (31, 16, 5) {real, imag} */,
  {32'h410ecb32, 32'hc05b263c} /* (31, 16, 4) {real, imag} */,
  {32'h424061b0, 32'hc19a23d2} /* (31, 16, 3) {real, imag} */,
  {32'h41b91719, 32'hc299ace6} /* (31, 16, 2) {real, imag} */,
  {32'h41f6979e, 32'hc16c7048} /* (31, 16, 1) {real, imag} */,
  {32'hc0efd7e7, 32'h4122cc3e} /* (31, 16, 0) {real, imag} */,
  {32'hc257d086, 32'hc22109b9} /* (31, 15, 31) {real, imag} */,
  {32'h4182232a, 32'hc0fce43f} /* (31, 15, 30) {real, imag} */,
  {32'h41a4fc56, 32'hbf4532f8} /* (31, 15, 29) {real, imag} */,
  {32'hc2220670, 32'h41832d86} /* (31, 15, 28) {real, imag} */,
  {32'h41accb58, 32'hc1086622} /* (31, 15, 27) {real, imag} */,
  {32'h4279d792, 32'h41a54b50} /* (31, 15, 26) {real, imag} */,
  {32'hc138aa56, 32'hc1827fb8} /* (31, 15, 25) {real, imag} */,
  {32'h421f596e, 32'h3fd63e30} /* (31, 15, 24) {real, imag} */,
  {32'hc11f0d53, 32'hc20a1459} /* (31, 15, 23) {real, imag} */,
  {32'h41b91b34, 32'h415f459b} /* (31, 15, 22) {real, imag} */,
  {32'h40b32f48, 32'hc13c36ff} /* (31, 15, 21) {real, imag} */,
  {32'h3f84e1f4, 32'h411666d4} /* (31, 15, 20) {real, imag} */,
  {32'h40eed376, 32'hc141fb16} /* (31, 15, 19) {real, imag} */,
  {32'hc0a1b1ce, 32'hc0e75863} /* (31, 15, 18) {real, imag} */,
  {32'hbe734580, 32'h3f960ff8} /* (31, 15, 17) {real, imag} */,
  {32'hc02ce960, 32'hc0b7e2b4} /* (31, 15, 16) {real, imag} */,
  {32'hbfbd3690, 32'h400d141c} /* (31, 15, 15) {real, imag} */,
  {32'hc15efb1b, 32'h41055e4a} /* (31, 15, 14) {real, imag} */,
  {32'h3f892e78, 32'h411c9a8e} /* (31, 15, 13) {real, imag} */,
  {32'hc1340926, 32'h4057d0c4} /* (31, 15, 12) {real, imag} */,
  {32'h413bad0a, 32'hc17b1543} /* (31, 15, 11) {real, imag} */,
  {32'h40f924de, 32'hc064fd74} /* (31, 15, 10) {real, imag} */,
  {32'hc10976b9, 32'h41a6338a} /* (31, 15, 9) {real, imag} */,
  {32'hc1d680bf, 32'hc224106e} /* (31, 15, 8) {real, imag} */,
  {32'h4101a2c8, 32'hc1921534} /* (31, 15, 7) {real, imag} */,
  {32'h4008c140, 32'h4194b2ac} /* (31, 15, 6) {real, imag} */,
  {32'hc21b85d8, 32'hc0dc5198} /* (31, 15, 5) {real, imag} */,
  {32'h41901655, 32'hc1483510} /* (31, 15, 4) {real, imag} */,
  {32'hc1961288, 32'h411295f2} /* (31, 15, 3) {real, imag} */,
  {32'hc0eafcfa, 32'h411c0698} /* (31, 15, 2) {real, imag} */,
  {32'hc125ef08, 32'h416780f5} /* (31, 15, 1) {real, imag} */,
  {32'hc284ef19, 32'hc12aa3ba} /* (31, 15, 0) {real, imag} */,
  {32'h428be489, 32'hc2516ef3} /* (31, 14, 31) {real, imag} */,
  {32'hc1b6d492, 32'h41ecca9e} /* (31, 14, 30) {real, imag} */,
  {32'hc13cf097, 32'hc248bc6c} /* (31, 14, 29) {real, imag} */,
  {32'hc09546a0, 32'hc228358e} /* (31, 14, 28) {real, imag} */,
  {32'hc19cfd9f, 32'h4096e4c6} /* (31, 14, 27) {real, imag} */,
  {32'hc1e540e4, 32'hbfea04f8} /* (31, 14, 26) {real, imag} */,
  {32'h41983a2e, 32'h4081111c} /* (31, 14, 25) {real, imag} */,
  {32'h41f89aca, 32'h424a80cf} /* (31, 14, 24) {real, imag} */,
  {32'hc21650d9, 32'hc179350f} /* (31, 14, 23) {real, imag} */,
  {32'h3f7e3f30, 32'hc0895292} /* (31, 14, 22) {real, imag} */,
  {32'h402e05ee, 32'h41b96590} /* (31, 14, 21) {real, imag} */,
  {32'h3ce8a900, 32'hc1748f6d} /* (31, 14, 20) {real, imag} */,
  {32'h41719f6d, 32'h4059c710} /* (31, 14, 19) {real, imag} */,
  {32'h3f8aa420, 32'hbf35f7f8} /* (31, 14, 18) {real, imag} */,
  {32'hc1814ffa, 32'hbfa45c0c} /* (31, 14, 17) {real, imag} */,
  {32'h40e99c08, 32'hc1432fe6} /* (31, 14, 16) {real, imag} */,
  {32'hc02945f4, 32'h4104fdea} /* (31, 14, 15) {real, imag} */,
  {32'hc11ea98a, 32'hc17f9220} /* (31, 14, 14) {real, imag} */,
  {32'h41367d5d, 32'h409a9158} /* (31, 14, 13) {real, imag} */,
  {32'hc178110c, 32'h402e68cc} /* (31, 14, 12) {real, imag} */,
  {32'hc045394e, 32'hc1c94fb0} /* (31, 14, 11) {real, imag} */,
  {32'hc1a544be, 32'hbe33c2c0} /* (31, 14, 10) {real, imag} */,
  {32'h420e531b, 32'h3f4338d0} /* (31, 14, 9) {real, imag} */,
  {32'hc08ff580, 32'hc14e2dbc} /* (31, 14, 8) {real, imag} */,
  {32'hc1b82442, 32'h42037826} /* (31, 14, 7) {real, imag} */,
  {32'hc122da1f, 32'h41ef14b8} /* (31, 14, 6) {real, imag} */,
  {32'hc218cbb4, 32'hc16fadd7} /* (31, 14, 5) {real, imag} */,
  {32'hc23d840e, 32'h41763211} /* (31, 14, 4) {real, imag} */,
  {32'h421b9850, 32'hbf9bb590} /* (31, 14, 3) {real, imag} */,
  {32'hc15d3084, 32'h41cdb03a} /* (31, 14, 2) {real, imag} */,
  {32'h42c4b779, 32'h420fe765} /* (31, 14, 1) {real, imag} */,
  {32'h42747193, 32'hc1ffb631} /* (31, 14, 0) {real, imag} */,
  {32'hc26401bd, 32'hc2933a7f} /* (31, 13, 31) {real, imag} */,
  {32'hc1bb3779, 32'h41eab69e} /* (31, 13, 30) {real, imag} */,
  {32'hc198cdd4, 32'h41ac950a} /* (31, 13, 29) {real, imag} */,
  {32'hc0db5110, 32'hc14e75b5} /* (31, 13, 28) {real, imag} */,
  {32'h410d0ad5, 32'hc1992611} /* (31, 13, 27) {real, imag} */,
  {32'h4293169d, 32'hc1c7ba9a} /* (31, 13, 26) {real, imag} */,
  {32'h42120d7c, 32'h429831c2} /* (31, 13, 25) {real, imag} */,
  {32'h4143b79d, 32'h41f06712} /* (31, 13, 24) {real, imag} */,
  {32'hc178b59e, 32'hc1886482} /* (31, 13, 23) {real, imag} */,
  {32'h41af7133, 32'hc1f1999f} /* (31, 13, 22) {real, imag} */,
  {32'hc01f1304, 32'h4038cf0c} /* (31, 13, 21) {real, imag} */,
  {32'hc14081e7, 32'hc041b49f} /* (31, 13, 20) {real, imag} */,
  {32'hc0bc6e92, 32'hbea3e460} /* (31, 13, 19) {real, imag} */,
  {32'hc103dc36, 32'hc1686a0d} /* (31, 13, 18) {real, imag} */,
  {32'hc02fd34a, 32'hc1404c78} /* (31, 13, 17) {real, imag} */,
  {32'hc0639600, 32'hc0de10ca} /* (31, 13, 16) {real, imag} */,
  {32'h41343bd6, 32'hc0d1e390} /* (31, 13, 15) {real, imag} */,
  {32'hc123d96a, 32'h3eec4ba0} /* (31, 13, 14) {real, imag} */,
  {32'hc1c6f232, 32'h410cae89} /* (31, 13, 13) {real, imag} */,
  {32'h41472753, 32'h4129a27a} /* (31, 13, 12) {real, imag} */,
  {32'h40cb2416, 32'h41b15d90} /* (31, 13, 11) {real, imag} */,
  {32'hc1a1407f, 32'hc1b821db} /* (31, 13, 10) {real, imag} */,
  {32'h41d5119d, 32'hc209b39c} /* (31, 13, 9) {real, imag} */,
  {32'hc100a85d, 32'hc16915e8} /* (31, 13, 8) {real, imag} */,
  {32'h405b5458, 32'hc11c4c70} /* (31, 13, 7) {real, imag} */,
  {32'h414a7fde, 32'hc1700fa8} /* (31, 13, 6) {real, imag} */,
  {32'hc21b6b67, 32'h4275d11c} /* (31, 13, 5) {real, imag} */,
  {32'hc2805749, 32'hc104308f} /* (31, 13, 4) {real, imag} */,
  {32'h42011367, 32'hc21d3626} /* (31, 13, 3) {real, imag} */,
  {32'hc006cdb8, 32'h41c5d4b2} /* (31, 13, 2) {real, imag} */,
  {32'h428dd743, 32'h428ef763} /* (31, 13, 1) {real, imag} */,
  {32'hc2436a57, 32'hc1083867} /* (31, 13, 0) {real, imag} */,
  {32'h42ca29b6, 32'h4218dc6d} /* (31, 12, 31) {real, imag} */,
  {32'h40113c88, 32'h40d8a20e} /* (31, 12, 30) {real, imag} */,
  {32'hc1dd4110, 32'hc1244324} /* (31, 12, 29) {real, imag} */,
  {32'hc1acd018, 32'h42140de8} /* (31, 12, 28) {real, imag} */,
  {32'h41112b06, 32'h428b6376} /* (31, 12, 27) {real, imag} */,
  {32'h3fa2166c, 32'hc2a25958} /* (31, 12, 26) {real, imag} */,
  {32'h402c5fe0, 32'hbfeb2ab8} /* (31, 12, 25) {real, imag} */,
  {32'h41b58b15, 32'hc1be5198} /* (31, 12, 24) {real, imag} */,
  {32'h403afe10, 32'hc1a57411} /* (31, 12, 23) {real, imag} */,
  {32'h41d5f800, 32'hc1801114} /* (31, 12, 22) {real, imag} */,
  {32'h41fdc0a6, 32'h41fba5a2} /* (31, 12, 21) {real, imag} */,
  {32'h41a316fe, 32'h41df073c} /* (31, 12, 20) {real, imag} */,
  {32'hc131b6d4, 32'hc124ab6e} /* (31, 12, 19) {real, imag} */,
  {32'hc1bd529d, 32'h4103340f} /* (31, 12, 18) {real, imag} */,
  {32'h41051c90, 32'h4167fe7f} /* (31, 12, 17) {real, imag} */,
  {32'hbfb5f100, 32'h4196331a} /* (31, 12, 16) {real, imag} */,
  {32'h40390b00, 32'h4045e794} /* (31, 12, 15) {real, imag} */,
  {32'hc1113626, 32'hc0fb7c56} /* (31, 12, 14) {real, imag} */,
  {32'h40c10178, 32'hc0defbdf} /* (31, 12, 13) {real, imag} */,
  {32'hc0ee6734, 32'h4194cecc} /* (31, 12, 12) {real, imag} */,
  {32'h3f35b5f0, 32'hc18ca44e} /* (31, 12, 11) {real, imag} */,
  {32'hc1a36bb4, 32'hc21a8b10} /* (31, 12, 10) {real, imag} */,
  {32'hbf697240, 32'hc1b534f7} /* (31, 12, 9) {real, imag} */,
  {32'hc1a4ec99, 32'h42053b22} /* (31, 12, 8) {real, imag} */,
  {32'hc1605df8, 32'h41a0daf6} /* (31, 12, 7) {real, imag} */,
  {32'h410e817c, 32'h41ab12e2} /* (31, 12, 6) {real, imag} */,
  {32'h423fe2fa, 32'hbffc48a0} /* (31, 12, 5) {real, imag} */,
  {32'hc141be9f, 32'h425c059c} /* (31, 12, 4) {real, imag} */,
  {32'h42734650, 32'hc0dca54b} /* (31, 12, 3) {real, imag} */,
  {32'hc24085c8, 32'h4115f4fd} /* (31, 12, 2) {real, imag} */,
  {32'h42324109, 32'h4198b334} /* (31, 12, 1) {real, imag} */,
  {32'hc3030c94, 32'hc2b3813a} /* (31, 12, 0) {real, imag} */,
  {32'h430d4d46, 32'hc2abe816} /* (31, 11, 31) {real, imag} */,
  {32'hc2997f3a, 32'h424b5417} /* (31, 11, 30) {real, imag} */,
  {32'hc236db60, 32'hc1a0b2bf} /* (31, 11, 29) {real, imag} */,
  {32'hc03fa890, 32'hc09299ea} /* (31, 11, 28) {real, imag} */,
  {32'hc29d399c, 32'h4299e792} /* (31, 11, 27) {real, imag} */,
  {32'hc13fcf11, 32'h42e98ab8} /* (31, 11, 26) {real, imag} */,
  {32'h4198998b, 32'h3f557520} /* (31, 11, 25) {real, imag} */,
  {32'h41a3f5e6, 32'h428d63d2} /* (31, 11, 24) {real, imag} */,
  {32'hc1948c71, 32'h41bacfde} /* (31, 11, 23) {real, imag} */,
  {32'hc126bfcf, 32'h41c5841d} /* (31, 11, 22) {real, imag} */,
  {32'hc0948dba, 32'hbebf8320} /* (31, 11, 21) {real, imag} */,
  {32'hc04d8f18, 32'h41a038e3} /* (31, 11, 20) {real, imag} */,
  {32'h3fc70094, 32'hc0af245a} /* (31, 11, 19) {real, imag} */,
  {32'hc1e80dcc, 32'hc008884a} /* (31, 11, 18) {real, imag} */,
  {32'h411e5df3, 32'hc1208dff} /* (31, 11, 17) {real, imag} */,
  {32'h4118115c, 32'h419a32ae} /* (31, 11, 16) {real, imag} */,
  {32'hbf850998, 32'h3fcc8a58} /* (31, 11, 15) {real, imag} */,
  {32'h412277d8, 32'hbec13430} /* (31, 11, 14) {real, imag} */,
  {32'hc14989d2, 32'h4086ba02} /* (31, 11, 13) {real, imag} */,
  {32'h4232e298, 32'hc1d49cbb} /* (31, 11, 12) {real, imag} */,
  {32'h41355a2d, 32'h3f71b090} /* (31, 11, 11) {real, imag} */,
  {32'hc1f7cdf0, 32'hc0ebc124} /* (31, 11, 10) {real, imag} */,
  {32'h42325744, 32'h41655f67} /* (31, 11, 9) {real, imag} */,
  {32'hc0e89990, 32'hc0c06070} /* (31, 11, 8) {real, imag} */,
  {32'h4180aecd, 32'hc21b8f00} /* (31, 11, 7) {real, imag} */,
  {32'hc0eaab3e, 32'h4285965c} /* (31, 11, 6) {real, imag} */,
  {32'hc1c9ba3e, 32'h4176e724} /* (31, 11, 5) {real, imag} */,
  {32'h42abc068, 32'h41265388} /* (31, 11, 4) {real, imag} */,
  {32'h4166200e, 32'h421f1c78} /* (31, 11, 3) {real, imag} */,
  {32'hc2e8f8aa, 32'h41964e22} /* (31, 11, 2) {real, imag} */,
  {32'h4323de24, 32'hc22fce6f} /* (31, 11, 1) {real, imag} */,
  {32'h42c9d5c6, 32'hc2b62806} /* (31, 11, 0) {real, imag} */,
  {32'hc2c259d2, 32'h40a70a08} /* (31, 10, 31) {real, imag} */,
  {32'h42f41fe5, 32'hc2134612} /* (31, 10, 30) {real, imag} */,
  {32'hc0a9ac52, 32'h42202885} /* (31, 10, 29) {real, imag} */,
  {32'hc09d5d6c, 32'h41fb0986} /* (31, 10, 28) {real, imag} */,
  {32'hc08d4008, 32'hc07c8ba0} /* (31, 10, 27) {real, imag} */,
  {32'h40672078, 32'hbf8f9f18} /* (31, 10, 26) {real, imag} */,
  {32'hc1d23304, 32'hc281202c} /* (31, 10, 25) {real, imag} */,
  {32'hc24bba98, 32'hc1bfc872} /* (31, 10, 24) {real, imag} */,
  {32'h414dfbf5, 32'hc1233f5c} /* (31, 10, 23) {real, imag} */,
  {32'hc1d02841, 32'h41135367} /* (31, 10, 22) {real, imag} */,
  {32'hc1f4f380, 32'hc1346e72} /* (31, 10, 21) {real, imag} */,
  {32'hc0d3590e, 32'h41fdd004} /* (31, 10, 20) {real, imag} */,
  {32'h40d55749, 32'hc18b1b98} /* (31, 10, 19) {real, imag} */,
  {32'h4181a6dd, 32'hc1aa68f6} /* (31, 10, 18) {real, imag} */,
  {32'h403f4d22, 32'h41144c4c} /* (31, 10, 17) {real, imag} */,
  {32'h411d6070, 32'hc0a12488} /* (31, 10, 16) {real, imag} */,
  {32'h410c61c0, 32'h405c9af0} /* (31, 10, 15) {real, imag} */,
  {32'h41838c15, 32'hc042c7a0} /* (31, 10, 14) {real, imag} */,
  {32'h41856903, 32'hc0b9be58} /* (31, 10, 13) {real, imag} */,
  {32'h417f8d1d, 32'h40586bbc} /* (31, 10, 12) {real, imag} */,
  {32'hc0ec2190, 32'h40d0ae84} /* (31, 10, 11) {real, imag} */,
  {32'h4127d2b2, 32'hc1c5cf92} /* (31, 10, 10) {real, imag} */,
  {32'h410c06f5, 32'h428c37f0} /* (31, 10, 9) {real, imag} */,
  {32'h4134666e, 32'hc25eddc1} /* (31, 10, 8) {real, imag} */,
  {32'h41d50370, 32'hc10024f4} /* (31, 10, 7) {real, imag} */,
  {32'hbffe5970, 32'hc1b84388} /* (31, 10, 6) {real, imag} */,
  {32'h422dc173, 32'h42ab2c3d} /* (31, 10, 5) {real, imag} */,
  {32'hc221dd6a, 32'h427e94ef} /* (31, 10, 4) {real, imag} */,
  {32'h41d9ee4a, 32'h41c6b9b6} /* (31, 10, 3) {real, imag} */,
  {32'h4122f028, 32'h42accc35} /* (31, 10, 2) {real, imag} */,
  {32'hc29a212a, 32'h42a3bd0a} /* (31, 10, 1) {real, imag} */,
  {32'hc2b2e1b0, 32'hc2a043ea} /* (31, 10, 0) {real, imag} */,
  {32'hc2a0c426, 32'hc2ab26da} /* (31, 9, 31) {real, imag} */,
  {32'h4376e0f2, 32'h42478e0c} /* (31, 9, 30) {real, imag} */,
  {32'hc3192ebc, 32'hc1672720} /* (31, 9, 29) {real, imag} */,
  {32'h4268751a, 32'h429abc69} /* (31, 9, 28) {real, imag} */,
  {32'h3e070100, 32'hc0aef894} /* (31, 9, 27) {real, imag} */,
  {32'h42a9e53c, 32'h42bd0633} /* (31, 9, 26) {real, imag} */,
  {32'hc03452c8, 32'hc1f7c38e} /* (31, 9, 25) {real, imag} */,
  {32'hc19b4f68, 32'hc2bf81fd} /* (31, 9, 24) {real, imag} */,
  {32'h410c5f44, 32'hc28447de} /* (31, 9, 23) {real, imag} */,
  {32'h418f8000, 32'h41c2f098} /* (31, 9, 22) {real, imag} */,
  {32'h4224f42e, 32'hc1724685} /* (31, 9, 21) {real, imag} */,
  {32'hc211c1f1, 32'hc1889200} /* (31, 9, 20) {real, imag} */,
  {32'hc2266924, 32'h40240468} /* (31, 9, 19) {real, imag} */,
  {32'h41cf82f3, 32'h41ad1621} /* (31, 9, 18) {real, imag} */,
  {32'hc1b63bba, 32'hc20382c4} /* (31, 9, 17) {real, imag} */,
  {32'h419e53ee, 32'h3e0e5880} /* (31, 9, 16) {real, imag} */,
  {32'hc20f37a3, 32'hc1b172c7} /* (31, 9, 15) {real, imag} */,
  {32'hc19cac8b, 32'h412eac5a} /* (31, 9, 14) {real, imag} */,
  {32'h418fd55f, 32'hbfa24870} /* (31, 9, 13) {real, imag} */,
  {32'h4207d7f9, 32'h3ee0f600} /* (31, 9, 12) {real, imag} */,
  {32'h417947c2, 32'hc14bcae7} /* (31, 9, 11) {real, imag} */,
  {32'h423eea94, 32'hbfc36a40} /* (31, 9, 10) {real, imag} */,
  {32'hc2c8a6cc, 32'hc22c60b6} /* (31, 9, 9) {real, imag} */,
  {32'h4288e82e, 32'hc2a20eb7} /* (31, 9, 8) {real, imag} */,
  {32'hc1cf393d, 32'hc26a14a7} /* (31, 9, 7) {real, imag} */,
  {32'hc1abecb7, 32'h41ea45b0} /* (31, 9, 6) {real, imag} */,
  {32'h42f9e722, 32'hc2271212} /* (31, 9, 5) {real, imag} */,
  {32'h42a7f8fb, 32'hc285a7ed} /* (31, 9, 4) {real, imag} */,
  {32'hc33ee058, 32'h4302d1be} /* (31, 9, 3) {real, imag} */,
  {32'h42e8eb63, 32'hc2dbc34a} /* (31, 9, 2) {real, imag} */,
  {32'hc31104d1, 32'h4245e2fc} /* (31, 9, 1) {real, imag} */,
  {32'hc29f7c78, 32'hc1756dc2} /* (31, 9, 0) {real, imag} */,
  {32'h4351bf0d, 32'hc3d6be97} /* (31, 8, 31) {real, imag} */,
  {32'hc1b675db, 32'h43267cfa} /* (31, 8, 30) {real, imag} */,
  {32'hc234e7b9, 32'hc15a2b83} /* (31, 8, 29) {real, imag} */,
  {32'hc2cbd00f, 32'h41258e8c} /* (31, 8, 28) {real, imag} */,
  {32'h414e5ebd, 32'h43867352} /* (31, 8, 27) {real, imag} */,
  {32'hbf013980, 32'h424930a8} /* (31, 8, 26) {real, imag} */,
  {32'hc25f742c, 32'hbf60d780} /* (31, 8, 25) {real, imag} */,
  {32'h4188680b, 32'h42c7f908} /* (31, 8, 24) {real, imag} */,
  {32'h426daa82, 32'hc1f8d261} /* (31, 8, 23) {real, imag} */,
  {32'hc2018337, 32'hc28348c5} /* (31, 8, 22) {real, imag} */,
  {32'hc149df06, 32'hc157c460} /* (31, 8, 21) {real, imag} */,
  {32'hc0c4af90, 32'hc21946a0} /* (31, 8, 20) {real, imag} */,
  {32'h3fd6ffe8, 32'h4133180f} /* (31, 8, 19) {real, imag} */,
  {32'h4061ead8, 32'h41bea27c} /* (31, 8, 18) {real, imag} */,
  {32'h4204c90e, 32'h415f0748} /* (31, 8, 17) {real, imag} */,
  {32'hc222c1c8, 32'hc168e528} /* (31, 8, 16) {real, imag} */,
  {32'h4184ae63, 32'h40c854f0} /* (31, 8, 15) {real, imag} */,
  {32'hc1810001, 32'h40f935f0} /* (31, 8, 14) {real, imag} */,
  {32'h4200cf0b, 32'hc1d7af76} /* (31, 8, 13) {real, imag} */,
  {32'hc1f49af8, 32'h41a96622} /* (31, 8, 12) {real, imag} */,
  {32'hc21999f8, 32'hc1dec7e0} /* (31, 8, 11) {real, imag} */,
  {32'h4245b411, 32'h411ff71a} /* (31, 8, 10) {real, imag} */,
  {32'hc27298d2, 32'hc07e6f78} /* (31, 8, 9) {real, imag} */,
  {32'hc270fbc2, 32'h428973c2} /* (31, 8, 8) {real, imag} */,
  {32'hc279b0c0, 32'hc2d77ba9} /* (31, 8, 7) {real, imag} */,
  {32'hc2ad6cd3, 32'hc171be52} /* (31, 8, 6) {real, imag} */,
  {32'hc004270c, 32'h429e8b02} /* (31, 8, 5) {real, imag} */,
  {32'h42dd95d9, 32'hc288f362} /* (31, 8, 4) {real, imag} */,
  {32'h41006e6c, 32'h41c3b9d8} /* (31, 8, 3) {real, imag} */,
  {32'hc13cf956, 32'h43a35b55} /* (31, 8, 2) {real, imag} */,
  {32'h42f439ae, 32'hc38bafb7} /* (31, 8, 1) {real, imag} */,
  {32'h42581380, 32'hc2bd6e45} /* (31, 8, 0) {real, imag} */,
  {32'hc305a924, 32'h437a1d6d} /* (31, 7, 31) {real, imag} */,
  {32'hc258d57d, 32'h42af4ae6} /* (31, 7, 30) {real, imag} */,
  {32'hc271b020, 32'hc2ab7657} /* (31, 7, 29) {real, imag} */,
  {32'hc2a39e7e, 32'hc2cde196} /* (31, 7, 28) {real, imag} */,
  {32'h41192e74, 32'h41b50ef0} /* (31, 7, 27) {real, imag} */,
  {32'h42a26a91, 32'h42365b0e} /* (31, 7, 26) {real, imag} */,
  {32'h4279ad66, 32'h42c38d46} /* (31, 7, 25) {real, imag} */,
  {32'h42884408, 32'hc249310f} /* (31, 7, 24) {real, imag} */,
  {32'h4202508c, 32'hc301773e} /* (31, 7, 23) {real, imag} */,
  {32'hc283a886, 32'h401db4d0} /* (31, 7, 22) {real, imag} */,
  {32'hc244f6ba, 32'h42199404} /* (31, 7, 21) {real, imag} */,
  {32'h40791388, 32'h418e11b0} /* (31, 7, 20) {real, imag} */,
  {32'hc205f04a, 32'h418b5588} /* (31, 7, 19) {real, imag} */,
  {32'h40ea08f0, 32'h41c3fe17} /* (31, 7, 18) {real, imag} */,
  {32'hc1dd60c5, 32'h41779052} /* (31, 7, 17) {real, imag} */,
  {32'hc1d26e54, 32'hc219d9da} /* (31, 7, 16) {real, imag} */,
  {32'h420372ce, 32'hc1c615df} /* (31, 7, 15) {real, imag} */,
  {32'h41a3d794, 32'hc216facc} /* (31, 7, 14) {real, imag} */,
  {32'hc186ad71, 32'h4099cf4e} /* (31, 7, 13) {real, imag} */,
  {32'h41fbb48b, 32'hc25c8d32} /* (31, 7, 12) {real, imag} */,
  {32'hc1bdbded, 32'h42805545} /* (31, 7, 11) {real, imag} */,
  {32'h40cd6864, 32'h42ca2050} /* (31, 7, 10) {real, imag} */,
  {32'h41c918d9, 32'h42193770} /* (31, 7, 9) {real, imag} */,
  {32'h4211c8a7, 32'h4207c3cb} /* (31, 7, 8) {real, imag} */,
  {32'hc15e9dc8, 32'h41f10092} /* (31, 7, 7) {real, imag} */,
  {32'h4220ac2e, 32'h42b65131} /* (31, 7, 6) {real, imag} */,
  {32'h424e39a6, 32'h42f25e30} /* (31, 7, 5) {real, imag} */,
  {32'hc30a1869, 32'hc3216f03} /* (31, 7, 4) {real, imag} */,
  {32'h420a4be4, 32'hc2d96061} /* (31, 7, 3) {real, imag} */,
  {32'h42ec2e76, 32'hc23cb59c} /* (31, 7, 2) {real, imag} */,
  {32'hc2d1b5e7, 32'hc30dfefb} /* (31, 7, 1) {real, imag} */,
  {32'h404b4720, 32'hc191c2c4} /* (31, 7, 0) {real, imag} */,
  {32'hc26c9f9a, 32'h433a6544} /* (31, 6, 31) {real, imag} */,
  {32'h417db064, 32'h430b50dc} /* (31, 6, 30) {real, imag} */,
  {32'h42f6a4f0, 32'h427c3286} /* (31, 6, 29) {real, imag} */,
  {32'h41b1a7cd, 32'hc298fcf5} /* (31, 6, 28) {real, imag} */,
  {32'hc1b7dbc4, 32'h428fe52c} /* (31, 6, 27) {real, imag} */,
  {32'h3f189d80, 32'h42bd28cb} /* (31, 6, 26) {real, imag} */,
  {32'h42b68656, 32'h42b64d0c} /* (31, 6, 25) {real, imag} */,
  {32'h420b55e6, 32'h42539e9a} /* (31, 6, 24) {real, imag} */,
  {32'hc2444cd8, 32'hc1d1a445} /* (31, 6, 23) {real, imag} */,
  {32'hc1873e14, 32'h421008d1} /* (31, 6, 22) {real, imag} */,
  {32'hc19959f2, 32'hc162bbc4} /* (31, 6, 21) {real, imag} */,
  {32'hc0c84a90, 32'hc1b45f6c} /* (31, 6, 20) {real, imag} */,
  {32'hc2a28fbc, 32'hc1b3100a} /* (31, 6, 19) {real, imag} */,
  {32'h419987ae, 32'h4206dec2} /* (31, 6, 18) {real, imag} */,
  {32'hc103930a, 32'hc1a094da} /* (31, 6, 17) {real, imag} */,
  {32'h41f8f9e1, 32'hc2709563} /* (31, 6, 16) {real, imag} */,
  {32'hc090536c, 32'hc0a2d018} /* (31, 6, 15) {real, imag} */,
  {32'hc197cf66, 32'h4202393a} /* (31, 6, 14) {real, imag} */,
  {32'hc1cbbdc2, 32'h419a98fa} /* (31, 6, 13) {real, imag} */,
  {32'hc2611ded, 32'hc0ca9ace} /* (31, 6, 12) {real, imag} */,
  {32'h41827b46, 32'h422ef4f5} /* (31, 6, 11) {real, imag} */,
  {32'h42d28e27, 32'h4215409d} /* (31, 6, 10) {real, imag} */,
  {32'h420a3330, 32'hc254ef42} /* (31, 6, 9) {real, imag} */,
  {32'h427f8872, 32'h424fa0d0} /* (31, 6, 8) {real, imag} */,
  {32'h417beff4, 32'h42d6dac6} /* (31, 6, 7) {real, imag} */,
  {32'hc3273dcc, 32'h4290a679} /* (31, 6, 6) {real, imag} */,
  {32'h42a02943, 32'h42c079d0} /* (31, 6, 5) {real, imag} */,
  {32'h4298287b, 32'hc2c5b1f5} /* (31, 6, 4) {real, imag} */,
  {32'hc315cf1e, 32'hc2f6145d} /* (31, 6, 3) {real, imag} */,
  {32'hc28683fe, 32'hc350a5a6} /* (31, 6, 2) {real, imag} */,
  {32'hc2b87dbb, 32'h41aa8d80} /* (31, 6, 1) {real, imag} */,
  {32'h42356e10, 32'hc2520e2b} /* (31, 6, 0) {real, imag} */,
  {32'hc2edad1a, 32'hc417e4f2} /* (31, 5, 31) {real, imag} */,
  {32'h42220ec4, 32'h4310471c} /* (31, 5, 30) {real, imag} */,
  {32'hc2c9ab72, 32'hc3533d66} /* (31, 5, 29) {real, imag} */,
  {32'h420e68d3, 32'hc2bc327c} /* (31, 5, 28) {real, imag} */,
  {32'hc21ce07a, 32'h4286928d} /* (31, 5, 27) {real, imag} */,
  {32'hc119c9b6, 32'hc2a7f44a} /* (31, 5, 26) {real, imag} */,
  {32'hc280c89a, 32'h41f0b104} /* (31, 5, 25) {real, imag} */,
  {32'h42e38956, 32'h42e62af0} /* (31, 5, 24) {real, imag} */,
  {32'hc1aed074, 32'hc21908a2} /* (31, 5, 23) {real, imag} */,
  {32'h415122d4, 32'h4105a8a0} /* (31, 5, 22) {real, imag} */,
  {32'hc1338068, 32'h42425166} /* (31, 5, 21) {real, imag} */,
  {32'h4224acd9, 32'hc29caf10} /* (31, 5, 20) {real, imag} */,
  {32'h411899db, 32'hc1335440} /* (31, 5, 19) {real, imag} */,
  {32'h414f8038, 32'hc1c396f3} /* (31, 5, 18) {real, imag} */,
  {32'hc2264529, 32'hbde0b000} /* (31, 5, 17) {real, imag} */,
  {32'hbd77e000, 32'h4157c280} /* (31, 5, 16) {real, imag} */,
  {32'h3f773ac0, 32'h40d45a40} /* (31, 5, 15) {real, imag} */,
  {32'hc1edcbec, 32'hc1eacc3d} /* (31, 5, 14) {real, imag} */,
  {32'h411844c5, 32'h42157db8} /* (31, 5, 13) {real, imag} */,
  {32'hc22aee67, 32'h428d0122} /* (31, 5, 12) {real, imag} */,
  {32'hc2cd146f, 32'h41e60dad} /* (31, 5, 11) {real, imag} */,
  {32'hc286184e, 32'hc15de598} /* (31, 5, 10) {real, imag} */,
  {32'hc23eb896, 32'h42af7f2b} /* (31, 5, 9) {real, imag} */,
  {32'hc27355cb, 32'hc237f4f7} /* (31, 5, 8) {real, imag} */,
  {32'h41ddec30, 32'hc326c512} /* (31, 5, 7) {real, imag} */,
  {32'hc227042c, 32'hbd302800} /* (31, 5, 6) {real, imag} */,
  {32'hc286b98b, 32'h4231356a} /* (31, 5, 5) {real, imag} */,
  {32'h42b183da, 32'hc16ac69c} /* (31, 5, 4) {real, imag} */,
  {32'hc2c8c026, 32'hc2c37758} /* (31, 5, 3) {real, imag} */,
  {32'hc36da8df, 32'h434d9682} /* (31, 5, 2) {real, imag} */,
  {32'h43c530a8, 32'hc3806910} /* (31, 5, 1) {real, imag} */,
  {32'h438ec484, 32'hc39e1a86} /* (31, 5, 0) {real, imag} */,
  {32'hc3d15336, 32'h437d8492} /* (31, 4, 31) {real, imag} */,
  {32'h438a39aa, 32'hc38c2e9e} /* (31, 4, 30) {real, imag} */,
  {32'hc1889cd4, 32'h42dcf5dc} /* (31, 4, 29) {real, imag} */,
  {32'hc1b93db8, 32'h4334def1} /* (31, 4, 28) {real, imag} */,
  {32'hc290a30c, 32'hc2806744} /* (31, 4, 27) {real, imag} */,
  {32'h410a0094, 32'hc2d7b0b4} /* (31, 4, 26) {real, imag} */,
  {32'hc1a58870, 32'hc278cb67} /* (31, 4, 25) {real, imag} */,
  {32'hc1376340, 32'hc2ac4057} /* (31, 4, 24) {real, imag} */,
  {32'hc2244a6c, 32'h42b0b00f} /* (31, 4, 23) {real, imag} */,
  {32'h42b23f76, 32'hc189654f} /* (31, 4, 22) {real, imag} */,
  {32'h42948f26, 32'h421c2af0} /* (31, 4, 21) {real, imag} */,
  {32'hc1c87f26, 32'h40becc7c} /* (31, 4, 20) {real, imag} */,
  {32'hc0b3b008, 32'h3fdbf580} /* (31, 4, 19) {real, imag} */,
  {32'h418d1c6c, 32'hc1effc70} /* (31, 4, 18) {real, imag} */,
  {32'h41abef1a, 32'hc031e3e0} /* (31, 4, 17) {real, imag} */,
  {32'hbf94b4c0, 32'h4101a990} /* (31, 4, 16) {real, imag} */,
  {32'hc23f732d, 32'hc04cc5a0} /* (31, 4, 15) {real, imag} */,
  {32'h42479c3a, 32'h428e29fc} /* (31, 4, 14) {real, imag} */,
  {32'h420df3d3, 32'hc1a9c358} /* (31, 4, 13) {real, imag} */,
  {32'hc29ad8fa, 32'hc221abac} /* (31, 4, 12) {real, imag} */,
  {32'h42ff44fe, 32'h42acdc58} /* (31, 4, 11) {real, imag} */,
  {32'hc1ac448a, 32'hc16daace} /* (31, 4, 10) {real, imag} */,
  {32'hbf980070, 32'h41c3d660} /* (31, 4, 9) {real, imag} */,
  {32'h429b8570, 32'h40fcd1a0} /* (31, 4, 8) {real, imag} */,
  {32'h428dcc60, 32'h42c59324} /* (31, 4, 7) {real, imag} */,
  {32'h42d70632, 32'h42a180fa} /* (31, 4, 6) {real, imag} */,
  {32'h4376bdd8, 32'hc29fc6ec} /* (31, 4, 5) {real, imag} */,
  {32'hc37eb99f, 32'hc2ef367e} /* (31, 4, 4) {real, imag} */,
  {32'hc301b1c4, 32'h3f38d000} /* (31, 4, 3) {real, imag} */,
  {32'h43508add, 32'hc3d3efe8} /* (31, 4, 2) {real, imag} */,
  {32'hc38635c2, 32'h4426166c} /* (31, 4, 1) {real, imag} */,
  {32'h4329cbe2, 32'h439ae198} /* (31, 4, 0) {real, imag} */,
  {32'hc3705718, 32'hc37e304e} /* (31, 3, 31) {real, imag} */,
  {32'h43ee3068, 32'h40599970} /* (31, 3, 30) {real, imag} */,
  {32'h429b1453, 32'hc20e843c} /* (31, 3, 29) {real, imag} */,
  {32'hc307109f, 32'h43752fe8} /* (31, 3, 28) {real, imag} */,
  {32'hc1a1f8c0, 32'hc35f28d8} /* (31, 3, 27) {real, imag} */,
  {32'hc17dc2fc, 32'hc2609c94} /* (31, 3, 26) {real, imag} */,
  {32'hc23a3d3e, 32'hc1fe7e48} /* (31, 3, 25) {real, imag} */,
  {32'h41d9430b, 32'h42e78a1e} /* (31, 3, 24) {real, imag} */,
  {32'h42370d09, 32'hc1ce1170} /* (31, 3, 23) {real, imag} */,
  {32'h429fe398, 32'h429ba928} /* (31, 3, 22) {real, imag} */,
  {32'hc2019c1d, 32'h40e47f00} /* (31, 3, 21) {real, imag} */,
  {32'hc2565714, 32'h403581a0} /* (31, 3, 20) {real, imag} */,
  {32'hc17adffe, 32'h425015dc} /* (31, 3, 19) {real, imag} */,
  {32'h41a0d6e8, 32'hc24e14a2} /* (31, 3, 18) {real, imag} */,
  {32'hc029237c, 32'hc0d10fc0} /* (31, 3, 17) {real, imag} */,
  {32'hc177bcea, 32'hc2781438} /* (31, 3, 16) {real, imag} */,
  {32'hc0f1af42, 32'hc1c178c0} /* (31, 3, 15) {real, imag} */,
  {32'h423fc7ec, 32'h43007baa} /* (31, 3, 14) {real, imag} */,
  {32'hc105f5fe, 32'hc128dc70} /* (31, 3, 13) {real, imag} */,
  {32'h41c53394, 32'h40cff450} /* (31, 3, 12) {real, imag} */,
  {32'hc196b940, 32'hc23dc13a} /* (31, 3, 11) {real, imag} */,
  {32'hc1cc66b6, 32'hc27662ec} /* (31, 3, 10) {real, imag} */,
  {32'h42abe8a6, 32'h42d2517a} /* (31, 3, 9) {real, imag} */,
  {32'hc26f8b98, 32'h42184463} /* (31, 3, 8) {real, imag} */,
  {32'h42ab5c71, 32'hc2897640} /* (31, 3, 7) {real, imag} */,
  {32'hc29afc8a, 32'hc144b580} /* (31, 3, 6) {real, imag} */,
  {32'hc3018fcd, 32'h421f6c28} /* (31, 3, 5) {real, imag} */,
  {32'hc28bc006, 32'hc32874b8} /* (31, 3, 4) {real, imag} */,
  {32'hc2960c13, 32'hc32bfd65} /* (31, 3, 3) {real, imag} */,
  {32'h434c77df, 32'h406b6af0} /* (31, 3, 2) {real, imag} */,
  {32'hc389bc6c, 32'h4405a2e2} /* (31, 3, 1) {real, imag} */,
  {32'h4210eb4c, 32'hc2cb9d44} /* (31, 3, 0) {real, imag} */,
  {32'hc30413af, 32'hc4efbcfe} /* (31, 2, 31) {real, imag} */,
  {32'h44094b88, 32'h4493f951} /* (31, 2, 30) {real, imag} */,
  {32'hc36e31a8, 32'hc2af3322} /* (31, 2, 29) {real, imag} */,
  {32'hc38f5bca, 32'hc214d0ac} /* (31, 2, 28) {real, imag} */,
  {32'h43421415, 32'h43a61052} /* (31, 2, 27) {real, imag} */,
  {32'h42a30198, 32'h42ba99ae} /* (31, 2, 26) {real, imag} */,
  {32'h42079018, 32'h41fca166} /* (31, 2, 25) {real, imag} */,
  {32'h4338413d, 32'h435cd90d} /* (31, 2, 24) {real, imag} */,
  {32'h413723f4, 32'hc303d722} /* (31, 2, 23) {real, imag} */,
  {32'hc0a8fc08, 32'hc1d53f6e} /* (31, 2, 22) {real, imag} */,
  {32'h41657cd4, 32'hc207e688} /* (31, 2, 21) {real, imag} */,
  {32'h412c6a84, 32'h4268c50e} /* (31, 2, 20) {real, imag} */,
  {32'h426850f8, 32'hc1f70c96} /* (31, 2, 19) {real, imag} */,
  {32'h4255873b, 32'hc188cc8c} /* (31, 2, 18) {real, imag} */,
  {32'h40aa0c68, 32'h41e5e2b0} /* (31, 2, 17) {real, imag} */,
  {32'h41b892d8, 32'h41ca4ef0} /* (31, 2, 16) {real, imag} */,
  {32'h41872d36, 32'hc1d0c4f0} /* (31, 2, 15) {real, imag} */,
  {32'hc0a274d8, 32'hc12c7268} /* (31, 2, 14) {real, imag} */,
  {32'hc0e7e6e0, 32'hc26a6ec9} /* (31, 2, 13) {real, imag} */,
  {32'h408d67e8, 32'h41bfac0c} /* (31, 2, 12) {real, imag} */,
  {32'hc2f1186c, 32'h4284745c} /* (31, 2, 11) {real, imag} */,
  {32'h41d3e0f2, 32'hc24e64f7} /* (31, 2, 10) {real, imag} */,
  {32'hc19a9206, 32'hc186b240} /* (31, 2, 9) {real, imag} */,
  {32'hc328047d, 32'h437c12e7} /* (31, 2, 8) {real, imag} */,
  {32'h42f8d7ac, 32'hc2ad9a66} /* (31, 2, 7) {real, imag} */,
  {32'hc249f078, 32'hc27a8add} /* (31, 2, 6) {real, imag} */,
  {32'hc359c9a3, 32'h43c7f1c0} /* (31, 2, 5) {real, imag} */,
  {32'h428d391a, 32'hc38655b2} /* (31, 2, 4) {real, imag} */,
  {32'hc36e81e8, 32'hc2808aa8} /* (31, 2, 3) {real, imag} */,
  {32'h4387c93c, 32'h445c1cbe} /* (31, 2, 2) {real, imag} */,
  {32'hc3b431c0, 32'hc4702c3c} /* (31, 2, 1) {real, imag} */,
  {32'h420c97bf, 32'hc470c0fc} /* (31, 2, 0) {real, imag} */,
  {32'h4400b8d5, 32'h44b1e7e4} /* (31, 1, 31) {real, imag} */,
  {32'hc2443648, 32'hc410fd6c} /* (31, 1, 30) {real, imag} */,
  {32'h422ca10b, 32'hc2856d84} /* (31, 1, 29) {real, imag} */,
  {32'hc382ae50, 32'h43e83337} /* (31, 1, 28) {real, imag} */,
  {32'hc2876293, 32'hc400fa9b} /* (31, 1, 27) {real, imag} */,
  {32'hc35f0ca4, 32'h423f58fc} /* (31, 1, 26) {real, imag} */,
  {32'h4185dfa4, 32'hc2c8961a} /* (31, 1, 25) {real, imag} */,
  {32'h40341800, 32'hc2f7fdda} /* (31, 1, 24) {real, imag} */,
  {32'hc1c4b314, 32'hc2b93c22} /* (31, 1, 23) {real, imag} */,
  {32'hc3320274, 32'hc03c0a80} /* (31, 1, 22) {real, imag} */,
  {32'hc2b83ee4, 32'hc31b97a4} /* (31, 1, 21) {real, imag} */,
  {32'h4291d4af, 32'h4264fe8c} /* (31, 1, 20) {real, imag} */,
  {32'hc1dfe9fe, 32'hc23eafaf} /* (31, 1, 19) {real, imag} */,
  {32'hc2fbf214, 32'hc28b41ac} /* (31, 1, 18) {real, imag} */,
  {32'hc093d580, 32'hc1165ab0} /* (31, 1, 17) {real, imag} */,
  {32'hc2282a3b, 32'h41106080} /* (31, 1, 16) {real, imag} */,
  {32'hc1c66fc0, 32'h41b2c118} /* (31, 1, 15) {real, imag} */,
  {32'h42620168, 32'hc2455168} /* (31, 1, 14) {real, imag} */,
  {32'h41ad7a16, 32'h41680adc} /* (31, 1, 13) {real, imag} */,
  {32'h42bd88cd, 32'h42393048} /* (31, 1, 12) {real, imag} */,
  {32'h432ba468, 32'hc2c51618} /* (31, 1, 11) {real, imag} */,
  {32'h41f0fa80, 32'hbf5b2a00} /* (31, 1, 10) {real, imag} */,
  {32'hc2db9d9d, 32'hc25e3d44} /* (31, 1, 9) {real, imag} */,
  {32'h4383edb8, 32'hc33e16fb} /* (31, 1, 8) {real, imag} */,
  {32'hc33da750, 32'h435765a7} /* (31, 1, 7) {real, imag} */,
  {32'h4273d8a0, 32'hc2916576} /* (31, 1, 6) {real, imag} */,
  {32'h42cb8555, 32'hc3d10912} /* (31, 1, 5) {real, imag} */,
  {32'h42452ff0, 32'h4295e8bc} /* (31, 1, 4) {real, imag} */,
  {32'h432748c3, 32'hc2aabca4} /* (31, 1, 3) {real, imag} */,
  {32'h44437dd2, 32'hc48d7892} /* (31, 1, 2) {real, imag} */,
  {32'hc45e807f, 32'h45051eba} /* (31, 1, 1) {real, imag} */,
  {32'hc232040d, 32'h44c01c98} /* (31, 1, 0) {real, imag} */,
  {32'h445bc1f9, 32'h445675ef} /* (31, 0, 31) {real, imag} */,
  {32'hc3d50e90, 32'hc2c58df6} /* (31, 0, 30) {real, imag} */,
  {32'h423a38f4, 32'hc286bc40} /* (31, 0, 29) {real, imag} */,
  {32'hc2e06a08, 32'hc30d5c72} /* (31, 0, 28) {real, imag} */,
  {32'h40be6a30, 32'hc3bfd37c} /* (31, 0, 27) {real, imag} */,
  {32'hc08f8df8, 32'h42c0b8a2} /* (31, 0, 26) {real, imag} */,
  {32'hc0ac0960, 32'hc1b68374} /* (31, 0, 25) {real, imag} */,
  {32'hc3899281, 32'hc1bc91ec} /* (31, 0, 24) {real, imag} */,
  {32'hc21f1a11, 32'hbffde300} /* (31, 0, 23) {real, imag} */,
  {32'h4154373c, 32'h41b547cc} /* (31, 0, 22) {real, imag} */,
  {32'hc1a615fa, 32'hc270ee88} /* (31, 0, 21) {real, imag} */,
  {32'hc2120f58, 32'h41464024} /* (31, 0, 20) {real, imag} */,
  {32'h41176424, 32'h41edb32f} /* (31, 0, 19) {real, imag} */,
  {32'hc1ff3ddc, 32'hc20bebe7} /* (31, 0, 18) {real, imag} */,
  {32'h41d87e6a, 32'hc283157d} /* (31, 0, 17) {real, imag} */,
  {32'hc1956bf6, 32'hc2a44970} /* (31, 0, 16) {real, imag} */,
  {32'hc1351dac, 32'hbe803b00} /* (31, 0, 15) {real, imag} */,
  {32'h42d50241, 32'hc11e3c64} /* (31, 0, 14) {real, imag} */,
  {32'hc159cafc, 32'h421c8662} /* (31, 0, 13) {real, imag} */,
  {32'hc1d84c51, 32'h41a1c50a} /* (31, 0, 12) {real, imag} */,
  {32'h40d0a398, 32'hc3176578} /* (31, 0, 11) {real, imag} */,
  {32'h42baf7b0, 32'hc2845a47} /* (31, 0, 10) {real, imag} */,
  {32'h41bca30e, 32'h411a0180} /* (31, 0, 9) {real, imag} */,
  {32'h42e3a46c, 32'h42595556} /* (31, 0, 8) {real, imag} */,
  {32'hc2ff74e2, 32'hc1950bdc} /* (31, 0, 7) {real, imag} */,
  {32'h4260fc19, 32'hc15582d0} /* (31, 0, 6) {real, imag} */,
  {32'h42842c5b, 32'hc3752670} /* (31, 0, 5) {real, imag} */,
  {32'h42f0c9cc, 32'hc26e3936} /* (31, 0, 4) {real, imag} */,
  {32'h4269853c, 32'h42319cdf} /* (31, 0, 3) {real, imag} */,
  {32'h43af9926, 32'hc3b5e602} /* (31, 0, 2) {real, imag} */,
  {32'hc4206ddd, 32'h44810077} /* (31, 0, 1) {real, imag} */,
  {32'h429ac1e8, 32'h445743c8} /* (31, 0, 0) {real, imag} */,
  {32'hc535cd5e, 32'hc550e473} /* (30, 31, 31) {real, imag} */,
  {32'h44ea9d8c, 32'h44a27ae8} /* (30, 31, 30) {real, imag} */,
  {32'hc314915b, 32'h4313d34a} /* (30, 31, 29) {real, imag} */,
  {32'hc3e05324, 32'hc35ea849} /* (30, 31, 28) {real, imag} */,
  {32'h44034d8e, 32'h440bc240} /* (30, 31, 27) {real, imag} */,
  {32'h42ff04f4, 32'h4149e850} /* (30, 31, 26) {real, imag} */,
  {32'hc35cb168, 32'hc2b74614} /* (30, 31, 25) {real, imag} */,
  {32'h44000f56, 32'h428d6e6a} /* (30, 31, 24) {real, imag} */,
  {32'h40f683f0, 32'hc190f330} /* (30, 31, 23) {real, imag} */,
  {32'h4303e908, 32'h42ba4ae6} /* (30, 31, 22) {real, imag} */,
  {32'h43348aa9, 32'h41935440} /* (30, 31, 21) {real, imag} */,
  {32'h4285ba76, 32'hc0122200} /* (30, 31, 20) {real, imag} */,
  {32'hc24a1bc6, 32'hc2e92971} /* (30, 31, 19) {real, imag} */,
  {32'h42daa5dc, 32'hc2880f20} /* (30, 31, 18) {real, imag} */,
  {32'hc12599c0, 32'h4214ded0} /* (30, 31, 17) {real, imag} */,
  {32'hc1f495a0, 32'h3eb71000} /* (30, 31, 16) {real, imag} */,
  {32'hbeed0800, 32'h41183ac0} /* (30, 31, 15) {real, imag} */,
  {32'hc2c8dfec, 32'h3f3cdfc0} /* (30, 31, 14) {real, imag} */,
  {32'hc1dffb5c, 32'hc234aa0a} /* (30, 31, 13) {real, imag} */,
  {32'hc1ecedd8, 32'hc0f741c0} /* (30, 31, 12) {real, imag} */,
  {32'hc283d576, 32'h438f4012} /* (30, 31, 11) {real, imag} */,
  {32'hc2d77f44, 32'hc2a65fbe} /* (30, 31, 10) {real, imag} */,
  {32'hc336faf0, 32'h430dc6d2} /* (30, 31, 9) {real, imag} */,
  {32'hc30f74cd, 32'h43558e1b} /* (30, 31, 8) {real, imag} */,
  {32'h42939891, 32'hc3478352} /* (30, 31, 7) {real, imag} */,
  {32'h43112d04, 32'h4374f8a7} /* (30, 31, 6) {real, imag} */,
  {32'h4363816a, 32'h44718c38} /* (30, 31, 5) {real, imag} */,
  {32'hc3dc86e2, 32'hc398e014} /* (30, 31, 4) {real, imag} */,
  {32'hc33a276d, 32'hc0a08ef0} /* (30, 31, 3) {real, imag} */,
  {32'h42ee0e68, 32'h44aaae7a} /* (30, 31, 2) {real, imag} */,
  {32'h42f86750, 32'hc529b903} /* (30, 31, 1) {real, imag} */,
  {32'hc444fd2f, 32'hc5165d50} /* (30, 31, 0) {real, imag} */,
  {32'hc1d752c0, 32'h4502118c} /* (30, 30, 31) {real, imag} */,
  {32'h42f4924e, 32'hc4d88acc} /* (30, 30, 30) {real, imag} */,
  {32'h427f2855, 32'h426102bb} /* (30, 30, 29) {real, imag} */,
  {32'h440941cd, 32'h444371a2} /* (30, 30, 28) {real, imag} */,
  {32'hc42d0160, 32'hc3a7ebff} /* (30, 30, 27) {real, imag} */,
  {32'hc229c644, 32'hc2cef88a} /* (30, 30, 26) {real, imag} */,
  {32'h417d2340, 32'h42d3eac6} /* (30, 30, 25) {real, imag} */,
  {32'hc35437c8, 32'hc32472d9} /* (30, 30, 24) {real, imag} */,
  {32'hc1d374dc, 32'h4299c1c2} /* (30, 30, 23) {real, imag} */,
  {32'h4260e2c8, 32'h42df0af2} /* (30, 30, 22) {real, imag} */,
  {32'hc34c73bc, 32'hc249b7f0} /* (30, 30, 21) {real, imag} */,
  {32'h41897b3c, 32'hc1aae894} /* (30, 30, 20) {real, imag} */,
  {32'h40cf13b8, 32'hbfc3a6e0} /* (30, 30, 19) {real, imag} */,
  {32'hc2c516ff, 32'hc14ef660} /* (30, 30, 18) {real, imag} */,
  {32'hc113da80, 32'h4289f61c} /* (30, 30, 17) {real, imag} */,
  {32'h416c4f00, 32'h42104af0} /* (30, 30, 16) {real, imag} */,
  {32'hc28a6250, 32'hbf837700} /* (30, 30, 15) {real, imag} */,
  {32'h429da34d, 32'hc28e0c74} /* (30, 30, 14) {real, imag} */,
  {32'hc1fe1406, 32'hc0aa9ec8} /* (30, 30, 13) {real, imag} */,
  {32'hc28cc899, 32'h429e415d} /* (30, 30, 12) {real, imag} */,
  {32'h43347ee8, 32'hc32d5de8} /* (30, 30, 11) {real, imag} */,
  {32'hc21ab112, 32'hc097bb28} /* (30, 30, 10) {real, imag} */,
  {32'hc2c692e9, 32'hc28a3f12} /* (30, 30, 9) {real, imag} */,
  {32'h438674f9, 32'hc3504f33} /* (30, 30, 8) {real, imag} */,
  {32'hc384c80a, 32'h439a4332} /* (30, 30, 7) {real, imag} */,
  {32'h4251e8b6, 32'hc344ec63} /* (30, 30, 6) {real, imag} */,
  {32'h433b54cc, 32'hc436aff8} /* (30, 30, 5) {real, imag} */,
  {32'hc4166c53, 32'h43a100cd} /* (30, 30, 4) {real, imag} */,
  {32'h43111e9e, 32'h4208e9f5} /* (30, 30, 3) {real, imag} */,
  {32'h434e8cc1, 32'hc507abd6} /* (30, 30, 2) {real, imag} */,
  {32'h44504766, 32'h4552372c} /* (30, 30, 1) {real, imag} */,
  {32'h440b7060, 32'h44a7e604} /* (30, 30, 0) {real, imag} */,
  {32'hc3f400a4, 32'hc39df32a} /* (30, 29, 31) {real, imag} */,
  {32'h44352fb9, 32'hc13b9de0} /* (30, 29, 30) {real, imag} */,
  {32'hc1db2dc5, 32'h42e4cca9} /* (30, 29, 29) {real, imag} */,
  {32'hc2161dc2, 32'h426bed58} /* (30, 29, 28) {real, imag} */,
  {32'hc3218b7a, 32'hc364fb5d} /* (30, 29, 27) {real, imag} */,
  {32'hc2b355fb, 32'h43030ae2} /* (30, 29, 26) {real, imag} */,
  {32'hc2605cc2, 32'hc2848912} /* (30, 29, 25) {real, imag} */,
  {32'h4318fe81, 32'h41c77a6a} /* (30, 29, 24) {real, imag} */,
  {32'hc2180585, 32'h4287be34} /* (30, 29, 23) {real, imag} */,
  {32'h428d4bef, 32'h42efb46c} /* (30, 29, 22) {real, imag} */,
  {32'hc238b2a0, 32'hc2edc01c} /* (30, 29, 21) {real, imag} */,
  {32'h41934b14, 32'hc15f4074} /* (30, 29, 20) {real, imag} */,
  {32'h41f78b43, 32'hc17896a8} /* (30, 29, 19) {real, imag} */,
  {32'h428cf004, 32'hc153c000} /* (30, 29, 18) {real, imag} */,
  {32'h40e9bca0, 32'h405fb680} /* (30, 29, 17) {real, imag} */,
  {32'hc2777611, 32'hc093b554} /* (30, 29, 16) {real, imag} */,
  {32'hbf8dd180, 32'h4186e470} /* (30, 29, 15) {real, imag} */,
  {32'hc0f16c38, 32'hc0835300} /* (30, 29, 14) {real, imag} */,
  {32'hc108beee, 32'h4246e10e} /* (30, 29, 13) {real, imag} */,
  {32'hc1935bd4, 32'h416cab7c} /* (30, 29, 12) {real, imag} */,
  {32'hc2239768, 32'h42c2bb68} /* (30, 29, 11) {real, imag} */,
  {32'hc31025b4, 32'hc277ac0b} /* (30, 29, 10) {real, imag} */,
  {32'hc314d4f1, 32'hc27311a9} /* (30, 29, 9) {real, imag} */,
  {32'h43148a29, 32'hc01ff6c0} /* (30, 29, 8) {real, imag} */,
  {32'hc047e840, 32'hc306bf7d} /* (30, 29, 7) {real, imag} */,
  {32'hc2e6903b, 32'hc1a7a94a} /* (30, 29, 6) {real, imag} */,
  {32'h425be0f6, 32'h437cc279} /* (30, 29, 5) {real, imag} */,
  {32'hc38652ad, 32'hc38ee5df} /* (30, 29, 4) {real, imag} */,
  {32'hc2a96350, 32'h40c90cd0} /* (30, 29, 3) {real, imag} */,
  {32'h440b30b7, 32'hc43bec5e} /* (30, 29, 2) {real, imag} */,
  {32'hc335e400, 32'h44344a9b} /* (30, 29, 1) {real, imag} */,
  {32'hc2829084, 32'h42084102} /* (30, 29, 0) {real, imag} */,
  {32'hc3f06a2b, 32'hc480ec20} /* (30, 28, 31) {real, imag} */,
  {32'h44263759, 32'h43e8793e} /* (30, 28, 30) {real, imag} */,
  {32'hc236d12d, 32'hc2f166d7} /* (30, 28, 29) {real, imag} */,
  {32'hc372ce66, 32'hc300ffd4} /* (30, 28, 28) {real, imag} */,
  {32'h4336ef7a, 32'hc279dcce} /* (30, 28, 27) {real, imag} */,
  {32'h406d4e20, 32'h428c759b} /* (30, 28, 26) {real, imag} */,
  {32'hc10807ba, 32'hc2bbc9fa} /* (30, 28, 25) {real, imag} */,
  {32'h4324bb09, 32'hc07beed0} /* (30, 28, 24) {real, imag} */,
  {32'h41f3947c, 32'hc12eb710} /* (30, 28, 23) {real, imag} */,
  {32'hc28aa077, 32'h42391356} /* (30, 28, 22) {real, imag} */,
  {32'hc0426530, 32'h408e0bb0} /* (30, 28, 21) {real, imag} */,
  {32'h42b9fad0, 32'h4244051a} /* (30, 28, 20) {real, imag} */,
  {32'h40cd5ada, 32'hc21455c8} /* (30, 28, 19) {real, imag} */,
  {32'h422c9ae9, 32'hc0859458} /* (30, 28, 18) {real, imag} */,
  {32'h41c00a6c, 32'h420ce950} /* (30, 28, 17) {real, imag} */,
  {32'h41b8f010, 32'h41c0fc28} /* (30, 28, 16) {real, imag} */,
  {32'hc283681b, 32'hc0fd2080} /* (30, 28, 15) {real, imag} */,
  {32'h415a3cdc, 32'h414915ec} /* (30, 28, 14) {real, imag} */,
  {32'h3f267730, 32'h4009e340} /* (30, 28, 13) {real, imag} */,
  {32'h422fdbb0, 32'h414d24f8} /* (30, 28, 12) {real, imag} */,
  {32'hc2aadc0e, 32'h433571c0} /* (30, 28, 11) {real, imag} */,
  {32'h4224a7d6, 32'hc2ccc689} /* (30, 28, 10) {real, imag} */,
  {32'hc2a80881, 32'hc2969d7c} /* (30, 28, 9) {real, imag} */,
  {32'hc0d46fa0, 32'h430187a7} /* (30, 28, 8) {real, imag} */,
  {32'hc28ecc47, 32'hc0b5bd00} /* (30, 28, 7) {real, imag} */,
  {32'hc30e7f8e, 32'hc2b71bd9} /* (30, 28, 6) {real, imag} */,
  {32'hc2902c7b, 32'h434257ba} /* (30, 28, 5) {real, imag} */,
  {32'hc2b81cbb, 32'hc3b18e05} /* (30, 28, 4) {real, imag} */,
  {32'h41238644, 32'h41e94cc4} /* (30, 28, 3) {real, imag} */,
  {32'h44075289, 32'h43d781f0} /* (30, 28, 2) {real, imag} */,
  {32'hc4142e20, 32'hc3478754} /* (30, 28, 1) {real, imag} */,
  {32'hc2ccc3d9, 32'hc34b0f31} /* (30, 28, 0) {real, imag} */,
  {32'h44073fac, 32'h43fd65db} /* (30, 27, 31) {real, imag} */,
  {32'hc324119d, 32'hc290588e} /* (30, 27, 30) {real, imag} */,
  {32'h42ad02e2, 32'h420044f4} /* (30, 27, 29) {real, imag} */,
  {32'h431a14bd, 32'h42e80a69} /* (30, 27, 28) {real, imag} */,
  {32'hc3c4e768, 32'hc3a726d8} /* (30, 27, 27) {real, imag} */,
  {32'hc2abd1c8, 32'h42e3a448} /* (30, 27, 26) {real, imag} */,
  {32'h42872f95, 32'hc080750c} /* (30, 27, 25) {real, imag} */,
  {32'hc308d338, 32'hc2a0bc11} /* (30, 27, 24) {real, imag} */,
  {32'h419b2f0c, 32'hc265f546} /* (30, 27, 23) {real, imag} */,
  {32'hc0d461d8, 32'h429c1cd8} /* (30, 27, 22) {real, imag} */,
  {32'hc2e95f5e, 32'hc1b4b37c} /* (30, 27, 21) {real, imag} */,
  {32'hc20d1eef, 32'hc2838256} /* (30, 27, 20) {real, imag} */,
  {32'h41e24444, 32'h41c47288} /* (30, 27, 19) {real, imag} */,
  {32'hc1d8253c, 32'h423a27f6} /* (30, 27, 18) {real, imag} */,
  {32'hc2050210, 32'h4201c9be} /* (30, 27, 17) {real, imag} */,
  {32'h411c84f0, 32'hc0c7ad40} /* (30, 27, 16) {real, imag} */,
  {32'h423659b8, 32'hc11533f8} /* (30, 27, 15) {real, imag} */,
  {32'h426a980e, 32'hc2460022} /* (30, 27, 14) {real, imag} */,
  {32'hc2120d2e, 32'h413361f0} /* (30, 27, 13) {real, imag} */,
  {32'hc1fe53be, 32'hc0337970} /* (30, 27, 12) {real, imag} */,
  {32'h41b72698, 32'hc31ad7da} /* (30, 27, 11) {real, imag} */,
  {32'h4218b85e, 32'hc2acb31a} /* (30, 27, 10) {real, imag} */,
  {32'hc25e3f3a, 32'h4186429b} /* (30, 27, 9) {real, imag} */,
  {32'h42672788, 32'hc2f41657} /* (30, 27, 8) {real, imag} */,
  {32'hc212f7f6, 32'h404bfca8} /* (30, 27, 7) {real, imag} */,
  {32'h428932ca, 32'hc2077585} /* (30, 27, 6) {real, imag} */,
  {32'h42e0f64a, 32'hc38c2b24} /* (30, 27, 5) {real, imag} */,
  {32'hc31f9d65, 32'h42edf1db} /* (30, 27, 4) {real, imag} */,
  {32'hc1a9bbf8, 32'hc2dd3276} /* (30, 27, 3) {real, imag} */,
  {32'hc29e0562, 32'hc39b9fa6} /* (30, 27, 2) {real, imag} */,
  {32'h439c9aa8, 32'h444bda3a} /* (30, 27, 1) {real, imag} */,
  {32'h43b3e0ba, 32'h440d0ebe} /* (30, 27, 0) {real, imag} */,
  {32'h4266f9b8, 32'h429fe056} /* (30, 26, 31) {real, imag} */,
  {32'h42e4231d, 32'hc33dd510} /* (30, 26, 30) {real, imag} */,
  {32'hc2c53ab4, 32'hc2841f25} /* (30, 26, 29) {real, imag} */,
  {32'h41aa2fde, 32'hc22c441f} /* (30, 26, 28) {real, imag} */,
  {32'h420778c7, 32'hc24cce52} /* (30, 26, 27) {real, imag} */,
  {32'hc291d2e7, 32'hc29c6dfa} /* (30, 26, 26) {real, imag} */,
  {32'h4257e242, 32'h41d5bb02} /* (30, 26, 25) {real, imag} */,
  {32'hc23ea4b8, 32'hc2caf836} /* (30, 26, 24) {real, imag} */,
  {32'h426cb950, 32'hc2305eb5} /* (30, 26, 23) {real, imag} */,
  {32'h40f0e514, 32'h42c39b07} /* (30, 26, 22) {real, imag} */,
  {32'hc185d116, 32'hc23171f8} /* (30, 26, 21) {real, imag} */,
  {32'h416e8b67, 32'h41d35656} /* (30, 26, 20) {real, imag} */,
  {32'hc265ba30, 32'hc19dc17a} /* (30, 26, 19) {real, imag} */,
  {32'h414b11b9, 32'h42080739} /* (30, 26, 18) {real, imag} */,
  {32'h413c6d3c, 32'hc0a11078} /* (30, 26, 17) {real, imag} */,
  {32'hc19adb9e, 32'hc10dd4fc} /* (30, 26, 16) {real, imag} */,
  {32'h40923857, 32'h414fc5cc} /* (30, 26, 15) {real, imag} */,
  {32'h40d320e2, 32'h40809e1a} /* (30, 26, 14) {real, imag} */,
  {32'h41e620cb, 32'h40905a47} /* (30, 26, 13) {real, imag} */,
  {32'hc1460155, 32'hc1fccf56} /* (30, 26, 12) {real, imag} */,
  {32'hc23fa2d1, 32'hc25273bc} /* (30, 26, 11) {real, imag} */,
  {32'h40deb9fc, 32'hc1af409c} /* (30, 26, 10) {real, imag} */,
  {32'hc15a81ee, 32'hc04eac50} /* (30, 26, 9) {real, imag} */,
  {32'hc2a1a9c2, 32'hc230456c} /* (30, 26, 8) {real, imag} */,
  {32'hc155c86a, 32'h421b2191} /* (30, 26, 7) {real, imag} */,
  {32'hc2716d2a, 32'hc1770220} /* (30, 26, 6) {real, imag} */,
  {32'hc284ce94, 32'h427cf65a} /* (30, 26, 5) {real, imag} */,
  {32'hc2746029, 32'hc265aafd} /* (30, 26, 4) {real, imag} */,
  {32'h41ac1bce, 32'h42684065} /* (30, 26, 3) {real, imag} */,
  {32'hc2995c37, 32'hc2ec7520} /* (30, 26, 2) {real, imag} */,
  {32'h428fd7fc, 32'hc26c843d} /* (30, 26, 1) {real, imag} */,
  {32'hc29dea26, 32'h428c6068} /* (30, 26, 0) {real, imag} */,
  {32'hc36fd513, 32'hc302e5ff} /* (30, 25, 31) {real, imag} */,
  {32'h4287b135, 32'h41ab2952} /* (30, 25, 30) {real, imag} */,
  {32'h4298b422, 32'h43550ebe} /* (30, 25, 29) {real, imag} */,
  {32'hc2700f04, 32'h40630dc6} /* (30, 25, 28) {real, imag} */,
  {32'h428c1f8c, 32'h42ae5ab1} /* (30, 25, 27) {real, imag} */,
  {32'hc22d6c51, 32'h4155f5e7} /* (30, 25, 26) {real, imag} */,
  {32'hc1284eb8, 32'hc3325ac3} /* (30, 25, 25) {real, imag} */,
  {32'h415594f0, 32'h4284e04c} /* (30, 25, 24) {real, imag} */,
  {32'hc1a827f4, 32'h4280c9ae} /* (30, 25, 23) {real, imag} */,
  {32'h41866b04, 32'hc1bde736} /* (30, 25, 22) {real, imag} */,
  {32'h425457e3, 32'hc286bd30} /* (30, 25, 21) {real, imag} */,
  {32'h41c1445a, 32'hc1b16f34} /* (30, 25, 20) {real, imag} */,
  {32'h4060bb3c, 32'h4168b740} /* (30, 25, 19) {real, imag} */,
  {32'hbf6d9400, 32'hc1dbe4c7} /* (30, 25, 18) {real, imag} */,
  {32'h41d01222, 32'hc175274c} /* (30, 25, 17) {real, imag} */,
  {32'hc0a4c510, 32'hc11eb480} /* (30, 25, 16) {real, imag} */,
  {32'h3fb90060, 32'h41555f3c} /* (30, 25, 15) {real, imag} */,
  {32'hc24bebae, 32'h415dc0aa} /* (30, 25, 14) {real, imag} */,
  {32'hc009e154, 32'hc1e5af00} /* (30, 25, 13) {real, imag} */,
  {32'hc207c762, 32'h41189ea6} /* (30, 25, 12) {real, imag} */,
  {32'h41e8bc02, 32'hc2bbabb6} /* (30, 25, 11) {real, imag} */,
  {32'hc0f37354, 32'h41c0124e} /* (30, 25, 10) {real, imag} */,
  {32'h42c6f857, 32'hc178de30} /* (30, 25, 9) {real, imag} */,
  {32'h425e6638, 32'h40e42340} /* (30, 25, 8) {real, imag} */,
  {32'hc26e6242, 32'h411d2530} /* (30, 25, 7) {real, imag} */,
  {32'h41612a03, 32'h41c7ca80} /* (30, 25, 6) {real, imag} */,
  {32'h4219960b, 32'h429064a5} /* (30, 25, 5) {real, imag} */,
  {32'hc1ed21cf, 32'h41141120} /* (30, 25, 4) {real, imag} */,
  {32'hc228be51, 32'hbe802000} /* (30, 25, 3) {real, imag} */,
  {32'h42e81867, 32'h42ba0e5a} /* (30, 25, 2) {real, imag} */,
  {32'hc18db408, 32'hc32b26e5} /* (30, 25, 1) {real, imag} */,
  {32'hc2e43bf9, 32'hc32e1050} /* (30, 25, 0) {real, imag} */,
  {32'h43901023, 32'h43243157} /* (30, 24, 31) {real, imag} */,
  {32'hc3152f81, 32'hc351d054} /* (30, 24, 30) {real, imag} */,
  {32'hc2eebe20, 32'hc28f2050} /* (30, 24, 29) {real, imag} */,
  {32'h42accfc2, 32'h43273daa} /* (30, 24, 28) {real, imag} */,
  {32'hc2576e3e, 32'hc315dee9} /* (30, 24, 27) {real, imag} */,
  {32'h3e520e00, 32'h40c633b8} /* (30, 24, 26) {real, imag} */,
  {32'hc2eb7692, 32'hc266dbe0} /* (30, 24, 25) {real, imag} */,
  {32'h42a58fd0, 32'hc0dd5e80} /* (30, 24, 24) {real, imag} */,
  {32'h426798c5, 32'h41e44078} /* (30, 24, 23) {real, imag} */,
  {32'hc0d429a0, 32'hc155b45c} /* (30, 24, 22) {real, imag} */,
  {32'hc231212e, 32'hc168aaa7} /* (30, 24, 21) {real, imag} */,
  {32'hc1e0cc30, 32'hc0c0fdf8} /* (30, 24, 20) {real, imag} */,
  {32'hc16a6c9b, 32'hbf5db2f0} /* (30, 24, 19) {real, imag} */,
  {32'h4121f701, 32'hc155b7d4} /* (30, 24, 18) {real, imag} */,
  {32'h4186fbd8, 32'h41c53c18} /* (30, 24, 17) {real, imag} */,
  {32'hc1feae98, 32'hc1cd6df6} /* (30, 24, 16) {real, imag} */,
  {32'hbf307700, 32'hc13181b0} /* (30, 24, 15) {real, imag} */,
  {32'h41d07c40, 32'hc14c796c} /* (30, 24, 14) {real, imag} */,
  {32'h40a198ea, 32'h41bff2a4} /* (30, 24, 13) {real, imag} */,
  {32'hc2075e9c, 32'hc1c401de} /* (30, 24, 12) {real, imag} */,
  {32'h41ee1014, 32'hc227141c} /* (30, 24, 11) {real, imag} */,
  {32'hc22c508c, 32'h418f452a} /* (30, 24, 10) {real, imag} */,
  {32'h4284f416, 32'hc1a8a870} /* (30, 24, 9) {real, imag} */,
  {32'hc2ab5d06, 32'hc3101e94} /* (30, 24, 8) {real, imag} */,
  {32'h42ff5bea, 32'hc1902a48} /* (30, 24, 7) {real, imag} */,
  {32'hc2ea0d5d, 32'hc1bdcb7a} /* (30, 24, 6) {real, imag} */,
  {32'hc1f8c5b4, 32'hc2870e92} /* (30, 24, 5) {real, imag} */,
  {32'h3fd68a80, 32'hc1c91c40} /* (30, 24, 4) {real, imag} */,
  {32'h4253555f, 32'h42d7e9f8} /* (30, 24, 3) {real, imag} */,
  {32'hc33f0c4f, 32'hc3d06838} /* (30, 24, 2) {real, imag} */,
  {32'h43b5c157, 32'h44112adc} /* (30, 24, 1) {real, imag} */,
  {32'h433dd339, 32'h430f6562} /* (30, 24, 0) {real, imag} */,
  {32'hc29451ae, 32'hc33904e8} /* (30, 23, 31) {real, imag} */,
  {32'h42ad8888, 32'hc2e01ff8} /* (30, 23, 30) {real, imag} */,
  {32'hc20fb737, 32'h41e857b9} /* (30, 23, 29) {real, imag} */,
  {32'hc2873486, 32'h42170552} /* (30, 23, 28) {real, imag} */,
  {32'hc2abb5f9, 32'h42237ff0} /* (30, 23, 27) {real, imag} */,
  {32'h4178b5e8, 32'h41592062} /* (30, 23, 26) {real, imag} */,
  {32'hc20a5f27, 32'h424c0c1a} /* (30, 23, 25) {real, imag} */,
  {32'hc15aed62, 32'hc1140442} /* (30, 23, 24) {real, imag} */,
  {32'h426f050b, 32'h41d67fb1} /* (30, 23, 23) {real, imag} */,
  {32'hc28e002f, 32'h425c61a8} /* (30, 23, 22) {real, imag} */,
  {32'hc1c7aa18, 32'hc17ab444} /* (30, 23, 21) {real, imag} */,
  {32'hc199486c, 32'h4019d0c8} /* (30, 23, 20) {real, imag} */,
  {32'h41c3632e, 32'hc1699866} /* (30, 23, 19) {real, imag} */,
  {32'hc20c1f7e, 32'hc0e1d778} /* (30, 23, 18) {real, imag} */,
  {32'h410ecd4d, 32'hc10bf496} /* (30, 23, 17) {real, imag} */,
  {32'hc1730038, 32'hc1672c50} /* (30, 23, 16) {real, imag} */,
  {32'h416ff52b, 32'h42005432} /* (30, 23, 15) {real, imag} */,
  {32'h422d80e2, 32'h41a1496e} /* (30, 23, 14) {real, imag} */,
  {32'hc07f0694, 32'hc21ae0b2} /* (30, 23, 13) {real, imag} */,
  {32'h4172a2c0, 32'h42175f02} /* (30, 23, 12) {real, imag} */,
  {32'h409fd91e, 32'h41e670be} /* (30, 23, 11) {real, imag} */,
  {32'hc1100568, 32'h416480a2} /* (30, 23, 10) {real, imag} */,
  {32'hc24c4c6f, 32'hc24c36e2} /* (30, 23, 9) {real, imag} */,
  {32'h4241bf96, 32'h426776c6} /* (30, 23, 8) {real, imag} */,
  {32'h41ce223e, 32'hc217bfcc} /* (30, 23, 7) {real, imag} */,
  {32'h426bfe36, 32'hc1d8d551} /* (30, 23, 6) {real, imag} */,
  {32'h4199915c, 32'h43359284} /* (30, 23, 5) {real, imag} */,
  {32'hc21c96d7, 32'hc1bdd2e2} /* (30, 23, 4) {real, imag} */,
  {32'hc29015e6, 32'hc2ab9c58} /* (30, 23, 3) {real, imag} */,
  {32'h433fd624, 32'hc32a173e} /* (30, 23, 2) {real, imag} */,
  {32'hc2f8a35a, 32'h435f6d6a} /* (30, 23, 1) {real, imag} */,
  {32'h424aa00c, 32'h420d744b} /* (30, 23, 0) {real, imag} */,
  {32'hc2baa7d5, 32'hc327cda6} /* (30, 22, 31) {real, imag} */,
  {32'h432f0482, 32'h41daf4d2} /* (30, 22, 30) {real, imag} */,
  {32'hc0b536f4, 32'h424c774e} /* (30, 22, 29) {real, imag} */,
  {32'hc2ba2af8, 32'h423be002} /* (30, 22, 28) {real, imag} */,
  {32'h3e391ac0, 32'hc1cd0e9e} /* (30, 22, 27) {real, imag} */,
  {32'h422292d6, 32'h4266c934} /* (30, 22, 26) {real, imag} */,
  {32'h415bbe62, 32'hc2ddf52c} /* (30, 22, 25) {real, imag} */,
  {32'hc24a2445, 32'hc21760e7} /* (30, 22, 24) {real, imag} */,
  {32'h42350a76, 32'hc27b559a} /* (30, 22, 23) {real, imag} */,
  {32'h42aa2bec, 32'h42018c54} /* (30, 22, 22) {real, imag} */,
  {32'h4024c698, 32'hc2100391} /* (30, 22, 21) {real, imag} */,
  {32'hc24553db, 32'hc0e65624} /* (30, 22, 20) {real, imag} */,
  {32'h41ecc631, 32'h41b38fcc} /* (30, 22, 19) {real, imag} */,
  {32'h41073b3a, 32'h4092f108} /* (30, 22, 18) {real, imag} */,
  {32'hc1e9fdbf, 32'h41769b22} /* (30, 22, 17) {real, imag} */,
  {32'hc1aec4c2, 32'hbf444240} /* (30, 22, 16) {real, imag} */,
  {32'hc1bdc029, 32'hc19d826d} /* (30, 22, 15) {real, imag} */,
  {32'h41c0c61b, 32'h412032ca} /* (30, 22, 14) {real, imag} */,
  {32'h41c8d53f, 32'h41d11e9c} /* (30, 22, 13) {real, imag} */,
  {32'hc19af9fa, 32'h41d53585} /* (30, 22, 12) {real, imag} */,
  {32'hc216e702, 32'h41a2d40e} /* (30, 22, 11) {real, imag} */,
  {32'hbfea4c20, 32'hc24c9420} /* (30, 22, 10) {real, imag} */,
  {32'hc260d6da, 32'hc220df5a} /* (30, 22, 9) {real, imag} */,
  {32'h4255b0d7, 32'h41954fd2} /* (30, 22, 8) {real, imag} */,
  {32'hbf8ef1ac, 32'h4159de60} /* (30, 22, 7) {real, imag} */,
  {32'h41fdd627, 32'hc26013e4} /* (30, 22, 6) {real, imag} */,
  {32'h41869264, 32'h42a18892} /* (30, 22, 5) {real, imag} */,
  {32'h41d3c7de, 32'hc246efe6} /* (30, 22, 4) {real, imag} */,
  {32'hc1e0982b, 32'hc2e47be9} /* (30, 22, 3) {real, imag} */,
  {32'h42f391fb, 32'h415bc58b} /* (30, 22, 2) {real, imag} */,
  {32'hc34aff5e, 32'hc281f45c} /* (30, 22, 1) {real, imag} */,
  {32'hc20f9265, 32'hc25f01b5} /* (30, 22, 0) {real, imag} */,
  {32'h437f268b, 32'h40d725a8} /* (30, 21, 31) {real, imag} */,
  {32'hc35abadc, 32'h42d3deda} /* (30, 21, 30) {real, imag} */,
  {32'hc2b1fdbe, 32'hc26f4b50} /* (30, 21, 29) {real, imag} */,
  {32'hc18591ee, 32'h41f35683} /* (30, 21, 28) {real, imag} */,
  {32'hc21a4298, 32'h410ac690} /* (30, 21, 27) {real, imag} */,
  {32'h42087ba0, 32'h418d4d40} /* (30, 21, 26) {real, imag} */,
  {32'h4067e5c0, 32'h422691ce} /* (30, 21, 25) {real, imag} */,
  {32'h40ff78c0, 32'hc1d1d204} /* (30, 21, 24) {real, imag} */,
  {32'hc217dfa5, 32'hc2911108} /* (30, 21, 23) {real, imag} */,
  {32'h42289506, 32'hbd11a500} /* (30, 21, 22) {real, imag} */,
  {32'hc1bcbc84, 32'h42680c92} /* (30, 21, 21) {real, imag} */,
  {32'hc1b214c2, 32'hc1c69456} /* (30, 21, 20) {real, imag} */,
  {32'h411a6802, 32'h4165c86e} /* (30, 21, 19) {real, imag} */,
  {32'h402c17e8, 32'hc1f8d454} /* (30, 21, 18) {real, imag} */,
  {32'h414e8726, 32'hc0c2d7d8} /* (30, 21, 17) {real, imag} */,
  {32'hc0e8ae80, 32'h414c01e0} /* (30, 21, 16) {real, imag} */,
  {32'h3fa159d0, 32'hc062bc10} /* (30, 21, 15) {real, imag} */,
  {32'h41943a03, 32'h41b19f74} /* (30, 21, 14) {real, imag} */,
  {32'hc1b2fa69, 32'h41976b8d} /* (30, 21, 13) {real, imag} */,
  {32'hc1c39266, 32'hc14c57b0} /* (30, 21, 12) {real, imag} */,
  {32'hc102d655, 32'hc210971c} /* (30, 21, 11) {real, imag} */,
  {32'h419161e5, 32'h4169e697} /* (30, 21, 10) {real, imag} */,
  {32'h42305ead, 32'h4229fd46} /* (30, 21, 9) {real, imag} */,
  {32'hc08def00, 32'h41910a5c} /* (30, 21, 8) {real, imag} */,
  {32'h42103c38, 32'hc0ea89a0} /* (30, 21, 7) {real, imag} */,
  {32'h42813fec, 32'hc2427f08} /* (30, 21, 6) {real, imag} */,
  {32'hc15a71d2, 32'h418c84fc} /* (30, 21, 5) {real, imag} */,
  {32'hc23f1ee5, 32'hc21c0493} /* (30, 21, 4) {real, imag} */,
  {32'h4023e340, 32'hc277a786} /* (30, 21, 3) {real, imag} */,
  {32'hc2fe1270, 32'hc31ed873} /* (30, 21, 2) {real, imag} */,
  {32'h43142643, 32'h42fd49c0} /* (30, 21, 1) {real, imag} */,
  {32'h4389ce5d, 32'h43778516} /* (30, 21, 0) {real, imag} */,
  {32'h418dbb10, 32'hc24edcce} /* (30, 20, 31) {real, imag} */,
  {32'hc168bfc4, 32'h420b29d9} /* (30, 20, 30) {real, imag} */,
  {32'hc22447cc, 32'hc2b9c513} /* (30, 20, 29) {real, imag} */,
  {32'hc1782abd, 32'h42292714} /* (30, 20, 28) {real, imag} */,
  {32'hc185177c, 32'h42873e2c} /* (30, 20, 27) {real, imag} */,
  {32'h421f481d, 32'h41fbad7e} /* (30, 20, 26) {real, imag} */,
  {32'hc050fca8, 32'h3fedfb68} /* (30, 20, 25) {real, imag} */,
  {32'h425d92be, 32'h4267b706} /* (30, 20, 24) {real, imag} */,
  {32'h416fa592, 32'h40cb4ac0} /* (30, 20, 23) {real, imag} */,
  {32'hc15cc9ad, 32'hc2277931} /* (30, 20, 22) {real, imag} */,
  {32'h4128b3b2, 32'hc1746ab6} /* (30, 20, 21) {real, imag} */,
  {32'hc19e9020, 32'h4173ed3c} /* (30, 20, 20) {real, imag} */,
  {32'h4193eb3e, 32'hc13aedce} /* (30, 20, 19) {real, imag} */,
  {32'hc1005a66, 32'h418b997e} /* (30, 20, 18) {real, imag} */,
  {32'hc091b126, 32'h40fca8c5} /* (30, 20, 17) {real, imag} */,
  {32'hbee326a0, 32'hc108a782} /* (30, 20, 16) {real, imag} */,
  {32'hc14593a3, 32'h416812a2} /* (30, 20, 15) {real, imag} */,
  {32'hbe506700, 32'hc188490a} /* (30, 20, 14) {real, imag} */,
  {32'hc1a30b8a, 32'h3edf8640} /* (30, 20, 13) {real, imag} */,
  {32'hc13541c5, 32'h3fe96030} /* (30, 20, 12) {real, imag} */,
  {32'h40ef1290, 32'h41373b0a} /* (30, 20, 11) {real, imag} */,
  {32'hc18a4af6, 32'hc1c51ec2} /* (30, 20, 10) {real, imag} */,
  {32'h40c84b5c, 32'hbeb72958} /* (30, 20, 9) {real, imag} */,
  {32'h422e814e, 32'hc080e754} /* (30, 20, 8) {real, imag} */,
  {32'hc21d679e, 32'h41a80a1c} /* (30, 20, 7) {real, imag} */,
  {32'h421db3c1, 32'h42806a92} /* (30, 20, 6) {real, imag} */,
  {32'hc1daf9d8, 32'hc224ce90} /* (30, 20, 5) {real, imag} */,
  {32'hc0ca665e, 32'h41889a34} /* (30, 20, 4) {real, imag} */,
  {32'h42204db8, 32'h42cb0d8d} /* (30, 20, 3) {real, imag} */,
  {32'h41b40982, 32'hc27805bf} /* (30, 20, 2) {real, imag} */,
  {32'hc1ab62a4, 32'hc2213c8a} /* (30, 20, 1) {real, imag} */,
  {32'hc1cefb2e, 32'hc0c52ea4} /* (30, 20, 0) {real, imag} */,
  {32'hc21c7d97, 32'h4113550c} /* (30, 19, 31) {real, imag} */,
  {32'hc20e4f1e, 32'h4167abe4} /* (30, 19, 30) {real, imag} */,
  {32'hbfac7780, 32'h41502be0} /* (30, 19, 29) {real, imag} */,
  {32'hc1d5883a, 32'h421ecb61} /* (30, 19, 28) {real, imag} */,
  {32'hc23a846c, 32'h400dae3e} /* (30, 19, 27) {real, imag} */,
  {32'h41b14bf2, 32'h41afa850} /* (30, 19, 26) {real, imag} */,
  {32'hbff48120, 32'hc28a2cf8} /* (30, 19, 25) {real, imag} */,
  {32'h40ad8211, 32'h41cc66da} /* (30, 19, 24) {real, imag} */,
  {32'h40c1d43a, 32'h401d8de4} /* (30, 19, 23) {real, imag} */,
  {32'hc0819c50, 32'hc0af7925} /* (30, 19, 22) {real, imag} */,
  {32'h4118ac56, 32'hc12867be} /* (30, 19, 21) {real, imag} */,
  {32'h3fe0b58c, 32'h41d4fb50} /* (30, 19, 20) {real, imag} */,
  {32'hc047586c, 32'hc12ea9fa} /* (30, 19, 19) {real, imag} */,
  {32'hc02baa00, 32'hc1ce3f2c} /* (30, 19, 18) {real, imag} */,
  {32'h405abb88, 32'h402d98d4} /* (30, 19, 17) {real, imag} */,
  {32'h40a59fea, 32'hc032be80} /* (30, 19, 16) {real, imag} */,
  {32'hc0190918, 32'hc11f43dc} /* (30, 19, 15) {real, imag} */,
  {32'hbf04cf80, 32'h4134fb20} /* (30, 19, 14) {real, imag} */,
  {32'hc08ba44a, 32'h40b181ff} /* (30, 19, 13) {real, imag} */,
  {32'h40c73917, 32'hc0b01e1a} /* (30, 19, 12) {real, imag} */,
  {32'hbecd9cc0, 32'hbfdec99c} /* (30, 19, 11) {real, imag} */,
  {32'hc084d18c, 32'h4182db12} /* (30, 19, 10) {real, imag} */,
  {32'hc19d8fe6, 32'h3f925a28} /* (30, 19, 9) {real, imag} */,
  {32'hc11bfbee, 32'hc18b2236} /* (30, 19, 8) {real, imag} */,
  {32'h420976df, 32'h41968840} /* (30, 19, 7) {real, imag} */,
  {32'hc147d7c5, 32'hc0a5688a} /* (30, 19, 6) {real, imag} */,
  {32'hc1c52af1, 32'h4156f4d8} /* (30, 19, 5) {real, imag} */,
  {32'h4124dbf4, 32'hc18e3978} /* (30, 19, 4) {real, imag} */,
  {32'hc1af012f, 32'hbfdb01f4} /* (30, 19, 3) {real, imag} */,
  {32'h4269bf58, 32'hc229cfc1} /* (30, 19, 2) {real, imag} */,
  {32'h3fd7c3a0, 32'h41ebf86a} /* (30, 19, 1) {real, imag} */,
  {32'h41027bfb, 32'hc225661a} /* (30, 19, 0) {real, imag} */,
  {32'h42bf9ba8, 32'hc1988f2a} /* (30, 18, 31) {real, imag} */,
  {32'hc2b727d4, 32'hc0d7ee10} /* (30, 18, 30) {real, imag} */,
  {32'hc1d74ed8, 32'h401a21d0} /* (30, 18, 29) {real, imag} */,
  {32'h42a251fd, 32'h42b12ff6} /* (30, 18, 28) {real, imag} */,
  {32'hc1b537e2, 32'h40ba9aea} /* (30, 18, 27) {real, imag} */,
  {32'hc1d81212, 32'hc02d2b4a} /* (30, 18, 26) {real, imag} */,
  {32'h423b57ea, 32'h410bbe92} /* (30, 18, 25) {real, imag} */,
  {32'hc162c96c, 32'h413b8c77} /* (30, 18, 24) {real, imag} */,
  {32'hc12f97a2, 32'h412f915e} /* (30, 18, 23) {real, imag} */,
  {32'h3e27c280, 32'h408c1b3a} /* (30, 18, 22) {real, imag} */,
  {32'h417de461, 32'h41d5c64f} /* (30, 18, 21) {real, imag} */,
  {32'h40cd082a, 32'hbf88d3c0} /* (30, 18, 20) {real, imag} */,
  {32'h40f15a48, 32'h3fa214f8} /* (30, 18, 19) {real, imag} */,
  {32'h410aabbc, 32'h408925b8} /* (30, 18, 18) {real, imag} */,
  {32'h41108258, 32'h411f102a} /* (30, 18, 17) {real, imag} */,
  {32'h40b77698, 32'hc1017d10} /* (30, 18, 16) {real, imag} */,
  {32'h40c15c00, 32'hc1400aba} /* (30, 18, 15) {real, imag} */,
  {32'hc0c93737, 32'hbf31b760} /* (30, 18, 14) {real, imag} */,
  {32'h411acfe8, 32'hc1abdf00} /* (30, 18, 13) {real, imag} */,
  {32'h41a1d6a8, 32'h409a8f90} /* (30, 18, 12) {real, imag} */,
  {32'h40a84b76, 32'h4126893a} /* (30, 18, 11) {real, imag} */,
  {32'hc13b8522, 32'h406f69d9} /* (30, 18, 10) {real, imag} */,
  {32'h4141b3fe, 32'h4100a0e2} /* (30, 18, 9) {real, imag} */,
  {32'h4083a498, 32'hc1a3313c} /* (30, 18, 8) {real, imag} */,
  {32'h3fddb050, 32'hc1d165dd} /* (30, 18, 7) {real, imag} */,
  {32'h42b231e0, 32'h411bb2a4} /* (30, 18, 6) {real, imag} */,
  {32'hc241a103, 32'hc0923ade} /* (30, 18, 5) {real, imag} */,
  {32'h424b4d3a, 32'hc15665b0} /* (30, 18, 4) {real, imag} */,
  {32'hc1fa3f1a, 32'h4245ef33} /* (30, 18, 3) {real, imag} */,
  {32'hc2cf0be4, 32'hc2309d06} /* (30, 18, 2) {real, imag} */,
  {32'h42ed5e2c, 32'h429de420} /* (30, 18, 1) {real, imag} */,
  {32'h42b8ee80, 32'hc16ab05a} /* (30, 18, 0) {real, imag} */,
  {32'hc28b13d8, 32'h42686974} /* (30, 17, 31) {real, imag} */,
  {32'h424e3094, 32'h422ded53} /* (30, 17, 30) {real, imag} */,
  {32'hc110e744, 32'hc20c909d} /* (30, 17, 29) {real, imag} */,
  {32'h424a6ea4, 32'h412c7503} /* (30, 17, 28) {real, imag} */,
  {32'hc0c4d4e2, 32'hc18c5fdf} /* (30, 17, 27) {real, imag} */,
  {32'hc2ad099e, 32'h40936fd2} /* (30, 17, 26) {real, imag} */,
  {32'h423a2378, 32'h41d861be} /* (30, 17, 25) {real, imag} */,
  {32'hc19cef42, 32'hc0d87504} /* (30, 17, 24) {real, imag} */,
  {32'h4153e97c, 32'h40ad8238} /* (30, 17, 23) {real, imag} */,
  {32'hbf7ddfa0, 32'h419a7406} /* (30, 17, 22) {real, imag} */,
  {32'h41674185, 32'hc16dc099} /* (30, 17, 21) {real, imag} */,
  {32'h419cac00, 32'hc076f37a} /* (30, 17, 20) {real, imag} */,
  {32'h4041344e, 32'h40baf1c8} /* (30, 17, 19) {real, imag} */,
  {32'hc0a266bf, 32'hc08fd91c} /* (30, 17, 18) {real, imag} */,
  {32'h410a6e46, 32'h40b992d4} /* (30, 17, 17) {real, imag} */,
  {32'hc02cbaa0, 32'h4091286b} /* (30, 17, 16) {real, imag} */,
  {32'h3fcbda30, 32'hc02c4b48} /* (30, 17, 15) {real, imag} */,
  {32'hc0916bbd, 32'hc04225d7} /* (30, 17, 14) {real, imag} */,
  {32'hc0a8be09, 32'h41186840} /* (30, 17, 13) {real, imag} */,
  {32'h40e76244, 32'h402cce56} /* (30, 17, 12) {real, imag} */,
  {32'h41336541, 32'hbffc9c38} /* (30, 17, 11) {real, imag} */,
  {32'h41af9a6d, 32'hc18f97ae} /* (30, 17, 10) {real, imag} */,
  {32'h41b6fad8, 32'hc1d95a70} /* (30, 17, 9) {real, imag} */,
  {32'h41879a94, 32'hc1269452} /* (30, 17, 8) {real, imag} */,
  {32'h401fbeb0, 32'hc10ab948} /* (30, 17, 7) {real, imag} */,
  {32'hc24d2cc7, 32'hc113145f} /* (30, 17, 6) {real, imag} */,
  {32'h41aa9ea2, 32'h41126878} /* (30, 17, 5) {real, imag} */,
  {32'hc0df42c0, 32'hc16e89d1} /* (30, 17, 4) {real, imag} */,
  {32'h41fa42b6, 32'hc2883d44} /* (30, 17, 3) {real, imag} */,
  {32'h41a3a000, 32'h42178ab5} /* (30, 17, 2) {real, imag} */,
  {32'hc1e19cca, 32'h42202236} /* (30, 17, 1) {real, imag} */,
  {32'hc231333e, 32'h4192da69} /* (30, 17, 0) {real, imag} */,
  {32'h3f9e5810, 32'hc18130c1} /* (30, 16, 31) {real, imag} */,
  {32'hc2076392, 32'h419de3d2} /* (30, 16, 30) {real, imag} */,
  {32'hc1cf7133, 32'hc19dbc54} /* (30, 16, 29) {real, imag} */,
  {32'h422bbcf2, 32'hc24741fe} /* (30, 16, 28) {real, imag} */,
  {32'h41eb2fb7, 32'hc0cbc738} /* (30, 16, 27) {real, imag} */,
  {32'h419dce61, 32'h416ad602} /* (30, 16, 26) {real, imag} */,
  {32'hc08f0be0, 32'h4004e262} /* (30, 16, 25) {real, imag} */,
  {32'hc0ea404e, 32'hc1858af1} /* (30, 16, 24) {real, imag} */,
  {32'h4133885d, 32'hc182e297} /* (30, 16, 23) {real, imag} */,
  {32'h41b94db1, 32'hc10198d4} /* (30, 16, 22) {real, imag} */,
  {32'hc14d2b06, 32'hc05605aa} /* (30, 16, 21) {real, imag} */,
  {32'hbee650c0, 32'h41555d4b} /* (30, 16, 20) {real, imag} */,
  {32'hc12a5e32, 32'h41c1c261} /* (30, 16, 19) {real, imag} */,
  {32'h3f95ae14, 32'hbfd9919c} /* (30, 16, 18) {real, imag} */,
  {32'hc139d611, 32'hc17d8d87} /* (30, 16, 17) {real, imag} */,
  {32'hc037c0c0, 32'hc0e494ad} /* (30, 16, 16) {real, imag} */,
  {32'hc08d928e, 32'hc0f72d5a} /* (30, 16, 15) {real, imag} */,
  {32'h410c6980, 32'hc0cbd145} /* (30, 16, 14) {real, imag} */,
  {32'hc11fb016, 32'h3f9a7120} /* (30, 16, 13) {real, imag} */,
  {32'hc08fda7c, 32'hc03d1a24} /* (30, 16, 12) {real, imag} */,
  {32'h4177ff2e, 32'hc132d880} /* (30, 16, 11) {real, imag} */,
  {32'hbf03c5e0, 32'hc21b2b71} /* (30, 16, 10) {real, imag} */,
  {32'h4144a3e1, 32'h40f0e445} /* (30, 16, 9) {real, imag} */,
  {32'h41efe47c, 32'h418c5e67} /* (30, 16, 8) {real, imag} */,
  {32'hc142ea0a, 32'hc1867e0a} /* (30, 16, 7) {real, imag} */,
  {32'hc21d8f6c, 32'hc12f8e7a} /* (30, 16, 6) {real, imag} */,
  {32'hc1a67f1f, 32'hc1da9012} /* (30, 16, 5) {real, imag} */,
  {32'h401aa1c0, 32'hc0d89d80} /* (30, 16, 4) {real, imag} */,
  {32'h41b78b31, 32'h408c2cc4} /* (30, 16, 3) {real, imag} */,
  {32'hc10c637a, 32'hbe944aa0} /* (30, 16, 2) {real, imag} */,
  {32'hc2334536, 32'h42268e82} /* (30, 16, 1) {real, imag} */,
  {32'hc2314a74, 32'h4192931c} /* (30, 16, 0) {real, imag} */,
  {32'h42d8b7bb, 32'h4208a035} /* (30, 15, 31) {real, imag} */,
  {32'hc2969dc8, 32'h40a64de6} /* (30, 15, 30) {real, imag} */,
  {32'h3f55eed0, 32'hc1ae4512} /* (30, 15, 29) {real, imag} */,
  {32'hc0a83a2e, 32'hc259a864} /* (30, 15, 28) {real, imag} */,
  {32'h41d506d2, 32'hbec4bc00} /* (30, 15, 27) {real, imag} */,
  {32'h41b499ad, 32'hc1c2db41} /* (30, 15, 26) {real, imag} */,
  {32'hc06d9d22, 32'h41a1f54d} /* (30, 15, 25) {real, imag} */,
  {32'h4183d676, 32'hc11eef2d} /* (30, 15, 24) {real, imag} */,
  {32'hc119a460, 32'h40c3a456} /* (30, 15, 23) {real, imag} */,
  {32'h41aaa4a6, 32'h40bd627a} /* (30, 15, 22) {real, imag} */,
  {32'hc0c64fd5, 32'hc10e91ee} /* (30, 15, 21) {real, imag} */,
  {32'hc043176c, 32'hbf751ce0} /* (30, 15, 20) {real, imag} */,
  {32'hc037e660, 32'hbfcf16d0} /* (30, 15, 19) {real, imag} */,
  {32'h404cf680, 32'h41953856} /* (30, 15, 18) {real, imag} */,
  {32'hc0e5b774, 32'hc1877c16} /* (30, 15, 17) {real, imag} */,
  {32'h40041880, 32'h412855ce} /* (30, 15, 16) {real, imag} */,
  {32'hc1077516, 32'h3ecd0760} /* (30, 15, 15) {real, imag} */,
  {32'hc1c0e9ca, 32'hc0c40ba4} /* (30, 15, 14) {real, imag} */,
  {32'h3fb63008, 32'hbf03d4a0} /* (30, 15, 13) {real, imag} */,
  {32'hc0ce7006, 32'h41921c9b} /* (30, 15, 12) {real, imag} */,
  {32'h4082ebeb, 32'hc1a2fd2f} /* (30, 15, 11) {real, imag} */,
  {32'h4196a946, 32'h4188e540} /* (30, 15, 10) {real, imag} */,
  {32'h41b616d6, 32'hc020d5dc} /* (30, 15, 9) {real, imag} */,
  {32'hc164169c, 32'hc16ec949} /* (30, 15, 8) {real, imag} */,
  {32'h3d6dd380, 32'hc24dc8c6} /* (30, 15, 7) {real, imag} */,
  {32'h4201d340, 32'h420abd32} /* (30, 15, 6) {real, imag} */,
  {32'hc16c4280, 32'hc1b40e34} /* (30, 15, 5) {real, imag} */,
  {32'h4202c30a, 32'h4243aa60} /* (30, 15, 4) {real, imag} */,
  {32'hc11ab296, 32'h403e9374} /* (30, 15, 3) {real, imag} */,
  {32'hc27f8f5f, 32'hc16a21e7} /* (30, 15, 2) {real, imag} */,
  {32'h4245332e, 32'hc1e047ba} /* (30, 15, 1) {real, imag} */,
  {32'h429e1a9c, 32'h422872dc} /* (30, 15, 0) {real, imag} */,
  {32'hc2cd7b7e, 32'h42eabfd3} /* (30, 14, 31) {real, imag} */,
  {32'h42198180, 32'hc2a04db1} /* (30, 14, 30) {real, imag} */,
  {32'h423d1730, 32'h41d9de6e} /* (30, 14, 29) {real, imag} */,
  {32'hc2900790, 32'h42f746ce} /* (30, 14, 28) {real, imag} */,
  {32'hc0896a54, 32'hc211a8ed} /* (30, 14, 27) {real, imag} */,
  {32'h41a51003, 32'hc1aa4b07} /* (30, 14, 26) {real, imag} */,
  {32'hc175f5c2, 32'hbfa0016c} /* (30, 14, 25) {real, imag} */,
  {32'h41ca4710, 32'hc259325e} /* (30, 14, 24) {real, imag} */,
  {32'h3fdda870, 32'h41506888} /* (30, 14, 23) {real, imag} */,
  {32'h409f489c, 32'hc12d9404} /* (30, 14, 22) {real, imag} */,
  {32'hbed7f310, 32'hc0b868f9} /* (30, 14, 21) {real, imag} */,
  {32'hc12bd637, 32'h3fcf9010} /* (30, 14, 20) {real, imag} */,
  {32'h413fa720, 32'h417fbf85} /* (30, 14, 19) {real, imag} */,
  {32'h4136a9ba, 32'h40420b1c} /* (30, 14, 18) {real, imag} */,
  {32'h40b6b285, 32'hc0ff774c} /* (30, 14, 17) {real, imag} */,
  {32'hc146f328, 32'hc0277508} /* (30, 14, 16) {real, imag} */,
  {32'hbfac7a54, 32'h40ed19d4} /* (30, 14, 15) {real, imag} */,
  {32'h411525c0, 32'hc10ca1ad} /* (30, 14, 14) {real, imag} */,
  {32'hc18d1994, 32'hbf1d4970} /* (30, 14, 13) {real, imag} */,
  {32'h4180b1be, 32'h41632266} /* (30, 14, 12) {real, imag} */,
  {32'h4145b670, 32'h405ef24e} /* (30, 14, 11) {real, imag} */,
  {32'hc16209c6, 32'hc1f479ba} /* (30, 14, 10) {real, imag} */,
  {32'h401de938, 32'hc20a4cba} /* (30, 14, 9) {real, imag} */,
  {32'h41822b3c, 32'hc11f6dd0} /* (30, 14, 8) {real, imag} */,
  {32'h419ab10b, 32'hc0a0bd0b} /* (30, 14, 7) {real, imag} */,
  {32'h4234eb86, 32'hc19b0419} /* (30, 14, 6) {real, imag} */,
  {32'h41f5e5bd, 32'h420eee69} /* (30, 14, 5) {real, imag} */,
  {32'h3f204700, 32'h420764cc} /* (30, 14, 4) {real, imag} */,
  {32'h41871741, 32'hc06e0244} /* (30, 14, 3) {real, imag} */,
  {32'h414058ae, 32'h41ee52e4} /* (30, 14, 2) {real, imag} */,
  {32'hc2936cda, 32'hc215fa9e} /* (30, 14, 1) {real, imag} */,
  {32'hc2a77c88, 32'hc228e8aa} /* (30, 14, 0) {real, imag} */,
  {32'h416edcd8, 32'hc1be4fd0} /* (30, 13, 31) {real, imag} */,
  {32'h3e912b90, 32'hc15aeada} /* (30, 13, 30) {real, imag} */,
  {32'hc1d56011, 32'hc0e8b270} /* (30, 13, 29) {real, imag} */,
  {32'h41e08c9e, 32'hc2954a4e} /* (30, 13, 28) {real, imag} */,
  {32'h411176f5, 32'hc24d6826} /* (30, 13, 27) {real, imag} */,
  {32'hc28fcadc, 32'hc294cd69} /* (30, 13, 26) {real, imag} */,
  {32'hc21337bd, 32'hbf92ce80} /* (30, 13, 25) {real, imag} */,
  {32'hc176a6f8, 32'h418d64d5} /* (30, 13, 24) {real, imag} */,
  {32'h41a40452, 32'hc182777f} /* (30, 13, 23) {real, imag} */,
  {32'h41282283, 32'hc1ecb167} /* (30, 13, 22) {real, imag} */,
  {32'h3dc54cc0, 32'h416c31d6} /* (30, 13, 21) {real, imag} */,
  {32'h41a7ac6c, 32'hbfa927fc} /* (30, 13, 20) {real, imag} */,
  {32'h3f8cc4a4, 32'h4018e2be} /* (30, 13, 19) {real, imag} */,
  {32'h418e1739, 32'h413f5a68} /* (30, 13, 18) {real, imag} */,
  {32'hbfa035e8, 32'h40d37944} /* (30, 13, 17) {real, imag} */,
  {32'h41919657, 32'hbc12c000} /* (30, 13, 16) {real, imag} */,
  {32'h40edcf4a, 32'hc017d888} /* (30, 13, 15) {real, imag} */,
  {32'hc101dde6, 32'hc1cf9884} /* (30, 13, 14) {real, imag} */,
  {32'h4006fafe, 32'hc0c5ac1d} /* (30, 13, 13) {real, imag} */,
  {32'hc1864210, 32'hc11dadd4} /* (30, 13, 12) {real, imag} */,
  {32'hc120c750, 32'h40ddda3c} /* (30, 13, 11) {real, imag} */,
  {32'hc10265eb, 32'h3f184260} /* (30, 13, 10) {real, imag} */,
  {32'h419c0716, 32'h4165da26} /* (30, 13, 9) {real, imag} */,
  {32'hc2043d48, 32'h40dab934} /* (30, 13, 8) {real, imag} */,
  {32'hc1ade94e, 32'hc2916be0} /* (30, 13, 7) {real, imag} */,
  {32'hc1cbf1b2, 32'h4220b54a} /* (30, 13, 6) {real, imag} */,
  {32'hc173cf1b, 32'h4242feb0} /* (30, 13, 5) {real, imag} */,
  {32'h41f93d06, 32'hc25e2a38} /* (30, 13, 4) {real, imag} */,
  {32'hc166517e, 32'h413fa0da} /* (30, 13, 3) {real, imag} */,
  {32'hc09dc0d1, 32'h41d03f37} /* (30, 13, 2) {real, imag} */,
  {32'h42852174, 32'hc2e13528} /* (30, 13, 1) {real, imag} */,
  {32'h4283b25b, 32'hc1b4f546} /* (30, 13, 0) {real, imag} */,
  {32'h429e6c41, 32'h41a1a41b} /* (30, 12, 31) {real, imag} */,
  {32'h4266d1a6, 32'hc0a5cf8a} /* (30, 12, 30) {real, imag} */,
  {32'hc029a338, 32'h416139e8} /* (30, 12, 29) {real, imag} */,
  {32'hc15346e7, 32'hc11ac8f0} /* (30, 12, 28) {real, imag} */,
  {32'h418f1630, 32'h42179563} /* (30, 12, 27) {real, imag} */,
  {32'hc1e182d4, 32'hc1e744bd} /* (30, 12, 26) {real, imag} */,
  {32'hc044c48c, 32'hc0198a20} /* (30, 12, 25) {real, imag} */,
  {32'h42226ba8, 32'h41a238c8} /* (30, 12, 24) {real, imag} */,
  {32'hc23b9a10, 32'h41e64ff6} /* (30, 12, 23) {real, imag} */,
  {32'hc129badf, 32'hc12c0cd8} /* (30, 12, 22) {real, imag} */,
  {32'h3f8957c8, 32'h401cae78} /* (30, 12, 21) {real, imag} */,
  {32'h4105b682, 32'h4209bc0b} /* (30, 12, 20) {real, imag} */,
  {32'h411abc1b, 32'hc05fb568} /* (30, 12, 19) {real, imag} */,
  {32'hc0706066, 32'h4184bdc0} /* (30, 12, 18) {real, imag} */,
  {32'hc1a9709e, 32'h41223beb} /* (30, 12, 17) {real, imag} */,
  {32'hc042deb8, 32'h3f052280} /* (30, 12, 16) {real, imag} */,
  {32'h3fd2e160, 32'hc00af3c4} /* (30, 12, 15) {real, imag} */,
  {32'hc0ac70eb, 32'h41d7f7ac} /* (30, 12, 14) {real, imag} */,
  {32'hc18e2508, 32'hc18972b7} /* (30, 12, 13) {real, imag} */,
  {32'hc1cee3a3, 32'h4149987c} /* (30, 12, 12) {real, imag} */,
  {32'h41468e33, 32'hc17bdaa6} /* (30, 12, 11) {real, imag} */,
  {32'h41580539, 32'hc214cb81} /* (30, 12, 10) {real, imag} */,
  {32'hc112c2d6, 32'h42ac6ac2} /* (30, 12, 9) {real, imag} */,
  {32'h411eb543, 32'hc14ede7c} /* (30, 12, 8) {real, imag} */,
  {32'hc1b844b6, 32'h41572328} /* (30, 12, 7) {real, imag} */,
  {32'h40058e7c, 32'hc259df1e} /* (30, 12, 6) {real, imag} */,
  {32'h3f9b2a58, 32'hc2017c31} /* (30, 12, 5) {real, imag} */,
  {32'hc1f2b55e, 32'hc212961c} /* (30, 12, 4) {real, imag} */,
  {32'h424e30c0, 32'hc226b801} /* (30, 12, 3) {real, imag} */,
  {32'hc240137a, 32'hc0b48c66} /* (30, 12, 2) {real, imag} */,
  {32'h41d62370, 32'h41ba7dc9} /* (30, 12, 1) {real, imag} */,
  {32'hc27a99f8, 32'hc299642f} /* (30, 12, 0) {real, imag} */,
  {32'hc337664b, 32'h4356faf2} /* (30, 11, 31) {real, imag} */,
  {32'h427b62cc, 32'hc2565ff9} /* (30, 11, 30) {real, imag} */,
  {32'hc22009f9, 32'hc2d2d85d} /* (30, 11, 29) {real, imag} */,
  {32'h42a62c8b, 32'h3f7b5de0} /* (30, 11, 28) {real, imag} */,
  {32'h426a9e68, 32'hc2931dde} /* (30, 11, 27) {real, imag} */,
  {32'h41d95e28, 32'h42849fb6} /* (30, 11, 26) {real, imag} */,
  {32'hc1f734af, 32'hc16060ba} /* (30, 11, 25) {real, imag} */,
  {32'hc032d8e0, 32'hc290e87e} /* (30, 11, 24) {real, imag} */,
  {32'h41630ade, 32'hc1b0570f} /* (30, 11, 23) {real, imag} */,
  {32'h41c8f378, 32'h41a618fa} /* (30, 11, 22) {real, imag} */,
  {32'h41426aaa, 32'hc23d529e} /* (30, 11, 21) {real, imag} */,
  {32'hc168fe80, 32'h4195082a} /* (30, 11, 20) {real, imag} */,
  {32'hc0fa2496, 32'hc04118c4} /* (30, 11, 19) {real, imag} */,
  {32'h402daac8, 32'hc0169d84} /* (30, 11, 18) {real, imag} */,
  {32'h41cca3a8, 32'h409bd22c} /* (30, 11, 17) {real, imag} */,
  {32'hc1eedc6a, 32'h41791388} /* (30, 11, 16) {real, imag} */,
  {32'hc0520d40, 32'hc08332cc} /* (30, 11, 15) {real, imag} */,
  {32'hc0ddc4f4, 32'h4120ba79} /* (30, 11, 14) {real, imag} */,
  {32'h41391205, 32'h3f151410} /* (30, 11, 13) {real, imag} */,
  {32'hc233fed2, 32'hbdf79380} /* (30, 11, 12) {real, imag} */,
  {32'h41d0bc03, 32'hc1d12ecb} /* (30, 11, 11) {real, imag} */,
  {32'h42519d12, 32'hc2bbb0d4} /* (30, 11, 10) {real, imag} */,
  {32'hc1cf93db, 32'hc208396a} /* (30, 11, 9) {real, imag} */,
  {32'h42896e33, 32'hc0b4d2f0} /* (30, 11, 8) {real, imag} */,
  {32'hc11f140a, 32'hc2386918} /* (30, 11, 7) {real, imag} */,
  {32'h4220c4ce, 32'h4244c9ef} /* (30, 11, 6) {real, imag} */,
  {32'h42d6ce88, 32'hc248f7a9} /* (30, 11, 5) {real, imag} */,
  {32'hc2124734, 32'hc2150820} /* (30, 11, 4) {real, imag} */,
  {32'hc18e8312, 32'hc26bfa12} /* (30, 11, 3) {real, imag} */,
  {32'h4319306d, 32'hc1b24cba} /* (30, 11, 2) {real, imag} */,
  {32'hc37ec771, 32'h430da39e} /* (30, 11, 1) {real, imag} */,
  {32'hc2e75818, 32'h437c5288} /* (30, 11, 0) {real, imag} */,
  {32'h434faa34, 32'h427ca70c} /* (30, 10, 31) {real, imag} */,
  {32'hc19e5354, 32'hc28a12b2} /* (30, 10, 30) {real, imag} */,
  {32'h42a4ca0b, 32'hc227fb86} /* (30, 10, 29) {real, imag} */,
  {32'hc23568ae, 32'hc155ab3a} /* (30, 10, 28) {real, imag} */,
  {32'hc18f940c, 32'h42b27dfe} /* (30, 10, 27) {real, imag} */,
  {32'hc17247a5, 32'h4266b4ff} /* (30, 10, 26) {real, imag} */,
  {32'h4235fd8e, 32'h4242482a} /* (30, 10, 25) {real, imag} */,
  {32'hc1d0fd6b, 32'h42727656} /* (30, 10, 24) {real, imag} */,
  {32'h3fdde7e0, 32'h3faa0c00} /* (30, 10, 23) {real, imag} */,
  {32'hc1bb6622, 32'hc1e0f066} /* (30, 10, 22) {real, imag} */,
  {32'hc258beb4, 32'hc1c6c376} /* (30, 10, 21) {real, imag} */,
  {32'hc1080a50, 32'h408e4ea5} /* (30, 10, 20) {real, imag} */,
  {32'h41f8c024, 32'hc0e8b832} /* (30, 10, 19) {real, imag} */,
  {32'h41b16540, 32'hc14af992} /* (30, 10, 18) {real, imag} */,
  {32'h41304c20, 32'hc1a27551} /* (30, 10, 17) {real, imag} */,
  {32'h41b7dceb, 32'h41d5859f} /* (30, 10, 16) {real, imag} */,
  {32'h40c40ea0, 32'h410f308e} /* (30, 10, 15) {real, imag} */,
  {32'hc1b3c318, 32'hc0ab4514} /* (30, 10, 14) {real, imag} */,
  {32'hc17fcb80, 32'hc1ecd942} /* (30, 10, 13) {real, imag} */,
  {32'hc2080f6d, 32'h41575e80} /* (30, 10, 12) {real, imag} */,
  {32'h416ea898, 32'h41fb4316} /* (30, 10, 11) {real, imag} */,
  {32'h421c3f11, 32'h4203d51d} /* (30, 10, 10) {real, imag} */,
  {32'hbfa6c240, 32'hc21d8bec} /* (30, 10, 9) {real, imag} */,
  {32'hc24d0a5a, 32'h41ffae8f} /* (30, 10, 8) {real, imag} */,
  {32'hc1b9911d, 32'hc17d8608} /* (30, 10, 7) {real, imag} */,
  {32'hc0fe8f1a, 32'hc2cee914} /* (30, 10, 6) {real, imag} */,
  {32'hc11d1f29, 32'hc282f3ca} /* (30, 10, 5) {real, imag} */,
  {32'h428fcb8b, 32'hc25086ec} /* (30, 10, 4) {real, imag} */,
  {32'h4204d820, 32'hc1eb3554} /* (30, 10, 3) {real, imag} */,
  {32'hc2b6092d, 32'h432dc03f} /* (30, 10, 2) {real, imag} */,
  {32'h428bfc50, 32'hc3192d8e} /* (30, 10, 1) {real, imag} */,
  {32'h428a570d, 32'hc13ebb66} /* (30, 10, 0) {real, imag} */,
  {32'h42a5c1ce, 32'h433e0d4f} /* (30, 9, 31) {real, imag} */,
  {32'hc348f286, 32'h4202ccce} /* (30, 9, 30) {real, imag} */,
  {32'h42a9d896, 32'hc09676bc} /* (30, 9, 29) {real, imag} */,
  {32'h4248504a, 32'hc27e38a7} /* (30, 9, 28) {real, imag} */,
  {32'hc23003e5, 32'h40db97c4} /* (30, 9, 27) {real, imag} */,
  {32'h42c49fbe, 32'h425751aa} /* (30, 9, 26) {real, imag} */,
  {32'h41a8918c, 32'hc196a786} /* (30, 9, 25) {real, imag} */,
  {32'hc1d87504, 32'h41ef0aff} /* (30, 9, 24) {real, imag} */,
  {32'h421f2a15, 32'hc1f1d3fc} /* (30, 9, 23) {real, imag} */,
  {32'hc220cbe4, 32'h429713d2} /* (30, 9, 22) {real, imag} */,
  {32'h41d18cd2, 32'h424118a4} /* (30, 9, 21) {real, imag} */,
  {32'hc2531de0, 32'hc229bd88} /* (30, 9, 20) {real, imag} */,
  {32'hc14cdf2c, 32'hc261574e} /* (30, 9, 19) {real, imag} */,
  {32'h414e6516, 32'hc204d180} /* (30, 9, 18) {real, imag} */,
  {32'h41a7e769, 32'hc0bc1703} /* (30, 9, 17) {real, imag} */,
  {32'h41cf1294, 32'h41114541} /* (30, 9, 16) {real, imag} */,
  {32'hc1978bf9, 32'h417a209e} /* (30, 9, 15) {real, imag} */,
  {32'hc105f056, 32'hc1bcd1c0} /* (30, 9, 14) {real, imag} */,
  {32'h42172379, 32'h421467e4} /* (30, 9, 13) {real, imag} */,
  {32'hc0f55a40, 32'hc1779a9a} /* (30, 9, 12) {real, imag} */,
  {32'hc2526777, 32'hc0713f78} /* (30, 9, 11) {real, imag} */,
  {32'hc1b291ab, 32'h428198ce} /* (30, 9, 10) {real, imag} */,
  {32'h42162f83, 32'hc1a86cda} /* (30, 9, 9) {real, imag} */,
  {32'hc2f2c975, 32'h4182410d} /* (30, 9, 8) {real, imag} */,
  {32'h4207d026, 32'hbfd47a40} /* (30, 9, 7) {real, imag} */,
  {32'h417b3df4, 32'hc23c593c} /* (30, 9, 6) {real, imag} */,
  {32'h42a42bba, 32'hc2836dae} /* (30, 9, 5) {real, imag} */,
  {32'h431b6ff6, 32'h4105b984} /* (30, 9, 4) {real, imag} */,
  {32'hc350f001, 32'h425e35ca} /* (30, 9, 3) {real, imag} */,
  {32'hc3266e86, 32'h412b2ce8} /* (30, 9, 2) {real, imag} */,
  {32'h43402ff3, 32'hc3398617} /* (30, 9, 1) {real, imag} */,
  {32'h41e289de, 32'hbdfce180} /* (30, 9, 0) {real, imag} */,
  {32'hc3adac72, 32'h443359a1} /* (30, 8, 31) {real, imag} */,
  {32'hc2a8daf2, 32'hc3b09143} /* (30, 8, 30) {real, imag} */,
  {32'hc3173aea, 32'hc20fb1c7} /* (30, 8, 29) {real, imag} */,
  {32'hc27457e3, 32'h41dafaa8} /* (30, 8, 28) {real, imag} */,
  {32'h42916811, 32'hc2654c6e} /* (30, 8, 27) {real, imag} */,
  {32'h402d6048, 32'h42dbba0d} /* (30, 8, 26) {real, imag} */,
  {32'hc2d5479e, 32'h422af68c} /* (30, 8, 25) {real, imag} */,
  {32'hc22042e1, 32'hc207c3c1} /* (30, 8, 24) {real, imag} */,
  {32'hbf0e9e30, 32'h428c7a80} /* (30, 8, 23) {real, imag} */,
  {32'h3e193600, 32'hc30b2cdc} /* (30, 8, 22) {real, imag} */,
  {32'hc15c77f8, 32'hc28ab257} /* (30, 8, 21) {real, imag} */,
  {32'hbf6fb240, 32'hc23f5f1c} /* (30, 8, 20) {real, imag} */,
  {32'h415ebbec, 32'hbeb65e00} /* (30, 8, 19) {real, imag} */,
  {32'h4164f979, 32'hbfc24240} /* (30, 8, 18) {real, imag} */,
  {32'h41e0f3a5, 32'hc14ee5a8} /* (30, 8, 17) {real, imag} */,
  {32'hc145a060, 32'h4020f100} /* (30, 8, 16) {real, imag} */,
  {32'hc0c43f54, 32'h4013cfa0} /* (30, 8, 15) {real, imag} */,
  {32'h40935fd2, 32'h3e328a00} /* (30, 8, 14) {real, imag} */,
  {32'h41725f5c, 32'h40525830} /* (30, 8, 13) {real, imag} */,
  {32'h41fdf99e, 32'h41aa7214} /* (30, 8, 12) {real, imag} */,
  {32'h4218a4ae, 32'hc1f05804} /* (30, 8, 11) {real, imag} */,
  {32'hc293459f, 32'hbeaced00} /* (30, 8, 10) {real, imag} */,
  {32'hc148a6a5, 32'h3ff7dee0} /* (30, 8, 9) {real, imag} */,
  {32'h4256f98b, 32'hc25e71c3} /* (30, 8, 8) {real, imag} */,
  {32'hc2aa0286, 32'hc1caab05} /* (30, 8, 7) {real, imag} */,
  {32'h4212a4b4, 32'hc2ab2067} /* (30, 8, 6) {real, imag} */,
  {32'h4332a462, 32'hc30ae316} /* (30, 8, 5) {real, imag} */,
  {32'hc26726cb, 32'h432a4501} /* (30, 8, 4) {real, imag} */,
  {32'h41a9e904, 32'h416add20} /* (30, 8, 3) {real, imag} */,
  {32'h42e7b864, 32'hc32540ea} /* (30, 8, 2) {real, imag} */,
  {32'hc361340c, 32'h43af5316} /* (30, 8, 1) {real, imag} */,
  {32'hc27c6876, 32'h43b86c38} /* (30, 8, 0) {real, imag} */,
  {32'h42fa430e, 32'hc2bd8edc} /* (30, 7, 31) {real, imag} */,
  {32'hc20f083d, 32'h4202339a} /* (30, 7, 30) {real, imag} */,
  {32'hc1935713, 32'hc24247da} /* (30, 7, 29) {real, imag} */,
  {32'hc22a150e, 32'h42b7d37b} /* (30, 7, 28) {real, imag} */,
  {32'h41c185d8, 32'h41f29f7e} /* (30, 7, 27) {real, imag} */,
  {32'h422f275c, 32'hc1955306} /* (30, 7, 26) {real, imag} */,
  {32'hc0fa38e6, 32'hc22d3d58} /* (30, 7, 25) {real, imag} */,
  {32'hc214511c, 32'h42968686} /* (30, 7, 24) {real, imag} */,
  {32'hc248cda5, 32'h41f5b2b7} /* (30, 7, 23) {real, imag} */,
  {32'h41ec98f6, 32'hc20313f4} /* (30, 7, 22) {real, imag} */,
  {32'hc0cdb394, 32'h40dfcd3c} /* (30, 7, 21) {real, imag} */,
  {32'hc10efc10, 32'hc18f10c3} /* (30, 7, 20) {real, imag} */,
  {32'h42024f1e, 32'hc2cf2e90} /* (30, 7, 19) {real, imag} */,
  {32'h41b6ff48, 32'h42491d60} /* (30, 7, 18) {real, imag} */,
  {32'hc18025dc, 32'h422601c8} /* (30, 7, 17) {real, imag} */,
  {32'h427ddeaa, 32'h420601bf} /* (30, 7, 16) {real, imag} */,
  {32'hc1135e08, 32'hc1b9ec84} /* (30, 7, 15) {real, imag} */,
  {32'h411d9759, 32'hc1a08ad0} /* (30, 7, 14) {real, imag} */,
  {32'hc2447e66, 32'hc0620b70} /* (30, 7, 13) {real, imag} */,
  {32'h413d4598, 32'h409ae8dc} /* (30, 7, 12) {real, imag} */,
  {32'h4087179c, 32'hc2348296} /* (30, 7, 11) {real, imag} */,
  {32'h40d32048, 32'h42253a7a} /* (30, 7, 10) {real, imag} */,
  {32'hc275dbf1, 32'h419c3e0f} /* (30, 7, 9) {real, imag} */,
  {32'hc2839ef4, 32'hc293757c} /* (30, 7, 8) {real, imag} */,
  {32'hc1a6753a, 32'hc099a804} /* (30, 7, 7) {real, imag} */,
  {32'hc3091135, 32'hc24048a9} /* (30, 7, 6) {real, imag} */,
  {32'hc2f13c02, 32'h42bee870} /* (30, 7, 5) {real, imag} */,
  {32'hc0f19b70, 32'h425ab0ea} /* (30, 7, 4) {real, imag} */,
  {32'hc1faec9b, 32'hc2a42d6b} /* (30, 7, 3) {real, imag} */,
  {32'hc24876a5, 32'hc0e384d0} /* (30, 7, 2) {real, imag} */,
  {32'h436f5f45, 32'hc2f9ba94} /* (30, 7, 1) {real, imag} */,
  {32'h434c8c52, 32'hc2c257c0} /* (30, 7, 0) {real, imag} */,
  {32'hc2f1fd13, 32'h4312a7d0} /* (30, 6, 31) {real, imag} */,
  {32'hc12cebbe, 32'hc2b8c494} /* (30, 6, 30) {real, imag} */,
  {32'hc20987f5, 32'hc2e1909e} /* (30, 6, 29) {real, imag} */,
  {32'hc35b0684, 32'h41cdde0a} /* (30, 6, 28) {real, imag} */,
  {32'h40a30c48, 32'hc2473f44} /* (30, 6, 27) {real, imag} */,
  {32'h433ffe4d, 32'hc29069ef} /* (30, 6, 26) {real, imag} */,
  {32'h41415fea, 32'hc1d2075b} /* (30, 6, 25) {real, imag} */,
  {32'h42b24902, 32'hc1e92cf6} /* (30, 6, 24) {real, imag} */,
  {32'hc195a43c, 32'hc2d9de23} /* (30, 6, 23) {real, imag} */,
  {32'h419677dc, 32'hc1746fa2} /* (30, 6, 22) {real, imag} */,
  {32'h41fe3364, 32'hc25dd87f} /* (30, 6, 21) {real, imag} */,
  {32'hc2132704, 32'h42177e49} /* (30, 6, 20) {real, imag} */,
  {32'hc1502b44, 32'hc21b272d} /* (30, 6, 19) {real, imag} */,
  {32'hbf5d3ab0, 32'hc20cc0e1} /* (30, 6, 18) {real, imag} */,
  {32'h419fe181, 32'hc1672778} /* (30, 6, 17) {real, imag} */,
  {32'h424725c8, 32'h41666cc6} /* (30, 6, 16) {real, imag} */,
  {32'hc1aee871, 32'hc14c7b80} /* (30, 6, 15) {real, imag} */,
  {32'hc19e8340, 32'hc116e484} /* (30, 6, 14) {real, imag} */,
  {32'h416102dc, 32'hc1b04966} /* (30, 6, 13) {real, imag} */,
  {32'h41cff8f1, 32'hc044d490} /* (30, 6, 12) {real, imag} */,
  {32'h41c2b8a8, 32'hc252ba5b} /* (30, 6, 11) {real, imag} */,
  {32'hc1dda1d8, 32'h4116cdc2} /* (30, 6, 10) {real, imag} */,
  {32'hc295bed5, 32'h427aa33a} /* (30, 6, 9) {real, imag} */,
  {32'hc2116c64, 32'hc2af178a} /* (30, 6, 8) {real, imag} */,
  {32'h41ed6965, 32'hc172c4f6} /* (30, 6, 7) {real, imag} */,
  {32'hc24f8864, 32'hbfb97c40} /* (30, 6, 6) {real, imag} */,
  {32'hc26ee071, 32'hc325f949} /* (30, 6, 5) {real, imag} */,
  {32'hc2840037, 32'h4285a730} /* (30, 6, 4) {real, imag} */,
  {32'h42fd0614, 32'h42547d8c} /* (30, 6, 3) {real, imag} */,
  {32'h424c1c4e, 32'hc32332a8} /* (30, 6, 2) {real, imag} */,
  {32'hc2049112, 32'h418215a0} /* (30, 6, 1) {real, imag} */,
  {32'h42474ea4, 32'hc25e7f2a} /* (30, 6, 0) {real, imag} */,
  {32'hc1d5a9a0, 32'h446606d8} /* (30, 5, 31) {real, imag} */,
  {32'hc30643fa, 32'hc3942bea} /* (30, 5, 30) {real, imag} */,
  {32'hc2b0f36e, 32'h427d6582} /* (30, 5, 29) {real, imag} */,
  {32'h4375339a, 32'h41f20a46} /* (30, 5, 28) {real, imag} */,
  {32'h434db3ea, 32'hc35e4b48} /* (30, 5, 27) {real, imag} */,
  {32'hc2ba3fe0, 32'hc29e51e2} /* (30, 5, 26) {real, imag} */,
  {32'hc2aaad71, 32'h42b666a4} /* (30, 5, 25) {real, imag} */,
  {32'hc2d56597, 32'hc22e74b2} /* (30, 5, 24) {real, imag} */,
  {32'h41601158, 32'h40185800} /* (30, 5, 23) {real, imag} */,
  {32'hc182a872, 32'hc3199ff4} /* (30, 5, 22) {real, imag} */,
  {32'hc2b563e2, 32'hc1da194a} /* (30, 5, 21) {real, imag} */,
  {32'hc191c01e, 32'hc1847e2e} /* (30, 5, 20) {real, imag} */,
  {32'h41ce867a, 32'hc22f5cfb} /* (30, 5, 19) {real, imag} */,
  {32'hc21087de, 32'h4200e9dd} /* (30, 5, 18) {real, imag} */,
  {32'hc10b2960, 32'h4082c438} /* (30, 5, 17) {real, imag} */,
  {32'hc2643512, 32'h41c21e70} /* (30, 5, 16) {real, imag} */,
  {32'h42424610, 32'hc090c038} /* (30, 5, 15) {real, imag} */,
  {32'h427ca22e, 32'h41901886} /* (30, 5, 14) {real, imag} */,
  {32'h4218609f, 32'h42356125} /* (30, 5, 13) {real, imag} */,
  {32'h41f2074a, 32'hc1dcde56} /* (30, 5, 12) {real, imag} */,
  {32'h42c33362, 32'h41d034f2} /* (30, 5, 11) {real, imag} */,
  {32'hc1d39fd6, 32'h41804570} /* (30, 5, 10) {real, imag} */,
  {32'h421342ce, 32'hc190a70c} /* (30, 5, 9) {real, imag} */,
  {32'h4154f618, 32'h4286b4dd} /* (30, 5, 8) {real, imag} */,
  {32'hc240ba0a, 32'h427752bf} /* (30, 5, 7) {real, imag} */,
  {32'h42cba9b0, 32'hc2609924} /* (30, 5, 6) {real, imag} */,
  {32'hc1b1b1c0, 32'hc358fed4} /* (30, 5, 5) {real, imag} */,
  {32'hc29caacc, 32'hc242db99} /* (30, 5, 4) {real, imag} */,
  {32'hc2c96c14, 32'h42dd4f9f} /* (30, 5, 3) {real, imag} */,
  {32'h4365869a, 32'hc356c668} /* (30, 5, 2) {real, imag} */,
  {32'hc4270033, 32'h44410574} /* (30, 5, 1) {real, imag} */,
  {32'hc3258e78, 32'h441f9ef6} /* (30, 5, 0) {real, imag} */,
  {32'h441a08e0, 32'hc3fddd74} /* (30, 4, 31) {real, imag} */,
  {32'hc401cb0d, 32'h44280d93} /* (30, 4, 30) {real, imag} */,
  {32'hc1af5a6a, 32'h41f39108} /* (30, 4, 29) {real, imag} */,
  {32'h4229d978, 32'hc370ce9c} /* (30, 4, 28) {real, imag} */,
  {32'h42c443d0, 32'h439627c9} /* (30, 4, 27) {real, imag} */,
  {32'h431df7ef, 32'hc20878b5} /* (30, 4, 26) {real, imag} */,
  {32'hc25711ee, 32'h4074e910} /* (30, 4, 25) {real, imag} */,
  {32'hc2293fc4, 32'h425f7698} /* (30, 4, 24) {real, imag} */,
  {32'hc3017fec, 32'hc2507801} /* (30, 4, 23) {real, imag} */,
  {32'hc220723c, 32'hc171a05c} /* (30, 4, 22) {real, imag} */,
  {32'h42d02030, 32'h430049b4} /* (30, 4, 21) {real, imag} */,
  {32'hc2d6df8c, 32'hc2a31e0c} /* (30, 4, 20) {real, imag} */,
  {32'hc155b052, 32'hc18c3480} /* (30, 4, 19) {real, imag} */,
  {32'hbffdb2e0, 32'h42a729c9} /* (30, 4, 18) {real, imag} */,
  {32'hc15e0c08, 32'hc2501f30} /* (30, 4, 17) {real, imag} */,
  {32'hc0bf27cc, 32'hc21a8148} /* (30, 4, 16) {real, imag} */,
  {32'h427f1042, 32'h41aac720} /* (30, 4, 15) {real, imag} */,
  {32'hc2b0e644, 32'h4202989e} /* (30, 4, 14) {real, imag} */,
  {32'h410048fa, 32'h405dedc0} /* (30, 4, 13) {real, imag} */,
  {32'h412c6b20, 32'hc22f2003} /* (30, 4, 12) {real, imag} */,
  {32'hc2141ca9, 32'hc1695b28} /* (30, 4, 11) {real, imag} */,
  {32'h43096fe9, 32'h42520a3b} /* (30, 4, 10) {real, imag} */,
  {32'h427ab29a, 32'h4213988b} /* (30, 4, 9) {real, imag} */,
  {32'hc2eeb37e, 32'h4321debf} /* (30, 4, 8) {real, imag} */,
  {32'h427c0ff6, 32'hc2b17366} /* (30, 4, 7) {real, imag} */,
  {32'h4161ad30, 32'h41f1f322} /* (30, 4, 6) {real, imag} */,
  {32'hc3949ecf, 32'h42851b33} /* (30, 4, 5) {real, imag} */,
  {32'h41abbfb1, 32'h428d0c11} /* (30, 4, 4) {real, imag} */,
  {32'h426e939f, 32'hc258aef8} /* (30, 4, 3) {real, imag} */,
  {32'hc3e2ee3b, 32'h44515d55} /* (30, 4, 2) {real, imag} */,
  {32'h43618f6e, 32'hc497ddf0} /* (30, 4, 1) {real, imag} */,
  {32'h40c9c47c, 32'hc3d13c11} /* (30, 4, 0) {real, imag} */,
  {32'h44129068, 32'h4417f8ec} /* (30, 3, 31) {real, imag} */,
  {32'hc41fb1a4, 32'hc31f25cc} /* (30, 3, 30) {real, imag} */,
  {32'h41ce3310, 32'hc254dfda} /* (30, 3, 29) {real, imag} */,
  {32'h43166d0a, 32'hc376549f} /* (30, 3, 28) {real, imag} */,
  {32'h42bbe6eb, 32'h431587f0} /* (30, 3, 27) {real, imag} */,
  {32'h42dc9fd8, 32'hc2d1fd88} /* (30, 3, 26) {real, imag} */,
  {32'hbfd97380, 32'hc1fa0100} /* (30, 3, 25) {real, imag} */,
  {32'hc33712ea, 32'h42f4e2b8} /* (30, 3, 24) {real, imag} */,
  {32'h42513125, 32'hc0aeb01c} /* (30, 3, 23) {real, imag} */,
  {32'h4316d8fe, 32'hc252c26f} /* (30, 3, 22) {real, imag} */,
  {32'hc0cf8e34, 32'h3fbb3640} /* (30, 3, 21) {real, imag} */,
  {32'hc212a288, 32'h429596f2} /* (30, 3, 20) {real, imag} */,
  {32'hc2d6742c, 32'h41dbaf80} /* (30, 3, 19) {real, imag} */,
  {32'hc2588b41, 32'hc1c6f5b0} /* (30, 3, 18) {real, imag} */,
  {32'h415f5bd0, 32'hc11b8064} /* (30, 3, 17) {real, imag} */,
  {32'hc1d7a2be, 32'h3fd33a80} /* (30, 3, 16) {real, imag} */,
  {32'h4139fff0, 32'hc21fd0c9} /* (30, 3, 15) {real, imag} */,
  {32'hc26f3b1f, 32'h41ecd2d0} /* (30, 3, 14) {real, imag} */,
  {32'hc1c28a98, 32'hc0efafc0} /* (30, 3, 13) {real, imag} */,
  {32'hc1a3c080, 32'h425f870c} /* (30, 3, 12) {real, imag} */,
  {32'h422cb8da, 32'hc2898de2} /* (30, 3, 11) {real, imag} */,
  {32'h4172a660, 32'h40ce0308} /* (30, 3, 10) {real, imag} */,
  {32'h4135396c, 32'hc0e5d0bc} /* (30, 3, 9) {real, imag} */,
  {32'hc124a1e8, 32'hc2eb6388} /* (30, 3, 8) {real, imag} */,
  {32'h43146677, 32'hc28d3ada} /* (30, 3, 7) {real, imag} */,
  {32'h426f982f, 32'h40a2c878} /* (30, 3, 6) {real, imag} */,
  {32'h414c7078, 32'h42620af7} /* (30, 3, 5) {real, imag} */,
  {32'h435a40d6, 32'h43b03350} /* (30, 3, 4) {real, imag} */,
  {32'h435501b9, 32'hc2906d1b} /* (30, 3, 3) {real, imag} */,
  {32'hc420e53a, 32'h4321ac7e} /* (30, 3, 2) {real, imag} */,
  {32'h43bf7302, 32'hc439e2e8} /* (30, 3, 1) {real, imag} */,
  {32'hc2de3172, 32'h4165d790} /* (30, 3, 0) {real, imag} */,
  {32'h4420accb, 32'h454a49df} /* (30, 2, 31) {real, imag} */,
  {32'hc48f84e8, 32'hc4ffa782} /* (30, 2, 30) {real, imag} */,
  {32'h42dffc3b, 32'h41b87a0e} /* (30, 2, 29) {real, imag} */,
  {32'h44192852, 32'h43926a80} /* (30, 2, 28) {real, imag} */,
  {32'hc3fe4407, 32'hc3872992} /* (30, 2, 27) {real, imag} */,
  {32'hc280071b, 32'hc2f4a9bc} /* (30, 2, 26) {real, imag} */,
  {32'h4399a97f, 32'h424fcd1e} /* (30, 2, 25) {real, imag} */,
  {32'hc41e7e61, 32'hc39704fc} /* (30, 2, 24) {real, imag} */,
  {32'hc1c3dc54, 32'hc271ac7e} /* (30, 2, 23) {real, imag} */,
  {32'h42652a7e, 32'hc0db2100} /* (30, 2, 22) {real, imag} */,
  {32'hc3805cd5, 32'hc1b88854} /* (30, 2, 21) {real, imag} */,
  {32'hc1027f60, 32'h42c591ae} /* (30, 2, 20) {real, imag} */,
  {32'hbfb487c0, 32'hc1902582} /* (30, 2, 19) {real, imag} */,
  {32'hc29567f0, 32'hc259a154} /* (30, 2, 18) {real, imag} */,
  {32'h42de1f3a, 32'hc14b7180} /* (30, 2, 17) {real, imag} */,
  {32'h4214d1ac, 32'hc27691b0} /* (30, 2, 16) {real, imag} */,
  {32'hc1c13a28, 32'h4232bfe0} /* (30, 2, 15) {real, imag} */,
  {32'h430765d0, 32'hc226bd2c} /* (30, 2, 14) {real, imag} */,
  {32'hc1307838, 32'h41dd66ea} /* (30, 2, 13) {real, imag} */,
  {32'h40af64c0, 32'h421d5574} /* (30, 2, 12) {real, imag} */,
  {32'h4322cd9c, 32'hc29e6a47} /* (30, 2, 11) {real, imag} */,
  {32'hc2ba0d4b, 32'h43156a19} /* (30, 2, 10) {real, imag} */,
  {32'hc29f9407, 32'h423fc222} /* (30, 2, 9) {real, imag} */,
  {32'h43653395, 32'hc3c3db1c} /* (30, 2, 8) {real, imag} */,
  {32'h4261e91e, 32'h42bdbe9f} /* (30, 2, 7) {real, imag} */,
  {32'h3f2b0f80, 32'h42c493aa} /* (30, 2, 6) {real, imag} */,
  {32'h440d4af3, 32'hc4111fd5} /* (30, 2, 5) {real, imag} */,
  {32'h426db4a8, 32'h441b221f} /* (30, 2, 4) {real, imag} */,
  {32'h42295796, 32'hc21cfb63} /* (30, 2, 3) {real, imag} */,
  {32'hc465d2b1, 32'hc4a671e6} /* (30, 2, 2) {real, imag} */,
  {32'h44236615, 32'h44de493e} /* (30, 2, 1) {real, imag} */,
  {32'h423a738c, 32'h44cde068} /* (30, 2, 0) {real, imag} */,
  {32'hc48f9594, 32'hc5214223} /* (30, 1, 31) {real, imag} */,
  {32'h4339b1d8, 32'h4477a464} /* (30, 1, 30) {real, imag} */,
  {32'h42f2449b, 32'h435fe64b} /* (30, 1, 29) {real, imag} */,
  {32'h43b1f020, 32'hc43d8e3f} /* (30, 1, 28) {real, imag} */,
  {32'h439993ea, 32'h448fe4ac} /* (30, 1, 27) {real, imag} */,
  {32'h43880448, 32'h430680db} /* (30, 1, 26) {real, imag} */,
  {32'hc3043199, 32'hc2eb5eba} /* (30, 1, 25) {real, imag} */,
  {32'h438f7ca2, 32'h431630d8} /* (30, 1, 24) {real, imag} */,
  {32'hc149fc2e, 32'h42cb6b52} /* (30, 1, 23) {real, imag} */,
  {32'h41700fb8, 32'hc11b6ff0} /* (30, 1, 22) {real, imag} */,
  {32'h4386d478, 32'h431a1dd8} /* (30, 1, 21) {real, imag} */,
  {32'hc154eca6, 32'h417c7af0} /* (30, 1, 20) {real, imag} */,
  {32'h40479920, 32'h42a78be6} /* (30, 1, 19) {real, imag} */,
  {32'h42e67c74, 32'hc1cecd08} /* (30, 1, 18) {real, imag} */,
  {32'hbf84d780, 32'h4108b740} /* (30, 1, 17) {real, imag} */,
  {32'h4176d240, 32'hc1d4e740} /* (30, 1, 16) {real, imag} */,
  {32'h427a7804, 32'h42042ef0} /* (30, 1, 15) {real, imag} */,
  {32'hc300f966, 32'hc233731c} /* (30, 1, 14) {real, imag} */,
  {32'h4171fb38, 32'hc207b4f1} /* (30, 1, 13) {real, imag} */,
  {32'hc14d603a, 32'hc22f69b4} /* (30, 1, 12) {real, imag} */,
  {32'hc2db0e2e, 32'h4312e070} /* (30, 1, 11) {real, imag} */,
  {32'h420eca06, 32'h42e146ee} /* (30, 1, 10) {real, imag} */,
  {32'hc229f10c, 32'h4198cb18} /* (30, 1, 9) {real, imag} */,
  {32'hc3d7245c, 32'h4392be8c} /* (30, 1, 8) {real, imag} */,
  {32'h43281887, 32'hc3087eff} /* (30, 1, 7) {real, imag} */,
  {32'h41502990, 32'h42845b7a} /* (30, 1, 6) {real, imag} */,
  {32'hc33815ed, 32'h4417d19a} /* (30, 1, 5) {real, imag} */,
  {32'h43749288, 32'hc2077330} /* (30, 1, 4) {real, imag} */,
  {32'h423fa34a, 32'h436f7131} /* (30, 1, 3) {real, imag} */,
  {32'hc49c278f, 32'h44efe52a} /* (30, 1, 2) {real, imag} */,
  {32'h449a8ca6, 32'hc57e51cd} /* (30, 1, 1) {real, imag} */,
  {32'hc3baea6e, 32'hc51dc3f4} /* (30, 1, 0) {real, imag} */,
  {32'hc4cff07a, 32'hc4b2125a} /* (30, 0, 31) {real, imag} */,
  {32'h444404b0, 32'h438b545d} /* (30, 0, 30) {real, imag} */,
  {32'h430c00ce, 32'h4341eae5} /* (30, 0, 29) {real, imag} */,
  {32'h433dad19, 32'h41b42216} /* (30, 0, 28) {real, imag} */,
  {32'h42c38d3c, 32'h43f507e0} /* (30, 0, 27) {real, imag} */,
  {32'hc2cfe556, 32'h427a6036} /* (30, 0, 26) {real, imag} */,
  {32'hc3cae62c, 32'h429552c5} /* (30, 0, 25) {real, imag} */,
  {32'h43acbdad, 32'hc276a2ae} /* (30, 0, 24) {real, imag} */,
  {32'h423864c0, 32'h42eac555} /* (30, 0, 23) {real, imag} */,
  {32'h428c045b, 32'hc27bd012} /* (30, 0, 22) {real, imag} */,
  {32'h42b0cc68, 32'hc0de7b70} /* (30, 0, 21) {real, imag} */,
  {32'h426a2688, 32'h42084516} /* (30, 0, 20) {real, imag} */,
  {32'hc2782e0f, 32'h426edb9a} /* (30, 0, 19) {real, imag} */,
  {32'hc1a7126c, 32'hc17d1f48} /* (30, 0, 18) {real, imag} */,
  {32'h418f8c50, 32'hc0e49340} /* (30, 0, 17) {real, imag} */,
  {32'hc1989560, 32'h41cb7780} /* (30, 0, 16) {real, imag} */,
  {32'h41ffb550, 32'hc239dfd8} /* (30, 0, 15) {real, imag} */,
  {32'hc1bf586c, 32'h4092fd90} /* (30, 0, 14) {real, imag} */,
  {32'h424340a5, 32'h41c16e8c} /* (30, 0, 13) {real, imag} */,
  {32'h42c660fc, 32'hc2f57d49} /* (30, 0, 12) {real, imag} */,
  {32'hc1ac7e70, 32'h42bac327} /* (30, 0, 11) {real, imag} */,
  {32'hc2180096, 32'h42b3be15} /* (30, 0, 10) {real, imag} */,
  {32'h4108f680, 32'h42b9d653} /* (30, 0, 9) {real, imag} */,
  {32'hc3636826, 32'h416d7678} /* (30, 0, 8) {real, imag} */,
  {32'h429edf80, 32'hc279e11a} /* (30, 0, 7) {real, imag} */,
  {32'hc1cc0ed0, 32'h42fda7a9} /* (30, 0, 6) {real, imag} */,
  {32'h42bef660, 32'h44027b6e} /* (30, 0, 5) {real, imag} */,
  {32'hc3e057a2, 32'hc1c906de} /* (30, 0, 4) {real, imag} */,
  {32'h41155278, 32'h432e916b} /* (30, 0, 3) {real, imag} */,
  {32'hc435d57c, 32'h44207178} /* (30, 0, 2) {real, imag} */,
  {32'h4470e104, 32'hc4ec0e8e} /* (30, 0, 1) {real, imag} */,
  {32'hc3b53fda, 32'hc4cad3ee} /* (30, 0, 0) {real, imag} */,
  {32'hc490dbee, 32'hc49f9f39} /* (29, 31, 31) {real, imag} */,
  {32'h443d8d10, 32'h43f3f585} /* (29, 31, 30) {real, imag} */,
  {32'h437c33fa, 32'hc2ecd2e0} /* (29, 31, 29) {real, imag} */,
  {32'h41c73958, 32'hc31cecfa} /* (29, 31, 28) {real, imag} */,
  {32'h4335198a, 32'h43905df3} /* (29, 31, 27) {real, imag} */,
  {32'hc30eebc3, 32'h42ca7150} /* (29, 31, 26) {real, imag} */,
  {32'hc2b4bb4c, 32'h431d7d20} /* (29, 31, 25) {real, imag} */,
  {32'h4327304c, 32'h416b47f8} /* (29, 31, 24) {real, imag} */,
  {32'h4311f08c, 32'hc185475c} /* (29, 31, 23) {real, imag} */,
  {32'hc22eff9c, 32'h4312eb82} /* (29, 31, 22) {real, imag} */,
  {32'h430c5e51, 32'h41d67054} /* (29, 31, 21) {real, imag} */,
  {32'h420290c7, 32'hc20fa2c4} /* (29, 31, 20) {real, imag} */,
  {32'hc2decf02, 32'h420c1d73} /* (29, 31, 19) {real, imag} */,
  {32'h4203b3a8, 32'hc276ad63} /* (29, 31, 18) {real, imag} */,
  {32'hc0c5df00, 32'h420106c4} /* (29, 31, 17) {real, imag} */,
  {32'h4232219c, 32'hc1efc280} /* (29, 31, 16) {real, imag} */,
  {32'hc1966280, 32'h420fadfc} /* (29, 31, 15) {real, imag} */,
  {32'hc2904f90, 32'h40b4e5d8} /* (29, 31, 14) {real, imag} */,
  {32'hc24cd8fc, 32'hc12a8b44} /* (29, 31, 13) {real, imag} */,
  {32'hc24d66e1, 32'hc253515c} /* (29, 31, 12) {real, imag} */,
  {32'hc14fa2b0, 32'h42cd8983} /* (29, 31, 11) {real, imag} */,
  {32'h4260c774, 32'hc28d70ef} /* (29, 31, 10) {real, imag} */,
  {32'h421398f6, 32'h41d6e6bc} /* (29, 31, 9) {real, imag} */,
  {32'hc2ad06e4, 32'h43227cf8} /* (29, 31, 8) {real, imag} */,
  {32'h4343b622, 32'hc246308e} /* (29, 31, 7) {real, imag} */,
  {32'hc20418dc, 32'h42a38482} /* (29, 31, 6) {real, imag} */,
  {32'h4317f194, 32'h43d51bf3} /* (29, 31, 5) {real, imag} */,
  {32'hc38630c0, 32'hc386405f} /* (29, 31, 4) {real, imag} */,
  {32'hc27a1988, 32'h4375788c} /* (29, 31, 3) {real, imag} */,
  {32'h435cca18, 32'h439c594f} /* (29, 31, 2) {real, imag} */,
  {32'hc2e9c6c8, 32'hc49561f5} /* (29, 31, 1) {real, imag} */,
  {32'hc3b9ef3e, 32'hc46e4f86} /* (29, 31, 0) {real, imag} */,
  {32'h3fbed500, 32'h44269688} /* (29, 30, 31) {real, imag} */,
  {32'hc11aed1c, 32'hc40fadbf} /* (29, 30, 30) {real, imag} */,
  {32'hc294d17f, 32'h429d4716} /* (29, 30, 29) {real, imag} */,
  {32'h4323a17e, 32'h4309011a} /* (29, 30, 28) {real, imag} */,
  {32'hc2cd7983, 32'hc331b72a} /* (29, 30, 27) {real, imag} */,
  {32'h417f00da, 32'h42028cfe} /* (29, 30, 26) {real, imag} */,
  {32'h42bb17dc, 32'h423e1ef0} /* (29, 30, 25) {real, imag} */,
  {32'hc0d1b190, 32'h3ffe5240} /* (29, 30, 24) {real, imag} */,
  {32'hc290b252, 32'hc1e40b90} /* (29, 30, 23) {real, imag} */,
  {32'h42836c33, 32'h427597c8} /* (29, 30, 22) {real, imag} */,
  {32'hc2364a56, 32'hc192abd4} /* (29, 30, 21) {real, imag} */,
  {32'h42726f92, 32'h42423112} /* (29, 30, 20) {real, imag} */,
  {32'hc068e3f0, 32'hc17b29b6} /* (29, 30, 19) {real, imag} */,
  {32'hc03c48a0, 32'h41aa31c0} /* (29, 30, 18) {real, imag} */,
  {32'hbff716c0, 32'h421abf14} /* (29, 30, 17) {real, imag} */,
  {32'h3f724500, 32'hc21c49ac} /* (29, 30, 16) {real, imag} */,
  {32'hc201c7b6, 32'h40f61460} /* (29, 30, 15) {real, imag} */,
  {32'h4132b4b0, 32'h41478200} /* (29, 30, 14) {real, imag} */,
  {32'h425e6a05, 32'hc196e3ed} /* (29, 30, 13) {real, imag} */,
  {32'hc1bc2c1b, 32'hc2693b0e} /* (29, 30, 12) {real, imag} */,
  {32'h42881bb5, 32'h42862667} /* (29, 30, 11) {real, imag} */,
  {32'hc314726c, 32'h41982ca4} /* (29, 30, 10) {real, imag} */,
  {32'hc275f065, 32'hc25e5328} /* (29, 30, 9) {real, imag} */,
  {32'h4256f266, 32'hc3216a1a} /* (29, 30, 8) {real, imag} */,
  {32'h4117a2e4, 32'hc079e800} /* (29, 30, 7) {real, imag} */,
  {32'h4232621e, 32'hc238be28} /* (29, 30, 6) {real, imag} */,
  {32'h42f3d155, 32'hc3565b26} /* (29, 30, 5) {real, imag} */,
  {32'hc35ca5ea, 32'h42b56009} /* (29, 30, 4) {real, imag} */,
  {32'h411cc4d8, 32'h42f3afae} /* (29, 30, 3) {real, imag} */,
  {32'hc2fe8570, 32'hc45151ab} /* (29, 30, 2) {real, imag} */,
  {32'h43f1cfbd, 32'h44a748c3} /* (29, 30, 1) {real, imag} */,
  {32'h4393e7b0, 32'h43da52de} /* (29, 30, 0) {real, imag} */,
  {32'hc34535c4, 32'hc21a0770} /* (29, 29, 31) {real, imag} */,
  {32'h4348cdb4, 32'hc342bc9b} /* (29, 29, 30) {real, imag} */,
  {32'hc20bbf00, 32'hc30e3076} /* (29, 29, 29) {real, imag} */,
  {32'hc2b4845c, 32'h438e6b02} /* (29, 29, 28) {real, imag} */,
  {32'hc27635fc, 32'hc31150e8} /* (29, 29, 27) {real, imag} */,
  {32'h42f12712, 32'hc277e2be} /* (29, 29, 26) {real, imag} */,
  {32'hc2d79894, 32'h4287ec15} /* (29, 29, 25) {real, imag} */,
  {32'h4151bf80, 32'hc2906aff} /* (29, 29, 24) {real, imag} */,
  {32'hc2e8a09f, 32'h40f6d5f4} /* (29, 29, 23) {real, imag} */,
  {32'h4269b175, 32'hc231e282} /* (29, 29, 22) {real, imag} */,
  {32'h40a12cec, 32'hc248b006} /* (29, 29, 21) {real, imag} */,
  {32'h426be6b6, 32'hc2753fc5} /* (29, 29, 20) {real, imag} */,
  {32'h41a80afc, 32'hc2155288} /* (29, 29, 19) {real, imag} */,
  {32'h4131e518, 32'h4201cb2e} /* (29, 29, 18) {real, imag} */,
  {32'hc21fb1be, 32'h4190bba0} /* (29, 29, 17) {real, imag} */,
  {32'h424e0df4, 32'h4214de02} /* (29, 29, 16) {real, imag} */,
  {32'h4249aeb8, 32'hc1d495b8} /* (29, 29, 15) {real, imag} */,
  {32'h425b19ea, 32'hc1bee993} /* (29, 29, 14) {real, imag} */,
  {32'hc2dfa02b, 32'hc1951d61} /* (29, 29, 13) {real, imag} */,
  {32'h41e5fa20, 32'hc17d17ec} /* (29, 29, 12) {real, imag} */,
  {32'h40d198ec, 32'h40af4acc} /* (29, 29, 11) {real, imag} */,
  {32'hc2269809, 32'h42823fdf} /* (29, 29, 10) {real, imag} */,
  {32'hc2e99b35, 32'hc1987b9d} /* (29, 29, 9) {real, imag} */,
  {32'h438ed91b, 32'hc248351e} /* (29, 29, 8) {real, imag} */,
  {32'hc280eaf8, 32'h4339c366} /* (29, 29, 7) {real, imag} */,
  {32'h431681a7, 32'hbf12b5c0} /* (29, 29, 6) {real, imag} */,
  {32'h429910a4, 32'h424c3bd0} /* (29, 29, 5) {real, imag} */,
  {32'hc2b75bd8, 32'hc0dc1cc0} /* (29, 29, 4) {real, imag} */,
  {32'hc0c1033c, 32'h40ead730} /* (29, 29, 3) {real, imag} */,
  {32'h418c6614, 32'hc3244571} /* (29, 29, 2) {real, imag} */,
  {32'hc26fe028, 32'h439a68c2} /* (29, 29, 1) {real, imag} */,
  {32'hc22ca1ac, 32'h433e3ef8} /* (29, 29, 0) {real, imag} */,
  {32'hc3739e1b, 32'hc398bea1} /* (29, 28, 31) {real, imag} */,
  {32'h43b6d26d, 32'h431d9ee4} /* (29, 28, 30) {real, imag} */,
  {32'h4301aa1c, 32'h4288865a} /* (29, 28, 29) {real, imag} */,
  {32'hc35ca69c, 32'hc2ff1557} /* (29, 28, 28) {real, imag} */,
  {32'h43202c9e, 32'h4215bdda} /* (29, 28, 27) {real, imag} */,
  {32'hc04da6a0, 32'hc28fc411} /* (29, 28, 26) {real, imag} */,
  {32'h42bad0a2, 32'h3fa167d0} /* (29, 28, 25) {real, imag} */,
  {32'h42a1d7cd, 32'h42ba1026} /* (29, 28, 24) {real, imag} */,
  {32'h429d16a2, 32'h4169d1fe} /* (29, 28, 23) {real, imag} */,
  {32'hc2a2b46d, 32'hc1b98a3e} /* (29, 28, 22) {real, imag} */,
  {32'h42583bbc, 32'hc2087adc} /* (29, 28, 21) {real, imag} */,
  {32'hbf5cf840, 32'h41c08c5e} /* (29, 28, 20) {real, imag} */,
  {32'h415b9b70, 32'h411d67b4} /* (29, 28, 19) {real, imag} */,
  {32'h423607bb, 32'h41e93018} /* (29, 28, 18) {real, imag} */,
  {32'h415c511a, 32'h425ca3e3} /* (29, 28, 17) {real, imag} */,
  {32'h4076f4a0, 32'hbff64100} /* (29, 28, 16) {real, imag} */,
  {32'h41894563, 32'hc1a377c6} /* (29, 28, 15) {real, imag} */,
  {32'h4142c1d4, 32'h418c8040} /* (29, 28, 14) {real, imag} */,
  {32'h409acb20, 32'hc181f396} /* (29, 28, 13) {real, imag} */,
  {32'h41c5716a, 32'hc2060a1b} /* (29, 28, 12) {real, imag} */,
  {32'hc1ba3ca0, 32'h424b4d88} /* (29, 28, 11) {real, imag} */,
  {32'hc2248982, 32'hc264840d} /* (29, 28, 10) {real, imag} */,
  {32'hc05011c0, 32'h422848f2} /* (29, 28, 9) {real, imag} */,
  {32'h427166da, 32'h417c37c0} /* (29, 28, 8) {real, imag} */,
  {32'h4295983a, 32'h4235f9b4} /* (29, 28, 7) {real, imag} */,
  {32'hc21004c2, 32'h42e1b6cb} /* (29, 28, 6) {real, imag} */,
  {32'h40ebaf40, 32'h432cc5a6} /* (29, 28, 5) {real, imag} */,
  {32'hbf9838c0, 32'hc2f03fbf} /* (29, 28, 4) {real, imag} */,
  {32'hc2c27495, 32'hc208deef} /* (29, 28, 3) {real, imag} */,
  {32'h43803921, 32'h434ba7fc} /* (29, 28, 2) {real, imag} */,
  {32'hc396a54a, 32'hc3319041} /* (29, 28, 1) {real, imag} */,
  {32'hc2962749, 32'hc3c7cf61} /* (29, 28, 0) {real, imag} */,
  {32'h43d2f20f, 32'h43268130} /* (29, 27, 31) {real, imag} */,
  {32'hc1f7e393, 32'hc31ea27c} /* (29, 27, 30) {real, imag} */,
  {32'hc2bafe02, 32'h41a51018} /* (29, 27, 29) {real, imag} */,
  {32'hc1cc8edb, 32'h4201246a} /* (29, 27, 28) {real, imag} */,
  {32'hc32e4aa7, 32'h42dc03ee} /* (29, 27, 27) {real, imag} */,
  {32'h42239d58, 32'hc294977b} /* (29, 27, 26) {real, imag} */,
  {32'h42f039ec, 32'hc14ec69e} /* (29, 27, 25) {real, imag} */,
  {32'hc2085e88, 32'hc271071b} /* (29, 27, 24) {real, imag} */,
  {32'h428ad328, 32'hc24e2b04} /* (29, 27, 23) {real, imag} */,
  {32'hc2664c4e, 32'hc2733bba} /* (29, 27, 22) {real, imag} */,
  {32'h410b4320, 32'h42609603} /* (29, 27, 21) {real, imag} */,
  {32'h41e7aa32, 32'hc24fdc4c} /* (29, 27, 20) {real, imag} */,
  {32'h40b65128, 32'h4032d840} /* (29, 27, 19) {real, imag} */,
  {32'hc23b65da, 32'h406dce04} /* (29, 27, 18) {real, imag} */,
  {32'hc1329818, 32'hc10828a0} /* (29, 27, 17) {real, imag} */,
  {32'hc18bc1c4, 32'hc2529c88} /* (29, 27, 16) {real, imag} */,
  {32'hbf81fb40, 32'hc1afa890} /* (29, 27, 15) {real, imag} */,
  {32'hc1f29a8d, 32'hc1c3e0b8} /* (29, 27, 14) {real, imag} */,
  {32'h427bd61b, 32'h40cdde00} /* (29, 27, 13) {real, imag} */,
  {32'h4213a2d3, 32'h418206e4} /* (29, 27, 12) {real, imag} */,
  {32'h421624b0, 32'hc21a92bd} /* (29, 27, 11) {real, imag} */,
  {32'hc21e19a6, 32'h40b0a254} /* (29, 27, 10) {real, imag} */,
  {32'h4221601f, 32'h41d69cbb} /* (29, 27, 9) {real, imag} */,
  {32'h42c3d770, 32'h42909d12} /* (29, 27, 8) {real, imag} */,
  {32'hc31764a0, 32'h4252af56} /* (29, 27, 7) {real, imag} */,
  {32'hc2af94e0, 32'h42288bce} /* (29, 27, 6) {real, imag} */,
  {32'hc21f8ef4, 32'hc335da33} /* (29, 27, 5) {real, imag} */,
  {32'h41871689, 32'h425cf160} /* (29, 27, 4) {real, imag} */,
  {32'hc16a5314, 32'hc2f876e0} /* (29, 27, 3) {real, imag} */,
  {32'hc294e3e9, 32'hc3652a78} /* (29, 27, 2) {real, imag} */,
  {32'h4306491a, 32'h43eace32} /* (29, 27, 1) {real, imag} */,
  {32'h430edccc, 32'h43705470} /* (29, 27, 0) {real, imag} */,
  {32'hc08bc390, 32'h4308a489} /* (29, 26, 31) {real, imag} */,
  {32'h423434a6, 32'h4320df64} /* (29, 26, 30) {real, imag} */,
  {32'h42a00ccf, 32'h41da2589} /* (29, 26, 29) {real, imag} */,
  {32'hc1fd37b9, 32'hc14c6382} /* (29, 26, 28) {real, imag} */,
  {32'hc25a6d3e, 32'h40aed530} /* (29, 26, 27) {real, imag} */,
  {32'hc28d582f, 32'hc1d92ee2} /* (29, 26, 26) {real, imag} */,
  {32'hc350e1a3, 32'hc2ee1f9e} /* (29, 26, 25) {real, imag} */,
  {32'h42037188, 32'h426a7fcc} /* (29, 26, 24) {real, imag} */,
  {32'hc1b46039, 32'h409d0640} /* (29, 26, 23) {real, imag} */,
  {32'hc18fca36, 32'h42030b17} /* (29, 26, 22) {real, imag} */,
  {32'hc1bd3dc2, 32'hc1b17498} /* (29, 26, 21) {real, imag} */,
  {32'hc28946a7, 32'hc1b56639} /* (29, 26, 20) {real, imag} */,
  {32'hc1bb5419, 32'hc11315fa} /* (29, 26, 19) {real, imag} */,
  {32'h4136db84, 32'h4055d9d0} /* (29, 26, 18) {real, imag} */,
  {32'hc15ba5e5, 32'h41f70bee} /* (29, 26, 17) {real, imag} */,
  {32'hc1ead7be, 32'h4189763a} /* (29, 26, 16) {real, imag} */,
  {32'h41605295, 32'h41ae6192} /* (29, 26, 15) {real, imag} */,
  {32'hc248af90, 32'hc1767674} /* (29, 26, 14) {real, imag} */,
  {32'h4229b7dc, 32'hc189972f} /* (29, 26, 13) {real, imag} */,
  {32'h4252bbe4, 32'h41c50423} /* (29, 26, 12) {real, imag} */,
  {32'h41bdaebc, 32'hc1c4bbce} /* (29, 26, 11) {real, imag} */,
  {32'h414e4240, 32'h42a5b3d6} /* (29, 26, 10) {real, imag} */,
  {32'hc001a938, 32'hc325ee80} /* (29, 26, 9) {real, imag} */,
  {32'h408d6e9c, 32'h4178f8e8} /* (29, 26, 8) {real, imag} */,
  {32'hc29a75da, 32'h4224d705} /* (29, 26, 7) {real, imag} */,
  {32'h428d53ff, 32'hc2e6ffca} /* (29, 26, 6) {real, imag} */,
  {32'h42029042, 32'h42fd7113} /* (29, 26, 5) {real, imag} */,
  {32'hc0a660d4, 32'h41e978d7} /* (29, 26, 4) {real, imag} */,
  {32'hc1a02d23, 32'h41374dde} /* (29, 26, 3) {real, imag} */,
  {32'h423c4596, 32'h429bf081} /* (29, 26, 2) {real, imag} */,
  {32'hc29e4cf5, 32'h4286638e} /* (29, 26, 1) {real, imag} */,
  {32'h422f9e37, 32'hc2b04e70} /* (29, 26, 0) {real, imag} */,
  {32'hc0e8fd34, 32'hc207fff5} /* (29, 25, 31) {real, imag} */,
  {32'h428712e4, 32'h423f3df0} /* (29, 25, 30) {real, imag} */,
  {32'h42ade4d2, 32'hc21fbdd8} /* (29, 25, 29) {real, imag} */,
  {32'hc2da0f3e, 32'hc2bba650} /* (29, 25, 28) {real, imag} */,
  {32'h42bfc94c, 32'hc29479b0} /* (29, 25, 27) {real, imag} */,
  {32'h41a91c79, 32'hc1e92690} /* (29, 25, 26) {real, imag} */,
  {32'hc2262d40, 32'h41e06cf5} /* (29, 25, 25) {real, imag} */,
  {32'h417e47f8, 32'h41d88c33} /* (29, 25, 24) {real, imag} */,
  {32'hc2803f6e, 32'h3f030f60} /* (29, 25, 23) {real, imag} */,
  {32'h42d30b97, 32'hc1bf68be} /* (29, 25, 22) {real, imag} */,
  {32'hc13af7e6, 32'hc1b63460} /* (29, 25, 21) {real, imag} */,
  {32'h41a59d9e, 32'h40f521c2} /* (29, 25, 20) {real, imag} */,
  {32'h42145ac8, 32'h41257040} /* (29, 25, 19) {real, imag} */,
  {32'hc2100f70, 32'hc106978a} /* (29, 25, 18) {real, imag} */,
  {32'h420bd6d2, 32'hc00b0c24} /* (29, 25, 17) {real, imag} */,
  {32'h408d7c2a, 32'hc13217b8} /* (29, 25, 16) {real, imag} */,
  {32'h41fa1d60, 32'h4181b31e} /* (29, 25, 15) {real, imag} */,
  {32'h4129e350, 32'hc24a54da} /* (29, 25, 14) {real, imag} */,
  {32'h41ae2193, 32'hc2880cb5} /* (29, 25, 13) {real, imag} */,
  {32'hc242e009, 32'h41f10370} /* (29, 25, 12) {real, imag} */,
  {32'hc24061f4, 32'hc09a3a4a} /* (29, 25, 11) {real, imag} */,
  {32'hc229c60e, 32'hbe0be000} /* (29, 25, 10) {real, imag} */,
  {32'h40c2a9a8, 32'h4233d7a6} /* (29, 25, 9) {real, imag} */,
  {32'hc2050816, 32'hc1cf8699} /* (29, 25, 8) {real, imag} */,
  {32'h422f0cc8, 32'h4200c0b2} /* (29, 25, 7) {real, imag} */,
  {32'h41681952, 32'hc2caecca} /* (29, 25, 6) {real, imag} */,
  {32'h4182bcda, 32'h41fed316} /* (29, 25, 5) {real, imag} */,
  {32'h42856c24, 32'hc2b1b920} /* (29, 25, 4) {real, imag} */,
  {32'h41deff9a, 32'hc27546aa} /* (29, 25, 3) {real, imag} */,
  {32'h3fed8a60, 32'h403b2208} /* (29, 25, 2) {real, imag} */,
  {32'h423076bc, 32'h4232ca43} /* (29, 25, 1) {real, imag} */,
  {32'h418387a8, 32'hc2eb6a65} /* (29, 25, 0) {real, imag} */,
  {32'h42e7b9a8, 32'h41132ad8} /* (29, 24, 31) {real, imag} */,
  {32'hc1af1fa2, 32'hc2be3ce8} /* (29, 24, 30) {real, imag} */,
  {32'hc2f808f4, 32'h42a44dbc} /* (29, 24, 29) {real, imag} */,
  {32'h420619a0, 32'hc2e4b3a3} /* (29, 24, 28) {real, imag} */,
  {32'hc1954455, 32'h4294b6ba} /* (29, 24, 27) {real, imag} */,
  {32'h3fca9440, 32'hc23b81b2} /* (29, 24, 26) {real, imag} */,
  {32'hc2a9ebe8, 32'h4139d652} /* (29, 24, 25) {real, imag} */,
  {32'hc2e1ea56, 32'h41ba126a} /* (29, 24, 24) {real, imag} */,
  {32'h41af1869, 32'h426d7f2e} /* (29, 24, 23) {real, imag} */,
  {32'hc0df400c, 32'hc2ca7580} /* (29, 24, 22) {real, imag} */,
  {32'hc2b4911c, 32'h4288fe0c} /* (29, 24, 21) {real, imag} */,
  {32'h4199747c, 32'h41b9a9c0} /* (29, 24, 20) {real, imag} */,
  {32'hc1dc8429, 32'hc02f686e} /* (29, 24, 19) {real, imag} */,
  {32'h403d8e10, 32'h412b3e47} /* (29, 24, 18) {real, imag} */,
  {32'h4003f905, 32'h412c3c2c} /* (29, 24, 17) {real, imag} */,
  {32'hc1972066, 32'hbffe8b00} /* (29, 24, 16) {real, imag} */,
  {32'h4081045e, 32'h41d57d22} /* (29, 24, 15) {real, imag} */,
  {32'h413f6402, 32'h414bce21} /* (29, 24, 14) {real, imag} */,
  {32'h41eab061, 32'hc139719c} /* (29, 24, 13) {real, imag} */,
  {32'hc0d10834, 32'hc0d67b40} /* (29, 24, 12) {real, imag} */,
  {32'hc2306cc4, 32'h41e50fca} /* (29, 24, 11) {real, imag} */,
  {32'hc0c157d4, 32'hc211af98} /* (29, 24, 10) {real, imag} */,
  {32'h41f6db09, 32'hbf2d2460} /* (29, 24, 9) {real, imag} */,
  {32'h41fe9020, 32'h4179c12c} /* (29, 24, 8) {real, imag} */,
  {32'h42e48f04, 32'h424fa266} /* (29, 24, 7) {real, imag} */,
  {32'h42ca45dd, 32'h41da6bbc} /* (29, 24, 6) {real, imag} */,
  {32'hc10c9246, 32'h4187d8fe} /* (29, 24, 5) {real, imag} */,
  {32'hc1bce2d3, 32'hc2019e9e} /* (29, 24, 4) {real, imag} */,
  {32'hc233f0ed, 32'h42289476} /* (29, 24, 3) {real, imag} */,
  {32'hc0105558, 32'hc3124676} /* (29, 24, 2) {real, imag} */,
  {32'h42cf3762, 32'h4322f266} /* (29, 24, 1) {real, imag} */,
  {32'h4295147a, 32'h42ea27f6} /* (29, 24, 0) {real, imag} */,
  {32'hc1a28894, 32'hc33f06c8} /* (29, 23, 31) {real, imag} */,
  {32'hc2665a42, 32'h4181fe32} /* (29, 23, 30) {real, imag} */,
  {32'h41b84d18, 32'h423e9d6e} /* (29, 23, 29) {real, imag} */,
  {32'hc19bf0e6, 32'hc25ecc94} /* (29, 23, 28) {real, imag} */,
  {32'hc2ddd7c6, 32'h42154068} /* (29, 23, 27) {real, imag} */,
  {32'hc24603f8, 32'h420e3438} /* (29, 23, 26) {real, imag} */,
  {32'h421173f5, 32'h4165eae5} /* (29, 23, 25) {real, imag} */,
  {32'h411f3d84, 32'hc1ede882} /* (29, 23, 24) {real, imag} */,
  {32'h410a7659, 32'h4222197c} /* (29, 23, 23) {real, imag} */,
  {32'h4205812a, 32'hc243e931} /* (29, 23, 22) {real, imag} */,
  {32'h41c46804, 32'hc103f459} /* (29, 23, 21) {real, imag} */,
  {32'h412f173d, 32'h40d687b8} /* (29, 23, 20) {real, imag} */,
  {32'hc1b03020, 32'h416ef376} /* (29, 23, 19) {real, imag} */,
  {32'hc1b41663, 32'h40c85a80} /* (29, 23, 18) {real, imag} */,
  {32'hc073f594, 32'hc097f1d8} /* (29, 23, 17) {real, imag} */,
  {32'hc0dde594, 32'hc0d32aec} /* (29, 23, 16) {real, imag} */,
  {32'hc1121583, 32'h3f49c540} /* (29, 23, 15) {real, imag} */,
  {32'h41cd9e79, 32'hc123f46c} /* (29, 23, 14) {real, imag} */,
  {32'hc1853528, 32'h426465c2} /* (29, 23, 13) {real, imag} */,
  {32'h41456739, 32'h42181171} /* (29, 23, 12) {real, imag} */,
  {32'hc1d3e2b4, 32'hc205e877} /* (29, 23, 11) {real, imag} */,
  {32'h41d9940a, 32'hc20d2a07} /* (29, 23, 10) {real, imag} */,
  {32'h41ad8804, 32'h41d3a513} /* (29, 23, 9) {real, imag} */,
  {32'hc15bbcbc, 32'hc1844f28} /* (29, 23, 8) {real, imag} */,
  {32'hc254eafd, 32'h41528f79} /* (29, 23, 7) {real, imag} */,
  {32'hc1e75c84, 32'h42a3f96a} /* (29, 23, 6) {real, imag} */,
  {32'h42a4cbc4, 32'h429d598e} /* (29, 23, 5) {real, imag} */,
  {32'h4238b899, 32'h431aa75f} /* (29, 23, 4) {real, imag} */,
  {32'hc3087acc, 32'hc226fbfa} /* (29, 23, 3) {real, imag} */,
  {32'h42a7e9ab, 32'hc1b47d80} /* (29, 23, 2) {real, imag} */,
  {32'hc27795e8, 32'h42ed6d13} /* (29, 23, 1) {real, imag} */,
  {32'h4234a610, 32'h420ac6de} /* (29, 23, 0) {real, imag} */,
  {32'hc2d3e324, 32'hc1897a88} /* (29, 22, 31) {real, imag} */,
  {32'h429f5756, 32'hc27b698b} /* (29, 22, 30) {real, imag} */,
  {32'h42a6c17b, 32'h42529d9c} /* (29, 22, 29) {real, imag} */,
  {32'h3f83c350, 32'hc048e4fc} /* (29, 22, 28) {real, imag} */,
  {32'h4180d284, 32'h42a307a4} /* (29, 22, 27) {real, imag} */,
  {32'h42083e74, 32'h42dd4fa1} /* (29, 22, 26) {real, imag} */,
  {32'h4166134f, 32'h421f5bae} /* (29, 22, 25) {real, imag} */,
  {32'hc251cbbe, 32'h4016e708} /* (29, 22, 24) {real, imag} */,
  {32'h4194554e, 32'h4149a738} /* (29, 22, 23) {real, imag} */,
  {32'hc1bad715, 32'h422013f4} /* (29, 22, 22) {real, imag} */,
  {32'hbf0cf880, 32'h4141f05e} /* (29, 22, 21) {real, imag} */,
  {32'hc1eec019, 32'hbfc6f190} /* (29, 22, 20) {real, imag} */,
  {32'hc1025e0a, 32'hc21b5d9a} /* (29, 22, 19) {real, imag} */,
  {32'hc12ebe65, 32'h40a2c992} /* (29, 22, 18) {real, imag} */,
  {32'h41b2c20f, 32'hc1456150} /* (29, 22, 17) {real, imag} */,
  {32'h40e29554, 32'h4130e058} /* (29, 22, 16) {real, imag} */,
  {32'hc14707f6, 32'h410c7012} /* (29, 22, 15) {real, imag} */,
  {32'h4092b83a, 32'hc087bc42} /* (29, 22, 14) {real, imag} */,
  {32'hc1953b51, 32'h417005ee} /* (29, 22, 13) {real, imag} */,
  {32'h40667548, 32'hc255fb72} /* (29, 22, 12) {real, imag} */,
  {32'hc244b1c8, 32'hc26334c8} /* (29, 22, 11) {real, imag} */,
  {32'h420c61c8, 32'h422c5cf8} /* (29, 22, 10) {real, imag} */,
  {32'hc1ab540c, 32'h4286bf25} /* (29, 22, 9) {real, imag} */,
  {32'h42e001b1, 32'hc1103712} /* (29, 22, 8) {real, imag} */,
  {32'h40eeecce, 32'h3fd13bd0} /* (29, 22, 7) {real, imag} */,
  {32'hc18a8b13, 32'h40cfc7b0} /* (29, 22, 6) {real, imag} */,
  {32'h41d927f0, 32'hc1d0c061} /* (29, 22, 5) {real, imag} */,
  {32'hc1977f49, 32'hc1b37f46} /* (29, 22, 4) {real, imag} */,
  {32'hc1fd9537, 32'hc196a8f3} /* (29, 22, 3) {real, imag} */,
  {32'h42a544ce, 32'hc29ceb6a} /* (29, 22, 2) {real, imag} */,
  {32'hc06ffc70, 32'hc17452f9} /* (29, 22, 1) {real, imag} */,
  {32'hc287fa7f, 32'h433ea4c6} /* (29, 22, 0) {real, imag} */,
  {32'h42cd8756, 32'hc225e6c8} /* (29, 21, 31) {real, imag} */,
  {32'hc2d5d38d, 32'hc1b33722} /* (29, 21, 30) {real, imag} */,
  {32'h41e6e7ba, 32'h41ae5c0b} /* (29, 21, 29) {real, imag} */,
  {32'h41c8cf8c, 32'h424da9f9} /* (29, 21, 28) {real, imag} */,
  {32'hc08fab06, 32'hc1dc678a} /* (29, 21, 27) {real, imag} */,
  {32'hc19d6f14, 32'h4270f351} /* (29, 21, 26) {real, imag} */,
  {32'h42856eb1, 32'hc1e8ee68} /* (29, 21, 25) {real, imag} */,
  {32'hc0639286, 32'h41a6c752} /* (29, 21, 24) {real, imag} */,
  {32'hc15c4fe4, 32'h418f7b70} /* (29, 21, 23) {real, imag} */,
  {32'hc21df5aa, 32'hc20c093f} /* (29, 21, 22) {real, imag} */,
  {32'hc21ac305, 32'h4089e864} /* (29, 21, 21) {real, imag} */,
  {32'hc15f32b2, 32'hbfb9fb48} /* (29, 21, 20) {real, imag} */,
  {32'h419881f2, 32'h41ad29dd} /* (29, 21, 19) {real, imag} */,
  {32'h40546434, 32'h41a272ce} /* (29, 21, 18) {real, imag} */,
  {32'hc11ad89a, 32'h40effd99} /* (29, 21, 17) {real, imag} */,
  {32'hbf903880, 32'h3fbcc784} /* (29, 21, 16) {real, imag} */,
  {32'hbf4bcce0, 32'h3fa80d74} /* (29, 21, 15) {real, imag} */,
  {32'h41dedd20, 32'hc1f0a776} /* (29, 21, 14) {real, imag} */,
  {32'hbf3f9810, 32'hc142a686} /* (29, 21, 13) {real, imag} */,
  {32'h40cfb02c, 32'hc0cf08c6} /* (29, 21, 12) {real, imag} */,
  {32'h42653e83, 32'hc1701b66} /* (29, 21, 11) {real, imag} */,
  {32'hc0b834b4, 32'h421c5c4b} /* (29, 21, 10) {real, imag} */,
  {32'hc0a4fc58, 32'h41ffaeca} /* (29, 21, 9) {real, imag} */,
  {32'hc12fec94, 32'h4267af67} /* (29, 21, 8) {real, imag} */,
  {32'hc2a63933, 32'hc16a0c95} /* (29, 21, 7) {real, imag} */,
  {32'hc24097d4, 32'h41958af6} /* (29, 21, 6) {real, imag} */,
  {32'hc15761bf, 32'hc0a98410} /* (29, 21, 5) {real, imag} */,
  {32'hc2150224, 32'h4155491c} /* (29, 21, 4) {real, imag} */,
  {32'hc23bf26b, 32'hc2a4e481} /* (29, 21, 3) {real, imag} */,
  {32'hc24e8c76, 32'hc24334b3} /* (29, 21, 2) {real, imag} */,
  {32'h42fa12d6, 32'h412b5500} /* (29, 21, 1) {real, imag} */,
  {32'h4211b222, 32'h4171d7c0} /* (29, 21, 0) {real, imag} */,
  {32'h41396734, 32'h425e7596} /* (29, 20, 31) {real, imag} */,
  {32'h41e83531, 32'h40338438} /* (29, 20, 30) {real, imag} */,
  {32'h40120fa8, 32'h4235a489} /* (29, 20, 29) {real, imag} */,
  {32'h42c8eef3, 32'hc04de800} /* (29, 20, 28) {real, imag} */,
  {32'hc286917c, 32'hc21f8de0} /* (29, 20, 27) {real, imag} */,
  {32'h3fbd9838, 32'hbf64c720} /* (29, 20, 26) {real, imag} */,
  {32'h4190e3af, 32'h4231611e} /* (29, 20, 25) {real, imag} */,
  {32'hc1c703ae, 32'h41bad1b5} /* (29, 20, 24) {real, imag} */,
  {32'h4023c2ce, 32'hc1c6adc6} /* (29, 20, 23) {real, imag} */,
  {32'h419981ef, 32'h414a317e} /* (29, 20, 22) {real, imag} */,
  {32'hc0ee0060, 32'hc17f0772} /* (29, 20, 21) {real, imag} */,
  {32'h40228de0, 32'hc238334c} /* (29, 20, 20) {real, imag} */,
  {32'h4003612c, 32'hc1469a32} /* (29, 20, 19) {real, imag} */,
  {32'h410b398a, 32'hbc752400} /* (29, 20, 18) {real, imag} */,
  {32'hc10bf942, 32'h3fcc3a78} /* (29, 20, 17) {real, imag} */,
  {32'h410c0ca4, 32'h415a8026} /* (29, 20, 16) {real, imag} */,
  {32'h417dedf6, 32'hc1cb082a} /* (29, 20, 15) {real, imag} */,
  {32'h40080dba, 32'h4060b44c} /* (29, 20, 14) {real, imag} */,
  {32'hc09b78f2, 32'h4213d1be} /* (29, 20, 13) {real, imag} */,
  {32'h415cc6a4, 32'h410441c0} /* (29, 20, 12) {real, imag} */,
  {32'h411bdf58, 32'hc1a1a365} /* (29, 20, 11) {real, imag} */,
  {32'hc10740f6, 32'hc0eb1c94} /* (29, 20, 10) {real, imag} */,
  {32'h411f6c2e, 32'hc1a91ce6} /* (29, 20, 9) {real, imag} */,
  {32'hc219ee7b, 32'h41b2fbcb} /* (29, 20, 8) {real, imag} */,
  {32'h40641cf2, 32'h413e7d90} /* (29, 20, 7) {real, imag} */,
  {32'h3ea43b80, 32'hc26dbe92} /* (29, 20, 6) {real, imag} */,
  {32'hc20d7132, 32'h4268b61a} /* (29, 20, 5) {real, imag} */,
  {32'hc1f1e924, 32'hc1ab2e68} /* (29, 20, 4) {real, imag} */,
  {32'hc22c2f9a, 32'h41c74696} /* (29, 20, 3) {real, imag} */,
  {32'h4243148a, 32'h42035dee} /* (29, 20, 2) {real, imag} */,
  {32'hbeb512f0, 32'hc1dcc26b} /* (29, 20, 1) {real, imag} */,
  {32'h40b96967, 32'hc11d3bc8} /* (29, 20, 0) {real, imag} */,
  {32'hc16f4dbc, 32'h41ebe85a} /* (29, 19, 31) {real, imag} */,
  {32'h428462ae, 32'h41eebb38} /* (29, 19, 30) {real, imag} */,
  {32'hc0b47044, 32'h3febd670} /* (29, 19, 29) {real, imag} */,
  {32'h41a1edb8, 32'hc23a414b} /* (29, 19, 28) {real, imag} */,
  {32'h41bab1ac, 32'h42304fca} /* (29, 19, 27) {real, imag} */,
  {32'hc1b7b730, 32'hc238687a} /* (29, 19, 26) {real, imag} */,
  {32'h41695c86, 32'hc19a929e} /* (29, 19, 25) {real, imag} */,
  {32'hc156f8d2, 32'h412c62ff} /* (29, 19, 24) {real, imag} */,
  {32'h40afec92, 32'h400b10a4} /* (29, 19, 23) {real, imag} */,
  {32'h41c246f8, 32'hc14c586f} /* (29, 19, 22) {real, imag} */,
  {32'hc1de2da7, 32'h41fcc16f} /* (29, 19, 21) {real, imag} */,
  {32'hc1afcb6c, 32'h40c25a14} /* (29, 19, 20) {real, imag} */,
  {32'h40ced592, 32'hc0e55c5d} /* (29, 19, 19) {real, imag} */,
  {32'h40d9d916, 32'hc053573c} /* (29, 19, 18) {real, imag} */,
  {32'hc056f0bc, 32'hc1596335} /* (29, 19, 17) {real, imag} */,
  {32'h40f0db4a, 32'hc1310cb4} /* (29, 19, 16) {real, imag} */,
  {32'h40d5701c, 32'h410e5495} /* (29, 19, 15) {real, imag} */,
  {32'hc09527ea, 32'h40034e04} /* (29, 19, 14) {real, imag} */,
  {32'hc176916b, 32'hc1a90857} /* (29, 19, 13) {real, imag} */,
  {32'hc162b714, 32'h4132f456} /* (29, 19, 12) {real, imag} */,
  {32'h418d752f, 32'hc0c1b39c} /* (29, 19, 11) {real, imag} */,
  {32'h4124e390, 32'h3fc19058} /* (29, 19, 10) {real, imag} */,
  {32'hc118861d, 32'hc196ab48} /* (29, 19, 9) {real, imag} */,
  {32'h41c45df1, 32'h410e4149} /* (29, 19, 8) {real, imag} */,
  {32'h41d626a3, 32'hc1511935} /* (29, 19, 7) {real, imag} */,
  {32'h425169ec, 32'h417c86ae} /* (29, 19, 6) {real, imag} */,
  {32'h40680950, 32'h40dc75ec} /* (29, 19, 5) {real, imag} */,
  {32'h4177eac5, 32'h418f5a0a} /* (29, 19, 4) {real, imag} */,
  {32'hc2023a9c, 32'hbfb8abf8} /* (29, 19, 3) {real, imag} */,
  {32'hc297a6c2, 32'hc127e60c} /* (29, 19, 2) {real, imag} */,
  {32'h41331ed4, 32'h4100da8d} /* (29, 19, 1) {real, imag} */,
  {32'hc1a83052, 32'hc212207f} /* (29, 19, 0) {real, imag} */,
  {32'h41b0cf88, 32'hc16be52e} /* (29, 18, 31) {real, imag} */,
  {32'hc28b8a44, 32'hc17c47fa} /* (29, 18, 30) {real, imag} */,
  {32'hc116552a, 32'h41bd0678} /* (29, 18, 29) {real, imag} */,
  {32'h41ae4b4b, 32'h4225ab92} /* (29, 18, 28) {real, imag} */,
  {32'hc251d2d0, 32'h420810b7} /* (29, 18, 27) {real, imag} */,
  {32'hc1376ab7, 32'h4236e5cf} /* (29, 18, 26) {real, imag} */,
  {32'hc10a7a09, 32'hc227c2cf} /* (29, 18, 25) {real, imag} */,
  {32'hc1456db2, 32'hc04add64} /* (29, 18, 24) {real, imag} */,
  {32'h41910ed2, 32'h40c75538} /* (29, 18, 23) {real, imag} */,
  {32'hbf861578, 32'hc1ef5290} /* (29, 18, 22) {real, imag} */,
  {32'hc0180bfa, 32'h414af27c} /* (29, 18, 21) {real, imag} */,
  {32'h400ace90, 32'h415e8bea} /* (29, 18, 20) {real, imag} */,
  {32'hc180ad16, 32'hc11f6a11} /* (29, 18, 19) {real, imag} */,
  {32'hc0ca0260, 32'h3fb6cf82} /* (29, 18, 18) {real, imag} */,
  {32'h40924bbc, 32'hc073414e} /* (29, 18, 17) {real, imag} */,
  {32'hc012eb52, 32'h409798ae} /* (29, 18, 16) {real, imag} */,
  {32'hc171396e, 32'h414bd9fe} /* (29, 18, 15) {real, imag} */,
  {32'hbff5a840, 32'h402a98a7} /* (29, 18, 14) {real, imag} */,
  {32'hc17edb84, 32'hc17b0a23} /* (29, 18, 13) {real, imag} */,
  {32'h41705754, 32'h3f4ba3f8} /* (29, 18, 12) {real, imag} */,
  {32'hbe1a6660, 32'hc1cb4818} /* (29, 18, 11) {real, imag} */,
  {32'h41c3de0a, 32'hc1063547} /* (29, 18, 10) {real, imag} */,
  {32'hc19bf01a, 32'hc1b0f807} /* (29, 18, 9) {real, imag} */,
  {32'h41e07071, 32'hc143ad2d} /* (29, 18, 8) {real, imag} */,
  {32'h41cba67c, 32'hc0eee748} /* (29, 18, 7) {real, imag} */,
  {32'h4148ac15, 32'h418adb1e} /* (29, 18, 6) {real, imag} */,
  {32'hc21e942c, 32'hc1799248} /* (29, 18, 5) {real, imag} */,
  {32'h418eb679, 32'h4181c231} /* (29, 18, 4) {real, imag} */,
  {32'hc0ccb23c, 32'h4106d499} /* (29, 18, 3) {real, imag} */,
  {32'hc235f922, 32'hc1c70217} /* (29, 18, 2) {real, imag} */,
  {32'h426bf1d0, 32'hc194f8ff} /* (29, 18, 1) {real, imag} */,
  {32'h412e4c7e, 32'h41754f6b} /* (29, 18, 0) {real, imag} */,
  {32'hc21bc6f6, 32'hc1e22126} /* (29, 17, 31) {real, imag} */,
  {32'h42cc239c, 32'hc1ba47f5} /* (29, 17, 30) {real, imag} */,
  {32'h3f085870, 32'hc1c00865} /* (29, 17, 29) {real, imag} */,
  {32'hc1370e89, 32'h41fba4ad} /* (29, 17, 28) {real, imag} */,
  {32'hc21e3a2e, 32'hc1d8efd7} /* (29, 17, 27) {real, imag} */,
  {32'h4193803a, 32'h402bc7e8} /* (29, 17, 26) {real, imag} */,
  {32'hc14f053f, 32'h414ab3ca} /* (29, 17, 25) {real, imag} */,
  {32'hc189de38, 32'hbfefaa58} /* (29, 17, 24) {real, imag} */,
  {32'h408459ad, 32'hc1965a47} /* (29, 17, 23) {real, imag} */,
  {32'hc119e5e2, 32'h40af48ac} /* (29, 17, 22) {real, imag} */,
  {32'h3fa28b28, 32'hc1f11a5b} /* (29, 17, 21) {real, imag} */,
  {32'h40d870d1, 32'h3f93ccb4} /* (29, 17, 20) {real, imag} */,
  {32'h411581d7, 32'h411bb4a1} /* (29, 17, 19) {real, imag} */,
  {32'h3f5cc040, 32'hc12472a0} /* (29, 17, 18) {real, imag} */,
  {32'h4037888a, 32'h401b6bef} /* (29, 17, 17) {real, imag} */,
  {32'hc117df17, 32'hc0434fa4} /* (29, 17, 16) {real, imag} */,
  {32'h40e70ac3, 32'hc077a49f} /* (29, 17, 15) {real, imag} */,
  {32'hc03e6330, 32'hc1187eea} /* (29, 17, 14) {real, imag} */,
  {32'hc12112b7, 32'hbfc5ae18} /* (29, 17, 13) {real, imag} */,
  {32'hc0aad153, 32'h4173c3ae} /* (29, 17, 12) {real, imag} */,
  {32'h41a4fefc, 32'h407934d8} /* (29, 17, 11) {real, imag} */,
  {32'hc2376fa4, 32'h41dac151} /* (29, 17, 10) {real, imag} */,
  {32'h40cda0d1, 32'h41280d06} /* (29, 17, 9) {real, imag} */,
  {32'hc1a5128c, 32'hc118aa35} /* (29, 17, 8) {real, imag} */,
  {32'hc04aad64, 32'hc1cdfab9} /* (29, 17, 7) {real, imag} */,
  {32'hc1daa758, 32'h419a75af} /* (29, 17, 6) {real, imag} */,
  {32'h401c06c8, 32'hbfcee030} /* (29, 17, 5) {real, imag} */,
  {32'hc18e27d9, 32'hc1061f1e} /* (29, 17, 4) {real, imag} */,
  {32'hc1ba49de, 32'hc19c4b9f} /* (29, 17, 3) {real, imag} */,
  {32'h428296a8, 32'hc1868343} /* (29, 17, 2) {real, imag} */,
  {32'hc205c3d2, 32'hc19d4324} /* (29, 17, 1) {real, imag} */,
  {32'hbf902698, 32'hc1600a85} /* (29, 17, 0) {real, imag} */,
  {32'hc0b43ffc, 32'h41c12f97} /* (29, 16, 31) {real, imag} */,
  {32'h419d2c51, 32'h4122a35e} /* (29, 16, 30) {real, imag} */,
  {32'hc20e4236, 32'hc14a1a5d} /* (29, 16, 29) {real, imag} */,
  {32'hc1e98968, 32'h421179a6} /* (29, 16, 28) {real, imag} */,
  {32'h40b545aa, 32'hc17ac034} /* (29, 16, 27) {real, imag} */,
  {32'h402f0676, 32'hc184355a} /* (29, 16, 26) {real, imag} */,
  {32'hc17075b8, 32'h40fc8bc4} /* (29, 16, 25) {real, imag} */,
  {32'h416bbcce, 32'h41538ad8} /* (29, 16, 24) {real, imag} */,
  {32'h403f123f, 32'h4007e4d2} /* (29, 16, 23) {real, imag} */,
  {32'hbf086600, 32'h40481378} /* (29, 16, 22) {real, imag} */,
  {32'hc1eeed08, 32'hc08856d8} /* (29, 16, 21) {real, imag} */,
  {32'hc139331e, 32'hc081cc74} /* (29, 16, 20) {real, imag} */,
  {32'hc0d158ba, 32'hc0d528c2} /* (29, 16, 19) {real, imag} */,
  {32'h40f5b383, 32'h411ea877} /* (29, 16, 18) {real, imag} */,
  {32'h413ffe27, 32'h3fd35518} /* (29, 16, 17) {real, imag} */,
  {32'h3fd1a9c8, 32'h405c7700} /* (29, 16, 16) {real, imag} */,
  {32'hbffacd48, 32'h403ed0c0} /* (29, 16, 15) {real, imag} */,
  {32'h4122937e, 32'hc0ae75e4} /* (29, 16, 14) {real, imag} */,
  {32'h40333a05, 32'hc0ba6856} /* (29, 16, 13) {real, imag} */,
  {32'hc0856fe5, 32'hc129079e} /* (29, 16, 12) {real, imag} */,
  {32'hc0e6fa9a, 32'h4111ab0c} /* (29, 16, 11) {real, imag} */,
  {32'hc125e91a, 32'hc1a2c417} /* (29, 16, 10) {real, imag} */,
  {32'h40886756, 32'hc0cb3669} /* (29, 16, 9) {real, imag} */,
  {32'h41fba7bf, 32'h41be59d0} /* (29, 16, 8) {real, imag} */,
  {32'hc1aebb2a, 32'hc1b31b3b} /* (29, 16, 7) {real, imag} */,
  {32'h4072a92a, 32'h4178a9f9} /* (29, 16, 6) {real, imag} */,
  {32'h414fe293, 32'h416d7850} /* (29, 16, 5) {real, imag} */,
  {32'h411c1ec0, 32'h400c4d38} /* (29, 16, 4) {real, imag} */,
  {32'h41eb0303, 32'hc22e40de} /* (29, 16, 3) {real, imag} */,
  {32'h40d90fac, 32'h3f128988} /* (29, 16, 2) {real, imag} */,
  {32'hc0af30b4, 32'h403c0a68} /* (29, 16, 1) {real, imag} */,
  {32'h41b74be6, 32'h423e92b2} /* (29, 16, 0) {real, imag} */,
  {32'h42a17b80, 32'h42277b2c} /* (29, 15, 31) {real, imag} */,
  {32'hc194af8a, 32'hc11fccb0} /* (29, 15, 30) {real, imag} */,
  {32'hc2808cc0, 32'hc1cee3a7} /* (29, 15, 29) {real, imag} */,
  {32'hc16145fe, 32'h40dc6f14} /* (29, 15, 28) {real, imag} */,
  {32'h41edb577, 32'h3fb3cbb0} /* (29, 15, 27) {real, imag} */,
  {32'h41943d4e, 32'h40061612} /* (29, 15, 26) {real, imag} */,
  {32'h41accfe0, 32'h3fcddd10} /* (29, 15, 25) {real, imag} */,
  {32'h419acc97, 32'hbf9c1128} /* (29, 15, 24) {real, imag} */,
  {32'h417e315c, 32'h408134fc} /* (29, 15, 23) {real, imag} */,
  {32'h4173307e, 32'h4148ef36} /* (29, 15, 22) {real, imag} */,
  {32'hc12c9d4b, 32'h41a118b5} /* (29, 15, 21) {real, imag} */,
  {32'hc1381afd, 32'hc196bb42} /* (29, 15, 20) {real, imag} */,
  {32'hc1547d2c, 32'hc18ef485} /* (29, 15, 19) {real, imag} */,
  {32'hc11b413a, 32'hc1013485} /* (29, 15, 18) {real, imag} */,
  {32'h40a68d4c, 32'hc0bb8be6} /* (29, 15, 17) {real, imag} */,
  {32'hc158cf85, 32'hbfc61e60} /* (29, 15, 16) {real, imag} */,
  {32'hc064c2f8, 32'hbfb26c18} /* (29, 15, 15) {real, imag} */,
  {32'hbcf44300, 32'h41904980} /* (29, 15, 14) {real, imag} */,
  {32'h3f2f2a00, 32'hc037837a} /* (29, 15, 13) {real, imag} */,
  {32'hc0caa182, 32'h40a21812} /* (29, 15, 12) {real, imag} */,
  {32'hbce35200, 32'h3fb9c150} /* (29, 15, 11) {real, imag} */,
  {32'hc1822c33, 32'hc16544aa} /* (29, 15, 10) {real, imag} */,
  {32'h405702ae, 32'h41872b81} /* (29, 15, 9) {real, imag} */,
  {32'hc15cde8a, 32'h419dec32} /* (29, 15, 8) {real, imag} */,
  {32'h418d532c, 32'h412d16ea} /* (29, 15, 7) {real, imag} */,
  {32'hc1001d20, 32'h417f6dbc} /* (29, 15, 6) {real, imag} */,
  {32'h4196c9f7, 32'hc1a85aa9} /* (29, 15, 5) {real, imag} */,
  {32'hc0950918, 32'h421799a4} /* (29, 15, 4) {real, imag} */,
  {32'hc17a73ae, 32'hc1275e32} /* (29, 15, 3) {real, imag} */,
  {32'hc189cdca, 32'hc13bd64e} /* (29, 15, 2) {real, imag} */,
  {32'h4182b63e, 32'hc1926500} /* (29, 15, 1) {real, imag} */,
  {32'hc2337e84, 32'hc1b18582} /* (29, 15, 0) {real, imag} */,
  {32'hc29e17f7, 32'h42428931} /* (29, 14, 31) {real, imag} */,
  {32'hc0dd0cc3, 32'hc2843c23} /* (29, 14, 30) {real, imag} */,
  {32'hc215aad1, 32'h4159017d} /* (29, 14, 29) {real, imag} */,
  {32'hc0841acc, 32'h41dbcd59} /* (29, 14, 28) {real, imag} */,
  {32'hbf141120, 32'hc0052af6} /* (29, 14, 27) {real, imag} */,
  {32'hc1b13a19, 32'hc028782a} /* (29, 14, 26) {real, imag} */,
  {32'h421feaac, 32'hc175da48} /* (29, 14, 25) {real, imag} */,
  {32'hc170f6b2, 32'hc246ecd2} /* (29, 14, 24) {real, imag} */,
  {32'h40f83344, 32'h41828025} /* (29, 14, 23) {real, imag} */,
  {32'h4116a772, 32'h419dfb7b} /* (29, 14, 22) {real, imag} */,
  {32'hc20ae42e, 32'h408f1050} /* (29, 14, 21) {real, imag} */,
  {32'hc0090b70, 32'h40a9df88} /* (29, 14, 20) {real, imag} */,
  {32'h41299ee2, 32'h4126a845} /* (29, 14, 19) {real, imag} */,
  {32'hc09bcb85, 32'h411176da} /* (29, 14, 18) {real, imag} */,
  {32'h40053f00, 32'h40b6b553} /* (29, 14, 17) {real, imag} */,
  {32'h413edba2, 32'h3ffc3de8} /* (29, 14, 16) {real, imag} */,
  {32'hc0b80e40, 32'h40b6b443} /* (29, 14, 15) {real, imag} */,
  {32'hc10f1944, 32'hc11a1a36} /* (29, 14, 14) {real, imag} */,
  {32'h414c26d4, 32'h4129770d} /* (29, 14, 13) {real, imag} */,
  {32'h413c64ec, 32'hc109d70a} /* (29, 14, 12) {real, imag} */,
  {32'h40da0040, 32'h41f6ff7c} /* (29, 14, 11) {real, imag} */,
  {32'h418a5067, 32'h41e6c589} /* (29, 14, 10) {real, imag} */,
  {32'hc24a3b22, 32'h4151a126} /* (29, 14, 9) {real, imag} */,
  {32'h421ffa6e, 32'hc10d7e40} /* (29, 14, 8) {real, imag} */,
  {32'h41901fbb, 32'h411ac518} /* (29, 14, 7) {real, imag} */,
  {32'hc0d6acbd, 32'h411db2c6} /* (29, 14, 6) {real, imag} */,
  {32'h420c26c6, 32'h3fd8433c} /* (29, 14, 5) {real, imag} */,
  {32'hc1dcd7e9, 32'h408277b8} /* (29, 14, 4) {real, imag} */,
  {32'hc11af6f4, 32'h4187687d} /* (29, 14, 3) {real, imag} */,
  {32'hc1060c31, 32'hc213f6f2} /* (29, 14, 2) {real, imag} */,
  {32'hc2592f62, 32'hc14525b0} /* (29, 14, 1) {real, imag} */,
  {32'hc28da347, 32'hc1964cbe} /* (29, 14, 0) {real, imag} */,
  {32'h42a66380, 32'hc23b228e} /* (29, 13, 31) {real, imag} */,
  {32'h40b77220, 32'h41880d4b} /* (29, 13, 30) {real, imag} */,
  {32'h4210456b, 32'h41c0fdfe} /* (29, 13, 29) {real, imag} */,
  {32'hc20550ac, 32'h41747700} /* (29, 13, 28) {real, imag} */,
  {32'hc0b7e9b4, 32'hc1ebdb76} /* (29, 13, 27) {real, imag} */,
  {32'hc1817b96, 32'hc1f4c927} /* (29, 13, 26) {real, imag} */,
  {32'hc18a5c5a, 32'h4164b474} /* (29, 13, 25) {real, imag} */,
  {32'hbff03200, 32'h419b8eeb} /* (29, 13, 24) {real, imag} */,
  {32'h42561cfd, 32'hc2095707} /* (29, 13, 23) {real, imag} */,
  {32'hc1a60419, 32'h4112f10a} /* (29, 13, 22) {real, imag} */,
  {32'hc12c6a38, 32'hc1c04750} /* (29, 13, 21) {real, imag} */,
  {32'hc12e40b4, 32'h40830360} /* (29, 13, 20) {real, imag} */,
  {32'hc0726c8e, 32'hc1a13f5b} /* (29, 13, 19) {real, imag} */,
  {32'h40d9bfea, 32'hc0317d1c} /* (29, 13, 18) {real, imag} */,
  {32'hbfd2abd0, 32'hc069dc7c} /* (29, 13, 17) {real, imag} */,
  {32'hbf19d340, 32'hc13a8abe} /* (29, 13, 16) {real, imag} */,
  {32'hc0f41ebc, 32'hc093ef56} /* (29, 13, 15) {real, imag} */,
  {32'hc0b9f1de, 32'hc0728a08} /* (29, 13, 14) {real, imag} */,
  {32'hc0105586, 32'hc16a14c6} /* (29, 13, 13) {real, imag} */,
  {32'hc17de3f4, 32'hbfdfb93a} /* (29, 13, 12) {real, imag} */,
  {32'hbf01bcf8, 32'h3fd34230} /* (29, 13, 11) {real, imag} */,
  {32'hc138b466, 32'hc11a1ff6} /* (29, 13, 10) {real, imag} */,
  {32'h41d2703e, 32'h420fc7c1} /* (29, 13, 9) {real, imag} */,
  {32'hc22cc102, 32'hc2606242} /* (29, 13, 8) {real, imag} */,
  {32'h40b4b850, 32'h419694b2} /* (29, 13, 7) {real, imag} */,
  {32'h41573000, 32'hc1bcb2bb} /* (29, 13, 6) {real, imag} */,
  {32'hc18de877, 32'hc0e7bb96} /* (29, 13, 5) {real, imag} */,
  {32'hc18ebc2c, 32'hc0842240} /* (29, 13, 4) {real, imag} */,
  {32'hc1b08511, 32'hc23a78f5} /* (29, 13, 3) {real, imag} */,
  {32'hc28caf72, 32'h41954501} /* (29, 13, 2) {real, imag} */,
  {32'hc0aee6d8, 32'h4095839c} /* (29, 13, 1) {real, imag} */,
  {32'hc1aa9dca, 32'hc209b4c2} /* (29, 13, 0) {real, imag} */,
  {32'hc275ba97, 32'hc282e989} /* (29, 12, 31) {real, imag} */,
  {32'hc2679357, 32'hc2160d4b} /* (29, 12, 30) {real, imag} */,
  {32'h42cbb245, 32'h42299bc2} /* (29, 12, 29) {real, imag} */,
  {32'h4152f407, 32'h41042d13} /* (29, 12, 28) {real, imag} */,
  {32'hbe166f00, 32'h40f3433e} /* (29, 12, 27) {real, imag} */,
  {32'hc0f5f32a, 32'h4155240e} /* (29, 12, 26) {real, imag} */,
  {32'h4287c204, 32'h41e62e40} /* (29, 12, 25) {real, imag} */,
  {32'h3f1fc740, 32'hc11ac4d3} /* (29, 12, 24) {real, imag} */,
  {32'h41249dfa, 32'h424daae6} /* (29, 12, 23) {real, imag} */,
  {32'hbf6c63c0, 32'h410e7468} /* (29, 12, 22) {real, imag} */,
  {32'h4159db49, 32'h4192ba30} /* (29, 12, 21) {real, imag} */,
  {32'h40956592, 32'h400aed1c} /* (29, 12, 20) {real, imag} */,
  {32'hc1d9960f, 32'h41ad5c78} /* (29, 12, 19) {real, imag} */,
  {32'h40b6adb4, 32'hc0d589d5} /* (29, 12, 18) {real, imag} */,
  {32'h3fc41ee8, 32'hc12d4dfe} /* (29, 12, 17) {real, imag} */,
  {32'h3f2994a0, 32'h401d9470} /* (29, 12, 16) {real, imag} */,
  {32'h3f74aed0, 32'hc19e8ed8} /* (29, 12, 15) {real, imag} */,
  {32'h40748478, 32'h4159223a} /* (29, 12, 14) {real, imag} */,
  {32'hc11cbc82, 32'h418fb57a} /* (29, 12, 13) {real, imag} */,
  {32'h4178b58d, 32'h41c53978} /* (29, 12, 12) {real, imag} */,
  {32'hc19bbc1c, 32'h404ed0bc} /* (29, 12, 11) {real, imag} */,
  {32'h41f453cb, 32'h3fd9dd04} /* (29, 12, 10) {real, imag} */,
  {32'h3f2c1e20, 32'hbf1ca020} /* (29, 12, 9) {real, imag} */,
  {32'h42417d35, 32'hc0292ebc} /* (29, 12, 8) {real, imag} */,
  {32'hc2d8ca08, 32'h42495334} /* (29, 12, 7) {real, imag} */,
  {32'h41cb6b9e, 32'hc117bdac} /* (29, 12, 6) {real, imag} */,
  {32'h420bb7e3, 32'h415c4991} /* (29, 12, 5) {real, imag} */,
  {32'h4141555f, 32'hc19a2bc2} /* (29, 12, 4) {real, imag} */,
  {32'hbe635e00, 32'hc174aa9a} /* (29, 12, 3) {real, imag} */,
  {32'h411cf7e4, 32'h424fb951} /* (29, 12, 2) {real, imag} */,
  {32'h415f142c, 32'hc1da0870} /* (29, 12, 1) {real, imag} */,
  {32'h423c8df4, 32'h42140b69} /* (29, 12, 0) {real, imag} */,
  {32'hc1ee0242, 32'h4218340d} /* (29, 11, 31) {real, imag} */,
  {32'h42634094, 32'hc2f53af5} /* (29, 11, 30) {real, imag} */,
  {32'h40f84228, 32'hc1b9b21c} /* (29, 11, 29) {real, imag} */,
  {32'hc29b5269, 32'hc29318c2} /* (29, 11, 28) {real, imag} */,
  {32'h4256309a, 32'h42149e23} /* (29, 11, 27) {real, imag} */,
  {32'hc1eff2ea, 32'h423d41b4} /* (29, 11, 26) {real, imag} */,
  {32'hc25d5aa3, 32'h422c7b75} /* (29, 11, 25) {real, imag} */,
  {32'h4238f2d2, 32'h42604cc0} /* (29, 11, 24) {real, imag} */,
  {32'h40704060, 32'h421106ba} /* (29, 11, 23) {real, imag} */,
  {32'h417859ce, 32'h415237ea} /* (29, 11, 22) {real, imag} */,
  {32'hc129a446, 32'hc212d836} /* (29, 11, 21) {real, imag} */,
  {32'h412e2100, 32'hc12afede} /* (29, 11, 20) {real, imag} */,
  {32'hc16a7b7a, 32'hc0925aea} /* (29, 11, 19) {real, imag} */,
  {32'hc1c82bd0, 32'hc0cd52dc} /* (29, 11, 18) {real, imag} */,
  {32'h412d5b48, 32'h41919e0f} /* (29, 11, 17) {real, imag} */,
  {32'h3f9de3e0, 32'hbee62900} /* (29, 11, 16) {real, imag} */,
  {32'hc0ec3d20, 32'hc16de1ae} /* (29, 11, 15) {real, imag} */,
  {32'hc204bfde, 32'h41a6a20b} /* (29, 11, 14) {real, imag} */,
  {32'h419ae9fb, 32'h40aba20a} /* (29, 11, 13) {real, imag} */,
  {32'hc08ddfe1, 32'h41f884e9} /* (29, 11, 12) {real, imag} */,
  {32'hc1d52a7d, 32'hbff7f640} /* (29, 11, 11) {real, imag} */,
  {32'h42080c22, 32'hc0996903} /* (29, 11, 10) {real, imag} */,
  {32'h4129fa38, 32'hc1b35a3c} /* (29, 11, 9) {real, imag} */,
  {32'hbf1e3700, 32'h40fde0dc} /* (29, 11, 8) {real, imag} */,
  {32'hc06b9e70, 32'h4151321b} /* (29, 11, 7) {real, imag} */,
  {32'h425c4067, 32'hc2861f04} /* (29, 11, 6) {real, imag} */,
  {32'hc210d74a, 32'h420b5067} /* (29, 11, 5) {real, imag} */,
  {32'h4287bb99, 32'hc0d5f778} /* (29, 11, 4) {real, imag} */,
  {32'h42b4224c, 32'hc102b159} /* (29, 11, 3) {real, imag} */,
  {32'h42950fb2, 32'hc2068f4e} /* (29, 11, 2) {real, imag} */,
  {32'hc2b8e774, 32'h423f7807} /* (29, 11, 1) {real, imag} */,
  {32'hc2b762d6, 32'h425f2424} /* (29, 11, 0) {real, imag} */,
  {32'h42c817ba, 32'hc23a4dc8} /* (29, 10, 31) {real, imag} */,
  {32'hc31ec78c, 32'h42fbe1ff} /* (29, 10, 30) {real, imag} */,
  {32'hbf584d80, 32'hc29075dc} /* (29, 10, 29) {real, imag} */,
  {32'h4235e2de, 32'hc3235727} /* (29, 10, 28) {real, imag} */,
  {32'hc2ac7088, 32'hc1b7fd9a} /* (29, 10, 27) {real, imag} */,
  {32'hc0bb8568, 32'h4143454e} /* (29, 10, 26) {real, imag} */,
  {32'hc2db9f34, 32'hc0db5ea6} /* (29, 10, 25) {real, imag} */,
  {32'h424bd0aa, 32'h416ea763} /* (29, 10, 24) {real, imag} */,
  {32'hc1b9da56, 32'h4115c860} /* (29, 10, 23) {real, imag} */,
  {32'hc116a544, 32'hc1b643f5} /* (29, 10, 22) {real, imag} */,
  {32'h424fba9a, 32'h41931ffc} /* (29, 10, 21) {real, imag} */,
  {32'hbff07ad8, 32'hc1a66749} /* (29, 10, 20) {real, imag} */,
  {32'hc15b5dfe, 32'h3e233180} /* (29, 10, 19) {real, imag} */,
  {32'hc20cc029, 32'hc19fa615} /* (29, 10, 18) {real, imag} */,
  {32'hc1054ade, 32'h3fdde958} /* (29, 10, 17) {real, imag} */,
  {32'hc1897b5c, 32'hc068cd00} /* (29, 10, 16) {real, imag} */,
  {32'hc11b3326, 32'h410f4595} /* (29, 10, 15) {real, imag} */,
  {32'h417d609c, 32'hc1915d0f} /* (29, 10, 14) {real, imag} */,
  {32'h420a354c, 32'h424c9b4e} /* (29, 10, 13) {real, imag} */,
  {32'hc0b4d242, 32'hc1b12439} /* (29, 10, 12) {real, imag} */,
  {32'hc1039e86, 32'hc1ecb538} /* (29, 10, 11) {real, imag} */,
  {32'h41d7238e, 32'h404a8508} /* (29, 10, 10) {real, imag} */,
  {32'h420e9fcf, 32'h4270bd0c} /* (29, 10, 9) {real, imag} */,
  {32'h41067ca8, 32'hc2046cd7} /* (29, 10, 8) {real, imag} */,
  {32'hc2910626, 32'h419fb762} /* (29, 10, 7) {real, imag} */,
  {32'hc24e9e8b, 32'hc0dbfeac} /* (29, 10, 6) {real, imag} */,
  {32'hc26fcb39, 32'h42622a63} /* (29, 10, 5) {real, imag} */,
  {32'hc165ca9e, 32'h42eafa26} /* (29, 10, 4) {real, imag} */,
  {32'h43193ed6, 32'h42c2956e} /* (29, 10, 3) {real, imag} */,
  {32'h42b70c3c, 32'h40a186d0} /* (29, 10, 2) {real, imag} */,
  {32'hc232449c, 32'h40f6292c} /* (29, 10, 1) {real, imag} */,
  {32'h42849f61, 32'hc278072a} /* (29, 10, 0) {real, imag} */,
  {32'h43388caf, 32'h429c9c56} /* (29, 9, 31) {real, imag} */,
  {32'hc24a2376, 32'h4205b718} /* (29, 9, 30) {real, imag} */,
  {32'h4237e092, 32'hc183dd1c} /* (29, 9, 29) {real, imag} */,
  {32'h426d8282, 32'h42185003} /* (29, 9, 28) {real, imag} */,
  {32'hc2e693d0, 32'h424a8502} /* (29, 9, 27) {real, imag} */,
  {32'h41848122, 32'h423ccd06} /* (29, 9, 26) {real, imag} */,
  {32'h40166744, 32'h40cb49e8} /* (29, 9, 25) {real, imag} */,
  {32'hc22bd04e, 32'hc0061c90} /* (29, 9, 24) {real, imag} */,
  {32'h425035ee, 32'h412b1165} /* (29, 9, 23) {real, imag} */,
  {32'hc1be23cc, 32'h4092a084} /* (29, 9, 22) {real, imag} */,
  {32'hc204fa0d, 32'h41a342cb} /* (29, 9, 21) {real, imag} */,
  {32'hbf9dcd68, 32'hc24335f8} /* (29, 9, 20) {real, imag} */,
  {32'h425de838, 32'h41d0cecf} /* (29, 9, 19) {real, imag} */,
  {32'hc0dd0820, 32'h415677b4} /* (29, 9, 18) {real, imag} */,
  {32'h414c947a, 32'hc22308e2} /* (29, 9, 17) {real, imag} */,
  {32'h40802860, 32'hc19c67ee} /* (29, 9, 16) {real, imag} */,
  {32'h420a37da, 32'hc0fa0df0} /* (29, 9, 15) {real, imag} */,
  {32'h413ed22e, 32'hc1acef00} /* (29, 9, 14) {real, imag} */,
  {32'hc1d4bf80, 32'hc1720502} /* (29, 9, 13) {real, imag} */,
  {32'h3e64adc0, 32'hc217f69c} /* (29, 9, 12) {real, imag} */,
  {32'hc1214a9c, 32'hc20e380c} /* (29, 9, 11) {real, imag} */,
  {32'h420a9b88, 32'h41d610bf} /* (29, 9, 10) {real, imag} */,
  {32'h40ea1370, 32'hbf51edb0} /* (29, 9, 9) {real, imag} */,
  {32'hc2644dc6, 32'h420fefb0} /* (29, 9, 8) {real, imag} */,
  {32'hc1d013f0, 32'hc28df7a0} /* (29, 9, 7) {real, imag} */,
  {32'hc27e768d, 32'hc13dca92} /* (29, 9, 6) {real, imag} */,
  {32'h42578040, 32'hc132cd32} /* (29, 9, 5) {real, imag} */,
  {32'hc240add6, 32'h4191f6cc} /* (29, 9, 4) {real, imag} */,
  {32'hc10562c8, 32'hbf0fccd0} /* (29, 9, 3) {real, imag} */,
  {32'hbfac9b80, 32'h42857be4} /* (29, 9, 2) {real, imag} */,
  {32'hc297e79a, 32'hc2a59518} /* (29, 9, 1) {real, imag} */,
  {32'h42258dbf, 32'hc25fe889} /* (29, 9, 0) {real, imag} */,
  {32'h418d1e08, 32'h438ab418} /* (29, 8, 31) {real, imag} */,
  {32'h418df328, 32'hc3666a17} /* (29, 8, 30) {real, imag} */,
  {32'hc33af478, 32'hc1bd16fe} /* (29, 8, 29) {real, imag} */,
  {32'h42b4b4a2, 32'h4247a290} /* (29, 8, 28) {real, imag} */,
  {32'hc2625e7e, 32'h42b82c5e} /* (29, 8, 27) {real, imag} */,
  {32'hc12b25b0, 32'h4202ade4} /* (29, 8, 26) {real, imag} */,
  {32'h4184e67a, 32'h4285a0af} /* (29, 8, 25) {real, imag} */,
  {32'hc27cb637, 32'h414aeeae} /* (29, 8, 24) {real, imag} */,
  {32'h41aeff89, 32'h42e89dc2} /* (29, 8, 23) {real, imag} */,
  {32'h420b67e4, 32'hc1429254} /* (29, 8, 22) {real, imag} */,
  {32'hc14a178c, 32'h422ca752} /* (29, 8, 21) {real, imag} */,
  {32'hc1abd35e, 32'h414f728b} /* (29, 8, 20) {real, imag} */,
  {32'h417a5bf8, 32'hc1c4ac58} /* (29, 8, 19) {real, imag} */,
  {32'h40c53c54, 32'hc145cd1c} /* (29, 8, 18) {real, imag} */,
  {32'h41caac78, 32'h40e43ec8} /* (29, 8, 17) {real, imag} */,
  {32'hc0ddf216, 32'hc09873b8} /* (29, 8, 16) {real, imag} */,
  {32'hc24bbbda, 32'h40a8d478} /* (29, 8, 15) {real, imag} */,
  {32'h4159a48a, 32'hc19185d6} /* (29, 8, 14) {real, imag} */,
  {32'hc215f490, 32'hc10874d1} /* (29, 8, 13) {real, imag} */,
  {32'hbfdbb580, 32'hc203720d} /* (29, 8, 12) {real, imag} */,
  {32'h42bb758e, 32'hc1a6649c} /* (29, 8, 11) {real, imag} */,
  {32'hc1463556, 32'h42c42f08} /* (29, 8, 10) {real, imag} */,
  {32'hc28a41fd, 32'hc214b17b} /* (29, 8, 9) {real, imag} */,
  {32'h4230a6bf, 32'h423a5244} /* (29, 8, 8) {real, imag} */,
  {32'h42b74bbe, 32'h423288d4} /* (29, 8, 7) {real, imag} */,
  {32'h42b5dad0, 32'h420d4bfe} /* (29, 8, 6) {real, imag} */,
  {32'h41331e4e, 32'hc3139231} /* (29, 8, 5) {real, imag} */,
  {32'hc1d981c1, 32'hc20cc7f4} /* (29, 8, 4) {real, imag} */,
  {32'h428dd0b8, 32'hc2cb8a1c} /* (29, 8, 3) {real, imag} */,
  {32'h42b02dba, 32'h426bdbd4} /* (29, 8, 2) {real, imag} */,
  {32'hc3128969, 32'h430a31a7} /* (29, 8, 1) {real, imag} */,
  {32'hbf8267b8, 32'h42d93bd0} /* (29, 8, 0) {real, imag} */,
  {32'h41e4c4c4, 32'hc2decd05} /* (29, 7, 31) {real, imag} */,
  {32'h4059aba0, 32'hc22159bb} /* (29, 7, 30) {real, imag} */,
  {32'h42e4fcf0, 32'h42a13a6c} /* (29, 7, 29) {real, imag} */,
  {32'h430aed18, 32'h42d6cd04} /* (29, 7, 28) {real, imag} */,
  {32'hc2639814, 32'hc23f6420} /* (29, 7, 27) {real, imag} */,
  {32'h41bf36a4, 32'h42223e90} /* (29, 7, 26) {real, imag} */,
  {32'h4158a14e, 32'h431122f2} /* (29, 7, 25) {real, imag} */,
  {32'hc13b918f, 32'h420cc103} /* (29, 7, 24) {real, imag} */,
  {32'hc1d08f05, 32'hc1d67b6c} /* (29, 7, 23) {real, imag} */,
  {32'hc22f05ad, 32'h41ac0b42} /* (29, 7, 22) {real, imag} */,
  {32'h41dbefbc, 32'hc23da241} /* (29, 7, 21) {real, imag} */,
  {32'h40287778, 32'h42819a86} /* (29, 7, 20) {real, imag} */,
  {32'h41ae0fb2, 32'hc11e18cc} /* (29, 7, 19) {real, imag} */,
  {32'hc1a43fc4, 32'hc1ad5425} /* (29, 7, 18) {real, imag} */,
  {32'hc0b14560, 32'h42422016} /* (29, 7, 17) {real, imag} */,
  {32'hc21510c5, 32'hc18836d0} /* (29, 7, 16) {real, imag} */,
  {32'h417f7af0, 32'h41bf5091} /* (29, 7, 15) {real, imag} */,
  {32'hc0faef70, 32'h40f654bc} /* (29, 7, 14) {real, imag} */,
  {32'h41354234, 32'h42086c03} /* (29, 7, 13) {real, imag} */,
  {32'hc1a084bb, 32'hc1da4da6} /* (29, 7, 12) {real, imag} */,
  {32'h42065ef2, 32'h418ba666} /* (29, 7, 11) {real, imag} */,
  {32'hc25d0e95, 32'hc24815d9} /* (29, 7, 10) {real, imag} */,
  {32'h421fffe0, 32'hc233d37e} /* (29, 7, 9) {real, imag} */,
  {32'h41b3f990, 32'h43152804} /* (29, 7, 8) {real, imag} */,
  {32'hc20930ea, 32'h4181bfb0} /* (29, 7, 7) {real, imag} */,
  {32'hc29e5214, 32'hc254c0d6} /* (29, 7, 6) {real, imag} */,
  {32'hc2b011ea, 32'hc230ef1a} /* (29, 7, 5) {real, imag} */,
  {32'h426199da, 32'hc2ad6164} /* (29, 7, 4) {real, imag} */,
  {32'h41fb7850, 32'h42702370} /* (29, 7, 3) {real, imag} */,
  {32'hc323fd6e, 32'hc28ab052} /* (29, 7, 2) {real, imag} */,
  {32'h42f87b13, 32'hc3330bb2} /* (29, 7, 1) {real, imag} */,
  {32'h42444c45, 32'hc344d689} /* (29, 7, 0) {real, imag} */,
  {32'h420cee83, 32'h41c69302} /* (29, 6, 31) {real, imag} */,
  {32'h41fbbe17, 32'h41b28af6} /* (29, 6, 30) {real, imag} */,
  {32'h42cad4e3, 32'h42044557} /* (29, 6, 29) {real, imag} */,
  {32'h425f7566, 32'hc2c1bc8b} /* (29, 6, 28) {real, imag} */,
  {32'h42731ee9, 32'hc1f67b6b} /* (29, 6, 27) {real, imag} */,
  {32'hc21f225c, 32'hc113d9f0} /* (29, 6, 26) {real, imag} */,
  {32'h428587df, 32'hc30383bb} /* (29, 6, 25) {real, imag} */,
  {32'hc214b644, 32'h4198993b} /* (29, 6, 24) {real, imag} */,
  {32'hc1af90d4, 32'h41256f98} /* (29, 6, 23) {real, imag} */,
  {32'hc05981f2, 32'hc2ae0626} /* (29, 6, 22) {real, imag} */,
  {32'h4120ab62, 32'hc15c8748} /* (29, 6, 21) {real, imag} */,
  {32'hc197c56d, 32'h41d7df98} /* (29, 6, 20) {real, imag} */,
  {32'hc232d10f, 32'h42774e1b} /* (29, 6, 19) {real, imag} */,
  {32'h41d4e705, 32'h41096a5d} /* (29, 6, 18) {real, imag} */,
  {32'h42093aa3, 32'h41866961} /* (29, 6, 17) {real, imag} */,
  {32'hc0ef9ea8, 32'h4156ffd0} /* (29, 6, 16) {real, imag} */,
  {32'h3fd42400, 32'h418d86db} /* (29, 6, 15) {real, imag} */,
  {32'hc1d9731d, 32'h41da4a30} /* (29, 6, 14) {real, imag} */,
  {32'hc20969b1, 32'h40b7be58} /* (29, 6, 13) {real, imag} */,
  {32'h40e172f4, 32'hc08188e6} /* (29, 6, 12) {real, imag} */,
  {32'hc230158c, 32'hc2b29ab7} /* (29, 6, 11) {real, imag} */,
  {32'h412f3f10, 32'h403f29f0} /* (29, 6, 10) {real, imag} */,
  {32'hc2e350d3, 32'h42ad6267} /* (29, 6, 9) {real, imag} */,
  {32'h42d37c60, 32'hc210501c} /* (29, 6, 8) {real, imag} */,
  {32'hc2c62343, 32'hc2d63e79} /* (29, 6, 7) {real, imag} */,
  {32'h4265c9d8, 32'hc31af928} /* (29, 6, 6) {real, imag} */,
  {32'h4251464b, 32'hc1b57e25} /* (29, 6, 5) {real, imag} */,
  {32'h42bc13b7, 32'hc227448a} /* (29, 6, 4) {real, imag} */,
  {32'h4215a302, 32'hc0edc3b8} /* (29, 6, 3) {real, imag} */,
  {32'hc25f40d4, 32'h425d5d05} /* (29, 6, 2) {real, imag} */,
  {32'hc09be3f0, 32'h42bf61cc} /* (29, 6, 1) {real, imag} */,
  {32'h427a2d6d, 32'h42cda874} /* (29, 6, 0) {real, imag} */,
  {32'hc1d5ee20, 32'h4390bc77} /* (29, 5, 31) {real, imag} */,
  {32'hc33421ab, 32'hc3124807} /* (29, 5, 30) {real, imag} */,
  {32'hc1933b19, 32'hc1f1b0dc} /* (29, 5, 29) {real, imag} */,
  {32'h42964e42, 32'h42d16195} /* (29, 5, 28) {real, imag} */,
  {32'hc30234f3, 32'hc324c7c0} /* (29, 5, 27) {real, imag} */,
  {32'h42108d38, 32'h42087de9} /* (29, 5, 26) {real, imag} */,
  {32'h42c6438e, 32'h41c362ae} /* (29, 5, 25) {real, imag} */,
  {32'h4282201a, 32'hc2b57d50} /* (29, 5, 24) {real, imag} */,
  {32'h41f7c75f, 32'h41a86f83} /* (29, 5, 23) {real, imag} */,
  {32'hc2499cf6, 32'hc13c8a24} /* (29, 5, 22) {real, imag} */,
  {32'hc11ffb60, 32'hc210ff11} /* (29, 5, 21) {real, imag} */,
  {32'hc1af5c54, 32'h4136ecd6} /* (29, 5, 20) {real, imag} */,
  {32'h41a80868, 32'h41c3eabd} /* (29, 5, 19) {real, imag} */,
  {32'hc1b5c9c6, 32'h41fccbf2} /* (29, 5, 18) {real, imag} */,
  {32'h41a0bed6, 32'hc1a7a2a6} /* (29, 5, 17) {real, imag} */,
  {32'hc175cf30, 32'h40e8dee0} /* (29, 5, 16) {real, imag} */,
  {32'h40e11f18, 32'hc217c565} /* (29, 5, 15) {real, imag} */,
  {32'h4194f382, 32'h40c26768} /* (29, 5, 14) {real, imag} */,
  {32'h4250f690, 32'hc1196b7a} /* (29, 5, 13) {real, imag} */,
  {32'hc1b20d1c, 32'h41be2121} /* (29, 5, 12) {real, imag} */,
  {32'hc20c0560, 32'hc1762245} /* (29, 5, 11) {real, imag} */,
  {32'hc184c455, 32'h42758861} /* (29, 5, 10) {real, imag} */,
  {32'h410f9626, 32'h425c5db4} /* (29, 5, 9) {real, imag} */,
  {32'hc1802457, 32'h4135ed80} /* (29, 5, 8) {real, imag} */,
  {32'h42771937, 32'hc2e4046c} /* (29, 5, 7) {real, imag} */,
  {32'hc2567fa4, 32'hc1e2442a} /* (29, 5, 6) {real, imag} */,
  {32'h4365269f, 32'hc2cfc9a4} /* (29, 5, 5) {real, imag} */,
  {32'hc29efca4, 32'h42c6cf33} /* (29, 5, 4) {real, imag} */,
  {32'hc1190572, 32'h4259c45e} /* (29, 5, 3) {real, imag} */,
  {32'h426d1aa1, 32'hc2de933e} /* (29, 5, 2) {real, imag} */,
  {32'hc34570e8, 32'h432fae1f} /* (29, 5, 1) {real, imag} */,
  {32'h42c5d6b2, 32'h43b26d66} /* (29, 5, 0) {real, imag} */,
  {32'h435352d9, 32'hc2ed73e2} /* (29, 4, 31) {real, imag} */,
  {32'hc37a30ec, 32'h43acdede} /* (29, 4, 30) {real, imag} */,
  {32'h40a10dc4, 32'h3f119940} /* (29, 4, 29) {real, imag} */,
  {32'h423c5c40, 32'hc244a3d0} /* (29, 4, 28) {real, imag} */,
  {32'hc28ad0b4, 32'hc1bdbd94} /* (29, 4, 27) {real, imag} */,
  {32'h43062036, 32'hc13f47ec} /* (29, 4, 26) {real, imag} */,
  {32'h42b069d2, 32'hc2591b66} /* (29, 4, 25) {real, imag} */,
  {32'hc118fdc0, 32'h428242da} /* (29, 4, 24) {real, imag} */,
  {32'h428ec202, 32'hc294b460} /* (29, 4, 23) {real, imag} */,
  {32'hc273b3eb, 32'hc29fc476} /* (29, 4, 22) {real, imag} */,
  {32'hc24cfbdb, 32'h4265a594} /* (29, 4, 21) {real, imag} */,
  {32'hc14fa033, 32'hc1df1f25} /* (29, 4, 20) {real, imag} */,
  {32'h41c760df, 32'hc19bacd7} /* (29, 4, 19) {real, imag} */,
  {32'hc1a77410, 32'h428350d4} /* (29, 4, 18) {real, imag} */,
  {32'hc154865a, 32'h4138f4e0} /* (29, 4, 17) {real, imag} */,
  {32'h3e516000, 32'h41c1b8c2} /* (29, 4, 16) {real, imag} */,
  {32'h420246c6, 32'hc1211c80} /* (29, 4, 15) {real, imag} */,
  {32'h42200990, 32'h4118001c} /* (29, 4, 14) {real, imag} */,
  {32'hc1562f1e, 32'hc2619bbe} /* (29, 4, 13) {real, imag} */,
  {32'hc151b681, 32'h40980f0c} /* (29, 4, 12) {real, imag} */,
  {32'hc275defd, 32'hc1bc7584} /* (29, 4, 11) {real, imag} */,
  {32'hc18d24ee, 32'h42dd50ba} /* (29, 4, 10) {real, imag} */,
  {32'hc210a5ec, 32'h4219c7fc} /* (29, 4, 9) {real, imag} */,
  {32'hc243e51b, 32'hc27804ad} /* (29, 4, 8) {real, imag} */,
  {32'hc1124630, 32'hc33c76e4} /* (29, 4, 7) {real, imag} */,
  {32'h4290c6d7, 32'hc2e99742} /* (29, 4, 6) {real, imag} */,
  {32'h42c67148, 32'hc24d7946} /* (29, 4, 5) {real, imag} */,
  {32'h42b2074c, 32'hc05a21f8} /* (29, 4, 4) {real, imag} */,
  {32'hc2237bb6, 32'h42e855ba} /* (29, 4, 3) {real, imag} */,
  {32'hc3120686, 32'h43af3ed8} /* (29, 4, 2) {real, imag} */,
  {32'h435e155f, 32'hc4036c94} /* (29, 4, 1) {real, imag} */,
  {32'h4332c5c4, 32'hc2b27564} /* (29, 4, 0) {real, imag} */,
  {32'h433b0260, 32'h43b692bb} /* (29, 3, 31) {real, imag} */,
  {32'hc39deaa4, 32'hc2efafe8} /* (29, 3, 30) {real, imag} */,
  {32'h416457d8, 32'hc1808490} /* (29, 3, 29) {real, imag} */,
  {32'h41af8a44, 32'hc2ca7ff7} /* (29, 3, 28) {real, imag} */,
  {32'hc33963ab, 32'h434f28cb} /* (29, 3, 27) {real, imag} */,
  {32'h421e944e, 32'hc1a0a336} /* (29, 3, 26) {real, imag} */,
  {32'h431f8208, 32'h41328a3c} /* (29, 3, 25) {real, imag} */,
  {32'hc264ae9a, 32'h42d04b00} /* (29, 3, 24) {real, imag} */,
  {32'h4291523a, 32'hc2d9491c} /* (29, 3, 23) {real, imag} */,
  {32'hc30f0812, 32'hc206334f} /* (29, 3, 22) {real, imag} */,
  {32'h4291561a, 32'h423518c0} /* (29, 3, 21) {real, imag} */,
  {32'hc1e5aac6, 32'hc1ab65c4} /* (29, 3, 20) {real, imag} */,
  {32'h42018940, 32'h3f704320} /* (29, 3, 19) {real, imag} */,
  {32'h415caf12, 32'hc08f064c} /* (29, 3, 18) {real, imag} */,
  {32'hc23bd913, 32'hc1a5a6f8} /* (29, 3, 17) {real, imag} */,
  {32'h41e3fcbc, 32'h41d0fbf4} /* (29, 3, 16) {real, imag} */,
  {32'h419e39e6, 32'hc18c56b8} /* (29, 3, 15) {real, imag} */,
  {32'hc23426b4, 32'hc1d4392d} /* (29, 3, 14) {real, imag} */,
  {32'hc21b9c84, 32'h41ac4697} /* (29, 3, 13) {real, imag} */,
  {32'h424acd2b, 32'h42b0fbe4} /* (29, 3, 12) {real, imag} */,
  {32'hc09bea18, 32'h4237e99a} /* (29, 3, 11) {real, imag} */,
  {32'h423a4e4a, 32'h42b3f0ac} /* (29, 3, 10) {real, imag} */,
  {32'h41efd600, 32'hc282d1f0} /* (29, 3, 9) {real, imag} */,
  {32'hc28d34ab, 32'h42fabd4c} /* (29, 3, 8) {real, imag} */,
  {32'h430edcd8, 32'h3f14bc40} /* (29, 3, 7) {real, imag} */,
  {32'hc0130960, 32'h42908352} /* (29, 3, 6) {real, imag} */,
  {32'hc3102551, 32'hc1ccfea8} /* (29, 3, 5) {real, imag} */,
  {32'h431c5d4a, 32'h41a923d0} /* (29, 3, 4) {real, imag} */,
  {32'h42543ba2, 32'hc2d3e996} /* (29, 3, 3) {real, imag} */,
  {32'hc3e09e62, 32'hc121c110} /* (29, 3, 2) {real, imag} */,
  {32'h4113e8a8, 32'hc39e6f1d} /* (29, 3, 1) {real, imag} */,
  {32'hc235478a, 32'h42926d07} /* (29, 3, 0) {real, imag} */,
  {32'h4346b570, 32'h44994ca2} /* (29, 2, 31) {real, imag} */,
  {32'hc40083f8, 32'hc4090cbf} /* (29, 2, 30) {real, imag} */,
  {32'h42ce2aab, 32'hc14ad61c} /* (29, 2, 29) {real, imag} */,
  {32'h433c83a0, 32'h419fef78} /* (29, 2, 28) {real, imag} */,
  {32'hc2c12646, 32'hc328baad} /* (29, 2, 27) {real, imag} */,
  {32'h4248bff0, 32'hc31a2b39} /* (29, 2, 26) {real, imag} */,
  {32'hc1f2596c, 32'hc2e34d2f} /* (29, 2, 25) {real, imag} */,
  {32'hc2bb9e2c, 32'hc33cf2d6} /* (29, 2, 24) {real, imag} */,
  {32'hc22e67a2, 32'hc2099ebb} /* (29, 2, 23) {real, imag} */,
  {32'hc1866ff0, 32'h417cff40} /* (29, 2, 22) {real, imag} */,
  {32'hc20305b8, 32'h41637f0c} /* (29, 2, 21) {real, imag} */,
  {32'hc19cf575, 32'h4194ad04} /* (29, 2, 20) {real, imag} */,
  {32'hc1ea09f3, 32'hc147619e} /* (29, 2, 19) {real, imag} */,
  {32'hc28c216e, 32'hc19fc5e8} /* (29, 2, 18) {real, imag} */,
  {32'hc1955c67, 32'hc24c5c7a} /* (29, 2, 17) {real, imag} */,
  {32'h4002aa00, 32'h3d0c0000} /* (29, 2, 16) {real, imag} */,
  {32'h4019f838, 32'h40e441d0} /* (29, 2, 15) {real, imag} */,
  {32'h41c5d356, 32'h424aac54} /* (29, 2, 14) {real, imag} */,
  {32'hc1a62403, 32'h4168924a} /* (29, 2, 13) {real, imag} */,
  {32'h4121cdda, 32'h420125aa} /* (29, 2, 12) {real, imag} */,
  {32'h42758d28, 32'hc2cf9f8c} /* (29, 2, 11) {real, imag} */,
  {32'hc1b1f798, 32'h429febae} /* (29, 2, 10) {real, imag} */,
  {32'h42bcfbff, 32'hc2fd7860} /* (29, 2, 9) {real, imag} */,
  {32'hc32c5786, 32'hc30d74c8} /* (29, 2, 8) {real, imag} */,
  {32'hc3173322, 32'h42d54875} /* (29, 2, 7) {real, imag} */,
  {32'hc211aa9c, 32'hc2a510d0} /* (29, 2, 6) {real, imag} */,
  {32'hc3266219, 32'hc34c42a7} /* (29, 2, 5) {real, imag} */,
  {32'h4224eae2, 32'h43ebc390} /* (29, 2, 4) {real, imag} */,
  {32'h426abfa6, 32'hc283af30} /* (29, 2, 3) {real, imag} */,
  {32'hc3b92a70, 32'hc41b7155} /* (29, 2, 2) {real, imag} */,
  {32'h4386b62e, 32'h4438dfd0} /* (29, 2, 1) {real, imag} */,
  {32'hc24383b0, 32'h444000c4} /* (29, 2, 0) {real, imag} */,
  {32'hc413db37, 32'hc42fc8ba} /* (29, 1, 31) {real, imag} */,
  {32'h42c41024, 32'h43d490cc} /* (29, 1, 30) {real, imag} */,
  {32'hc2f741e3, 32'h427883e4} /* (29, 1, 29) {real, imag} */,
  {32'h426cf194, 32'hc3484a69} /* (29, 1, 28) {real, imag} */,
  {32'h4362772c, 32'h4389fb8a} /* (29, 1, 27) {real, imag} */,
  {32'hc08bdd50, 32'h42a0a354} /* (29, 1, 26) {real, imag} */,
  {32'hc1f0d0fa, 32'hc345a00c} /* (29, 1, 25) {real, imag} */,
  {32'h4299005c, 32'h42dbc563} /* (29, 1, 24) {real, imag} */,
  {32'h40a00cb8, 32'hc2ef47f0} /* (29, 1, 23) {real, imag} */,
  {32'h4287fa64, 32'h420096ba} /* (29, 1, 22) {real, imag} */,
  {32'h4300eb3a, 32'h4336d1ee} /* (29, 1, 21) {real, imag} */,
  {32'hc143ca46, 32'hc19624f3} /* (29, 1, 20) {real, imag} */,
  {32'hc157b482, 32'hc21169f7} /* (29, 1, 19) {real, imag} */,
  {32'h42b71b25, 32'h42475e64} /* (29, 1, 18) {real, imag} */,
  {32'h41700bfc, 32'hc1625b80} /* (29, 1, 17) {real, imag} */,
  {32'h41715e44, 32'h423f3618} /* (29, 1, 16) {real, imag} */,
  {32'h42452447, 32'h40882d00} /* (29, 1, 15) {real, imag} */,
  {32'hc2c587d5, 32'h41bb3c98} /* (29, 1, 14) {real, imag} */,
  {32'h417e001e, 32'h415c94bc} /* (29, 1, 13) {real, imag} */,
  {32'h41eedfc1, 32'h41efbf23} /* (29, 1, 12) {real, imag} */,
  {32'hc1e0473c, 32'h421af7f2} /* (29, 1, 11) {real, imag} */,
  {32'h414395b0, 32'hbfc13540} /* (29, 1, 10) {real, imag} */,
  {32'h428ca284, 32'h41847ca0} /* (29, 1, 9) {real, imag} */,
  {32'hc3102c5c, 32'hc01ab560} /* (29, 1, 8) {real, imag} */,
  {32'h42454553, 32'hc2b71530} /* (29, 1, 7) {real, imag} */,
  {32'h42955a09, 32'h42c55144} /* (29, 1, 6) {real, imag} */,
  {32'hc33a1b36, 32'h43b8baaa} /* (29, 1, 5) {real, imag} */,
  {32'hc29b7a82, 32'hc37ebbff} /* (29, 1, 4) {real, imag} */,
  {32'h437d3044, 32'h4379e8f7} /* (29, 1, 3) {real, imag} */,
  {32'hc3c5f1ad, 32'h4444bcfa} /* (29, 1, 2) {real, imag} */,
  {32'h438b212e, 32'hc4ca2031} /* (29, 1, 1) {real, imag} */,
  {32'hc307e6ed, 32'hc47244dc} /* (29, 1, 0) {real, imag} */,
  {32'hc40eb485, 32'hc409e052} /* (29, 0, 31) {real, imag} */,
  {32'h434e934c, 32'h42071224} /* (29, 0, 30) {real, imag} */,
  {32'hc311781a, 32'h43792164} /* (29, 0, 29) {real, imag} */,
  {32'h43372f4a, 32'h41fc1c81} /* (29, 0, 28) {real, imag} */,
  {32'h4395434c, 32'h4364d05f} /* (29, 0, 27) {real, imag} */,
  {32'hc3547680, 32'hc2681938} /* (29, 0, 26) {real, imag} */,
  {32'hc31ec62a, 32'h4332fd1a} /* (29, 0, 25) {real, imag} */,
  {32'h42e56964, 32'h41e0a3d8} /* (29, 0, 24) {real, imag} */,
  {32'h41d12fd5, 32'h422c796e} /* (29, 0, 23) {real, imag} */,
  {32'h4301800e, 32'hc29d42b4} /* (29, 0, 22) {real, imag} */,
  {32'h4277e490, 32'hc1ee88e6} /* (29, 0, 21) {real, imag} */,
  {32'hc2d18f99, 32'hc08b0f18} /* (29, 0, 20) {real, imag} */,
  {32'hc181a72a, 32'hc29dc86d} /* (29, 0, 19) {real, imag} */,
  {32'h422c18a3, 32'hc2a6ac24} /* (29, 0, 18) {real, imag} */,
  {32'hc2280867, 32'hc1629ea6} /* (29, 0, 17) {real, imag} */,
  {32'hc13646c8, 32'h421b86b4} /* (29, 0, 16) {real, imag} */,
  {32'hc1690f1c, 32'h4201531a} /* (29, 0, 15) {real, imag} */,
  {32'h40f00918, 32'h423c0ce8} /* (29, 0, 14) {real, imag} */,
  {32'hc0cb6f38, 32'h4195d12c} /* (29, 0, 13) {real, imag} */,
  {32'h424214b6, 32'hc2725419} /* (29, 0, 12) {real, imag} */,
  {32'hc1155080, 32'h428487f6} /* (29, 0, 11) {real, imag} */,
  {32'h42162baa, 32'hc2846b08} /* (29, 0, 10) {real, imag} */,
  {32'h41c4c22d, 32'hc2b3fec3} /* (29, 0, 9) {real, imag} */,
  {32'hc2e257d6, 32'hc28073c2} /* (29, 0, 8) {real, imag} */,
  {32'h42da2024, 32'hc28ea669} /* (29, 0, 7) {real, imag} */,
  {32'hc2cfc59c, 32'h4277bc00} /* (29, 0, 6) {real, imag} */,
  {32'h42bb0b1e, 32'h438131fd} /* (29, 0, 5) {real, imag} */,
  {32'hc37d26c0, 32'h41919b99} /* (29, 0, 4) {real, imag} */,
  {32'hc33eb7a6, 32'h41e8afc0} /* (29, 0, 3) {real, imag} */,
  {32'hc364a3a4, 32'h43612c2f} /* (29, 0, 2) {real, imag} */,
  {32'h43ea177a, 32'hc42cf7a2} /* (29, 0, 1) {real, imag} */,
  {32'hc35da878, 32'hc3e39f5c} /* (29, 0, 0) {real, imag} */,
  {32'hc48513ed, 32'hc451fb6d} /* (28, 31, 31) {real, imag} */,
  {32'h445fd3a6, 32'h4368218a} /* (28, 31, 30) {real, imag} */,
  {32'hc213a924, 32'h432c0029} /* (28, 31, 29) {real, imag} */,
  {32'hc221809b, 32'h416d77c8} /* (28, 31, 28) {real, imag} */,
  {32'h4380b248, 32'h43208d62} /* (28, 31, 27) {real, imag} */,
  {32'h42f6f576, 32'hc29b6962} /* (28, 31, 26) {real, imag} */,
  {32'hc1c76b14, 32'h40e401d4} /* (28, 31, 25) {real, imag} */,
  {32'h433c3915, 32'h410f8560} /* (28, 31, 24) {real, imag} */,
  {32'h428076e7, 32'hc2a40421} /* (28, 31, 23) {real, imag} */,
  {32'hc23af6c4, 32'h4268f83d} /* (28, 31, 22) {real, imag} */,
  {32'h42897bf3, 32'h41a34d00} /* (28, 31, 21) {real, imag} */,
  {32'hbf9bd7e0, 32'h427854dc} /* (28, 31, 20) {real, imag} */,
  {32'hc1981388, 32'h4154f7dc} /* (28, 31, 19) {real, imag} */,
  {32'h40ac85e0, 32'hc208e3d6} /* (28, 31, 18) {real, imag} */,
  {32'hc22ec200, 32'h421d2702} /* (28, 31, 17) {real, imag} */,
  {32'h424af840, 32'hc1b6bf80} /* (28, 31, 16) {real, imag} */,
  {32'hc18d8c20, 32'h410868f8} /* (28, 31, 15) {real, imag} */,
  {32'hc2a6409a, 32'hc0c98150} /* (28, 31, 14) {real, imag} */,
  {32'hc21824d6, 32'hc173f114} /* (28, 31, 13) {real, imag} */,
  {32'h42e1514a, 32'hc203cac8} /* (28, 31, 12) {real, imag} */,
  {32'hc364b8de, 32'h43129b63} /* (28, 31, 11) {real, imag} */,
  {32'h41686ba0, 32'hc236185d} /* (28, 31, 10) {real, imag} */,
  {32'h4105c998, 32'hc1541c58} /* (28, 31, 9) {real, imag} */,
  {32'hc2b01946, 32'h433bfc2a} /* (28, 31, 8) {real, imag} */,
  {32'h4300b8bc, 32'hc1b01ae5} /* (28, 31, 7) {real, imag} */,
  {32'hc2dbaf48, 32'hc2a3e556} /* (28, 31, 6) {real, imag} */,
  {32'h4331077c, 32'h43e08325} /* (28, 31, 5) {real, imag} */,
  {32'hc260ad09, 32'hc37f9fd8} /* (28, 31, 4) {real, imag} */,
  {32'hc171be28, 32'hc302885f} /* (28, 31, 3) {real, imag} */,
  {32'h432f9d72, 32'h43cf50f3} /* (28, 31, 2) {real, imag} */,
  {32'hc21772e0, 32'hc458d853} /* (28, 31, 1) {real, imag} */,
  {32'hc4187fe4, 32'hc4335fe0} /* (28, 31, 0) {real, imag} */,
  {32'h42ded3d6, 32'h44219004} /* (28, 30, 31) {real, imag} */,
  {32'hc0d94ba0, 32'hc40b0116} /* (28, 30, 30) {real, imag} */,
  {32'h426704e9, 32'h42ee9807} /* (28, 30, 29) {real, imag} */,
  {32'hc2202d16, 32'h4347adf6} /* (28, 30, 28) {real, imag} */,
  {32'hc333c5dc, 32'hc3402cb6} /* (28, 30, 27) {real, imag} */,
  {32'hc28f3f24, 32'h41e6b50e} /* (28, 30, 26) {real, imag} */,
  {32'h42b66e31, 32'h4183c5d2} /* (28, 30, 25) {real, imag} */,
  {32'hc2b9f1ce, 32'hc32b0f20} /* (28, 30, 24) {real, imag} */,
  {32'hc2a4985f, 32'hc1c35f9a} /* (28, 30, 23) {real, imag} */,
  {32'h3f6bdf80, 32'h42666b70} /* (28, 30, 22) {real, imag} */,
  {32'hc28c1c13, 32'hc0abad80} /* (28, 30, 21) {real, imag} */,
  {32'h40b3865c, 32'h424f6d0b} /* (28, 30, 20) {real, imag} */,
  {32'h41181756, 32'h41b076fe} /* (28, 30, 19) {real, imag} */,
  {32'hc22e2507, 32'hc28269a2} /* (28, 30, 18) {real, imag} */,
  {32'hc1bcb0d8, 32'h41c08c0c} /* (28, 30, 17) {real, imag} */,
  {32'hc223f8d4, 32'hc1e3caa0} /* (28, 30, 16) {real, imag} */,
  {32'hc0f61ca0, 32'h3c22a000} /* (28, 30, 15) {real, imag} */,
  {32'h4170319c, 32'h40c3af98} /* (28, 30, 14) {real, imag} */,
  {32'h408f6f9c, 32'hc0eded76} /* (28, 30, 13) {real, imag} */,
  {32'hc2125cf0, 32'h41d237ea} /* (28, 30, 12) {real, imag} */,
  {32'h42b59bdb, 32'hc28f6174} /* (28, 30, 11) {real, imag} */,
  {32'hc2eb4c5e, 32'hc19deb00} /* (28, 30, 10) {real, imag} */,
  {32'h426dfbaa, 32'hc1e0ed6a} /* (28, 30, 9) {real, imag} */,
  {32'h423ef19b, 32'hc35ab78a} /* (28, 30, 8) {real, imag} */,
  {32'h41a5f234, 32'h426c1119} /* (28, 30, 7) {real, imag} */,
  {32'hc28ab4f8, 32'h42918d04} /* (28, 30, 6) {real, imag} */,
  {32'h42986463, 32'hc34622dc} /* (28, 30, 5) {real, imag} */,
  {32'hc2b91d45, 32'h438a876f} /* (28, 30, 4) {real, imag} */,
  {32'h42821580, 32'h432da934} /* (28, 30, 3) {real, imag} */,
  {32'hc33ec105, 32'hc4495bc2} /* (28, 30, 2) {real, imag} */,
  {32'h43f08c8a, 32'h448965da} /* (28, 30, 1) {real, imag} */,
  {32'h439cd4c0, 32'h440c71b3} /* (28, 30, 0) {real, imag} */,
  {32'hc384a7bc, 32'h41c1d010} /* (28, 29, 31) {real, imag} */,
  {32'h43260ce4, 32'h41b18c98} /* (28, 29, 30) {real, imag} */,
  {32'hc30ff4fc, 32'hc090f940} /* (28, 29, 29) {real, imag} */,
  {32'h426def32, 32'h413ddf32} /* (28, 29, 28) {real, imag} */,
  {32'h422d7c0f, 32'hc2ba5224} /* (28, 29, 27) {real, imag} */,
  {32'h41f1c324, 32'hc3117148} /* (28, 29, 26) {real, imag} */,
  {32'hc318712c, 32'hc3105535} /* (28, 29, 25) {real, imag} */,
  {32'h40e33f68, 32'h40fd9b1c} /* (28, 29, 24) {real, imag} */,
  {32'h424013b4, 32'h42621aec} /* (28, 29, 23) {real, imag} */,
  {32'hc1c21d7e, 32'h42a6689b} /* (28, 29, 22) {real, imag} */,
  {32'h40478b68, 32'hc228211f} /* (28, 29, 21) {real, imag} */,
  {32'h400e5930, 32'h426928f6} /* (28, 29, 20) {real, imag} */,
  {32'hc263e17a, 32'hc166ba3a} /* (28, 29, 19) {real, imag} */,
  {32'hc149de1e, 32'hc2043e8c} /* (28, 29, 18) {real, imag} */,
  {32'hc113e884, 32'hc0f01be0} /* (28, 29, 17) {real, imag} */,
  {32'hc0dc4390, 32'hc249baad} /* (28, 29, 16) {real, imag} */,
  {32'hc21474e9, 32'h42798708} /* (28, 29, 15) {real, imag} */,
  {32'h41fa612f, 32'hc2073940} /* (28, 29, 14) {real, imag} */,
  {32'h4234c688, 32'hc1a5a17b} /* (28, 29, 13) {real, imag} */,
  {32'hc2ad3ee4, 32'hc243f376} /* (28, 29, 12) {real, imag} */,
  {32'h42122ca4, 32'h42affebe} /* (28, 29, 11) {real, imag} */,
  {32'hc1dd359e, 32'hc2631d4e} /* (28, 29, 10) {real, imag} */,
  {32'hc2ef3c6c, 32'hc0e227d0} /* (28, 29, 9) {real, imag} */,
  {32'h41ac8d74, 32'hc22ec4f6} /* (28, 29, 8) {real, imag} */,
  {32'h42564e04, 32'h42657b43} /* (28, 29, 7) {real, imag} */,
  {32'h3fb42200, 32'h421a6814} /* (28, 29, 6) {real, imag} */,
  {32'h4287aa9a, 32'hc2da851c} /* (28, 29, 5) {real, imag} */,
  {32'hc280f7d0, 32'h4295e026} /* (28, 29, 4) {real, imag} */,
  {32'h42167406, 32'hc2cf41fe} /* (28, 29, 3) {real, imag} */,
  {32'h437fe440, 32'hc33d60c8} /* (28, 29, 2) {real, imag} */,
  {32'h41ec92b0, 32'h43a0893f} /* (28, 29, 1) {real, imag} */,
  {32'h41ef2aaa, 32'h4193afc6} /* (28, 29, 0) {real, imag} */,
  {32'hc39f7cc5, 32'hc3f6cfa4} /* (28, 28, 31) {real, imag} */,
  {32'h439e3b3e, 32'h42ac0b71} /* (28, 28, 30) {real, imag} */,
  {32'hc26352aa, 32'hc2d0f913} /* (28, 28, 29) {real, imag} */,
  {32'hc2d345e9, 32'h41ec51c4} /* (28, 28, 28) {real, imag} */,
  {32'h4044aea8, 32'h4196d934} /* (28, 28, 27) {real, imag} */,
  {32'h42a9e92c, 32'h42c4f558} /* (28, 28, 26) {real, imag} */,
  {32'hc2a9a5e2, 32'hc1e9115c} /* (28, 28, 25) {real, imag} */,
  {32'h427a8e60, 32'h404e67f0} /* (28, 28, 24) {real, imag} */,
  {32'h42a8b910, 32'hc29d0343} /* (28, 28, 23) {real, imag} */,
  {32'h419d79c4, 32'h4223ae70} /* (28, 28, 22) {real, imag} */,
  {32'h42359af6, 32'hc17a0752} /* (28, 28, 21) {real, imag} */,
  {32'hc147e068, 32'h412f92e4} /* (28, 28, 20) {real, imag} */,
  {32'h429c8fd1, 32'hc1a127b6} /* (28, 28, 19) {real, imag} */,
  {32'h41854db4, 32'h41a27f84} /* (28, 28, 18) {real, imag} */,
  {32'h41489a6e, 32'h3f384580} /* (28, 28, 17) {real, imag} */,
  {32'h41279da8, 32'h4139a79c} /* (28, 28, 16) {real, imag} */,
  {32'hc1c74447, 32'h40e89c90} /* (28, 28, 15) {real, imag} */,
  {32'hc12498e8, 32'hc16fbd1c} /* (28, 28, 14) {real, imag} */,
  {32'hc2048fbe, 32'hc276738b} /* (28, 28, 13) {real, imag} */,
  {32'h3d0ea800, 32'hc1978172} /* (28, 28, 12) {real, imag} */,
  {32'h421955d6, 32'h4243cc94} /* (28, 28, 11) {real, imag} */,
  {32'hc1e8ff88, 32'hc1e2df88} /* (28, 28, 10) {real, imag} */,
  {32'h42bd93b8, 32'h4236749e} /* (28, 28, 9) {real, imag} */,
  {32'hc1c737c0, 32'h41eda3b6} /* (28, 28, 8) {real, imag} */,
  {32'hc2d7fd16, 32'h408284b8} /* (28, 28, 7) {real, imag} */,
  {32'h428959f0, 32'hc294aaaa} /* (28, 28, 6) {real, imag} */,
  {32'hc0d48644, 32'h43020d26} /* (28, 28, 5) {real, imag} */,
  {32'hc3971dfc, 32'hc32bed84} /* (28, 28, 4) {real, imag} */,
  {32'hc29059ab, 32'h42e1e375} /* (28, 28, 3) {real, imag} */,
  {32'h4385594a, 32'hc2703c55} /* (28, 28, 2) {real, imag} */,
  {32'hc399286f, 32'hc3598428} /* (28, 28, 1) {real, imag} */,
  {32'hc306c1a6, 32'hc28ad316} /* (28, 28, 0) {real, imag} */,
  {32'h438ab83c, 32'h42fc39d6} /* (28, 27, 31) {real, imag} */,
  {32'hc2db163e, 32'hc2cf12ff} /* (28, 27, 30) {real, imag} */,
  {32'hc2bc84de, 32'hc1a7aad2} /* (28, 27, 29) {real, imag} */,
  {32'hc29623ad, 32'hc20d019c} /* (28, 27, 28) {real, imag} */,
  {32'h3f33a880, 32'hc19b8ee6} /* (28, 27, 27) {real, imag} */,
  {32'hc227c962, 32'hc34f2845} /* (28, 27, 26) {real, imag} */,
  {32'h4218aeea, 32'h41049670} /* (28, 27, 25) {real, imag} */,
  {32'h4189fe78, 32'h429ccfb2} /* (28, 27, 24) {real, imag} */,
  {32'hc28f2edc, 32'h40ecf378} /* (28, 27, 23) {real, imag} */,
  {32'h412e98e9, 32'h42d17d84} /* (28, 27, 22) {real, imag} */,
  {32'hc20deb09, 32'hc13c62d2} /* (28, 27, 21) {real, imag} */,
  {32'h40c8a97c, 32'hc09d3a18} /* (28, 27, 20) {real, imag} */,
  {32'h4215e6c7, 32'h40b1aa4a} /* (28, 27, 19) {real, imag} */,
  {32'h41290abc, 32'h40d3fcec} /* (28, 27, 18) {real, imag} */,
  {32'h4109b428, 32'h408ed78c} /* (28, 27, 17) {real, imag} */,
  {32'h419ed534, 32'h410bb9b8} /* (28, 27, 16) {real, imag} */,
  {32'hc1561608, 32'hbeb9acc0} /* (28, 27, 15) {real, imag} */,
  {32'h418da94a, 32'hc1cba59b} /* (28, 27, 14) {real, imag} */,
  {32'h42a84158, 32'h41854ff6} /* (28, 27, 13) {real, imag} */,
  {32'h400446b8, 32'h424f8c76} /* (28, 27, 12) {real, imag} */,
  {32'hc1cdb396, 32'hc24dd29e} /* (28, 27, 11) {real, imag} */,
  {32'hc167a3e7, 32'h417a58b0} /* (28, 27, 10) {real, imag} */,
  {32'h422b8d42, 32'h41d0d9ae} /* (28, 27, 9) {real, imag} */,
  {32'hc1cf3ff0, 32'h4247541b} /* (28, 27, 8) {real, imag} */,
  {32'hc2d18537, 32'h42f23c86} /* (28, 27, 7) {real, imag} */,
  {32'hc15eb798, 32'h406fb080} /* (28, 27, 6) {real, imag} */,
  {32'hc25b46a0, 32'hc3001300} /* (28, 27, 5) {real, imag} */,
  {32'h4319bfa6, 32'h4280b2c4} /* (28, 27, 4) {real, imag} */,
  {32'h426f58ec, 32'h4186933a} /* (28, 27, 3) {real, imag} */,
  {32'hc133e8fc, 32'hc27b6a22} /* (28, 27, 2) {real, imag} */,
  {32'h425783fc, 32'h4336db67} /* (28, 27, 1) {real, imag} */,
  {32'h431c8412, 32'h4308ac3a} /* (28, 27, 0) {real, imag} */,
  {32'hc1d52714, 32'h42944c32} /* (28, 26, 31) {real, imag} */,
  {32'hc2adf448, 32'h42f36825} /* (28, 26, 30) {real, imag} */,
  {32'h411bd762, 32'hc22cf3f3} /* (28, 26, 29) {real, imag} */,
  {32'h423e2fba, 32'h415b5630} /* (28, 26, 28) {real, imag} */,
  {32'h42477ec8, 32'hc21f8df9} /* (28, 26, 27) {real, imag} */,
  {32'hc0adf3e0, 32'h42d7f3ed} /* (28, 26, 26) {real, imag} */,
  {32'hbfd1d7d0, 32'h4231bc1a} /* (28, 26, 25) {real, imag} */,
  {32'h41fbd9c4, 32'hc2470b49} /* (28, 26, 24) {real, imag} */,
  {32'h42781e54, 32'h42129546} /* (28, 26, 23) {real, imag} */,
  {32'hc1618134, 32'hc23f84bf} /* (28, 26, 22) {real, imag} */,
  {32'hc24a516c, 32'h41925cee} /* (28, 26, 21) {real, imag} */,
  {32'hc1ec4be3, 32'hc21be1aa} /* (28, 26, 20) {real, imag} */,
  {32'hc137a7be, 32'h41fa011e} /* (28, 26, 19) {real, imag} */,
  {32'hc1b657f6, 32'hc1890cb6} /* (28, 26, 18) {real, imag} */,
  {32'h3e9f1700, 32'hc18e8912} /* (28, 26, 17) {real, imag} */,
  {32'h411f34d2, 32'hbef64100} /* (28, 26, 16) {real, imag} */,
  {32'h41b2d392, 32'hc0e59752} /* (28, 26, 15) {real, imag} */,
  {32'h413d102c, 32'hc0806566} /* (28, 26, 14) {real, imag} */,
  {32'h4197c325, 32'h41ecbc2e} /* (28, 26, 13) {real, imag} */,
  {32'h40381078, 32'h42b81b75} /* (28, 26, 12) {real, imag} */,
  {32'h424be4e2, 32'h420c0734} /* (28, 26, 11) {real, imag} */,
  {32'hc1fdeb46, 32'h42cba27a} /* (28, 26, 10) {real, imag} */,
  {32'h428f11fe, 32'h417275e6} /* (28, 26, 9) {real, imag} */,
  {32'h42c1b707, 32'h41f8391a} /* (28, 26, 8) {real, imag} */,
  {32'hc0fa15a4, 32'hc294c585} /* (28, 26, 7) {real, imag} */,
  {32'hc2577456, 32'hc229c3a2} /* (28, 26, 6) {real, imag} */,
  {32'hc2a0cc4a, 32'h4190c484} /* (28, 26, 5) {real, imag} */,
  {32'hc27eb666, 32'hc2a4f044} /* (28, 26, 4) {real, imag} */,
  {32'hc16f7136, 32'h426558a7} /* (28, 26, 3) {real, imag} */,
  {32'hc31e71ee, 32'hc2b8b38b} /* (28, 26, 2) {real, imag} */,
  {32'hc2d55c7b, 32'hc00a9750} /* (28, 26, 1) {real, imag} */,
  {32'hc25f8326, 32'h42f3a05f} /* (28, 26, 0) {real, imag} */,
  {32'hc36aa675, 32'h41be47cc} /* (28, 25, 31) {real, imag} */,
  {32'h4316ec3e, 32'hc1025e60} /* (28, 25, 30) {real, imag} */,
  {32'hc297e01a, 32'h4247858e} /* (28, 25, 29) {real, imag} */,
  {32'hc1757094, 32'h428a2517} /* (28, 25, 28) {real, imag} */,
  {32'hc2245b4e, 32'hc3081135} /* (28, 25, 27) {real, imag} */,
  {32'hc30e4d3c, 32'hc28562d6} /* (28, 25, 26) {real, imag} */,
  {32'h4305089d, 32'h42621c4c} /* (28, 25, 25) {real, imag} */,
  {32'hc0137cc0, 32'hc23766b0} /* (28, 25, 24) {real, imag} */,
  {32'h41f2e272, 32'h413dfefe} /* (28, 25, 23) {real, imag} */,
  {32'hc29db9b0, 32'hc2732022} /* (28, 25, 22) {real, imag} */,
  {32'h422a2a2a, 32'h422fd104} /* (28, 25, 21) {real, imag} */,
  {32'hc162c673, 32'h419f06b6} /* (28, 25, 20) {real, imag} */,
  {32'h41d1828e, 32'h3f4c77e0} /* (28, 25, 19) {real, imag} */,
  {32'h420d2124, 32'hc1cdf778} /* (28, 25, 18) {real, imag} */,
  {32'hc197ca50, 32'h41962801} /* (28, 25, 17) {real, imag} */,
  {32'h420a683f, 32'h419dc170} /* (28, 25, 16) {real, imag} */,
  {32'h41c126fc, 32'h4166606a} /* (28, 25, 15) {real, imag} */,
  {32'hc1aa7d3f, 32'hbf3e0100} /* (28, 25, 14) {real, imag} */,
  {32'hc0e688c8, 32'h426bd32e} /* (28, 25, 13) {real, imag} */,
  {32'h4215b438, 32'hc217359f} /* (28, 25, 12) {real, imag} */,
  {32'hc1006864, 32'h40e42a24} /* (28, 25, 11) {real, imag} */,
  {32'hc127a66c, 32'h40e0a1b0} /* (28, 25, 10) {real, imag} */,
  {32'h42acb57e, 32'hc2599f78} /* (28, 25, 9) {real, imag} */,
  {32'hc1233be8, 32'h41c59b88} /* (28, 25, 8) {real, imag} */,
  {32'hc26da894, 32'h4287fc2a} /* (28, 25, 7) {real, imag} */,
  {32'hc2939b44, 32'h420f8e54} /* (28, 25, 6) {real, imag} */,
  {32'hc1940c3e, 32'h4329599b} /* (28, 25, 5) {real, imag} */,
  {32'h4260141d, 32'hc2a1dd69} /* (28, 25, 4) {real, imag} */,
  {32'hc281e9be, 32'hc296d199} /* (28, 25, 3) {real, imag} */,
  {32'h42782954, 32'h42daf5ce} /* (28, 25, 2) {real, imag} */,
  {32'h41f39528, 32'hc30a9b04} /* (28, 25, 1) {real, imag} */,
  {32'hc29a4abe, 32'hc2b7b3c5} /* (28, 25, 0) {real, imag} */,
  {32'h439af01f, 32'h42cf3f30} /* (28, 24, 31) {real, imag} */,
  {32'hc2dd296c, 32'hc31fc012} /* (28, 24, 30) {real, imag} */,
  {32'hc1bf5f6e, 32'hc1d97164} /* (28, 24, 29) {real, imag} */,
  {32'h42f70dbb, 32'hc224669f} /* (28, 24, 28) {real, imag} */,
  {32'hc26e5782, 32'h432d9a5a} /* (28, 24, 27) {real, imag} */,
  {32'hc2bbaa15, 32'h420b434a} /* (28, 24, 26) {real, imag} */,
  {32'h42c36c0a, 32'hc2a5fd58} /* (28, 24, 25) {real, imag} */,
  {32'hc1536f94, 32'h4006c0d0} /* (28, 24, 24) {real, imag} */,
  {32'h420f5203, 32'h4127e3f8} /* (28, 24, 23) {real, imag} */,
  {32'hc207adaf, 32'hc119c556} /* (28, 24, 22) {real, imag} */,
  {32'hc1a06aec, 32'hc19a8202} /* (28, 24, 21) {real, imag} */,
  {32'hc2020bec, 32'h4274b0d3} /* (28, 24, 20) {real, imag} */,
  {32'hc2030436, 32'hc143c17c} /* (28, 24, 19) {real, imag} */,
  {32'h4222344d, 32'h415dcd87} /* (28, 24, 18) {real, imag} */,
  {32'h41f5275a, 32'h40602830} /* (28, 24, 17) {real, imag} */,
  {32'hc080fddc, 32'h41edf01a} /* (28, 24, 16) {real, imag} */,
  {32'hbf518b40, 32'hc001a570} /* (28, 24, 15) {real, imag} */,
  {32'hc16ad8ec, 32'h3f37ad90} /* (28, 24, 14) {real, imag} */,
  {32'hc1cf8500, 32'hc1500814} /* (28, 24, 13) {real, imag} */,
  {32'hc01c9d38, 32'hc1f1ced6} /* (28, 24, 12) {real, imag} */,
  {32'hc250756e, 32'hc2658679} /* (28, 24, 11) {real, imag} */,
  {32'h41be5ffc, 32'h41d30b35} /* (28, 24, 10) {real, imag} */,
  {32'h426429c5, 32'hc23b7c14} /* (28, 24, 9) {real, imag} */,
  {32'h423d2c6c, 32'hc0b22b48} /* (28, 24, 8) {real, imag} */,
  {32'h428e2e12, 32'h4292bc18} /* (28, 24, 7) {real, imag} */,
  {32'h41038688, 32'hc2706a4a} /* (28, 24, 6) {real, imag} */,
  {32'h42a905fb, 32'hc2f9fe90} /* (28, 24, 5) {real, imag} */,
  {32'h42e1ab45, 32'h42866790} /* (28, 24, 4) {real, imag} */,
  {32'hc2e5a048, 32'hc32e30d6} /* (28, 24, 3) {real, imag} */,
  {32'hc2b44780, 32'hc3001234} /* (28, 24, 2) {real, imag} */,
  {32'h43589cf6, 32'h434ac724} /* (28, 24, 1) {real, imag} */,
  {32'h4261f0f6, 32'h41eaf0ce} /* (28, 24, 0) {real, imag} */,
  {32'hc32aab20, 32'h420034d4} /* (28, 23, 31) {real, imag} */,
  {32'h42760ab6, 32'h420d5d08} /* (28, 23, 30) {real, imag} */,
  {32'hc2e669b5, 32'hc24ed022} /* (28, 23, 29) {real, imag} */,
  {32'hc209b9d6, 32'hc266601e} /* (28, 23, 28) {real, imag} */,
  {32'hc19a46c2, 32'hc1b28daf} /* (28, 23, 27) {real, imag} */,
  {32'h430d5354, 32'h42cbda98} /* (28, 23, 26) {real, imag} */,
  {32'hc0c58ee8, 32'hc2985ea8} /* (28, 23, 25) {real, imag} */,
  {32'hc2a8d5c2, 32'hc27a09af} /* (28, 23, 24) {real, imag} */,
  {32'hc1ae5a1a, 32'hc1f2c6e0} /* (28, 23, 23) {real, imag} */,
  {32'h422cc62a, 32'hc18c1ebd} /* (28, 23, 22) {real, imag} */,
  {32'h410780ae, 32'hc17e4332} /* (28, 23, 21) {real, imag} */,
  {32'h415125bc, 32'hc20f3090} /* (28, 23, 20) {real, imag} */,
  {32'h419eea4b, 32'hc15c881f} /* (28, 23, 19) {real, imag} */,
  {32'hc146c3a7, 32'h4150492d} /* (28, 23, 18) {real, imag} */,
  {32'h4182397f, 32'hc047fc24} /* (28, 23, 17) {real, imag} */,
  {32'h41712584, 32'h410cb538} /* (28, 23, 16) {real, imag} */,
  {32'h40ee16ec, 32'h418d4094} /* (28, 23, 15) {real, imag} */,
  {32'hc08c4532, 32'h4123d5dd} /* (28, 23, 14) {real, imag} */,
  {32'hc10aa946, 32'h41043679} /* (28, 23, 13) {real, imag} */,
  {32'hbf862a60, 32'hc0c151c2} /* (28, 23, 12) {real, imag} */,
  {32'h425e337a, 32'hc0e392a4} /* (28, 23, 11) {real, imag} */,
  {32'hc12bfd8e, 32'hc1d120ab} /* (28, 23, 10) {real, imag} */,
  {32'h4214d184, 32'hbfe4e540} /* (28, 23, 9) {real, imag} */,
  {32'h424ae03d, 32'h417ac66c} /* (28, 23, 8) {real, imag} */,
  {32'h422ee460, 32'h42163e2b} /* (28, 23, 7) {real, imag} */,
  {32'hc1874724, 32'h40e8df40} /* (28, 23, 6) {real, imag} */,
  {32'h424cee6b, 32'h422be578} /* (28, 23, 5) {real, imag} */,
  {32'hc328a928, 32'hc2a36873} /* (28, 23, 4) {real, imag} */,
  {32'h41363098, 32'h42270eb4} /* (28, 23, 3) {real, imag} */,
  {32'h428158d7, 32'hc28cd807} /* (28, 23, 2) {real, imag} */,
  {32'h4200df26, 32'h428a5565} /* (28, 23, 1) {real, imag} */,
  {32'hc241c04d, 32'h42625f0a} /* (28, 23, 0) {real, imag} */,
  {32'h410d952a, 32'hc09b664c} /* (28, 22, 31) {real, imag} */,
  {32'h43025771, 32'hc108a3d8} /* (28, 22, 30) {real, imag} */,
  {32'h42917ebc, 32'h423a0ff0} /* (28, 22, 29) {real, imag} */,
  {32'h42285058, 32'h4281e748} /* (28, 22, 28) {real, imag} */,
  {32'h421c5fcb, 32'hc219da17} /* (28, 22, 27) {real, imag} */,
  {32'hc21e2d45, 32'hc24bcc55} /* (28, 22, 26) {real, imag} */,
  {32'hc23658bb, 32'h4110c934} /* (28, 22, 25) {real, imag} */,
  {32'h4275dfd7, 32'h427cae09} /* (28, 22, 24) {real, imag} */,
  {32'h429f1636, 32'h4229b038} /* (28, 22, 23) {real, imag} */,
  {32'hc1937b72, 32'h3f49ab10} /* (28, 22, 22) {real, imag} */,
  {32'hc1a4a1d6, 32'hc0ebfbc6} /* (28, 22, 21) {real, imag} */,
  {32'hc1e550de, 32'hc19c9728} /* (28, 22, 20) {real, imag} */,
  {32'hc00e278c, 32'hc169e5c4} /* (28, 22, 19) {real, imag} */,
  {32'hc1203884, 32'h41a4c168} /* (28, 22, 18) {real, imag} */,
  {32'hc1fd8eb5, 32'hc02159e8} /* (28, 22, 17) {real, imag} */,
  {32'hc1084450, 32'h4151a6e0} /* (28, 22, 16) {real, imag} */,
  {32'h40d5e2e4, 32'hbedb1dc0} /* (28, 22, 15) {real, imag} */,
  {32'hc0240bf0, 32'hc14af578} /* (28, 22, 14) {real, imag} */,
  {32'h4082d8d6, 32'hc11d0b9e} /* (28, 22, 13) {real, imag} */,
  {32'h4152bfcc, 32'hc1c87cbc} /* (28, 22, 12) {real, imag} */,
  {32'h421159a1, 32'h41a8d722} /* (28, 22, 11) {real, imag} */,
  {32'hc0cc7a06, 32'h404d5cbc} /* (28, 22, 10) {real, imag} */,
  {32'h41d55c9e, 32'h42cab916} /* (28, 22, 9) {real, imag} */,
  {32'h4164b454, 32'h40046b90} /* (28, 22, 8) {real, imag} */,
  {32'hc21f5925, 32'hc241eda9} /* (28, 22, 7) {real, imag} */,
  {32'hc29661a0, 32'hc27a6443} /* (28, 22, 6) {real, imag} */,
  {32'hc1dd4042, 32'hc1a3569a} /* (28, 22, 5) {real, imag} */,
  {32'hc15dbf3a, 32'hc0a11f88} /* (28, 22, 4) {real, imag} */,
  {32'h42779b88, 32'h4194ba08} /* (28, 22, 3) {real, imag} */,
  {32'h4235c455, 32'hc2eb84b0} /* (28, 22, 2) {real, imag} */,
  {32'hc257de16, 32'h42619c18} /* (28, 22, 1) {real, imag} */,
  {32'hc2b398d0, 32'h409a872c} /* (28, 22, 0) {real, imag} */,
  {32'h431e31ae, 32'h41349cb6} /* (28, 21, 31) {real, imag} */,
  {32'h4186f4e4, 32'h42e556c3} /* (28, 21, 30) {real, imag} */,
  {32'h42bab4df, 32'hc122b6f5} /* (28, 21, 29) {real, imag} */,
  {32'hc02c2870, 32'hc1873b06} /* (28, 21, 28) {real, imag} */,
  {32'hc2c7d1a3, 32'h420dba6b} /* (28, 21, 27) {real, imag} */,
  {32'hc16f6492, 32'h4231f25c} /* (28, 21, 26) {real, imag} */,
  {32'hc1907aec, 32'h415a62de} /* (28, 21, 25) {real, imag} */,
  {32'hc1d42712, 32'hc185c662} /* (28, 21, 24) {real, imag} */,
  {32'hc19f2d31, 32'hc1ae3dff} /* (28, 21, 23) {real, imag} */,
  {32'hc11d3c06, 32'hc243c104} /* (28, 21, 22) {real, imag} */,
  {32'h418fa62a, 32'h409906da} /* (28, 21, 21) {real, imag} */,
  {32'h3e7e5840, 32'hbeb09ec0} /* (28, 21, 20) {real, imag} */,
  {32'hc1c817af, 32'hc0cb48b2} /* (28, 21, 19) {real, imag} */,
  {32'hc1a0b5a8, 32'h4154300e} /* (28, 21, 18) {real, imag} */,
  {32'h40c08274, 32'hc1a9633f} /* (28, 21, 17) {real, imag} */,
  {32'h412e8200, 32'h413e5bbb} /* (28, 21, 16) {real, imag} */,
  {32'hc164df12, 32'h40dd0df3} /* (28, 21, 15) {real, imag} */,
  {32'h410e5edc, 32'hc162f55e} /* (28, 21, 14) {real, imag} */,
  {32'hc2007186, 32'h419582de} /* (28, 21, 13) {real, imag} */,
  {32'hc1faf00c, 32'hc23236ba} /* (28, 21, 12) {real, imag} */,
  {32'hc1b22704, 32'h41064e55} /* (28, 21, 11) {real, imag} */,
  {32'h422d1540, 32'h4128e39e} /* (28, 21, 10) {real, imag} */,
  {32'hc2008a9a, 32'hc1921163} /* (28, 21, 9) {real, imag} */,
  {32'h40f1fdaa, 32'hc238bd51} /* (28, 21, 8) {real, imag} */,
  {32'hc0c2ee5e, 32'h42142022} /* (28, 21, 7) {real, imag} */,
  {32'h4232c6ce, 32'h41a1320d} /* (28, 21, 6) {real, imag} */,
  {32'h408e0db0, 32'h41ad1626} /* (28, 21, 5) {real, imag} */,
  {32'h42238715, 32'h409eef0e} /* (28, 21, 4) {real, imag} */,
  {32'hc2009342, 32'hc21c7290} /* (28, 21, 3) {real, imag} */,
  {32'hc2d435e9, 32'h4216f782} /* (28, 21, 2) {real, imag} */,
  {32'h4283bb7c, 32'h41d5b101} /* (28, 21, 1) {real, imag} */,
  {32'h42379e16, 32'h41a870ba} /* (28, 21, 0) {real, imag} */,
  {32'hc131b634, 32'h41540cb4} /* (28, 20, 31) {real, imag} */,
  {32'h42098d7f, 32'h4268ec54} /* (28, 20, 30) {real, imag} */,
  {32'hc1d23143, 32'h41cf7982} /* (28, 20, 29) {real, imag} */,
  {32'h421b8e9e, 32'hc1ce89d4} /* (28, 20, 28) {real, imag} */,
  {32'hc1aebde7, 32'hbf3042c0} /* (28, 20, 27) {real, imag} */,
  {32'hbe680d00, 32'hc21f3c63} /* (28, 20, 26) {real, imag} */,
  {32'hc20da6d2, 32'hc2406320} /* (28, 20, 25) {real, imag} */,
  {32'hc2101e47, 32'h4225fba8} /* (28, 20, 24) {real, imag} */,
  {32'hc2731cc2, 32'hbf86c658} /* (28, 20, 23) {real, imag} */,
  {32'hc19350e2, 32'h40fe7a2c} /* (28, 20, 22) {real, imag} */,
  {32'hc150d738, 32'h41d315ca} /* (28, 20, 21) {real, imag} */,
  {32'h416405ed, 32'h410f672d} /* (28, 20, 20) {real, imag} */,
  {32'hc1eaf478, 32'hc0811c2c} /* (28, 20, 19) {real, imag} */,
  {32'h401d5798, 32'hc11aaf2f} /* (28, 20, 18) {real, imag} */,
  {32'h40d695a4, 32'hc0b13f36} /* (28, 20, 17) {real, imag} */,
  {32'hc02076a8, 32'hc03fd65c} /* (28, 20, 16) {real, imag} */,
  {32'h40705870, 32'hbfe72508} /* (28, 20, 15) {real, imag} */,
  {32'h41e5678d, 32'h41724e03} /* (28, 20, 14) {real, imag} */,
  {32'hc006a634, 32'hc11f7d80} /* (28, 20, 13) {real, imag} */,
  {32'hc1003407, 32'h41d3e6f2} /* (28, 20, 12) {real, imag} */,
  {32'h3d7f0a80, 32'hc1d256b2} /* (28, 20, 11) {real, imag} */,
  {32'h4128bde7, 32'hc241e6a8} /* (28, 20, 10) {real, imag} */,
  {32'hc1a79967, 32'hc1c4fd78} /* (28, 20, 9) {real, imag} */,
  {32'hc178f61f, 32'hc08cbf60} /* (28, 20, 8) {real, imag} */,
  {32'h408baf7c, 32'hc1eda0b8} /* (28, 20, 7) {real, imag} */,
  {32'h4296cbba, 32'h422f654d} /* (28, 20, 6) {real, imag} */,
  {32'h41d9b28d, 32'h4284b788} /* (28, 20, 5) {real, imag} */,
  {32'h41af7860, 32'hc1194121} /* (28, 20, 4) {real, imag} */,
  {32'h418dba75, 32'hc1be85c2} /* (28, 20, 3) {real, imag} */,
  {32'h4138b9c4, 32'hc1ca5db5} /* (28, 20, 2) {real, imag} */,
  {32'hc2406b13, 32'h4284a56e} /* (28, 20, 1) {real, imag} */,
  {32'hc206e686, 32'h41a8e6b4} /* (28, 20, 0) {real, imag} */,
  {32'hc1507e0f, 32'hc29913a3} /* (28, 19, 31) {real, imag} */,
  {32'h42053c1a, 32'hc20deb67} /* (28, 19, 30) {real, imag} */,
  {32'hc15e242d, 32'hc1b1fa38} /* (28, 19, 29) {real, imag} */,
  {32'hc195d6e6, 32'hc1e71617} /* (28, 19, 28) {real, imag} */,
  {32'h3ed73680, 32'h42253773} /* (28, 19, 27) {real, imag} */,
  {32'h41151454, 32'hc228c8a4} /* (28, 19, 26) {real, imag} */,
  {32'h3f906948, 32'hc1c7a6cd} /* (28, 19, 25) {real, imag} */,
  {32'h4104b47a, 32'h42761f4c} /* (28, 19, 24) {real, imag} */,
  {32'h414c0efb, 32'hc1893ce7} /* (28, 19, 23) {real, imag} */,
  {32'h41e5a762, 32'h4186f0d0} /* (28, 19, 22) {real, imag} */,
  {32'hc044f5e0, 32'hc18f237c} /* (28, 19, 21) {real, imag} */,
  {32'hc0916d0a, 32'h407c1d70} /* (28, 19, 20) {real, imag} */,
  {32'hc1ab32f0, 32'h410afdeb} /* (28, 19, 19) {real, imag} */,
  {32'hc10c1c3d, 32'hc10e365a} /* (28, 19, 18) {real, imag} */,
  {32'hbfdbc7e0, 32'h3fa11cf8} /* (28, 19, 17) {real, imag} */,
  {32'hc09dfff0, 32'hbf696e80} /* (28, 19, 16) {real, imag} */,
  {32'h410b33e2, 32'h4095e072} /* (28, 19, 15) {real, imag} */,
  {32'hc14eadb9, 32'h40c8ab7c} /* (28, 19, 14) {real, imag} */,
  {32'h41bc0950, 32'hbfa35d58} /* (28, 19, 13) {real, imag} */,
  {32'h41402f1f, 32'hc1a59862} /* (28, 19, 12) {real, imag} */,
  {32'h408fa300, 32'h40ebd20c} /* (28, 19, 11) {real, imag} */,
  {32'hc09ff11a, 32'hc09eec46} /* (28, 19, 10) {real, imag} */,
  {32'h41b56de6, 32'h417fa6b2} /* (28, 19, 9) {real, imag} */,
  {32'hc1b22519, 32'hc10f2562} /* (28, 19, 8) {real, imag} */,
  {32'hc1b83b94, 32'hc20b708c} /* (28, 19, 7) {real, imag} */,
  {32'h42366ab3, 32'hc134a2a3} /* (28, 19, 6) {real, imag} */,
  {32'h42377ed7, 32'h3fcb9860} /* (28, 19, 5) {real, imag} */,
  {32'h41a44e0c, 32'hc245e86c} /* (28, 19, 4) {real, imag} */,
  {32'hc15c857b, 32'hc20b36d0} /* (28, 19, 3) {real, imag} */,
  {32'hc1621ad9, 32'h4258a92b} /* (28, 19, 2) {real, imag} */,
  {32'hc1a87538, 32'hc232f62f} /* (28, 19, 1) {real, imag} */,
  {32'hc28f88db, 32'h422572f1} /* (28, 19, 0) {real, imag} */,
  {32'h42542fee, 32'hc1ddf8c0} /* (28, 18, 31) {real, imag} */,
  {32'hc210f74a, 32'h42852984} /* (28, 18, 30) {real, imag} */,
  {32'hc17e4aaa, 32'hc103a61c} /* (28, 18, 29) {real, imag} */,
  {32'h422bea1e, 32'h410219a2} /* (28, 18, 28) {real, imag} */,
  {32'hc18e4bce, 32'h40242894} /* (28, 18, 27) {real, imag} */,
  {32'h414800a6, 32'hc1c66292} /* (28, 18, 26) {real, imag} */,
  {32'hc1a0dd64, 32'h41bea639} /* (28, 18, 25) {real, imag} */,
  {32'h4125bd17, 32'hc1d5ce8f} /* (28, 18, 24) {real, imag} */,
  {32'hc0ac0f5a, 32'h41a30709} /* (28, 18, 23) {real, imag} */,
  {32'h40779cfc, 32'h3ea15e80} /* (28, 18, 22) {real, imag} */,
  {32'h4122b004, 32'h4159f99a} /* (28, 18, 21) {real, imag} */,
  {32'hbf197d90, 32'hc11f3b4e} /* (28, 18, 20) {real, imag} */,
  {32'hbfd04fb8, 32'hbff2c760} /* (28, 18, 19) {real, imag} */,
  {32'hc0e08806, 32'hc110a293} /* (28, 18, 18) {real, imag} */,
  {32'hbf556610, 32'h40f8d043} /* (28, 18, 17) {real, imag} */,
  {32'hbfc024e4, 32'hc10743f1} /* (28, 18, 16) {real, imag} */,
  {32'h40c1c102, 32'hc0a10d9d} /* (28, 18, 15) {real, imag} */,
  {32'hc032db64, 32'hc183d7be} /* (28, 18, 14) {real, imag} */,
  {32'h408e093c, 32'h41b71026} /* (28, 18, 13) {real, imag} */,
  {32'hc19edacc, 32'h4063cfec} /* (28, 18, 12) {real, imag} */,
  {32'h3ff9a24c, 32'h4142dad4} /* (28, 18, 11) {real, imag} */,
  {32'hbf7bdc90, 32'h41c35459} /* (28, 18, 10) {real, imag} */,
  {32'hbfe08756, 32'hc14fb89a} /* (28, 18, 9) {real, imag} */,
  {32'h41eed788, 32'h41b2c833} /* (28, 18, 8) {real, imag} */,
  {32'h41d8d510, 32'hc1cd0771} /* (28, 18, 7) {real, imag} */,
  {32'h41a37259, 32'hc161ef0b} /* (28, 18, 6) {real, imag} */,
  {32'hc16b4bb4, 32'hc1b9e8f4} /* (28, 18, 5) {real, imag} */,
  {32'h41785d5a, 32'h41eae925} /* (28, 18, 4) {real, imag} */,
  {32'h4029f1b6, 32'h412e54d8} /* (28, 18, 3) {real, imag} */,
  {32'h40e4ffec, 32'hc11c618c} /* (28, 18, 2) {real, imag} */,
  {32'h42aa78b1, 32'h3f0c4480} /* (28, 18, 1) {real, imag} */,
  {32'h41601858, 32'hc1bc2bb8} /* (28, 18, 0) {real, imag} */,
  {32'hc27e1c20, 32'hc1b7d518} /* (28, 17, 31) {real, imag} */,
  {32'h41f88291, 32'hc16abbf8} /* (28, 17, 30) {real, imag} */,
  {32'hc206d180, 32'hc1e10f8c} /* (28, 17, 29) {real, imag} */,
  {32'h40f1cbc6, 32'hc21d48af} /* (28, 17, 28) {real, imag} */,
  {32'h4234854b, 32'h418bfc5e} /* (28, 17, 27) {real, imag} */,
  {32'h41d1a697, 32'hc093d6ec} /* (28, 17, 26) {real, imag} */,
  {32'h3e98e140, 32'h41e7d810} /* (28, 17, 25) {real, imag} */,
  {32'h409209a6, 32'h40e2d1dc} /* (28, 17, 24) {real, imag} */,
  {32'h40e91896, 32'h4198c08e} /* (28, 17, 23) {real, imag} */,
  {32'h4098faa6, 32'hc0e24f9e} /* (28, 17, 22) {real, imag} */,
  {32'hc1d3849a, 32'hc104588e} /* (28, 17, 21) {real, imag} */,
  {32'hc110c6c6, 32'hc136043a} /* (28, 17, 20) {real, imag} */,
  {32'hbebc2210, 32'h3f869b30} /* (28, 17, 19) {real, imag} */,
  {32'h40f60c0c, 32'hbf12c578} /* (28, 17, 18) {real, imag} */,
  {32'hc0051bac, 32'hbfb68f86} /* (28, 17, 17) {real, imag} */,
  {32'h3f695a00, 32'hc0c137ee} /* (28, 17, 16) {real, imag} */,
  {32'h409a3646, 32'h4070f963} /* (28, 17, 15) {real, imag} */,
  {32'hbfbe5c20, 32'hc0a1de45} /* (28, 17, 14) {real, imag} */,
  {32'hc0d8cabf, 32'hc0a83e98} /* (28, 17, 13) {real, imag} */,
  {32'h4108599e, 32'h4033a55e} /* (28, 17, 12) {real, imag} */,
  {32'hc1eac92a, 32'hc05864fe} /* (28, 17, 11) {real, imag} */,
  {32'h41d5293c, 32'h413905d5} /* (28, 17, 10) {real, imag} */,
  {32'h420730b9, 32'h418ecd84} /* (28, 17, 9) {real, imag} */,
  {32'h41ef7a36, 32'h42463678} /* (28, 17, 8) {real, imag} */,
  {32'h4215e1ce, 32'hc0e53a18} /* (28, 17, 7) {real, imag} */,
  {32'hc0ee8574, 32'hc1ffe3e1} /* (28, 17, 6) {real, imag} */,
  {32'hbfe86f20, 32'h4097b5a6} /* (28, 17, 5) {real, imag} */,
  {32'hc211a4cb, 32'h41f35d76} /* (28, 17, 4) {real, imag} */,
  {32'hc23499d8, 32'h418cd228} /* (28, 17, 3) {real, imag} */,
  {32'hbe279900, 32'hc2219a16} /* (28, 17, 2) {real, imag} */,
  {32'hc1cd36ec, 32'hc1404281} /* (28, 17, 1) {real, imag} */,
  {32'hc18e07ce, 32'h4075556c} /* (28, 17, 0) {real, imag} */,
  {32'h41d840dd, 32'hc02b7111} /* (28, 16, 31) {real, imag} */,
  {32'h409f5fda, 32'hc1d08f45} /* (28, 16, 30) {real, imag} */,
  {32'hc215d25d, 32'h402f2c28} /* (28, 16, 29) {real, imag} */,
  {32'h41145f97, 32'h4231f3b8} /* (28, 16, 28) {real, imag} */,
  {32'hc1d7413b, 32'hc1b462c7} /* (28, 16, 27) {real, imag} */,
  {32'h4184f2a9, 32'h42066b95} /* (28, 16, 26) {real, imag} */,
  {32'h418ca150, 32'h410c4ecf} /* (28, 16, 25) {real, imag} */,
  {32'hc0c5f988, 32'h411e7454} /* (28, 16, 24) {real, imag} */,
  {32'hc11c7eb1, 32'hc0c372da} /* (28, 16, 23) {real, imag} */,
  {32'hc1684eea, 32'hbed9d108} /* (28, 16, 22) {real, imag} */,
  {32'hc048c4e2, 32'hc15feb16} /* (28, 16, 21) {real, imag} */,
  {32'hc1114f35, 32'h40978e6a} /* (28, 16, 20) {real, imag} */,
  {32'h41f43630, 32'hbeb01d40} /* (28, 16, 19) {real, imag} */,
  {32'hc04d1943, 32'hc0dd7bf4} /* (28, 16, 18) {real, imag} */,
  {32'hc0d63fa3, 32'hc042e35f} /* (28, 16, 17) {real, imag} */,
  {32'h414b95f8, 32'h3f880160} /* (28, 16, 16) {real, imag} */,
  {32'hc0296902, 32'hc05772cd} /* (28, 16, 15) {real, imag} */,
  {32'hc0d17064, 32'hc08a4414} /* (28, 16, 14) {real, imag} */,
  {32'hc0c015a6, 32'hc1445a24} /* (28, 16, 13) {real, imag} */,
  {32'h408336c4, 32'h4099201e} /* (28, 16, 12) {real, imag} */,
  {32'h412e77b8, 32'hc08680c4} /* (28, 16, 11) {real, imag} */,
  {32'hc10630a0, 32'hc0cd8e90} /* (28, 16, 10) {real, imag} */,
  {32'hc1b880b4, 32'hc127b853} /* (28, 16, 9) {real, imag} */,
  {32'hc0cc0988, 32'hc1db2132} /* (28, 16, 8) {real, imag} */,
  {32'hc12bea6a, 32'hc18b3990} /* (28, 16, 7) {real, imag} */,
  {32'h40c3ba59, 32'hc1bc9ed2} /* (28, 16, 6) {real, imag} */,
  {32'hc258f2c6, 32'h403f4ab8} /* (28, 16, 5) {real, imag} */,
  {32'hc0bd3bc4, 32'h4215f2c0} /* (28, 16, 4) {real, imag} */,
  {32'h418492bc, 32'hc1e2cf56} /* (28, 16, 3) {real, imag} */,
  {32'h4189ff48, 32'h41b007eb} /* (28, 16, 2) {real, imag} */,
  {32'h41eae03b, 32'hc0b18aa2} /* (28, 16, 1) {real, imag} */,
  {32'h4148e448, 32'hc26c5683} /* (28, 16, 0) {real, imag} */,
  {32'h40a52472, 32'hc14aacef} /* (28, 15, 31) {real, imag} */,
  {32'h412951e5, 32'hc13ce4f8} /* (28, 15, 30) {real, imag} */,
  {32'h3fbbdecc, 32'hc283c130} /* (28, 15, 29) {real, imag} */,
  {32'h41988a52, 32'h414dcc02} /* (28, 15, 28) {real, imag} */,
  {32'h41f2bc76, 32'hc05600f8} /* (28, 15, 27) {real, imag} */,
  {32'h414a740c, 32'h423ac4f4} /* (28, 15, 26) {real, imag} */,
  {32'hc0cb1b59, 32'h418c32bc} /* (28, 15, 25) {real, imag} */,
  {32'hc11e6645, 32'hc1e8647d} /* (28, 15, 24) {real, imag} */,
  {32'h402ebb25, 32'hc135c6ef} /* (28, 15, 23) {real, imag} */,
  {32'hc0026d34, 32'hc04f15fc} /* (28, 15, 22) {real, imag} */,
  {32'hc1146371, 32'hbde79880} /* (28, 15, 21) {real, imag} */,
  {32'h41bafeb5, 32'h404deaf4} /* (28, 15, 20) {real, imag} */,
  {32'hc109d352, 32'h41a2af53} /* (28, 15, 19) {real, imag} */,
  {32'h40aeb2ea, 32'h40d541ea} /* (28, 15, 18) {real, imag} */,
  {32'h3f885f60, 32'hc14c98b2} /* (28, 15, 17) {real, imag} */,
  {32'hc075b496, 32'hbf5edc80} /* (28, 15, 16) {real, imag} */,
  {32'h40df1c8c, 32'hc05de1b0} /* (28, 15, 15) {real, imag} */,
  {32'h4154ba55, 32'h3fc9d1f0} /* (28, 15, 14) {real, imag} */,
  {32'h41010a84, 32'h40900d84} /* (28, 15, 13) {real, imag} */,
  {32'hc147f59e, 32'hc191e5ee} /* (28, 15, 12) {real, imag} */,
  {32'h41e0f5c4, 32'hc13a5376} /* (28, 15, 11) {real, imag} */,
  {32'hc0bf989e, 32'h3eb96a60} /* (28, 15, 10) {real, imag} */,
  {32'hc115b7eb, 32'hc11569bb} /* (28, 15, 9) {real, imag} */,
  {32'hc15e0af7, 32'hc1de61a7} /* (28, 15, 8) {real, imag} */,
  {32'hc11c1abe, 32'h420059d8} /* (28, 15, 7) {real, imag} */,
  {32'hc1947571, 32'h412421ae} /* (28, 15, 6) {real, imag} */,
  {32'hc12ba6bd, 32'h41d78fff} /* (28, 15, 5) {real, imag} */,
  {32'h410dc397, 32'h417df720} /* (28, 15, 4) {real, imag} */,
  {32'hc1873f22, 32'h42449480} /* (28, 15, 3) {real, imag} */,
  {32'h40a0d90a, 32'h40a878a7} /* (28, 15, 2) {real, imag} */,
  {32'h42141b30, 32'hc21346f8} /* (28, 15, 1) {real, imag} */,
  {32'hc150c096, 32'h420dec9c} /* (28, 15, 0) {real, imag} */,
  {32'hc288b9a8, 32'h40b6c586} /* (28, 14, 31) {real, imag} */,
  {32'h419882e0, 32'h41438b20} /* (28, 14, 30) {real, imag} */,
  {32'h40f18352, 32'h418a8004} /* (28, 14, 29) {real, imag} */,
  {32'h41e4f0b6, 32'hc10d15ea} /* (28, 14, 28) {real, imag} */,
  {32'hc12e0e42, 32'h406d72df} /* (28, 14, 27) {real, imag} */,
  {32'h425fe590, 32'hc23c1499} /* (28, 14, 26) {real, imag} */,
  {32'hc2085c10, 32'hbea2df90} /* (28, 14, 25) {real, imag} */,
  {32'hc1b941a2, 32'h419d422e} /* (28, 14, 24) {real, imag} */,
  {32'h412e2cb6, 32'h40f2d43e} /* (28, 14, 23) {real, imag} */,
  {32'h4112257c, 32'h4199eb18} /* (28, 14, 22) {real, imag} */,
  {32'hc10a6d14, 32'h40eb4c34} /* (28, 14, 21) {real, imag} */,
  {32'h412850f2, 32'h4101127e} /* (28, 14, 20) {real, imag} */,
  {32'h411d3a4f, 32'hc0a3ae9f} /* (28, 14, 19) {real, imag} */,
  {32'hc0b56c80, 32'h41211f10} /* (28, 14, 18) {real, imag} */,
  {32'hc04f7c82, 32'h40f6afa2} /* (28, 14, 17) {real, imag} */,
  {32'hc04f9d48, 32'h409366b2} /* (28, 14, 16) {real, imag} */,
  {32'hc13ab164, 32'hc11cf10d} /* (28, 14, 15) {real, imag} */,
  {32'h40182838, 32'h3fe049f0} /* (28, 14, 14) {real, imag} */,
  {32'hc0b86cea, 32'hbbb54400} /* (28, 14, 13) {real, imag} */,
  {32'hc05f970e, 32'h3c90d300} /* (28, 14, 12) {real, imag} */,
  {32'h4149e050, 32'hc09195a6} /* (28, 14, 11) {real, imag} */,
  {32'hc234699a, 32'hc1b26794} /* (28, 14, 10) {real, imag} */,
  {32'h401c9bd0, 32'hc17b59b9} /* (28, 14, 9) {real, imag} */,
  {32'hc1f81cac, 32'hc1a10a3a} /* (28, 14, 8) {real, imag} */,
  {32'h41a750f4, 32'h40f3aa25} /* (28, 14, 7) {real, imag} */,
  {32'h42135220, 32'hc1955e4a} /* (28, 14, 6) {real, imag} */,
  {32'h41f48f75, 32'hc021e45d} /* (28, 14, 5) {real, imag} */,
  {32'h41e44f1a, 32'h41e933a5} /* (28, 14, 4) {real, imag} */,
  {32'h409eb44a, 32'hc194d078} /* (28, 14, 3) {real, imag} */,
  {32'h41e8b6e4, 32'hc2564630} /* (28, 14, 2) {real, imag} */,
  {32'h4212e12b, 32'h4209ead3} /* (28, 14, 1) {real, imag} */,
  {32'hc243eff4, 32'h42043efe} /* (28, 14, 0) {real, imag} */,
  {32'h41aa9332, 32'h408b32b8} /* (28, 13, 31) {real, imag} */,
  {32'hc1f86896, 32'h4238eb5a} /* (28, 13, 30) {real, imag} */,
  {32'h4246fa06, 32'h402aeb1c} /* (28, 13, 29) {real, imag} */,
  {32'hc0d6e870, 32'hc0104da8} /* (28, 13, 28) {real, imag} */,
  {32'h41a01ff9, 32'h413762b0} /* (28, 13, 27) {real, imag} */,
  {32'h40326250, 32'hc108f108} /* (28, 13, 26) {real, imag} */,
  {32'hbfb1d7ec, 32'h4204b992} /* (28, 13, 25) {real, imag} */,
  {32'h41619611, 32'h40df9b08} /* (28, 13, 24) {real, imag} */,
  {32'hc188e456, 32'hc08758bb} /* (28, 13, 23) {real, imag} */,
  {32'hc2214259, 32'h3fe0eb30} /* (28, 13, 22) {real, imag} */,
  {32'hc1fd7c1e, 32'hc15023d4} /* (28, 13, 21) {real, imag} */,
  {32'h40b5da12, 32'hc13b02e8} /* (28, 13, 20) {real, imag} */,
  {32'hc15f99d6, 32'h4171bbac} /* (28, 13, 19) {real, imag} */,
  {32'hbe961460, 32'h41a3f522} /* (28, 13, 18) {real, imag} */,
  {32'h40ae6b86, 32'h41711fa6} /* (28, 13, 17) {real, imag} */,
  {32'h4126a8f8, 32'hc11b06d7} /* (28, 13, 16) {real, imag} */,
  {32'h3e194bd0, 32'h4131b462} /* (28, 13, 15) {real, imag} */,
  {32'hc08209d2, 32'hc086843c} /* (28, 13, 14) {real, imag} */,
  {32'h40b92ff4, 32'hbfe7b114} /* (28, 13, 13) {real, imag} */,
  {32'hc0f03c42, 32'h41205d44} /* (28, 13, 12) {real, imag} */,
  {32'hc1290814, 32'h40a8cffc} /* (28, 13, 11) {real, imag} */,
  {32'h41d118e7, 32'h41f8ccc9} /* (28, 13, 10) {real, imag} */,
  {32'hc18d205a, 32'hc02e136a} /* (28, 13, 9) {real, imag} */,
  {32'h421cabe7, 32'hc1a35310} /* (28, 13, 8) {real, imag} */,
  {32'h40eb0031, 32'h41c9082f} /* (28, 13, 7) {real, imag} */,
  {32'h42120d58, 32'hc090f261} /* (28, 13, 6) {real, imag} */,
  {32'hc08f9185, 32'h425235de} /* (28, 13, 5) {real, imag} */,
  {32'hc2395ece, 32'hc268e54c} /* (28, 13, 4) {real, imag} */,
  {32'h4206eb2a, 32'h41e45c0a} /* (28, 13, 3) {real, imag} */,
  {32'hc24b999d, 32'hc1834668} /* (28, 13, 2) {real, imag} */,
  {32'hc1337084, 32'hc21453bb} /* (28, 13, 1) {real, imag} */,
  {32'h424382bd, 32'hc0e21602} /* (28, 13, 0) {real, imag} */,
  {32'hc2004123, 32'h413b3934} /* (28, 12, 31) {real, imag} */,
  {32'h430d5c10, 32'hc079bdcd} /* (28, 12, 30) {real, imag} */,
  {32'hc073f1f0, 32'hc23019a4} /* (28, 12, 29) {real, imag} */,
  {32'hc1aab72f, 32'hc1321fdc} /* (28, 12, 28) {real, imag} */,
  {32'hc1f68674, 32'hc2b45424} /* (28, 12, 27) {real, imag} */,
  {32'h419b597e, 32'hc15bacdd} /* (28, 12, 26) {real, imag} */,
  {32'h41b01484, 32'h42047006} /* (28, 12, 25) {real, imag} */,
  {32'hc24ec5aa, 32'hc0edc880} /* (28, 12, 24) {real, imag} */,
  {32'h4071a473, 32'h41c5f7b0} /* (28, 12, 23) {real, imag} */,
  {32'h4015456e, 32'h4230ed9a} /* (28, 12, 22) {real, imag} */,
  {32'hc1419aec, 32'hc2384e1a} /* (28, 12, 21) {real, imag} */,
  {32'hc0e0893e, 32'h41837368} /* (28, 12, 20) {real, imag} */,
  {32'h408a02d6, 32'h4127b1b6} /* (28, 12, 19) {real, imag} */,
  {32'hc104b614, 32'h4167fe0a} /* (28, 12, 18) {real, imag} */,
  {32'hc1029be2, 32'hc1871f2b} /* (28, 12, 17) {real, imag} */,
  {32'h3fc467e0, 32'hc0c13ff8} /* (28, 12, 16) {real, imag} */,
  {32'hc0e8a2f4, 32'h4142592a} /* (28, 12, 15) {real, imag} */,
  {32'hc051dd90, 32'h413080ae} /* (28, 12, 14) {real, imag} */,
  {32'hc19f6952, 32'hbf151d20} /* (28, 12, 13) {real, imag} */,
  {32'hc0101ff8, 32'hc172fa44} /* (28, 12, 12) {real, imag} */,
  {32'h411e010e, 32'h40d2891c} /* (28, 12, 11) {real, imag} */,
  {32'h40adc74d, 32'h40d0b220} /* (28, 12, 10) {real, imag} */,
  {32'hc015c80b, 32'hc1e374ee} /* (28, 12, 9) {real, imag} */,
  {32'h420f2090, 32'h41f8b868} /* (28, 12, 8) {real, imag} */,
  {32'h41878914, 32'hc129b9fe} /* (28, 12, 7) {real, imag} */,
  {32'h40d077fd, 32'hc1494ba5} /* (28, 12, 6) {real, imag} */,
  {32'h411dcef1, 32'h4249ddb8} /* (28, 12, 5) {real, imag} */,
  {32'hc0e3dbfb, 32'hc1e777c8} /* (28, 12, 4) {real, imag} */,
  {32'hc2402bfb, 32'hc1985ccf} /* (28, 12, 3) {real, imag} */,
  {32'h3fded940, 32'hbe32de70} /* (28, 12, 2) {real, imag} */,
  {32'h422882d7, 32'hc1baf9d6} /* (28, 12, 1) {real, imag} */,
  {32'h420bfdc7, 32'h41b33d36} /* (28, 12, 0) {real, imag} */,
  {32'h40e5028c, 32'h428c3900} /* (28, 11, 31) {real, imag} */,
  {32'h42e971b9, 32'hc20eb975} /* (28, 11, 30) {real, imag} */,
  {32'h41f2c277, 32'h423b4a5e} /* (28, 11, 29) {real, imag} */,
  {32'h40fcfd4b, 32'h412424f7} /* (28, 11, 28) {real, imag} */,
  {32'hc1a23467, 32'hc2956090} /* (28, 11, 27) {real, imag} */,
  {32'h423a3a0e, 32'hc1b85cde} /* (28, 11, 26) {real, imag} */,
  {32'hc18eae0a, 32'h4234d8f0} /* (28, 11, 25) {real, imag} */,
  {32'h41a494a2, 32'h417a7876} /* (28, 11, 24) {real, imag} */,
  {32'h41d6d7bc, 32'hc1847f15} /* (28, 11, 23) {real, imag} */,
  {32'hc1ab1dd5, 32'h41ee88fa} /* (28, 11, 22) {real, imag} */,
  {32'h41185294, 32'hc166ec66} /* (28, 11, 21) {real, imag} */,
  {32'h40f88ec1, 32'h3f4ea8b0} /* (28, 11, 20) {real, imag} */,
  {32'hc1570cc2, 32'hc08884b8} /* (28, 11, 19) {real, imag} */,
  {32'h413ce3ac, 32'h3f5786d0} /* (28, 11, 18) {real, imag} */,
  {32'hc10e0bb6, 32'h40dbcb92} /* (28, 11, 17) {real, imag} */,
  {32'h41a1ea46, 32'h411f3cd4} /* (28, 11, 16) {real, imag} */,
  {32'h40e624a4, 32'h40583d4c} /* (28, 11, 15) {real, imag} */,
  {32'hc0b8a038, 32'h4002403c} /* (28, 11, 14) {real, imag} */,
  {32'hbf78c720, 32'hc1a41826} /* (28, 11, 13) {real, imag} */,
  {32'h413a7344, 32'hc11ee2c7} /* (28, 11, 12) {real, imag} */,
  {32'h41147e2c, 32'h419d9009} /* (28, 11, 11) {real, imag} */,
  {32'hc2184bce, 32'h41c76892} /* (28, 11, 10) {real, imag} */,
  {32'hc1605a04, 32'hc06a90c8} /* (28, 11, 9) {real, imag} */,
  {32'hc1d85dd6, 32'h41f0b739} /* (28, 11, 8) {real, imag} */,
  {32'hc1cfc34c, 32'hc20eb656} /* (28, 11, 7) {real, imag} */,
  {32'h420ad97a, 32'h41160b03} /* (28, 11, 6) {real, imag} */,
  {32'h41e6b351, 32'hc21cb460} /* (28, 11, 5) {real, imag} */,
  {32'h4109132b, 32'h42013432} /* (28, 11, 4) {real, imag} */,
  {32'hc29fb8a7, 32'hc28d10e9} /* (28, 11, 3) {real, imag} */,
  {32'h43189d6c, 32'hc1fbbc26} /* (28, 11, 2) {real, imag} */,
  {32'hc255d4f2, 32'h4191e996} /* (28, 11, 1) {real, imag} */,
  {32'hc2cb9d0a, 32'h42463f29} /* (28, 11, 0) {real, imag} */,
  {32'hc201589e, 32'hc2563cf6} /* (28, 10, 31) {real, imag} */,
  {32'hc2640ef3, 32'h42f5b14c} /* (28, 10, 30) {real, imag} */,
  {32'hc2934b9f, 32'hc28f9f5a} /* (28, 10, 29) {real, imag} */,
  {32'hc26be6b0, 32'hc20871e9} /* (28, 10, 28) {real, imag} */,
  {32'hc0f8a7e4, 32'hc1175a5a} /* (28, 10, 27) {real, imag} */,
  {32'hc1724fc0, 32'hc13753dc} /* (28, 10, 26) {real, imag} */,
  {32'h41b4ac0b, 32'hc1d714bf} /* (28, 10, 25) {real, imag} */,
  {32'hc1895b70, 32'hc140f97a} /* (28, 10, 24) {real, imag} */,
  {32'h41fb33c4, 32'hc213743c} /* (28, 10, 23) {real, imag} */,
  {32'hc175994c, 32'h3f5b5680} /* (28, 10, 22) {real, imag} */,
  {32'hc15bc12e, 32'h40fcb0bc} /* (28, 10, 21) {real, imag} */,
  {32'h40187f38, 32'hc1de2e0a} /* (28, 10, 20) {real, imag} */,
  {32'h411353bc, 32'hc113b242} /* (28, 10, 19) {real, imag} */,
  {32'hc12ede21, 32'hc078a218} /* (28, 10, 18) {real, imag} */,
  {32'hbf822258, 32'h40fd5574} /* (28, 10, 17) {real, imag} */,
  {32'hc181c392, 32'h41a68d0e} /* (28, 10, 16) {real, imag} */,
  {32'hc10ea253, 32'hc16121fa} /* (28, 10, 15) {real, imag} */,
  {32'hc14196b7, 32'h4148a786} /* (28, 10, 14) {real, imag} */,
  {32'h4253918d, 32'hc1876a83} /* (28, 10, 13) {real, imag} */,
  {32'h41f4c5b1, 32'h410344c5} /* (28, 10, 12) {real, imag} */,
  {32'hc1b5a9b5, 32'hc1fab617} /* (28, 10, 11) {real, imag} */,
  {32'h4195a14a, 32'h40779420} /* (28, 10, 10) {real, imag} */,
  {32'h418dae5e, 32'hc2245d06} /* (28, 10, 9) {real, imag} */,
  {32'hbff10bc0, 32'h3d81ed00} /* (28, 10, 8) {real, imag} */,
  {32'h428c022b, 32'hc2561d96} /* (28, 10, 7) {real, imag} */,
  {32'h3f44a3e8, 32'h426cc109} /* (28, 10, 6) {real, imag} */,
  {32'hc23d1ad6, 32'h41dc7101} /* (28, 10, 5) {real, imag} */,
  {32'hc23d7614, 32'hc21a4f13} /* (28, 10, 4) {real, imag} */,
  {32'hc05000a0, 32'h4202cafc} /* (28, 10, 3) {real, imag} */,
  {32'hc27a8547, 32'h428b1f18} /* (28, 10, 2) {real, imag} */,
  {32'h418b3818, 32'hc2d55529} /* (28, 10, 1) {real, imag} */,
  {32'h42b30e7e, 32'h42dfaae8} /* (28, 10, 0) {real, imag} */,
  {32'h42226929, 32'hc26ab84a} /* (28, 9, 31) {real, imag} */,
  {32'hc3226a58, 32'hc1eef744} /* (28, 9, 30) {real, imag} */,
  {32'hc1fc65ce, 32'h42b374cf} /* (28, 9, 29) {real, imag} */,
  {32'h42c776d6, 32'hc2357a41} /* (28, 9, 28) {real, imag} */,
  {32'h4243ab66, 32'h42bdbd60} /* (28, 9, 27) {real, imag} */,
  {32'h42789e1f, 32'hc2a07470} /* (28, 9, 26) {real, imag} */,
  {32'hc223309f, 32'hc291d9b8} /* (28, 9, 25) {real, imag} */,
  {32'h412bf2c0, 32'hc1891008} /* (28, 9, 24) {real, imag} */,
  {32'hc1953d96, 32'hc0739440} /* (28, 9, 23) {real, imag} */,
  {32'h429f30f0, 32'h41907dfc} /* (28, 9, 22) {real, imag} */,
  {32'h41e9fbb3, 32'h4241b27d} /* (28, 9, 21) {real, imag} */,
  {32'h41268776, 32'hc20fdc26} /* (28, 9, 20) {real, imag} */,
  {32'hc12ef932, 32'hbfbbf9a0} /* (28, 9, 19) {real, imag} */,
  {32'hc03988b8, 32'h41a7b4ce} /* (28, 9, 18) {real, imag} */,
  {32'hc105dcba, 32'h41822020} /* (28, 9, 17) {real, imag} */,
  {32'h407542e8, 32'h416f97d0} /* (28, 9, 16) {real, imag} */,
  {32'hc11a236e, 32'hc0b943ba} /* (28, 9, 15) {real, imag} */,
  {32'hbf951ad0, 32'hc16ad95c} /* (28, 9, 14) {real, imag} */,
  {32'h41fe2813, 32'h3e96bc00} /* (28, 9, 13) {real, imag} */,
  {32'h41572cd2, 32'hc15ea8f6} /* (28, 9, 12) {real, imag} */,
  {32'hc2056647, 32'hc1a99456} /* (28, 9, 11) {real, imag} */,
  {32'hc1ffe78e, 32'h42156806} /* (28, 9, 10) {real, imag} */,
  {32'h3fb4f0e8, 32'hc22ab5d6} /* (28, 9, 9) {real, imag} */,
  {32'h424cb445, 32'hc01f5c7c} /* (28, 9, 8) {real, imag} */,
  {32'hc2248615, 32'hc1bc9d74} /* (28, 9, 7) {real, imag} */,
  {32'hc1a4d14a, 32'h41a7a880} /* (28, 9, 6) {real, imag} */,
  {32'hc289c221, 32'hc2c5b894} /* (28, 9, 5) {real, imag} */,
  {32'h429efbca, 32'hc2164b17} /* (28, 9, 4) {real, imag} */,
  {32'hc0f876b2, 32'h40a07070} /* (28, 9, 3) {real, imag} */,
  {32'hc23d0820, 32'h43017c20} /* (28, 9, 2) {real, imag} */,
  {32'h422695b5, 32'hc13bb026} /* (28, 9, 1) {real, imag} */,
  {32'h424592d8, 32'hc25c403c} /* (28, 9, 0) {real, imag} */,
  {32'hc29bd6d8, 32'h4383e95e} /* (28, 8, 31) {real, imag} */,
  {32'hc2c484fb, 32'hc344d7f0} /* (28, 8, 30) {real, imag} */,
  {32'h41e50378, 32'hc28ebdf2} /* (28, 8, 29) {real, imag} */,
  {32'hc0b2077e, 32'h4186f740} /* (28, 8, 28) {real, imag} */,
  {32'h4204296c, 32'hc0ec8f70} /* (28, 8, 27) {real, imag} */,
  {32'hc29f4e7a, 32'hc2c8aaf7} /* (28, 8, 26) {real, imag} */,
  {32'h41331794, 32'h41f4005e} /* (28, 8, 25) {real, imag} */,
  {32'hc2c3a590, 32'hc23c876e} /* (28, 8, 24) {real, imag} */,
  {32'h423faf7a, 32'h41aeda98} /* (28, 8, 23) {real, imag} */,
  {32'h41c15c7d, 32'hc2a9de3f} /* (28, 8, 22) {real, imag} */,
  {32'hc14af67c, 32'hc1c0482c} /* (28, 8, 21) {real, imag} */,
  {32'hc18978ea, 32'h42bf2922} /* (28, 8, 20) {real, imag} */,
  {32'hc18b76bd, 32'h3f9c78d0} /* (28, 8, 19) {real, imag} */,
  {32'hc184372a, 32'h413c4c38} /* (28, 8, 18) {real, imag} */,
  {32'h408f5d09, 32'hc140265a} /* (28, 8, 17) {real, imag} */,
  {32'h411d78c0, 32'h40668a60} /* (28, 8, 16) {real, imag} */,
  {32'h40de2a27, 32'hc1561e36} /* (28, 8, 15) {real, imag} */,
  {32'hc196f95e, 32'hc14dc088} /* (28, 8, 14) {real, imag} */,
  {32'hc106ebea, 32'hc13016ca} /* (28, 8, 13) {real, imag} */,
  {32'hc040799c, 32'h4244d5f4} /* (28, 8, 12) {real, imag} */,
  {32'h404ff190, 32'h4068a700} /* (28, 8, 11) {real, imag} */,
  {32'h41d9b6d9, 32'h41a1be3c} /* (28, 8, 10) {real, imag} */,
  {32'h420f86ce, 32'h41fdab14} /* (28, 8, 9) {real, imag} */,
  {32'h41c1a968, 32'hc2a96aad} /* (28, 8, 8) {real, imag} */,
  {32'h41f1b55c, 32'h428d67fa} /* (28, 8, 7) {real, imag} */,
  {32'h41e7528d, 32'hc238c7da} /* (28, 8, 6) {real, imag} */,
  {32'h422641c0, 32'h42cb73ae} /* (28, 8, 5) {real, imag} */,
  {32'hc19a78aa, 32'h42694a9e} /* (28, 8, 4) {real, imag} */,
  {32'hc2fb657a, 32'hc1823571} /* (28, 8, 3) {real, imag} */,
  {32'h42d50679, 32'hc26886ca} /* (28, 8, 2) {real, imag} */,
  {32'hc274d560, 32'h4360fa30} /* (28, 8, 1) {real, imag} */,
  {32'hc2cba094, 32'h436f9798} /* (28, 8, 0) {real, imag} */,
  {32'hc287ace6, 32'h42138cf1} /* (28, 7, 31) {real, imag} */,
  {32'h42d5bbc0, 32'hc1e5d76c} /* (28, 7, 30) {real, imag} */,
  {32'hc1c280e4, 32'hc1a5ce92} /* (28, 7, 29) {real, imag} */,
  {32'hc283e131, 32'h42fedf5c} /* (28, 7, 28) {real, imag} */,
  {32'hc26943b4, 32'hc16ec56c} /* (28, 7, 27) {real, imag} */,
  {32'h42a59a06, 32'h42490a1f} /* (28, 7, 26) {real, imag} */,
  {32'hc0c0cd3c, 32'hc1daccb4} /* (28, 7, 25) {real, imag} */,
  {32'h430ff3c0, 32'hc13b9f02} /* (28, 7, 24) {real, imag} */,
  {32'hc1be918c, 32'hc22ef9ee} /* (28, 7, 23) {real, imag} */,
  {32'h3fa8fbb8, 32'h41ad29c4} /* (28, 7, 22) {real, imag} */,
  {32'hc1fee72c, 32'hc1360cbc} /* (28, 7, 21) {real, imag} */,
  {32'hc271a2bb, 32'h418be916} /* (28, 7, 20) {real, imag} */,
  {32'h4145b2ff, 32'hc207670f} /* (28, 7, 19) {real, imag} */,
  {32'hc19fce6f, 32'hc1ea2b3c} /* (28, 7, 18) {real, imag} */,
  {32'h4169dd21, 32'hc1e575d0} /* (28, 7, 17) {real, imag} */,
  {32'hc1cf3363, 32'hc1a1f68e} /* (28, 7, 16) {real, imag} */,
  {32'hc169ee65, 32'h40ab893e} /* (28, 7, 15) {real, imag} */,
  {32'h41fbb96d, 32'h419ad70c} /* (28, 7, 14) {real, imag} */,
  {32'h421c7a89, 32'hc0440310} /* (28, 7, 13) {real, imag} */,
  {32'hc1c0ab52, 32'h416d6fc3} /* (28, 7, 12) {real, imag} */,
  {32'h426cf6a8, 32'h41a76526} /* (28, 7, 11) {real, imag} */,
  {32'h41aa5edc, 32'hc19ec5ce} /* (28, 7, 10) {real, imag} */,
  {32'hc2523aa0, 32'h423fe946} /* (28, 7, 9) {real, imag} */,
  {32'hc1009df8, 32'h420270ce} /* (28, 7, 8) {real, imag} */,
  {32'hc1b3fbf0, 32'hc28d2a4b} /* (28, 7, 7) {real, imag} */,
  {32'hc2269843, 32'hc14c2780} /* (28, 7, 6) {real, imag} */,
  {32'hc13a5468, 32'hc2e10de4} /* (28, 7, 5) {real, imag} */,
  {32'h42ff0b43, 32'h42850522} /* (28, 7, 4) {real, imag} */,
  {32'hc20d1d39, 32'h42adcdc0} /* (28, 7, 3) {real, imag} */,
  {32'hc323431a, 32'hc3541684} /* (28, 7, 2) {real, imag} */,
  {32'hc228ecfb, 32'h4117ffab} /* (28, 7, 1) {real, imag} */,
  {32'h41d42437, 32'hc1a7e1b6} /* (28, 7, 0) {real, imag} */,
  {32'h4303049c, 32'h418e8568} /* (28, 6, 31) {real, imag} */,
  {32'hc32f2c4a, 32'hc20caf86} /* (28, 6, 30) {real, imag} */,
  {32'hc2a64d34, 32'hc211e968} /* (28, 6, 29) {real, imag} */,
  {32'h422e3535, 32'h43087a24} /* (28, 6, 28) {real, imag} */,
  {32'h431805b6, 32'h419c79b8} /* (28, 6, 27) {real, imag} */,
  {32'hc288be23, 32'h43301496} /* (28, 6, 26) {real, imag} */,
  {32'h42398278, 32'h4206b4e1} /* (28, 6, 25) {real, imag} */,
  {32'h4153c086, 32'hc2fe3c62} /* (28, 6, 24) {real, imag} */,
  {32'hc2098e74, 32'h41a1a230} /* (28, 6, 23) {real, imag} */,
  {32'hc24fade6, 32'h41ecd0db} /* (28, 6, 22) {real, imag} */,
  {32'h409c4360, 32'h42a1b896} /* (28, 6, 21) {real, imag} */,
  {32'h3fc68b68, 32'h41da01b8} /* (28, 6, 20) {real, imag} */,
  {32'hc1b83df6, 32'h41582e02} /* (28, 6, 19) {real, imag} */,
  {32'h41483250, 32'hc21092be} /* (28, 6, 18) {real, imag} */,
  {32'hc1c1ea18, 32'h41e6fb50} /* (28, 6, 17) {real, imag} */,
  {32'h40235d40, 32'h4146ef24} /* (28, 6, 16) {real, imag} */,
  {32'h41987420, 32'h41000410} /* (28, 6, 15) {real, imag} */,
  {32'h420c9b02, 32'h4200760a} /* (28, 6, 14) {real, imag} */,
  {32'hc1b11aae, 32'hc2499172} /* (28, 6, 13) {real, imag} */,
  {32'hbeb190a0, 32'hbf843080} /* (28, 6, 12) {real, imag} */,
  {32'h4244950e, 32'h3f975880} /* (28, 6, 11) {real, imag} */,
  {32'hc1159660, 32'h41c88e45} /* (28, 6, 10) {real, imag} */,
  {32'h42d1f914, 32'hbe94fc80} /* (28, 6, 9) {real, imag} */,
  {32'h421334bc, 32'hc2093238} /* (28, 6, 8) {real, imag} */,
  {32'hbfc5d470, 32'h41ddead0} /* (28, 6, 7) {real, imag} */,
  {32'h41ee4528, 32'h43143e2e} /* (28, 6, 6) {real, imag} */,
  {32'h4269c1df, 32'h4296d57e} /* (28, 6, 5) {real, imag} */,
  {32'h42c3a942, 32'hc1a1b694} /* (28, 6, 4) {real, imag} */,
  {32'hc19b614a, 32'h4266197e} /* (28, 6, 3) {real, imag} */,
  {32'h4253c317, 32'hc156a488} /* (28, 6, 2) {real, imag} */,
  {32'h42a0e1c2, 32'h431f9cfa} /* (28, 6, 1) {real, imag} */,
  {32'hc2c4f972, 32'hc2bb9902} /* (28, 6, 0) {real, imag} */,
  {32'h43ce41d8, 32'h43b4d8cc} /* (28, 5, 31) {real, imag} */,
  {32'hc259c804, 32'hc336cf6a} /* (28, 5, 30) {real, imag} */,
  {32'h405af558, 32'h4294c7c9} /* (28, 5, 29) {real, imag} */,
  {32'hc228ae92, 32'hc22bbf90} /* (28, 5, 28) {real, imag} */,
  {32'hc265fc1e, 32'hc2b95de6} /* (28, 5, 27) {real, imag} */,
  {32'h4206a2c7, 32'h42f1ec7e} /* (28, 5, 26) {real, imag} */,
  {32'hc2e753bb, 32'h42653f26} /* (28, 5, 25) {real, imag} */,
  {32'h427cb314, 32'h424b9c3f} /* (28, 5, 24) {real, imag} */,
  {32'hc1f83f24, 32'hc2405159} /* (28, 5, 23) {real, imag} */,
  {32'hbfd5ceb0, 32'hc0b31bf8} /* (28, 5, 22) {real, imag} */,
  {32'hc21a4f88, 32'hc2a0e766} /* (28, 5, 21) {real, imag} */,
  {32'hc0d44234, 32'hc13d89af} /* (28, 5, 20) {real, imag} */,
  {32'h4219822d, 32'hc1957af9} /* (28, 5, 19) {real, imag} */,
  {32'hc196a0d9, 32'hc185c7f2} /* (28, 5, 18) {real, imag} */,
  {32'hc22410c4, 32'hc082d3a4} /* (28, 5, 17) {real, imag} */,
  {32'h401a9888, 32'h41990478} /* (28, 5, 16) {real, imag} */,
  {32'h41026610, 32'h40178f48} /* (28, 5, 15) {real, imag} */,
  {32'h403a6e38, 32'h41448595} /* (28, 5, 14) {real, imag} */,
  {32'hc22f3ad7, 32'h41f19f73} /* (28, 5, 13) {real, imag} */,
  {32'hc1eb5237, 32'h422c107c} /* (28, 5, 12) {real, imag} */,
  {32'hc1b57205, 32'h420c2c37} /* (28, 5, 11) {real, imag} */,
  {32'h3fcc9790, 32'hc20a9feb} /* (28, 5, 10) {real, imag} */,
  {32'hc2035136, 32'h41995a1a} /* (28, 5, 9) {real, imag} */,
  {32'h41d00de0, 32'h4126fd2c} /* (28, 5, 8) {real, imag} */,
  {32'hc2cf902d, 32'h4181ab5c} /* (28, 5, 7) {real, imag} */,
  {32'h425a23f5, 32'hc2e6e3d4} /* (28, 5, 6) {real, imag} */,
  {32'h42ceb339, 32'h420cdd4b} /* (28, 5, 5) {real, imag} */,
  {32'hc25ef40c, 32'h42df9942} /* (28, 5, 4) {real, imag} */,
  {32'hc1af0b55, 32'hc2e93b77} /* (28, 5, 3) {real, imag} */,
  {32'h43178ee4, 32'hc333ba46} /* (28, 5, 2) {real, imag} */,
  {32'hc3273919, 32'h43d50744} /* (28, 5, 1) {real, imag} */,
  {32'hc24073f8, 32'h438dfd5c} /* (28, 5, 0) {real, imag} */,
  {32'h42b24026, 32'hc361d018} /* (28, 4, 31) {real, imag} */,
  {32'hc29ab660, 32'h43162c14} /* (28, 4, 30) {real, imag} */,
  {32'h428ee2ef, 32'hc3229676} /* (28, 4, 29) {real, imag} */,
  {32'h4292d2dd, 32'hc3865b51} /* (28, 4, 28) {real, imag} */,
  {32'h40b58230, 32'h4338bc7c} /* (28, 4, 27) {real, imag} */,
  {32'h422993dc, 32'hc20f6df9} /* (28, 4, 26) {real, imag} */,
  {32'hc18ae93d, 32'h428066c6} /* (28, 4, 25) {real, imag} */,
  {32'h42ba5a9b, 32'hc0f38fb0} /* (28, 4, 24) {real, imag} */,
  {32'hc181d12b, 32'h41ac50c2} /* (28, 4, 23) {real, imag} */,
  {32'hc1d99a7e, 32'h40d74e88} /* (28, 4, 22) {real, imag} */,
  {32'hc206815f, 32'h42a5fba8} /* (28, 4, 21) {real, imag} */,
  {32'h3effea40, 32'h401ff480} /* (28, 4, 20) {real, imag} */,
  {32'hc1fdd090, 32'h4176d4fc} /* (28, 4, 19) {real, imag} */,
  {32'h42b5fc4c, 32'hc25f6674} /* (28, 4, 18) {real, imag} */,
  {32'h40647a38, 32'hc24c7a16} /* (28, 4, 17) {real, imag} */,
  {32'h411b8058, 32'h4148aeb0} /* (28, 4, 16) {real, imag} */,
  {32'h41fdb649, 32'hc05ccaa0} /* (28, 4, 15) {real, imag} */,
  {32'hc1c3b16e, 32'h4092e704} /* (28, 4, 14) {real, imag} */,
  {32'hc27a9974, 32'h42197b39} /* (28, 4, 13) {real, imag} */,
  {32'h420c7af0, 32'hc0e99160} /* (28, 4, 12) {real, imag} */,
  {32'h4229afe5, 32'hc190aaf2} /* (28, 4, 11) {real, imag} */,
  {32'h4314f5f8, 32'h41bd9372} /* (28, 4, 10) {real, imag} */,
  {32'hc0686298, 32'hbf301250} /* (28, 4, 9) {real, imag} */,
  {32'hc12d8028, 32'h4208c266} /* (28, 4, 8) {real, imag} */,
  {32'h4226ae7e, 32'hc202837b} /* (28, 4, 7) {real, imag} */,
  {32'hc21b4e12, 32'hc1680ec4} /* (28, 4, 6) {real, imag} */,
  {32'hc352178a, 32'h41ddfa60} /* (28, 4, 5) {real, imag} */,
  {32'hbf309880, 32'hc1c50254} /* (28, 4, 4) {real, imag} */,
  {32'hc2881e6d, 32'h426de8d8} /* (28, 4, 3) {real, imag} */,
  {32'hc39cdeb8, 32'h43a45102} /* (28, 4, 2) {real, imag} */,
  {32'h42c9ca8e, 32'hc3dc9988} /* (28, 4, 1) {real, imag} */,
  {32'h42c6aa05, 32'hc39b0ace} /* (28, 4, 0) {real, imag} */,
  {32'h43e1f68e, 32'h433763de} /* (28, 3, 31) {real, imag} */,
  {32'hc39ba0b6, 32'h40dba610} /* (28, 3, 30) {real, imag} */,
  {32'h431b7be8, 32'hc02b47a0} /* (28, 3, 29) {real, imag} */,
  {32'hbfe73540, 32'hc2819b4e} /* (28, 3, 28) {real, imag} */,
  {32'h429db742, 32'h424c48df} /* (28, 3, 27) {real, imag} */,
  {32'hc2d664c7, 32'h42a5ac4e} /* (28, 3, 26) {real, imag} */,
  {32'hc2f56f56, 32'hc2687492} /* (28, 3, 25) {real, imag} */,
  {32'hc325f113, 32'h42c0a2eb} /* (28, 3, 24) {real, imag} */,
  {32'hc2b16f2b, 32'h413b5068} /* (28, 3, 23) {real, imag} */,
  {32'h40ef2e90, 32'hc115f158} /* (28, 3, 22) {real, imag} */,
  {32'h4219ca86, 32'h40a611e2} /* (28, 3, 21) {real, imag} */,
  {32'hc198d6ca, 32'hbffda130} /* (28, 3, 20) {real, imag} */,
  {32'h423a48d8, 32'hc1be3026} /* (28, 3, 19) {real, imag} */,
  {32'h4125d8ba, 32'h41af0b98} /* (28, 3, 18) {real, imag} */,
  {32'h4281d867, 32'h40af5030} /* (28, 3, 17) {real, imag} */,
  {32'hc1b62730, 32'h40f2518e} /* (28, 3, 16) {real, imag} */,
  {32'h408d0090, 32'h41bfdd4c} /* (28, 3, 15) {real, imag} */,
  {32'h4061fe98, 32'hc19c6e38} /* (28, 3, 14) {real, imag} */,
  {32'hc0972e20, 32'hc1d21fe2} /* (28, 3, 13) {real, imag} */,
  {32'h40768790, 32'h41aecaf5} /* (28, 3, 12) {real, imag} */,
  {32'h4269e49a, 32'hc096f9de} /* (28, 3, 11) {real, imag} */,
  {32'hc23dceee, 32'h429ca1fb} /* (28, 3, 10) {real, imag} */,
  {32'h40d78100, 32'h42a93f6b} /* (28, 3, 9) {real, imag} */,
  {32'h414b1530, 32'hc2c74cf9} /* (28, 3, 8) {real, imag} */,
  {32'hc33cf209, 32'hc24f2ef6} /* (28, 3, 7) {real, imag} */,
  {32'hc2b7b41b, 32'h42a7ffb8} /* (28, 3, 6) {real, imag} */,
  {32'hc2961198, 32'hc2dd3458} /* (28, 3, 5) {real, imag} */,
  {32'hc31b6fa6, 32'h42c95cf0} /* (28, 3, 4) {real, imag} */,
  {32'h429929c6, 32'hc3586d70} /* (28, 3, 3) {real, imag} */,
  {32'hc3446ffa, 32'h435276ca} /* (28, 3, 2) {real, imag} */,
  {32'h4332816c, 32'hc3ff804d} /* (28, 3, 1) {real, imag} */,
  {32'h433b49b4, 32'hc1de5d40} /* (28, 3, 0) {real, imag} */,
  {32'h4373e313, 32'h448d7812} /* (28, 2, 31) {real, imag} */,
  {32'hc3c13411, 32'hc43a9ae3} /* (28, 2, 30) {real, imag} */,
  {32'h4288ccbc, 32'h42d5c679} /* (28, 2, 29) {real, imag} */,
  {32'h4385d968, 32'h432ceafa} /* (28, 2, 28) {real, imag} */,
  {32'hc210219a, 32'h424e84f8} /* (28, 2, 27) {real, imag} */,
  {32'h405f9280, 32'hc0d557e8} /* (28, 2, 26) {real, imag} */,
  {32'hc1b4b366, 32'h42a3aaba} /* (28, 2, 25) {real, imag} */,
  {32'hc2eb876c, 32'hc30021a8} /* (28, 2, 24) {real, imag} */,
  {32'h427af963, 32'h42c90d8e} /* (28, 2, 23) {real, imag} */,
  {32'h42b69c78, 32'hc2682cad} /* (28, 2, 22) {real, imag} */,
  {32'hc2a064e4, 32'hc24b3df4} /* (28, 2, 21) {real, imag} */,
  {32'h41eac62c, 32'hc1f772ef} /* (28, 2, 20) {real, imag} */,
  {32'h4222a99f, 32'hbf12a920} /* (28, 2, 19) {real, imag} */,
  {32'hc28388b0, 32'h422625f4} /* (28, 2, 18) {real, imag} */,
  {32'h40f4ed98, 32'hc10e1a88} /* (28, 2, 17) {real, imag} */,
  {32'hc2517374, 32'h423f56f0} /* (28, 2, 16) {real, imag} */,
  {32'h4211dfe5, 32'h41ec6444} /* (28, 2, 15) {real, imag} */,
  {32'h40407f80, 32'hc251f7d4} /* (28, 2, 14) {real, imag} */,
  {32'h41b2888e, 32'h41373fbe} /* (28, 2, 13) {real, imag} */,
  {32'hc2003ec2, 32'hbf616320} /* (28, 2, 12) {real, imag} */,
  {32'h42636bff, 32'hc2f16a3e} /* (28, 2, 11) {real, imag} */,
  {32'h41b104c2, 32'hc2145f23} /* (28, 2, 10) {real, imag} */,
  {32'h42551531, 32'hc1dfb258} /* (28, 2, 9) {real, imag} */,
  {32'hc0ac7a00, 32'hc2ca5304} /* (28, 2, 8) {real, imag} */,
  {32'hc2ad75f8, 32'h42a3fab6} /* (28, 2, 7) {real, imag} */,
  {32'h430475c6, 32'h42144bbd} /* (28, 2, 6) {real, imag} */,
  {32'hc0e3bce0, 32'hc3a3ca80} /* (28, 2, 5) {real, imag} */,
  {32'h43740485, 32'h439364a7} /* (28, 2, 4) {real, imag} */,
  {32'hc2082f83, 32'hc2660626} /* (28, 2, 3) {real, imag} */,
  {32'hc32b445e, 32'hc3afc3ae} /* (28, 2, 2) {real, imag} */,
  {32'h43432aff, 32'h441c75af} /* (28, 2, 1) {real, imag} */,
  {32'h42a873ca, 32'h441b8361} /* (28, 2, 0) {real, imag} */,
  {32'hc3cb1df0, 32'hc4782d1c} /* (28, 1, 31) {real, imag} */,
  {32'h41784f50, 32'h43d81cb3} /* (28, 1, 30) {real, imag} */,
  {32'h428514ef, 32'hc22b73c3} /* (28, 1, 29) {real, imag} */,
  {32'hc29ba728, 32'hc2dcff02} /* (28, 1, 28) {real, imag} */,
  {32'h439330a4, 32'h43a0450b} /* (28, 1, 27) {real, imag} */,
  {32'hc08c6aa8, 32'h42c3cefc} /* (28, 1, 26) {real, imag} */,
  {32'hc245e962, 32'h42446086} /* (28, 1, 25) {real, imag} */,
  {32'h42e04cd0, 32'h4290370e} /* (28, 1, 24) {real, imag} */,
  {32'h421267e4, 32'h424f4ba2} /* (28, 1, 23) {real, imag} */,
  {32'hc2daf00a, 32'hc2ea97f7} /* (28, 1, 22) {real, imag} */,
  {32'h432b5207, 32'hc1c9ac80} /* (28, 1, 21) {real, imag} */,
  {32'hc17c5010, 32'hc2322201} /* (28, 1, 20) {real, imag} */,
  {32'h41d9c5a2, 32'h422971b0} /* (28, 1, 19) {real, imag} */,
  {32'h3e926600, 32'h42bc7b95} /* (28, 1, 18) {real, imag} */,
  {32'hc20d08ec, 32'hbfc07500} /* (28, 1, 17) {real, imag} */,
  {32'hc22d8e4c, 32'h4147e880} /* (28, 1, 16) {real, imag} */,
  {32'hc140d650, 32'h4190ca90} /* (28, 1, 15) {real, imag} */,
  {32'hc291813e, 32'hc192f1f4} /* (28, 1, 14) {real, imag} */,
  {32'h40ddcc28, 32'hc0963270} /* (28, 1, 13) {real, imag} */,
  {32'hc01f3560, 32'hc292c754} /* (28, 1, 12) {real, imag} */,
  {32'hc2986a52, 32'h41c60220} /* (28, 1, 11) {real, imag} */,
  {32'hc1a3b448, 32'hc10f9e08} /* (28, 1, 10) {real, imag} */,
  {32'h42776204, 32'hc2e8d155} /* (28, 1, 9) {real, imag} */,
  {32'hc31ba9a4, 32'h42ed08fa} /* (28, 1, 8) {real, imag} */,
  {32'h42f6ba1f, 32'hc29f12ff} /* (28, 1, 7) {real, imag} */,
  {32'h4211754b, 32'h42f5da0c} /* (28, 1, 6) {real, imag} */,
  {32'h4113f2c0, 32'h4357d8f6} /* (28, 1, 5) {real, imag} */,
  {32'h42edb640, 32'hc32257ff} /* (28, 1, 4) {real, imag} */,
  {32'h4281b961, 32'h43062f9d} /* (28, 1, 3) {real, imag} */,
  {32'hc3b38e34, 32'h444d263e} /* (28, 1, 2) {real, imag} */,
  {32'h42bcfbde, 32'hc4bb28fa} /* (28, 1, 1) {real, imag} */,
  {32'hc39c767e, 32'hc43b3ea5} /* (28, 1, 0) {real, imag} */,
  {32'hc42bf624, 32'hc3ccd967} /* (28, 0, 31) {real, imag} */,
  {32'h437725c6, 32'hc1c318cb} /* (28, 0, 30) {real, imag} */,
  {32'h429d0aa4, 32'h4322791b} /* (28, 0, 29) {real, imag} */,
  {32'h42754747, 32'hc2b13347} /* (28, 0, 28) {real, imag} */,
  {32'h41329750, 32'h43187eb1} /* (28, 0, 27) {real, imag} */,
  {32'hc222c951, 32'h429fb892} /* (28, 0, 26) {real, imag} */,
  {32'hc30e61f0, 32'h423353b6} /* (28, 0, 25) {real, imag} */,
  {32'h42ea2170, 32'h417f0be0} /* (28, 0, 24) {real, imag} */,
  {32'h430b83f2, 32'hc299802f} /* (28, 0, 23) {real, imag} */,
  {32'hbccb5000, 32'h42cc627c} /* (28, 0, 22) {real, imag} */,
  {32'h42770dd3, 32'h420fc4d3} /* (28, 0, 21) {real, imag} */,
  {32'hc08333dc, 32'h41316e76} /* (28, 0, 20) {real, imag} */,
  {32'hc0f1b178, 32'h428c06a6} /* (28, 0, 19) {real, imag} */,
  {32'h421b0ebc, 32'h4127d330} /* (28, 0, 18) {real, imag} */,
  {32'h41aa29bc, 32'h4137d618} /* (28, 0, 17) {real, imag} */,
  {32'h420191b2, 32'h414d3fd0} /* (28, 0, 16) {real, imag} */,
  {32'hc21c7caa, 32'hc183608c} /* (28, 0, 15) {real, imag} */,
  {32'hc2c221a6, 32'h41d5fd12} /* (28, 0, 14) {real, imag} */,
  {32'hc0e360a8, 32'hc091b990} /* (28, 0, 13) {real, imag} */,
  {32'h41a397ed, 32'h4096216b} /* (28, 0, 12) {real, imag} */,
  {32'h4155b9cc, 32'h42f4933e} /* (28, 0, 11) {real, imag} */,
  {32'h42a47e98, 32'h41c650e6} /* (28, 0, 10) {real, imag} */,
  {32'hc300b2a8, 32'h43253aa0} /* (28, 0, 9) {real, imag} */,
  {32'hc247e0dc, 32'h42a2d840} /* (28, 0, 8) {real, imag} */,
  {32'h430e97b6, 32'hc2ab2bc3} /* (28, 0, 7) {real, imag} */,
  {32'h42ab15ba, 32'hbf8befe0} /* (28, 0, 6) {real, imag} */,
  {32'h4326fd99, 32'h433667ff} /* (28, 0, 5) {real, imag} */,
  {32'hc274b3bf, 32'h42cde885} /* (28, 0, 4) {real, imag} */,
  {32'h41984c66, 32'hc2bcfcfa} /* (28, 0, 3) {real, imag} */,
  {32'hc364ea90, 32'h4236a84a} /* (28, 0, 2) {real, imag} */,
  {32'h436f90fe, 32'hc440bafc} /* (28, 0, 1) {real, imag} */,
  {32'hc38faec1, 32'hc3fc1558} /* (28, 0, 0) {real, imag} */,
  {32'h440461d6, 32'h434e64b6} /* (27, 31, 31) {real, imag} */,
  {32'hc3e6bf56, 32'hc356dabe} /* (27, 31, 30) {real, imag} */,
  {32'hc1e8e8c1, 32'h4286a82e} /* (27, 31, 29) {real, imag} */,
  {32'h425a5e39, 32'h42c803c2} /* (27, 31, 28) {real, imag} */,
  {32'hc2ae8ca8, 32'hbec75300} /* (27, 31, 27) {real, imag} */,
  {32'h4257f1a2, 32'h41a6c558} /* (27, 31, 26) {real, imag} */,
  {32'h41acc7a2, 32'hc2a2aba2} /* (27, 31, 25) {real, imag} */,
  {32'hc2806f9f, 32'h4236711a} /* (27, 31, 24) {real, imag} */,
  {32'hc2aea70e, 32'h41c6fc7e} /* (27, 31, 23) {real, imag} */,
  {32'h4259ef1e, 32'hc14e307c} /* (27, 31, 22) {real, imag} */,
  {32'hc29d621e, 32'h41aa5e41} /* (27, 31, 21) {real, imag} */,
  {32'h4048e3f0, 32'hc272b7bc} /* (27, 31, 20) {real, imag} */,
  {32'hc0ff7524, 32'hbf0a7610} /* (27, 31, 19) {real, imag} */,
  {32'hc173c038, 32'h41bbb46c} /* (27, 31, 18) {real, imag} */,
  {32'hbffa4f00, 32'h417778bc} /* (27, 31, 17) {real, imag} */,
  {32'hc1c75d9c, 32'h4018c680} /* (27, 31, 16) {real, imag} */,
  {32'hc23af630, 32'hc1763e7c} /* (27, 31, 15) {real, imag} */,
  {32'h42d6c6d5, 32'h41d2adc4} /* (27, 31, 14) {real, imag} */,
  {32'hc122cc32, 32'h4094a6ee} /* (27, 31, 13) {real, imag} */,
  {32'hc20ea159, 32'h415769b8} /* (27, 31, 12) {real, imag} */,
  {32'h420d1c6b, 32'hc23de90c} /* (27, 31, 11) {real, imag} */,
  {32'h42595bd2, 32'hc2133520} /* (27, 31, 10) {real, imag} */,
  {32'h41bd035e, 32'h4226eed5} /* (27, 31, 9) {real, imag} */,
  {32'hc23ad242, 32'hc29dedbd} /* (27, 31, 8) {real, imag} */,
  {32'hc23a5f53, 32'h4155821c} /* (27, 31, 7) {real, imag} */,
  {32'hc22861da, 32'h41a8f57a} /* (27, 31, 6) {real, imag} */,
  {32'hc31c8194, 32'hc2f1c7d9} /* (27, 31, 5) {real, imag} */,
  {32'h430bc1e0, 32'hc1a06704} /* (27, 31, 4) {real, imag} */,
  {32'h4224ff22, 32'hc2a3cef2} /* (27, 31, 3) {real, imag} */,
  {32'hc27eaecc, 32'hc240c3fe} /* (27, 31, 2) {real, imag} */,
  {32'h4320da77, 32'h43c1e99f} /* (27, 31, 1) {real, imag} */,
  {32'h4353ff34, 32'h43a57171} /* (27, 31, 0) {real, imag} */,
  {32'hc2adf6df, 32'hc35bd8db} /* (27, 30, 31) {real, imag} */,
  {32'h4281d011, 32'h43c8341a} /* (27, 30, 30) {real, imag} */,
  {32'hc2215075, 32'hc3355913} /* (27, 30, 29) {real, imag} */,
  {32'hc345f579, 32'hc22f003d} /* (27, 30, 28) {real, imag} */,
  {32'h434c4078, 32'h41bb9c20} /* (27, 30, 27) {real, imag} */,
  {32'hc27d70ea, 32'hc2a056c4} /* (27, 30, 26) {real, imag} */,
  {32'h40681a30, 32'hc2df5dc2} /* (27, 30, 25) {real, imag} */,
  {32'h42866316, 32'h42945528} /* (27, 30, 24) {real, imag} */,
  {32'hc2638def, 32'h42102053} /* (27, 30, 23) {real, imag} */,
  {32'h4108ea48, 32'h422afe2c} /* (27, 30, 22) {real, imag} */,
  {32'h420d6422, 32'h4218da4c} /* (27, 30, 21) {real, imag} */,
  {32'hc166d6f2, 32'hc11e1588} /* (27, 30, 20) {real, imag} */,
  {32'hc05c442c, 32'h3f70af20} /* (27, 30, 19) {real, imag} */,
  {32'h4155fdde, 32'h4114db38} /* (27, 30, 18) {real, imag} */,
  {32'h40413420, 32'hbea6be00} /* (27, 30, 17) {real, imag} */,
  {32'hc1faa73a, 32'hc223a7bc} /* (27, 30, 16) {real, imag} */,
  {32'h4288a1a9, 32'h4172b570} /* (27, 30, 15) {real, imag} */,
  {32'hc1eedeef, 32'h40cbe550} /* (27, 30, 14) {real, imag} */,
  {32'h407d83cc, 32'hc1e0be71} /* (27, 30, 13) {real, imag} */,
  {32'hc1da6339, 32'h428d242c} /* (27, 30, 12) {real, imag} */,
  {32'h41e4a494, 32'hc0539c60} /* (27, 30, 11) {real, imag} */,
  {32'hc228baca, 32'h42391302} /* (27, 30, 10) {real, imag} */,
  {32'h41f2d7ee, 32'h427ec599} /* (27, 30, 9) {real, imag} */,
  {32'h409ffdec, 32'hc2e022f4} /* (27, 30, 8) {real, imag} */,
  {32'hc26976c3, 32'hc26063f1} /* (27, 30, 7) {real, imag} */,
  {32'h4195e634, 32'h42c454b4} /* (27, 30, 6) {real, imag} */,
  {32'h42c14481, 32'h43548160} /* (27, 30, 5) {real, imag} */,
  {32'h43371c57, 32'hc3139417} /* (27, 30, 4) {real, imag} */,
  {32'hc27abbe1, 32'hc2e5bf2a} /* (27, 30, 3) {real, imag} */,
  {32'h42bcf0f3, 32'h4401952d} /* (27, 30, 2) {real, imag} */,
  {32'hc357ae3c, 32'hc4143def} /* (27, 30, 1) {real, imag} */,
  {32'hc21ddad9, 32'hc1f015d5} /* (27, 30, 0) {real, imag} */,
  {32'h43d1102e, 32'h41b7530c} /* (27, 29, 31) {real, imag} */,
  {32'hc304c7a4, 32'hc29be739} /* (27, 29, 30) {real, imag} */,
  {32'h42fefb3e, 32'h4114f4e0} /* (27, 29, 29) {real, imag} */,
  {32'h404cb7f8, 32'hc2fb19e0} /* (27, 29, 28) {real, imag} */,
  {32'h43227f8a, 32'h4281f623} /* (27, 29, 27) {real, imag} */,
  {32'h409ad4d0, 32'hc2cb195c} /* (27, 29, 26) {real, imag} */,
  {32'hc1726298, 32'hc0322440} /* (27, 29, 25) {real, imag} */,
  {32'h4285b44c, 32'h41bc930e} /* (27, 29, 24) {real, imag} */,
  {32'h40e5be54, 32'h41009c88} /* (27, 29, 23) {real, imag} */,
  {32'h424f3390, 32'h416cb5dc} /* (27, 29, 22) {real, imag} */,
  {32'h41aaaa2c, 32'h41bedcf6} /* (27, 29, 21) {real, imag} */,
  {32'h420f51fa, 32'h42a748da} /* (27, 29, 20) {real, imag} */,
  {32'h41b566f8, 32'hc128627e} /* (27, 29, 19) {real, imag} */,
  {32'h425f345a, 32'hc0658ebe} /* (27, 29, 18) {real, imag} */,
  {32'hc2059fac, 32'hc171782a} /* (27, 29, 17) {real, imag} */,
  {32'hc1d1ab22, 32'hc219d1ff} /* (27, 29, 16) {real, imag} */,
  {32'hc028abc0, 32'hc1f64437} /* (27, 29, 15) {real, imag} */,
  {32'hc247b03e, 32'hbd9b7bc0} /* (27, 29, 14) {real, imag} */,
  {32'h41e27920, 32'h41f7ac51} /* (27, 29, 13) {real, imag} */,
  {32'hc07b9674, 32'h422ba3ad} /* (27, 29, 12) {real, imag} */,
  {32'h41dbcf98, 32'h40d97908} /* (27, 29, 11) {real, imag} */,
  {32'h4201ac9c, 32'h42437d77} /* (27, 29, 10) {real, imag} */,
  {32'h42785a66, 32'hc27e6784} /* (27, 29, 9) {real, imag} */,
  {32'hc2301685, 32'hc26cb333} /* (27, 29, 8) {real, imag} */,
  {32'h3f1ced40, 32'hc2cb1523} /* (27, 29, 7) {real, imag} */,
  {32'hc2929f59, 32'h42997b10} /* (27, 29, 6) {real, imag} */,
  {32'hc1702660, 32'hc2e97d99} /* (27, 29, 5) {real, imag} */,
  {32'h422b9366, 32'h419112ca} /* (27, 29, 4) {real, imag} */,
  {32'h41af2f88, 32'hc2dafb24} /* (27, 29, 3) {real, imag} */,
  {32'hc29b11af, 32'h42987b23} /* (27, 29, 2) {real, imag} */,
  {32'hc33eb8cf, 32'hc1ac4df6} /* (27, 29, 1) {real, imag} */,
  {32'hc2f20340, 32'hc2837f8a} /* (27, 29, 0) {real, imag} */,
  {32'h43157c1a, 32'h424ff6f9} /* (27, 28, 31) {real, imag} */,
  {32'hc354d6e3, 32'hc256a8b4} /* (27, 28, 30) {real, imag} */,
  {32'h3ecc61c0, 32'hc22af086} /* (27, 28, 29) {real, imag} */,
  {32'hc258118d, 32'hc22398f0} /* (27, 28, 28) {real, imag} */,
  {32'hc1cb7f50, 32'hc1b1c9fe} /* (27, 28, 27) {real, imag} */,
  {32'hc30726f0, 32'hc11995b0} /* (27, 28, 26) {real, imag} */,
  {32'h41ba3dfb, 32'h41d6a434} /* (27, 28, 25) {real, imag} */,
  {32'hc2191f35, 32'hc06276c0} /* (27, 28, 24) {real, imag} */,
  {32'hc23f09b6, 32'h4286df63} /* (27, 28, 23) {real, imag} */,
  {32'hc166d420, 32'h41bee1f9} /* (27, 28, 22) {real, imag} */,
  {32'h420c114c, 32'hc207003e} /* (27, 28, 21) {real, imag} */,
  {32'h4131b618, 32'hc1f64dae} /* (27, 28, 20) {real, imag} */,
  {32'h4261365c, 32'h415cbfc8} /* (27, 28, 19) {real, imag} */,
  {32'hc2502c74, 32'hc1c21798} /* (27, 28, 18) {real, imag} */,
  {32'hc0fad9f8, 32'h418f55ea} /* (27, 28, 17) {real, imag} */,
  {32'h406077c0, 32'h4183918a} /* (27, 28, 16) {real, imag} */,
  {32'hc0fec0d8, 32'hc208da43} /* (27, 28, 15) {real, imag} */,
  {32'hc0e505e0, 32'hc0f8ab80} /* (27, 28, 14) {real, imag} */,
  {32'h40083ec8, 32'hc21d539c} /* (27, 28, 13) {real, imag} */,
  {32'hc10a5d80, 32'hc1ae9722} /* (27, 28, 12) {real, imag} */,
  {32'hc15def12, 32'hc237db26} /* (27, 28, 11) {real, imag} */,
  {32'h40c74940, 32'h41eff6f9} /* (27, 28, 10) {real, imag} */,
  {32'hc21a3bbe, 32'hc1efd857} /* (27, 28, 9) {real, imag} */,
  {32'hc2497ae5, 32'hc25b17e4} /* (27, 28, 8) {real, imag} */,
  {32'h4288b46d, 32'hc30cc50e} /* (27, 28, 7) {real, imag} */,
  {32'h418aa15c, 32'h433592c5} /* (27, 28, 6) {real, imag} */,
  {32'h42da8550, 32'h423950e1} /* (27, 28, 5) {real, imag} */,
  {32'h4302c0a7, 32'h42f167f4} /* (27, 28, 4) {real, imag} */,
  {32'hc1b0ad47, 32'h41a3fd99} /* (27, 28, 3) {real, imag} */,
  {32'hc37ee45d, 32'h433e6ad0} /* (27, 28, 2) {real, imag} */,
  {32'h427b100a, 32'h41214214} /* (27, 28, 1) {real, imag} */,
  {32'h4379e00b, 32'h42801dfe} /* (27, 28, 0) {real, imag} */,
  {32'hc33e63ee, 32'hc3169d31} /* (27, 27, 31) {real, imag} */,
  {32'hc2e593d0, 32'hc13fccb1} /* (27, 27, 30) {real, imag} */,
  {32'hc1a9f50c, 32'hc1df377a} /* (27, 27, 29) {real, imag} */,
  {32'hbfbba5a0, 32'h42fdd4cc} /* (27, 27, 28) {real, imag} */,
  {32'h4248208e, 32'h42849050} /* (27, 27, 27) {real, imag} */,
  {32'h42c5e500, 32'h40b7f790} /* (27, 27, 26) {real, imag} */,
  {32'h42c2341f, 32'hc258c4be} /* (27, 27, 25) {real, imag} */,
  {32'hc13b32a4, 32'hc03ce310} /* (27, 27, 24) {real, imag} */,
  {32'hc203d425, 32'h40fb0ecc} /* (27, 27, 23) {real, imag} */,
  {32'hc095d9d8, 32'hc0bdbe4a} /* (27, 27, 22) {real, imag} */,
  {32'h422f3980, 32'hc151b87c} /* (27, 27, 21) {real, imag} */,
  {32'hc1f4ff38, 32'h40ef6fac} /* (27, 27, 20) {real, imag} */,
  {32'hc1cbd79b, 32'hc20f9955} /* (27, 27, 19) {real, imag} */,
  {32'hc1d9fd5d, 32'hc2342ced} /* (27, 27, 18) {real, imag} */,
  {32'h416a9ca6, 32'h412ddc14} /* (27, 27, 17) {real, imag} */,
  {32'hc11f2270, 32'h40efe100} /* (27, 27, 16) {real, imag} */,
  {32'hc0e9adfc, 32'hc11868a4} /* (27, 27, 15) {real, imag} */,
  {32'hc1bc1b75, 32'h3f034cc0} /* (27, 27, 14) {real, imag} */,
  {32'h3e970bc0, 32'hc1bc4e22} /* (27, 27, 13) {real, imag} */,
  {32'h40f00500, 32'h41508fd6} /* (27, 27, 12) {real, imag} */,
  {32'hc10a30ee, 32'h42274159} /* (27, 27, 11) {real, imag} */,
  {32'h424d72c9, 32'hc20d2f55} /* (27, 27, 10) {real, imag} */,
  {32'h421d66e3, 32'hc277c35e} /* (27, 27, 9) {real, imag} */,
  {32'h42cbdf46, 32'h42b1f924} /* (27, 27, 8) {real, imag} */,
  {32'h4291f24d, 32'h40f5cfb4} /* (27, 27, 7) {real, imag} */,
  {32'h4141e5f4, 32'hc28ec96f} /* (27, 27, 6) {real, imag} */,
  {32'hc1674a76, 32'h4218a405} /* (27, 27, 5) {real, imag} */,
  {32'hc2ac6e46, 32'hc15a97c0} /* (27, 27, 4) {real, imag} */,
  {32'h42aa6349, 32'hc283ca92} /* (27, 27, 3) {real, imag} */,
  {32'h42857742, 32'h40d88382} /* (27, 27, 2) {real, imag} */,
  {32'hc281fdef, 32'hc263789c} /* (27, 27, 1) {real, imag} */,
  {32'hc361851f, 32'hc2c1ffb6} /* (27, 27, 0) {real, imag} */,
  {32'hc3189ef0, 32'h4132b830} /* (27, 26, 31) {real, imag} */,
  {32'h429c4240, 32'hc2279cd5} /* (27, 26, 30) {real, imag} */,
  {32'hc11bfbed, 32'h42a3ec3a} /* (27, 26, 29) {real, imag} */,
  {32'hc2299de3, 32'hc207c03a} /* (27, 26, 28) {real, imag} */,
  {32'hc2a0f7b3, 32'hc0b1cbf6} /* (27, 26, 27) {real, imag} */,
  {32'h42b17f84, 32'h429e6544} /* (27, 26, 26) {real, imag} */,
  {32'hc23ab2dd, 32'h40c5ffbe} /* (27, 26, 25) {real, imag} */,
  {32'h4296f84e, 32'hc276296f} /* (27, 26, 24) {real, imag} */,
  {32'h41af0daa, 32'hc0c8827a} /* (27, 26, 23) {real, imag} */,
  {32'h42c4ba34, 32'h421911ce} /* (27, 26, 22) {real, imag} */,
  {32'hbfc87dc8, 32'h428c3801} /* (27, 26, 21) {real, imag} */,
  {32'h4133cbda, 32'hc1820551} /* (27, 26, 20) {real, imag} */,
  {32'hc19c07f4, 32'h42133156} /* (27, 26, 19) {real, imag} */,
  {32'h411ff960, 32'h40ce9cc8} /* (27, 26, 18) {real, imag} */,
  {32'hc1a0b6af, 32'h404c3d50} /* (27, 26, 17) {real, imag} */,
  {32'h40bd364c, 32'hc25d4a78} /* (27, 26, 16) {real, imag} */,
  {32'hc17a2536, 32'h4243cbab} /* (27, 26, 15) {real, imag} */,
  {32'hc24a6c0b, 32'h400323f0} /* (27, 26, 14) {real, imag} */,
  {32'hc18d8aa8, 32'h40e5b824} /* (27, 26, 13) {real, imag} */,
  {32'h41c45d23, 32'hc1ef8d4f} /* (27, 26, 12) {real, imag} */,
  {32'h41f5aa1e, 32'h41470f50} /* (27, 26, 11) {real, imag} */,
  {32'h4145cd8c, 32'h41c08da8} /* (27, 26, 10) {real, imag} */,
  {32'h421f5790, 32'h417ac8e7} /* (27, 26, 9) {real, imag} */,
  {32'h41d7caa2, 32'h41a34e02} /* (27, 26, 8) {real, imag} */,
  {32'hc2833c9e, 32'h3fc55ad8} /* (27, 26, 7) {real, imag} */,
  {32'hc1d12776, 32'h4163497c} /* (27, 26, 6) {real, imag} */,
  {32'h41a64e84, 32'h414b69a3} /* (27, 26, 5) {real, imag} */,
  {32'hc22c496f, 32'hc2c412c7} /* (27, 26, 4) {real, imag} */,
  {32'h40cb1f12, 32'h41b23813} /* (27, 26, 3) {real, imag} */,
  {32'h421643f4, 32'h42ad6d76} /* (27, 26, 2) {real, imag} */,
  {32'h418046b4, 32'hc314ce31} /* (27, 26, 1) {real, imag} */,
  {32'h4184ae53, 32'h421f18ce} /* (27, 26, 0) {real, imag} */,
  {32'h43435270, 32'h42bdec69} /* (27, 25, 31) {real, imag} */,
  {32'hc2ae4a4a, 32'hc22f6797} /* (27, 25, 30) {real, imag} */,
  {32'h42943a46, 32'h41d94b34} /* (27, 25, 29) {real, imag} */,
  {32'hc1540939, 32'hc2fdac48} /* (27, 25, 28) {real, imag} */,
  {32'hc22714bb, 32'h426b8fec} /* (27, 25, 27) {real, imag} */,
  {32'h428df186, 32'hc30bc5f5} /* (27, 25, 26) {real, imag} */,
  {32'hc2d64901, 32'h410e4604} /* (27, 25, 25) {real, imag} */,
  {32'hc28db922, 32'hc257d5a6} /* (27, 25, 24) {real, imag} */,
  {32'h4288fcd9, 32'h41d805b4} /* (27, 25, 23) {real, imag} */,
  {32'h418f13e7, 32'h4151fb00} /* (27, 25, 22) {real, imag} */,
  {32'h411ea9b5, 32'hc291d3d6} /* (27, 25, 21) {real, imag} */,
  {32'h410e2e54, 32'h3fbea360} /* (27, 25, 20) {real, imag} */,
  {32'h421eb368, 32'hc16f5f74} /* (27, 25, 19) {real, imag} */,
  {32'hbfe0c410, 32'h41504639} /* (27, 25, 18) {real, imag} */,
  {32'h3f555380, 32'h417e3bac} /* (27, 25, 17) {real, imag} */,
  {32'hc1e429d9, 32'h4115d6f8} /* (27, 25, 16) {real, imag} */,
  {32'h418dea1c, 32'hc1dace3e} /* (27, 25, 15) {real, imag} */,
  {32'hc1d5d361, 32'hc19fa4dc} /* (27, 25, 14) {real, imag} */,
  {32'hc21d4748, 32'h41a7591a} /* (27, 25, 13) {real, imag} */,
  {32'h4135ff6c, 32'hc2214337} /* (27, 25, 12) {real, imag} */,
  {32'hc2146361, 32'h42390346} /* (27, 25, 11) {real, imag} */,
  {32'hc1c311d7, 32'hc21ad2f5} /* (27, 25, 10) {real, imag} */,
  {32'hc1a0f03b, 32'hc2b3e79e} /* (27, 25, 9) {real, imag} */,
  {32'h42d77162, 32'h42ca7321} /* (27, 25, 8) {real, imag} */,
  {32'h4311e7db, 32'hc28fd714} /* (27, 25, 7) {real, imag} */,
  {32'h421ae930, 32'hc03ace00} /* (27, 25, 6) {real, imag} */,
  {32'h42d4ee56, 32'hc06e9ca0} /* (27, 25, 5) {real, imag} */,
  {32'hc1a7726c, 32'hc1e80466} /* (27, 25, 4) {real, imag} */,
  {32'hc23d7d8b, 32'h42b1539d} /* (27, 25, 3) {real, imag} */,
  {32'hc1f78042, 32'h41e6f84a} /* (27, 25, 2) {real, imag} */,
  {32'hbfaef3c0, 32'h42bf3525} /* (27, 25, 1) {real, imag} */,
  {32'hc288a5c1, 32'hc1369a30} /* (27, 25, 0) {real, imag} */,
  {32'hc287a8b9, 32'hc120d410} /* (27, 24, 31) {real, imag} */,
  {32'hc282b0fa, 32'h41da510b} /* (27, 24, 30) {real, imag} */,
  {32'h3fb5c7a0, 32'h422525e2} /* (27, 24, 29) {real, imag} */,
  {32'hc2b94d3b, 32'hc208eab5} /* (27, 24, 28) {real, imag} */,
  {32'hc2099d42, 32'hc10aa619} /* (27, 24, 27) {real, imag} */,
  {32'hc283c939, 32'hc220553a} /* (27, 24, 26) {real, imag} */,
  {32'h41f60890, 32'h41c02e8d} /* (27, 24, 25) {real, imag} */,
  {32'h40472380, 32'hc1d72de8} /* (27, 24, 24) {real, imag} */,
  {32'h4213ef06, 32'hc190864f} /* (27, 24, 23) {real, imag} */,
  {32'hc1e2ad8d, 32'hc1bc9e20} /* (27, 24, 22) {real, imag} */,
  {32'h418ce2ca, 32'h4224f210} /* (27, 24, 21) {real, imag} */,
  {32'hc1ad59bb, 32'hc07b1ad8} /* (27, 24, 20) {real, imag} */,
  {32'hc0a42aa8, 32'h4160487c} /* (27, 24, 19) {real, imag} */,
  {32'h4204d2f0, 32'h401475f6} /* (27, 24, 18) {real, imag} */,
  {32'h3fa6b0b0, 32'h3fc1be40} /* (27, 24, 17) {real, imag} */,
  {32'h417237c8, 32'hc1b3e313} /* (27, 24, 16) {real, imag} */,
  {32'hc129333e, 32'hc1b9f8c4} /* (27, 24, 15) {real, imag} */,
  {32'hc1915f2c, 32'hc1732926} /* (27, 24, 14) {real, imag} */,
  {32'hc1477d3c, 32'hc1a5cef0} /* (27, 24, 13) {real, imag} */,
  {32'h41c4a2eb, 32'hc1cebc43} /* (27, 24, 12) {real, imag} */,
  {32'h41800e44, 32'h4254570a} /* (27, 24, 11) {real, imag} */,
  {32'hc277e2f0, 32'hc239d6f2} /* (27, 24, 10) {real, imag} */,
  {32'hc097c1c4, 32'h4222dfc8} /* (27, 24, 9) {real, imag} */,
  {32'h42c23854, 32'h42971b08} /* (27, 24, 8) {real, imag} */,
  {32'h42ce2114, 32'h416badea} /* (27, 24, 7) {real, imag} */,
  {32'hc1e5b411, 32'h42869efa} /* (27, 24, 6) {real, imag} */,
  {32'h421a2c9e, 32'hc1beb3bc} /* (27, 24, 5) {real, imag} */,
  {32'hc22ab7ea, 32'hc20dd6cf} /* (27, 24, 4) {real, imag} */,
  {32'h41eb28d2, 32'h423e4fde} /* (27, 24, 3) {real, imag} */,
  {32'h4231ea65, 32'hc11a6006} /* (27, 24, 2) {real, imag} */,
  {32'hc24ddfec, 32'hc30b1077} /* (27, 24, 1) {real, imag} */,
  {32'hc2b53461, 32'hc11b7f82} /* (27, 24, 0) {real, imag} */,
  {32'hc22872c1, 32'hc29fd4c3} /* (27, 23, 31) {real, imag} */,
  {32'h41ddc05a, 32'h42a675be} /* (27, 23, 30) {real, imag} */,
  {32'h4223ac22, 32'h42a3671f} /* (27, 23, 29) {real, imag} */,
  {32'h429aca3f, 32'h41910ac0} /* (27, 23, 28) {real, imag} */,
  {32'h4216bf28, 32'hc09a33bc} /* (27, 23, 27) {real, imag} */,
  {32'hc1a28200, 32'hc290e347} /* (27, 23, 26) {real, imag} */,
  {32'h428a8987, 32'hc2302983} /* (27, 23, 25) {real, imag} */,
  {32'hc1695ad4, 32'h411c2498} /* (27, 23, 24) {real, imag} */,
  {32'h3fb9bdd0, 32'h4095846c} /* (27, 23, 23) {real, imag} */,
  {32'hc1c159b4, 32'h40fb4dfc} /* (27, 23, 22) {real, imag} */,
  {32'h415c4f08, 32'h411bb682} /* (27, 23, 21) {real, imag} */,
  {32'h4189bda1, 32'hc0971b28} /* (27, 23, 20) {real, imag} */,
  {32'hc1345e18, 32'h415dab1e} /* (27, 23, 19) {real, imag} */,
  {32'h41a17a12, 32'h412b0134} /* (27, 23, 18) {real, imag} */,
  {32'hc1e610fe, 32'h4205860d} /* (27, 23, 17) {real, imag} */,
  {32'h41b47e78, 32'hc166ccb0} /* (27, 23, 16) {real, imag} */,
  {32'hc1d52b76, 32'hc16b72fc} /* (27, 23, 15) {real, imag} */,
  {32'hc0fb6978, 32'h41cd6f72} /* (27, 23, 14) {real, imag} */,
  {32'h40db56d0, 32'hc1b07989} /* (27, 23, 13) {real, imag} */,
  {32'hc1ff57b7, 32'hc18ddc3a} /* (27, 23, 12) {real, imag} */,
  {32'h42403b46, 32'hc203b502} /* (27, 23, 11) {real, imag} */,
  {32'h425f2208, 32'hc20fa734} /* (27, 23, 10) {real, imag} */,
  {32'hc1b8742f, 32'hc0af4728} /* (27, 23, 9) {real, imag} */,
  {32'hc143f394, 32'hc0ba8ca9} /* (27, 23, 8) {real, imag} */,
  {32'hc13db7e6, 32'h413f4e4c} /* (27, 23, 7) {real, imag} */,
  {32'hc2b036df, 32'h4246ef6a} /* (27, 23, 6) {real, imag} */,
  {32'hc28b3866, 32'hc25eb5f6} /* (27, 23, 5) {real, imag} */,
  {32'hc11cde78, 32'h42489b50} /* (27, 23, 4) {real, imag} */,
  {32'hc1393d3a, 32'hc2054e12} /* (27, 23, 3) {real, imag} */,
  {32'hc2b91e6a, 32'hc1bdb18a} /* (27, 23, 2) {real, imag} */,
  {32'h431189c3, 32'hc284f3e5} /* (27, 23, 1) {real, imag} */,
  {32'hc298775e, 32'hc1496648} /* (27, 23, 0) {real, imag} */,
  {32'h42abd910, 32'h4225679c} /* (27, 22, 31) {real, imag} */,
  {32'h422b4941, 32'hc0690f30} /* (27, 22, 30) {real, imag} */,
  {32'hc20247d3, 32'h410eeb34} /* (27, 22, 29) {real, imag} */,
  {32'h41cb8478, 32'h412d2eca} /* (27, 22, 28) {real, imag} */,
  {32'h4115755c, 32'hc27e9391} /* (27, 22, 27) {real, imag} */,
  {32'hc2265e07, 32'h4254b02e} /* (27, 22, 26) {real, imag} */,
  {32'hc17736c2, 32'hc0a8f950} /* (27, 22, 25) {real, imag} */,
  {32'h4284a290, 32'hc195edee} /* (27, 22, 24) {real, imag} */,
  {32'hc23e3b68, 32'h42261e6f} /* (27, 22, 23) {real, imag} */,
  {32'hc1c6ffd4, 32'h422d9dee} /* (27, 22, 22) {real, imag} */,
  {32'h41e6eed2, 32'h4188c17b} /* (27, 22, 21) {real, imag} */,
  {32'hc0e93548, 32'hc114f7fc} /* (27, 22, 20) {real, imag} */,
  {32'hc1f45967, 32'hbfb98388} /* (27, 22, 19) {real, imag} */,
  {32'h405165cc, 32'h3e842ba0} /* (27, 22, 18) {real, imag} */,
  {32'hc024d786, 32'hc1f7e79d} /* (27, 22, 17) {real, imag} */,
  {32'h412a87f8, 32'h4206a288} /* (27, 22, 16) {real, imag} */,
  {32'hc09438c3, 32'h3fc56630} /* (27, 22, 15) {real, imag} */,
  {32'h41183eb9, 32'hc09a298a} /* (27, 22, 14) {real, imag} */,
  {32'h41885949, 32'hc1c339e6} /* (27, 22, 13) {real, imag} */,
  {32'hc1cb4ab8, 32'h400b14c0} /* (27, 22, 12) {real, imag} */,
  {32'h410cb52d, 32'hc0561348} /* (27, 22, 11) {real, imag} */,
  {32'hc140f90c, 32'h41247b48} /* (27, 22, 10) {real, imag} */,
  {32'hc10b234a, 32'hc21e6b35} /* (27, 22, 9) {real, imag} */,
  {32'hc0a07ec0, 32'h4215063c} /* (27, 22, 8) {real, imag} */,
  {32'h42121abe, 32'hc0bc8cb0} /* (27, 22, 7) {real, imag} */,
  {32'hc06ebe80, 32'h408c8750} /* (27, 22, 6) {real, imag} */,
  {32'hc120c952, 32'hc15baa6c} /* (27, 22, 5) {real, imag} */,
  {32'h42791048, 32'hc259c0e2} /* (27, 22, 4) {real, imag} */,
  {32'h41b1985f, 32'h429aae78} /* (27, 22, 3) {real, imag} */,
  {32'hc08401e8, 32'h4203eaa5} /* (27, 22, 2) {real, imag} */,
  {32'hc2aa4e50, 32'hc151e152} /* (27, 22, 1) {real, imag} */,
  {32'h43030176, 32'hc2b92a64} /* (27, 22, 0) {real, imag} */,
  {32'hc236c863, 32'h422bf990} /* (27, 21, 31) {real, imag} */,
  {32'hc1de4097, 32'h41c601fa} /* (27, 21, 30) {real, imag} */,
  {32'h3f1cfb50, 32'h3f7e8620} /* (27, 21, 29) {real, imag} */,
  {32'hc0dcadbc, 32'hc2294075} /* (27, 21, 28) {real, imag} */,
  {32'h41d7193d, 32'hc02fb1d4} /* (27, 21, 27) {real, imag} */,
  {32'h425b225a, 32'h42382d75} /* (27, 21, 26) {real, imag} */,
  {32'hc1b91051, 32'h4133d34f} /* (27, 21, 25) {real, imag} */,
  {32'h4031b338, 32'hc15767fe} /* (27, 21, 24) {real, imag} */,
  {32'hbe57eb80, 32'h4292f808} /* (27, 21, 23) {real, imag} */,
  {32'hc2264d5c, 32'h4132bfda} /* (27, 21, 22) {real, imag} */,
  {32'h41070a84, 32'hc24fa8be} /* (27, 21, 21) {real, imag} */,
  {32'h40f16e33, 32'h401bf2d8} /* (27, 21, 20) {real, imag} */,
  {32'h416d5484, 32'hc0e8475b} /* (27, 21, 19) {real, imag} */,
  {32'h41168dcf, 32'hbf946800} /* (27, 21, 18) {real, imag} */,
  {32'hc0fce7a3, 32'h41c4b4de} /* (27, 21, 17) {real, imag} */,
  {32'h41004d4e, 32'h40453ae0} /* (27, 21, 16) {real, imag} */,
  {32'h40ea0225, 32'hc0d4f100} /* (27, 21, 15) {real, imag} */,
  {32'hc1229ce1, 32'h41a90c4a} /* (27, 21, 14) {real, imag} */,
  {32'h4182c355, 32'h3e29e060} /* (27, 21, 13) {real, imag} */,
  {32'h417fe532, 32'hc121f23a} /* (27, 21, 12) {real, imag} */,
  {32'h409cdaa0, 32'h41bf4efc} /* (27, 21, 11) {real, imag} */,
  {32'h4148b4a0, 32'h404bc518} /* (27, 21, 10) {real, imag} */,
  {32'h416e9592, 32'h405c4970} /* (27, 21, 9) {real, imag} */,
  {32'hc218dbb6, 32'h405d8d78} /* (27, 21, 8) {real, imag} */,
  {32'hc1fbbca9, 32'h4111271f} /* (27, 21, 7) {real, imag} */,
  {32'hc17a4600, 32'h420c0887} /* (27, 21, 6) {real, imag} */,
  {32'h428546ef, 32'hbfcef328} /* (27, 21, 5) {real, imag} */,
  {32'hc21cde74, 32'hc21d66db} /* (27, 21, 4) {real, imag} */,
  {32'hc113fadf, 32'h4204445a} /* (27, 21, 3) {real, imag} */,
  {32'h4217ff9e, 32'hc2774973} /* (27, 21, 2) {real, imag} */,
  {32'h42690c89, 32'hc116d3ec} /* (27, 21, 1) {real, imag} */,
  {32'hc27a006c, 32'hc2720b92} /* (27, 21, 0) {real, imag} */,
  {32'h4209c586, 32'h4114b129} /* (27, 20, 31) {real, imag} */,
  {32'hc1a6ba6f, 32'hc20b4443} /* (27, 20, 30) {real, imag} */,
  {32'hc084d89c, 32'hc147d7fb} /* (27, 20, 29) {real, imag} */,
  {32'hc184258b, 32'h418784bd} /* (27, 20, 28) {real, imag} */,
  {32'hbfaa8e50, 32'h42589cea} /* (27, 20, 27) {real, imag} */,
  {32'hc21835e2, 32'h409e26cc} /* (27, 20, 26) {real, imag} */,
  {32'h42414dd3, 32'hc208447c} /* (27, 20, 25) {real, imag} */,
  {32'h40ef5c94, 32'hc194d30e} /* (27, 20, 24) {real, imag} */,
  {32'h417e8c23, 32'hc136d282} /* (27, 20, 23) {real, imag} */,
  {32'h408af8c2, 32'h40c408d0} /* (27, 20, 22) {real, imag} */,
  {32'hc204aeda, 32'hc18968a3} /* (27, 20, 21) {real, imag} */,
  {32'hc14ba351, 32'h3fea0ea4} /* (27, 20, 20) {real, imag} */,
  {32'h3deafea0, 32'h41604dcd} /* (27, 20, 19) {real, imag} */,
  {32'h41471e86, 32'hc18dd6e4} /* (27, 20, 18) {real, imag} */,
  {32'h4075bd42, 32'hbf5e9170} /* (27, 20, 17) {real, imag} */,
  {32'h403fdf88, 32'h404865f4} /* (27, 20, 16) {real, imag} */,
  {32'h40add3e1, 32'hc1a05884} /* (27, 20, 15) {real, imag} */,
  {32'hbfda39ac, 32'h41017236} /* (27, 20, 14) {real, imag} */,
  {32'h40bf8916, 32'hc0d161d6} /* (27, 20, 13) {real, imag} */,
  {32'h41150217, 32'hbefe9150} /* (27, 20, 12) {real, imag} */,
  {32'h403c6b18, 32'h41c91b8f} /* (27, 20, 11) {real, imag} */,
  {32'hc1a18a12, 32'h40b74378} /* (27, 20, 10) {real, imag} */,
  {32'h41aca40e, 32'h41d608f3} /* (27, 20, 9) {real, imag} */,
  {32'h4229003a, 32'hc1c292c6} /* (27, 20, 8) {real, imag} */,
  {32'h40c7da78, 32'hc1cf477a} /* (27, 20, 7) {real, imag} */,
  {32'hc1b83d23, 32'hc208059c} /* (27, 20, 6) {real, imag} */,
  {32'h42291522, 32'hc1d25b3d} /* (27, 20, 5) {real, imag} */,
  {32'hc1b83ded, 32'h41e98477} /* (27, 20, 4) {real, imag} */,
  {32'hc1967712, 32'h421fa8eb} /* (27, 20, 3) {real, imag} */,
  {32'hc2300b8c, 32'h423d68f9} /* (27, 20, 2) {real, imag} */,
  {32'hc2063a4c, 32'h41880942} /* (27, 20, 1) {real, imag} */,
  {32'h426a3a66, 32'h41dd8460} /* (27, 20, 0) {real, imag} */,
  {32'hc1eeb720, 32'hc1d75d61} /* (27, 19, 31) {real, imag} */,
  {32'h40a4fc2c, 32'h41d8c436} /* (27, 19, 30) {real, imag} */,
  {32'h423ddde5, 32'hc19497e8} /* (27, 19, 29) {real, imag} */,
  {32'h40fcc967, 32'hc1210f74} /* (27, 19, 28) {real, imag} */,
  {32'h41f5d285, 32'h40347fc0} /* (27, 19, 27) {real, imag} */,
  {32'hc1cbe076, 32'hc1e97f34} /* (27, 19, 26) {real, imag} */,
  {32'h41a78db4, 32'hc04f9028} /* (27, 19, 25) {real, imag} */,
  {32'h419b7c00, 32'h4217fb96} /* (27, 19, 24) {real, imag} */,
  {32'h416720b2, 32'hc0c201ec} /* (27, 19, 23) {real, imag} */,
  {32'h3f1c3070, 32'h413fbf48} /* (27, 19, 22) {real, imag} */,
  {32'h411e3590, 32'hc0d09338} /* (27, 19, 21) {real, imag} */,
  {32'hc05bb776, 32'hc14c9842} /* (27, 19, 20) {real, imag} */,
  {32'hc14b5cca, 32'h41001794} /* (27, 19, 19) {real, imag} */,
  {32'hc056fa21, 32'h4200a5bf} /* (27, 19, 18) {real, imag} */,
  {32'h4060f484, 32'hc0ef78fb} /* (27, 19, 17) {real, imag} */,
  {32'h3f0dd680, 32'h40442d40} /* (27, 19, 16) {real, imag} */,
  {32'h40f6b2ae, 32'hc00053be} /* (27, 19, 15) {real, imag} */,
  {32'hc114ceb2, 32'hc12ee45b} /* (27, 19, 14) {real, imag} */,
  {32'hbeca2050, 32'h40136e52} /* (27, 19, 13) {real, imag} */,
  {32'h41637722, 32'h4080f538} /* (27, 19, 12) {real, imag} */,
  {32'hc1b08b15, 32'hc1a3a3d0} /* (27, 19, 11) {real, imag} */,
  {32'h419f075a, 32'hc23bd273} /* (27, 19, 10) {real, imag} */,
  {32'hc1983655, 32'h42236ce6} /* (27, 19, 9) {real, imag} */,
  {32'h41026563, 32'h4091f78c} /* (27, 19, 8) {real, imag} */,
  {32'h41d09fc8, 32'h420a63b6} /* (27, 19, 7) {real, imag} */,
  {32'h420fc01c, 32'hc106bf7c} /* (27, 19, 6) {real, imag} */,
  {32'hc23d7d10, 32'h41e3ebda} /* (27, 19, 5) {real, imag} */,
  {32'h4067799e, 32'h41c5243a} /* (27, 19, 4) {real, imag} */,
  {32'h425b6cb7, 32'hc1a11434} /* (27, 19, 3) {real, imag} */,
  {32'hc07c7b2f, 32'hc1fb40c6} /* (27, 19, 2) {real, imag} */,
  {32'h40bf36d0, 32'h42169cb4} /* (27, 19, 1) {real, imag} */,
  {32'hc23d9c75, 32'hc24cccd4} /* (27, 19, 0) {real, imag} */,
  {32'hc271c8d4, 32'hc1433f56} /* (27, 18, 31) {real, imag} */,
  {32'h428ad44d, 32'hc1c45782} /* (27, 18, 30) {real, imag} */,
  {32'h417e169a, 32'h40db7af8} /* (27, 18, 29) {real, imag} */,
  {32'hc23595d8, 32'h41b69a20} /* (27, 18, 28) {real, imag} */,
  {32'h401a1428, 32'hc22d1bc9} /* (27, 18, 27) {real, imag} */,
  {32'h40aaa800, 32'hc1ab5de5} /* (27, 18, 26) {real, imag} */,
  {32'hc0af8c74, 32'hc19b983e} /* (27, 18, 25) {real, imag} */,
  {32'h41bf3aed, 32'hc1580c70} /* (27, 18, 24) {real, imag} */,
  {32'hc085b06b, 32'hc2075c86} /* (27, 18, 23) {real, imag} */,
  {32'h41427e86, 32'hc17ee842} /* (27, 18, 22) {real, imag} */,
  {32'hc1b973c1, 32'h41b17ade} /* (27, 18, 21) {real, imag} */,
  {32'h41802c31, 32'h4134460e} /* (27, 18, 20) {real, imag} */,
  {32'h410275f8, 32'hc11d6759} /* (27, 18, 19) {real, imag} */,
  {32'h402f6868, 32'h412972ec} /* (27, 18, 18) {real, imag} */,
  {32'hc0e9ba44, 32'h407a02e2} /* (27, 18, 17) {real, imag} */,
  {32'h409862bc, 32'hc125a508} /* (27, 18, 16) {real, imag} */,
  {32'h411c014a, 32'h41837ca7} /* (27, 18, 15) {real, imag} */,
  {32'h4026e228, 32'h4127c0ce} /* (27, 18, 14) {real, imag} */,
  {32'h3fe9c1c0, 32'h3ff80b96} /* (27, 18, 13) {real, imag} */,
  {32'h3eb651c0, 32'h4180d5e0} /* (27, 18, 12) {real, imag} */,
  {32'h419f7efb, 32'h40c67806} /* (27, 18, 11) {real, imag} */,
  {32'hc194f7c3, 32'hc1129f3a} /* (27, 18, 10) {real, imag} */,
  {32'h410989ee, 32'hc1b07a2b} /* (27, 18, 9) {real, imag} */,
  {32'hc18dc809, 32'h41adfaa6} /* (27, 18, 8) {real, imag} */,
  {32'hc2281234, 32'h4221ae54} /* (27, 18, 7) {real, imag} */,
  {32'hc222cb11, 32'hc177a8c2} /* (27, 18, 6) {real, imag} */,
  {32'hc26088a4, 32'h410d6594} /* (27, 18, 5) {real, imag} */,
  {32'hc198886d, 32'hc0fd2e6e} /* (27, 18, 4) {real, imag} */,
  {32'hc1f7a89b, 32'hc1bc544c} /* (27, 18, 3) {real, imag} */,
  {32'hc0eab31c, 32'hc120b72d} /* (27, 18, 2) {real, imag} */,
  {32'hc1c945a5, 32'hc0f29997} /* (27, 18, 1) {real, imag} */,
  {32'h41a88a61, 32'hc202ee7b} /* (27, 18, 0) {real, imag} */,
  {32'h41f730f2, 32'hc14d3bcd} /* (27, 17, 31) {real, imag} */,
  {32'hc1b2b146, 32'h4149bf5c} /* (27, 17, 30) {real, imag} */,
  {32'hc15ea388, 32'hbf811a10} /* (27, 17, 29) {real, imag} */,
  {32'h4169e481, 32'hc097fd57} /* (27, 17, 28) {real, imag} */,
  {32'h40d2f6a0, 32'hc14067fc} /* (27, 17, 27) {real, imag} */,
  {32'h3fff4e4c, 32'h413fdc01} /* (27, 17, 26) {real, imag} */,
  {32'h40dfef6c, 32'h3dad6860} /* (27, 17, 25) {real, imag} */,
  {32'hc212a1c2, 32'hbf0ab660} /* (27, 17, 24) {real, imag} */,
  {32'hc058ae27, 32'hc055ed03} /* (27, 17, 23) {real, imag} */,
  {32'h41df66a5, 32'h419a8138} /* (27, 17, 22) {real, imag} */,
  {32'h406e78e4, 32'hc1037866} /* (27, 17, 21) {real, imag} */,
  {32'hc080f7e2, 32'hc1ac8568} /* (27, 17, 20) {real, imag} */,
  {32'h40d1ea71, 32'hc11e48ca} /* (27, 17, 19) {real, imag} */,
  {32'h3fa56e80, 32'hc122d969} /* (27, 17, 18) {real, imag} */,
  {32'h409884aa, 32'hc0a6dd98} /* (27, 17, 17) {real, imag} */,
  {32'hc0f2cef8, 32'hc166e9f8} /* (27, 17, 16) {real, imag} */,
  {32'h4116b1ff, 32'h40f4090e} /* (27, 17, 15) {real, imag} */,
  {32'hc1253cfa, 32'h3f4fd5f0} /* (27, 17, 14) {real, imag} */,
  {32'hc1571246, 32'h40cefd05} /* (27, 17, 13) {real, imag} */,
  {32'h409bceb4, 32'h3f3875b0} /* (27, 17, 12) {real, imag} */,
  {32'h402f8754, 32'h40765b92} /* (27, 17, 11) {real, imag} */,
  {32'h416aec7e, 32'hc18be0c6} /* (27, 17, 10) {real, imag} */,
  {32'h4135db4a, 32'hbfc34082} /* (27, 17, 9) {real, imag} */,
  {32'hc20a5fd8, 32'h405752c8} /* (27, 17, 8) {real, imag} */,
  {32'hc1d33275, 32'h40dca238} /* (27, 17, 7) {real, imag} */,
  {32'hc07f051e, 32'hc16f0443} /* (27, 17, 6) {real, imag} */,
  {32'hc224cf7a, 32'hc1477ec0} /* (27, 17, 5) {real, imag} */,
  {32'hc10b8a43, 32'h414ee416} /* (27, 17, 4) {real, imag} */,
  {32'h3e8db3b0, 32'h409eee26} /* (27, 17, 3) {real, imag} */,
  {32'hc0e3285e, 32'hc293c4a2} /* (27, 17, 2) {real, imag} */,
  {32'hc16017bc, 32'h413022eb} /* (27, 17, 1) {real, imag} */,
  {32'h4274ec83, 32'hc2a1a6d9} /* (27, 17, 0) {real, imag} */,
  {32'hc1be37e6, 32'hc1a1c1cb} /* (27, 16, 31) {real, imag} */,
  {32'hc1b59cc8, 32'h419d03d6} /* (27, 16, 30) {real, imag} */,
  {32'hc08ae172, 32'hc2029d88} /* (27, 16, 29) {real, imag} */,
  {32'h40d374e2, 32'h40f658e8} /* (27, 16, 28) {real, imag} */,
  {32'hbfa1ebd9, 32'hc07550c8} /* (27, 16, 27) {real, imag} */,
  {32'hc170de74, 32'hc05bfffd} /* (27, 16, 26) {real, imag} */,
  {32'h414a93f0, 32'hc1394ea6} /* (27, 16, 25) {real, imag} */,
  {32'h41074b54, 32'h411cc9b2} /* (27, 16, 24) {real, imag} */,
  {32'h419f9ca3, 32'hc1bdea5a} /* (27, 16, 23) {real, imag} */,
  {32'hc0b96cf9, 32'h4171a1f8} /* (27, 16, 22) {real, imag} */,
  {32'h4160a14c, 32'h411af68e} /* (27, 16, 21) {real, imag} */,
  {32'h40af7b6c, 32'hbf995a34} /* (27, 16, 20) {real, imag} */,
  {32'h40d2e928, 32'hc021528c} /* (27, 16, 19) {real, imag} */,
  {32'hc09101fc, 32'hc0fe2742} /* (27, 16, 18) {real, imag} */,
  {32'hbe59b240, 32'h40c3f829} /* (27, 16, 17) {real, imag} */,
  {32'hc0ab79e8, 32'h412f2dcd} /* (27, 16, 16) {real, imag} */,
  {32'h405f9a74, 32'hbe125da0} /* (27, 16, 15) {real, imag} */,
  {32'h4043b950, 32'hc032b9a4} /* (27, 16, 14) {real, imag} */,
  {32'hc19668a2, 32'h3f8246c8} /* (27, 16, 13) {real, imag} */,
  {32'hc1f16725, 32'hc107737a} /* (27, 16, 12) {real, imag} */,
  {32'hc1088114, 32'h410e9a0a} /* (27, 16, 11) {real, imag} */,
  {32'h4158893e, 32'h414d014a} /* (27, 16, 10) {real, imag} */,
  {32'hbf42dd60, 32'hbf925908} /* (27, 16, 9) {real, imag} */,
  {32'hc0146068, 32'hc2237d60} /* (27, 16, 8) {real, imag} */,
  {32'h410b222c, 32'h40576712} /* (27, 16, 7) {real, imag} */,
  {32'h4070f3fa, 32'h3fff73ca} /* (27, 16, 6) {real, imag} */,
  {32'h3f95d467, 32'hc1a87dc3} /* (27, 16, 5) {real, imag} */,
  {32'hc1849f0a, 32'hc1e059b0} /* (27, 16, 4) {real, imag} */,
  {32'h40894628, 32'h41ee4633} /* (27, 16, 3) {real, imag} */,
  {32'h3ac3c000, 32'hc03679c8} /* (27, 16, 2) {real, imag} */,
  {32'h3fc732d8, 32'hc16da2f2} /* (27, 16, 1) {real, imag} */,
  {32'h417d0344, 32'hbdcb1c80} /* (27, 16, 0) {real, imag} */,
  {32'hc2385235, 32'hc08be574} /* (27, 15, 31) {real, imag} */,
  {32'hc042ec1a, 32'hc183531a} /* (27, 15, 30) {real, imag} */,
  {32'hc141c98b, 32'hc10849e5} /* (27, 15, 29) {real, imag} */,
  {32'h40d01288, 32'h41602bac} /* (27, 15, 28) {real, imag} */,
  {32'h3fe31780, 32'hc08f0dc2} /* (27, 15, 27) {real, imag} */,
  {32'hc09c3052, 32'hc1c72f6e} /* (27, 15, 26) {real, imag} */,
  {32'hc1b88880, 32'h411284cc} /* (27, 15, 25) {real, imag} */,
  {32'h3e5afdc0, 32'hbf6d5460} /* (27, 15, 24) {real, imag} */,
  {32'hc151f81e, 32'h4120b66c} /* (27, 15, 23) {real, imag} */,
  {32'hc15b06c4, 32'hc11ae462} /* (27, 15, 22) {real, imag} */,
  {32'h409817a8, 32'hbf386db0} /* (27, 15, 21) {real, imag} */,
  {32'hc11b0c50, 32'hc087addc} /* (27, 15, 20) {real, imag} */,
  {32'hc03d958d, 32'hc12a5e7c} /* (27, 15, 19) {real, imag} */,
  {32'hc1477736, 32'hc16a0e03} /* (27, 15, 18) {real, imag} */,
  {32'h3f8ce238, 32'hbeeba5c0} /* (27, 15, 17) {real, imag} */,
  {32'h4118497a, 32'h40dbc5d0} /* (27, 15, 16) {real, imag} */,
  {32'hc02d9a4c, 32'h40463598} /* (27, 15, 15) {real, imag} */,
  {32'hc085b550, 32'hbdd7f380} /* (27, 15, 14) {real, imag} */,
  {32'h40bdda0c, 32'h3eb755c0} /* (27, 15, 13) {real, imag} */,
  {32'hbf5b8078, 32'hc0ff717e} /* (27, 15, 12) {real, imag} */,
  {32'h403084a0, 32'h41b1e54a} /* (27, 15, 11) {real, imag} */,
  {32'h4124ce02, 32'h40f60bec} /* (27, 15, 10) {real, imag} */,
  {32'hc10d2972, 32'hc1399f30} /* (27, 15, 9) {real, imag} */,
  {32'h41e40cb8, 32'h4107d9d8} /* (27, 15, 8) {real, imag} */,
  {32'hc1dd6cd8, 32'h40dd4599} /* (27, 15, 7) {real, imag} */,
  {32'hc1acb186, 32'hc2184b0e} /* (27, 15, 6) {real, imag} */,
  {32'h42893b5c, 32'hc0543f65} /* (27, 15, 5) {real, imag} */,
  {32'hc1d85aca, 32'hc1916f54} /* (27, 15, 4) {real, imag} */,
  {32'h4119e4a5, 32'hbfec6e2a} /* (27, 15, 3) {real, imag} */,
  {32'hc144fa32, 32'h42024792} /* (27, 15, 2) {real, imag} */,
  {32'hbfc2b4e0, 32'h4238746a} /* (27, 15, 1) {real, imag} */,
  {32'h3f336c58, 32'h41196b2a} /* (27, 15, 0) {real, imag} */,
  {32'hbf5f2358, 32'hc28a24e4} /* (27, 14, 31) {real, imag} */,
  {32'hc19aa6bd, 32'h420aa28e} /* (27, 14, 30) {real, imag} */,
  {32'h414c5552, 32'h416a758e} /* (27, 14, 29) {real, imag} */,
  {32'hc1778a13, 32'h427b9a17} /* (27, 14, 28) {real, imag} */,
  {32'hc10eb16a, 32'h40659e4a} /* (27, 14, 27) {real, imag} */,
  {32'h421c1709, 32'h422ea242} /* (27, 14, 26) {real, imag} */,
  {32'hc2209ff9, 32'h4181354a} /* (27, 14, 25) {real, imag} */,
  {32'hc1a51eac, 32'hc1df73b4} /* (27, 14, 24) {real, imag} */,
  {32'h410a6fd5, 32'hc0f6ab62} /* (27, 14, 23) {real, imag} */,
  {32'h41160a3c, 32'hc21503bf} /* (27, 14, 22) {real, imag} */,
  {32'h4131a0d1, 32'h3e2ff160} /* (27, 14, 21) {real, imag} */,
  {32'h40a8ea5e, 32'h41b11ece} /* (27, 14, 20) {real, imag} */,
  {32'h40f470a7, 32'h41186616} /* (27, 14, 19) {real, imag} */,
  {32'hc0f72706, 32'h404ce638} /* (27, 14, 18) {real, imag} */,
  {32'h407a342e, 32'hc0a08620} /* (27, 14, 17) {real, imag} */,
  {32'hc0699f72, 32'h3fa4c778} /* (27, 14, 16) {real, imag} */,
  {32'h40f53763, 32'h414e3cbc} /* (27, 14, 15) {real, imag} */,
  {32'hc04918dc, 32'hc0328958} /* (27, 14, 14) {real, imag} */,
  {32'h4112b06e, 32'hc09166ec} /* (27, 14, 13) {real, imag} */,
  {32'h40d4a77c, 32'h41d83d38} /* (27, 14, 12) {real, imag} */,
  {32'h4168ef17, 32'hc0e7bb01} /* (27, 14, 11) {real, imag} */,
  {32'h42260c27, 32'h41c5315d} /* (27, 14, 10) {real, imag} */,
  {32'hc1f4c7fc, 32'hc10e4a67} /* (27, 14, 9) {real, imag} */,
  {32'hc101cc2c, 32'hbf0cafb0} /* (27, 14, 8) {real, imag} */,
  {32'h417ed071, 32'h40cb7ac6} /* (27, 14, 7) {real, imag} */,
  {32'h410074bd, 32'hc0f1ee7c} /* (27, 14, 6) {real, imag} */,
  {32'h41fb5b2b, 32'h3e242720} /* (27, 14, 5) {real, imag} */,
  {32'hc11a7875, 32'h41407624} /* (27, 14, 4) {real, imag} */,
  {32'h41ce82e7, 32'h4284162e} /* (27, 14, 3) {real, imag} */,
  {32'h3e96ab80, 32'hc2961075} /* (27, 14, 2) {real, imag} */,
  {32'hc103a35c, 32'h419d35d1} /* (27, 14, 1) {real, imag} */,
  {32'h40d3c717, 32'hc1bf5986} /* (27, 14, 0) {real, imag} */,
  {32'h42080834, 32'h41713f5a} /* (27, 13, 31) {real, imag} */,
  {32'h413fa9cd, 32'h41729d78} /* (27, 13, 30) {real, imag} */,
  {32'hc22229b8, 32'hc07a81f8} /* (27, 13, 29) {real, imag} */,
  {32'h42696148, 32'hc0e75d83} /* (27, 13, 28) {real, imag} */,
  {32'hc2a36170, 32'h41735890} /* (27, 13, 27) {real, imag} */,
  {32'h40f2226c, 32'h403d473c} /* (27, 13, 26) {real, imag} */,
  {32'hc1467a1a, 32'hc19c30ae} /* (27, 13, 25) {real, imag} */,
  {32'hc204192e, 32'h4141a90c} /* (27, 13, 24) {real, imag} */,
  {32'hc1c0be85, 32'hc1c1eaac} /* (27, 13, 23) {real, imag} */,
  {32'h41e4293b, 32'h41678a76} /* (27, 13, 22) {real, imag} */,
  {32'hc199ff5b, 32'hc0302474} /* (27, 13, 21) {real, imag} */,
  {32'hc043e89e, 32'hc172e542} /* (27, 13, 20) {real, imag} */,
  {32'h407d0bc4, 32'hc19562d1} /* (27, 13, 19) {real, imag} */,
  {32'h40436a5a, 32'hc1227c04} /* (27, 13, 18) {real, imag} */,
  {32'hc121ab96, 32'h40be0252} /* (27, 13, 17) {real, imag} */,
  {32'h4154af20, 32'h40e4fac2} /* (27, 13, 16) {real, imag} */,
  {32'hc06a4150, 32'hc15ba4df} /* (27, 13, 15) {real, imag} */,
  {32'hc1120456, 32'hc0396cee} /* (27, 13, 14) {real, imag} */,
  {32'h4065a85c, 32'hc114474a} /* (27, 13, 13) {real, imag} */,
  {32'hc06aba3e, 32'h4009c59e} /* (27, 13, 12) {real, imag} */,
  {32'h41ccd305, 32'h41934924} /* (27, 13, 11) {real, imag} */,
  {32'h410d00be, 32'hc104f360} /* (27, 13, 10) {real, imag} */,
  {32'h417ec856, 32'h42139c2e} /* (27, 13, 9) {real, imag} */,
  {32'h40d15ed0, 32'h3f300ec0} /* (27, 13, 8) {real, imag} */,
  {32'h423ea288, 32'h421f04f5} /* (27, 13, 7) {real, imag} */,
  {32'hc1e4d8f7, 32'hc19985b2} /* (27, 13, 6) {real, imag} */,
  {32'h41fa98e1, 32'h41badc3e} /* (27, 13, 5) {real, imag} */,
  {32'hc20cca6e, 32'h41015664} /* (27, 13, 4) {real, imag} */,
  {32'hc2000af0, 32'h41b8a0e5} /* (27, 13, 3) {real, imag} */,
  {32'h418ebc06, 32'hc1f4a9ea} /* (27, 13, 2) {real, imag} */,
  {32'hc10b0af9, 32'h40d25bf0} /* (27, 13, 1) {real, imag} */,
  {32'hc234e37c, 32'h404f699c} /* (27, 13, 0) {real, imag} */,
  {32'h41ab26b3, 32'h422df8a6} /* (27, 12, 31) {real, imag} */,
  {32'hc0a03d16, 32'hc0c57970} /* (27, 12, 30) {real, imag} */,
  {32'h4222ef4a, 32'hc1c0fd9a} /* (27, 12, 29) {real, imag} */,
  {32'hc29ff198, 32'hc267f0e4} /* (27, 12, 28) {real, imag} */,
  {32'hc1980a6d, 32'h4215433d} /* (27, 12, 27) {real, imag} */,
  {32'h422e4839, 32'hc1672653} /* (27, 12, 26) {real, imag} */,
  {32'h40f02eee, 32'h426de3d5} /* (27, 12, 25) {real, imag} */,
  {32'hc0c68c4a, 32'hc10142cb} /* (27, 12, 24) {real, imag} */,
  {32'h42311b64, 32'h419410ca} /* (27, 12, 23) {real, imag} */,
  {32'hc1703634, 32'h418609d8} /* (27, 12, 22) {real, imag} */,
  {32'h418c88de, 32'h419c4d8c} /* (27, 12, 21) {real, imag} */,
  {32'h401190cc, 32'hbe72b980} /* (27, 12, 20) {real, imag} */,
  {32'hc1976583, 32'h408c4ea4} /* (27, 12, 19) {real, imag} */,
  {32'hc18654a4, 32'hc0de997e} /* (27, 12, 18) {real, imag} */,
  {32'hc12dad96, 32'h411ad150} /* (27, 12, 17) {real, imag} */,
  {32'h409afc9c, 32'hc0f323c4} /* (27, 12, 16) {real, imag} */,
  {32'h40791d36, 32'h40a40d00} /* (27, 12, 15) {real, imag} */,
  {32'hc0279a3c, 32'hc08e1fe2} /* (27, 12, 14) {real, imag} */,
  {32'hc119c6c8, 32'h400e3650} /* (27, 12, 13) {real, imag} */,
  {32'h412a01d3, 32'hc1dcdc62} /* (27, 12, 12) {real, imag} */,
  {32'hc080d81a, 32'h4130f0fa} /* (27, 12, 11) {real, imag} */,
  {32'h411ee774, 32'h420de55b} /* (27, 12, 10) {real, imag} */,
  {32'hc13cde58, 32'h420f4c95} /* (27, 12, 9) {real, imag} */,
  {32'h4182676a, 32'hc119ddfb} /* (27, 12, 8) {real, imag} */,
  {32'h3e9cdc20, 32'hc0839458} /* (27, 12, 7) {real, imag} */,
  {32'hc25f70d1, 32'hbd24f100} /* (27, 12, 6) {real, imag} */,
  {32'hc25b8076, 32'h423a1ef3} /* (27, 12, 5) {real, imag} */,
  {32'h423f5e01, 32'h42033124} /* (27, 12, 4) {real, imag} */,
  {32'hc1a9c614, 32'hc135fd83} /* (27, 12, 3) {real, imag} */,
  {32'h4137ae95, 32'h41fca544} /* (27, 12, 2) {real, imag} */,
  {32'h422ac6d8, 32'h422c003a} /* (27, 12, 1) {real, imag} */,
  {32'h4239fd00, 32'h41bfd97c} /* (27, 12, 0) {real, imag} */,
  {32'hbf9efe60, 32'hc29d6962} /* (27, 11, 31) {real, imag} */,
  {32'hc1489a30, 32'hc1e59765} /* (27, 11, 30) {real, imag} */,
  {32'h41a4d93e, 32'hc106740e} /* (27, 11, 29) {real, imag} */,
  {32'hc1e77460, 32'hc2682b8e} /* (27, 11, 28) {real, imag} */,
  {32'hc1bdb58d, 32'h42b170a3} /* (27, 11, 27) {real, imag} */,
  {32'hc03642ec, 32'h418095b8} /* (27, 11, 26) {real, imag} */,
  {32'h3f2c0288, 32'hc2a6ce54} /* (27, 11, 25) {real, imag} */,
  {32'hbf973328, 32'h420c67e1} /* (27, 11, 24) {real, imag} */,
  {32'h4171e8d0, 32'h41cf5aeb} /* (27, 11, 23) {real, imag} */,
  {32'hc110ea18, 32'h40c1ecdc} /* (27, 11, 22) {real, imag} */,
  {32'h41378fcc, 32'h41aa9380} /* (27, 11, 21) {real, imag} */,
  {32'h409a71b2, 32'h3fbc46e8} /* (27, 11, 20) {real, imag} */,
  {32'h41d13bf3, 32'hc17fd8dc} /* (27, 11, 19) {real, imag} */,
  {32'h41d16aec, 32'h413148d4} /* (27, 11, 18) {real, imag} */,
  {32'hc11a0f62, 32'hbe9c7fe0} /* (27, 11, 17) {real, imag} */,
  {32'hbf9d8d00, 32'hc1b20dfa} /* (27, 11, 16) {real, imag} */,
  {32'hc0c48b3d, 32'h419cb6da} /* (27, 11, 15) {real, imag} */,
  {32'hc1131ae8, 32'h41955686} /* (27, 11, 14) {real, imag} */,
  {32'hc1327272, 32'hc1c7516e} /* (27, 11, 13) {real, imag} */,
  {32'hc1c01e28, 32'h400f1f9c} /* (27, 11, 12) {real, imag} */,
  {32'h40b0a2b8, 32'hc1e9f294} /* (27, 11, 11) {real, imag} */,
  {32'hc22bb352, 32'hc22dc3ba} /* (27, 11, 10) {real, imag} */,
  {32'h40b00e35, 32'hc2222a24} /* (27, 11, 9) {real, imag} */,
  {32'hc184f04e, 32'h40d95326} /* (27, 11, 8) {real, imag} */,
  {32'h4136632a, 32'hbfe86260} /* (27, 11, 7) {real, imag} */,
  {32'h418e77f2, 32'h3f163d70} /* (27, 11, 6) {real, imag} */,
  {32'hc2372034, 32'hc160bce0} /* (27, 11, 5) {real, imag} */,
  {32'h42dfb864, 32'hc13596a8} /* (27, 11, 4) {real, imag} */,
  {32'h41cd5280, 32'hc1f64f6d} /* (27, 11, 3) {real, imag} */,
  {32'hc1d73ea6, 32'hc2250068} /* (27, 11, 2) {real, imag} */,
  {32'h42034e15, 32'hc033d090} /* (27, 11, 1) {real, imag} */,
  {32'h41c8f1b3, 32'hc2b0baaa} /* (27, 11, 0) {real, imag} */,
  {32'hc2a0e4b3, 32'h422d7689} /* (27, 10, 31) {real, imag} */,
  {32'hc08bc6f8, 32'hc219e14c} /* (27, 10, 30) {real, imag} */,
  {32'hc22f0380, 32'hc184f5d0} /* (27, 10, 29) {real, imag} */,
  {32'h4224ff5e, 32'hc2063f81} /* (27, 10, 28) {real, imag} */,
  {32'h4274999a, 32'hc17ea65e} /* (27, 10, 27) {real, imag} */,
  {32'hc1efcb06, 32'hc078b072} /* (27, 10, 26) {real, imag} */,
  {32'h41f0b1c7, 32'hc24c2358} /* (27, 10, 25) {real, imag} */,
  {32'hc2158f5d, 32'h41829078} /* (27, 10, 24) {real, imag} */,
  {32'hc17d6b16, 32'h420d9c0b} /* (27, 10, 23) {real, imag} */,
  {32'h42258418, 32'hc1f6ac0a} /* (27, 10, 22) {real, imag} */,
  {32'hc012b140, 32'h4217fec2} /* (27, 10, 21) {real, imag} */,
  {32'h41316b03, 32'h4138d334} /* (27, 10, 20) {real, imag} */,
  {32'h3fd4fcb0, 32'h41526390} /* (27, 10, 19) {real, imag} */,
  {32'hc0508ac0, 32'hc08b00b0} /* (27, 10, 18) {real, imag} */,
  {32'h4137e060, 32'hc1ed3151} /* (27, 10, 17) {real, imag} */,
  {32'hbfb886f0, 32'h4098b3e0} /* (27, 10, 16) {real, imag} */,
  {32'h3e03d000, 32'h415ebe66} /* (27, 10, 15) {real, imag} */,
  {32'h40db2ce0, 32'h404a6210} /* (27, 10, 14) {real, imag} */,
  {32'h41a33a69, 32'hc0cd5610} /* (27, 10, 13) {real, imag} */,
  {32'hc22bc93e, 32'hc1085c10} /* (27, 10, 12) {real, imag} */,
  {32'h41d27a33, 32'hc1872c4a} /* (27, 10, 11) {real, imag} */,
  {32'hc067f488, 32'h40d79028} /* (27, 10, 10) {real, imag} */,
  {32'h41143e76, 32'h3fd1c660} /* (27, 10, 9) {real, imag} */,
  {32'hc12e06cf, 32'hc229de50} /* (27, 10, 8) {real, imag} */,
  {32'h42a44b78, 32'h4216436c} /* (27, 10, 7) {real, imag} */,
  {32'hc28f926c, 32'hc167ab24} /* (27, 10, 6) {real, imag} */,
  {32'h41ac3770, 32'hc18831ad} /* (27, 10, 5) {real, imag} */,
  {32'hc195b5f2, 32'h4252f9e3} /* (27, 10, 4) {real, imag} */,
  {32'hc2a261e3, 32'h42c7b439} /* (27, 10, 3) {real, imag} */,
  {32'hc29ec0b2, 32'hc2a35c64} /* (27, 10, 2) {real, imag} */,
  {32'h42c3a8e9, 32'h429d4a72} /* (27, 10, 1) {real, imag} */,
  {32'hc243d364, 32'h4287d7dd} /* (27, 10, 0) {real, imag} */,
  {32'hc23fb772, 32'h425dd7bb} /* (27, 9, 31) {real, imag} */,
  {32'h42268b19, 32'h42b31e5c} /* (27, 9, 30) {real, imag} */,
  {32'h42814634, 32'h40a02580} /* (27, 9, 29) {real, imag} */,
  {32'hc2535846, 32'hc2c884b1} /* (27, 9, 28) {real, imag} */,
  {32'hc1788e70, 32'hc2a43a7b} /* (27, 9, 27) {real, imag} */,
  {32'hc29965fc, 32'hc2bfe2d4} /* (27, 9, 26) {real, imag} */,
  {32'h4251041a, 32'h4240c4c2} /* (27, 9, 25) {real, imag} */,
  {32'h41bbff75, 32'hc2228d56} /* (27, 9, 24) {real, imag} */,
  {32'h424240bb, 32'h41e430c4} /* (27, 9, 23) {real, imag} */,
  {32'h4156cd5c, 32'h4089a28c} /* (27, 9, 22) {real, imag} */,
  {32'hc23592da, 32'hc1ea8a98} /* (27, 9, 21) {real, imag} */,
  {32'h418177b6, 32'h40e19748} /* (27, 9, 20) {real, imag} */,
  {32'h4135a5a0, 32'h4171ee6a} /* (27, 9, 19) {real, imag} */,
  {32'hc10cd778, 32'hc0eef115} /* (27, 9, 18) {real, imag} */,
  {32'h42500a7e, 32'h4140a10b} /* (27, 9, 17) {real, imag} */,
  {32'hc2600372, 32'h413695ee} /* (27, 9, 16) {real, imag} */,
  {32'hc0c16780, 32'hc1b35102} /* (27, 9, 15) {real, imag} */,
  {32'h41a0f378, 32'hc104da26} /* (27, 9, 14) {real, imag} */,
  {32'h41dc11be, 32'h415e106a} /* (27, 9, 13) {real, imag} */,
  {32'hc1a8c23a, 32'h40c20d70} /* (27, 9, 12) {real, imag} */,
  {32'hc0b69df8, 32'h427e49c6} /* (27, 9, 11) {real, imag} */,
  {32'hc0468c20, 32'hc176d026} /* (27, 9, 10) {real, imag} */,
  {32'hc1c449e6, 32'h422cead6} /* (27, 9, 9) {real, imag} */,
  {32'hc1e4bd9b, 32'hc17c9af6} /* (27, 9, 8) {real, imag} */,
  {32'hc2151514, 32'hc1aacfac} /* (27, 9, 7) {real, imag} */,
  {32'h4190f4b9, 32'hc23af000} /* (27, 9, 6) {real, imag} */,
  {32'h42d34d3c, 32'h42893c01} /* (27, 9, 5) {real, imag} */,
  {32'hc2a38f21, 32'h413768a8} /* (27, 9, 4) {real, imag} */,
  {32'hc1874c51, 32'hc2d960be} /* (27, 9, 3) {real, imag} */,
  {32'hc1b15afe, 32'h4282eec6} /* (27, 9, 2) {real, imag} */,
  {32'h41295400, 32'hbf3b6e40} /* (27, 9, 1) {real, imag} */,
  {32'hc18047cc, 32'h41813c0b} /* (27, 9, 0) {real, imag} */,
  {32'h421afb32, 32'hc344cd78} /* (27, 8, 31) {real, imag} */,
  {32'hc1b265a1, 32'h42aba9de} /* (27, 8, 30) {real, imag} */,
  {32'h4312ab17, 32'h41d46e00} /* (27, 8, 29) {real, imag} */,
  {32'hc2ad7dfc, 32'h428fa744} /* (27, 8, 28) {real, imag} */,
  {32'h42da7af8, 32'hc1d93c40} /* (27, 8, 27) {real, imag} */,
  {32'hc1775a0c, 32'h4243788c} /* (27, 8, 26) {real, imag} */,
  {32'hc0bc94dc, 32'hc20735da} /* (27, 8, 25) {real, imag} */,
  {32'h42d707e1, 32'h42703d62} /* (27, 8, 24) {real, imag} */,
  {32'h4239ac79, 32'h417a644f} /* (27, 8, 23) {real, imag} */,
  {32'hc0e83cc8, 32'h41d6e28c} /* (27, 8, 22) {real, imag} */,
  {32'hbfa7fce0, 32'hc135cbb5} /* (27, 8, 21) {real, imag} */,
  {32'hc2155c5f, 32'hc198f36b} /* (27, 8, 20) {real, imag} */,
  {32'h418b3e10, 32'h4188f1ed} /* (27, 8, 19) {real, imag} */,
  {32'hc0e64d93, 32'hc11a9acb} /* (27, 8, 18) {real, imag} */,
  {32'hc175e20e, 32'h40afdc20} /* (27, 8, 17) {real, imag} */,
  {32'hc1c0bf92, 32'h403b8520} /* (27, 8, 16) {real, imag} */,
  {32'h41da320f, 32'hc1140ed8} /* (27, 8, 15) {real, imag} */,
  {32'hc0063386, 32'hc0d44f1a} /* (27, 8, 14) {real, imag} */,
  {32'h4117b219, 32'hc11df366} /* (27, 8, 13) {real, imag} */,
  {32'h420805b5, 32'hc1f8ee35} /* (27, 8, 12) {real, imag} */,
  {32'h42aa02fa, 32'h41aade94} /* (27, 8, 11) {real, imag} */,
  {32'hc2982b3e, 32'hc281ed6b} /* (27, 8, 10) {real, imag} */,
  {32'hc2078337, 32'hc212c20b} /* (27, 8, 9) {real, imag} */,
  {32'hc20ed91e, 32'h41ac073d} /* (27, 8, 8) {real, imag} */,
  {32'hc288fa1f, 32'h3f76aa20} /* (27, 8, 7) {real, imag} */,
  {32'h429fd6b6, 32'hc2a558ac} /* (27, 8, 6) {real, imag} */,
  {32'hc1fcf01e, 32'hc1918a88} /* (27, 8, 5) {real, imag} */,
  {32'hc27b1a59, 32'hc1d53a1e} /* (27, 8, 4) {real, imag} */,
  {32'hc28c506e, 32'h42b94b86} /* (27, 8, 3) {real, imag} */,
  {32'h4241da96, 32'h4267b0cd} /* (27, 8, 2) {real, imag} */,
  {32'hc0d6d278, 32'hc0c7d1c0} /* (27, 8, 1) {real, imag} */,
  {32'h4153d1f0, 32'hc2da59b5} /* (27, 8, 0) {real, imag} */,
  {32'h414cfe84, 32'hc2a16e56} /* (27, 7, 31) {real, imag} */,
  {32'h43155144, 32'hc1666c74} /* (27, 7, 30) {real, imag} */,
  {32'h4283e204, 32'hc282c90a} /* (27, 7, 29) {real, imag} */,
  {32'hc1a3ad9a, 32'h428afa08} /* (27, 7, 28) {real, imag} */,
  {32'hbe15d280, 32'hc2641f60} /* (27, 7, 27) {real, imag} */,
  {32'hc25bd20e, 32'hc0e0b2d4} /* (27, 7, 26) {real, imag} */,
  {32'hc27efa9a, 32'hc1af7956} /* (27, 7, 25) {real, imag} */,
  {32'h42989889, 32'hc1b52b65} /* (27, 7, 24) {real, imag} */,
  {32'h4197a494, 32'hc1ff7110} /* (27, 7, 23) {real, imag} */,
  {32'hc112b758, 32'h41dd2e79} /* (27, 7, 22) {real, imag} */,
  {32'h4226787a, 32'hc272fb4b} /* (27, 7, 21) {real, imag} */,
  {32'h4210ca0c, 32'h420fe470} /* (27, 7, 20) {real, imag} */,
  {32'hc1a2ced2, 32'h423b36fe} /* (27, 7, 19) {real, imag} */,
  {32'h405966f4, 32'hbe58a300} /* (27, 7, 18) {real, imag} */,
  {32'h3f405320, 32'h420d756f} /* (27, 7, 17) {real, imag} */,
  {32'hc25c2296, 32'h4001b7c0} /* (27, 7, 16) {real, imag} */,
  {32'h41ab41db, 32'h41e7dcb6} /* (27, 7, 15) {real, imag} */,
  {32'h41d18a32, 32'h4198470e} /* (27, 7, 14) {real, imag} */,
  {32'h41a9c2aa, 32'h40443268} /* (27, 7, 13) {real, imag} */,
  {32'h41e09c88, 32'hc1be8ee5} /* (27, 7, 12) {real, imag} */,
  {32'hc1432538, 32'hc2347a9b} /* (27, 7, 11) {real, imag} */,
  {32'hc16c7ef8, 32'hbf2a83a0} /* (27, 7, 10) {real, imag} */,
  {32'h3e1347c0, 32'hc0c16a76} /* (27, 7, 9) {real, imag} */,
  {32'h41f3a273, 32'hc1e7f7f3} /* (27, 7, 8) {real, imag} */,
  {32'hc26e15f0, 32'hc0563b5c} /* (27, 7, 7) {real, imag} */,
  {32'hc2100202, 32'hc1324d8e} /* (27, 7, 6) {real, imag} */,
  {32'h419452b7, 32'h4266e760} /* (27, 7, 5) {real, imag} */,
  {32'h42357c21, 32'hc25c9e4e} /* (27, 7, 4) {real, imag} */,
  {32'h424c9cdc, 32'h429271d6} /* (27, 7, 3) {real, imag} */,
  {32'h430cea6a, 32'hc2b22532} /* (27, 7, 2) {real, imag} */,
  {32'hc228d8b8, 32'h42e6b882} /* (27, 7, 1) {real, imag} */,
  {32'hc25ef592, 32'h42dcaba8} /* (27, 7, 0) {real, imag} */,
  {32'hc31b1ff5, 32'hc2d742e8} /* (27, 6, 31) {real, imag} */,
  {32'hc291e5b2, 32'h4188b289} /* (27, 6, 30) {real, imag} */,
  {32'hc3001eaa, 32'hc13a0ffa} /* (27, 6, 29) {real, imag} */,
  {32'h428f12d2, 32'hc0f2e1c0} /* (27, 6, 28) {real, imag} */,
  {32'h433e7806, 32'h41b52e24} /* (27, 6, 27) {real, imag} */,
  {32'h42a5fd80, 32'h428cebd4} /* (27, 6, 26) {real, imag} */,
  {32'h423342fd, 32'hc2d536d7} /* (27, 6, 25) {real, imag} */,
  {32'hc1cc40c6, 32'hc1ce200e} /* (27, 6, 24) {real, imag} */,
  {32'hc233db96, 32'h3ff336f0} /* (27, 6, 23) {real, imag} */,
  {32'h42b416d6, 32'h41c1a6db} /* (27, 6, 22) {real, imag} */,
  {32'hc1b4fb3c, 32'h40137af0} /* (27, 6, 21) {real, imag} */,
  {32'h41a27b3c, 32'hc0b2fb9f} /* (27, 6, 20) {real, imag} */,
  {32'h41965251, 32'hc192e5e1} /* (27, 6, 19) {real, imag} */,
  {32'hc0e09c94, 32'hc158bb20} /* (27, 6, 18) {real, imag} */,
  {32'hc1c09ee9, 32'hc1e251c1} /* (27, 6, 17) {real, imag} */,
  {32'h41303d9c, 32'hc1384968} /* (27, 6, 16) {real, imag} */,
  {32'h41e4cd49, 32'h41eaf739} /* (27, 6, 15) {real, imag} */,
  {32'hc1743bce, 32'hc253dd84} /* (27, 6, 14) {real, imag} */,
  {32'h3f5b19a0, 32'hc17824da} /* (27, 6, 13) {real, imag} */,
  {32'hc22e00b4, 32'hc19d33f0} /* (27, 6, 12) {real, imag} */,
  {32'h424647ee, 32'h41eca200} /* (27, 6, 11) {real, imag} */,
  {32'hc0c8fbc0, 32'h4194f2e7} /* (27, 6, 10) {real, imag} */,
  {32'hc2c8b871, 32'h40638dc8} /* (27, 6, 9) {real, imag} */,
  {32'h42a86614, 32'h43076c94} /* (27, 6, 8) {real, imag} */,
  {32'hc1fb28aa, 32'hc2879ca7} /* (27, 6, 7) {real, imag} */,
  {32'h4211c384, 32'hc2bf80a0} /* (27, 6, 6) {real, imag} */,
  {32'h41aafabc, 32'hc2e093ed} /* (27, 6, 5) {real, imag} */,
  {32'hc2148a32, 32'hc23693e0} /* (27, 6, 4) {real, imag} */,
  {32'h422ccc02, 32'h42321e9c} /* (27, 6, 3) {real, imag} */,
  {32'h418609e2, 32'h3f1b73a0} /* (27, 6, 2) {real, imag} */,
  {32'hc30a64fb, 32'hc23e21f4} /* (27, 6, 1) {real, imag} */,
  {32'h42004719, 32'hc3166abc} /* (27, 6, 0) {real, imag} */,
  {32'h4287507e, 32'hc331a3aa} /* (27, 5, 31) {real, imag} */,
  {32'h43320891, 32'h4320e1c0} /* (27, 5, 30) {real, imag} */,
  {32'hc3017d2a, 32'h42e33386} /* (27, 5, 29) {real, imag} */,
  {32'hc124d726, 32'h42619df8} /* (27, 5, 28) {real, imag} */,
  {32'h430e3698, 32'hc1c34550} /* (27, 5, 27) {real, imag} */,
  {32'h4222bde3, 32'hc25e7e1c} /* (27, 5, 26) {real, imag} */,
  {32'hc14cdc82, 32'hc2a246dc} /* (27, 5, 25) {real, imag} */,
  {32'hc1c10a2a, 32'hc0660930} /* (27, 5, 24) {real, imag} */,
  {32'hc27b881f, 32'h41e98b43} /* (27, 5, 23) {real, imag} */,
  {32'h4185b29c, 32'h40eab918} /* (27, 5, 22) {real, imag} */,
  {32'h41092884, 32'h4136533a} /* (27, 5, 21) {real, imag} */,
  {32'h420ca000, 32'hc1823d8c} /* (27, 5, 20) {real, imag} */,
  {32'h416b246e, 32'hc0ec4c98} /* (27, 5, 19) {real, imag} */,
  {32'h41e1b198, 32'h4209cec5} /* (27, 5, 18) {real, imag} */,
  {32'h41828b46, 32'h412c13cc} /* (27, 5, 17) {real, imag} */,
  {32'h41f5e250, 32'hc1a4bed0} /* (27, 5, 16) {real, imag} */,
  {32'hc1af52aa, 32'hbf58c7b8} /* (27, 5, 15) {real, imag} */,
  {32'hc212cde6, 32'hc0923948} /* (27, 5, 14) {real, imag} */,
  {32'h4080a13c, 32'h420598ad} /* (27, 5, 13) {real, imag} */,
  {32'h424d52c2, 32'hc28c7dce} /* (27, 5, 12) {real, imag} */,
  {32'h412d6664, 32'h3ce24c00} /* (27, 5, 11) {real, imag} */,
  {32'h423ccd13, 32'h42933232} /* (27, 5, 10) {real, imag} */,
  {32'h41db6c82, 32'h4219163c} /* (27, 5, 9) {real, imag} */,
  {32'hc16f0a8c, 32'hc2c3169a} /* (27, 5, 8) {real, imag} */,
  {32'h42398e6e, 32'hc2591f58} /* (27, 5, 7) {real, imag} */,
  {32'hc1689fc0, 32'h42f63d12} /* (27, 5, 6) {real, imag} */,
  {32'h42755a28, 32'h42c39152} /* (27, 5, 5) {real, imag} */,
  {32'h41097efe, 32'hc1940334} /* (27, 5, 4) {real, imag} */,
  {32'h42137f6a, 32'hc1a86d46} /* (27, 5, 3) {real, imag} */,
  {32'hc1e5a9e8, 32'h4281f73a} /* (27, 5, 2) {real, imag} */,
  {32'hc370a6ff, 32'hc3443386} /* (27, 5, 1) {real, imag} */,
  {32'hc2e78040, 32'hc2838146} /* (27, 5, 0) {real, imag} */,
  {32'hc340c2b3, 32'h42e0cabd} /* (27, 4, 31) {real, imag} */,
  {32'h42d3e678, 32'hc2e34fec} /* (27, 4, 30) {real, imag} */,
  {32'h41d0a523, 32'hc2e9ffbf} /* (27, 4, 29) {real, imag} */,
  {32'hc28147fe, 32'h431dcaba} /* (27, 4, 28) {real, imag} */,
  {32'hc1583ec2, 32'hc2395a6e} /* (27, 4, 27) {real, imag} */,
  {32'hc284d238, 32'hc2934035} /* (27, 4, 26) {real, imag} */,
  {32'h41a06e97, 32'h4297e94a} /* (27, 4, 25) {real, imag} */,
  {32'hc2a70200, 32'hc29b1048} /* (27, 4, 24) {real, imag} */,
  {32'hc1b50152, 32'hc293be70} /* (27, 4, 23) {real, imag} */,
  {32'h4295c1fd, 32'h421efad6} /* (27, 4, 22) {real, imag} */,
  {32'h3f9c7ae0, 32'h40e11ae4} /* (27, 4, 21) {real, imag} */,
  {32'hc1f19ab0, 32'hc18e5bc2} /* (27, 4, 20) {real, imag} */,
  {32'hc140ac96, 32'hc224a900} /* (27, 4, 19) {real, imag} */,
  {32'hc18fdad2, 32'h413d3ee0} /* (27, 4, 18) {real, imag} */,
  {32'h422a10e8, 32'hbf456600} /* (27, 4, 17) {real, imag} */,
  {32'h416e2d9c, 32'h42218666} /* (27, 4, 16) {real, imag} */,
  {32'hc1868660, 32'hc2192c00} /* (27, 4, 15) {real, imag} */,
  {32'hc106e7ac, 32'hc25f0068} /* (27, 4, 14) {real, imag} */,
  {32'h4180a853, 32'h3f9a40c0} /* (27, 4, 13) {real, imag} */,
  {32'h3f8e2ab8, 32'h41c2fdfe} /* (27, 4, 12) {real, imag} */,
  {32'hc218b2ea, 32'h41df2051} /* (27, 4, 11) {real, imag} */,
  {32'hc27de46e, 32'hbfe13490} /* (27, 4, 10) {real, imag} */,
  {32'h42815194, 32'h4215cf26} /* (27, 4, 9) {real, imag} */,
  {32'h4167d100, 32'h41e6e4c5} /* (27, 4, 8) {real, imag} */,
  {32'h41b9f53d, 32'hbf9ca760} /* (27, 4, 7) {real, imag} */,
  {32'h418a7d73, 32'h431bf20a} /* (27, 4, 6) {real, imag} */,
  {32'h426b421c, 32'hc2688192} /* (27, 4, 5) {real, imag} */,
  {32'hc0baa148, 32'h421eed78} /* (27, 4, 4) {real, imag} */,
  {32'hc238f45e, 32'hc2b3c671} /* (27, 4, 3) {real, imag} */,
  {32'hc303df64, 32'hc353003e} /* (27, 4, 2) {real, imag} */,
  {32'hc0151840, 32'h438f4d38} /* (27, 4, 1) {real, imag} */,
  {32'h427d5679, 32'hc306af4e} /* (27, 4, 0) {real, imag} */,
  {32'hc3955e5a, 32'hc27a46da} /* (27, 3, 31) {real, imag} */,
  {32'h4360a5ef, 32'h42dad565} /* (27, 3, 30) {real, imag} */,
  {32'h428aff1e, 32'hc20bd3f9} /* (27, 3, 29) {real, imag} */,
  {32'h42d843f7, 32'h42ed8a2c} /* (27, 3, 28) {real, imag} */,
  {32'hc2b02f43, 32'hc2fb630f} /* (27, 3, 27) {real, imag} */,
  {32'hc2c7d4fa, 32'h4228472c} /* (27, 3, 26) {real, imag} */,
  {32'h422d30ba, 32'hc289c2c6} /* (27, 3, 25) {real, imag} */,
  {32'h42b3bb84, 32'hc31b80f4} /* (27, 3, 24) {real, imag} */,
  {32'h42bd1a46, 32'h416c2044} /* (27, 3, 23) {real, imag} */,
  {32'hc2b74aa4, 32'h42390bd8} /* (27, 3, 22) {real, imag} */,
  {32'h4029f148, 32'h418cdc68} /* (27, 3, 21) {real, imag} */,
  {32'hc22dbb70, 32'hc1491614} /* (27, 3, 20) {real, imag} */,
  {32'h41ef00fc, 32'h42253cf1} /* (27, 3, 19) {real, imag} */,
  {32'h4226dc80, 32'hc1cd5ace} /* (27, 3, 18) {real, imag} */,
  {32'h42084600, 32'h4106d35a} /* (27, 3, 17) {real, imag} */,
  {32'hc1534500, 32'h41918a8c} /* (27, 3, 16) {real, imag} */,
  {32'hc1e977a0, 32'hc1d2c9a3} /* (27, 3, 15) {real, imag} */,
  {32'hc21daa88, 32'hc197254e} /* (27, 3, 14) {real, imag} */,
  {32'hbffe7aa8, 32'hc20399d5} /* (27, 3, 13) {real, imag} */,
  {32'h41ebc1b8, 32'h42a6b640} /* (27, 3, 12) {real, imag} */,
  {32'h410fe4d6, 32'h41a07a6c} /* (27, 3, 11) {real, imag} */,
  {32'hc20024a7, 32'hc1a5c3f5} /* (27, 3, 10) {real, imag} */,
  {32'hc0f7ada0, 32'hc2da3f0a} /* (27, 3, 9) {real, imag} */,
  {32'hc24aef9c, 32'hc28d20bb} /* (27, 3, 8) {real, imag} */,
  {32'hc28990cb, 32'h43205fca} /* (27, 3, 7) {real, imag} */,
  {32'h43047121, 32'hc30d7ca5} /* (27, 3, 6) {real, imag} */,
  {32'hc1167d68, 32'h42c09aa1} /* (27, 3, 5) {real, imag} */,
  {32'hc2a78ec3, 32'h418d736a} /* (27, 3, 4) {real, imag} */,
  {32'h41262e60, 32'hc109d284} /* (27, 3, 3) {real, imag} */,
  {32'h43001353, 32'hc2cf5c0d} /* (27, 3, 2) {real, imag} */,
  {32'hc28aed16, 32'h42f8f5f3} /* (27, 3, 1) {real, imag} */,
  {32'h42fe71f2, 32'h43127e04} /* (27, 3, 0) {real, imag} */,
  {32'hc3c6580c, 32'hc3eb8fac} /* (27, 2, 31) {real, imag} */,
  {32'h433bdbe6, 32'h4387a5d4} /* (27, 2, 30) {real, imag} */,
  {32'hc33ce760, 32'hc306cc46} /* (27, 2, 29) {real, imag} */,
  {32'hc336f44c, 32'hc1fb52a2} /* (27, 2, 28) {real, imag} */,
  {32'h4288c4be, 32'h41ec2dfc} /* (27, 2, 27) {real, imag} */,
  {32'h43249a2a, 32'h41cc0767} /* (27, 2, 26) {real, imag} */,
  {32'hc32af61c, 32'h42353dbc} /* (27, 2, 25) {real, imag} */,
  {32'h43056d15, 32'hbfd109a0} /* (27, 2, 24) {real, imag} */,
  {32'h42d92ae5, 32'hc28c3b64} /* (27, 2, 23) {real, imag} */,
  {32'h41beff79, 32'hc0ce1330} /* (27, 2, 22) {real, imag} */,
  {32'h420f8866, 32'hc2516900} /* (27, 2, 21) {real, imag} */,
  {32'h419586b6, 32'h4088a9b8} /* (27, 2, 20) {real, imag} */,
  {32'h40ce7328, 32'hc21a37aa} /* (27, 2, 19) {real, imag} */,
  {32'h4192076e, 32'hc211aaf4} /* (27, 2, 18) {real, imag} */,
  {32'hc1822974, 32'h4216859a} /* (27, 2, 17) {real, imag} */,
  {32'h412b3344, 32'hc1abb700} /* (27, 2, 16) {real, imag} */,
  {32'h415a2988, 32'hc0cdeed0} /* (27, 2, 15) {real, imag} */,
  {32'h423f1e55, 32'h4249b884} /* (27, 2, 14) {real, imag} */,
  {32'hc201a987, 32'h409c07dc} /* (27, 2, 13) {real, imag} */,
  {32'hbfb35b20, 32'hc1822f56} /* (27, 2, 12) {real, imag} */,
  {32'hc101b790, 32'hbff7e270} /* (27, 2, 11) {real, imag} */,
  {32'h42017588, 32'hc1ca96e2} /* (27, 2, 10) {real, imag} */,
  {32'hc224c0fa, 32'hc1e36db2} /* (27, 2, 9) {real, imag} */,
  {32'h417951a0, 32'hc29701fa} /* (27, 2, 8) {real, imag} */,
  {32'hc2904ed7, 32'hc245db4a} /* (27, 2, 7) {real, imag} */,
  {32'h42ae94ba, 32'hc29f0c2a} /* (27, 2, 6) {real, imag} */,
  {32'hc2aa3c02, 32'h43342666} /* (27, 2, 5) {real, imag} */,
  {32'hc25c2912, 32'hc3036a50} /* (27, 2, 4) {real, imag} */,
  {32'h41415538, 32'h418b3b8a} /* (27, 2, 3) {real, imag} */,
  {32'h436d2e56, 32'h43bd57a2} /* (27, 2, 2) {real, imag} */,
  {32'hc32cca40, 32'hc3adf63e} /* (27, 2, 1) {real, imag} */,
  {32'h42a57824, 32'hc3f147f2} /* (27, 2, 0) {real, imag} */,
  {32'h43f060e9, 32'h439f2673} /* (27, 1, 31) {real, imag} */,
  {32'hc3086fde, 32'hc30a2284} /* (27, 1, 30) {real, imag} */,
  {32'h425d397e, 32'h422007ea} /* (27, 1, 29) {real, imag} */,
  {32'h42dde68b, 32'h4095fb40} /* (27, 1, 28) {real, imag} */,
  {32'hc3744681, 32'hc3074182} /* (27, 1, 27) {real, imag} */,
  {32'hc2378eed, 32'hbc58d600} /* (27, 1, 26) {real, imag} */,
  {32'hc1813d64, 32'h433d4310} /* (27, 1, 25) {real, imag} */,
  {32'hc2d25e04, 32'hc25e7b18} /* (27, 1, 24) {real, imag} */,
  {32'hc19226db, 32'h409ae570} /* (27, 1, 23) {real, imag} */,
  {32'h418fc7e6, 32'h4117f8aa} /* (27, 1, 22) {real, imag} */,
  {32'hc209fb35, 32'hc099c858} /* (27, 1, 21) {real, imag} */,
  {32'hc174d0bc, 32'h424da9c6} /* (27, 1, 20) {real, imag} */,
  {32'h41252162, 32'hc1403bb0} /* (27, 1, 19) {real, imag} */,
  {32'h408597ac, 32'hc216732a} /* (27, 1, 18) {real, imag} */,
  {32'h40820010, 32'hc1f3b11c} /* (27, 1, 17) {real, imag} */,
  {32'h41bd6c58, 32'h4120dca0} /* (27, 1, 16) {real, imag} */,
  {32'hc1a7155c, 32'hc22e4da2} /* (27, 1, 15) {real, imag} */,
  {32'h420f734e, 32'h4264c6da} /* (27, 1, 14) {real, imag} */,
  {32'h421604a0, 32'h42159cdc} /* (27, 1, 13) {real, imag} */,
  {32'h41810b3e, 32'h4173e7e0} /* (27, 1, 12) {real, imag} */,
  {32'hc11f606c, 32'hc28f8c80} /* (27, 1, 11) {real, imag} */,
  {32'h40b726d6, 32'hc1082ca2} /* (27, 1, 10) {real, imag} */,
  {32'hc1b1b013, 32'hc250c456} /* (27, 1, 9) {real, imag} */,
  {32'h420257e9, 32'hc34eb418} /* (27, 1, 8) {real, imag} */,
  {32'h42bb9bb1, 32'h42e08685} /* (27, 1, 7) {real, imag} */,
  {32'h42b75f92, 32'hc01f574a} /* (27, 1, 6) {real, imag} */,
  {32'hc21abb4c, 32'hc26dbd5b} /* (27, 1, 5) {real, imag} */,
  {32'hc1fcd254, 32'h42b1f187} /* (27, 1, 4) {real, imag} */,
  {32'hbf7aaca0, 32'hc362b010} /* (27, 1, 3) {real, imag} */,
  {32'h43403fe4, 32'hc3bd6940} /* (27, 1, 2) {real, imag} */,
  {32'h416c05a0, 32'h441e81ae} /* (27, 1, 1) {real, imag} */,
  {32'h4324ff25, 32'h4405c81c} /* (27, 1, 0) {real, imag} */,
  {32'h43cd35fa, 32'h427b25ec} /* (27, 0, 31) {real, imag} */,
  {32'hc376bdef, 32'hc2a54a12} /* (27, 0, 30) {real, imag} */,
  {32'h423d9aa1, 32'hc2fd8eae} /* (27, 0, 29) {real, imag} */,
  {32'h419d89bd, 32'hc10c4644} /* (27, 0, 28) {real, imag} */,
  {32'h42245372, 32'hc1c9b2ec} /* (27, 0, 27) {real, imag} */,
  {32'h42663ac0, 32'hc1cc8226} /* (27, 0, 26) {real, imag} */,
  {32'hc23e221a, 32'hc2357c78} /* (27, 0, 25) {real, imag} */,
  {32'hc2cd4224, 32'hc2687d7e} /* (27, 0, 24) {real, imag} */,
  {32'hc256ff66, 32'h4212a288} /* (27, 0, 23) {real, imag} */,
  {32'hc2b985ef, 32'hc0d78f7a} /* (27, 0, 22) {real, imag} */,
  {32'hc1beab88, 32'h41804f14} /* (27, 0, 21) {real, imag} */,
  {32'h4202f33e, 32'h4282a394} /* (27, 0, 20) {real, imag} */,
  {32'h42541543, 32'h42444b02} /* (27, 0, 19) {real, imag} */,
  {32'hc18c9a99, 32'hc20cd645} /* (27, 0, 18) {real, imag} */,
  {32'hc0623a20, 32'hc111a210} /* (27, 0, 17) {real, imag} */,
  {32'h427b7f55, 32'h41885630} /* (27, 0, 16) {real, imag} */,
  {32'hc01bd8e0, 32'hc1e37448} /* (27, 0, 15) {real, imag} */,
  {32'h426e4290, 32'hc105bb2c} /* (27, 0, 14) {real, imag} */,
  {32'h40e02348, 32'hc1f92c35} /* (27, 0, 13) {real, imag} */,
  {32'hc0befcdc, 32'h42b51744} /* (27, 0, 12) {real, imag} */,
  {32'hc09fb744, 32'hc281ea35} /* (27, 0, 11) {real, imag} */,
  {32'hc2a21d07, 32'h41bbd486} /* (27, 0, 10) {real, imag} */,
  {32'hc2e3fe1f, 32'h411c4a18} /* (27, 0, 9) {real, imag} */,
  {32'h41ca093e, 32'h43193bac} /* (27, 0, 8) {real, imag} */,
  {32'hc2289cf2, 32'h4276fb3e} /* (27, 0, 7) {real, imag} */,
  {32'hc25651e8, 32'h41fc5ebe} /* (27, 0, 6) {real, imag} */,
  {32'h412ecb27, 32'hc34b0f12} /* (27, 0, 5) {real, imag} */,
  {32'h41b36217, 32'hc302e6d2} /* (27, 0, 4) {real, imag} */,
  {32'hc2c82050, 32'h4212d538} /* (27, 0, 3) {real, imag} */,
  {32'h42a3fd42, 32'hc3082617} /* (27, 0, 2) {real, imag} */,
  {32'h40cbd800, 32'h43ec2d52} /* (27, 0, 1) {real, imag} */,
  {32'h42339501, 32'h43abdc1f} /* (27, 0, 0) {real, imag} */,
  {32'h4260623a, 32'hc2447569} /* (26, 31, 31) {real, imag} */,
  {32'hc2e3f0d6, 32'hc2191e73} /* (26, 31, 30) {real, imag} */,
  {32'hc225668a, 32'hc21376d9} /* (26, 31, 29) {real, imag} */,
  {32'h42aff948, 32'hc13c3748} /* (26, 31, 28) {real, imag} */,
  {32'h422c7d79, 32'hc1aff4bb} /* (26, 31, 27) {real, imag} */,
  {32'hc23c03d2, 32'h41e5cf5e} /* (26, 31, 26) {real, imag} */,
  {32'hc272f64e, 32'h416471c2} /* (26, 31, 25) {real, imag} */,
  {32'hc2416d4a, 32'hc0475e70} /* (26, 31, 24) {real, imag} */,
  {32'h3fe99ca0, 32'hc0d8961c} /* (26, 31, 23) {real, imag} */,
  {32'hc11ca024, 32'h4198d40c} /* (26, 31, 22) {real, imag} */,
  {32'hc215eb68, 32'hc1befa81} /* (26, 31, 21) {real, imag} */,
  {32'hc21d42c4, 32'h42007c40} /* (26, 31, 20) {real, imag} */,
  {32'hc1bde8de, 32'hc2bb54ba} /* (26, 31, 19) {real, imag} */,
  {32'h3ff499c0, 32'h428fe486} /* (26, 31, 18) {real, imag} */,
  {32'h41921392, 32'hc14ed93d} /* (26, 31, 17) {real, imag} */,
  {32'hc1d5eaa0, 32'hbdaa9600} /* (26, 31, 16) {real, imag} */,
  {32'h418658ec, 32'hc1098775} /* (26, 31, 15) {real, imag} */,
  {32'h42852a29, 32'hc1771c68} /* (26, 31, 14) {real, imag} */,
  {32'hc155981d, 32'hc18289aa} /* (26, 31, 13) {real, imag} */,
  {32'h42311a0c, 32'hc297b78c} /* (26, 31, 12) {real, imag} */,
  {32'hc26d79a0, 32'hc102faf6} /* (26, 31, 11) {real, imag} */,
  {32'h42aad628, 32'hc1caea08} /* (26, 31, 10) {real, imag} */,
  {32'hc2917c3c, 32'h42853760} /* (26, 31, 9) {real, imag} */,
  {32'hc009d408, 32'h42d2c038} /* (26, 31, 8) {real, imag} */,
  {32'hc1eef420, 32'h40a76024} /* (26, 31, 7) {real, imag} */,
  {32'h42933236, 32'h4249d34d} /* (26, 31, 6) {real, imag} */,
  {32'h417a47fd, 32'h41110fbe} /* (26, 31, 5) {real, imag} */,
  {32'h42f408bc, 32'hc2e1420f} /* (26, 31, 4) {real, imag} */,
  {32'hc214c978, 32'h42eb21c4} /* (26, 31, 3) {real, imag} */,
  {32'hc1e23970, 32'h426c1f83} /* (26, 31, 2) {real, imag} */,
  {32'hc23ff09e, 32'h422c33c1} /* (26, 31, 1) {real, imag} */,
  {32'h43122fee, 32'h42e849be} /* (26, 31, 0) {real, imag} */,
  {32'hc2d26b99, 32'hc23c7acf} /* (26, 30, 31) {real, imag} */,
  {32'hc26c4dd5, 32'h42d1db66} /* (26, 30, 30) {real, imag} */,
  {32'h42dac500, 32'h42e76ad3} /* (26, 30, 29) {real, imag} */,
  {32'h419e7310, 32'hc29ee298} /* (26, 30, 28) {real, imag} */,
  {32'hc2cfb777, 32'hc28e1df0} /* (26, 30, 27) {real, imag} */,
  {32'h4281c4de, 32'hc28a2b50} /* (26, 30, 26) {real, imag} */,
  {32'hc27dec04, 32'hc292f83c} /* (26, 30, 25) {real, imag} */,
  {32'h42977da9, 32'hc2246654} /* (26, 30, 24) {real, imag} */,
  {32'hc2531c96, 32'h3f3db9c0} /* (26, 30, 23) {real, imag} */,
  {32'hc18f947c, 32'h41a6a17d} /* (26, 30, 22) {real, imag} */,
  {32'hbfb02790, 32'hc136d754} /* (26, 30, 21) {real, imag} */,
  {32'hc1d0bde6, 32'hc23891a2} /* (26, 30, 20) {real, imag} */,
  {32'hc0e98a01, 32'hc16e7bac} /* (26, 30, 19) {real, imag} */,
  {32'h40429c24, 32'h41eb8254} /* (26, 30, 18) {real, imag} */,
  {32'h3f8cde40, 32'hc16c059f} /* (26, 30, 17) {real, imag} */,
  {32'h41411802, 32'hc172c070} /* (26, 30, 16) {real, imag} */,
  {32'h413eaec8, 32'h4018e8bc} /* (26, 30, 15) {real, imag} */,
  {32'hc08c10ae, 32'hc101c624} /* (26, 30, 14) {real, imag} */,
  {32'h418ed2f0, 32'h413ae314} /* (26, 30, 13) {real, imag} */,
  {32'h40c59928, 32'hc22d6ecc} /* (26, 30, 12) {real, imag} */,
  {32'hc18c666b, 32'h4291750e} /* (26, 30, 11) {real, imag} */,
  {32'h3f906708, 32'h4284a5ad} /* (26, 30, 10) {real, imag} */,
  {32'hc0ec1490, 32'hc2b8577a} /* (26, 30, 9) {real, imag} */,
  {32'hc2e3ccfb, 32'hc2ccca32} /* (26, 30, 8) {real, imag} */,
  {32'h42f2b610, 32'h4196b6aa} /* (26, 30, 7) {real, imag} */,
  {32'hc2b5e7be, 32'hc16ad552} /* (26, 30, 6) {real, imag} */,
  {32'hc25ee3ba, 32'hc2afa5e0} /* (26, 30, 5) {real, imag} */,
  {32'hc2c387e4, 32'h4316fa48} /* (26, 30, 4) {real, imag} */,
  {32'hc2d45f46, 32'h41d27284} /* (26, 30, 3) {real, imag} */,
  {32'h42540cc7, 32'h41ab0530} /* (26, 30, 2) {real, imag} */,
  {32'h43af149e, 32'hc18bba5a} /* (26, 30, 1) {real, imag} */,
  {32'hc28e0b78, 32'h43175ed3} /* (26, 30, 0) {real, imag} */,
  {32'h42ebc970, 32'h42e98624} /* (26, 29, 31) {real, imag} */,
  {32'h42c676c8, 32'hc0af4f60} /* (26, 29, 30) {real, imag} */,
  {32'hc309090d, 32'hc290bfdc} /* (26, 29, 29) {real, imag} */,
  {32'h426b347c, 32'h419a20dd} /* (26, 29, 28) {real, imag} */,
  {32'h41ac4fd3, 32'h432ebce2} /* (26, 29, 27) {real, imag} */,
  {32'hc22e6112, 32'hc1690934} /* (26, 29, 26) {real, imag} */,
  {32'hc213abc2, 32'h41b5b836} /* (26, 29, 25) {real, imag} */,
  {32'hc213ab2a, 32'h41166848} /* (26, 29, 24) {real, imag} */,
  {32'hc1a38678, 32'h418d467b} /* (26, 29, 23) {real, imag} */,
  {32'hbfdc4f5c, 32'h41619944} /* (26, 29, 22) {real, imag} */,
  {32'hbfb72950, 32'h4229f424} /* (26, 29, 21) {real, imag} */,
  {32'hc226fb8c, 32'h411103da} /* (26, 29, 20) {real, imag} */,
  {32'h40082330, 32'h416df6fa} /* (26, 29, 19) {real, imag} */,
  {32'h41682d7a, 32'h4261ff0e} /* (26, 29, 18) {real, imag} */,
  {32'hbf3e6df0, 32'hc1869516} /* (26, 29, 17) {real, imag} */,
  {32'h4229e246, 32'hc1ec15e5} /* (26, 29, 16) {real, imag} */,
  {32'h4111c86f, 32'hc1a6aac6} /* (26, 29, 15) {real, imag} */,
  {32'hc013fb68, 32'h41eb94bd} /* (26, 29, 14) {real, imag} */,
  {32'h41fcfa3e, 32'hc1075b22} /* (26, 29, 13) {real, imag} */,
  {32'hc20db5dc, 32'hc140d1e4} /* (26, 29, 12) {real, imag} */,
  {32'h423e5436, 32'hc2db04fa} /* (26, 29, 11) {real, imag} */,
  {32'h41228590, 32'h42c42d18} /* (26, 29, 10) {real, imag} */,
  {32'h420fba3e, 32'h42833de6} /* (26, 29, 9) {real, imag} */,
  {32'h411356de, 32'h4061f910} /* (26, 29, 8) {real, imag} */,
  {32'h41017fc0, 32'h42c1df84} /* (26, 29, 7) {real, imag} */,
  {32'h420c531e, 32'hc2a6fc22} /* (26, 29, 6) {real, imag} */,
  {32'hc0f58ca4, 32'h421440b0} /* (26, 29, 5) {real, imag} */,
  {32'h41c9e5ff, 32'hc218fe28} /* (26, 29, 4) {real, imag} */,
  {32'h41b41e92, 32'hc1e243ef} /* (26, 29, 3) {real, imag} */,
  {32'h428e4d50, 32'h428bd5e0} /* (26, 29, 2) {real, imag} */,
  {32'h42444c7b, 32'hc3237084} /* (26, 29, 1) {real, imag} */,
  {32'hc229a806, 32'hc2b0b47b} /* (26, 29, 0) {real, imag} */,
  {32'h42dd784e, 32'hc2254986} /* (26, 28, 31) {real, imag} */,
  {32'hc22ac43d, 32'hc2579d14} /* (26, 28, 30) {real, imag} */,
  {32'hc2ab4e68, 32'h4331afff} /* (26, 28, 29) {real, imag} */,
  {32'h4239e960, 32'h428ea0ea} /* (26, 28, 28) {real, imag} */,
  {32'h41c54052, 32'hc25d93d8} /* (26, 28, 27) {real, imag} */,
  {32'h41eac780, 32'h4241e630} /* (26, 28, 26) {real, imag} */,
  {32'hc2a0f24e, 32'h40079110} /* (26, 28, 25) {real, imag} */,
  {32'hc285cb5a, 32'hc11fda22} /* (26, 28, 24) {real, imag} */,
  {32'hc2e5606c, 32'hc257b180} /* (26, 28, 23) {real, imag} */,
  {32'h42589a55, 32'h419d4a88} /* (26, 28, 22) {real, imag} */,
  {32'h421351d7, 32'hc1423576} /* (26, 28, 21) {real, imag} */,
  {32'hc1b8ec48, 32'hc0808ce2} /* (26, 28, 20) {real, imag} */,
  {32'hc1075ba6, 32'h41064e4a} /* (26, 28, 19) {real, imag} */,
  {32'hbf7ce080, 32'hc0174f28} /* (26, 28, 18) {real, imag} */,
  {32'h40e169d4, 32'hc1404662} /* (26, 28, 17) {real, imag} */,
  {32'h41108dc0, 32'h41db0863} /* (26, 28, 16) {real, imag} */,
  {32'hc2155fae, 32'h3f766520} /* (26, 28, 15) {real, imag} */,
  {32'h40678628, 32'h405f3918} /* (26, 28, 14) {real, imag} */,
  {32'h41ced14d, 32'hc24b17da} /* (26, 28, 13) {real, imag} */,
  {32'h42407ba0, 32'hc17f1209} /* (26, 28, 12) {real, imag} */,
  {32'hc2627cc5, 32'hc1c72b6d} /* (26, 28, 11) {real, imag} */,
  {32'h4263207f, 32'hc2376048} /* (26, 28, 10) {real, imag} */,
  {32'hc23c6664, 32'hc2c2c2ea} /* (26, 28, 9) {real, imag} */,
  {32'h420ce118, 32'h420b9304} /* (26, 28, 8) {real, imag} */,
  {32'hc2b623b0, 32'hc20b8f0c} /* (26, 28, 7) {real, imag} */,
  {32'hbf4ce240, 32'h42f7e02a} /* (26, 28, 6) {real, imag} */,
  {32'h4268e591, 32'h4277ea18} /* (26, 28, 5) {real, imag} */,
  {32'hc30159db, 32'hc2efa052} /* (26, 28, 4) {real, imag} */,
  {32'h419294a8, 32'h432c0177} /* (26, 28, 3) {real, imag} */,
  {32'h400b7010, 32'h4162b146} /* (26, 28, 2) {real, imag} */,
  {32'h40877600, 32'hc2b81bc7} /* (26, 28, 1) {real, imag} */,
  {32'h42c38022, 32'h4228419a} /* (26, 28, 0) {real, imag} */,
  {32'h42bfeb8f, 32'h42c29cdf} /* (26, 27, 31) {real, imag} */,
  {32'hc2205d04, 32'h42e86110} /* (26, 27, 30) {real, imag} */,
  {32'hc16481e8, 32'hbf9b7420} /* (26, 27, 29) {real, imag} */,
  {32'h426788e6, 32'hc2290fe2} /* (26, 27, 28) {real, imag} */,
  {32'h41bd86ff, 32'h41b4abe6} /* (26, 27, 27) {real, imag} */,
  {32'h41d6b857, 32'h4073f814} /* (26, 27, 26) {real, imag} */,
  {32'h4243dd9d, 32'hc2f12435} /* (26, 27, 25) {real, imag} */,
  {32'hc1d8e977, 32'h411c1c3a} /* (26, 27, 24) {real, imag} */,
  {32'hc111ca10, 32'h42cff635} /* (26, 27, 23) {real, imag} */,
  {32'hc292584a, 32'hc2295872} /* (26, 27, 22) {real, imag} */,
  {32'h421beab1, 32'hc10ebf72} /* (26, 27, 21) {real, imag} */,
  {32'hc286df67, 32'h409dfbb8} /* (26, 27, 20) {real, imag} */,
  {32'h4234c79a, 32'hc18db1dc} /* (26, 27, 19) {real, imag} */,
  {32'h40676b38, 32'hc1756850} /* (26, 27, 18) {real, imag} */,
  {32'hbe433100, 32'hc20c8df0} /* (26, 27, 17) {real, imag} */,
  {32'hc26ffccb, 32'h41c2e535} /* (26, 27, 16) {real, imag} */,
  {32'hc0e1bfd8, 32'h4227a95c} /* (26, 27, 15) {real, imag} */,
  {32'h41ad58d7, 32'h40a0a990} /* (26, 27, 14) {real, imag} */,
  {32'h3f90d150, 32'h41532609} /* (26, 27, 13) {real, imag} */,
  {32'h41de92dd, 32'h422aa107} /* (26, 27, 12) {real, imag} */,
  {32'hc261e69f, 32'h4283a256} /* (26, 27, 11) {real, imag} */,
  {32'h3de72a00, 32'h420ca8f0} /* (26, 27, 10) {real, imag} */,
  {32'hc1efff84, 32'h42628746} /* (26, 27, 9) {real, imag} */,
  {32'hc2a7d867, 32'h41f1c5a1} /* (26, 27, 8) {real, imag} */,
  {32'hc2402c61, 32'h422441e6} /* (26, 27, 7) {real, imag} */,
  {32'hc242ce9a, 32'hc0e1a486} /* (26, 27, 6) {real, imag} */,
  {32'h42087ace, 32'h42761671} /* (26, 27, 5) {real, imag} */,
  {32'h40b6f10c, 32'hc35146d2} /* (26, 27, 4) {real, imag} */,
  {32'hc3163404, 32'hc28809c8} /* (26, 27, 3) {real, imag} */,
  {32'h42e9e222, 32'hc0514020} /* (26, 27, 2) {real, imag} */,
  {32'h419b29a8, 32'hc2098b82} /* (26, 27, 1) {real, imag} */,
  {32'hc308eb55, 32'hc26885aa} /* (26, 27, 0) {real, imag} */,
  {32'h42119b48, 32'hc25bc8d4} /* (26, 26, 31) {real, imag} */,
  {32'h41a51704, 32'hc244e8b0} /* (26, 26, 30) {real, imag} */,
  {32'h41c53223, 32'h429e151c} /* (26, 26, 29) {real, imag} */,
  {32'hc25df43e, 32'h4286c054} /* (26, 26, 28) {real, imag} */,
  {32'hc2064e81, 32'hc30739f8} /* (26, 26, 27) {real, imag} */,
  {32'hc1c30c06, 32'hc2237c70} /* (26, 26, 26) {real, imag} */,
  {32'h42670961, 32'h43316e6d} /* (26, 26, 25) {real, imag} */,
  {32'hc28999fc, 32'h41fbfb56} /* (26, 26, 24) {real, imag} */,
  {32'h42721b14, 32'h42389764} /* (26, 26, 23) {real, imag} */,
  {32'hc2c0e773, 32'hc2b2d320} /* (26, 26, 22) {real, imag} */,
  {32'hc200b5e7, 32'hc09115e6} /* (26, 26, 21) {real, imag} */,
  {32'h404a72c8, 32'h414adc4e} /* (26, 26, 20) {real, imag} */,
  {32'h41c476bf, 32'h40abd580} /* (26, 26, 19) {real, imag} */,
  {32'hc145f0fe, 32'hc14faf9a} /* (26, 26, 18) {real, imag} */,
  {32'hc1a07e4b, 32'hc199a21e} /* (26, 26, 17) {real, imag} */,
  {32'hc0996ee0, 32'hc22c2606} /* (26, 26, 16) {real, imag} */,
  {32'h41c2e145, 32'h412ec0c0} /* (26, 26, 15) {real, imag} */,
  {32'hc1120dce, 32'hc2533594} /* (26, 26, 14) {real, imag} */,
  {32'hc07265a8, 32'h41fae874} /* (26, 26, 13) {real, imag} */,
  {32'hc225396a, 32'h4280809e} /* (26, 26, 12) {real, imag} */,
  {32'h41f15bd2, 32'hc1cd33ca} /* (26, 26, 11) {real, imag} */,
  {32'h4092b110, 32'hc0cef738} /* (26, 26, 10) {real, imag} */,
  {32'hc2ab5b8e, 32'hc173e778} /* (26, 26, 9) {real, imag} */,
  {32'h41db0eba, 32'hc0cc79b8} /* (26, 26, 8) {real, imag} */,
  {32'h4256737f, 32'h4227b29c} /* (26, 26, 7) {real, imag} */,
  {32'h417aa350, 32'h41c292ad} /* (26, 26, 6) {real, imag} */,
  {32'h4284b822, 32'h429f5801} /* (26, 26, 5) {real, imag} */,
  {32'h42846d7f, 32'hc2c51222} /* (26, 26, 4) {real, imag} */,
  {32'h424b6a2e, 32'h41a44e2e} /* (26, 26, 3) {real, imag} */,
  {32'hc31e4a78, 32'h42893876} /* (26, 26, 2) {real, imag} */,
  {32'hc1c9df17, 32'h41c353d1} /* (26, 26, 1) {real, imag} */,
  {32'hc1828be5, 32'h42b96d73} /* (26, 26, 0) {real, imag} */,
  {32'h4187725e, 32'h423f52d4} /* (26, 25, 31) {real, imag} */,
  {32'hc2ca080a, 32'hc26d98b9} /* (26, 25, 30) {real, imag} */,
  {32'h432ff37a, 32'hc2361c5c} /* (26, 25, 29) {real, imag} */,
  {32'h433eb0f2, 32'h420df073} /* (26, 25, 28) {real, imag} */,
  {32'hc27779f8, 32'hc1455fbc} /* (26, 25, 27) {real, imag} */,
  {32'h40e5318c, 32'hc1bd8107} /* (26, 25, 26) {real, imag} */,
  {32'hc04c7820, 32'hc0087100} /* (26, 25, 25) {real, imag} */,
  {32'hc225dd62, 32'h41ec1a9a} /* (26, 25, 24) {real, imag} */,
  {32'h4248c47a, 32'h411b41a6} /* (26, 25, 23) {real, imag} */,
  {32'h4280c76a, 32'h421d68fa} /* (26, 25, 22) {real, imag} */,
  {32'hc23d20d2, 32'h40a3589c} /* (26, 25, 21) {real, imag} */,
  {32'hc215ec18, 32'h41a3238c} /* (26, 25, 20) {real, imag} */,
  {32'hc203ed54, 32'hbf8fa970} /* (26, 25, 19) {real, imag} */,
  {32'hc1c1ffa4, 32'h41e6e782} /* (26, 25, 18) {real, imag} */,
  {32'hc2087cb6, 32'h41f5cd3d} /* (26, 25, 17) {real, imag} */,
  {32'h41816112, 32'hc1c87ed0} /* (26, 25, 16) {real, imag} */,
  {32'hc256b416, 32'hc14376de} /* (26, 25, 15) {real, imag} */,
  {32'hbf75e780, 32'hc019ccb0} /* (26, 25, 14) {real, imag} */,
  {32'h414c7fd2, 32'hc14fb80a} /* (26, 25, 13) {real, imag} */,
  {32'hc1cb8e45, 32'h4192904e} /* (26, 25, 12) {real, imag} */,
  {32'h429055bf, 32'h4149890a} /* (26, 25, 11) {real, imag} */,
  {32'h42170309, 32'hc0a8f324} /* (26, 25, 10) {real, imag} */,
  {32'hc21eae62, 32'h40b2f81c} /* (26, 25, 9) {real, imag} */,
  {32'hc240aa32, 32'hc0293890} /* (26, 25, 8) {real, imag} */,
  {32'h42f3d8ad, 32'h4188ff2c} /* (26, 25, 7) {real, imag} */,
  {32'h412ec9ee, 32'hc2aab129} /* (26, 25, 6) {real, imag} */,
  {32'hc2875496, 32'h42941e70} /* (26, 25, 5) {real, imag} */,
  {32'h42bfbf37, 32'h41870928} /* (26, 25, 4) {real, imag} */,
  {32'h425040b6, 32'hc269904e} /* (26, 25, 3) {real, imag} */,
  {32'h42d2b656, 32'h430fa3e3} /* (26, 25, 2) {real, imag} */,
  {32'h42284d05, 32'hc319927f} /* (26, 25, 1) {real, imag} */,
  {32'hc27e4799, 32'h4320e77e} /* (26, 25, 0) {real, imag} */,
  {32'hc214e660, 32'hc2d48b86} /* (26, 24, 31) {real, imag} */,
  {32'h40b4b8a4, 32'hc21f11e6} /* (26, 24, 30) {real, imag} */,
  {32'hc1fc565c, 32'h428ab0ab} /* (26, 24, 29) {real, imag} */,
  {32'hc2e09564, 32'h41fdcfd2} /* (26, 24, 28) {real, imag} */,
  {32'hc281fe04, 32'h407bac38} /* (26, 24, 27) {real, imag} */,
  {32'hc199189e, 32'hc253e1c2} /* (26, 24, 26) {real, imag} */,
  {32'h425f49a1, 32'h4012c5b0} /* (26, 24, 25) {real, imag} */,
  {32'h422c8408, 32'h424d9504} /* (26, 24, 24) {real, imag} */,
  {32'h41529356, 32'hc21755cd} /* (26, 24, 23) {real, imag} */,
  {32'hc20c5d71, 32'h4123b456} /* (26, 24, 22) {real, imag} */,
  {32'hc13e747b, 32'h419b7443} /* (26, 24, 21) {real, imag} */,
  {32'h4158dac4, 32'h42469841} /* (26, 24, 20) {real, imag} */,
  {32'hc099d3ea, 32'hc265fe89} /* (26, 24, 19) {real, imag} */,
  {32'hc1c68f59, 32'hc0397688} /* (26, 24, 18) {real, imag} */,
  {32'h3fb26478, 32'h4133f3a2} /* (26, 24, 17) {real, imag} */,
  {32'h40a3f5f2, 32'h411e5361} /* (26, 24, 16) {real, imag} */,
  {32'h412ac0a9, 32'hc125986a} /* (26, 24, 15) {real, imag} */,
  {32'hc163d5c2, 32'h40812b64} /* (26, 24, 14) {real, imag} */,
  {32'hc1da6072, 32'h41df0fce} /* (26, 24, 13) {real, imag} */,
  {32'hbfc33be0, 32'h4155d4fc} /* (26, 24, 12) {real, imag} */,
  {32'hc19f6622, 32'h411f5cde} /* (26, 24, 11) {real, imag} */,
  {32'hc1c68ca4, 32'hc202907c} /* (26, 24, 10) {real, imag} */,
  {32'h4283870c, 32'h42a6d8ac} /* (26, 24, 9) {real, imag} */,
  {32'h414953f9, 32'hc2572838} /* (26, 24, 8) {real, imag} */,
  {32'hc16f857c, 32'h42327045} /* (26, 24, 7) {real, imag} */,
  {32'hc22cb0f4, 32'hc2d3964b} /* (26, 24, 6) {real, imag} */,
  {32'hc2b5375e, 32'h4256744e} /* (26, 24, 5) {real, imag} */,
  {32'hc2963a28, 32'h42a24dea} /* (26, 24, 4) {real, imag} */,
  {32'hc22af958, 32'hc2ad91af} /* (26, 24, 3) {real, imag} */,
  {32'h426ac824, 32'h42174136} /* (26, 24, 2) {real, imag} */,
  {32'h41097408, 32'hc28de07e} /* (26, 24, 1) {real, imag} */,
  {32'h41289979, 32'h41ad9432} /* (26, 24, 0) {real, imag} */,
  {32'hc183475f, 32'hc09c6268} /* (26, 23, 31) {real, imag} */,
  {32'h42b8a5b3, 32'hc09bb5e8} /* (26, 23, 30) {real, imag} */,
  {32'h42c29c13, 32'hc24c7a6f} /* (26, 23, 29) {real, imag} */,
  {32'hc22905b7, 32'h42048bff} /* (26, 23, 28) {real, imag} */,
  {32'h415f4492, 32'hc20943a8} /* (26, 23, 27) {real, imag} */,
  {32'h415c0455, 32'hc2128d59} /* (26, 23, 26) {real, imag} */,
  {32'h42a0191d, 32'h4284e012} /* (26, 23, 25) {real, imag} */,
  {32'h41a7b55a, 32'hc08e6db6} /* (26, 23, 24) {real, imag} */,
  {32'h42952965, 32'h41c3be68} /* (26, 23, 23) {real, imag} */,
  {32'hc080177c, 32'h402d89b8} /* (26, 23, 22) {real, imag} */,
  {32'h3fef2eb0, 32'hc1ce570b} /* (26, 23, 21) {real, imag} */,
  {32'h41b400a8, 32'h40238258} /* (26, 23, 20) {real, imag} */,
  {32'h41955121, 32'hc16ef8e0} /* (26, 23, 19) {real, imag} */,
  {32'h3edb5300, 32'h4215726e} /* (26, 23, 18) {real, imag} */,
  {32'h41bdb757, 32'hc06c07b0} /* (26, 23, 17) {real, imag} */,
  {32'h40e27bc2, 32'hc08a4090} /* (26, 23, 16) {real, imag} */,
  {32'h4131824e, 32'hc153d1fa} /* (26, 23, 15) {real, imag} */,
  {32'h4098b2e0, 32'h411cfbb2} /* (26, 23, 14) {real, imag} */,
  {32'hc0f3e2eb, 32'h41b3910c} /* (26, 23, 13) {real, imag} */,
  {32'hc1aa6fb2, 32'hc1d69c70} /* (26, 23, 12) {real, imag} */,
  {32'h410e042a, 32'h419af177} /* (26, 23, 11) {real, imag} */,
  {32'hc2472b68, 32'h41488658} /* (26, 23, 10) {real, imag} */,
  {32'h41a17bc8, 32'h40f30f50} /* (26, 23, 9) {real, imag} */,
  {32'h427475bb, 32'hc07229d4} /* (26, 23, 8) {real, imag} */,
  {32'h4186dc30, 32'hc2b06e72} /* (26, 23, 7) {real, imag} */,
  {32'h4186d1a8, 32'hc132337d} /* (26, 23, 6) {real, imag} */,
  {32'h42997bbc, 32'hc20fcbfe} /* (26, 23, 5) {real, imag} */,
  {32'hc1953b48, 32'hbffbc018} /* (26, 23, 4) {real, imag} */,
  {32'hc2e81231, 32'hc256c047} /* (26, 23, 3) {real, imag} */,
  {32'hbfaa2900, 32'h42db4d8a} /* (26, 23, 2) {real, imag} */,
  {32'hc2013952, 32'hc24eb2f1} /* (26, 23, 1) {real, imag} */,
  {32'hc0fbbd82, 32'hc3395994} /* (26, 23, 0) {real, imag} */,
  {32'h413f051a, 32'hc24865cb} /* (26, 22, 31) {real, imag} */,
  {32'hc0fd86f2, 32'h403ecd88} /* (26, 22, 30) {real, imag} */,
  {32'hbf42f200, 32'hc1e41352} /* (26, 22, 29) {real, imag} */,
  {32'h42b8dde9, 32'hc1a6b685} /* (26, 22, 28) {real, imag} */,
  {32'h41ab43d6, 32'h4285ec51} /* (26, 22, 27) {real, imag} */,
  {32'h423c1cdf, 32'hc2743f75} /* (26, 22, 26) {real, imag} */,
  {32'hc203ced0, 32'hc1b511ab} /* (26, 22, 25) {real, imag} */,
  {32'h418e80f2, 32'hc20a51fc} /* (26, 22, 24) {real, imag} */,
  {32'hc1797458, 32'h421bdf7c} /* (26, 22, 23) {real, imag} */,
  {32'h41047e84, 32'h400d3380} /* (26, 22, 22) {real, imag} */,
  {32'hc237df3a, 32'hc20090bf} /* (26, 22, 21) {real, imag} */,
  {32'hc18f362a, 32'h41c8c63e} /* (26, 22, 20) {real, imag} */,
  {32'h41e96710, 32'hc161270f} /* (26, 22, 19) {real, imag} */,
  {32'hc1d81998, 32'hc1952004} /* (26, 22, 18) {real, imag} */,
  {32'hc04a096e, 32'h40de6360} /* (26, 22, 17) {real, imag} */,
  {32'h40eb98aa, 32'hbf5fbde0} /* (26, 22, 16) {real, imag} */,
  {32'h40f84749, 32'hc204ca97} /* (26, 22, 15) {real, imag} */,
  {32'h40d90170, 32'h3e6a7b00} /* (26, 22, 14) {real, imag} */,
  {32'hc0cd87b8, 32'h41a019d8} /* (26, 22, 13) {real, imag} */,
  {32'hc112c9b3, 32'h41bc608c} /* (26, 22, 12) {real, imag} */,
  {32'hc1408108, 32'h41b450ac} /* (26, 22, 11) {real, imag} */,
  {32'h41be711a, 32'hc22fc3c4} /* (26, 22, 10) {real, imag} */,
  {32'h419eefd4, 32'hc1d729a9} /* (26, 22, 9) {real, imag} */,
  {32'h3e82ac20, 32'h420e5d9c} /* (26, 22, 8) {real, imag} */,
  {32'hc2562338, 32'hc1b0ba1b} /* (26, 22, 7) {real, imag} */,
  {32'hc209529d, 32'h419e9736} /* (26, 22, 6) {real, imag} */,
  {32'hc1c4e156, 32'hc26de349} /* (26, 22, 5) {real, imag} */,
  {32'hc1d3e85c, 32'h425dd996} /* (26, 22, 4) {real, imag} */,
  {32'hc28cb46a, 32'hc1a2f1b2} /* (26, 22, 3) {real, imag} */,
  {32'h4179cd7f, 32'hc1925a4f} /* (26, 22, 2) {real, imag} */,
  {32'hc1d1bff3, 32'hc261965d} /* (26, 22, 1) {real, imag} */,
  {32'h41b9564c, 32'h424eb4ac} /* (26, 22, 0) {real, imag} */,
  {32'hc13e2d48, 32'hc176331c} /* (26, 21, 31) {real, imag} */,
  {32'h4293f748, 32'hc209ceec} /* (26, 21, 30) {real, imag} */,
  {32'h41d893ba, 32'h4263c94c} /* (26, 21, 29) {real, imag} */,
  {32'hc2162de4, 32'hc184fd20} /* (26, 21, 28) {real, imag} */,
  {32'h40ed4230, 32'hc20da45a} /* (26, 21, 27) {real, imag} */,
  {32'h41771e02, 32'hc1d944ed} /* (26, 21, 26) {real, imag} */,
  {32'hc24b8699, 32'h420f4e66} /* (26, 21, 25) {real, imag} */,
  {32'hc16bc3d9, 32'hc122952d} /* (26, 21, 24) {real, imag} */,
  {32'h3fbce820, 32'h4145e589} /* (26, 21, 23) {real, imag} */,
  {32'hc116dd80, 32'h41855b18} /* (26, 21, 22) {real, imag} */,
  {32'hc0656b20, 32'hc140796e} /* (26, 21, 21) {real, imag} */,
  {32'h415fb4ca, 32'hc17167ef} /* (26, 21, 20) {real, imag} */,
  {32'hc030255e, 32'hc19142c9} /* (26, 21, 19) {real, imag} */,
  {32'hbf5d0960, 32'hc13f1f2d} /* (26, 21, 18) {real, imag} */,
  {32'h41a775f0, 32'h3fa04438} /* (26, 21, 17) {real, imag} */,
  {32'hbff95ce0, 32'hc18d1cbf} /* (26, 21, 16) {real, imag} */,
  {32'hc1076944, 32'h419d52ec} /* (26, 21, 15) {real, imag} */,
  {32'h40e1f08c, 32'hc19c3d74} /* (26, 21, 14) {real, imag} */,
  {32'h4128e212, 32'h41004b3e} /* (26, 21, 13) {real, imag} */,
  {32'hc172f7a4, 32'hc1870d34} /* (26, 21, 12) {real, imag} */,
  {32'hc2010ecd, 32'h416612a4} /* (26, 21, 11) {real, imag} */,
  {32'h413d6020, 32'h41f7d282} /* (26, 21, 10) {real, imag} */,
  {32'h416eb5e0, 32'hc1943fd0} /* (26, 21, 9) {real, imag} */,
  {32'h41ea9d2a, 32'hc1f6580e} /* (26, 21, 8) {real, imag} */,
  {32'hc21a0703, 32'hc233c666} /* (26, 21, 7) {real, imag} */,
  {32'h41fac49f, 32'h42a693f9} /* (26, 21, 6) {real, imag} */,
  {32'hc2a99b41, 32'h41c32cfc} /* (26, 21, 5) {real, imag} */,
  {32'hc1807e04, 32'hc1e15780} /* (26, 21, 4) {real, imag} */,
  {32'h40ef1ac8, 32'hbfc0e390} /* (26, 21, 3) {real, imag} */,
  {32'h415990ee, 32'h426c1a90} /* (26, 21, 2) {real, imag} */,
  {32'h412c10ac, 32'h42a3ac4a} /* (26, 21, 1) {real, imag} */,
  {32'h422620e7, 32'hc246efc8} /* (26, 21, 0) {real, imag} */,
  {32'hc23da4af, 32'h4164b551} /* (26, 20, 31) {real, imag} */,
  {32'h4186f4c8, 32'hc102cf7b} /* (26, 20, 30) {real, imag} */,
  {32'hc00ca68c, 32'hbfea9ef4} /* (26, 20, 29) {real, imag} */,
  {32'hc2229ce1, 32'h41659d6a} /* (26, 20, 28) {real, imag} */,
  {32'h42573e90, 32'hc0a3f87e} /* (26, 20, 27) {real, imag} */,
  {32'hc1c7436e, 32'h41077f7c} /* (26, 20, 26) {real, imag} */,
  {32'hc1019732, 32'hc1fc381c} /* (26, 20, 25) {real, imag} */,
  {32'hc1152b7c, 32'hbf1270e0} /* (26, 20, 24) {real, imag} */,
  {32'h408e3309, 32'h403e6c2e} /* (26, 20, 23) {real, imag} */,
  {32'h40b507be, 32'h422b9231} /* (26, 20, 22) {real, imag} */,
  {32'h417cb3fe, 32'hc162cdc0} /* (26, 20, 21) {real, imag} */,
  {32'hc0e4d248, 32'hc112580c} /* (26, 20, 20) {real, imag} */,
  {32'h41836dc1, 32'h411238cf} /* (26, 20, 19) {real, imag} */,
  {32'hc008f010, 32'hbefe9060} /* (26, 20, 18) {real, imag} */,
  {32'h3f119a28, 32'hc09a3e6c} /* (26, 20, 17) {real, imag} */,
  {32'hc0ba3c00, 32'hbf548fb0} /* (26, 20, 16) {real, imag} */,
  {32'hc0364d4a, 32'hc1577c76} /* (26, 20, 15) {real, imag} */,
  {32'h41085110, 32'hc167cc37} /* (26, 20, 14) {real, imag} */,
  {32'h41a6c263, 32'hc16d98b1} /* (26, 20, 13) {real, imag} */,
  {32'h41134b02, 32'hc0058276} /* (26, 20, 12) {real, imag} */,
  {32'hc111ea22, 32'h405f1a62} /* (26, 20, 11) {real, imag} */,
  {32'h41f62828, 32'hc15efbc4} /* (26, 20, 10) {real, imag} */,
  {32'h4199fc12, 32'h4023d712} /* (26, 20, 9) {real, imag} */,
  {32'h41a71704, 32'h41848805} /* (26, 20, 8) {real, imag} */,
  {32'h41bf89e5, 32'hc24ea302} /* (26, 20, 7) {real, imag} */,
  {32'h417f7943, 32'h42287cdd} /* (26, 20, 6) {real, imag} */,
  {32'h41c204d9, 32'hc18d0740} /* (26, 20, 5) {real, imag} */,
  {32'h40125490, 32'hc1fa1f57} /* (26, 20, 4) {real, imag} */,
  {32'hc197c00c, 32'h408fc7d1} /* (26, 20, 3) {real, imag} */,
  {32'hc294b178, 32'h420df868} /* (26, 20, 2) {real, imag} */,
  {32'hc201ae65, 32'hc0e7e292} /* (26, 20, 1) {real, imag} */,
  {32'hc20c524c, 32'h4160aa61} /* (26, 20, 0) {real, imag} */,
  {32'h40c71b38, 32'h4240b519} /* (26, 19, 31) {real, imag} */,
  {32'hc21b61be, 32'h4026cb60} /* (26, 19, 30) {real, imag} */,
  {32'hc21db5dc, 32'h40c6c256} /* (26, 19, 29) {real, imag} */,
  {32'h422d30c2, 32'hc0e31ce2} /* (26, 19, 28) {real, imag} */,
  {32'hc2445918, 32'h41e7137b} /* (26, 19, 27) {real, imag} */,
  {32'hc16358b6, 32'hc20c171c} /* (26, 19, 26) {real, imag} */,
  {32'hc21d6a50, 32'h41ee3594} /* (26, 19, 25) {real, imag} */,
  {32'h4104d511, 32'hc1a1e879} /* (26, 19, 24) {real, imag} */,
  {32'h40c98e21, 32'h401b17b0} /* (26, 19, 23) {real, imag} */,
  {32'hbfd68a60, 32'hc197cfca} /* (26, 19, 22) {real, imag} */,
  {32'hc0f9cd83, 32'hbfaf9830} /* (26, 19, 21) {real, imag} */,
  {32'hc183a5d3, 32'h4188a9a9} /* (26, 19, 20) {real, imag} */,
  {32'h40d3f4a2, 32'h412c7f70} /* (26, 19, 19) {real, imag} */,
  {32'h4122f548, 32'hc210303a} /* (26, 19, 18) {real, imag} */,
  {32'h4087a8c0, 32'h4153534e} /* (26, 19, 17) {real, imag} */,
  {32'hc0126594, 32'h412f926c} /* (26, 19, 16) {real, imag} */,
  {32'h40658608, 32'hbf331ed8} /* (26, 19, 15) {real, imag} */,
  {32'h410936e6, 32'hc050a428} /* (26, 19, 14) {real, imag} */,
  {32'hc1a2fb9e, 32'h40ba56df} /* (26, 19, 13) {real, imag} */,
  {32'h40a63700, 32'h415583ec} /* (26, 19, 12) {real, imag} */,
  {32'h41505c16, 32'hc1912d59} /* (26, 19, 11) {real, imag} */,
  {32'hbf8b7aa0, 32'hc097f196} /* (26, 19, 10) {real, imag} */,
  {32'h40af1335, 32'h41a47c80} /* (26, 19, 9) {real, imag} */,
  {32'h411249a5, 32'h3fdeb6d0} /* (26, 19, 8) {real, imag} */,
  {32'hbe99ba40, 32'h413d1eb4} /* (26, 19, 7) {real, imag} */,
  {32'hc223ed5e, 32'h41ad90bc} /* (26, 19, 6) {real, imag} */,
  {32'h41a6ac1d, 32'h41d89cad} /* (26, 19, 5) {real, imag} */,
  {32'h4042d200, 32'h418364e6} /* (26, 19, 4) {real, imag} */,
  {32'h4214fe54, 32'h3f9b84a0} /* (26, 19, 3) {real, imag} */,
  {32'hc099c210, 32'hc19d2b86} /* (26, 19, 2) {real, imag} */,
  {32'h42480a73, 32'h426a39cd} /* (26, 19, 1) {real, imag} */,
  {32'hc05bdacc, 32'h418f2b5a} /* (26, 19, 0) {real, imag} */,
  {32'hc119fa9c, 32'h4117ba4c} /* (26, 18, 31) {real, imag} */,
  {32'h41ed8804, 32'hc17c1898} /* (26, 18, 30) {real, imag} */,
  {32'h416128bb, 32'h40d71be4} /* (26, 18, 29) {real, imag} */,
  {32'hc148379e, 32'hc008b600} /* (26, 18, 28) {real, imag} */,
  {32'h41ababf6, 32'hc25036d2} /* (26, 18, 27) {real, imag} */,
  {32'hc2289127, 32'hc1496db8} /* (26, 18, 26) {real, imag} */,
  {32'h41264102, 32'h40eb842c} /* (26, 18, 25) {real, imag} */,
  {32'hc08b6284, 32'hc201d4fa} /* (26, 18, 24) {real, imag} */,
  {32'h4175c0a8, 32'hc0de9e91} /* (26, 18, 23) {real, imag} */,
  {32'h412b32b6, 32'hc16597f8} /* (26, 18, 22) {real, imag} */,
  {32'hc0e1c6f2, 32'hc0e65a54} /* (26, 18, 21) {real, imag} */,
  {32'hc0cfca67, 32'hc0d9b356} /* (26, 18, 20) {real, imag} */,
  {32'hc09780de, 32'hc0a6246c} /* (26, 18, 19) {real, imag} */,
  {32'h413a2095, 32'hc0af8b14} /* (26, 18, 18) {real, imag} */,
  {32'hbff103d0, 32'h40b6cdaf} /* (26, 18, 17) {real, imag} */,
  {32'hc086c878, 32'hc0fde238} /* (26, 18, 16) {real, imag} */,
  {32'h403b7110, 32'hc0ca9773} /* (26, 18, 15) {real, imag} */,
  {32'hc0f98a8e, 32'h415d6c1e} /* (26, 18, 14) {real, imag} */,
  {32'hc15545b7, 32'h40fe6bd0} /* (26, 18, 13) {real, imag} */,
  {32'hc144604e, 32'h411500d3} /* (26, 18, 12) {real, imag} */,
  {32'h40966b12, 32'hc1a49049} /* (26, 18, 11) {real, imag} */,
  {32'hc126de8a, 32'h40ab65f4} /* (26, 18, 10) {real, imag} */,
  {32'h4142826a, 32'h4191674a} /* (26, 18, 9) {real, imag} */,
  {32'hc20c1a88, 32'h4198bba6} /* (26, 18, 8) {real, imag} */,
  {32'hc114a320, 32'h3ff21718} /* (26, 18, 7) {real, imag} */,
  {32'hbf168a80, 32'hc24053fa} /* (26, 18, 6) {real, imag} */,
  {32'hc0c79162, 32'hc162a9a6} /* (26, 18, 5) {real, imag} */,
  {32'hbf2b8338, 32'hc18e1e4a} /* (26, 18, 4) {real, imag} */,
  {32'hc14755ad, 32'hc0a182d8} /* (26, 18, 3) {real, imag} */,
  {32'hc082780e, 32'hc21c8d8a} /* (26, 18, 2) {real, imag} */,
  {32'hc2530567, 32'h418f442b} /* (26, 18, 1) {real, imag} */,
  {32'hc22f52d0, 32'hc21b6ef3} /* (26, 18, 0) {real, imag} */,
  {32'hc18befaa, 32'h418a5b20} /* (26, 17, 31) {real, imag} */,
  {32'hbf82b4d8, 32'hc0d98412} /* (26, 17, 30) {real, imag} */,
  {32'h4255bdae, 32'hbffd8510} /* (26, 17, 29) {real, imag} */,
  {32'hc200d902, 32'hc1fba1b1} /* (26, 17, 28) {real, imag} */,
  {32'h3ece4060, 32'h41d04560} /* (26, 17, 27) {real, imag} */,
  {32'hbfbcc630, 32'hc1304fd8} /* (26, 17, 26) {real, imag} */,
  {32'h412913bc, 32'h41db9d80} /* (26, 17, 25) {real, imag} */,
  {32'hc18c7536, 32'h418ad62c} /* (26, 17, 24) {real, imag} */,
  {32'hc1e20432, 32'hc1a6e910} /* (26, 17, 23) {real, imag} */,
  {32'h4166b148, 32'hc1c13187} /* (26, 17, 22) {real, imag} */,
  {32'hc17e2cc7, 32'hbf520568} /* (26, 17, 21) {real, imag} */,
  {32'h4007007a, 32'hbef6ec48} /* (26, 17, 20) {real, imag} */,
  {32'h408a9780, 32'hc0e810d4} /* (26, 17, 19) {real, imag} */,
  {32'hc069f374, 32'h40a5ce86} /* (26, 17, 18) {real, imag} */,
  {32'h3e3696c8, 32'h40f0d662} /* (26, 17, 17) {real, imag} */,
  {32'h40ca4c90, 32'hc0845dba} /* (26, 17, 16) {real, imag} */,
  {32'hc0752ca4, 32'hbf96b1e8} /* (26, 17, 15) {real, imag} */,
  {32'hc1418b27, 32'h4076bd75} /* (26, 17, 14) {real, imag} */,
  {32'hbfda4b70, 32'hc1543e1a} /* (26, 17, 13) {real, imag} */,
  {32'hbfd3e9ec, 32'hbed97638} /* (26, 17, 12) {real, imag} */,
  {32'hc1ad1484, 32'h40366042} /* (26, 17, 11) {real, imag} */,
  {32'hc089c6d8, 32'h41052632} /* (26, 17, 10) {real, imag} */,
  {32'h40423790, 32'h41010c8c} /* (26, 17, 9) {real, imag} */,
  {32'hc211f80b, 32'h41d6a0ae} /* (26, 17, 8) {real, imag} */,
  {32'h4188da16, 32'h41fef4d2} /* (26, 17, 7) {real, imag} */,
  {32'h41b741dd, 32'hc1c07592} /* (26, 17, 6) {real, imag} */,
  {32'hc1cc0352, 32'h41e5b734} /* (26, 17, 5) {real, imag} */,
  {32'h4050f418, 32'hc1b39769} /* (26, 17, 4) {real, imag} */,
  {32'h408fd580, 32'h422a151c} /* (26, 17, 3) {real, imag} */,
  {32'h418d945c, 32'hc1b1dda0} /* (26, 17, 2) {real, imag} */,
  {32'h41a2c8dc, 32'h41f8a322} /* (26, 17, 1) {real, imag} */,
  {32'h424f5c0a, 32'hc19a0b2c} /* (26, 17, 0) {real, imag} */,
  {32'h3d413300, 32'h41b9bdbe} /* (26, 16, 31) {real, imag} */,
  {32'h40123690, 32'hc1a9e6fd} /* (26, 16, 30) {real, imag} */,
  {32'h4151f9e0, 32'h413c0d61} /* (26, 16, 29) {real, imag} */,
  {32'hc21c2c6a, 32'hbff527f6} /* (26, 16, 28) {real, imag} */,
  {32'hc184fc11, 32'hc1d6ad2e} /* (26, 16, 27) {real, imag} */,
  {32'hc0c97820, 32'h4181506a} /* (26, 16, 26) {real, imag} */,
  {32'h4012cb78, 32'h40961285} /* (26, 16, 25) {real, imag} */,
  {32'hc000e898, 32'h3ff4ec40} /* (26, 16, 24) {real, imag} */,
  {32'hc1237472, 32'hc144038a} /* (26, 16, 23) {real, imag} */,
  {32'hbf8a0d58, 32'h41961cce} /* (26, 16, 22) {real, imag} */,
  {32'h400c70aa, 32'hc0709516} /* (26, 16, 21) {real, imag} */,
  {32'hc0fbb58a, 32'hc11a90b1} /* (26, 16, 20) {real, imag} */,
  {32'h410af18a, 32'h40a1df41} /* (26, 16, 19) {real, imag} */,
  {32'h40eb3790, 32'h417b0781} /* (26, 16, 18) {real, imag} */,
  {32'hc00c13c8, 32'h4057b0a2} /* (26, 16, 17) {real, imag} */,
  {32'h3faa1378, 32'h40d4346c} /* (26, 16, 16) {real, imag} */,
  {32'h413c23c3, 32'hc0babb2d} /* (26, 16, 15) {real, imag} */,
  {32'h410a61c1, 32'h4121fee1} /* (26, 16, 14) {real, imag} */,
  {32'h40c95dcb, 32'hc005494a} /* (26, 16, 13) {real, imag} */,
  {32'h413ea319, 32'hbf9111a8} /* (26, 16, 12) {real, imag} */,
  {32'h407386c6, 32'hc1256ba0} /* (26, 16, 11) {real, imag} */,
  {32'h40394bde, 32'hbeaeab60} /* (26, 16, 10) {real, imag} */,
  {32'h403dfa79, 32'hbf1b2688} /* (26, 16, 9) {real, imag} */,
  {32'h413cddab, 32'h41491a27} /* (26, 16, 8) {real, imag} */,
  {32'h40826815, 32'h4115cde4} /* (26, 16, 7) {real, imag} */,
  {32'hc104e18a, 32'hc1a078a6} /* (26, 16, 6) {real, imag} */,
  {32'hc16248e3, 32'h4190443a} /* (26, 16, 5) {real, imag} */,
  {32'hc1706239, 32'h400f233b} /* (26, 16, 4) {real, imag} */,
  {32'h41a8a990, 32'hc10afacb} /* (26, 16, 3) {real, imag} */,
  {32'h419166f2, 32'hc11bff94} /* (26, 16, 2) {real, imag} */,
  {32'h413bf624, 32'h41674e94} /* (26, 16, 1) {real, imag} */,
  {32'h411a2890, 32'hc1085827} /* (26, 16, 0) {real, imag} */,
  {32'hc13b5b70, 32'hc05611cc} /* (26, 15, 31) {real, imag} */,
  {32'hc2a9b2e7, 32'hc147a2c0} /* (26, 15, 30) {real, imag} */,
  {32'h41b878df, 32'hc2191acc} /* (26, 15, 29) {real, imag} */,
  {32'h42001f9c, 32'h40318b98} /* (26, 15, 28) {real, imag} */,
  {32'hc1b95272, 32'h4158e390} /* (26, 15, 27) {real, imag} */,
  {32'hc09eed94, 32'hc158bff6} /* (26, 15, 26) {real, imag} */,
  {32'hc19c85a0, 32'hc1ac41d6} /* (26, 15, 25) {real, imag} */,
  {32'hc10a6b86, 32'h41ad256c} /* (26, 15, 24) {real, imag} */,
  {32'h3f78e998, 32'h40e25e4b} /* (26, 15, 23) {real, imag} */,
  {32'hc1bf2ffb, 32'h419a68e0} /* (26, 15, 22) {real, imag} */,
  {32'h3cf11680, 32'hbf9ea7f0} /* (26, 15, 21) {real, imag} */,
  {32'hbfe3d600, 32'hc0b8dddf} /* (26, 15, 20) {real, imag} */,
  {32'hc109b1c9, 32'h40ff2e6c} /* (26, 15, 19) {real, imag} */,
  {32'h41050039, 32'h40475622} /* (26, 15, 18) {real, imag} */,
  {32'h412e3afe, 32'h405e903c} /* (26, 15, 17) {real, imag} */,
  {32'hc1922365, 32'hc02e5bb8} /* (26, 15, 16) {real, imag} */,
  {32'hbfb5093c, 32'h40e678e2} /* (26, 15, 15) {real, imag} */,
  {32'h3fcdde08, 32'hc1419a84} /* (26, 15, 14) {real, imag} */,
  {32'hc0c7c5b2, 32'h4125c086} /* (26, 15, 13) {real, imag} */,
  {32'h4101317c, 32'h40ba55bf} /* (26, 15, 12) {real, imag} */,
  {32'hc0a808a6, 32'hc14e678d} /* (26, 15, 11) {real, imag} */,
  {32'hc1041fc2, 32'h3c6d6c00} /* (26, 15, 10) {real, imag} */,
  {32'h41814287, 32'hc0f92471} /* (26, 15, 9) {real, imag} */,
  {32'h3f27dbd8, 32'hc13f08cc} /* (26, 15, 8) {real, imag} */,
  {32'h40834240, 32'hc1255ebd} /* (26, 15, 7) {real, imag} */,
  {32'hc20e75b8, 32'h418bde26} /* (26, 15, 6) {real, imag} */,
  {32'hc18f0a32, 32'h41ae0ce6} /* (26, 15, 5) {real, imag} */,
  {32'hc1ca69f3, 32'hc1b5eab9} /* (26, 15, 4) {real, imag} */,
  {32'hc113b21a, 32'hc06c0548} /* (26, 15, 3) {real, imag} */,
  {32'h42744d39, 32'hc2226a93} /* (26, 15, 2) {real, imag} */,
  {32'h415f48a4, 32'hc0b19582} /* (26, 15, 1) {real, imag} */,
  {32'hc219bc38, 32'h4087fb3e} /* (26, 15, 0) {real, imag} */,
  {32'h40c7ad68, 32'hc1ff702d} /* (26, 14, 31) {real, imag} */,
  {32'hc12143e6, 32'hc0d6bc9a} /* (26, 14, 30) {real, imag} */,
  {32'h418117b8, 32'h426696b5} /* (26, 14, 29) {real, imag} */,
  {32'hc261e6f3, 32'hc0f5a56c} /* (26, 14, 28) {real, imag} */,
  {32'hbfd70228, 32'hc17286d2} /* (26, 14, 27) {real, imag} */,
  {32'h420784ea, 32'hc1db4d76} /* (26, 14, 26) {real, imag} */,
  {32'h42137ffe, 32'hc142253e} /* (26, 14, 25) {real, imag} */,
  {32'h3e47d1b0, 32'hc197d943} /* (26, 14, 24) {real, imag} */,
  {32'hc0858bae, 32'hc18adbc2} /* (26, 14, 23) {real, imag} */,
  {32'hc193392a, 32'hc1c7005c} /* (26, 14, 22) {real, imag} */,
  {32'h40d705c2, 32'hbfc95a38} /* (26, 14, 21) {real, imag} */,
  {32'hbfeb7e7c, 32'h40805530} /* (26, 14, 20) {real, imag} */,
  {32'h4011f3f4, 32'h408b3437} /* (26, 14, 19) {real, imag} */,
  {32'h40ca4000, 32'hc12a867e} /* (26, 14, 18) {real, imag} */,
  {32'hc1460540, 32'hbf530638} /* (26, 14, 17) {real, imag} */,
  {32'hc0553879, 32'hbfc6a078} /* (26, 14, 16) {real, imag} */,
  {32'hc0acc128, 32'h3fc54c64} /* (26, 14, 15) {real, imag} */,
  {32'hc17d7b08, 32'h3f08bc58} /* (26, 14, 14) {real, imag} */,
  {32'h408d4446, 32'h4121f078} /* (26, 14, 13) {real, imag} */,
  {32'hc0946a59, 32'h415047d0} /* (26, 14, 12) {real, imag} */,
  {32'hc0ed9b5e, 32'hc1032581} /* (26, 14, 11) {real, imag} */,
  {32'h40d9dc32, 32'h40f3d0ce} /* (26, 14, 10) {real, imag} */,
  {32'hc1fc4ea8, 32'h4021e0f0} /* (26, 14, 9) {real, imag} */,
  {32'h402c5493, 32'hc0f26703} /* (26, 14, 8) {real, imag} */,
  {32'h405c4660, 32'hc13bdbc2} /* (26, 14, 7) {real, imag} */,
  {32'hc1dc80e7, 32'h41c833d2} /* (26, 14, 6) {real, imag} */,
  {32'hbf548e10, 32'hc0e23758} /* (26, 14, 5) {real, imag} */,
  {32'hc1f89222, 32'hc1e0ef95} /* (26, 14, 4) {real, imag} */,
  {32'h41fbde78, 32'hc24a1547} /* (26, 14, 3) {real, imag} */,
  {32'hc112a992, 32'hc0c5103c} /* (26, 14, 2) {real, imag} */,
  {32'hc23c4a9a, 32'h414d4a36} /* (26, 14, 1) {real, imag} */,
  {32'h40125edb, 32'h41731ee3} /* (26, 14, 0) {real, imag} */,
  {32'hc17230a4, 32'hbeca32c0} /* (26, 13, 31) {real, imag} */,
  {32'h41bf82b4, 32'hc1d7c55e} /* (26, 13, 30) {real, imag} */,
  {32'hc1df0e7d, 32'hc012b80e} /* (26, 13, 29) {real, imag} */,
  {32'hc09d98e8, 32'h41db4702} /* (26, 13, 28) {real, imag} */,
  {32'h41cab528, 32'h417cd26a} /* (26, 13, 27) {real, imag} */,
  {32'hc1bf08b2, 32'hc132b384} /* (26, 13, 26) {real, imag} */,
  {32'hc14dc91a, 32'h40d01877} /* (26, 13, 25) {real, imag} */,
  {32'h41103959, 32'hc1374d1d} /* (26, 13, 24) {real, imag} */,
  {32'h4215ad9a, 32'h41400c4e} /* (26, 13, 23) {real, imag} */,
  {32'h41c1f9fb, 32'h414715fe} /* (26, 13, 22) {real, imag} */,
  {32'hc0b78f55, 32'hc1645195} /* (26, 13, 21) {real, imag} */,
  {32'hc1b24be0, 32'h3e8a32e0} /* (26, 13, 20) {real, imag} */,
  {32'hc10b9deb, 32'h406a2fba} /* (26, 13, 19) {real, imag} */,
  {32'hc0de3ff3, 32'h41748a00} /* (26, 13, 18) {real, imag} */,
  {32'hc1470003, 32'h40cbee2e} /* (26, 13, 17) {real, imag} */,
  {32'h3fa2feb4, 32'hbfa66560} /* (26, 13, 16) {real, imag} */,
  {32'h40ce7c12, 32'hc042608c} /* (26, 13, 15) {real, imag} */,
  {32'hbf699bd8, 32'hc123805a} /* (26, 13, 14) {real, imag} */,
  {32'h4118f005, 32'h416fe5d2} /* (26, 13, 13) {real, imag} */,
  {32'h4013e250, 32'h416da261} /* (26, 13, 12) {real, imag} */,
  {32'h400eb97e, 32'h417413cf} /* (26, 13, 11) {real, imag} */,
  {32'hc098197c, 32'hc143c06e} /* (26, 13, 10) {real, imag} */,
  {32'hc19357e3, 32'hc0438646} /* (26, 13, 9) {real, imag} */,
  {32'h41d076b6, 32'h4118d537} /* (26, 13, 8) {real, imag} */,
  {32'hc241c624, 32'h40e8d12f} /* (26, 13, 7) {real, imag} */,
  {32'hc1b7556e, 32'hc13ed610} /* (26, 13, 6) {real, imag} */,
  {32'hc097f55e, 32'h401a2ad2} /* (26, 13, 5) {real, imag} */,
  {32'hc1a95114, 32'h41c90d62} /* (26, 13, 4) {real, imag} */,
  {32'hc1a974ef, 32'hc1665680} /* (26, 13, 3) {real, imag} */,
  {32'h41031037, 32'h4211440f} /* (26, 13, 2) {real, imag} */,
  {32'hc1a0fbba, 32'hc270d058} /* (26, 13, 1) {real, imag} */,
  {32'hc0fbe02b, 32'h41e9a8fb} /* (26, 13, 0) {real, imag} */,
  {32'h411ee0b5, 32'h41ab4a8a} /* (26, 12, 31) {real, imag} */,
  {32'h41cf7632, 32'hc0c924e0} /* (26, 12, 30) {real, imag} */,
  {32'hc20de510, 32'hc1f94920} /* (26, 12, 29) {real, imag} */,
  {32'hc207d209, 32'hc21e093b} /* (26, 12, 28) {real, imag} */,
  {32'hc1958a48, 32'h4215a820} /* (26, 12, 27) {real, imag} */,
  {32'hc2102dc8, 32'hc199e48a} /* (26, 12, 26) {real, imag} */,
  {32'h3f79d7b4, 32'h41895e89} /* (26, 12, 25) {real, imag} */,
  {32'hc202a464, 32'hc12146d2} /* (26, 12, 24) {real, imag} */,
  {32'h4187b037, 32'h4194f67c} /* (26, 12, 23) {real, imag} */,
  {32'h416d3e10, 32'h414d1dc1} /* (26, 12, 22) {real, imag} */,
  {32'h41ab91ca, 32'hc19293be} /* (26, 12, 21) {real, imag} */,
  {32'hc1797c05, 32'h4133e90e} /* (26, 12, 20) {real, imag} */,
  {32'h41913f12, 32'h4085da36} /* (26, 12, 19) {real, imag} */,
  {32'hbf384df0, 32'hc0faf81c} /* (26, 12, 18) {real, imag} */,
  {32'h4102d6a7, 32'hc184e030} /* (26, 12, 17) {real, imag} */,
  {32'hc0ae2081, 32'hc185aff5} /* (26, 12, 16) {real, imag} */,
  {32'hbeacfba0, 32'hbff91868} /* (26, 12, 15) {real, imag} */,
  {32'hc02ab504, 32'hc1a7c965} /* (26, 12, 14) {real, imag} */,
  {32'h40bd49b4, 32'h40f97f9e} /* (26, 12, 13) {real, imag} */,
  {32'h41a41dc6, 32'hc06ce4f8} /* (26, 12, 12) {real, imag} */,
  {32'hc1503954, 32'h414a7b86} /* (26, 12, 11) {real, imag} */,
  {32'h41990576, 32'h41de342a} /* (26, 12, 10) {real, imag} */,
  {32'hc1ad2659, 32'hc195b48c} /* (26, 12, 9) {real, imag} */,
  {32'h41d71189, 32'h425713d6} /* (26, 12, 8) {real, imag} */,
  {32'h3f39bf94, 32'hc118fe06} /* (26, 12, 7) {real, imag} */,
  {32'h4128a822, 32'h40a425f6} /* (26, 12, 6) {real, imag} */,
  {32'hc03dd4a0, 32'hc1e4a9ac} /* (26, 12, 5) {real, imag} */,
  {32'hc0d304b8, 32'h4199be90} /* (26, 12, 4) {real, imag} */,
  {32'hc054a280, 32'h42248600} /* (26, 12, 3) {real, imag} */,
  {32'h427271e7, 32'hc2398b82} /* (26, 12, 2) {real, imag} */,
  {32'hc2233f85, 32'hc1b7ac02} /* (26, 12, 1) {real, imag} */,
  {32'h41577cce, 32'hc215fa5e} /* (26, 12, 0) {real, imag} */,
  {32'hc2968d6b, 32'hc1a8cfe2} /* (26, 11, 31) {real, imag} */,
  {32'h4298f8f4, 32'h41af4a50} /* (26, 11, 30) {real, imag} */,
  {32'h42226d00, 32'h41884b24} /* (26, 11, 29) {real, imag} */,
  {32'hc1ccbde0, 32'h423ffe70} /* (26, 11, 28) {real, imag} */,
  {32'hc2542c33, 32'hc04e42b6} /* (26, 11, 27) {real, imag} */,
  {32'hc1c415ee, 32'hc0b9f336} /* (26, 11, 26) {real, imag} */,
  {32'hc1f81566, 32'h4228bf94} /* (26, 11, 25) {real, imag} */,
  {32'h41cb676c, 32'hc0e1dacc} /* (26, 11, 24) {real, imag} */,
  {32'h410c7567, 32'hc1ba68e6} /* (26, 11, 23) {real, imag} */,
  {32'h4091c660, 32'h412257f8} /* (26, 11, 22) {real, imag} */,
  {32'hc1659695, 32'hc170b3a8} /* (26, 11, 21) {real, imag} */,
  {32'hc1cc63eb, 32'h41a86d87} /* (26, 11, 20) {real, imag} */,
  {32'h4021568e, 32'h41c46570} /* (26, 11, 19) {real, imag} */,
  {32'hc0fee6d0, 32'hc16346a6} /* (26, 11, 18) {real, imag} */,
  {32'h4112e040, 32'hc0bba838} /* (26, 11, 17) {real, imag} */,
  {32'hc097c06e, 32'h412c2a7e} /* (26, 11, 16) {real, imag} */,
  {32'hc0e11018, 32'hc1b00549} /* (26, 11, 15) {real, imag} */,
  {32'h40c3b2b8, 32'hbf39eee0} /* (26, 11, 14) {real, imag} */,
  {32'hc1705f64, 32'h41d54e64} /* (26, 11, 13) {real, imag} */,
  {32'hc08e50e4, 32'h41999b45} /* (26, 11, 12) {real, imag} */,
  {32'hc1837386, 32'hc19eec9c} /* (26, 11, 11) {real, imag} */,
  {32'hc129f2ec, 32'hc128bd1e} /* (26, 11, 10) {real, imag} */,
  {32'h418bf4c6, 32'h427d8c55} /* (26, 11, 9) {real, imag} */,
  {32'h418d9d90, 32'h420e6d0a} /* (26, 11, 8) {real, imag} */,
  {32'h4019be70, 32'hc1c92498} /* (26, 11, 7) {real, imag} */,
  {32'hc2293dc5, 32'hc1cb339a} /* (26, 11, 6) {real, imag} */,
  {32'hc0f7d478, 32'h410141de} /* (26, 11, 5) {real, imag} */,
  {32'h41834714, 32'h42830d8d} /* (26, 11, 4) {real, imag} */,
  {32'hc29232b5, 32'hc168c1c8} /* (26, 11, 3) {real, imag} */,
  {32'hc18a85c7, 32'h41387600} /* (26, 11, 2) {real, imag} */,
  {32'h41f8cd3d, 32'hc20d78b9} /* (26, 11, 1) {real, imag} */,
  {32'h4208fc03, 32'h40e202b4} /* (26, 11, 0) {real, imag} */,
  {32'hc15b1f3e, 32'hc1ec4997} /* (26, 10, 31) {real, imag} */,
  {32'hc245e786, 32'hc1c10a3e} /* (26, 10, 30) {real, imag} */,
  {32'h42a729f0, 32'hc0369920} /* (26, 10, 29) {real, imag} */,
  {32'hc0bb991f, 32'hc186e5f0} /* (26, 10, 28) {real, imag} */,
  {32'hc1c8f7f3, 32'hc295019a} /* (26, 10, 27) {real, imag} */,
  {32'hc10d2e6c, 32'h42adbade} /* (26, 10, 26) {real, imag} */,
  {32'hc20233a1, 32'hc2172bda} /* (26, 10, 25) {real, imag} */,
  {32'h42ac6fa0, 32'h41ffcfe7} /* (26, 10, 24) {real, imag} */,
  {32'h41b4ca56, 32'hc0e462a8} /* (26, 10, 23) {real, imag} */,
  {32'h40dd7920, 32'hc232c7ef} /* (26, 10, 22) {real, imag} */,
  {32'hc11e4370, 32'h3fd9ca00} /* (26, 10, 21) {real, imag} */,
  {32'h41877c89, 32'h401a9afc} /* (26, 10, 20) {real, imag} */,
  {32'hc14f513f, 32'h4083a01a} /* (26, 10, 19) {real, imag} */,
  {32'h40cf952e, 32'h40c9f704} /* (26, 10, 18) {real, imag} */,
  {32'hbf289340, 32'h42075783} /* (26, 10, 17) {real, imag} */,
  {32'h41c08d50, 32'hc0d20cec} /* (26, 10, 16) {real, imag} */,
  {32'hbfb1ea68, 32'hc0341b70} /* (26, 10, 15) {real, imag} */,
  {32'h40b7caba, 32'hc181d5f3} /* (26, 10, 14) {real, imag} */,
  {32'hc138dc99, 32'h3fefbba8} /* (26, 10, 13) {real, imag} */,
  {32'h4121b2fe, 32'h40600d8c} /* (26, 10, 12) {real, imag} */,
  {32'hc14b0a88, 32'hc110aea0} /* (26, 10, 11) {real, imag} */,
  {32'hc1b3f50c, 32'h417bec4c} /* (26, 10, 10) {real, imag} */,
  {32'hc0d01e12, 32'h41b0fa8c} /* (26, 10, 9) {real, imag} */,
  {32'h42140b48, 32'hc281ae7c} /* (26, 10, 8) {real, imag} */,
  {32'hbf107710, 32'h418fe5a6} /* (26, 10, 7) {real, imag} */,
  {32'h4299b7c0, 32'h41802f6a} /* (26, 10, 6) {real, imag} */,
  {32'h418711b7, 32'h40117f70} /* (26, 10, 5) {real, imag} */,
  {32'hc1a6fda8, 32'h4290dd06} /* (26, 10, 4) {real, imag} */,
  {32'h4287a710, 32'hc24b4500} /* (26, 10, 3) {real, imag} */,
  {32'hc19c66d4, 32'hc1bafe50} /* (26, 10, 2) {real, imag} */,
  {32'h3e066a40, 32'h40d8f8e4} /* (26, 10, 1) {real, imag} */,
  {32'hc2779628, 32'h4206d598} /* (26, 10, 0) {real, imag} */,
  {32'h413979d7, 32'hc15f8708} /* (26, 9, 31) {real, imag} */,
  {32'hc077e100, 32'h42bb98c4} /* (26, 9, 30) {real, imag} */,
  {32'hbfea0980, 32'hc275c726} /* (26, 9, 29) {real, imag} */,
  {32'hc262df7a, 32'hc1dc433e} /* (26, 9, 28) {real, imag} */,
  {32'h4212e484, 32'hc2972ea4} /* (26, 9, 27) {real, imag} */,
  {32'h420f9f26, 32'h41683e12} /* (26, 9, 26) {real, imag} */,
  {32'h409eb520, 32'hc22a549e} /* (26, 9, 25) {real, imag} */,
  {32'hc2178af0, 32'hc1022b3f} /* (26, 9, 24) {real, imag} */,
  {32'hc11c9600, 32'h41eda931} /* (26, 9, 23) {real, imag} */,
  {32'h41b1d1d6, 32'h423e7abd} /* (26, 9, 22) {real, imag} */,
  {32'h41322559, 32'hc222aec9} /* (26, 9, 21) {real, imag} */,
  {32'h41b1cca2, 32'h41a322a9} /* (26, 9, 20) {real, imag} */,
  {32'hc0fea95c, 32'hc112d3a2} /* (26, 9, 19) {real, imag} */,
  {32'hc14fe07d, 32'h42125f5a} /* (26, 9, 18) {real, imag} */,
  {32'hc138cea5, 32'h40d9f39c} /* (26, 9, 17) {real, imag} */,
  {32'hc1f42998, 32'h41e1f767} /* (26, 9, 16) {real, imag} */,
  {32'hc1809284, 32'h40d5942c} /* (26, 9, 15) {real, imag} */,
  {32'h418caf36, 32'hc175046e} /* (26, 9, 14) {real, imag} */,
  {32'hc04233c0, 32'h41462a54} /* (26, 9, 13) {real, imag} */,
  {32'hc19e9d8e, 32'h40f44fd4} /* (26, 9, 12) {real, imag} */,
  {32'h4159e161, 32'hc20ec2f3} /* (26, 9, 11) {real, imag} */,
  {32'hc164e3d1, 32'hc2402d41} /* (26, 9, 10) {real, imag} */,
  {32'h4288e649, 32'hc15737b2} /* (26, 9, 9) {real, imag} */,
  {32'hc1229aa2, 32'h41df03ba} /* (26, 9, 8) {real, imag} */,
  {32'h4258e3ba, 32'h405ada10} /* (26, 9, 7) {real, imag} */,
  {32'h40787598, 32'hc28438eb} /* (26, 9, 6) {real, imag} */,
  {32'h417e619a, 32'h4191177b} /* (26, 9, 5) {real, imag} */,
  {32'h41d1ed85, 32'h41eda8ae} /* (26, 9, 4) {real, imag} */,
  {32'h425579e8, 32'h4162adb0} /* (26, 9, 3) {real, imag} */,
  {32'h42470d92, 32'h41ef6203} /* (26, 9, 2) {real, imag} */,
  {32'h4185f0a2, 32'h4172ae30} /* (26, 9, 1) {real, imag} */,
  {32'h424c1824, 32'h422ecf4f} /* (26, 9, 0) {real, imag} */,
  {32'hc1e7e766, 32'h4165aa3b} /* (26, 8, 31) {real, imag} */,
  {32'hc2fc998d, 32'hc318ec84} /* (26, 8, 30) {real, imag} */,
  {32'hc0df9bae, 32'h42aa83d6} /* (26, 8, 29) {real, imag} */,
  {32'h41d7bdde, 32'hc257a92d} /* (26, 8, 28) {real, imag} */,
  {32'hc170cd47, 32'hc0b80fa3} /* (26, 8, 27) {real, imag} */,
  {32'hc27a5b1b, 32'h42b1e84c} /* (26, 8, 26) {real, imag} */,
  {32'h41136e60, 32'hc01e5714} /* (26, 8, 25) {real, imag} */,
  {32'hc2a1b808, 32'h3ff00528} /* (26, 8, 24) {real, imag} */,
  {32'h41418810, 32'h41b55fe7} /* (26, 8, 23) {real, imag} */,
  {32'h41f5fd79, 32'hc1f8c743} /* (26, 8, 22) {real, imag} */,
  {32'hc1f2d7ac, 32'h42381544} /* (26, 8, 21) {real, imag} */,
  {32'h41f3c880, 32'h4166fca2} /* (26, 8, 20) {real, imag} */,
  {32'hc0ca55fa, 32'hc16de18b} /* (26, 8, 19) {real, imag} */,
  {32'h40f85e40, 32'h420a6f1b} /* (26, 8, 18) {real, imag} */,
  {32'h40677198, 32'hc12d9229} /* (26, 8, 17) {real, imag} */,
  {32'hc16071a0, 32'hc1b73d10} /* (26, 8, 16) {real, imag} */,
  {32'hc160ed1e, 32'h41adf7d4} /* (26, 8, 15) {real, imag} */,
  {32'h41f29448, 32'h419947ee} /* (26, 8, 14) {real, imag} */,
  {32'hc1f51bb6, 32'hc1c0b3b6} /* (26, 8, 13) {real, imag} */,
  {32'hc1426ec8, 32'h4190c439} /* (26, 8, 12) {real, imag} */,
  {32'hc1af8542, 32'h4212fc30} /* (26, 8, 11) {real, imag} */,
  {32'hc16534a2, 32'h426184c2} /* (26, 8, 10) {real, imag} */,
  {32'h4262f0c0, 32'h41f26245} /* (26, 8, 9) {real, imag} */,
  {32'h41a8cf63, 32'hc1deb2a0} /* (26, 8, 8) {real, imag} */,
  {32'h42ca4292, 32'hc1c1de4a} /* (26, 8, 7) {real, imag} */,
  {32'h416efac4, 32'h40e01280} /* (26, 8, 6) {real, imag} */,
  {32'hc219819d, 32'hc1253e8e} /* (26, 8, 5) {real, imag} */,
  {32'h42803c72, 32'h41c1b276} /* (26, 8, 4) {real, imag} */,
  {32'hc02f21e4, 32'h42968b92} /* (26, 8, 3) {real, imag} */,
  {32'h4289f37d, 32'h433115ec} /* (26, 8, 2) {real, imag} */,
  {32'hc269a40f, 32'hc225184d} /* (26, 8, 1) {real, imag} */,
  {32'h42d9646a, 32'hc21537ae} /* (26, 8, 0) {real, imag} */,
  {32'h4290dbe5, 32'h42d4311a} /* (26, 7, 31) {real, imag} */,
  {32'hc22b36ca, 32'h417a0c52} /* (26, 7, 30) {real, imag} */,
  {32'h3f8f31be, 32'h423315b1} /* (26, 7, 29) {real, imag} */,
  {32'hc29730f2, 32'h428ffcf7} /* (26, 7, 28) {real, imag} */,
  {32'h40f98bae, 32'hc294cf7c} /* (26, 7, 27) {real, imag} */,
  {32'hc2015e6e, 32'h423eebad} /* (26, 7, 26) {real, imag} */,
  {32'h41c9045e, 32'hc1d2925a} /* (26, 7, 25) {real, imag} */,
  {32'hc2b2c89e, 32'h41914844} /* (26, 7, 24) {real, imag} */,
  {32'h41240930, 32'h40387ea8} /* (26, 7, 23) {real, imag} */,
  {32'hc0c7a228, 32'hc2099ea9} /* (26, 7, 22) {real, imag} */,
  {32'h4225e9dd, 32'h4252800e} /* (26, 7, 21) {real, imag} */,
  {32'hc1dae4e6, 32'hbf8c75e8} /* (26, 7, 20) {real, imag} */,
  {32'hc0ce3368, 32'h41f320ba} /* (26, 7, 19) {real, imag} */,
  {32'hc1eebd94, 32'hc1b37099} /* (26, 7, 18) {real, imag} */,
  {32'h413ac133, 32'hc1a44f58} /* (26, 7, 17) {real, imag} */,
  {32'hc1a2fee8, 32'hc1a637bc} /* (26, 7, 16) {real, imag} */,
  {32'hc088d7c6, 32'h422a8ef6} /* (26, 7, 15) {real, imag} */,
  {32'hbf963920, 32'h421773c5} /* (26, 7, 14) {real, imag} */,
  {32'hc127d15e, 32'h40232a10} /* (26, 7, 13) {real, imag} */,
  {32'h414d73e3, 32'h3f149fb0} /* (26, 7, 12) {real, imag} */,
  {32'h4202cb83, 32'hc184b4d4} /* (26, 7, 11) {real, imag} */,
  {32'hc21472d7, 32'hc10423ff} /* (26, 7, 10) {real, imag} */,
  {32'hc142bcce, 32'hc1326232} /* (26, 7, 9) {real, imag} */,
  {32'h41afb220, 32'hc283e461} /* (26, 7, 8) {real, imag} */,
  {32'hc0fe183a, 32'h4267669b} /* (26, 7, 7) {real, imag} */,
  {32'hc1dd482c, 32'h429a0e5a} /* (26, 7, 6) {real, imag} */,
  {32'h41a224e4, 32'hc144f6e0} /* (26, 7, 5) {real, imag} */,
  {32'h41b22baa, 32'hc1163c08} /* (26, 7, 4) {real, imag} */,
  {32'h406976e9, 32'hc321862d} /* (26, 7, 3) {real, imag} */,
  {32'hc12390fc, 32'hc1d26e05} /* (26, 7, 2) {real, imag} */,
  {32'h42aa7709, 32'h42c14bde} /* (26, 7, 1) {real, imag} */,
  {32'hc23b07fc, 32'h42a2e485} /* (26, 7, 0) {real, imag} */,
  {32'h427a3128, 32'h42083bad} /* (26, 6, 31) {real, imag} */,
  {32'hc2b59c57, 32'hc0f4acea} /* (26, 6, 30) {real, imag} */,
  {32'h4324ddae, 32'h3ff8b7e0} /* (26, 6, 29) {real, imag} */,
  {32'h420a23e3, 32'hc2d8333a} /* (26, 6, 28) {real, imag} */,
  {32'h42869f14, 32'hc0fe4670} /* (26, 6, 27) {real, imag} */,
  {32'h42d90949, 32'hc28f9681} /* (26, 6, 26) {real, imag} */,
  {32'hc2394ebf, 32'h42ff4abf} /* (26, 6, 25) {real, imag} */,
  {32'hc20ec687, 32'h4191a1c6} /* (26, 6, 24) {real, imag} */,
  {32'h3fe32f10, 32'hc06a0388} /* (26, 6, 23) {real, imag} */,
  {32'hc21eb608, 32'h41659fb7} /* (26, 6, 22) {real, imag} */,
  {32'h42042a32, 32'hc1485b60} /* (26, 6, 21) {real, imag} */,
  {32'h411de987, 32'h416aa8b8} /* (26, 6, 20) {real, imag} */,
  {32'hc21843fb, 32'h419d34a2} /* (26, 6, 19) {real, imag} */,
  {32'h40238b10, 32'h41a74cc0} /* (26, 6, 18) {real, imag} */,
  {32'hc12b63c2, 32'h3f164430} /* (26, 6, 17) {real, imag} */,
  {32'h41b8166a, 32'h3ed4d300} /* (26, 6, 16) {real, imag} */,
  {32'hc0bdb42c, 32'hc18399e6} /* (26, 6, 15) {real, imag} */,
  {32'h412df428, 32'h40c2056c} /* (26, 6, 14) {real, imag} */,
  {32'hc1e04672, 32'hc283b14c} /* (26, 6, 13) {real, imag} */,
  {32'h415d4c39, 32'h4195cbc4} /* (26, 6, 12) {real, imag} */,
  {32'hc0b10acc, 32'h415d211c} /* (26, 6, 11) {real, imag} */,
  {32'hc252ec50, 32'hc09da8de} /* (26, 6, 10) {real, imag} */,
  {32'h425657a6, 32'hc253df2a} /* (26, 6, 9) {real, imag} */,
  {32'h40ea1318, 32'hc2c128c0} /* (26, 6, 8) {real, imag} */,
  {32'h425ee2f9, 32'h41d166f4} /* (26, 6, 7) {real, imag} */,
  {32'h4190adfc, 32'hc209f1c4} /* (26, 6, 6) {real, imag} */,
  {32'hc1b1a13e, 32'h4102ed64} /* (26, 6, 5) {real, imag} */,
  {32'hc1159794, 32'h42d03152} /* (26, 6, 4) {real, imag} */,
  {32'hc1d2a23c, 32'hc2da16d0} /* (26, 6, 3) {real, imag} */,
  {32'hc17194e8, 32'hc1c4dbda} /* (26, 6, 2) {real, imag} */,
  {32'h42da9978, 32'h42c265b2} /* (26, 6, 1) {real, imag} */,
  {32'h41d6bc66, 32'hc31b2bca} /* (26, 6, 0) {real, imag} */,
  {32'hc2a0a33a, 32'h4276cb6e} /* (26, 5, 31) {real, imag} */,
  {32'h41c75d9c, 32'hc0b71fc8} /* (26, 5, 30) {real, imag} */,
  {32'hc2187d72, 32'hc1e07773} /* (26, 5, 29) {real, imag} */,
  {32'hc275136c, 32'h41c8c574} /* (26, 5, 28) {real, imag} */,
  {32'h40d6b1cc, 32'h4309dc09} /* (26, 5, 27) {real, imag} */,
  {32'h411ce41f, 32'hc10067bc} /* (26, 5, 26) {real, imag} */,
  {32'h423822e2, 32'hc0a5c04c} /* (26, 5, 25) {real, imag} */,
  {32'hc0fc1cd8, 32'h42804dea} /* (26, 5, 24) {real, imag} */,
  {32'h413d0f29, 32'h425ccf55} /* (26, 5, 23) {real, imag} */,
  {32'hc28a68b6, 32'hc1a591b6} /* (26, 5, 22) {real, imag} */,
  {32'h41fe7363, 32'hc1864e74} /* (26, 5, 21) {real, imag} */,
  {32'h42aaa99b, 32'hc1f30d90} /* (26, 5, 20) {real, imag} */,
  {32'hc1c76df0, 32'h419a16b9} /* (26, 5, 19) {real, imag} */,
  {32'h40642ce8, 32'hc1a1822e} /* (26, 5, 18) {real, imag} */,
  {32'hc12d7ad3, 32'hc19ee658} /* (26, 5, 17) {real, imag} */,
  {32'hc193ee7e, 32'h41e43e68} /* (26, 5, 16) {real, imag} */,
  {32'hc025a974, 32'hc07ec15c} /* (26, 5, 15) {real, imag} */,
  {32'h41228fa6, 32'hc1984156} /* (26, 5, 14) {real, imag} */,
  {32'h41c60ab0, 32'h4286e72b} /* (26, 5, 13) {real, imag} */,
  {32'h41d413fb, 32'h419726c8} /* (26, 5, 12) {real, imag} */,
  {32'hbffa6910, 32'h40f12150} /* (26, 5, 11) {real, imag} */,
  {32'h427b2514, 32'hc1f34150} /* (26, 5, 10) {real, imag} */,
  {32'h3fb7aa48, 32'hc0a40e38} /* (26, 5, 9) {real, imag} */,
  {32'h42972646, 32'h428b8f1e} /* (26, 5, 8) {real, imag} */,
  {32'hc29e69a5, 32'hc1d16dec} /* (26, 5, 7) {real, imag} */,
  {32'h40f337ce, 32'hc125f060} /* (26, 5, 6) {real, imag} */,
  {32'hc20b6906, 32'hc064e840} /* (26, 5, 5) {real, imag} */,
  {32'hc2e2e0ac, 32'h41afaa8c} /* (26, 5, 4) {real, imag} */,
  {32'hc11b62e0, 32'hc256204c} /* (26, 5, 3) {real, imag} */,
  {32'h4303b26a, 32'h42883f88} /* (26, 5, 2) {real, imag} */,
  {32'hc1c5ea26, 32'hc25649e4} /* (26, 5, 1) {real, imag} */,
  {32'h403e130c, 32'h42ce318e} /* (26, 5, 0) {real, imag} */,
  {32'hc2c8dad6, 32'hc22437b3} /* (26, 4, 31) {real, imag} */,
  {32'h430227c8, 32'hc2c2c969} /* (26, 4, 30) {real, imag} */,
  {32'h42ebfbc2, 32'hc23a55ef} /* (26, 4, 29) {real, imag} */,
  {32'h42b28f7d, 32'hc254c42b} /* (26, 4, 28) {real, imag} */,
  {32'h3e3afe00, 32'h42b4ff5e} /* (26, 4, 27) {real, imag} */,
  {32'hc219c3b7, 32'h431c1902} /* (26, 4, 26) {real, imag} */,
  {32'h43179d7b, 32'h41e1ddb0} /* (26, 4, 25) {real, imag} */,
  {32'h4282780d, 32'hc12cf85a} /* (26, 4, 24) {real, imag} */,
  {32'h41a2a30e, 32'hc231c96c} /* (26, 4, 23) {real, imag} */,
  {32'h4145462c, 32'hc2339e90} /* (26, 4, 22) {real, imag} */,
  {32'hc25b5d1e, 32'hc23fefcf} /* (26, 4, 21) {real, imag} */,
  {32'h425516f2, 32'h42846188} /* (26, 4, 20) {real, imag} */,
  {32'hc1fbb801, 32'h42a5fa92} /* (26, 4, 19) {real, imag} */,
  {32'h41e74c3e, 32'h40b81578} /* (26, 4, 18) {real, imag} */,
  {32'h41ec1d88, 32'h40bd94b0} /* (26, 4, 17) {real, imag} */,
  {32'hc162c786, 32'h41a2825c} /* (26, 4, 16) {real, imag} */,
  {32'hc1ee6b6c, 32'h4236ea68} /* (26, 4, 15) {real, imag} */,
  {32'h411502dc, 32'h40c67ef0} /* (26, 4, 14) {real, imag} */,
  {32'hc27a62d8, 32'hc1c585b2} /* (26, 4, 13) {real, imag} */,
  {32'h421a8aca, 32'h41a418d5} /* (26, 4, 12) {real, imag} */,
  {32'hc0e070d0, 32'hc2130ba5} /* (26, 4, 11) {real, imag} */,
  {32'h4089f588, 32'hc18d73ab} /* (26, 4, 10) {real, imag} */,
  {32'hc14b9fa4, 32'h41caaa41} /* (26, 4, 9) {real, imag} */,
  {32'h42ad103f, 32'h419cf149} /* (26, 4, 8) {real, imag} */,
  {32'h42862526, 32'hc27b3c7c} /* (26, 4, 7) {real, imag} */,
  {32'hc3094143, 32'hc19a9290} /* (26, 4, 6) {real, imag} */,
  {32'h42d41ead, 32'hc28eb16a} /* (26, 4, 5) {real, imag} */,
  {32'h41bf32f4, 32'h4298c523} /* (26, 4, 4) {real, imag} */,
  {32'h432e323b, 32'h42dbbc22} /* (26, 4, 3) {real, imag} */,
  {32'hc31603de, 32'hc14fc6a8} /* (26, 4, 2) {real, imag} */,
  {32'hc2bc2d1a, 32'h42d46abe} /* (26, 4, 1) {real, imag} */,
  {32'h418ff82f, 32'hc16d1a00} /* (26, 4, 0) {real, imag} */,
  {32'h4267e0bb, 32'hc116f520} /* (26, 3, 31) {real, imag} */,
  {32'hc27942cb, 32'hc32b75f6} /* (26, 3, 30) {real, imag} */,
  {32'h424e64fd, 32'hc30b930d} /* (26, 3, 29) {real, imag} */,
  {32'hc29c1125, 32'h411f9a06} /* (26, 3, 28) {real, imag} */,
  {32'hc283e50d, 32'h430eb8cc} /* (26, 3, 27) {real, imag} */,
  {32'h41cf05e8, 32'hc23893eb} /* (26, 3, 26) {real, imag} */,
  {32'h4216b603, 32'h420a58d7} /* (26, 3, 25) {real, imag} */,
  {32'h430b83f1, 32'hc141393c} /* (26, 3, 24) {real, imag} */,
  {32'h4190fd00, 32'h4218b7db} /* (26, 3, 23) {real, imag} */,
  {32'hc21c87df, 32'hc0c00d9c} /* (26, 3, 22) {real, imag} */,
  {32'h41ecc7f8, 32'h42b3e3ee} /* (26, 3, 21) {real, imag} */,
  {32'h427175f0, 32'hc1942454} /* (26, 3, 20) {real, imag} */,
  {32'hc1d9206a, 32'hc195b173} /* (26, 3, 19) {real, imag} */,
  {32'hc213b9e3, 32'hc2462d6f} /* (26, 3, 18) {real, imag} */,
  {32'h4161ef60, 32'hc18423c2} /* (26, 3, 17) {real, imag} */,
  {32'h41981d48, 32'h416e20c0} /* (26, 3, 16) {real, imag} */,
  {32'h41b50ec8, 32'h41820322} /* (26, 3, 15) {real, imag} */,
  {32'h4236a2d9, 32'hc14424ec} /* (26, 3, 14) {real, imag} */,
  {32'h4280b83a, 32'hc1dc0a11} /* (26, 3, 13) {real, imag} */,
  {32'h40cf4e00, 32'hc25224ee} /* (26, 3, 12) {real, imag} */,
  {32'h42957154, 32'h42adf11e} /* (26, 3, 11) {real, imag} */,
  {32'hc1a804ca, 32'h41e50a87} /* (26, 3, 10) {real, imag} */,
  {32'hc2a9c4c3, 32'h4298a246} /* (26, 3, 9) {real, imag} */,
  {32'hc196c656, 32'hc277e689} /* (26, 3, 8) {real, imag} */,
  {32'hc29da278, 32'hbeab6e80} /* (26, 3, 7) {real, imag} */,
  {32'h413b0eb7, 32'hc26a95e9} /* (26, 3, 6) {real, imag} */,
  {32'hc1596b68, 32'h424ffc16} /* (26, 3, 5) {real, imag} */,
  {32'hc2a104c9, 32'hc1ff8df9} /* (26, 3, 4) {real, imag} */,
  {32'h43137c73, 32'hc1f2db98} /* (26, 3, 3) {real, imag} */,
  {32'h4272ae35, 32'hc305d78c} /* (26, 3, 2) {real, imag} */,
  {32'hc1dd365a, 32'h432ad81c} /* (26, 3, 1) {real, imag} */,
  {32'h4326ee31, 32'h4381c499} /* (26, 3, 0) {real, imag} */,
  {32'hc303c69d, 32'hc26fbfcc} /* (26, 2, 31) {real, imag} */,
  {32'h431c9cab, 32'h43468f0c} /* (26, 2, 30) {real, imag} */,
  {32'hc271957a, 32'hc3271b62} /* (26, 2, 29) {real, imag} */,
  {32'h424ccdd4, 32'h431abf3f} /* (26, 2, 28) {real, imag} */,
  {32'hc308ad48, 32'hc2f6a060} /* (26, 2, 27) {real, imag} */,
  {32'h41ac2c82, 32'h42dc7962} /* (26, 2, 26) {real, imag} */,
  {32'h4118ec0a, 32'h411d7e22} /* (26, 2, 25) {real, imag} */,
  {32'h422fca05, 32'hc28f1703} /* (26, 2, 24) {real, imag} */,
  {32'h41be1ae8, 32'hbe88d080} /* (26, 2, 23) {real, imag} */,
  {32'hc2d11bfc, 32'h423123ee} /* (26, 2, 22) {real, imag} */,
  {32'h41481a1e, 32'hc013c090} /* (26, 2, 21) {real, imag} */,
  {32'h40d9d4b0, 32'h4248bc37} /* (26, 2, 20) {real, imag} */,
  {32'hc05b52e0, 32'hc17439a6} /* (26, 2, 19) {real, imag} */,
  {32'hbec337e0, 32'h4087b930} /* (26, 2, 18) {real, imag} */,
  {32'hc207a8a4, 32'hc1a0a31d} /* (26, 2, 17) {real, imag} */,
  {32'hc142977c, 32'h410f9ce5} /* (26, 2, 16) {real, imag} */,
  {32'hc1a6bd99, 32'h4106b126} /* (26, 2, 15) {real, imag} */,
  {32'hc18a2c88, 32'h40e42b00} /* (26, 2, 14) {real, imag} */,
  {32'h40f4e900, 32'h423d9284} /* (26, 2, 13) {real, imag} */,
  {32'hc2b33d81, 32'hc2657099} /* (26, 2, 12) {real, imag} */,
  {32'h3eb19cc0, 32'hc1e9d8ec} /* (26, 2, 11) {real, imag} */,
  {32'hc26b8b98, 32'hbeb1b800} /* (26, 2, 10) {real, imag} */,
  {32'hc2aac1f8, 32'h420df8c7} /* (26, 2, 9) {real, imag} */,
  {32'h4055b010, 32'hc280e5f5} /* (26, 2, 8) {real, imag} */,
  {32'hc1011cf2, 32'hc13c8158} /* (26, 2, 7) {real, imag} */,
  {32'hc25575f7, 32'h41b103ea} /* (26, 2, 6) {real, imag} */,
  {32'h413fa3e8, 32'h41d0f7b0} /* (26, 2, 5) {real, imag} */,
  {32'hc28a67bc, 32'hc2b98626} /* (26, 2, 4) {real, imag} */,
  {32'h43011daa, 32'h41f9ae84} /* (26, 2, 3) {real, imag} */,
  {32'h43019375, 32'hc1cbc0d0} /* (26, 2, 2) {real, imag} */,
  {32'h4343ff21, 32'hc2165ac8} /* (26, 2, 1) {real, imag} */,
  {32'hc2a9ccda, 32'h41ffc3ac} /* (26, 2, 0) {real, imag} */,
  {32'hc11e9c5c, 32'h421dae86} /* (26, 1, 31) {real, imag} */,
  {32'h4329e720, 32'hc3048c46} /* (26, 1, 30) {real, imag} */,
  {32'h417d1ae0, 32'h4346ae4b} /* (26, 1, 29) {real, imag} */,
  {32'hc308893e, 32'hc342d98b} /* (26, 1, 28) {real, imag} */,
  {32'h4219c744, 32'hc262d42a} /* (26, 1, 27) {real, imag} */,
  {32'hc2939ef8, 32'h42c4e475} /* (26, 1, 26) {real, imag} */,
  {32'hc2628391, 32'hc2a78f95} /* (26, 1, 25) {real, imag} */,
  {32'h41bfc8a0, 32'h4200fc9e} /* (26, 1, 24) {real, imag} */,
  {32'h42b4689b, 32'hc24eab70} /* (26, 1, 23) {real, imag} */,
  {32'hc228b494, 32'hc153b20c} /* (26, 1, 22) {real, imag} */,
  {32'hc2809a5c, 32'hc0256578} /* (26, 1, 21) {real, imag} */,
  {32'h4295daa0, 32'hc23e729b} /* (26, 1, 20) {real, imag} */,
  {32'hc19097d4, 32'hc18e7a80} /* (26, 1, 19) {real, imag} */,
  {32'h41afb06c, 32'h41d6d750} /* (26, 1, 18) {real, imag} */,
  {32'h412d7dd2, 32'h40369c30} /* (26, 1, 17) {real, imag} */,
  {32'hc02dc500, 32'hc0cf959c} /* (26, 1, 16) {real, imag} */,
  {32'hc0f0e674, 32'h423f0933} /* (26, 1, 15) {real, imag} */,
  {32'h408b75b0, 32'hc0719e40} /* (26, 1, 14) {real, imag} */,
  {32'h425f0898, 32'hc27b5aa0} /* (26, 1, 13) {real, imag} */,
  {32'hc12ee552, 32'h425e6bd7} /* (26, 1, 12) {real, imag} */,
  {32'hc1c13c55, 32'hc200ae90} /* (26, 1, 11) {real, imag} */,
  {32'hc27e0c18, 32'hc1be40d6} /* (26, 1, 10) {real, imag} */,
  {32'h4284c2c1, 32'h40253b28} /* (26, 1, 9) {real, imag} */,
  {32'hc292d368, 32'h425bf6e2} /* (26, 1, 8) {real, imag} */,
  {32'h42a5fbd2, 32'hc218b9a0} /* (26, 1, 7) {real, imag} */,
  {32'hc18df0c8, 32'h42a58267} /* (26, 1, 6) {real, imag} */,
  {32'hc118ef4a, 32'hc1c616cb} /* (26, 1, 5) {real, imag} */,
  {32'hc1e3de64, 32'hc3144d31} /* (26, 1, 4) {real, imag} */,
  {32'h43894f81, 32'hc21e08c4} /* (26, 1, 3) {real, imag} */,
  {32'hc1cd20b4, 32'h42811892} /* (26, 1, 2) {real, imag} */,
  {32'hc2ba0944, 32'h423ee0cc} /* (26, 1, 1) {real, imag} */,
  {32'hc3445530, 32'h41254cf2} /* (26, 1, 0) {real, imag} */,
  {32'h42a2d7b4, 32'hc1da6e2c} /* (26, 0, 31) {real, imag} */,
  {32'h43032f8c, 32'hc3190e1a} /* (26, 0, 30) {real, imag} */,
  {32'h40bb580c, 32'hc248509a} /* (26, 0, 29) {real, imag} */,
  {32'hc28643ce, 32'h42e9fe29} /* (26, 0, 28) {real, imag} */,
  {32'hc2206d6c, 32'h42c191f8} /* (26, 0, 27) {real, imag} */,
  {32'hc16fcdc3, 32'hc237dc02} /* (26, 0, 26) {real, imag} */,
  {32'h430f513c, 32'h428418f9} /* (26, 0, 25) {real, imag} */,
  {32'hc200407b, 32'h41b1c3d6} /* (26, 0, 24) {real, imag} */,
  {32'hc1cdb552, 32'h420ef86e} /* (26, 0, 23) {real, imag} */,
  {32'hc1edf7b0, 32'h4282d82a} /* (26, 0, 22) {real, imag} */,
  {32'h417d39d2, 32'h42992cf0} /* (26, 0, 21) {real, imag} */,
  {32'h411a783a, 32'h421c3bf8} /* (26, 0, 20) {real, imag} */,
  {32'hc28754ee, 32'h421f5bf5} /* (26, 0, 19) {real, imag} */,
  {32'h41eb8440, 32'hc25a9b0a} /* (26, 0, 18) {real, imag} */,
  {32'hc13c41e9, 32'h4158cf82} /* (26, 0, 17) {real, imag} */,
  {32'hc12f5960, 32'hc2413338} /* (26, 0, 16) {real, imag} */,
  {32'hc21ef45a, 32'hc0b98b44} /* (26, 0, 15) {real, imag} */,
  {32'hc20b356e, 32'hc095610c} /* (26, 0, 14) {real, imag} */,
  {32'h41720f14, 32'hc1e8650e} /* (26, 0, 13) {real, imag} */,
  {32'h41ac2b19, 32'hc0ec76c0} /* (26, 0, 12) {real, imag} */,
  {32'hc18fe117, 32'h414143fc} /* (26, 0, 11) {real, imag} */,
  {32'h4238e124, 32'hc22cb708} /* (26, 0, 10) {real, imag} */,
  {32'hc23b7fa3, 32'hc1bdcd57} /* (26, 0, 9) {real, imag} */,
  {32'hc1d6dc20, 32'h43042b3b} /* (26, 0, 8) {real, imag} */,
  {32'h4216a6b1, 32'h4228c00e} /* (26, 0, 7) {real, imag} */,
  {32'h40ad4b82, 32'hc245f82a} /* (26, 0, 6) {real, imag} */,
  {32'h42f2124e, 32'hc3668418} /* (26, 0, 5) {real, imag} */,
  {32'hc1ede04a, 32'h42cf0dfb} /* (26, 0, 4) {real, imag} */,
  {32'h406c0b08, 32'hbfa35f10} /* (26, 0, 3) {real, imag} */,
  {32'hc31994a6, 32'h419f5cf8} /* (26, 0, 2) {real, imag} */,
  {32'h41765170, 32'hc3033c94} /* (26, 0, 1) {real, imag} */,
  {32'h43269c08, 32'hc3154c58} /* (26, 0, 0) {real, imag} */,
  {32'h42ec4ca6, 32'h42c32d6d} /* (25, 31, 31) {real, imag} */,
  {32'hc2a0358f, 32'hc301b7aa} /* (25, 31, 30) {real, imag} */,
  {32'hc02d1b90, 32'h42fd06ee} /* (25, 31, 29) {real, imag} */,
  {32'h3f9e3700, 32'hc02f0630} /* (25, 31, 28) {real, imag} */,
  {32'hc1b061d8, 32'h42117e2c} /* (25, 31, 27) {real, imag} */,
  {32'h42c3709e, 32'h43353dff} /* (25, 31, 26) {real, imag} */,
  {32'h3f800a10, 32'hc23c20ce} /* (25, 31, 25) {real, imag} */,
  {32'hc208bac0, 32'h40f9aa44} /* (25, 31, 24) {real, imag} */,
  {32'h41483e92, 32'h40025520} /* (25, 31, 23) {real, imag} */,
  {32'hc29aed44, 32'h41e7ce1c} /* (25, 31, 22) {real, imag} */,
  {32'hc1b01b7c, 32'h4274c4d6} /* (25, 31, 21) {real, imag} */,
  {32'h3f78e9a0, 32'hc1ce10f1} /* (25, 31, 20) {real, imag} */,
  {32'h41dab7ba, 32'hc12684a7} /* (25, 31, 19) {real, imag} */,
  {32'h402a5078, 32'h41eea7ea} /* (25, 31, 18) {real, imag} */,
  {32'hc141eed4, 32'hc15ea396} /* (25, 31, 17) {real, imag} */,
  {32'h41428859, 32'h4110be90} /* (25, 31, 16) {real, imag} */,
  {32'hc11750b0, 32'hc1af309d} /* (25, 31, 15) {real, imag} */,
  {32'hc21dd2d8, 32'hc191527e} /* (25, 31, 14) {real, imag} */,
  {32'h41b77432, 32'h4222f05a} /* (25, 31, 13) {real, imag} */,
  {32'hc1f47c65, 32'hc20c0adc} /* (25, 31, 12) {real, imag} */,
  {32'hc2220bea, 32'h41fc9ccc} /* (25, 31, 11) {real, imag} */,
  {32'hc2ce2264, 32'hc200ba76} /* (25, 31, 10) {real, imag} */,
  {32'h4219c5d6, 32'h42e27a43} /* (25, 31, 9) {real, imag} */,
  {32'h41a2d690, 32'h423f3b32} /* (25, 31, 8) {real, imag} */,
  {32'h42407654, 32'hc3062b76} /* (25, 31, 7) {real, imag} */,
  {32'h41eb5192, 32'hc1b31e20} /* (25, 31, 6) {real, imag} */,
  {32'h42931f80, 32'hc32b2d34} /* (25, 31, 5) {real, imag} */,
  {32'h42d027e4, 32'h42071b6c} /* (25, 31, 4) {real, imag} */,
  {32'h411ad04c, 32'hc2547754} /* (25, 31, 3) {real, imag} */,
  {32'hc31d11ac, 32'hc2ea6605} /* (25, 31, 2) {real, imag} */,
  {32'h4034e640, 32'h433ecf0a} /* (25, 31, 1) {real, imag} */,
  {32'h41b99dbc, 32'hc2b71f40} /* (25, 31, 0) {real, imag} */,
  {32'hc1bb9d90, 32'hc237db81} /* (25, 30, 31) {real, imag} */,
  {32'hc2c99cb9, 32'h428b8c5b} /* (25, 30, 30) {real, imag} */,
  {32'h42cd81c2, 32'h4100a6a8} /* (25, 30, 29) {real, imag} */,
  {32'h421fc913, 32'h41e1c354} /* (25, 30, 28) {real, imag} */,
  {32'h42c5d0da, 32'h4227de53} /* (25, 30, 27) {real, imag} */,
  {32'hc2343a4c, 32'hc20ce592} /* (25, 30, 26) {real, imag} */,
  {32'h41e3c286, 32'h4031fd80} /* (25, 30, 25) {real, imag} */,
  {32'h4202cffd, 32'hbfb76c80} /* (25, 30, 24) {real, imag} */,
  {32'h42b8c266, 32'hc0ce0ed4} /* (25, 30, 23) {real, imag} */,
  {32'hc2958478, 32'h3f9ee308} /* (25, 30, 22) {real, imag} */,
  {32'hc2bf9607, 32'h4220dc4c} /* (25, 30, 21) {real, imag} */,
  {32'h4200f1e0, 32'hc1393ab8} /* (25, 30, 20) {real, imag} */,
  {32'hc0cdc688, 32'hc109f74c} /* (25, 30, 19) {real, imag} */,
  {32'h41cfccf3, 32'hc0a22870} /* (25, 30, 18) {real, imag} */,
  {32'hbfa204a0, 32'hc06c4238} /* (25, 30, 17) {real, imag} */,
  {32'h40ce8078, 32'h41a397d6} /* (25, 30, 16) {real, imag} */,
  {32'h4153272c, 32'hc259f6e0} /* (25, 30, 15) {real, imag} */,
  {32'h40b57d54, 32'h41df3f04} /* (25, 30, 14) {real, imag} */,
  {32'hc0d34908, 32'hc18e99e2} /* (25, 30, 13) {real, imag} */,
  {32'h420adb56, 32'hc1595080} /* (25, 30, 12) {real, imag} */,
  {32'hc275f3da, 32'h412258c2} /* (25, 30, 11) {real, imag} */,
  {32'hc213f83b, 32'hc1a25ab4} /* (25, 30, 10) {real, imag} */,
  {32'h421dada7, 32'hc16759f6} /* (25, 30, 9) {real, imag} */,
  {32'h420d7d67, 32'h42e409c4} /* (25, 30, 8) {real, imag} */,
  {32'h410ec2df, 32'hc2a3d740} /* (25, 30, 7) {real, imag} */,
  {32'hc20e291c, 32'hc1a8fb68} /* (25, 30, 6) {real, imag} */,
  {32'hc296a798, 32'hc2507405} /* (25, 30, 5) {real, imag} */,
  {32'h42d09552, 32'h430b6f48} /* (25, 30, 4) {real, imag} */,
  {32'hc334bebd, 32'h43105a04} /* (25, 30, 3) {real, imag} */,
  {32'hc241b95e, 32'h431b23dc} /* (25, 30, 2) {real, imag} */,
  {32'hc2929622, 32'hc296d9d6} /* (25, 30, 1) {real, imag} */,
  {32'hc1ce5884, 32'hc296d556} /* (25, 30, 0) {real, imag} */,
  {32'h42c4aa18, 32'hc1b14728} /* (25, 29, 31) {real, imag} */,
  {32'h4224fc64, 32'h422e8cd2} /* (25, 29, 30) {real, imag} */,
  {32'h431b503a, 32'hc0837770} /* (25, 29, 29) {real, imag} */,
  {32'h42c9a06e, 32'h405bfb30} /* (25, 29, 28) {real, imag} */,
  {32'hc27fd0fa, 32'h42ded6f2} /* (25, 29, 27) {real, imag} */,
  {32'hc28e97ee, 32'hc28995a0} /* (25, 29, 26) {real, imag} */,
  {32'hc2db5520, 32'hc1721377} /* (25, 29, 25) {real, imag} */,
  {32'h410367c6, 32'hc1d88aa6} /* (25, 29, 24) {real, imag} */,
  {32'h40fc1a6c, 32'h42a45821} /* (25, 29, 23) {real, imag} */,
  {32'h412e9182, 32'h420e196f} /* (25, 29, 22) {real, imag} */,
  {32'h4242b5d0, 32'h40b7b212} /* (25, 29, 21) {real, imag} */,
  {32'h4194d8c8, 32'h42444cd2} /* (25, 29, 20) {real, imag} */,
  {32'hc0341bc0, 32'hc0a1d470} /* (25, 29, 19) {real, imag} */,
  {32'hc29191ea, 32'h41be09c5} /* (25, 29, 18) {real, imag} */,
  {32'h418d29a0, 32'h40be3104} /* (25, 29, 17) {real, imag} */,
  {32'hc146bcb4, 32'h410877e4} /* (25, 29, 16) {real, imag} */,
  {32'hc126d720, 32'h4161a9ba} /* (25, 29, 15) {real, imag} */,
  {32'h417b285e, 32'h4129b086} /* (25, 29, 14) {real, imag} */,
  {32'hc136f168, 32'hc262535e} /* (25, 29, 13) {real, imag} */,
  {32'h426d1722, 32'h42b77543} /* (25, 29, 12) {real, imag} */,
  {32'hc0a66624, 32'h41a67e48} /* (25, 29, 11) {real, imag} */,
  {32'hc16e62ae, 32'hc21032db} /* (25, 29, 10) {real, imag} */,
  {32'h41f59291, 32'hc2ab50b3} /* (25, 29, 9) {real, imag} */,
  {32'h423091da, 32'h40f51d78} /* (25, 29, 8) {real, imag} */,
  {32'h421a004b, 32'h41ac9004} /* (25, 29, 7) {real, imag} */,
  {32'h42111a89, 32'h42851798} /* (25, 29, 6) {real, imag} */,
  {32'h4048ad38, 32'h424bc853} /* (25, 29, 5) {real, imag} */,
  {32'hc151b128, 32'h428d6148} /* (25, 29, 4) {real, imag} */,
  {32'hc05ba800, 32'hc329be72} /* (25, 29, 3) {real, imag} */,
  {32'h40b27b18, 32'hc29ea427} /* (25, 29, 2) {real, imag} */,
  {32'hc3201888, 32'h42f8eeee} /* (25, 29, 1) {real, imag} */,
  {32'h42d417a4, 32'hc143a364} /* (25, 29, 0) {real, imag} */,
  {32'hc1398d50, 32'hc2845640} /* (25, 28, 31) {real, imag} */,
  {32'h42377488, 32'h434348cd} /* (25, 28, 30) {real, imag} */,
  {32'hc2a1a316, 32'hc2adbab6} /* (25, 28, 29) {real, imag} */,
  {32'h43125308, 32'h3df5f800} /* (25, 28, 28) {real, imag} */,
  {32'h4205512d, 32'hc210005c} /* (25, 28, 27) {real, imag} */,
  {32'h4196a86e, 32'hc26d9b96} /* (25, 28, 26) {real, imag} */,
  {32'hc2a0453f, 32'h420d4fa2} /* (25, 28, 25) {real, imag} */,
  {32'h4284a245, 32'hc2809042} /* (25, 28, 24) {real, imag} */,
  {32'hc21f7322, 32'h424490d4} /* (25, 28, 23) {real, imag} */,
  {32'h40e2dc9a, 32'h41ccdcca} /* (25, 28, 22) {real, imag} */,
  {32'h41b64fbc, 32'hc24da62d} /* (25, 28, 21) {real, imag} */,
  {32'h41c7de24, 32'h4203a2fd} /* (25, 28, 20) {real, imag} */,
  {32'hc284e363, 32'h41824ace} /* (25, 28, 19) {real, imag} */,
  {32'h40f4f8d6, 32'hc2120ba5} /* (25, 28, 18) {real, imag} */,
  {32'h40af059e, 32'h3ffd78b8} /* (25, 28, 17) {real, imag} */,
  {32'h40d56778, 32'hc0edf990} /* (25, 28, 16) {real, imag} */,
  {32'hc0830b72, 32'h418f1e90} /* (25, 28, 15) {real, imag} */,
  {32'hc16ee2ab, 32'hc2598035} /* (25, 28, 14) {real, imag} */,
  {32'hc1ab9bbf, 32'h4030f5d0} /* (25, 28, 13) {real, imag} */,
  {32'h41070858, 32'hc0746d50} /* (25, 28, 12) {real, imag} */,
  {32'hc28f57b6, 32'h421ecf2f} /* (25, 28, 11) {real, imag} */,
  {32'hc19e21d6, 32'hc29b51f6} /* (25, 28, 10) {real, imag} */,
  {32'hbfb2c4d0, 32'hbecb5b00} /* (25, 28, 9) {real, imag} */,
  {32'h428bc923, 32'hc24f6af5} /* (25, 28, 8) {real, imag} */,
  {32'h41bc0f8d, 32'hc245dfec} /* (25, 28, 7) {real, imag} */,
  {32'hc22b3f4f, 32'hc25f8920} /* (25, 28, 6) {real, imag} */,
  {32'h42cfacde, 32'h42a65582} /* (25, 28, 5) {real, imag} */,
  {32'hc281663d, 32'hc2b6e1fd} /* (25, 28, 4) {real, imag} */,
  {32'hc1cbb34b, 32'h428d1142} /* (25, 28, 3) {real, imag} */,
  {32'h42bc43dc, 32'h42f78532} /* (25, 28, 2) {real, imag} */,
  {32'h423a873a, 32'h4252407e} /* (25, 28, 1) {real, imag} */,
  {32'hc18193fa, 32'hc2860847} /* (25, 28, 0) {real, imag} */,
  {32'hc257cfd4, 32'h41c12c68} /* (25, 27, 31) {real, imag} */,
  {32'hc2a949ee, 32'hc2a82804} /* (25, 27, 30) {real, imag} */,
  {32'hc1e4439a, 32'h42a45bb0} /* (25, 27, 29) {real, imag} */,
  {32'h421b1c45, 32'hc2524124} /* (25, 27, 28) {real, imag} */,
  {32'hc1c15832, 32'hc203d18a} /* (25, 27, 27) {real, imag} */,
  {32'hc27e0bc2, 32'hc1830c45} /* (25, 27, 26) {real, imag} */,
  {32'h42806e24, 32'h42987fd0} /* (25, 27, 25) {real, imag} */,
  {32'h418ed835, 32'hc220e866} /* (25, 27, 24) {real, imag} */,
  {32'h4020e7d0, 32'hc2910c2c} /* (25, 27, 23) {real, imag} */,
  {32'hc12d6317, 32'hc2d46114} /* (25, 27, 22) {real, imag} */,
  {32'hbf78fe00, 32'h423d919a} /* (25, 27, 21) {real, imag} */,
  {32'h410d3fb4, 32'h41ced78c} /* (25, 27, 20) {real, imag} */,
  {32'h418ada58, 32'h41898e7a} /* (25, 27, 19) {real, imag} */,
  {32'h4187ac8c, 32'hc0b9ecd0} /* (25, 27, 18) {real, imag} */,
  {32'h41b023d6, 32'h414f0be8} /* (25, 27, 17) {real, imag} */,
  {32'h41b24586, 32'hc0333840} /* (25, 27, 16) {real, imag} */,
  {32'h4049c6a0, 32'hc16721e4} /* (25, 27, 15) {real, imag} */,
  {32'h42620042, 32'hc1a895d4} /* (25, 27, 14) {real, imag} */,
  {32'hc285f885, 32'hc11e6e5b} /* (25, 27, 13) {real, imag} */,
  {32'hc200db85, 32'h41308654} /* (25, 27, 12) {real, imag} */,
  {32'hc211b5f2, 32'h41895634} /* (25, 27, 11) {real, imag} */,
  {32'h4158062f, 32'hc0e599f8} /* (25, 27, 10) {real, imag} */,
  {32'h428eddf4, 32'hc2896408} /* (25, 27, 9) {real, imag} */,
  {32'hc09ce4dc, 32'h41fc68d8} /* (25, 27, 8) {real, imag} */,
  {32'h4272f743, 32'hc2f32c4c} /* (25, 27, 7) {real, imag} */,
  {32'hc2bb0187, 32'hc1882309} /* (25, 27, 6) {real, imag} */,
  {32'h4302bb40, 32'h429b068b} /* (25, 27, 5) {real, imag} */,
  {32'h41cda316, 32'h4246900c} /* (25, 27, 4) {real, imag} */,
  {32'h420ec3b9, 32'hc14589c4} /* (25, 27, 3) {real, imag} */,
  {32'hc0b50ee8, 32'hc3412296} /* (25, 27, 2) {real, imag} */,
  {32'h422886c4, 32'hc214b73f} /* (25, 27, 1) {real, imag} */,
  {32'h42088cda, 32'h432f2893} /* (25, 27, 0) {real, imag} */,
  {32'h42e4fb1e, 32'hc2518146} /* (25, 26, 31) {real, imag} */,
  {32'hc2130494, 32'h42acdcd0} /* (25, 26, 30) {real, imag} */,
  {32'hc0e85604, 32'h41400248} /* (25, 26, 29) {real, imag} */,
  {32'h4232be16, 32'hc11eb7a4} /* (25, 26, 28) {real, imag} */,
  {32'hc23ad454, 32'h420b2df2} /* (25, 26, 27) {real, imag} */,
  {32'hc11be3b2, 32'h41209d97} /* (25, 26, 26) {real, imag} */,
  {32'hc16f5c30, 32'h4250142a} /* (25, 26, 25) {real, imag} */,
  {32'hc255f4c8, 32'hc23d67af} /* (25, 26, 24) {real, imag} */,
  {32'h41d3dcf4, 32'h424c4746} /* (25, 26, 23) {real, imag} */,
  {32'h41694d62, 32'h41287e03} /* (25, 26, 22) {real, imag} */,
  {32'hbe469f00, 32'hc2475580} /* (25, 26, 21) {real, imag} */,
  {32'h3e4336e0, 32'h418abf6e} /* (25, 26, 20) {real, imag} */,
  {32'h40668f18, 32'hc239c0e8} /* (25, 26, 19) {real, imag} */,
  {32'h41384b1a, 32'h40b378dc} /* (25, 26, 18) {real, imag} */,
  {32'h40c2a1bc, 32'hc0cbe7e4} /* (25, 26, 17) {real, imag} */,
  {32'h40906562, 32'h41010908} /* (25, 26, 16) {real, imag} */,
  {32'hc03f2688, 32'hc1a5723f} /* (25, 26, 15) {real, imag} */,
  {32'hc07f5098, 32'h40ce5994} /* (25, 26, 14) {real, imag} */,
  {32'hc1740330, 32'h41f0bbb8} /* (25, 26, 13) {real, imag} */,
  {32'h4049a1e2, 32'h41b2387c} /* (25, 26, 12) {real, imag} */,
  {32'h4229f85e, 32'hc245ca18} /* (25, 26, 11) {real, imag} */,
  {32'hc27f4c3c, 32'hc1d438c8} /* (25, 26, 10) {real, imag} */,
  {32'h4233a1e8, 32'hbec671c0} /* (25, 26, 9) {real, imag} */,
  {32'hc1f40c7f, 32'hc1a30c7a} /* (25, 26, 8) {real, imag} */,
  {32'h428c2edb, 32'h418c1e8c} /* (25, 26, 7) {real, imag} */,
  {32'hc228169c, 32'hbf3b9ad0} /* (25, 26, 6) {real, imag} */,
  {32'hc270be24, 32'hc28fb517} /* (25, 26, 5) {real, imag} */,
  {32'h41333f76, 32'hc22cba60} /* (25, 26, 4) {real, imag} */,
  {32'h417ac1a4, 32'hc2af5495} /* (25, 26, 3) {real, imag} */,
  {32'h42eb1db2, 32'hc1696b34} /* (25, 26, 2) {real, imag} */,
  {32'hc24d8314, 32'h42552aee} /* (25, 26, 1) {real, imag} */,
  {32'hc107f0f1, 32'h41b4e87a} /* (25, 26, 0) {real, imag} */,
  {32'h427f4b9e, 32'h41eed3ae} /* (25, 25, 31) {real, imag} */,
  {32'h420c1205, 32'hc21cf3ac} /* (25, 25, 30) {real, imag} */,
  {32'hc2a5015f, 32'hc18069fc} /* (25, 25, 29) {real, imag} */,
  {32'hc1d655d2, 32'h41cc4223} /* (25, 25, 28) {real, imag} */,
  {32'h412c1ada, 32'hc2a2b879} /* (25, 25, 27) {real, imag} */,
  {32'h406f2bc0, 32'hc2517588} /* (25, 25, 26) {real, imag} */,
  {32'h4239b460, 32'hbffe3740} /* (25, 25, 25) {real, imag} */,
  {32'h416b99c5, 32'h42048056} /* (25, 25, 24) {real, imag} */,
  {32'hc20bf601, 32'h425cde86} /* (25, 25, 23) {real, imag} */,
  {32'hc06f3960, 32'h408f0e54} /* (25, 25, 22) {real, imag} */,
  {32'hbf820b48, 32'hc15dde48} /* (25, 25, 21) {real, imag} */,
  {32'hc18d6ff6, 32'hc0c42a1b} /* (25, 25, 20) {real, imag} */,
  {32'h41b8cc51, 32'h4147207c} /* (25, 25, 19) {real, imag} */,
  {32'hbf9028a8, 32'h4136ab2a} /* (25, 25, 18) {real, imag} */,
  {32'h416fd351, 32'hc1844b7d} /* (25, 25, 17) {real, imag} */,
  {32'h411b2104, 32'hbe2d2480} /* (25, 25, 16) {real, imag} */,
  {32'h415651e9, 32'h40ff13f0} /* (25, 25, 15) {real, imag} */,
  {32'hc0730b3c, 32'hc1dce655} /* (25, 25, 14) {real, imag} */,
  {32'hc12127da, 32'h40c90980} /* (25, 25, 13) {real, imag} */,
  {32'h42135472, 32'h415cd62c} /* (25, 25, 12) {real, imag} */,
  {32'h41f25708, 32'hc238cf61} /* (25, 25, 11) {real, imag} */,
  {32'h421f2f5c, 32'h41fc6e57} /* (25, 25, 10) {real, imag} */,
  {32'h4109a35d, 32'hc1dc2670} /* (25, 25, 9) {real, imag} */,
  {32'hc1169533, 32'h410bb20e} /* (25, 25, 8) {real, imag} */,
  {32'h40a086c0, 32'h426dc29c} /* (25, 25, 7) {real, imag} */,
  {32'hc260250e, 32'h3f9e5ab0} /* (25, 25, 6) {real, imag} */,
  {32'hc1d4d63f, 32'hc1786768} /* (25, 25, 5) {real, imag} */,
  {32'h41865250, 32'hc19fd755} /* (25, 25, 4) {real, imag} */,
  {32'h4290d327, 32'hc2a2cbdf} /* (25, 25, 3) {real, imag} */,
  {32'h4241133b, 32'hc2a99d5e} /* (25, 25, 2) {real, imag} */,
  {32'h419f8a0f, 32'h418baff2} /* (25, 25, 1) {real, imag} */,
  {32'hc26c780b, 32'h41ff7e4b} /* (25, 25, 0) {real, imag} */,
  {32'hc26b92eb, 32'h42939665} /* (25, 24, 31) {real, imag} */,
  {32'hc1b16025, 32'h426afe4a} /* (25, 24, 30) {real, imag} */,
  {32'hbee1ab80, 32'hc0924bf0} /* (25, 24, 29) {real, imag} */,
  {32'h427ae4b4, 32'hc21683d8} /* (25, 24, 28) {real, imag} */,
  {32'hc2216e82, 32'hc1cfe117} /* (25, 24, 27) {real, imag} */,
  {32'h41fe6904, 32'hc17803b0} /* (25, 24, 26) {real, imag} */,
  {32'h42a4c1d5, 32'hc14f3adb} /* (25, 24, 25) {real, imag} */,
  {32'h413b9776, 32'h4091299a} /* (25, 24, 24) {real, imag} */,
  {32'h4270a90d, 32'hc251f2ac} /* (25, 24, 23) {real, imag} */,
  {32'h41bf8104, 32'h4209a6a6} /* (25, 24, 22) {real, imag} */,
  {32'h429716a8, 32'hc0e6d094} /* (25, 24, 21) {real, imag} */,
  {32'hc2353cdf, 32'hc0101984} /* (25, 24, 20) {real, imag} */,
  {32'hc04ac420, 32'h413944ad} /* (25, 24, 19) {real, imag} */,
  {32'hc0bc2c00, 32'hc164a4ec} /* (25, 24, 18) {real, imag} */,
  {32'hc0cbc1b2, 32'h41dfff51} /* (25, 24, 17) {real, imag} */,
  {32'hbf9ff068, 32'h417f6078} /* (25, 24, 16) {real, imag} */,
  {32'hc1dab7a8, 32'hc091f1ac} /* (25, 24, 15) {real, imag} */,
  {32'hc0980da0, 32'h411ef33e} /* (25, 24, 14) {real, imag} */,
  {32'h41a36af4, 32'hc0bdb83a} /* (25, 24, 13) {real, imag} */,
  {32'h40c49170, 32'h411e8159} /* (25, 24, 12) {real, imag} */,
  {32'hc1501102, 32'hc04d86f8} /* (25, 24, 11) {real, imag} */,
  {32'hc1ccf904, 32'h422194ce} /* (25, 24, 10) {real, imag} */,
  {32'hc28dbcb1, 32'h417e8498} /* (25, 24, 9) {real, imag} */,
  {32'hc1e1205f, 32'hc1679929} /* (25, 24, 8) {real, imag} */,
  {32'hc23c6546, 32'h41195a2d} /* (25, 24, 7) {real, imag} */,
  {32'h41490317, 32'h42b23c74} /* (25, 24, 6) {real, imag} */,
  {32'h421e587a, 32'hc28795e1} /* (25, 24, 5) {real, imag} */,
  {32'hc15d0036, 32'hc2a4e5a2} /* (25, 24, 4) {real, imag} */,
  {32'h42c2a9c4, 32'h40edf230} /* (25, 24, 3) {real, imag} */,
  {32'hc20e0fe0, 32'hc1ad1850} /* (25, 24, 2) {real, imag} */,
  {32'hc0d96468, 32'hc1f39e8f} /* (25, 24, 1) {real, imag} */,
  {32'h41a40ae6, 32'hc2d0a42f} /* (25, 24, 0) {real, imag} */,
  {32'h421071f3, 32'hc206df18} /* (25, 23, 31) {real, imag} */,
  {32'h4309ecae, 32'hc10d9412} /* (25, 23, 30) {real, imag} */,
  {32'h3fb493a8, 32'hc1686ada} /* (25, 23, 29) {real, imag} */,
  {32'hc1bcd469, 32'hc1db5a9e} /* (25, 23, 28) {real, imag} */,
  {32'hc04abb94, 32'h40de5dec} /* (25, 23, 27) {real, imag} */,
  {32'hc1dde8a4, 32'h4294ffb4} /* (25, 23, 26) {real, imag} */,
  {32'hc22bc2da, 32'hc2c96720} /* (25, 23, 25) {real, imag} */,
  {32'h4203f548, 32'hc1ae53c3} /* (25, 23, 24) {real, imag} */,
  {32'hc0f99b0e, 32'h42732a5f} /* (25, 23, 23) {real, imag} */,
  {32'h421fa698, 32'hc248883c} /* (25, 23, 22) {real, imag} */,
  {32'hc1ddeb6e, 32'h414b1e71} /* (25, 23, 21) {real, imag} */,
  {32'h41561d57, 32'hc09a434a} /* (25, 23, 20) {real, imag} */,
  {32'h41b48e4a, 32'h40a6e8f7} /* (25, 23, 19) {real, imag} */,
  {32'h40a1e674, 32'hc140654a} /* (25, 23, 18) {real, imag} */,
  {32'h4088190a, 32'h41213ed9} /* (25, 23, 17) {real, imag} */,
  {32'h4090844e, 32'h414320b6} /* (25, 23, 16) {real, imag} */,
  {32'hc1109bfd, 32'hc191198c} /* (25, 23, 15) {real, imag} */,
  {32'h4108f466, 32'h41958cdd} /* (25, 23, 14) {real, imag} */,
  {32'h41902bca, 32'h418e58fb} /* (25, 23, 13) {real, imag} */,
  {32'hc14b462b, 32'hc08bab3a} /* (25, 23, 12) {real, imag} */,
  {32'hc21fadc1, 32'hc1628df9} /* (25, 23, 11) {real, imag} */,
  {32'h422ee60a, 32'hc20556fa} /* (25, 23, 10) {real, imag} */,
  {32'h4192d288, 32'h40fd97f8} /* (25, 23, 9) {real, imag} */,
  {32'hbdc69700, 32'h4201620a} /* (25, 23, 8) {real, imag} */,
  {32'h42919728, 32'hc1668744} /* (25, 23, 7) {real, imag} */,
  {32'hc204cbb8, 32'hc0ebb6f8} /* (25, 23, 6) {real, imag} */,
  {32'hc1a39764, 32'h422f0e74} /* (25, 23, 5) {real, imag} */,
  {32'h424df3b6, 32'h40c4ce78} /* (25, 23, 4) {real, imag} */,
  {32'hc191d520, 32'hc1eb6f4f} /* (25, 23, 3) {real, imag} */,
  {32'h420ebf6e, 32'hc137fa26} /* (25, 23, 2) {real, imag} */,
  {32'h41b07eb6, 32'h42238d28} /* (25, 23, 1) {real, imag} */,
  {32'hc1cc05fe, 32'hc28e87bd} /* (25, 23, 0) {real, imag} */,
  {32'h41464c86, 32'h41d1b83a} /* (25, 22, 31) {real, imag} */,
  {32'h425648a0, 32'hc2721f69} /* (25, 22, 30) {real, imag} */,
  {32'hc0f42ee6, 32'h428b5120} /* (25, 22, 29) {real, imag} */,
  {32'hc229186a, 32'h411de6da} /* (25, 22, 28) {real, imag} */,
  {32'hc1e6b2c4, 32'hc1e7bd35} /* (25, 22, 27) {real, imag} */,
  {32'hc1b66044, 32'hc20a3632} /* (25, 22, 26) {real, imag} */,
  {32'h41b7e89b, 32'hbe8e2200} /* (25, 22, 25) {real, imag} */,
  {32'hc135ac8a, 32'hc1a77e04} /* (25, 22, 24) {real, imag} */,
  {32'hbfe71dac, 32'h4165e120} /* (25, 22, 23) {real, imag} */,
  {32'h40bdb44c, 32'h41f397e8} /* (25, 22, 22) {real, imag} */,
  {32'hc0bddab8, 32'hc01f5428} /* (25, 22, 21) {real, imag} */,
  {32'h41e2f00a, 32'h414cc1ab} /* (25, 22, 20) {real, imag} */,
  {32'hc02d47d8, 32'hc17400ed} /* (25, 22, 19) {real, imag} */,
  {32'hc04a10dc, 32'h412ec5b1} /* (25, 22, 18) {real, imag} */,
  {32'hc112e8f6, 32'hc08d8d1a} /* (25, 22, 17) {real, imag} */,
  {32'hbfc3f680, 32'h4010a4e8} /* (25, 22, 16) {real, imag} */,
  {32'hbef57d20, 32'h41a23cb2} /* (25, 22, 15) {real, imag} */,
  {32'h40822a82, 32'h403eb824} /* (25, 22, 14) {real, imag} */,
  {32'hc21168a4, 32'hc10147b9} /* (25, 22, 13) {real, imag} */,
  {32'hc1d8c330, 32'hc0d941ee} /* (25, 22, 12) {real, imag} */,
  {32'hc1fda5f8, 32'hc1a87907} /* (25, 22, 11) {real, imag} */,
  {32'h421f5a86, 32'h418e4fb4} /* (25, 22, 10) {real, imag} */,
  {32'hc12d5906, 32'h422fd236} /* (25, 22, 9) {real, imag} */,
  {32'h41ba5a0b, 32'hc20baa91} /* (25, 22, 8) {real, imag} */,
  {32'h420644bb, 32'h4243903a} /* (25, 22, 7) {real, imag} */,
  {32'h41738338, 32'hc286653c} /* (25, 22, 6) {real, imag} */,
  {32'h415a5624, 32'hc22088ea} /* (25, 22, 5) {real, imag} */,
  {32'hc2864941, 32'h417d2920} /* (25, 22, 4) {real, imag} */,
  {32'hc1f677c4, 32'hc2781b2c} /* (25, 22, 3) {real, imag} */,
  {32'hc20bc30e, 32'h428b9e77} /* (25, 22, 2) {real, imag} */,
  {32'h40a5aee5, 32'h42021231} /* (25, 22, 1) {real, imag} */,
  {32'h4209ecc9, 32'hc0d3563c} /* (25, 22, 0) {real, imag} */,
  {32'hc29fe0a6, 32'h4250b715} /* (25, 21, 31) {real, imag} */,
  {32'h42832628, 32'h4203d6d8} /* (25, 21, 30) {real, imag} */,
  {32'hc1ae79d7, 32'hc20513d0} /* (25, 21, 29) {real, imag} */,
  {32'hc1b77c58, 32'h413f2d26} /* (25, 21, 28) {real, imag} */,
  {32'hc0fe1ec0, 32'h41985eb8} /* (25, 21, 27) {real, imag} */,
  {32'hc21decbc, 32'hc2165c94} /* (25, 21, 26) {real, imag} */,
  {32'h42773daf, 32'hc105a6a2} /* (25, 21, 25) {real, imag} */,
  {32'h41353d8a, 32'h3e8c5340} /* (25, 21, 24) {real, imag} */,
  {32'hc20aa1cc, 32'hc1653036} /* (25, 21, 23) {real, imag} */,
  {32'hc20a479b, 32'h4121e14a} /* (25, 21, 22) {real, imag} */,
  {32'hc18af38e, 32'h40e1466e} /* (25, 21, 21) {real, imag} */,
  {32'h3ff9418c, 32'h4143cfbc} /* (25, 21, 20) {real, imag} */,
  {32'h414929c4, 32'h420758b6} /* (25, 21, 19) {real, imag} */,
  {32'h41ac02e0, 32'h3f860d24} /* (25, 21, 18) {real, imag} */,
  {32'hc0a36d12, 32'hc183f6ac} /* (25, 21, 17) {real, imag} */,
  {32'h41535fb0, 32'h41197b58} /* (25, 21, 16) {real, imag} */,
  {32'hbf1507f0, 32'h3fd16780} /* (25, 21, 15) {real, imag} */,
  {32'hc0d59bbe, 32'h412a0768} /* (25, 21, 14) {real, imag} */,
  {32'hc11c3938, 32'hc1787e07} /* (25, 21, 13) {real, imag} */,
  {32'h408cbe81, 32'hc19eb756} /* (25, 21, 12) {real, imag} */,
  {32'h40ce0f8a, 32'h400ce7ec} /* (25, 21, 11) {real, imag} */,
  {32'h4149d95c, 32'h40a23d40} /* (25, 21, 10) {real, imag} */,
  {32'hc15cbff7, 32'h426039e0} /* (25, 21, 9) {real, imag} */,
  {32'hc0c15564, 32'h42161ba8} /* (25, 21, 8) {real, imag} */,
  {32'h41e34c9e, 32'h42073c0e} /* (25, 21, 7) {real, imag} */,
  {32'hc00d2d20, 32'h41a22810} /* (25, 21, 6) {real, imag} */,
  {32'h427facfe, 32'hc28678a0} /* (25, 21, 5) {real, imag} */,
  {32'hc08ab05a, 32'hc13c0940} /* (25, 21, 4) {real, imag} */,
  {32'hc253a9bc, 32'hc206cdd6} /* (25, 21, 3) {real, imag} */,
  {32'hc225b693, 32'h42563358} /* (25, 21, 2) {real, imag} */,
  {32'hc2106d0f, 32'hc0973178} /* (25, 21, 1) {real, imag} */,
  {32'hc1997b94, 32'h41ca784a} /* (25, 21, 0) {real, imag} */,
  {32'hc132c174, 32'hc1f35055} /* (25, 20, 31) {real, imag} */,
  {32'hc18685e2, 32'h413f578e} /* (25, 20, 30) {real, imag} */,
  {32'h4097e842, 32'hc09dd7a4} /* (25, 20, 29) {real, imag} */,
  {32'hc1477f41, 32'h40fa4344} /* (25, 20, 28) {real, imag} */,
  {32'h424619f2, 32'hc1f3df9d} /* (25, 20, 27) {real, imag} */,
  {32'h403d907f, 32'h4106ec94} /* (25, 20, 26) {real, imag} */,
  {32'hc1f558c6, 32'h4176552a} /* (25, 20, 25) {real, imag} */,
  {32'h408e0880, 32'h4253d7d0} /* (25, 20, 24) {real, imag} */,
  {32'h422341af, 32'hc1ca6a0e} /* (25, 20, 23) {real, imag} */,
  {32'hc18737f2, 32'hc1247dba} /* (25, 20, 22) {real, imag} */,
  {32'hbf2c3e30, 32'hc0fe3314} /* (25, 20, 21) {real, imag} */,
  {32'hc0ad03e7, 32'hc15363c6} /* (25, 20, 20) {real, imag} */,
  {32'h40c4423a, 32'h40ec548c} /* (25, 20, 19) {real, imag} */,
  {32'hc13a5c22, 32'h410b8b6a} /* (25, 20, 18) {real, imag} */,
  {32'h4038baa7, 32'h411554b3} /* (25, 20, 17) {real, imag} */,
  {32'hc088c7c9, 32'h40b29969} /* (25, 20, 16) {real, imag} */,
  {32'hc11f7176, 32'h41724445} /* (25, 20, 15) {real, imag} */,
  {32'h40b8b38f, 32'h41504a16} /* (25, 20, 14) {real, imag} */,
  {32'h41b3a38a, 32'h413a431e} /* (25, 20, 13) {real, imag} */,
  {32'h4023482c, 32'h40c1880c} /* (25, 20, 12) {real, imag} */,
  {32'h41bb9888, 32'hc22928ac} /* (25, 20, 11) {real, imag} */,
  {32'h412208a8, 32'hc0d65558} /* (25, 20, 10) {real, imag} */,
  {32'h41c31cfa, 32'hbf096b40} /* (25, 20, 9) {real, imag} */,
  {32'hc1bf43fa, 32'hc1a3e45f} /* (25, 20, 8) {real, imag} */,
  {32'hc16921ab, 32'h41aeab3b} /* (25, 20, 7) {real, imag} */,
  {32'hc02be621, 32'h429011e6} /* (25, 20, 6) {real, imag} */,
  {32'hc1a679fc, 32'hc1a6285d} /* (25, 20, 5) {real, imag} */,
  {32'hbfa2dde8, 32'h4272c9d6} /* (25, 20, 4) {real, imag} */,
  {32'hc1350c9f, 32'hc2338304} /* (25, 20, 3) {real, imag} */,
  {32'hc12b2f51, 32'h41a7233b} /* (25, 20, 2) {real, imag} */,
  {32'h406347d1, 32'h420a4c24} /* (25, 20, 1) {real, imag} */,
  {32'hc08d5fa9, 32'h4182a865} /* (25, 20, 0) {real, imag} */,
  {32'h42519686, 32'h4132c424} /* (25, 19, 31) {real, imag} */,
  {32'h41a223df, 32'hc11bd6d4} /* (25, 19, 30) {real, imag} */,
  {32'h3f2571c0, 32'h40b210a8} /* (25, 19, 29) {real, imag} */,
  {32'hc0f9cf4e, 32'hc1ac378a} /* (25, 19, 28) {real, imag} */,
  {32'h4191bd6d, 32'h3f743810} /* (25, 19, 27) {real, imag} */,
  {32'hc1654d40, 32'h42898520} /* (25, 19, 26) {real, imag} */,
  {32'hc1da2e8d, 32'hc19a3778} /* (25, 19, 25) {real, imag} */,
  {32'hc112860a, 32'h3f94e868} /* (25, 19, 24) {real, imag} */,
  {32'h40a60f57, 32'hc1d48ac8} /* (25, 19, 23) {real, imag} */,
  {32'h412961e4, 32'hc130c468} /* (25, 19, 22) {real, imag} */,
  {32'h418b5156, 32'hc084f2a6} /* (25, 19, 21) {real, imag} */,
  {32'h40a5b1f4, 32'hc0c90ef1} /* (25, 19, 20) {real, imag} */,
  {32'h410f7879, 32'h4133a649} /* (25, 19, 19) {real, imag} */,
  {32'hc11a9baf, 32'h41840ce2} /* (25, 19, 18) {real, imag} */,
  {32'h3f175e30, 32'hc1990c9d} /* (25, 19, 17) {real, imag} */,
  {32'h416f8d12, 32'hc04e5450} /* (25, 19, 16) {real, imag} */,
  {32'hc08e18ae, 32'hbf1f35e0} /* (25, 19, 15) {real, imag} */,
  {32'hbfd237c8, 32'hc18ec0e0} /* (25, 19, 14) {real, imag} */,
  {32'hbf968858, 32'h412be53f} /* (25, 19, 13) {real, imag} */,
  {32'hc0f56f70, 32'hc1aa9e37} /* (25, 19, 12) {real, imag} */,
  {32'h400eb9ce, 32'h4198cc38} /* (25, 19, 11) {real, imag} */,
  {32'h40b32e5c, 32'hc15f6ea4} /* (25, 19, 10) {real, imag} */,
  {32'h3ebbd510, 32'hc121c649} /* (25, 19, 9) {real, imag} */,
  {32'h41f14d17, 32'h3f8d61e8} /* (25, 19, 8) {real, imag} */,
  {32'hc0df32f4, 32'hc033a518} /* (25, 19, 7) {real, imag} */,
  {32'hc1a5f45c, 32'h41696172} /* (25, 19, 6) {real, imag} */,
  {32'h4212bdee, 32'hc0dddebe} /* (25, 19, 5) {real, imag} */,
  {32'hc1f28e8c, 32'h41902c30} /* (25, 19, 4) {real, imag} */,
  {32'hc239f36f, 32'h422490c1} /* (25, 19, 3) {real, imag} */,
  {32'h419b3421, 32'hc1597868} /* (25, 19, 2) {real, imag} */,
  {32'hc058fa28, 32'hc0f45ea1} /* (25, 19, 1) {real, imag} */,
  {32'hc1f70753, 32'h422c9a11} /* (25, 19, 0) {real, imag} */,
  {32'hc22e08ed, 32'hc180c167} /* (25, 18, 31) {real, imag} */,
  {32'hc132fd1e, 32'hc1ffebd2} /* (25, 18, 30) {real, imag} */,
  {32'h417bb0b4, 32'hc04320c8} /* (25, 18, 29) {real, imag} */,
  {32'hc08d8e1d, 32'hc1674fb2} /* (25, 18, 28) {real, imag} */,
  {32'h403fcb94, 32'hc09d404c} /* (25, 18, 27) {real, imag} */,
  {32'h42385d2a, 32'h419c2af6} /* (25, 18, 26) {real, imag} */,
  {32'h4208560c, 32'h410016d6} /* (25, 18, 25) {real, imag} */,
  {32'hc151ada6, 32'h408ab3ce} /* (25, 18, 24) {real, imag} */,
  {32'hc0c08bb3, 32'h413fb15d} /* (25, 18, 23) {real, imag} */,
  {32'h413a9d48, 32'h4146375a} /* (25, 18, 22) {real, imag} */,
  {32'h409561fd, 32'h40a8ddbe} /* (25, 18, 21) {real, imag} */,
  {32'h415595bc, 32'hc0ae2c18} /* (25, 18, 20) {real, imag} */,
  {32'hc0e1b57b, 32'hc0cc6c00} /* (25, 18, 19) {real, imag} */,
  {32'hc030ff27, 32'hc0896d3e} /* (25, 18, 18) {real, imag} */,
  {32'hbf836628, 32'h40d076fa} /* (25, 18, 17) {real, imag} */,
  {32'h404f32a8, 32'hbfc312be} /* (25, 18, 16) {real, imag} */,
  {32'h411c646d, 32'h3e1b2330} /* (25, 18, 15) {real, imag} */,
  {32'h4114781e, 32'hc071f0cc} /* (25, 18, 14) {real, imag} */,
  {32'h406a78de, 32'h4028b758} /* (25, 18, 13) {real, imag} */,
  {32'h4031a9e2, 32'h4103c4b3} /* (25, 18, 12) {real, imag} */,
  {32'hc0e748ef, 32'hc14c7fb7} /* (25, 18, 11) {real, imag} */,
  {32'hc024dd30, 32'h414cc514} /* (25, 18, 10) {real, imag} */,
  {32'hc074d97a, 32'hc0a73736} /* (25, 18, 9) {real, imag} */,
  {32'hc08f6c55, 32'hc189893a} /* (25, 18, 8) {real, imag} */,
  {32'h41a18061, 32'h41a78726} /* (25, 18, 7) {real, imag} */,
  {32'hc2203bb6, 32'hc18f6946} /* (25, 18, 6) {real, imag} */,
  {32'h41ebe758, 32'h42690348} /* (25, 18, 5) {real, imag} */,
  {32'hc123bc98, 32'h41e66a87} /* (25, 18, 4) {real, imag} */,
  {32'h41d8efae, 32'hc19096ec} /* (25, 18, 3) {real, imag} */,
  {32'h40e75274, 32'hc17f58d4} /* (25, 18, 2) {real, imag} */,
  {32'hc0a15f08, 32'h40291268} /* (25, 18, 1) {real, imag} */,
  {32'hc18343da, 32'hbfae7c96} /* (25, 18, 0) {real, imag} */,
  {32'h4097b2e2, 32'h424448a0} /* (25, 17, 31) {real, imag} */,
  {32'h41225b68, 32'h41aae998} /* (25, 17, 30) {real, imag} */,
  {32'h41531d94, 32'h40c61a7f} /* (25, 17, 29) {real, imag} */,
  {32'h40ffb521, 32'h420a7c80} /* (25, 17, 28) {real, imag} */,
  {32'h407edaab, 32'hc1eb28f2} /* (25, 17, 27) {real, imag} */,
  {32'hbfa17af2, 32'hc1195baa} /* (25, 17, 26) {real, imag} */,
  {32'h41cf5895, 32'hc1d433f7} /* (25, 17, 25) {real, imag} */,
  {32'hbf16d348, 32'h41b7b59a} /* (25, 17, 24) {real, imag} */,
  {32'h41470582, 32'hc1941c50} /* (25, 17, 23) {real, imag} */,
  {32'hc19ba644, 32'h40c1f99d} /* (25, 17, 22) {real, imag} */,
  {32'hc0066470, 32'hc117aec8} /* (25, 17, 21) {real, imag} */,
  {32'hc0c21327, 32'h4059148d} /* (25, 17, 20) {real, imag} */,
  {32'h3fb5a56a, 32'hc0c4de1e} /* (25, 17, 19) {real, imag} */,
  {32'hc1066d24, 32'h3d0d35c0} /* (25, 17, 18) {real, imag} */,
  {32'h40087c21, 32'h4016b3b0} /* (25, 17, 17) {real, imag} */,
  {32'hbeccff00, 32'hbfc665cc} /* (25, 17, 16) {real, imag} */,
  {32'h40a87fe4, 32'h3fd77380} /* (25, 17, 15) {real, imag} */,
  {32'h40e83486, 32'hc03c7d07} /* (25, 17, 14) {real, imag} */,
  {32'h40614ad5, 32'hbea097b8} /* (25, 17, 13) {real, imag} */,
  {32'hc07498de, 32'hc061fe1b} /* (25, 17, 12) {real, imag} */,
  {32'h417e1bcc, 32'h41029608} /* (25, 17, 11) {real, imag} */,
  {32'h40061aec, 32'hc1961dd2} /* (25, 17, 10) {real, imag} */,
  {32'h4124468a, 32'h413b7f93} /* (25, 17, 9) {real, imag} */,
  {32'hc14e0228, 32'hc1729f5d} /* (25, 17, 8) {real, imag} */,
  {32'h4229e9ea, 32'hc0f4fca4} /* (25, 17, 7) {real, imag} */,
  {32'hbf21dc74, 32'h41a70ee8} /* (25, 17, 6) {real, imag} */,
  {32'h3d5688c0, 32'hc1be419a} /* (25, 17, 5) {real, imag} */,
  {32'hc0449e66, 32'hc1f8d28b} /* (25, 17, 4) {real, imag} */,
  {32'hc090f35c, 32'hc10ddba0} /* (25, 17, 3) {real, imag} */,
  {32'hc1c9ded2, 32'h413d252c} /* (25, 17, 2) {real, imag} */,
  {32'h41915150, 32'h417fdabe} /* (25, 17, 1) {real, imag} */,
  {32'hc242537e, 32'h41506eac} /* (25, 17, 0) {real, imag} */,
  {32'hc21d34ec, 32'h41af7c39} /* (25, 16, 31) {real, imag} */,
  {32'hc200bf14, 32'h3f9f3090} /* (25, 16, 30) {real, imag} */,
  {32'h40990980, 32'h411c1b51} /* (25, 16, 29) {real, imag} */,
  {32'hc03d91e0, 32'hc151143e} /* (25, 16, 28) {real, imag} */,
  {32'h412776c3, 32'hc158a8a7} /* (25, 16, 27) {real, imag} */,
  {32'h40cdb740, 32'hc1056348} /* (25, 16, 26) {real, imag} */,
  {32'hc1f0ae1f, 32'hbdbca480} /* (25, 16, 25) {real, imag} */,
  {32'h400e2e1c, 32'hc18bdcbf} /* (25, 16, 24) {real, imag} */,
  {32'h3fce3244, 32'hc1b60bca} /* (25, 16, 23) {real, imag} */,
  {32'hc10c9cfb, 32'h419e4024} /* (25, 16, 22) {real, imag} */,
  {32'hc0974d89, 32'hc17db782} /* (25, 16, 21) {real, imag} */,
  {32'h3fd67760, 32'hbfb69a2c} /* (25, 16, 20) {real, imag} */,
  {32'h3ec79a50, 32'h41082e0f} /* (25, 16, 19) {real, imag} */,
  {32'hc01ffe86, 32'h408abb2a} /* (25, 16, 18) {real, imag} */,
  {32'h4021af00, 32'h3f5a0760} /* (25, 16, 17) {real, imag} */,
  {32'hbfc845e4, 32'h4081be89} /* (25, 16, 16) {real, imag} */,
  {32'hc1033058, 32'hbfc63230} /* (25, 16, 15) {real, imag} */,
  {32'hc0b22a11, 32'h40d0947c} /* (25, 16, 14) {real, imag} */,
  {32'h40d1ecb1, 32'h414200c5} /* (25, 16, 13) {real, imag} */,
  {32'hc119c612, 32'h40cf9697} /* (25, 16, 12) {real, imag} */,
  {32'h40d8de7d, 32'hc1031862} /* (25, 16, 11) {real, imag} */,
  {32'h40ad1108, 32'hc055b618} /* (25, 16, 10) {real, imag} */,
  {32'hc0412746, 32'h40be53b2} /* (25, 16, 9) {real, imag} */,
  {32'h41652113, 32'hc020a5da} /* (25, 16, 8) {real, imag} */,
  {32'h4106ceca, 32'h412d097d} /* (25, 16, 7) {real, imag} */,
  {32'hc1db20f8, 32'h418308b9} /* (25, 16, 6) {real, imag} */,
  {32'hc123cb31, 32'h3f1ef800} /* (25, 16, 5) {real, imag} */,
  {32'h4230059c, 32'hbedaa3f0} /* (25, 16, 4) {real, imag} */,
  {32'h41e0bd04, 32'h4196f108} /* (25, 16, 3) {real, imag} */,
  {32'hc1d802f9, 32'h41c4a0c9} /* (25, 16, 2) {real, imag} */,
  {32'h41c0646b, 32'hc197ea6d} /* (25, 16, 1) {real, imag} */,
  {32'h40eb4281, 32'hbf1f9838} /* (25, 16, 0) {real, imag} */,
  {32'hbbe05800, 32'hc190e75f} /* (25, 15, 31) {real, imag} */,
  {32'h41374eaa, 32'h42300c54} /* (25, 15, 30) {real, imag} */,
  {32'h414ed295, 32'h411240aa} /* (25, 15, 29) {real, imag} */,
  {32'hc159ef72, 32'h40a165dc} /* (25, 15, 28) {real, imag} */,
  {32'hc15b83e6, 32'hbff4229c} /* (25, 15, 27) {real, imag} */,
  {32'hc2041c38, 32'hc1d95f1d} /* (25, 15, 26) {real, imag} */,
  {32'hc08521a4, 32'h40dcee66} /* (25, 15, 25) {real, imag} */,
  {32'hc0909acf, 32'hc1241016} /* (25, 15, 24) {real, imag} */,
  {32'hc0d204d6, 32'hc1a1095c} /* (25, 15, 23) {real, imag} */,
  {32'h3facade4, 32'hc092fc3b} /* (25, 15, 22) {real, imag} */,
  {32'h3fdbc7d0, 32'h410f9574} /* (25, 15, 21) {real, imag} */,
  {32'hc0a18cce, 32'h40447582} /* (25, 15, 20) {real, imag} */,
  {32'h418b1ba8, 32'h411c67d6} /* (25, 15, 19) {real, imag} */,
  {32'h40ac3c6a, 32'hc156353e} /* (25, 15, 18) {real, imag} */,
  {32'h40d6d114, 32'hc115b193} /* (25, 15, 17) {real, imag} */,
  {32'h40df8410, 32'h4002c896} /* (25, 15, 16) {real, imag} */,
  {32'hc02da927, 32'hc084df4a} /* (25, 15, 15) {real, imag} */,
  {32'h40d5e168, 32'hbe949dc0} /* (25, 15, 14) {real, imag} */,
  {32'hc0ef5cb4, 32'hc11d6c8c} /* (25, 15, 13) {real, imag} */,
  {32'h4085c93e, 32'hc04d0cc2} /* (25, 15, 12) {real, imag} */,
  {32'hc1babd79, 32'h3df79dc0} /* (25, 15, 11) {real, imag} */,
  {32'hc0d832c7, 32'h4117d63e} /* (25, 15, 10) {real, imag} */,
  {32'hc0910012, 32'h409c610a} /* (25, 15, 9) {real, imag} */,
  {32'h412cec1e, 32'h41be9519} /* (25, 15, 8) {real, imag} */,
  {32'h407a2283, 32'h418f0d40} /* (25, 15, 7) {real, imag} */,
  {32'h41d63e51, 32'hc1b6a2bf} /* (25, 15, 6) {real, imag} */,
  {32'h408bfabd, 32'hbff5de14} /* (25, 15, 5) {real, imag} */,
  {32'h40a6571c, 32'hc13fc3ea} /* (25, 15, 4) {real, imag} */,
  {32'hc149b631, 32'hc0c9ff78} /* (25, 15, 3) {real, imag} */,
  {32'h404d5714, 32'h4043d5d0} /* (25, 15, 2) {real, imag} */,
  {32'h410b9d8d, 32'h4167df12} /* (25, 15, 1) {real, imag} */,
  {32'hc257425c, 32'hc16b1de2} /* (25, 15, 0) {real, imag} */,
  {32'hc18209a1, 32'hc108090b} /* (25, 14, 31) {real, imag} */,
  {32'h4102e660, 32'hc1bb8cc6} /* (25, 14, 30) {real, imag} */,
  {32'hc22bc885, 32'h40ab8bb2} /* (25, 14, 29) {real, imag} */,
  {32'hc1fb1faa, 32'h41a8577a} /* (25, 14, 28) {real, imag} */,
  {32'hc025a000, 32'hc05dddc0} /* (25, 14, 27) {real, imag} */,
  {32'hc1652818, 32'h41b1cde7} /* (25, 14, 26) {real, imag} */,
  {32'h40295806, 32'hc22278bc} /* (25, 14, 25) {real, imag} */,
  {32'h4195979c, 32'hc1b77cc4} /* (25, 14, 24) {real, imag} */,
  {32'h41b7fda4, 32'h40a65fb2} /* (25, 14, 23) {real, imag} */,
  {32'h412a14a3, 32'hc11b51be} /* (25, 14, 22) {real, imag} */,
  {32'h413b3802, 32'h40554970} /* (25, 14, 21) {real, imag} */,
  {32'h4126917d, 32'hc0d7f5bb} /* (25, 14, 20) {real, imag} */,
  {32'h4127e961, 32'h40113914} /* (25, 14, 19) {real, imag} */,
  {32'h4197a04f, 32'hc01e2b37} /* (25, 14, 18) {real, imag} */,
  {32'hc11c4bc4, 32'h400a1302} /* (25, 14, 17) {real, imag} */,
  {32'hc0ac5870, 32'hc096e536} /* (25, 14, 16) {real, imag} */,
  {32'hbfb434dc, 32'hc0be55f3} /* (25, 14, 15) {real, imag} */,
  {32'h3f528d40, 32'hbfa7533e} /* (25, 14, 14) {real, imag} */,
  {32'h40f81326, 32'h40d7296e} /* (25, 14, 13) {real, imag} */,
  {32'h3fe42df8, 32'h4047d40e} /* (25, 14, 12) {real, imag} */,
  {32'h40c2c2f8, 32'hc0bd9220} /* (25, 14, 11) {real, imag} */,
  {32'hbe9415a0, 32'h42062254} /* (25, 14, 10) {real, imag} */,
  {32'hc10f17d4, 32'hc121df35} /* (25, 14, 9) {real, imag} */,
  {32'hc05d6616, 32'hc1d576b0} /* (25, 14, 8) {real, imag} */,
  {32'h40c4a63d, 32'h3df38d00} /* (25, 14, 7) {real, imag} */,
  {32'hc1ffdc58, 32'h4018a818} /* (25, 14, 6) {real, imag} */,
  {32'hc23faaf0, 32'hc25a1ba8} /* (25, 14, 5) {real, imag} */,
  {32'h41a947b6, 32'hc19c2932} /* (25, 14, 4) {real, imag} */,
  {32'h41598294, 32'hc1c68324} /* (25, 14, 3) {real, imag} */,
  {32'hc22ae0da, 32'h40f35afc} /* (25, 14, 2) {real, imag} */,
  {32'hc1af1ec9, 32'hc1c0255a} /* (25, 14, 1) {real, imag} */,
  {32'h4202ef90, 32'hc1510d35} /* (25, 14, 0) {real, imag} */,
  {32'h41bcdb89, 32'h407735d0} /* (25, 13, 31) {real, imag} */,
  {32'h418841e6, 32'h425ec246} /* (25, 13, 30) {real, imag} */,
  {32'hc19edd5b, 32'hc1f3db93} /* (25, 13, 29) {real, imag} */,
  {32'hc05f7d84, 32'hc11b5e6e} /* (25, 13, 28) {real, imag} */,
  {32'hc1933174, 32'h41061dc2} /* (25, 13, 27) {real, imag} */,
  {32'h41050300, 32'hc204e286} /* (25, 13, 26) {real, imag} */,
  {32'h40cf8030, 32'hc0d65270} /* (25, 13, 25) {real, imag} */,
  {32'hc1303685, 32'h40e322b8} /* (25, 13, 24) {real, imag} */,
  {32'h402fd160, 32'h409417f0} /* (25, 13, 23) {real, imag} */,
  {32'h40aa2224, 32'hc0b500dc} /* (25, 13, 22) {real, imag} */,
  {32'h416520de, 32'hc17e570c} /* (25, 13, 21) {real, imag} */,
  {32'h42235bdc, 32'hbf812cec} /* (25, 13, 20) {real, imag} */,
  {32'hc014c6c1, 32'hc13b1b70} /* (25, 13, 19) {real, imag} */,
  {32'h3f6c77d0, 32'hbf8fc6a0} /* (25, 13, 18) {real, imag} */,
  {32'hbf2f4a20, 32'h41348e84} /* (25, 13, 17) {real, imag} */,
  {32'h408acda9, 32'h41418a22} /* (25, 13, 16) {real, imag} */,
  {32'hc0f5daaa, 32'hc0f87738} /* (25, 13, 15) {real, imag} */,
  {32'hc10b8159, 32'hbf2b8a80} /* (25, 13, 14) {real, imag} */,
  {32'hc0281d6f, 32'hbfa205e0} /* (25, 13, 13) {real, imag} */,
  {32'hc02ad348, 32'h412bbe82} /* (25, 13, 12) {real, imag} */,
  {32'hc0f638f9, 32'h40867e48} /* (25, 13, 11) {real, imag} */,
  {32'h41b9ca15, 32'hc17ec4a2} /* (25, 13, 10) {real, imag} */,
  {32'h41740484, 32'hc146f3b4} /* (25, 13, 9) {real, imag} */,
  {32'hbfb6c768, 32'h40747f04} /* (25, 13, 8) {real, imag} */,
  {32'hc205acbb, 32'hc28d99c3} /* (25, 13, 7) {real, imag} */,
  {32'hc1308444, 32'h4123ae5a} /* (25, 13, 6) {real, imag} */,
  {32'hc108efcd, 32'h4119acbe} /* (25, 13, 5) {real, imag} */,
  {32'hc129950f, 32'hc1f39df1} /* (25, 13, 4) {real, imag} */,
  {32'hc196a22b, 32'hc1eaf3fb} /* (25, 13, 3) {real, imag} */,
  {32'h429642f4, 32'h41962253} /* (25, 13, 2) {real, imag} */,
  {32'h41414b46, 32'h420c11d3} /* (25, 13, 1) {real, imag} */,
  {32'h40d46383, 32'h41022a6a} /* (25, 13, 0) {real, imag} */,
  {32'hc1679247, 32'h420c3ba4} /* (25, 12, 31) {real, imag} */,
  {32'h424bf022, 32'hc169eaf1} /* (25, 12, 30) {real, imag} */,
  {32'hc1b75b20, 32'h407a0924} /* (25, 12, 29) {real, imag} */,
  {32'h407a50c1, 32'h423ecd2c} /* (25, 12, 28) {real, imag} */,
  {32'h40c499a8, 32'h41354124} /* (25, 12, 27) {real, imag} */,
  {32'hc23aff74, 32'h4064533c} /* (25, 12, 26) {real, imag} */,
  {32'h41988034, 32'hc233ee16} /* (25, 12, 25) {real, imag} */,
  {32'hc2033bdf, 32'h41028fa6} /* (25, 12, 24) {real, imag} */,
  {32'hc20947c0, 32'hc1e21120} /* (25, 12, 23) {real, imag} */,
  {32'hc0595f16, 32'hc159b743} /* (25, 12, 22) {real, imag} */,
  {32'hc187e802, 32'hc142cdcc} /* (25, 12, 21) {real, imag} */,
  {32'hc13ffbba, 32'h421457f8} /* (25, 12, 20) {real, imag} */,
  {32'hc12c8284, 32'h410fb72c} /* (25, 12, 19) {real, imag} */,
  {32'hc045881c, 32'hc0bac1fe} /* (25, 12, 18) {real, imag} */,
  {32'hbfbb182a, 32'h40c8690c} /* (25, 12, 17) {real, imag} */,
  {32'h41084df8, 32'hbf972d18} /* (25, 12, 16) {real, imag} */,
  {32'hc10d8517, 32'h4123b082} /* (25, 12, 15) {real, imag} */,
  {32'hc003cafc, 32'hc1947e8e} /* (25, 12, 14) {real, imag} */,
  {32'h4063e8b2, 32'h3fb37864} /* (25, 12, 13) {real, imag} */,
  {32'hc1e75bf7, 32'hc16993a8} /* (25, 12, 12) {real, imag} */,
  {32'h4135c048, 32'hbef3fb80} /* (25, 12, 11) {real, imag} */,
  {32'h4146250c, 32'hc211e0ae} /* (25, 12, 10) {real, imag} */,
  {32'h40355ddc, 32'h40411b44} /* (25, 12, 9) {real, imag} */,
  {32'h4121c44d, 32'hc256f7e6} /* (25, 12, 8) {real, imag} */,
  {32'hc0b6f48a, 32'h41521a50} /* (25, 12, 7) {real, imag} */,
  {32'hc1b82773, 32'hc197b022} /* (25, 12, 6) {real, imag} */,
  {32'h41c898ac, 32'hc036c530} /* (25, 12, 5) {real, imag} */,
  {32'h40223b87, 32'h422c1cca} /* (25, 12, 4) {real, imag} */,
  {32'h41db934c, 32'hc1a5bafc} /* (25, 12, 3) {real, imag} */,
  {32'hc0e53b70, 32'hc16012ef} /* (25, 12, 2) {real, imag} */,
  {32'h3fb45098, 32'h40bf9ee0} /* (25, 12, 1) {real, imag} */,
  {32'h41bd79a6, 32'hc1c422de} /* (25, 12, 0) {real, imag} */,
  {32'hc191ecc0, 32'h4152ac54} /* (25, 11, 31) {real, imag} */,
  {32'h41d11d1c, 32'h4116652e} /* (25, 11, 30) {real, imag} */,
  {32'hc24db34c, 32'h405e71b0} /* (25, 11, 29) {real, imag} */,
  {32'h421e94a9, 32'hc0f163f8} /* (25, 11, 28) {real, imag} */,
  {32'hc0784ce0, 32'h41dcdf56} /* (25, 11, 27) {real, imag} */,
  {32'h4211bbfb, 32'h41c02740} /* (25, 11, 26) {real, imag} */,
  {32'h422ef9db, 32'hc09cd8ac} /* (25, 11, 25) {real, imag} */,
  {32'hc1d24664, 32'h413e5e10} /* (25, 11, 24) {real, imag} */,
  {32'h422df75c, 32'hc0970444} /* (25, 11, 23) {real, imag} */,
  {32'h40b2c3a8, 32'h418ead9e} /* (25, 11, 22) {real, imag} */,
  {32'hc1a4f2b5, 32'h4116265c} /* (25, 11, 21) {real, imag} */,
  {32'hc1a05a5c, 32'hc18387d3} /* (25, 11, 20) {real, imag} */,
  {32'hc1211072, 32'h40af68fa} /* (25, 11, 19) {real, imag} */,
  {32'hc18bc499, 32'h41a9aeb6} /* (25, 11, 18) {real, imag} */,
  {32'hc025ff78, 32'hc1b7fd0e} /* (25, 11, 17) {real, imag} */,
  {32'hc0cbf4ad, 32'h4148b5a6} /* (25, 11, 16) {real, imag} */,
  {32'hc16c958a, 32'h40549410} /* (25, 11, 15) {real, imag} */,
  {32'h413043d8, 32'hc073704c} /* (25, 11, 14) {real, imag} */,
  {32'h41731dea, 32'h410c2253} /* (25, 11, 13) {real, imag} */,
  {32'hc1269b35, 32'h41a355f7} /* (25, 11, 12) {real, imag} */,
  {32'h4203e164, 32'hc0af216d} /* (25, 11, 11) {real, imag} */,
  {32'h40606448, 32'hc1c693c6} /* (25, 11, 10) {real, imag} */,
  {32'h4186fa85, 32'h42422324} /* (25, 11, 9) {real, imag} */,
  {32'hc2006ffa, 32'hc1888868} /* (25, 11, 8) {real, imag} */,
  {32'hc13c6b9f, 32'hc1f8d717} /* (25, 11, 7) {real, imag} */,
  {32'h41adffae, 32'h40c86820} /* (25, 11, 6) {real, imag} */,
  {32'hc28d2ca1, 32'h3fedaab8} /* (25, 11, 5) {real, imag} */,
  {32'h41810960, 32'hc22de64e} /* (25, 11, 4) {real, imag} */,
  {32'hc16d7a7e, 32'h421ab8a1} /* (25, 11, 3) {real, imag} */,
  {32'hc1e02568, 32'h3f7cea08} /* (25, 11, 2) {real, imag} */,
  {32'h427bf42c, 32'h42615415} /* (25, 11, 1) {real, imag} */,
  {32'hc07693e6, 32'h4123c16e} /* (25, 11, 0) {real, imag} */,
  {32'h401143f8, 32'hc183fc17} /* (25, 10, 31) {real, imag} */,
  {32'h40503338, 32'hc2f6855a} /* (25, 10, 30) {real, imag} */,
  {32'hc1498eb4, 32'hc1de6402} /* (25, 10, 29) {real, imag} */,
  {32'h41d462ac, 32'hc28fa563} /* (25, 10, 28) {real, imag} */,
  {32'hc02e6930, 32'h4199e17a} /* (25, 10, 27) {real, imag} */,
  {32'h421f7257, 32'h41ee52a3} /* (25, 10, 26) {real, imag} */,
  {32'h3ec05b20, 32'h426f7462} /* (25, 10, 25) {real, imag} */,
  {32'h3ffe81b8, 32'h41660e61} /* (25, 10, 24) {real, imag} */,
  {32'h42426510, 32'h42667f5d} /* (25, 10, 23) {real, imag} */,
  {32'hc243d6f2, 32'hc19594f8} /* (25, 10, 22) {real, imag} */,
  {32'hc0ac810a, 32'h402d7188} /* (25, 10, 21) {real, imag} */,
  {32'h4183a155, 32'hbe3d6940} /* (25, 10, 20) {real, imag} */,
  {32'hc0e810d8, 32'hc1a48c80} /* (25, 10, 19) {real, imag} */,
  {32'hc186a09e, 32'hc07b62a4} /* (25, 10, 18) {real, imag} */,
  {32'h4094a736, 32'hc1027d02} /* (25, 10, 17) {real, imag} */,
  {32'h4123e542, 32'hc1b6a0f2} /* (25, 10, 16) {real, imag} */,
  {32'hc101b3c9, 32'hc08fb663} /* (25, 10, 15) {real, imag} */,
  {32'h405b7ee4, 32'hc13075b9} /* (25, 10, 14) {real, imag} */,
  {32'hc18872ea, 32'h41d273e4} /* (25, 10, 13) {real, imag} */,
  {32'h415190d0, 32'hc1df94ac} /* (25, 10, 12) {real, imag} */,
  {32'h412e3329, 32'h41ded282} /* (25, 10, 11) {real, imag} */,
  {32'hc17104f6, 32'hc1240c76} /* (25, 10, 10) {real, imag} */,
  {32'hc13232c6, 32'hc236c8e3} /* (25, 10, 9) {real, imag} */,
  {32'h4030f55c, 32'h4205d1bd} /* (25, 10, 8) {real, imag} */,
  {32'hbfd4ca58, 32'h409cf54c} /* (25, 10, 7) {real, imag} */,
  {32'hc24a98cd, 32'h42237f2e} /* (25, 10, 6) {real, imag} */,
  {32'hc22fb103, 32'hc18806e2} /* (25, 10, 5) {real, imag} */,
  {32'h4265006e, 32'hc231950f} /* (25, 10, 4) {real, imag} */,
  {32'hc2855a22, 32'hc27597e1} /* (25, 10, 3) {real, imag} */,
  {32'h4216fea4, 32'h42acad50} /* (25, 10, 2) {real, imag} */,
  {32'h421f3f3e, 32'h426ed494} /* (25, 10, 1) {real, imag} */,
  {32'h40d33650, 32'h41f09cea} /* (25, 10, 0) {real, imag} */,
  {32'h427d2728, 32'hc2978a5a} /* (25, 9, 31) {real, imag} */,
  {32'h420f2ce9, 32'hc16e6737} /* (25, 9, 30) {real, imag} */,
  {32'hc1186be6, 32'h401b5740} /* (25, 9, 29) {real, imag} */,
  {32'hc199a36b, 32'h40089cf0} /* (25, 9, 28) {real, imag} */,
  {32'h41ead40b, 32'hc1413283} /* (25, 9, 27) {real, imag} */,
  {32'hc0eb92f2, 32'hc19ed8e7} /* (25, 9, 26) {real, imag} */,
  {32'hc0b0552e, 32'h4294778c} /* (25, 9, 25) {real, imag} */,
  {32'h421de295, 32'hc00d2f6c} /* (25, 9, 24) {real, imag} */,
  {32'h40fba7f8, 32'hc0a3e70a} /* (25, 9, 23) {real, imag} */,
  {32'hc12559a0, 32'hc184d80a} /* (25, 9, 22) {real, imag} */,
  {32'h4102469a, 32'hc178a527} /* (25, 9, 21) {real, imag} */,
  {32'hc0abbfec, 32'hc0601960} /* (25, 9, 20) {real, imag} */,
  {32'hc2349329, 32'hbf5ef600} /* (25, 9, 19) {real, imag} */,
  {32'hc11fb214, 32'h4118058f} /* (25, 9, 18) {real, imag} */,
  {32'h3fa17294, 32'h403c59c8} /* (25, 9, 17) {real, imag} */,
  {32'h410b89ff, 32'h3fef0d10} /* (25, 9, 16) {real, imag} */,
  {32'h411cbc1e, 32'hc1b00191} /* (25, 9, 15) {real, imag} */,
  {32'h406ca8b0, 32'hc1d61990} /* (25, 9, 14) {real, imag} */,
  {32'h41f8dfda, 32'h410d7c3c} /* (25, 9, 13) {real, imag} */,
  {32'hc18a0fc3, 32'h40def6e4} /* (25, 9, 12) {real, imag} */,
  {32'hc05427f8, 32'hc163bbdd} /* (25, 9, 11) {real, imag} */,
  {32'h427b5c34, 32'h419d5bb4} /* (25, 9, 10) {real, imag} */,
  {32'hc285a116, 32'hc20efad0} /* (25, 9, 9) {real, imag} */,
  {32'h41afd0a8, 32'h41a22fe2} /* (25, 9, 8) {real, imag} */,
  {32'h40077794, 32'h41c4ee5e} /* (25, 9, 7) {real, imag} */,
  {32'hc200d712, 32'h428f58a0} /* (25, 9, 6) {real, imag} */,
  {32'hc26aa0b8, 32'hc1f4b758} /* (25, 9, 5) {real, imag} */,
  {32'h428b9538, 32'hc239c86d} /* (25, 9, 4) {real, imag} */,
  {32'h3fb2e890, 32'h42cf3024} /* (25, 9, 3) {real, imag} */,
  {32'h42a02f5c, 32'h4229ce20} /* (25, 9, 2) {real, imag} */,
  {32'hc265ace8, 32'hc28fe8c4} /* (25, 9, 1) {real, imag} */,
  {32'hc176a613, 32'h418fc4f7} /* (25, 9, 0) {real, imag} */,
  {32'hc1eae67b, 32'hc237ca37} /* (25, 8, 31) {real, imag} */,
  {32'hc27fb875, 32'hc10b3ec2} /* (25, 8, 30) {real, imag} */,
  {32'h42947456, 32'h41e79b40} /* (25, 8, 29) {real, imag} */,
  {32'hc24593dd, 32'hc25c64e2} /* (25, 8, 28) {real, imag} */,
  {32'hc24a916b, 32'hc122c0a4} /* (25, 8, 27) {real, imag} */,
  {32'hc1c341e8, 32'hc232fcfe} /* (25, 8, 26) {real, imag} */,
  {32'h42b37c96, 32'h4241bb7d} /* (25, 8, 25) {real, imag} */,
  {32'hc1f6decc, 32'h41b4c59e} /* (25, 8, 24) {real, imag} */,
  {32'hc270cc7b, 32'h41927864} /* (25, 8, 23) {real, imag} */,
  {32'hc26dad7a, 32'h4283cc07} /* (25, 8, 22) {real, imag} */,
  {32'h4099eb20, 32'h41bd183c} /* (25, 8, 21) {real, imag} */,
  {32'hc1513b32, 32'hc2543b4a} /* (25, 8, 20) {real, imag} */,
  {32'h419e365b, 32'h418980e4} /* (25, 8, 19) {real, imag} */,
  {32'h3f3c3870, 32'hbee79ec0} /* (25, 8, 18) {real, imag} */,
  {32'h41395d76, 32'hc1c56554} /* (25, 8, 17) {real, imag} */,
  {32'h401dec7c, 32'hc0579d10} /* (25, 8, 16) {real, imag} */,
  {32'hc0e59f5c, 32'hc015dd50} /* (25, 8, 15) {real, imag} */,
  {32'hbf4ddeb0, 32'h421a2d9c} /* (25, 8, 14) {real, imag} */,
  {32'h410a1572, 32'hc0906702} /* (25, 8, 13) {real, imag} */,
  {32'h41041412, 32'hc202cb76} /* (25, 8, 12) {real, imag} */,
  {32'h3f796d00, 32'hc0d9e252} /* (25, 8, 11) {real, imag} */,
  {32'hc205980e, 32'hc1c12809} /* (25, 8, 10) {real, imag} */,
  {32'h40cae838, 32'h3f2ba2c0} /* (25, 8, 9) {real, imag} */,
  {32'hc1187ed8, 32'h41a2b7e6} /* (25, 8, 8) {real, imag} */,
  {32'h432a4379, 32'h40e4bb80} /* (25, 8, 7) {real, imag} */,
  {32'h4251bb2a, 32'h41f05af8} /* (25, 8, 6) {real, imag} */,
  {32'h42aa5a32, 32'hc28006c4} /* (25, 8, 5) {real, imag} */,
  {32'h425a8ee7, 32'h40ab6b4c} /* (25, 8, 4) {real, imag} */,
  {32'h41982cc1, 32'hc2959514} /* (25, 8, 3) {real, imag} */,
  {32'h3f856060, 32'hc2632b5c} /* (25, 8, 2) {real, imag} */,
  {32'hc296c00e, 32'h422d0075} /* (25, 8, 1) {real, imag} */,
  {32'h40ef6634, 32'h42d34e44} /* (25, 8, 0) {real, imag} */,
  {32'hc299cf30, 32'hc056cec8} /* (25, 7, 31) {real, imag} */,
  {32'hc236cce5, 32'hc243c267} /* (25, 7, 30) {real, imag} */,
  {32'hc1556069, 32'hc1ed471c} /* (25, 7, 29) {real, imag} */,
  {32'h429f1629, 32'hc2eb6efb} /* (25, 7, 28) {real, imag} */,
  {32'hc29e2c88, 32'h40645d50} /* (25, 7, 27) {real, imag} */,
  {32'h428fea0e, 32'hc29a135d} /* (25, 7, 26) {real, imag} */,
  {32'hc15c1146, 32'hc23cd596} /* (25, 7, 25) {real, imag} */,
  {32'hc1834ad8, 32'h41fd22d3} /* (25, 7, 24) {real, imag} */,
  {32'h415ae816, 32'hc1936bde} /* (25, 7, 23) {real, imag} */,
  {32'h423d4089, 32'hc24717d2} /* (25, 7, 22) {real, imag} */,
  {32'hc206b1a4, 32'h418276a0} /* (25, 7, 21) {real, imag} */,
  {32'h421bca2e, 32'hc21cd278} /* (25, 7, 20) {real, imag} */,
  {32'h416e76c5, 32'h42089d01} /* (25, 7, 19) {real, imag} */,
  {32'h40f26ba2, 32'hbee16480} /* (25, 7, 18) {real, imag} */,
  {32'h42005d48, 32'hc0c38ae8} /* (25, 7, 17) {real, imag} */,
  {32'h41edae04, 32'hc13cf1da} /* (25, 7, 16) {real, imag} */,
  {32'hc1035790, 32'hc1e032ca} /* (25, 7, 15) {real, imag} */,
  {32'h40b5ac6e, 32'h4207406f} /* (25, 7, 14) {real, imag} */,
  {32'hc2356a36, 32'h4193d2da} /* (25, 7, 13) {real, imag} */,
  {32'hc1ae0547, 32'h419156b5} /* (25, 7, 12) {real, imag} */,
  {32'h3f61a680, 32'hc027d27c} /* (25, 7, 11) {real, imag} */,
  {32'hc21af501, 32'h4132321c} /* (25, 7, 10) {real, imag} */,
  {32'h419109e6, 32'h421f407e} /* (25, 7, 9) {real, imag} */,
  {32'hc203a5b2, 32'hc21cd770} /* (25, 7, 8) {real, imag} */,
  {32'hc2306ade, 32'h409eae44} /* (25, 7, 7) {real, imag} */,
  {32'h42340359, 32'h41f5e4bb} /* (25, 7, 6) {real, imag} */,
  {32'h3f8f0a40, 32'hc261e623} /* (25, 7, 5) {real, imag} */,
  {32'hc2bf39c3, 32'h42a8b5ad} /* (25, 7, 4) {real, imag} */,
  {32'h4223c2f3, 32'hc20ad4c0} /* (25, 7, 3) {real, imag} */,
  {32'hc215e339, 32'hc1ee9bce} /* (25, 7, 2) {real, imag} */,
  {32'h42c43d52, 32'hc22bf0ae} /* (25, 7, 1) {real, imag} */,
  {32'h425a7054, 32'h41b9784f} /* (25, 7, 0) {real, imag} */,
  {32'hc19cbba0, 32'hc184ceee} /* (25, 6, 31) {real, imag} */,
  {32'h4046c018, 32'hc0d9cb12} /* (25, 6, 30) {real, imag} */,
  {32'hc280c5b4, 32'hc20db107} /* (25, 6, 29) {real, imag} */,
  {32'hc1e75c92, 32'h42e4088b} /* (25, 6, 28) {real, imag} */,
  {32'h42816bda, 32'h3f8f9c40} /* (25, 6, 27) {real, imag} */,
  {32'h41df320b, 32'hc226fde3} /* (25, 6, 26) {real, imag} */,
  {32'hc2b54a0d, 32'hc19cc3cc} /* (25, 6, 25) {real, imag} */,
  {32'h40aabe58, 32'hc20a5222} /* (25, 6, 24) {real, imag} */,
  {32'hc27f006a, 32'h3fcc7968} /* (25, 6, 23) {real, imag} */,
  {32'hbf25cfc0, 32'hc1ae1cfc} /* (25, 6, 22) {real, imag} */,
  {32'hc150162d, 32'hc20d12b2} /* (25, 6, 21) {real, imag} */,
  {32'hc1402b94, 32'h422fc7c6} /* (25, 6, 20) {real, imag} */,
  {32'h427330cf, 32'h41a4d12c} /* (25, 6, 19) {real, imag} */,
  {32'h41f51d8f, 32'hc1745dbe} /* (25, 6, 18) {real, imag} */,
  {32'hc0e0b3de, 32'hc0fbf010} /* (25, 6, 17) {real, imag} */,
  {32'hc1878b4f, 32'h41abac9c} /* (25, 6, 16) {real, imag} */,
  {32'h4076497c, 32'hc1238cf8} /* (25, 6, 15) {real, imag} */,
  {32'hc1b0d4eb, 32'hc201336e} /* (25, 6, 14) {real, imag} */,
  {32'hc1d7bd56, 32'h3f886178} /* (25, 6, 13) {real, imag} */,
  {32'h42660b4d, 32'h41aab17d} /* (25, 6, 12) {real, imag} */,
  {32'hc0a5739a, 32'h4266bede} /* (25, 6, 11) {real, imag} */,
  {32'hc25ca0fe, 32'h427232ce} /* (25, 6, 10) {real, imag} */,
  {32'h4082287c, 32'hc1f51a9a} /* (25, 6, 9) {real, imag} */,
  {32'hc1def2a6, 32'hbe3b5080} /* (25, 6, 8) {real, imag} */,
  {32'h4271fd86, 32'h4202f060} /* (25, 6, 7) {real, imag} */,
  {32'hc26fe55a, 32'h424d8461} /* (25, 6, 6) {real, imag} */,
  {32'hc2580094, 32'h428eba4f} /* (25, 6, 5) {real, imag} */,
  {32'hc2a9d5e6, 32'h411e60d8} /* (25, 6, 4) {real, imag} */,
  {32'h41dc204e, 32'hc2208c7f} /* (25, 6, 3) {real, imag} */,
  {32'hc0f49bfc, 32'h41c17162} /* (25, 6, 2) {real, imag} */,
  {32'hc2a1af88, 32'hc2bdc484} /* (25, 6, 1) {real, imag} */,
  {32'hbf4b3fa0, 32'hc14411b0} /* (25, 6, 0) {real, imag} */,
  {32'hc2cfc38b, 32'h42abfb7e} /* (25, 5, 31) {real, imag} */,
  {32'hc2da62d7, 32'h428327c2} /* (25, 5, 30) {real, imag} */,
  {32'hc126ab4c, 32'hc28e5514} /* (25, 5, 29) {real, imag} */,
  {32'hc291bc22, 32'hc3134a4b} /* (25, 5, 28) {real, imag} */,
  {32'hc2822d1e, 32'hc131db3e} /* (25, 5, 27) {real, imag} */,
  {32'h42dc0e4a, 32'h430d2646} /* (25, 5, 26) {real, imag} */,
  {32'h418142f8, 32'hc233bf5b} /* (25, 5, 25) {real, imag} */,
  {32'hc0846494, 32'hc28ed6a1} /* (25, 5, 24) {real, imag} */,
  {32'h427f6004, 32'h41a39232} /* (25, 5, 23) {real, imag} */,
  {32'hc268f056, 32'hc23d28d4} /* (25, 5, 22) {real, imag} */,
  {32'h42033086, 32'h41921d41} /* (25, 5, 21) {real, imag} */,
  {32'hc1d75934, 32'hc20e7bef} /* (25, 5, 20) {real, imag} */,
  {32'hc1c4a5ba, 32'h41768c32} /* (25, 5, 19) {real, imag} */,
  {32'h3f4a2680, 32'h4025178c} /* (25, 5, 18) {real, imag} */,
  {32'h410f59bc, 32'h4045de97} /* (25, 5, 17) {real, imag} */,
  {32'hc12b6be0, 32'h412c3294} /* (25, 5, 16) {real, imag} */,
  {32'hc048d2ae, 32'h3fedb66e} /* (25, 5, 15) {real, imag} */,
  {32'h423194da, 32'h40c49de6} /* (25, 5, 14) {real, imag} */,
  {32'h411a0fa4, 32'h414239da} /* (25, 5, 13) {real, imag} */,
  {32'hc1c9395e, 32'hc1a67e4e} /* (25, 5, 12) {real, imag} */,
  {32'hc202909e, 32'h41c0db73} /* (25, 5, 11) {real, imag} */,
  {32'h3e93c1c0, 32'h4134f4f0} /* (25, 5, 10) {real, imag} */,
  {32'h42061de4, 32'hc2f06502} /* (25, 5, 9) {real, imag} */,
  {32'hc220fb88, 32'hc0f09de0} /* (25, 5, 8) {real, imag} */,
  {32'h413dc588, 32'hc2398dfb} /* (25, 5, 7) {real, imag} */,
  {32'h40cdc388, 32'h41887530} /* (25, 5, 6) {real, imag} */,
  {32'h411238c0, 32'hc2762e4e} /* (25, 5, 5) {real, imag} */,
  {32'hc0f50088, 32'h431f07f5} /* (25, 5, 4) {real, imag} */,
  {32'h42151427, 32'h4290869c} /* (25, 5, 3) {real, imag} */,
  {32'h41cfab74, 32'hc24ec8b8} /* (25, 5, 2) {real, imag} */,
  {32'hc2a4955d, 32'hc2b88ce6} /* (25, 5, 1) {real, imag} */,
  {32'h42cfe4fb, 32'hc2d265b8} /* (25, 5, 0) {real, imag} */,
  {32'hc1ea1817, 32'h42095a17} /* (25, 4, 31) {real, imag} */,
  {32'h3ea56780, 32'h42603a77} /* (25, 4, 30) {real, imag} */,
  {32'h41abd557, 32'hc2265b1b} /* (25, 4, 29) {real, imag} */,
  {32'h426be228, 32'h40c927a5} /* (25, 4, 28) {real, imag} */,
  {32'hc22e2681, 32'hc25c61ea} /* (25, 4, 27) {real, imag} */,
  {32'hc20a1dcd, 32'h43129870} /* (25, 4, 26) {real, imag} */,
  {32'hc10bcf98, 32'h4120ff16} /* (25, 4, 25) {real, imag} */,
  {32'hc20ba47a, 32'h4195a532} /* (25, 4, 24) {real, imag} */,
  {32'h42140cba, 32'h42527130} /* (25, 4, 23) {real, imag} */,
  {32'h41998901, 32'hc23267f2} /* (25, 4, 22) {real, imag} */,
  {32'h42538a42, 32'h4249b8a3} /* (25, 4, 21) {real, imag} */,
  {32'hc0b139ea, 32'hc15a33dc} /* (25, 4, 20) {real, imag} */,
  {32'h40817ace, 32'hc22c6fcb} /* (25, 4, 19) {real, imag} */,
  {32'hc11f25c4, 32'hc106fb52} /* (25, 4, 18) {real, imag} */,
  {32'hc0b5c55c, 32'hbfe8aa68} /* (25, 4, 17) {real, imag} */,
  {32'hc19b683d, 32'hc2064a2f} /* (25, 4, 16) {real, imag} */,
  {32'h41256228, 32'hc178d9c5} /* (25, 4, 15) {real, imag} */,
  {32'hc16e6ba4, 32'h41846977} /* (25, 4, 14) {real, imag} */,
  {32'h41b44b6c, 32'h41c5b182} /* (25, 4, 13) {real, imag} */,
  {32'hc2026253, 32'hc16d58c8} /* (25, 4, 12) {real, imag} */,
  {32'hc250b300, 32'hc184f71a} /* (25, 4, 11) {real, imag} */,
  {32'h42a5998a, 32'h414ecbf8} /* (25, 4, 10) {real, imag} */,
  {32'h42621612, 32'h40d7d64c} /* (25, 4, 9) {real, imag} */,
  {32'hc28568e7, 32'hc2a05d36} /* (25, 4, 8) {real, imag} */,
  {32'h4194a884, 32'hc26bf5b8} /* (25, 4, 7) {real, imag} */,
  {32'hbf83d580, 32'hc2bf9a90} /* (25, 4, 6) {real, imag} */,
  {32'hc2b6c438, 32'h40f5a364} /* (25, 4, 5) {real, imag} */,
  {32'h4302fbd8, 32'h408ec4ed} /* (25, 4, 4) {real, imag} */,
  {32'h419ec4f5, 32'h42c51aba} /* (25, 4, 3) {real, imag} */,
  {32'hc1efba06, 32'hc237189d} /* (25, 4, 2) {real, imag} */,
  {32'hc1d7a605, 32'hc297f762} /* (25, 4, 1) {real, imag} */,
  {32'h41bbfffd, 32'h4300b0e1} /* (25, 4, 0) {real, imag} */,
  {32'hc21aa320, 32'hc1f0a477} /* (25, 3, 31) {real, imag} */,
  {32'h41c08108, 32'h4217dfad} /* (25, 3, 30) {real, imag} */,
  {32'h41d70a8a, 32'hbdfa7400} /* (25, 3, 29) {real, imag} */,
  {32'hc2822eea, 32'h420c4ef4} /* (25, 3, 28) {real, imag} */,
  {32'hc1d6f958, 32'hc324e052} /* (25, 3, 27) {real, imag} */,
  {32'hc29071e1, 32'h40cb1190} /* (25, 3, 26) {real, imag} */,
  {32'h42566eca, 32'hc2b9e12f} /* (25, 3, 25) {real, imag} */,
  {32'h4207ff32, 32'hc1d423bb} /* (25, 3, 24) {real, imag} */,
  {32'hc2348ffc, 32'h42721f52} /* (25, 3, 23) {real, imag} */,
  {32'hc0c124c4, 32'hc1f5fb5c} /* (25, 3, 22) {real, imag} */,
  {32'hc1d4bb24, 32'hc243d6f3} /* (25, 3, 21) {real, imag} */,
  {32'hc0da6a94, 32'hc24148a0} /* (25, 3, 20) {real, imag} */,
  {32'hc0c24206, 32'hc1bf0f38} /* (25, 3, 19) {real, imag} */,
  {32'hbf8af560, 32'h4241f156} /* (25, 3, 18) {real, imag} */,
  {32'hc1abdf74, 32'hc1a54e5f} /* (25, 3, 17) {real, imag} */,
  {32'h41ce1470, 32'hc1375d30} /* (25, 3, 16) {real, imag} */,
  {32'h4124b718, 32'hbfe6b870} /* (25, 3, 15) {real, imag} */,
  {32'hc16da4dc, 32'h41bc094c} /* (25, 3, 14) {real, imag} */,
  {32'hc012bc4c, 32'hc1dc3b72} /* (25, 3, 13) {real, imag} */,
  {32'hc128797e, 32'hbe073680} /* (25, 3, 12) {real, imag} */,
  {32'h40391620, 32'h41408f40} /* (25, 3, 11) {real, imag} */,
  {32'hc224beae, 32'h42a31d1d} /* (25, 3, 10) {real, imag} */,
  {32'h42136ca8, 32'hc197544c} /* (25, 3, 9) {real, imag} */,
  {32'h417702b2, 32'hbe8fd3c0} /* (25, 3, 8) {real, imag} */,
  {32'hc2abbda9, 32'hc194f54c} /* (25, 3, 7) {real, imag} */,
  {32'h4142861a, 32'hc2fe8193} /* (25, 3, 6) {real, imag} */,
  {32'h430d5c06, 32'h41a8d59c} /* (25, 3, 5) {real, imag} */,
  {32'hc269018a, 32'h41ff5687} /* (25, 3, 4) {real, imag} */,
  {32'hc28fefb0, 32'h41c6b946} /* (25, 3, 3) {real, imag} */,
  {32'hc305a3ec, 32'h413fda7c} /* (25, 3, 2) {real, imag} */,
  {32'h416bafb6, 32'hc2371e30} /* (25, 3, 1) {real, imag} */,
  {32'hc311304e, 32'hc27b8224} /* (25, 3, 0) {real, imag} */,
  {32'h42dcf233, 32'hc2f28c85} /* (25, 2, 31) {real, imag} */,
  {32'h41623297, 32'hc3105f48} /* (25, 2, 30) {real, imag} */,
  {32'h42b6a7b6, 32'h4285fd2b} /* (25, 2, 29) {real, imag} */,
  {32'hc2b23317, 32'h43008d76} /* (25, 2, 28) {real, imag} */,
  {32'h41419120, 32'h418057b0} /* (25, 2, 27) {real, imag} */,
  {32'hc3267c09, 32'hc043fa14} /* (25, 2, 26) {real, imag} */,
  {32'hc2590a1c, 32'hc220e17f} /* (25, 2, 25) {real, imag} */,
  {32'h41edcde6, 32'h419cfd8f} /* (25, 2, 24) {real, imag} */,
  {32'h41f3924e, 32'hc117a2dc} /* (25, 2, 23) {real, imag} */,
  {32'h4286b0c6, 32'h426345cf} /* (25, 2, 22) {real, imag} */,
  {32'h3fffd500, 32'hc145317c} /* (25, 2, 21) {real, imag} */,
  {32'hc106cc9f, 32'h40f10980} /* (25, 2, 20) {real, imag} */,
  {32'hc0bd04aa, 32'h3f867000} /* (25, 2, 19) {real, imag} */,
  {32'h426b3047, 32'hc0f3842c} /* (25, 2, 18) {real, imag} */,
  {32'h41a7a674, 32'hc1ee0ad7} /* (25, 2, 17) {real, imag} */,
  {32'h419f6ae8, 32'hc1441bf8} /* (25, 2, 16) {real, imag} */,
  {32'h41d8d4b4, 32'h41d63f87} /* (25, 2, 15) {real, imag} */,
  {32'hc1009174, 32'hc0723658} /* (25, 2, 14) {real, imag} */,
  {32'hc14c8b73, 32'hc19d8cc0} /* (25, 2, 13) {real, imag} */,
  {32'hc189cd80, 32'hc295ae08} /* (25, 2, 12) {real, imag} */,
  {32'hc1a05e2d, 32'hc2237fa7} /* (25, 2, 11) {real, imag} */,
  {32'hc266c332, 32'hc29aaa75} /* (25, 2, 10) {real, imag} */,
  {32'hc225a0f1, 32'h428d376c} /* (25, 2, 9) {real, imag} */,
  {32'h427be559, 32'h421925dc} /* (25, 2, 8) {real, imag} */,
  {32'hc2f26f72, 32'h4298d1e2} /* (25, 2, 7) {real, imag} */,
  {32'h42ce9746, 32'hc10acb25} /* (25, 2, 6) {real, imag} */,
  {32'h4241a6a2, 32'hc194124a} /* (25, 2, 5) {real, imag} */,
  {32'hc1f40e94, 32'h42801cc9} /* (25, 2, 4) {real, imag} */,
  {32'h41df9a5e, 32'h42e133ab} /* (25, 2, 3) {real, imag} */,
  {32'hc1d1a5fa, 32'h41170d60} /* (25, 2, 2) {real, imag} */,
  {32'hc238847a, 32'hc1ea0a7c} /* (25, 2, 1) {real, imag} */,
  {32'hc2a16148, 32'hc354609c} /* (25, 2, 0) {real, imag} */,
  {32'hc230f503, 32'hc2826233} /* (25, 1, 31) {real, imag} */,
  {32'h41e0acf0, 32'hc3187d83} /* (25, 1, 30) {real, imag} */,
  {32'hbe41a400, 32'h4277a3e8} /* (25, 1, 29) {real, imag} */,
  {32'hc30c4383, 32'h42fe5df2} /* (25, 1, 28) {real, imag} */,
  {32'hc2b453ba, 32'hc1ace108} /* (25, 1, 27) {real, imag} */,
  {32'h421d6edc, 32'hc28cf708} /* (25, 1, 26) {real, imag} */,
  {32'hc28cd32c, 32'h410cf255} /* (25, 1, 25) {real, imag} */,
  {32'hc17aa620, 32'hc1de1d9a} /* (25, 1, 24) {real, imag} */,
  {32'h40cf1460, 32'hc20bc873} /* (25, 1, 23) {real, imag} */,
  {32'hc25f00a4, 32'h417cb691} /* (25, 1, 22) {real, imag} */,
  {32'hc201637c, 32'hc228f2a6} /* (25, 1, 21) {real, imag} */,
  {32'hc1aeed44, 32'hc10f0ae9} /* (25, 1, 20) {real, imag} */,
  {32'h41a469f8, 32'hc19ea475} /* (25, 1, 19) {real, imag} */,
  {32'h4208b74b, 32'hc1c72c8e} /* (25, 1, 18) {real, imag} */,
  {32'h4141fbbc, 32'hc03c1d68} /* (25, 1, 17) {real, imag} */,
  {32'h4152a5cc, 32'h40670cc0} /* (25, 1, 16) {real, imag} */,
  {32'h4155160c, 32'h41789016} /* (25, 1, 15) {real, imag} */,
  {32'h41b5fa3c, 32'h4108c14c} /* (25, 1, 14) {real, imag} */,
  {32'h41e2a200, 32'h41bc2a93} /* (25, 1, 13) {real, imag} */,
  {32'h40fb79d0, 32'hc215248c} /* (25, 1, 12) {real, imag} */,
  {32'h4197413f, 32'hc175de9c} /* (25, 1, 11) {real, imag} */,
  {32'h426562bc, 32'h410ef3d7} /* (25, 1, 10) {real, imag} */,
  {32'hc300646a, 32'h40de7ad6} /* (25, 1, 9) {real, imag} */,
  {32'h4296102e, 32'h41ea4e42} /* (25, 1, 8) {real, imag} */,
  {32'hc130e090, 32'hc102357b} /* (25, 1, 7) {real, imag} */,
  {32'hc173b40e, 32'hc2e5a7f4} /* (25, 1, 6) {real, imag} */,
  {32'h4272dda8, 32'hc2ceb144} /* (25, 1, 5) {real, imag} */,
  {32'h41825a50, 32'h430a016b} /* (25, 1, 4) {real, imag} */,
  {32'hc363ad8c, 32'h420570c0} /* (25, 1, 3) {real, imag} */,
  {32'h42f87328, 32'hc2a2f56c} /* (25, 1, 2) {real, imag} */,
  {32'h42b5c584, 32'h431eda18} /* (25, 1, 1) {real, imag} */,
  {32'hc2b84076, 32'h42a83466} /* (25, 1, 0) {real, imag} */,
  {32'h4279f326, 32'hc2282e00} /* (25, 0, 31) {real, imag} */,
  {32'hc21f9641, 32'h430aaf2c} /* (25, 0, 30) {real, imag} */,
  {32'h42a7b584, 32'hc228b502} /* (25, 0, 29) {real, imag} */,
  {32'h42ff8c9c, 32'hc2d8b34b} /* (25, 0, 28) {real, imag} */,
  {32'hc2c6a598, 32'h4107117c} /* (25, 0, 27) {real, imag} */,
  {32'h42ba96ff, 32'h4192b732} /* (25, 0, 26) {real, imag} */,
  {32'hc1b3f908, 32'h428b7d76} /* (25, 0, 25) {real, imag} */,
  {32'h42549b79, 32'h41e28376} /* (25, 0, 24) {real, imag} */,
  {32'hc0fb13b8, 32'hc2717f6b} /* (25, 0, 23) {real, imag} */,
  {32'hc07023e0, 32'h42075368} /* (25, 0, 22) {real, imag} */,
  {32'hc261731e, 32'h4204d8b2} /* (25, 0, 21) {real, imag} */,
  {32'h40b57ab0, 32'h42a929be} /* (25, 0, 20) {real, imag} */,
  {32'hc1f1789a, 32'hc25d05e1} /* (25, 0, 19) {real, imag} */,
  {32'h418a6950, 32'h412bb3ec} /* (25, 0, 18) {real, imag} */,
  {32'hc18bd962, 32'h41e29123} /* (25, 0, 17) {real, imag} */,
  {32'hc1afc62c, 32'h41c81116} /* (25, 0, 16) {real, imag} */,
  {32'hc2089208, 32'hc26f62b2} /* (25, 0, 15) {real, imag} */,
  {32'hc0e631b8, 32'h408de388} /* (25, 0, 14) {real, imag} */,
  {32'h4201ffd5, 32'hc00f7f30} /* (25, 0, 13) {real, imag} */,
  {32'h41fa7b08, 32'hc1a7b956} /* (25, 0, 12) {real, imag} */,
  {32'h41ca0604, 32'h41daec3d} /* (25, 0, 11) {real, imag} */,
  {32'hc2aa586f, 32'h3ebfe9c0} /* (25, 0, 10) {real, imag} */,
  {32'hc204bddb, 32'h41543624} /* (25, 0, 9) {real, imag} */,
  {32'h4223400b, 32'hc28f8840} /* (25, 0, 8) {real, imag} */,
  {32'h4183d19c, 32'h3e4bf100} /* (25, 0, 7) {real, imag} */,
  {32'h42f4548f, 32'h422fb117} /* (25, 0, 6) {real, imag} */,
  {32'hc1c76b98, 32'hc2c7ff14} /* (25, 0, 5) {real, imag} */,
  {32'hc23de0d1, 32'hc318a2ff} /* (25, 0, 4) {real, imag} */,
  {32'hc21b49ee, 32'hc22476e2} /* (25, 0, 3) {real, imag} */,
  {32'hc191f5cc, 32'hc1fc1190} /* (25, 0, 2) {real, imag} */,
  {32'hbe8f3380, 32'hc2a86026} /* (25, 0, 1) {real, imag} */,
  {32'hc0f50dc8, 32'h431453f1} /* (25, 0, 0) {real, imag} */,
  {32'hc4313580, 32'hc3216347} /* (24, 31, 31) {real, imag} */,
  {32'h43f48a1b, 32'h4282d6c2} /* (24, 31, 30) {real, imag} */,
  {32'h4234954a, 32'hc245f0d7} /* (24, 31, 29) {real, imag} */,
  {32'h4205f8fa, 32'h43236678} /* (24, 31, 28) {real, imag} */,
  {32'h434bd740, 32'h419dcd9c} /* (24, 31, 27) {real, imag} */,
  {32'h4243b905, 32'hc2248400} /* (24, 31, 26) {real, imag} */,
  {32'hc3215287, 32'h41c1ac90} /* (24, 31, 25) {real, imag} */,
  {32'h42fbacfd, 32'hc1466820} /* (24, 31, 24) {real, imag} */,
  {32'h3f997d60, 32'h427b58d0} /* (24, 31, 23) {real, imag} */,
  {32'hbf1b39c0, 32'hc2592a1c} /* (24, 31, 22) {real, imag} */,
  {32'h413f431c, 32'hc1b422d2} /* (24, 31, 21) {real, imag} */,
  {32'hc22706c3, 32'h42a30ef6} /* (24, 31, 20) {real, imag} */,
  {32'hc1b42600, 32'hc09ecb4c} /* (24, 31, 19) {real, imag} */,
  {32'h41678a78, 32'hc1719124} /* (24, 31, 18) {real, imag} */,
  {32'h4020b400, 32'hc15a0b40} /* (24, 31, 17) {real, imag} */,
  {32'h40ab6220, 32'hbff8b480} /* (24, 31, 16) {real, imag} */,
  {32'h40f0be00, 32'hc0e40e40} /* (24, 31, 15) {real, imag} */,
  {32'h41fa4d1c, 32'h41715b24} /* (24, 31, 14) {real, imag} */,
  {32'hc24a363c, 32'hc09e383c} /* (24, 31, 13) {real, imag} */,
  {32'hc2366bad, 32'h42306e39} /* (24, 31, 12) {real, imag} */,
  {32'hc1c31106, 32'h42d52058} /* (24, 31, 11) {real, imag} */,
  {32'hc24a442d, 32'hc158ba80} /* (24, 31, 10) {real, imag} */,
  {32'hc022dbb0, 32'hc2549d80} /* (24, 31, 9) {real, imag} */,
  {32'hc1ccea3c, 32'h42f46810} /* (24, 31, 8) {real, imag} */,
  {32'hc30e31fd, 32'hc11eb520} /* (24, 31, 7) {real, imag} */,
  {32'hc2603869, 32'hc266a1e0} /* (24, 31, 6) {real, imag} */,
  {32'h42c84090, 32'h42f42c6f} /* (24, 31, 5) {real, imag} */,
  {32'hc2619988, 32'h42488f35} /* (24, 31, 4) {real, imag} */,
  {32'h40e25fcc, 32'hc24f5e9d} /* (24, 31, 3) {real, imag} */,
  {32'hc1e35c30, 32'h43487fc7} /* (24, 31, 2) {real, imag} */,
  {32'hc3a97cdc, 32'hc3ef71d8} /* (24, 31, 1) {real, imag} */,
  {32'hc3835188, 32'hc3a391f8} /* (24, 31, 0) {real, imag} */,
  {32'h439cc651, 32'h43a23a85} /* (24, 30, 31) {real, imag} */,
  {32'hc295c910, 32'hc3117414} /* (24, 30, 30) {real, imag} */,
  {32'h4172692c, 32'h42505156} /* (24, 30, 29) {real, imag} */,
  {32'h431d287b, 32'h431793b3} /* (24, 30, 28) {real, imag} */,
  {32'hc31aaca2, 32'h42514d8c} /* (24, 30, 27) {real, imag} */,
  {32'h4294515e, 32'hc1516a1a} /* (24, 30, 26) {real, imag} */,
  {32'h41c003d7, 32'h41201158} /* (24, 30, 25) {real, imag} */,
  {32'hc302524c, 32'hc1fffc14} /* (24, 30, 24) {real, imag} */,
  {32'hc25e4638, 32'hc0fb36d0} /* (24, 30, 23) {real, imag} */,
  {32'hc19b4e91, 32'h4184dee9} /* (24, 30, 22) {real, imag} */,
  {32'hc297fb54, 32'h42869a5e} /* (24, 30, 21) {real, imag} */,
  {32'hc1b73dbb, 32'h408970d8} /* (24, 30, 20) {real, imag} */,
  {32'hc07baee0, 32'h41e8c454} /* (24, 30, 19) {real, imag} */,
  {32'hc21b1bcb, 32'hc18c7f6c} /* (24, 30, 18) {real, imag} */,
  {32'hbcab3000, 32'hc21cd500} /* (24, 30, 17) {real, imag} */,
  {32'hc19d1f50, 32'hbfeef380} /* (24, 30, 16) {real, imag} */,
  {32'hc21cb4aa, 32'hc1358e42} /* (24, 30, 15) {real, imag} */,
  {32'hc0e3c328, 32'hc0a10d90} /* (24, 30, 14) {real, imag} */,
  {32'hc1b79892, 32'h411ea2f3} /* (24, 30, 13) {real, imag} */,
  {32'h41835735, 32'h41cfeb76} /* (24, 30, 12) {real, imag} */,
  {32'h40113e50, 32'hc12f9d40} /* (24, 30, 11) {real, imag} */,
  {32'h41cac527, 32'h40622378} /* (24, 30, 10) {real, imag} */,
  {32'h415485c2, 32'hc1cc55cc} /* (24, 30, 9) {real, imag} */,
  {32'h3ea52b00, 32'hc2eca7a3} /* (24, 30, 8) {real, imag} */,
  {32'h420e8564, 32'h41e47d54} /* (24, 30, 7) {real, imag} */,
  {32'hc1ef4267, 32'hc256f146} /* (24, 30, 6) {real, imag} */,
  {32'hc18c42d4, 32'h41425716} /* (24, 30, 5) {real, imag} */,
  {32'hc206e064, 32'h420fa7dc} /* (24, 30, 4) {real, imag} */,
  {32'hc229269e, 32'h42b1f4f1} /* (24, 30, 3) {real, imag} */,
  {32'hc38b5d14, 32'hc3a6623d} /* (24, 30, 2) {real, imag} */,
  {32'h43ec60dd, 32'h43a3915d} /* (24, 30, 1) {real, imag} */,
  {32'h439f12bb, 32'h434ab2e5} /* (24, 30, 0) {real, imag} */,
  {32'hc31b9b82, 32'hc1d86e54} /* (24, 29, 31) {real, imag} */,
  {32'h431a5ab8, 32'hc1c2288c} /* (24, 29, 30) {real, imag} */,
  {32'h421abb78, 32'h41760221} /* (24, 29, 29) {real, imag} */,
  {32'h42655dc1, 32'h423038ac} /* (24, 29, 28) {real, imag} */,
  {32'h420e52dc, 32'hc1bb442d} /* (24, 29, 27) {real, imag} */,
  {32'hc26bd1f4, 32'hc22cfb82} /* (24, 29, 26) {real, imag} */,
  {32'hc1189e24, 32'h42b58a0a} /* (24, 29, 25) {real, imag} */,
  {32'h42294e9f, 32'hc2a30b08} /* (24, 29, 24) {real, imag} */,
  {32'hc2bb2927, 32'hc2adc707} /* (24, 29, 23) {real, imag} */,
  {32'h421c98df, 32'h424872c4} /* (24, 29, 22) {real, imag} */,
  {32'h42169d26, 32'h41c7cc70} /* (24, 29, 21) {real, imag} */,
  {32'h41e84b5c, 32'h41d5d845} /* (24, 29, 20) {real, imag} */,
  {32'hc1f2870c, 32'h41a1cd8a} /* (24, 29, 19) {real, imag} */,
  {32'hc1add719, 32'h40d40a90} /* (24, 29, 18) {real, imag} */,
  {32'hc0f603ce, 32'h41ef5961} /* (24, 29, 17) {real, imag} */,
  {32'h411d05ac, 32'hc217e272} /* (24, 29, 16) {real, imag} */,
  {32'hc21ccd00, 32'h4114ad9a} /* (24, 29, 15) {real, imag} */,
  {32'h3fb413d0, 32'hc224eec6} /* (24, 29, 14) {real, imag} */,
  {32'hc23ec5d6, 32'h4202b6a5} /* (24, 29, 13) {real, imag} */,
  {32'h4233fb08, 32'h41c42d83} /* (24, 29, 12) {real, imag} */,
  {32'h420abe06, 32'hc2017ebc} /* (24, 29, 11) {real, imag} */,
  {32'h429abe98, 32'hc1b17968} /* (24, 29, 10) {real, imag} */,
  {32'hc04da3a0, 32'hc0f27100} /* (24, 29, 9) {real, imag} */,
  {32'hc1facf7a, 32'h42ccd6ee} /* (24, 29, 8) {real, imag} */,
  {32'hc1f763fc, 32'hc235d019} /* (24, 29, 7) {real, imag} */,
  {32'hc21af31e, 32'hc291e48f} /* (24, 29, 6) {real, imag} */,
  {32'hc1eebb00, 32'h41c1fdc7} /* (24, 29, 5) {real, imag} */,
  {32'hc2ec0b64, 32'hc23c5698} /* (24, 29, 4) {real, imag} */,
  {32'h4301d463, 32'h40c0294e} /* (24, 29, 3) {real, imag} */,
  {32'h4268dcd8, 32'hc27af75e} /* (24, 29, 2) {real, imag} */,
  {32'hc2883d50, 32'h43227250} /* (24, 29, 1) {real, imag} */,
  {32'hc2843b3c, 32'h4278795a} /* (24, 29, 0) {real, imag} */,
  {32'hc357030a, 32'hc2c03634} /* (24, 28, 31) {real, imag} */,
  {32'h434b5179, 32'h428137a6} /* (24, 28, 30) {real, imag} */,
  {32'h41ebffde, 32'hc25ebeab} /* (24, 28, 29) {real, imag} */,
  {32'hc27347f0, 32'h433785ca} /* (24, 28, 28) {real, imag} */,
  {32'h42299cff, 32'hc04cdf3e} /* (24, 28, 27) {real, imag} */,
  {32'h425920ba, 32'h42bf7271} /* (24, 28, 26) {real, imag} */,
  {32'hc313c194, 32'hc1a04418} /* (24, 28, 25) {real, imag} */,
  {32'h429a4c05, 32'h42f6bff0} /* (24, 28, 24) {real, imag} */,
  {32'hc26e023c, 32'hc21b456d} /* (24, 28, 23) {real, imag} */,
  {32'h40ba8f9c, 32'h42738494} /* (24, 28, 22) {real, imag} */,
  {32'hc192852e, 32'h422cb05c} /* (24, 28, 21) {real, imag} */,
  {32'h4064a024, 32'hc21026d2} /* (24, 28, 20) {real, imag} */,
  {32'hc246ccce, 32'hc22317ea} /* (24, 28, 19) {real, imag} */,
  {32'hc1abead2, 32'hc1a06d7a} /* (24, 28, 18) {real, imag} */,
  {32'hc0037800, 32'h41720e66} /* (24, 28, 17) {real, imag} */,
  {32'h41fc2685, 32'h413b59b6} /* (24, 28, 16) {real, imag} */,
  {32'hc14007a0, 32'hc1c7bf45} /* (24, 28, 15) {real, imag} */,
  {32'h42242e99, 32'hc1a9ff2e} /* (24, 28, 14) {real, imag} */,
  {32'h41ac3504, 32'h402bab88} /* (24, 28, 13) {real, imag} */,
  {32'hc16f0afd, 32'hbfd80d40} /* (24, 28, 12) {real, imag} */,
  {32'h422d980d, 32'hc161765e} /* (24, 28, 11) {real, imag} */,
  {32'h40fa7cdc, 32'h40f2d930} /* (24, 28, 10) {real, imag} */,
  {32'hc2159e20, 32'h41a098b0} /* (24, 28, 9) {real, imag} */,
  {32'h4231d532, 32'h409d84c8} /* (24, 28, 8) {real, imag} */,
  {32'h42a315c7, 32'h42077653} /* (24, 28, 7) {real, imag} */,
  {32'hc22a9146, 32'h429d1a73} /* (24, 28, 6) {real, imag} */,
  {32'h41a24a4e, 32'h402e3ada} /* (24, 28, 5) {real, imag} */,
  {32'hc19bd3e8, 32'hc1ed35d0} /* (24, 28, 4) {real, imag} */,
  {32'h427994fb, 32'h4242dfcb} /* (24, 28, 3) {real, imag} */,
  {32'h4347cff7, 32'h4167bea4} /* (24, 28, 2) {real, imag} */,
  {32'hc2bcbd9f, 32'h42b806ce} /* (24, 28, 1) {real, imag} */,
  {32'hc1b477cf, 32'h419436ed} /* (24, 28, 0) {real, imag} */,
  {32'h429ff62f, 32'hc223f96a} /* (24, 27, 31) {real, imag} */,
  {32'hc28e355c, 32'h428335f3} /* (24, 27, 30) {real, imag} */,
  {32'h4261348c, 32'h425c8906} /* (24, 27, 29) {real, imag} */,
  {32'h427fb484, 32'hc2fdc3ea} /* (24, 27, 28) {real, imag} */,
  {32'h42be695a, 32'hc2914fbd} /* (24, 27, 27) {real, imag} */,
  {32'hc234e071, 32'hbec280e0} /* (24, 27, 26) {real, imag} */,
  {32'h40fce990, 32'hc20fd000} /* (24, 27, 25) {real, imag} */,
  {32'hc1d4f721, 32'hc1149f8a} /* (24, 27, 24) {real, imag} */,
  {32'hc209780a, 32'hc02b6217} /* (24, 27, 23) {real, imag} */,
  {32'h41305d72, 32'h419a795c} /* (24, 27, 22) {real, imag} */,
  {32'h426c5d1d, 32'h42075eab} /* (24, 27, 21) {real, imag} */,
  {32'h418239d2, 32'hc0bee264} /* (24, 27, 20) {real, imag} */,
  {32'hc1b792a6, 32'h421cb29f} /* (24, 27, 19) {real, imag} */,
  {32'hc13ae7e8, 32'h421ba846} /* (24, 27, 18) {real, imag} */,
  {32'h4209ac5e, 32'hc16189e0} /* (24, 27, 17) {real, imag} */,
  {32'h40fdcf70, 32'hc14f4100} /* (24, 27, 16) {real, imag} */,
  {32'hc1062daa, 32'h3fd6e380} /* (24, 27, 15) {real, imag} */,
  {32'h4140f5b8, 32'hc14e38fa} /* (24, 27, 14) {real, imag} */,
  {32'hc1555828, 32'hc19a7fb0} /* (24, 27, 13) {real, imag} */,
  {32'hc15c88c3, 32'hc14d045a} /* (24, 27, 12) {real, imag} */,
  {32'hc1b6bef6, 32'h40a00c8a} /* (24, 27, 11) {real, imag} */,
  {32'hc0b23544, 32'hc275521a} /* (24, 27, 10) {real, imag} */,
  {32'h41b45bac, 32'h3fd39b32} /* (24, 27, 9) {real, imag} */,
  {32'h4208b99a, 32'h41b97843} /* (24, 27, 8) {real, imag} */,
  {32'h423c137c, 32'h421bb7a4} /* (24, 27, 7) {real, imag} */,
  {32'h421a3f53, 32'h406a7894} /* (24, 27, 6) {real, imag} */,
  {32'h421526bc, 32'hc26bd36a} /* (24, 27, 5) {real, imag} */,
  {32'h42bcf31e, 32'hc0bbb398} /* (24, 27, 4) {real, imag} */,
  {32'h41c046a9, 32'h4168c066} /* (24, 27, 3) {real, imag} */,
  {32'hc2bf1f12, 32'hc287b3e3} /* (24, 27, 2) {real, imag} */,
  {32'h42ee5e3b, 32'h43390852} /* (24, 27, 1) {real, imag} */,
  {32'h432e1eac, 32'h42a147a2} /* (24, 27, 0) {real, imag} */,
  {32'h428f939a, 32'hc182bf92} /* (24, 26, 31) {real, imag} */,
  {32'h41b80334, 32'h418e5b32} /* (24, 26, 30) {real, imag} */,
  {32'hc23e4158, 32'hc2aea4d6} /* (24, 26, 29) {real, imag} */,
  {32'h40554fe8, 32'h415b733a} /* (24, 26, 28) {real, imag} */,
  {32'h4223f851, 32'h4216182e} /* (24, 26, 27) {real, imag} */,
  {32'hc2449e06, 32'h41aa8e3e} /* (24, 26, 26) {real, imag} */,
  {32'hc26d95d8, 32'hc22657a6} /* (24, 26, 25) {real, imag} */,
  {32'hc24e4518, 32'h42a69b9a} /* (24, 26, 24) {real, imag} */,
  {32'h40db210e, 32'h42aaf63a} /* (24, 26, 23) {real, imag} */,
  {32'hc1e86803, 32'hc12af14c} /* (24, 26, 22) {real, imag} */,
  {32'h40a70466, 32'hc1eb94e7} /* (24, 26, 21) {real, imag} */,
  {32'h41f04c91, 32'h41a66fa6} /* (24, 26, 20) {real, imag} */,
  {32'hc111f26b, 32'h41b1e7c6} /* (24, 26, 19) {real, imag} */,
  {32'h404f2e84, 32'hbfefffb8} /* (24, 26, 18) {real, imag} */,
  {32'h40ec0508, 32'h4023d580} /* (24, 26, 17) {real, imag} */,
  {32'hc162fe1b, 32'h4135b414} /* (24, 26, 16) {real, imag} */,
  {32'h4245dc67, 32'hc19a6a68} /* (24, 26, 15) {real, imag} */,
  {32'h4070ce9c, 32'h41dc05a4} /* (24, 26, 14) {real, imag} */,
  {32'hc15aad03, 32'h41504dd4} /* (24, 26, 13) {real, imag} */,
  {32'h40aefd9c, 32'h4208796e} /* (24, 26, 12) {real, imag} */,
  {32'hc1319235, 32'h40357ac8} /* (24, 26, 11) {real, imag} */,
  {32'h418e9949, 32'hc198be8e} /* (24, 26, 10) {real, imag} */,
  {32'h41967af4, 32'hc1aa04aa} /* (24, 26, 9) {real, imag} */,
  {32'h411f2506, 32'h41da051a} /* (24, 26, 8) {real, imag} */,
  {32'h42b29774, 32'hc1ffab29} /* (24, 26, 7) {real, imag} */,
  {32'hc1ecb41c, 32'h42912e6c} /* (24, 26, 6) {real, imag} */,
  {32'hc25a0c09, 32'hc252e16e} /* (24, 26, 5) {real, imag} */,
  {32'hc26a1e48, 32'hc23f4ef0} /* (24, 26, 4) {real, imag} */,
  {32'h42c46c78, 32'h42b232b6} /* (24, 26, 3) {real, imag} */,
  {32'h42a7c062, 32'hc286cc9a} /* (24, 26, 2) {real, imag} */,
  {32'h430454e9, 32'h421d5d33} /* (24, 26, 1) {real, imag} */,
  {32'hc13c72d9, 32'h42997dd2} /* (24, 26, 0) {real, imag} */,
  {32'h4232d6e3, 32'h432115f5} /* (24, 25, 31) {real, imag} */,
  {32'h3f003d80, 32'h40b5d82a} /* (24, 25, 30) {real, imag} */,
  {32'hc2bc07ad, 32'hc2a0b01d} /* (24, 25, 29) {real, imag} */,
  {32'hc1c53914, 32'hc26ac514} /* (24, 25, 28) {real, imag} */,
  {32'h42834172, 32'hc267f041} /* (24, 25, 27) {real, imag} */,
  {32'hc24ef330, 32'hc1597440} /* (24, 25, 26) {real, imag} */,
  {32'hc2146562, 32'hc2282370} /* (24, 25, 25) {real, imag} */,
  {32'h410c9297, 32'hc2b7d7cf} /* (24, 25, 24) {real, imag} */,
  {32'h41a1d4ec, 32'h4200bb78} /* (24, 25, 23) {real, imag} */,
  {32'h401ffe08, 32'hc0d838fd} /* (24, 25, 22) {real, imag} */,
  {32'h424a3e95, 32'h40efc252} /* (24, 25, 21) {real, imag} */,
  {32'hc0bce188, 32'hc0da6c8c} /* (24, 25, 20) {real, imag} */,
  {32'hc1ee42fd, 32'h4189774d} /* (24, 25, 19) {real, imag} */,
  {32'h41dea41e, 32'hc18b848a} /* (24, 25, 18) {real, imag} */,
  {32'hc028efd0, 32'h40b98fa8} /* (24, 25, 17) {real, imag} */,
  {32'h40afa420, 32'hc0a2dd88} /* (24, 25, 16) {real, imag} */,
  {32'h4113d6dc, 32'hc19c1352} /* (24, 25, 15) {real, imag} */,
  {32'h3ffb0c60, 32'h41c31e02} /* (24, 25, 14) {real, imag} */,
  {32'h402defc8, 32'hbdcbe500} /* (24, 25, 13) {real, imag} */,
  {32'h40fc1854, 32'h3f55b5e0} /* (24, 25, 12) {real, imag} */,
  {32'hc2166b53, 32'hc1f5dd58} /* (24, 25, 11) {real, imag} */,
  {32'h422f10c6, 32'h413b7e06} /* (24, 25, 10) {real, imag} */,
  {32'hc10a1d6d, 32'h40b3f560} /* (24, 25, 9) {real, imag} */,
  {32'hc1a990c0, 32'h4186e93c} /* (24, 25, 8) {real, imag} */,
  {32'h3fadb390, 32'hc27a5ed4} /* (24, 25, 7) {real, imag} */,
  {32'h41eb30e8, 32'h42402643} /* (24, 25, 6) {real, imag} */,
  {32'hc20cb2c1, 32'h4088a1f8} /* (24, 25, 5) {real, imag} */,
  {32'h41c22aac, 32'hc150d1b6} /* (24, 25, 4) {real, imag} */,
  {32'hc290b20f, 32'h417d7c28} /* (24, 25, 3) {real, imag} */,
  {32'hc0cd717e, 32'h41abf0a2} /* (24, 25, 2) {real, imag} */,
  {32'hc2e0d0ac, 32'h423a4477} /* (24, 25, 1) {real, imag} */,
  {32'h423ead20, 32'hc2b1346e} /* (24, 25, 0) {real, imag} */,
  {32'h41d0da43, 32'hc20d6531} /* (24, 24, 31) {real, imag} */,
  {32'hc34cca1c, 32'hc0ecca48} /* (24, 24, 30) {real, imag} */,
  {32'hc0de06d0, 32'h4222d355} /* (24, 24, 29) {real, imag} */,
  {32'h42909f43, 32'h4311f9ca} /* (24, 24, 28) {real, imag} */,
  {32'h41fe6b80, 32'h42046440} /* (24, 24, 27) {real, imag} */,
  {32'h421ff534, 32'h42085d2a} /* (24, 24, 26) {real, imag} */,
  {32'hc238652b, 32'hc13db594} /* (24, 24, 25) {real, imag} */,
  {32'hc1a40a50, 32'h424e9d0a} /* (24, 24, 24) {real, imag} */,
  {32'h4294239a, 32'h423de149} /* (24, 24, 23) {real, imag} */,
  {32'h42325bf2, 32'hc22ef87a} /* (24, 24, 22) {real, imag} */,
  {32'hc24d66f4, 32'h40239e38} /* (24, 24, 21) {real, imag} */,
  {32'h409777fc, 32'hc051ef9c} /* (24, 24, 20) {real, imag} */,
  {32'hc15c4704, 32'h409b75dc} /* (24, 24, 19) {real, imag} */,
  {32'hc1faa60c, 32'hc2377312} /* (24, 24, 18) {real, imag} */,
  {32'h419e967b, 32'h3ffc8080} /* (24, 24, 17) {real, imag} */,
  {32'h4173fc7c, 32'h42088aca} /* (24, 24, 16) {real, imag} */,
  {32'hc10fdf7e, 32'hbf8de700} /* (24, 24, 15) {real, imag} */,
  {32'h4108df88, 32'hc0160a00} /* (24, 24, 14) {real, imag} */,
  {32'hc0b2e290, 32'h413863ee} /* (24, 24, 13) {real, imag} */,
  {32'hc147606e, 32'hc0fa9cf2} /* (24, 24, 12) {real, imag} */,
  {32'h41e62d29, 32'hc1f4a4db} /* (24, 24, 11) {real, imag} */,
  {32'hc0a1585c, 32'hc265d3ca} /* (24, 24, 10) {real, imag} */,
  {32'hc1659144, 32'h42477157} /* (24, 24, 9) {real, imag} */,
  {32'hc2085151, 32'h41d6785c} /* (24, 24, 8) {real, imag} */,
  {32'h3e586100, 32'h42a30582} /* (24, 24, 7) {real, imag} */,
  {32'hc1b0eac9, 32'h42527212} /* (24, 24, 6) {real, imag} */,
  {32'hc1add5de, 32'h41839993} /* (24, 24, 5) {real, imag} */,
  {32'h42b7142b, 32'h42a9aeb0} /* (24, 24, 4) {real, imag} */,
  {32'h4247e383, 32'h42a5dad2} /* (24, 24, 3) {real, imag} */,
  {32'h41f19fc4, 32'hc23e492f} /* (24, 24, 2) {real, imag} */,
  {32'h429e88be, 32'h41c8c846} /* (24, 24, 1) {real, imag} */,
  {32'h426f2b45, 32'hc167523f} /* (24, 24, 0) {real, imag} */,
  {32'hc214c43d, 32'h408ea624} /* (24, 23, 31) {real, imag} */,
  {32'hc0f24de1, 32'hc1146df4} /* (24, 23, 30) {real, imag} */,
  {32'h42802a0b, 32'h42ac41ea} /* (24, 23, 29) {real, imag} */,
  {32'hc21e7769, 32'hc26a0318} /* (24, 23, 28) {real, imag} */,
  {32'hc1823921, 32'h4189184e} /* (24, 23, 27) {real, imag} */,
  {32'hc1cf5313, 32'hc128f4f2} /* (24, 23, 26) {real, imag} */,
  {32'hc084e101, 32'hc088aef9} /* (24, 23, 25) {real, imag} */,
  {32'h418af769, 32'h418da96e} /* (24, 23, 24) {real, imag} */,
  {32'hc21fb036, 32'hc1e62902} /* (24, 23, 23) {real, imag} */,
  {32'h410ef536, 32'hc1d20ff9} /* (24, 23, 22) {real, imag} */,
  {32'hc0a373a0, 32'h41664917} /* (24, 23, 21) {real, imag} */,
  {32'h420410f1, 32'hc19feadf} /* (24, 23, 20) {real, imag} */,
  {32'h41fdd08c, 32'h400bfd38} /* (24, 23, 19) {real, imag} */,
  {32'h3e49b380, 32'h409f9914} /* (24, 23, 18) {real, imag} */,
  {32'h4183c82e, 32'hc1944432} /* (24, 23, 17) {real, imag} */,
  {32'hc07bad50, 32'h4122a102} /* (24, 23, 16) {real, imag} */,
  {32'h41a2ab2a, 32'hc0563c84} /* (24, 23, 15) {real, imag} */,
  {32'hc196478f, 32'h3f9417b0} /* (24, 23, 14) {real, imag} */,
  {32'h41bc2054, 32'hc215ddb2} /* (24, 23, 13) {real, imag} */,
  {32'h411a7718, 32'hc0c31374} /* (24, 23, 12) {real, imag} */,
  {32'hc193ca10, 32'h412946f7} /* (24, 23, 11) {real, imag} */,
  {32'h409da6b4, 32'hc0c719a4} /* (24, 23, 10) {real, imag} */,
  {32'h41995e5b, 32'h421a2e93} /* (24, 23, 9) {real, imag} */,
  {32'hc0c19d2c, 32'hc1d1a810} /* (24, 23, 8) {real, imag} */,
  {32'h4148d430, 32'h408c0b4f} /* (24, 23, 7) {real, imag} */,
  {32'h417bcace, 32'hc245f398} /* (24, 23, 6) {real, imag} */,
  {32'h419ab56f, 32'hc1f32cec} /* (24, 23, 5) {real, imag} */,
  {32'hc279e7af, 32'h420475f8} /* (24, 23, 4) {real, imag} */,
  {32'h41836ff4, 32'h41f6c203} /* (24, 23, 3) {real, imag} */,
  {32'hc1256978, 32'h429f1ed6} /* (24, 23, 2) {real, imag} */,
  {32'hc26f0cf7, 32'h424c1c16} /* (24, 23, 1) {real, imag} */,
  {32'hc26bee84, 32'h42084316} /* (24, 23, 0) {real, imag} */,
  {32'hc1aaa4cf, 32'hc21718a4} /* (24, 22, 31) {real, imag} */,
  {32'h428d31e5, 32'h3eb72640} /* (24, 22, 30) {real, imag} */,
  {32'hc25dba6a, 32'h4128c09e} /* (24, 22, 29) {real, imag} */,
  {32'hc0e709d4, 32'h407f4c74} /* (24, 22, 28) {real, imag} */,
  {32'h41585a60, 32'hc0843a28} /* (24, 22, 27) {real, imag} */,
  {32'hc1e232d8, 32'h42133d87} /* (24, 22, 26) {real, imag} */,
  {32'hbf67f090, 32'h41fbef28} /* (24, 22, 25) {real, imag} */,
  {32'hc1d5cddc, 32'hc1328a00} /* (24, 22, 24) {real, imag} */,
  {32'h418e60d4, 32'hc0375aba} /* (24, 22, 23) {real, imag} */,
  {32'h42070832, 32'h41812024} /* (24, 22, 22) {real, imag} */,
  {32'h413a8d64, 32'h40042ac4} /* (24, 22, 21) {real, imag} */,
  {32'hc1543bca, 32'hbfb2a32e} /* (24, 22, 20) {real, imag} */,
  {32'h3f8f9528, 32'hc1a620e8} /* (24, 22, 19) {real, imag} */,
  {32'hc150f670, 32'hc01ae49c} /* (24, 22, 18) {real, imag} */,
  {32'h413e805e, 32'h40e54d9d} /* (24, 22, 17) {real, imag} */,
  {32'hbffc9b60, 32'h402accf9} /* (24, 22, 16) {real, imag} */,
  {32'h40bf94b4, 32'h40f39835} /* (24, 22, 15) {real, imag} */,
  {32'h3f864080, 32'h40c6701e} /* (24, 22, 14) {real, imag} */,
  {32'h41884b38, 32'hc17f6ec4} /* (24, 22, 13) {real, imag} */,
  {32'hc0982cd4, 32'hc065fc7f} /* (24, 22, 12) {real, imag} */,
  {32'h418b5ca8, 32'h405a751c} /* (24, 22, 11) {real, imag} */,
  {32'h40714bf4, 32'h40a9de56} /* (24, 22, 10) {real, imag} */,
  {32'hc1dca146, 32'h417a51de} /* (24, 22, 9) {real, imag} */,
  {32'h4162b68c, 32'h40b19a08} /* (24, 22, 8) {real, imag} */,
  {32'hbf3e5950, 32'h40671080} /* (24, 22, 7) {real, imag} */,
  {32'hc0877956, 32'hbf8ce5e0} /* (24, 22, 6) {real, imag} */,
  {32'h40899600, 32'h41da3243} /* (24, 22, 5) {real, imag} */,
  {32'hc1bbdc9d, 32'hc1c3926c} /* (24, 22, 4) {real, imag} */,
  {32'h40e86664, 32'hc0c110b4} /* (24, 22, 3) {real, imag} */,
  {32'h40ba3b70, 32'hc229394e} /* (24, 22, 2) {real, imag} */,
  {32'hc27c76e2, 32'h4296ae3c} /* (24, 22, 1) {real, imag} */,
  {32'hc22c02fe, 32'hbfe51cae} /* (24, 22, 0) {real, imag} */,
  {32'h418703ff, 32'hc1a1334a} /* (24, 21, 31) {real, imag} */,
  {32'hc22713f8, 32'h4281d91e} /* (24, 21, 30) {real, imag} */,
  {32'h41bd987f, 32'h422fa454} /* (24, 21, 29) {real, imag} */,
  {32'h42063513, 32'h41efebdf} /* (24, 21, 28) {real, imag} */,
  {32'hc1f931a4, 32'hc137917a} /* (24, 21, 27) {real, imag} */,
  {32'h42020966, 32'h41168eae} /* (24, 21, 26) {real, imag} */,
  {32'hc21d48c2, 32'hc1a6cf54} /* (24, 21, 25) {real, imag} */,
  {32'hc1db142e, 32'h41d0fafd} /* (24, 21, 24) {real, imag} */,
  {32'h419e3051, 32'h41821352} /* (24, 21, 23) {real, imag} */,
  {32'hc21175c0, 32'hc1cc521b} /* (24, 21, 22) {real, imag} */,
  {32'hc0cdff41, 32'hc1c2d84b} /* (24, 21, 21) {real, imag} */,
  {32'hc16ddf97, 32'h3f53f920} /* (24, 21, 20) {real, imag} */,
  {32'hc19d83a1, 32'h41316945} /* (24, 21, 19) {real, imag} */,
  {32'h409878db, 32'h41a6fd97} /* (24, 21, 18) {real, imag} */,
  {32'h3f6c92c0, 32'hc11c6d25} /* (24, 21, 17) {real, imag} */,
  {32'h40341658, 32'hc079f678} /* (24, 21, 16) {real, imag} */,
  {32'hc1239268, 32'hbfd372f8} /* (24, 21, 15) {real, imag} */,
  {32'hc0864485, 32'hc0ae282c} /* (24, 21, 14) {real, imag} */,
  {32'h40cee79c, 32'h40b1d0ba} /* (24, 21, 13) {real, imag} */,
  {32'h404b911c, 32'hc187fb37} /* (24, 21, 12) {real, imag} */,
  {32'hc025a0ce, 32'hc14687b2} /* (24, 21, 11) {real, imag} */,
  {32'h418960eb, 32'hc12231a2} /* (24, 21, 10) {real, imag} */,
  {32'hc0886ff4, 32'h41716185} /* (24, 21, 9) {real, imag} */,
  {32'h4012716c, 32'hc1c6dfb7} /* (24, 21, 8) {real, imag} */,
  {32'hc1b328c5, 32'h41991faa} /* (24, 21, 7) {real, imag} */,
  {32'h41fa886b, 32'hc1579606} /* (24, 21, 6) {real, imag} */,
  {32'hc155e544, 32'h424917fa} /* (24, 21, 5) {real, imag} */,
  {32'h4164fb11, 32'h4262c010} /* (24, 21, 4) {real, imag} */,
  {32'h3eaf0cc0, 32'hc18fc4f0} /* (24, 21, 3) {real, imag} */,
  {32'h41880a27, 32'hc1635e0c} /* (24, 21, 2) {real, imag} */,
  {32'h429d84ea, 32'hc20f4b96} /* (24, 21, 1) {real, imag} */,
  {32'h420471a4, 32'hc26fcce2} /* (24, 21, 0) {real, imag} */,
  {32'hc1921fea, 32'h40c421f8} /* (24, 20, 31) {real, imag} */,
  {32'hc1402fa5, 32'h409a1ef8} /* (24, 20, 30) {real, imag} */,
  {32'h3f241e60, 32'h41ee5a05} /* (24, 20, 29) {real, imag} */,
  {32'hc18a7f14, 32'hc1d2f634} /* (24, 20, 28) {real, imag} */,
  {32'h41cb7d0e, 32'h420ff9a2} /* (24, 20, 27) {real, imag} */,
  {32'h40ca51b0, 32'h418a8d50} /* (24, 20, 26) {real, imag} */,
  {32'h4216fa63, 32'hc2312785} /* (24, 20, 25) {real, imag} */,
  {32'h40a22de8, 32'hc2619ecd} /* (24, 20, 24) {real, imag} */,
  {32'h40cfd2bf, 32'h4116b8b6} /* (24, 20, 23) {real, imag} */,
  {32'hc1df7235, 32'hbfa37cc0} /* (24, 20, 22) {real, imag} */,
  {32'hc0158832, 32'hc13e71ca} /* (24, 20, 21) {real, imag} */,
  {32'h40824c0c, 32'hbf58ff60} /* (24, 20, 20) {real, imag} */,
  {32'hc0ce7142, 32'h41447b40} /* (24, 20, 19) {real, imag} */,
  {32'hc10a3fbf, 32'h400d0968} /* (24, 20, 18) {real, imag} */,
  {32'h3eff6ae0, 32'h41cfdb9d} /* (24, 20, 17) {real, imag} */,
  {32'h40edc20c, 32'hc11b84b1} /* (24, 20, 16) {real, imag} */,
  {32'h4101374a, 32'hc0406880} /* (24, 20, 15) {real, imag} */,
  {32'hc1798f57, 32'h410e90b8} /* (24, 20, 14) {real, imag} */,
  {32'h417c1b13, 32'h405e9780} /* (24, 20, 13) {real, imag} */,
  {32'hc063b189, 32'h4114f922} /* (24, 20, 12) {real, imag} */,
  {32'hc16031f6, 32'h41a9996b} /* (24, 20, 11) {real, imag} */,
  {32'h413f6296, 32'h419c8c09} /* (24, 20, 10) {real, imag} */,
  {32'hc151ea42, 32'h40af584c} /* (24, 20, 9) {real, imag} */,
  {32'h41e45c8a, 32'h411ad8bc} /* (24, 20, 8) {real, imag} */,
  {32'hbe9a3f80, 32'h4125b840} /* (24, 20, 7) {real, imag} */,
  {32'hc1d7f7e4, 32'hc19e31f4} /* (24, 20, 6) {real, imag} */,
  {32'h40c50e02, 32'h41e9018c} /* (24, 20, 5) {real, imag} */,
  {32'hc02f7040, 32'h4271c85c} /* (24, 20, 4) {real, imag} */,
  {32'hc233bc92, 32'hc1c22a4b} /* (24, 20, 3) {real, imag} */,
  {32'hbcb99200, 32'h423970a7} /* (24, 20, 2) {real, imag} */,
  {32'hc14843c0, 32'hc21a4967} /* (24, 20, 1) {real, imag} */,
  {32'hc099af14, 32'hc1b00fc2} /* (24, 20, 0) {real, imag} */,
  {32'hc162e619, 32'hc2010d49} /* (24, 19, 31) {real, imag} */,
  {32'h3fda86c4, 32'h41ba8134} /* (24, 19, 30) {real, imag} */,
  {32'hc1b079cb, 32'hc1442bad} /* (24, 19, 29) {real, imag} */,
  {32'hc086df60, 32'h422a4926} /* (24, 19, 28) {real, imag} */,
  {32'h4113554c, 32'hc20b3c7b} /* (24, 19, 27) {real, imag} */,
  {32'h4151b8f8, 32'hc1c5a717} /* (24, 19, 26) {real, imag} */,
  {32'h40a6aa29, 32'h4133ffc6} /* (24, 19, 25) {real, imag} */,
  {32'h41f7882c, 32'h41117be8} /* (24, 19, 24) {real, imag} */,
  {32'h41c8e5ff, 32'hc0b14246} /* (24, 19, 23) {real, imag} */,
  {32'h41275956, 32'h40532b12} /* (24, 19, 22) {real, imag} */,
  {32'hc1d9fd8b, 32'h41a1f9cc} /* (24, 19, 21) {real, imag} */,
  {32'h41453827, 32'h3f14c420} /* (24, 19, 20) {real, imag} */,
  {32'h3f418990, 32'h3fa5bcfc} /* (24, 19, 19) {real, imag} */,
  {32'h3eba3eb0, 32'h41027b3e} /* (24, 19, 18) {real, imag} */,
  {32'h4002edef, 32'h40f45a78} /* (24, 19, 17) {real, imag} */,
  {32'hc11f0618, 32'hc0b59704} /* (24, 19, 16) {real, imag} */,
  {32'h41040869, 32'hbfc64790} /* (24, 19, 15) {real, imag} */,
  {32'h4155e340, 32'h400605c0} /* (24, 19, 14) {real, imag} */,
  {32'hc0aa939e, 32'hc14cdc7a} /* (24, 19, 13) {real, imag} */,
  {32'h40e83df6, 32'h41273106} /* (24, 19, 12) {real, imag} */,
  {32'h40d5362c, 32'h419f7e34} /* (24, 19, 11) {real, imag} */,
  {32'hc093f70c, 32'h4169bcb0} /* (24, 19, 10) {real, imag} */,
  {32'hc1b03ff9, 32'hc1e5d0cc} /* (24, 19, 9) {real, imag} */,
  {32'hc1b19cb6, 32'hc07bed86} /* (24, 19, 8) {real, imag} */,
  {32'hc11edd2a, 32'hc1d0e1c7} /* (24, 19, 7) {real, imag} */,
  {32'h3e6c3e00, 32'hc1839141} /* (24, 19, 6) {real, imag} */,
  {32'h4180902c, 32'hbfca81e0} /* (24, 19, 5) {real, imag} */,
  {32'h41af21ab, 32'hc1854a5f} /* (24, 19, 4) {real, imag} */,
  {32'h41d59035, 32'hc1c557cc} /* (24, 19, 3) {real, imag} */,
  {32'hc12e494e, 32'h421750f6} /* (24, 19, 2) {real, imag} */,
  {32'hc1d83a5a, 32'hc215055d} /* (24, 19, 1) {real, imag} */,
  {32'h3fbc0a20, 32'h42224e86} /* (24, 19, 0) {real, imag} */,
  {32'h41f3128d, 32'hc1c4ee75} /* (24, 18, 31) {real, imag} */,
  {32'hc0feb759, 32'h3fe07268} /* (24, 18, 30) {real, imag} */,
  {32'hc061955d, 32'hc10a0f84} /* (24, 18, 29) {real, imag} */,
  {32'h41d2c031, 32'hc1477fea} /* (24, 18, 28) {real, imag} */,
  {32'hbfc27310, 32'hc1093ae4} /* (24, 18, 27) {real, imag} */,
  {32'hc07b7e04, 32'h41f99b42} /* (24, 18, 26) {real, imag} */,
  {32'h4145a374, 32'h41748a1c} /* (24, 18, 25) {real, imag} */,
  {32'hc1846240, 32'h41d054fd} /* (24, 18, 24) {real, imag} */,
  {32'hc0da3414, 32'h41a0f259} /* (24, 18, 23) {real, imag} */,
  {32'h40f0aa2a, 32'hc0f071e7} /* (24, 18, 22) {real, imag} */,
  {32'h3f29b718, 32'hc17d5fdc} /* (24, 18, 21) {real, imag} */,
  {32'h3fd9541c, 32'hc0909f24} /* (24, 18, 20) {real, imag} */,
  {32'h404eb26c, 32'h3fd9fbe0} /* (24, 18, 19) {real, imag} */,
  {32'h409b80fb, 32'hc111e92b} /* (24, 18, 18) {real, imag} */,
  {32'hc097c7f4, 32'h40bc556a} /* (24, 18, 17) {real, imag} */,
  {32'hc093f579, 32'h41286e2a} /* (24, 18, 16) {real, imag} */,
  {32'hc0f4bfa0, 32'hc114eca1} /* (24, 18, 15) {real, imag} */,
  {32'h40ca09c1, 32'h416421bf} /* (24, 18, 14) {real, imag} */,
  {32'hbf0d9378, 32'h4039bdc0} /* (24, 18, 13) {real, imag} */,
  {32'hc110e09c, 32'hc1478326} /* (24, 18, 12) {real, imag} */,
  {32'h40d39037, 32'hc12adca0} /* (24, 18, 11) {real, imag} */,
  {32'hc17821d3, 32'h411023d2} /* (24, 18, 10) {real, imag} */,
  {32'h41839055, 32'hc0d8446b} /* (24, 18, 9) {real, imag} */,
  {32'h40d73c75, 32'hc134c7d2} /* (24, 18, 8) {real, imag} */,
  {32'h415a5e08, 32'hc1d6e2b2} /* (24, 18, 7) {real, imag} */,
  {32'hc1dd6808, 32'hc173ff7c} /* (24, 18, 6) {real, imag} */,
  {32'h41f76f53, 32'h40dddf1f} /* (24, 18, 5) {real, imag} */,
  {32'hc1496cc2, 32'h424d0d5c} /* (24, 18, 4) {real, imag} */,
  {32'hc0c58366, 32'h4210eb5c} /* (24, 18, 3) {real, imag} */,
  {32'hc1b99da9, 32'hc18ecf38} /* (24, 18, 2) {real, imag} */,
  {32'h3fa79be0, 32'hc1b37e89} /* (24, 18, 1) {real, imag} */,
  {32'h41a308de, 32'hc1582664} /* (24, 18, 0) {real, imag} */,
  {32'hc055f7c7, 32'hc1146eaa} /* (24, 17, 31) {real, imag} */,
  {32'h405a7f66, 32'hc1f1b20d} /* (24, 17, 30) {real, imag} */,
  {32'hc0d4d636, 32'h41e17f58} /* (24, 17, 29) {real, imag} */,
  {32'hc15c6804, 32'hc1cd6c62} /* (24, 17, 28) {real, imag} */,
  {32'hc18dee47, 32'hc0ced654} /* (24, 17, 27) {real, imag} */,
  {32'h414d84d6, 32'hc1459d94} /* (24, 17, 26) {real, imag} */,
  {32'hc043f600, 32'h404bf93c} /* (24, 17, 25) {real, imag} */,
  {32'hc13daf6a, 32'hc0518c86} /* (24, 17, 24) {real, imag} */,
  {32'hc08b396f, 32'h40b28ff5} /* (24, 17, 23) {real, imag} */,
  {32'hc0038f1e, 32'h40a0a550} /* (24, 17, 22) {real, imag} */,
  {32'h3fed3bee, 32'hbfdff588} /* (24, 17, 21) {real, imag} */,
  {32'hc152f9d7, 32'h416eb843} /* (24, 17, 20) {real, imag} */,
  {32'h401c4169, 32'hc0597c12} /* (24, 17, 19) {real, imag} */,
  {32'hbf2820bc, 32'h407db138} /* (24, 17, 18) {real, imag} */,
  {32'hbfae6070, 32'hc09ad7e7} /* (24, 17, 17) {real, imag} */,
  {32'hc06a3228, 32'hbfaf57d0} /* (24, 17, 16) {real, imag} */,
  {32'hc08f3ed3, 32'hbf8fd7bc} /* (24, 17, 15) {real, imag} */,
  {32'hbfa16456, 32'hc01cb6b8} /* (24, 17, 14) {real, imag} */,
  {32'hc052448f, 32'hbf4a04d8} /* (24, 17, 13) {real, imag} */,
  {32'h400cf738, 32'hbf61a720} /* (24, 17, 12) {real, imag} */,
  {32'hc00495f7, 32'h4086c153} /* (24, 17, 11) {real, imag} */,
  {32'hc1711fc4, 32'h41243a27} /* (24, 17, 10) {real, imag} */,
  {32'h3fcc31c8, 32'h4171da6c} /* (24, 17, 9) {real, imag} */,
  {32'h40a855cc, 32'h4119cc5e} /* (24, 17, 8) {real, imag} */,
  {32'hc178eece, 32'h41a87026} /* (24, 17, 7) {real, imag} */,
  {32'hbf4d7d18, 32'hc14637ec} /* (24, 17, 6) {real, imag} */,
  {32'hc18d2795, 32'h41453d6e} /* (24, 17, 5) {real, imag} */,
  {32'h4132d9bc, 32'hc1727728} /* (24, 17, 4) {real, imag} */,
  {32'h4177e15f, 32'h3f903068} /* (24, 17, 3) {real, imag} */,
  {32'h41021c84, 32'hc20d57fe} /* (24, 17, 2) {real, imag} */,
  {32'h3f3394b4, 32'h420b3d4c} /* (24, 17, 1) {real, imag} */,
  {32'h413d8438, 32'h421842f6} /* (24, 17, 0) {real, imag} */,
  {32'hc12471c8, 32'hc097550a} /* (24, 16, 31) {real, imag} */,
  {32'h416bba63, 32'h413c9bcc} /* (24, 16, 30) {real, imag} */,
  {32'h42040668, 32'hc1e3452f} /* (24, 16, 29) {real, imag} */,
  {32'h41aeeac7, 32'hc1dacb80} /* (24, 16, 28) {real, imag} */,
  {32'h41db203a, 32'hc11a41b8} /* (24, 16, 27) {real, imag} */,
  {32'hc1af3914, 32'hc1d53874} /* (24, 16, 26) {real, imag} */,
  {32'h410c0b27, 32'hc0c6f97a} /* (24, 16, 25) {real, imag} */,
  {32'h41cf76bf, 32'hc119627b} /* (24, 16, 24) {real, imag} */,
  {32'hbf7beafc, 32'h40d818df} /* (24, 16, 23) {real, imag} */,
  {32'hc180e715, 32'hc01ababc} /* (24, 16, 22) {real, imag} */,
  {32'hc08c106d, 32'h3fae2a78} /* (24, 16, 21) {real, imag} */,
  {32'h3fb3b61d, 32'hc0bb79d0} /* (24, 16, 20) {real, imag} */,
  {32'h408c2f40, 32'hc05c08de} /* (24, 16, 19) {real, imag} */,
  {32'hbfa38060, 32'h3ffaf5ae} /* (24, 16, 18) {real, imag} */,
  {32'hbe845280, 32'h4015b99a} /* (24, 16, 17) {real, imag} */,
  {32'h4101c616, 32'hc02bde80} /* (24, 16, 16) {real, imag} */,
  {32'h4092b1d8, 32'hbf871208} /* (24, 16, 15) {real, imag} */,
  {32'hc167915e, 32'hc022ce3b} /* (24, 16, 14) {real, imag} */,
  {32'hbf2c37a0, 32'hc0ad6d3d} /* (24, 16, 13) {real, imag} */,
  {32'h40256686, 32'h41204904} /* (24, 16, 12) {real, imag} */,
  {32'hc09e7bbd, 32'hc1339f6a} /* (24, 16, 11) {real, imag} */,
  {32'hc0928cdc, 32'hbfd6aff8} /* (24, 16, 10) {real, imag} */,
  {32'hc0805cac, 32'hc0e39349} /* (24, 16, 9) {real, imag} */,
  {32'hc0fbbdc4, 32'h4175f4bd} /* (24, 16, 8) {real, imag} */,
  {32'h41502127, 32'hc1bb28d6} /* (24, 16, 7) {real, imag} */,
  {32'h41be5b06, 32'h3ff556f8} /* (24, 16, 6) {real, imag} */,
  {32'hc197168c, 32'h41b92494} /* (24, 16, 5) {real, imag} */,
  {32'hc1c2d565, 32'hbfcd6960} /* (24, 16, 4) {real, imag} */,
  {32'hc1dd8a4d, 32'hc17330c2} /* (24, 16, 3) {real, imag} */,
  {32'hc19cc32a, 32'h4153f86c} /* (24, 16, 2) {real, imag} */,
  {32'hc240205c, 32'h410d2635} /* (24, 16, 1) {real, imag} */,
  {32'hc10c24ea, 32'h4259fe04} /* (24, 16, 0) {real, imag} */,
  {32'h4227ae1a, 32'hc0766cd3} /* (24, 15, 31) {real, imag} */,
  {32'hc1521a5c, 32'h403ea4c5} /* (24, 15, 30) {real, imag} */,
  {32'hc2135806, 32'h417abb4e} /* (24, 15, 29) {real, imag} */,
  {32'hc0f11418, 32'hc1fbcd3f} /* (24, 15, 28) {real, imag} */,
  {32'h41d3601e, 32'h41382dbd} /* (24, 15, 27) {real, imag} */,
  {32'h40fdc078, 32'hc160e626} /* (24, 15, 26) {real, imag} */,
  {32'h419dc977, 32'h40960203} /* (24, 15, 25) {real, imag} */,
  {32'hc1121a02, 32'h41b7f29a} /* (24, 15, 24) {real, imag} */,
  {32'h3f11b3bc, 32'h3ecc9d60} /* (24, 15, 23) {real, imag} */,
  {32'h40f09aae, 32'hc18e7886} /* (24, 15, 22) {real, imag} */,
  {32'hc12be95e, 32'hc0d7b906} /* (24, 15, 21) {real, imag} */,
  {32'h4091c62c, 32'h40ac3b25} /* (24, 15, 20) {real, imag} */,
  {32'h40c1d0f1, 32'h40468f68} /* (24, 15, 19) {real, imag} */,
  {32'h3e4cafc0, 32'hbe8ea698} /* (24, 15, 18) {real, imag} */,
  {32'hbdf05c80, 32'h4116f39c} /* (24, 15, 17) {real, imag} */,
  {32'hc006e07c, 32'h4039e62b} /* (24, 15, 16) {real, imag} */,
  {32'h3d8ba980, 32'h3fd9bca4} /* (24, 15, 15) {real, imag} */,
  {32'h4062714c, 32'hc0665429} /* (24, 15, 14) {real, imag} */,
  {32'h3fd0c0d4, 32'h410ad0b0} /* (24, 15, 13) {real, imag} */,
  {32'hc15c9e12, 32'h40532c5a} /* (24, 15, 12) {real, imag} */,
  {32'hbf892684, 32'hc0dda896} /* (24, 15, 11) {real, imag} */,
  {32'h40b78f7e, 32'hc16b5c2c} /* (24, 15, 10) {real, imag} */,
  {32'hc09c779a, 32'hc1de68a6} /* (24, 15, 9) {real, imag} */,
  {32'h4037c1f2, 32'hc1e69b56} /* (24, 15, 8) {real, imag} */,
  {32'hc06976d8, 32'h412fd4f0} /* (24, 15, 7) {real, imag} */,
  {32'hc181dd1f, 32'hc21a823a} /* (24, 15, 6) {real, imag} */,
  {32'h40a64806, 32'hc20f1c74} /* (24, 15, 5) {real, imag} */,
  {32'h3fd6f9a8, 32'hc01c5178} /* (24, 15, 4) {real, imag} */,
  {32'h40cce620, 32'h41002af0} /* (24, 15, 3) {real, imag} */,
  {32'hc0ad943c, 32'h40e179cc} /* (24, 15, 2) {real, imag} */,
  {32'hc175211d, 32'h41356120} /* (24, 15, 1) {real, imag} */,
  {32'hc0657634, 32'hc11ba82d} /* (24, 15, 0) {real, imag} */,
  {32'hc155ace6, 32'h4219da77} /* (24, 14, 31) {real, imag} */,
  {32'h41066044, 32'h40672d20} /* (24, 14, 30) {real, imag} */,
  {32'hc1809946, 32'h40cc47b8} /* (24, 14, 29) {real, imag} */,
  {32'h4209d4fc, 32'hc1130592} /* (24, 14, 28) {real, imag} */,
  {32'hc14bcd0e, 32'h412bcad3} /* (24, 14, 27) {real, imag} */,
  {32'hc21c6187, 32'h3f932e86} /* (24, 14, 26) {real, imag} */,
  {32'h4105939e, 32'hc18bae30} /* (24, 14, 25) {real, imag} */,
  {32'h41d43ebe, 32'hc080adc2} /* (24, 14, 24) {real, imag} */,
  {32'h42109259, 32'hc08a7f08} /* (24, 14, 23) {real, imag} */,
  {32'hbe7e7840, 32'h3edd3eb0} /* (24, 14, 22) {real, imag} */,
  {32'hc0f1fc50, 32'h419d0d40} /* (24, 14, 21) {real, imag} */,
  {32'h40f3b505, 32'hc0e9a5c3} /* (24, 14, 20) {real, imag} */,
  {32'hc03b07fa, 32'hc080ad46} /* (24, 14, 19) {real, imag} */,
  {32'hc006208a, 32'h4115df52} /* (24, 14, 18) {real, imag} */,
  {32'hc0cddbbd, 32'hc059533c} /* (24, 14, 17) {real, imag} */,
  {32'h40f6b66c, 32'h4090de70} /* (24, 14, 16) {real, imag} */,
  {32'h3f4d9d38, 32'hbf345e70} /* (24, 14, 15) {real, imag} */,
  {32'h4012d046, 32'h3e8469d0} /* (24, 14, 14) {real, imag} */,
  {32'hbf8375b5, 32'h40aaffca} /* (24, 14, 13) {real, imag} */,
  {32'h4151514e, 32'h4193030b} /* (24, 14, 12) {real, imag} */,
  {32'h40e064fe, 32'h4174dbdf} /* (24, 14, 11) {real, imag} */,
  {32'hc14bc3a5, 32'hc11526b4} /* (24, 14, 10) {real, imag} */,
  {32'h415bb775, 32'h41c1f97e} /* (24, 14, 9) {real, imag} */,
  {32'h41853804, 32'h3e3d0a40} /* (24, 14, 8) {real, imag} */,
  {32'h41543c22, 32'hc1e477b4} /* (24, 14, 7) {real, imag} */,
  {32'hc18cf122, 32'h40157761} /* (24, 14, 6) {real, imag} */,
  {32'hc103763a, 32'h412202d5} /* (24, 14, 5) {real, imag} */,
  {32'h404cd6a8, 32'hc17fab6e} /* (24, 14, 4) {real, imag} */,
  {32'hc118e334, 32'hc258facb} /* (24, 14, 3) {real, imag} */,
  {32'h4156a0a4, 32'hc1bb9cbc} /* (24, 14, 2) {real, imag} */,
  {32'hc18ab8bb, 32'hc11969e5} /* (24, 14, 1) {real, imag} */,
  {32'hc2125064, 32'h410c4b1a} /* (24, 14, 0) {real, imag} */,
  {32'hc1b0b318, 32'h4218c34e} /* (24, 13, 31) {real, imag} */,
  {32'h41d4654a, 32'h4200040a} /* (24, 13, 30) {real, imag} */,
  {32'h40c437cf, 32'h41691a96} /* (24, 13, 29) {real, imag} */,
  {32'h40a8c084, 32'hc1cde036} /* (24, 13, 28) {real, imag} */,
  {32'h42201622, 32'h40b54548} /* (24, 13, 27) {real, imag} */,
  {32'h4158028e, 32'h421252e4} /* (24, 13, 26) {real, imag} */,
  {32'hbff180a0, 32'hc18ac6b1} /* (24, 13, 25) {real, imag} */,
  {32'hc114fa66, 32'h41d5229a} /* (24, 13, 24) {real, imag} */,
  {32'hc0d2f225, 32'hc0d41cda} /* (24, 13, 23) {real, imag} */,
  {32'hc167c457, 32'hc0ab68b0} /* (24, 13, 22) {real, imag} */,
  {32'hc1520a26, 32'h3f9f7a91} /* (24, 13, 21) {real, imag} */,
  {32'hc188e292, 32'h3ff40620} /* (24, 13, 20) {real, imag} */,
  {32'h41a060f3, 32'hc0f5c8ab} /* (24, 13, 19) {real, imag} */,
  {32'hc0c4855c, 32'h410209e4} /* (24, 13, 18) {real, imag} */,
  {32'h3de2d620, 32'hc0582426} /* (24, 13, 17) {real, imag} */,
  {32'h40591664, 32'hc07ff618} /* (24, 13, 16) {real, imag} */,
  {32'hbe488810, 32'hc0da474b} /* (24, 13, 15) {real, imag} */,
  {32'hc0b14610, 32'hc08e1473} /* (24, 13, 14) {real, imag} */,
  {32'h40a28c19, 32'h416b8db4} /* (24, 13, 13) {real, imag} */,
  {32'h419008b4, 32'hc1a4a892} /* (24, 13, 12) {real, imag} */,
  {32'h41dea603, 32'hc019658c} /* (24, 13, 11) {real, imag} */,
  {32'h3ffe3de8, 32'hc0f42928} /* (24, 13, 10) {real, imag} */,
  {32'h40666696, 32'h41107077} /* (24, 13, 9) {real, imag} */,
  {32'h41cde4cf, 32'h40a8d67e} /* (24, 13, 8) {real, imag} */,
  {32'h41a9f47e, 32'hc1972a23} /* (24, 13, 7) {real, imag} */,
  {32'hc1bdbb63, 32'hc0958edc} /* (24, 13, 6) {real, imag} */,
  {32'hc098218c, 32'hc085d2b6} /* (24, 13, 5) {real, imag} */,
  {32'h41f63d7b, 32'hc15ed370} /* (24, 13, 4) {real, imag} */,
  {32'h41486506, 32'h41b5cce9} /* (24, 13, 3) {real, imag} */,
  {32'h41a920d2, 32'hbe692980} /* (24, 13, 2) {real, imag} */,
  {32'hc1c2280a, 32'hc24bb5ee} /* (24, 13, 1) {real, imag} */,
  {32'h42006c71, 32'h413709a5} /* (24, 13, 0) {real, imag} */,
  {32'h3f4960a0, 32'h4058d224} /* (24, 12, 31) {real, imag} */,
  {32'hc1be29e2, 32'hc1387901} /* (24, 12, 30) {real, imag} */,
  {32'hc1bf319a, 32'hc2242599} /* (24, 12, 29) {real, imag} */,
  {32'hc1ac41f7, 32'h422c708e} /* (24, 12, 28) {real, imag} */,
  {32'hc1b0b77d, 32'h41e9cc4a} /* (24, 12, 27) {real, imag} */,
  {32'hc1837b13, 32'hc2172fb7} /* (24, 12, 26) {real, imag} */,
  {32'h413c603a, 32'h41769f2c} /* (24, 12, 25) {real, imag} */,
  {32'h414b4310, 32'h421f4efc} /* (24, 12, 24) {real, imag} */,
  {32'hbefb2850, 32'h419de2cf} /* (24, 12, 23) {real, imag} */,
  {32'hc0e243cc, 32'h40bf5bc2} /* (24, 12, 22) {real, imag} */,
  {32'hc164e9fa, 32'h418951ff} /* (24, 12, 21) {real, imag} */,
  {32'h40d8c79c, 32'h3fae9db4} /* (24, 12, 20) {real, imag} */,
  {32'h40474bd1, 32'h41191b84} /* (24, 12, 19) {real, imag} */,
  {32'h4052bd2c, 32'h41625476} /* (24, 12, 18) {real, imag} */,
  {32'h3f01ad10, 32'hc14e77ab} /* (24, 12, 17) {real, imag} */,
  {32'hc132bd45, 32'hc0b4c28c} /* (24, 12, 16) {real, imag} */,
  {32'hc0eef50a, 32'hc10fc261} /* (24, 12, 15) {real, imag} */,
  {32'h418bb020, 32'h40493570} /* (24, 12, 14) {real, imag} */,
  {32'h4112e3d2, 32'h40e0ea48} /* (24, 12, 13) {real, imag} */,
  {32'hc08c4234, 32'hc0d53659} /* (24, 12, 12) {real, imag} */,
  {32'hc03eb0e0, 32'hc133ae44} /* (24, 12, 11) {real, imag} */,
  {32'h42083634, 32'hc18975fe} /* (24, 12, 10) {real, imag} */,
  {32'h412273ce, 32'h41364586} /* (24, 12, 9) {real, imag} */,
  {32'h412a10c8, 32'h4116bf3d} /* (24, 12, 8) {real, imag} */,
  {32'hc0b64dcc, 32'hc22ce671} /* (24, 12, 7) {real, imag} */,
  {32'h418b7903, 32'h41152907} /* (24, 12, 6) {real, imag} */,
  {32'hc1b3ea0f, 32'hc16ccb7d} /* (24, 12, 5) {real, imag} */,
  {32'hc1d5dc1f, 32'h41bcfd71} /* (24, 12, 4) {real, imag} */,
  {32'hc0c5a17c, 32'hc1d9b3da} /* (24, 12, 3) {real, imag} */,
  {32'h419a92d6, 32'h420d3ba6} /* (24, 12, 2) {real, imag} */,
  {32'h420b80dc, 32'h41cd948e} /* (24, 12, 1) {real, imag} */,
  {32'hc1a8f996, 32'h42436a96} /* (24, 12, 0) {real, imag} */,
  {32'h41ed1330, 32'h4222bb48} /* (24, 11, 31) {real, imag} */,
  {32'h402d1858, 32'hc1d2bbac} /* (24, 11, 30) {real, imag} */,
  {32'hc1aa676e, 32'h40a6fdf8} /* (24, 11, 29) {real, imag} */,
  {32'h3f99f5c0, 32'h42204229} /* (24, 11, 28) {real, imag} */,
  {32'h4152ea33, 32'h3f2f23a0} /* (24, 11, 27) {real, imag} */,
  {32'hc07f6e90, 32'hc22e7e7a} /* (24, 11, 26) {real, imag} */,
  {32'hc1f11dc1, 32'h4113ea3a} /* (24, 11, 25) {real, imag} */,
  {32'hc18b5a4e, 32'h418f6977} /* (24, 11, 24) {real, imag} */,
  {32'h41cb2f3f, 32'h40701562} /* (24, 11, 23) {real, imag} */,
  {32'h41266e6e, 32'h3f4d1cd0} /* (24, 11, 22) {real, imag} */,
  {32'h419a990e, 32'hc2196bb4} /* (24, 11, 21) {real, imag} */,
  {32'hc10f83e0, 32'hbf5fd1a0} /* (24, 11, 20) {real, imag} */,
  {32'hc0dac656, 32'h4149b3d8} /* (24, 11, 19) {real, imag} */,
  {32'h3fed5cb4, 32'hbf9ca684} /* (24, 11, 18) {real, imag} */,
  {32'hbffe0f5a, 32'hc0065b56} /* (24, 11, 17) {real, imag} */,
  {32'h411ece31, 32'h3f978a0c} /* (24, 11, 16) {real, imag} */,
  {32'h40a2ac56, 32'hc0a3ece5} /* (24, 11, 15) {real, imag} */,
  {32'h3fb95fac, 32'hbd486180} /* (24, 11, 14) {real, imag} */,
  {32'h40984b32, 32'hc00784d2} /* (24, 11, 13) {real, imag} */,
  {32'hc1c6ef2a, 32'hc138c5be} /* (24, 11, 12) {real, imag} */,
  {32'h416568ad, 32'hbfa15d90} /* (24, 11, 11) {real, imag} */,
  {32'hc11c9f9e, 32'h41a0c3b8} /* (24, 11, 10) {real, imag} */,
  {32'h3f903270, 32'hc1280104} /* (24, 11, 9) {real, imag} */,
  {32'hc004b076, 32'h412d715a} /* (24, 11, 8) {real, imag} */,
  {32'h41a8a873, 32'h41c6728f} /* (24, 11, 7) {real, imag} */,
  {32'hc0a8008e, 32'hc0f4bc14} /* (24, 11, 6) {real, imag} */,
  {32'hc1bcd526, 32'h419ebfd7} /* (24, 11, 5) {real, imag} */,
  {32'hc28b21b5, 32'hc2a060de} /* (24, 11, 4) {real, imag} */,
  {32'h4238ccc1, 32'hc0342c2d} /* (24, 11, 3) {real, imag} */,
  {32'h41f5ce3b, 32'hc1a12178} /* (24, 11, 2) {real, imag} */,
  {32'hc2037628, 32'h41e6960d} /* (24, 11, 1) {real, imag} */,
  {32'hc11c1fd3, 32'h402aedfa} /* (24, 11, 0) {real, imag} */,
  {32'h42cfaf59, 32'hc1d4407a} /* (24, 10, 31) {real, imag} */,
  {32'hc20fd719, 32'h42b3bd62} /* (24, 10, 30) {real, imag} */,
  {32'hc249460c, 32'h41a5b249} /* (24, 10, 29) {real, imag} */,
  {32'h424c77a8, 32'hc234e15e} /* (24, 10, 28) {real, imag} */,
  {32'hc1ab7e32, 32'h42a41555} /* (24, 10, 27) {real, imag} */,
  {32'hc210bda5, 32'h417ebd69} /* (24, 10, 26) {real, imag} */,
  {32'hc1ec384e, 32'hc18ee337} /* (24, 10, 25) {real, imag} */,
  {32'h41ea5818, 32'hc033ae88} /* (24, 10, 24) {real, imag} */,
  {32'h4188950e, 32'hc1a24b6f} /* (24, 10, 23) {real, imag} */,
  {32'hc1ee17fc, 32'h42261f18} /* (24, 10, 22) {real, imag} */,
  {32'h41aa6279, 32'h3f0523f8} /* (24, 10, 21) {real, imag} */,
  {32'h41bdc3c0, 32'hbf3c6ce0} /* (24, 10, 20) {real, imag} */,
  {32'hbfe6dfe4, 32'hbf8d6c98} /* (24, 10, 19) {real, imag} */,
  {32'hc0e0690e, 32'h4094e560} /* (24, 10, 18) {real, imag} */,
  {32'h3f7971e0, 32'h414144ac} /* (24, 10, 17) {real, imag} */,
  {32'hc14588a8, 32'h4197b7e2} /* (24, 10, 16) {real, imag} */,
  {32'h40e36254, 32'h419af9e2} /* (24, 10, 15) {real, imag} */,
  {32'hc165cb9f, 32'hc012f760} /* (24, 10, 14) {real, imag} */,
  {32'h40ccde8f, 32'hc0f392aa} /* (24, 10, 13) {real, imag} */,
  {32'h415e4724, 32'hc1d15763} /* (24, 10, 12) {real, imag} */,
  {32'hbec03ec0, 32'h40d0970f} /* (24, 10, 11) {real, imag} */,
  {32'h4179c5d9, 32'hc1a5dd0a} /* (24, 10, 10) {real, imag} */,
  {32'h4163e38b, 32'h41247942} /* (24, 10, 9) {real, imag} */,
  {32'hc1838028, 32'h40c17210} /* (24, 10, 8) {real, imag} */,
  {32'hc18ac4ea, 32'h41dcd86d} /* (24, 10, 7) {real, imag} */,
  {32'hc18f587e, 32'h41787f55} /* (24, 10, 6) {real, imag} */,
  {32'hc07232b0, 32'hc2c63d7b} /* (24, 10, 5) {real, imag} */,
  {32'h4286430c, 32'hc1695e22} /* (24, 10, 4) {real, imag} */,
  {32'h4205d47c, 32'hc0ca6260} /* (24, 10, 3) {real, imag} */,
  {32'h4226af7d, 32'hc0868868} /* (24, 10, 2) {real, imag} */,
  {32'hc1ca73a4, 32'h4192aabe} /* (24, 10, 1) {real, imag} */,
  {32'hc23beeae, 32'hc28c4c20} /* (24, 10, 0) {real, imag} */,
  {32'h3f222060, 32'h42101cd8} /* (24, 9, 31) {real, imag} */,
  {32'h41c992d3, 32'hc2bf68a9} /* (24, 9, 30) {real, imag} */,
  {32'hc1c86444, 32'hc23709a9} /* (24, 9, 29) {real, imag} */,
  {32'h40b726f0, 32'hc23df9be} /* (24, 9, 28) {real, imag} */,
  {32'hc22ebd77, 32'h422dbb4a} /* (24, 9, 27) {real, imag} */,
  {32'hc185bbdc, 32'h4187ef8f} /* (24, 9, 26) {real, imag} */,
  {32'h4122a364, 32'hc22d8d92} /* (24, 9, 25) {real, imag} */,
  {32'hc1e2ada5, 32'h41de6900} /* (24, 9, 24) {real, imag} */,
  {32'hc1fa917d, 32'h4175593a} /* (24, 9, 23) {real, imag} */,
  {32'hc0a8846e, 32'hc16816c4} /* (24, 9, 22) {real, imag} */,
  {32'h410f1e36, 32'hc1e9493a} /* (24, 9, 21) {real, imag} */,
  {32'h41d258ea, 32'hc194fd62} /* (24, 9, 20) {real, imag} */,
  {32'hc1a3a69a, 32'hc12e8856} /* (24, 9, 19) {real, imag} */,
  {32'hc1b3fee7, 32'h42598a9e} /* (24, 9, 18) {real, imag} */,
  {32'hc0274878, 32'hc1ed0923} /* (24, 9, 17) {real, imag} */,
  {32'hc1598689, 32'hc025c5f0} /* (24, 9, 16) {real, imag} */,
  {32'hbf9c9bc0, 32'hc130cc5a} /* (24, 9, 15) {real, imag} */,
  {32'h41a9cbed, 32'hc095d290} /* (24, 9, 14) {real, imag} */,
  {32'hc24db555, 32'hc13f1ce2} /* (24, 9, 13) {real, imag} */,
  {32'h4104fda4, 32'hc1b9d412} /* (24, 9, 12) {real, imag} */,
  {32'h40a621cc, 32'hc213137b} /* (24, 9, 11) {real, imag} */,
  {32'hc1560787, 32'hc17c38b8} /* (24, 9, 10) {real, imag} */,
  {32'h40d812cc, 32'h41ebe703} /* (24, 9, 9) {real, imag} */,
  {32'hc1118e6e, 32'h410758a8} /* (24, 9, 8) {real, imag} */,
  {32'h4200288a, 32'h41b995c4} /* (24, 9, 7) {real, imag} */,
  {32'h417ba8a9, 32'h4141b4ca} /* (24, 9, 6) {real, imag} */,
  {32'h4082bc10, 32'h414f56b8} /* (24, 9, 5) {real, imag} */,
  {32'h422d04e8, 32'hc088b4e0} /* (24, 9, 4) {real, imag} */,
  {32'h414221b8, 32'hc24f2795} /* (24, 9, 3) {real, imag} */,
  {32'hc1bf2361, 32'h429d4d69} /* (24, 9, 2) {real, imag} */,
  {32'hc1d1aa47, 32'h42ad844a} /* (24, 9, 1) {real, imag} */,
  {32'hc0c281ba, 32'hc2c1d8a8} /* (24, 9, 0) {real, imag} */,
  {32'h400a16f8, 32'h43294d79} /* (24, 8, 31) {real, imag} */,
  {32'hc2cd8a2c, 32'hc3160bc6} /* (24, 8, 30) {real, imag} */,
  {32'h428e993a, 32'h42aa9d28} /* (24, 8, 29) {real, imag} */,
  {32'h42306d2f, 32'hc2e936fc} /* (24, 8, 28) {real, imag} */,
  {32'hc2137dcd, 32'hc2108789} /* (24, 8, 27) {real, imag} */,
  {32'h42208904, 32'hc0804de0} /* (24, 8, 26) {real, imag} */,
  {32'hc27647ce, 32'h4141c431} /* (24, 8, 25) {real, imag} */,
  {32'hc2a97062, 32'h4002b59a} /* (24, 8, 24) {real, imag} */,
  {32'h414d02e0, 32'hbeb118c0} /* (24, 8, 23) {real, imag} */,
  {32'hc1a0ab22, 32'h4163e99a} /* (24, 8, 22) {real, imag} */,
  {32'hc09d5c21, 32'h40999134} /* (24, 8, 21) {real, imag} */,
  {32'h41998c81, 32'hc119e8c6} /* (24, 8, 20) {real, imag} */,
  {32'hc12b8438, 32'hc17a1912} /* (24, 8, 19) {real, imag} */,
  {32'h411ccf5e, 32'h405d1eb0} /* (24, 8, 18) {real, imag} */,
  {32'h412d183d, 32'h3ffa7cac} /* (24, 8, 17) {real, imag} */,
  {32'hbea2f600, 32'hc17dc31a} /* (24, 8, 16) {real, imag} */,
  {32'hc074543c, 32'h4179a50a} /* (24, 8, 15) {real, imag} */,
  {32'h4121bf6a, 32'h41923866} /* (24, 8, 14) {real, imag} */,
  {32'h41b0672c, 32'h41edd74f} /* (24, 8, 13) {real, imag} */,
  {32'h40f292b0, 32'h4144f32e} /* (24, 8, 12) {real, imag} */,
  {32'h40f7f897, 32'h41a6466f} /* (24, 8, 11) {real, imag} */,
  {32'h41685a74, 32'hc17dc720} /* (24, 8, 10) {real, imag} */,
  {32'hc1af7f08, 32'h423ce6aa} /* (24, 8, 9) {real, imag} */,
  {32'h420485c0, 32'h41365f68} /* (24, 8, 8) {real, imag} */,
  {32'hc2a99553, 32'h40bc7d36} /* (24, 8, 7) {real, imag} */,
  {32'h40b5cbe0, 32'hc2270d86} /* (24, 8, 6) {real, imag} */,
  {32'h40a6abd0, 32'hc29e2490} /* (24, 8, 5) {real, imag} */,
  {32'h42332f05, 32'hc194ec20} /* (24, 8, 4) {real, imag} */,
  {32'hc2c04b40, 32'h4220f050} /* (24, 8, 3) {real, imag} */,
  {32'hc115f1c4, 32'hc28e6564} /* (24, 8, 2) {real, imag} */,
  {32'h427e1188, 32'h431da0a1} /* (24, 8, 1) {real, imag} */,
  {32'h42883bf6, 32'h41eb84f1} /* (24, 8, 0) {real, imag} */,
  {32'hc23ee345, 32'h41b28804} /* (24, 7, 31) {real, imag} */,
  {32'h4240a155, 32'h42eb0cb7} /* (24, 7, 30) {real, imag} */,
  {32'h427059b8, 32'hc210220e} /* (24, 7, 29) {real, imag} */,
  {32'hc25d543c, 32'hc28d45ec} /* (24, 7, 28) {real, imag} */,
  {32'hc1310274, 32'hc2b22213} /* (24, 7, 27) {real, imag} */,
  {32'h41a5284a, 32'hc2a9ccd5} /* (24, 7, 26) {real, imag} */,
  {32'h4276d96e, 32'h4281fd65} /* (24, 7, 25) {real, imag} */,
  {32'h4288010c, 32'h41d1bdb9} /* (24, 7, 24) {real, imag} */,
  {32'h423df1ad, 32'hc1b3fb34} /* (24, 7, 23) {real, imag} */,
  {32'hc12b41c6, 32'hc24fc0fe} /* (24, 7, 22) {real, imag} */,
  {32'hc18348cc, 32'hc1193f92} /* (24, 7, 21) {real, imag} */,
  {32'hc1dd5002, 32'h423daee9} /* (24, 7, 20) {real, imag} */,
  {32'h4139572c, 32'hc08ce9cc} /* (24, 7, 19) {real, imag} */,
  {32'hc0b04fbe, 32'h40948e74} /* (24, 7, 18) {real, imag} */,
  {32'hc13dc232, 32'h410df0ec} /* (24, 7, 17) {real, imag} */,
  {32'h3f25fe20, 32'hc1ade55e} /* (24, 7, 16) {real, imag} */,
  {32'hc0af7d4c, 32'hc0a8a514} /* (24, 7, 15) {real, imag} */,
  {32'h41c291e4, 32'hc187569d} /* (24, 7, 14) {real, imag} */,
  {32'hc14e3644, 32'hc1cd2879} /* (24, 7, 13) {real, imag} */,
  {32'hc0c3d700, 32'h4141887c} /* (24, 7, 12) {real, imag} */,
  {32'h41094f69, 32'hc1a55771} /* (24, 7, 11) {real, imag} */,
  {32'h4236f2d8, 32'hc1eb0e28} /* (24, 7, 10) {real, imag} */,
  {32'hc1b9559e, 32'h40ce2238} /* (24, 7, 9) {real, imag} */,
  {32'hc19870c5, 32'h420c10b2} /* (24, 7, 8) {real, imag} */,
  {32'h41cc1a9f, 32'hc0a1a4ec} /* (24, 7, 7) {real, imag} */,
  {32'hc2bfd08a, 32'hc2315e5e} /* (24, 7, 6) {real, imag} */,
  {32'h4226bce5, 32'h42b7cdd3} /* (24, 7, 5) {real, imag} */,
  {32'h419472d9, 32'h41a5b038} /* (24, 7, 4) {real, imag} */,
  {32'hc2cc5516, 32'h40fa43f4} /* (24, 7, 3) {real, imag} */,
  {32'hc1bb003a, 32'hc1b08edc} /* (24, 7, 2) {real, imag} */,
  {32'h42257077, 32'h400aba38} /* (24, 7, 1) {real, imag} */,
  {32'hc23a2ade, 32'hc2f3bed4} /* (24, 7, 0) {real, imag} */,
  {32'hc2d156a4, 32'hc2112804} /* (24, 6, 31) {real, imag} */,
  {32'hbf395c60, 32'h4307ecc8} /* (24, 6, 30) {real, imag} */,
  {32'h4258d32d, 32'hc1e69999} /* (24, 6, 29) {real, imag} */,
  {32'h42c03230, 32'h42fcbf34} /* (24, 6, 28) {real, imag} */,
  {32'h42dcaf76, 32'h41efcde0} /* (24, 6, 27) {real, imag} */,
  {32'hc298110f, 32'h41ab0742} /* (24, 6, 26) {real, imag} */,
  {32'hc19bc11b, 32'h428e4dbc} /* (24, 6, 25) {real, imag} */,
  {32'hc25e7616, 32'hc212b9a2} /* (24, 6, 24) {real, imag} */,
  {32'hc1f4b3d2, 32'hc1ae4b26} /* (24, 6, 23) {real, imag} */,
  {32'hc16b3910, 32'hc22efd18} /* (24, 6, 22) {real, imag} */,
  {32'h413cb83a, 32'hc16efa4e} /* (24, 6, 21) {real, imag} */,
  {32'hc0e30984, 32'hc1dda56c} /* (24, 6, 20) {real, imag} */,
  {32'h424f5a3c, 32'h421b3040} /* (24, 6, 19) {real, imag} */,
  {32'hc1f1ebbf, 32'hc18f998a} /* (24, 6, 18) {real, imag} */,
  {32'h412920b2, 32'h409a6a14} /* (24, 6, 17) {real, imag} */,
  {32'hc01612b0, 32'hc08feb3a} /* (24, 6, 16) {real, imag} */,
  {32'h4114d6de, 32'hc1ad7bb1} /* (24, 6, 15) {real, imag} */,
  {32'h415cbe66, 32'hbf0671c0} /* (24, 6, 14) {real, imag} */,
  {32'h41ba1fd8, 32'hc00dbe58} /* (24, 6, 13) {real, imag} */,
  {32'h416c6d22, 32'h4185cf78} /* (24, 6, 12) {real, imag} */,
  {32'hc2854355, 32'h41a35809} /* (24, 6, 11) {real, imag} */,
  {32'hc22a8e2e, 32'h425a4c80} /* (24, 6, 10) {real, imag} */,
  {32'h40901166, 32'h416e5ca4} /* (24, 6, 9) {real, imag} */,
  {32'hc193adcd, 32'h40264f18} /* (24, 6, 8) {real, imag} */,
  {32'hbf8a6940, 32'h42b27ad0} /* (24, 6, 7) {real, imag} */,
  {32'h41ce4340, 32'hc21eb387} /* (24, 6, 6) {real, imag} */,
  {32'h41008ce0, 32'hc2d456ac} /* (24, 6, 5) {real, imag} */,
  {32'h427a2418, 32'h41904e32} /* (24, 6, 4) {real, imag} */,
  {32'h429b7592, 32'hc1e017f9} /* (24, 6, 3) {real, imag} */,
  {32'h41b6bed3, 32'h413cc094} /* (24, 6, 2) {real, imag} */,
  {32'h419d8c26, 32'hc2a99431} /* (24, 6, 1) {real, imag} */,
  {32'hc28caeb0, 32'hc10d48e9} /* (24, 6, 0) {real, imag} */,
  {32'h42696196, 32'h42b69e98} /* (24, 5, 31) {real, imag} */,
  {32'hc253b0ca, 32'hc2b26ddc} /* (24, 5, 30) {real, imag} */,
  {32'h41b1f7b2, 32'h41257f1e} /* (24, 5, 29) {real, imag} */,
  {32'h424a3536, 32'hc13c6a9c} /* (24, 5, 28) {real, imag} */,
  {32'hc289fa0e, 32'h420570e3} /* (24, 5, 27) {real, imag} */,
  {32'hc1ebacbe, 32'h41ed3dd4} /* (24, 5, 26) {real, imag} */,
  {32'h4270b5e3, 32'h41c3fcb9} /* (24, 5, 25) {real, imag} */,
  {32'hc1dbb600, 32'hc1c00a36} /* (24, 5, 24) {real, imag} */,
  {32'h41462c66, 32'hbff5edc8} /* (24, 5, 23) {real, imag} */,
  {32'hbf799470, 32'hc0839e7d} /* (24, 5, 22) {real, imag} */,
  {32'h41234873, 32'h423372ee} /* (24, 5, 21) {real, imag} */,
  {32'hc1b5a9f7, 32'h41056e10} /* (24, 5, 20) {real, imag} */,
  {32'hc0994038, 32'hc11b4984} /* (24, 5, 19) {real, imag} */,
  {32'hc196f8a3, 32'h41a6af55} /* (24, 5, 18) {real, imag} */,
  {32'hc0f541e9, 32'hc125b7aa} /* (24, 5, 17) {real, imag} */,
  {32'h41c4836e, 32'h4256b5fa} /* (24, 5, 16) {real, imag} */,
  {32'hc0ee0ca9, 32'hc1d3779f} /* (24, 5, 15) {real, imag} */,
  {32'hc18bd2cd, 32'h41a1b507} /* (24, 5, 14) {real, imag} */,
  {32'hc2824a00, 32'hc0b24264} /* (24, 5, 13) {real, imag} */,
  {32'h423ef5b4, 32'h40ba8e10} /* (24, 5, 12) {real, imag} */,
  {32'h41aabec6, 32'hc0f5ee30} /* (24, 5, 11) {real, imag} */,
  {32'hc13893c7, 32'hbe8f9d70} /* (24, 5, 10) {real, imag} */,
  {32'h41688116, 32'h41875d24} /* (24, 5, 9) {real, imag} */,
  {32'h42779066, 32'hc2332e6d} /* (24, 5, 8) {real, imag} */,
  {32'hc28d5ad3, 32'h420d851b} /* (24, 5, 7) {real, imag} */,
  {32'h41bba392, 32'h409e5190} /* (24, 5, 6) {real, imag} */,
  {32'h4202e055, 32'h404cb670} /* (24, 5, 5) {real, imag} */,
  {32'h42a24525, 32'hc2c69a94} /* (24, 5, 4) {real, imag} */,
  {32'h40a15212, 32'h3f0b3a00} /* (24, 5, 3) {real, imag} */,
  {32'h41fdf38c, 32'hc2bc3380} /* (24, 5, 2) {real, imag} */,
  {32'hc2498d3e, 32'h41d4dc76} /* (24, 5, 1) {real, imag} */,
  {32'h41c1ab32, 32'h42929991} /* (24, 5, 0) {real, imag} */,
  {32'hc02d9b10, 32'hc2951729} /* (24, 4, 31) {real, imag} */,
  {32'h4210eeda, 32'h432f9cbb} /* (24, 4, 30) {real, imag} */,
  {32'h421519bb, 32'hc3111a58} /* (24, 4, 29) {real, imag} */,
  {32'hc256a5fc, 32'hbffd90e0} /* (24, 4, 28) {real, imag} */,
  {32'h411584d4, 32'hc3363cf8} /* (24, 4, 27) {real, imag} */,
  {32'h41dea777, 32'h41704430} /* (24, 4, 26) {real, imag} */,
  {32'h42066ff2, 32'h402e94a0} /* (24, 4, 25) {real, imag} */,
  {32'h4262a30c, 32'hc1c807d1} /* (24, 4, 24) {real, imag} */,
  {32'h41c761d4, 32'hc1a15eb3} /* (24, 4, 23) {real, imag} */,
  {32'h40f40074, 32'hc225a804} /* (24, 4, 22) {real, imag} */,
  {32'hc167e050, 32'hc128e38c} /* (24, 4, 21) {real, imag} */,
  {32'hc11afb55, 32'h41a907ba} /* (24, 4, 20) {real, imag} */,
  {32'h412eae60, 32'hc1690f32} /* (24, 4, 19) {real, imag} */,
  {32'hc1b25dfe, 32'h41ea47a3} /* (24, 4, 18) {real, imag} */,
  {32'hc11cceb9, 32'h41bfdd70} /* (24, 4, 17) {real, imag} */,
  {32'h408da71c, 32'hc14063fe} /* (24, 4, 16) {real, imag} */,
  {32'h40c32c1e, 32'h40edfd20} /* (24, 4, 15) {real, imag} */,
  {32'hc03b7150, 32'h42124f36} /* (24, 4, 14) {real, imag} */,
  {32'h419366c8, 32'hc1c886af} /* (24, 4, 13) {real, imag} */,
  {32'hc1865bf2, 32'hc19d2302} /* (24, 4, 12) {real, imag} */,
  {32'hc2818b92, 32'h4299272c} /* (24, 4, 11) {real, imag} */,
  {32'h42002b24, 32'h41326cbc} /* (24, 4, 10) {real, imag} */,
  {32'hc2d8f711, 32'h422af942} /* (24, 4, 9) {real, imag} */,
  {32'h4106a922, 32'h409ab754} /* (24, 4, 8) {real, imag} */,
  {32'h419c011b, 32'hc3037fdc} /* (24, 4, 7) {real, imag} */,
  {32'h41633fe6, 32'hc164e30c} /* (24, 4, 6) {real, imag} */,
  {32'h420e3495, 32'h40fd4e50} /* (24, 4, 5) {real, imag} */,
  {32'h42bc900c, 32'hc2ed015a} /* (24, 4, 4) {real, imag} */,
  {32'hc201e9d5, 32'hc30e46a4} /* (24, 4, 3) {real, imag} */,
  {32'hc2821360, 32'h4330f383} /* (24, 4, 2) {real, imag} */,
  {32'hc25a57ad, 32'hc35baea4} /* (24, 4, 1) {real, imag} */,
  {32'hc08d35bc, 32'hc1d48d9d} /* (24, 4, 0) {real, imag} */,
  {32'h43101fff, 32'hc19d0d6e} /* (24, 3, 31) {real, imag} */,
  {32'hc270f4b2, 32'hc25a3bc7} /* (24, 3, 30) {real, imag} */,
  {32'hc2a6f816, 32'h4346c4e4} /* (24, 3, 29) {real, imag} */,
  {32'h4222bfff, 32'hc33c18ba} /* (24, 3, 28) {real, imag} */,
  {32'h428f55ea, 32'hbf8d1cc0} /* (24, 3, 27) {real, imag} */,
  {32'h42cfefac, 32'hc29edd44} /* (24, 3, 26) {real, imag} */,
  {32'hc237adf0, 32'h41b0985a} /* (24, 3, 25) {real, imag} */,
  {32'hc22e1450, 32'h429ef616} /* (24, 3, 24) {real, imag} */,
  {32'h41a8b8af, 32'h4264496f} /* (24, 3, 23) {real, imag} */,
  {32'h428ead30, 32'h3fb42ab0} /* (24, 3, 22) {real, imag} */,
  {32'hc25662df, 32'hc221d8d2} /* (24, 3, 21) {real, imag} */,
  {32'hc0587b88, 32'h420419a8} /* (24, 3, 20) {real, imag} */,
  {32'hc1ccacfe, 32'hc134c978} /* (24, 3, 19) {real, imag} */,
  {32'hc22e575b, 32'hc1fac21f} /* (24, 3, 18) {real, imag} */,
  {32'h40028320, 32'h4199cea6} /* (24, 3, 17) {real, imag} */,
  {32'hc17474e4, 32'h41292e52} /* (24, 3, 16) {real, imag} */,
  {32'h419988c8, 32'h4225bc15} /* (24, 3, 15) {real, imag} */,
  {32'h40866b40, 32'hc22c8c76} /* (24, 3, 14) {real, imag} */,
  {32'hc22a7df5, 32'h41b44c9c} /* (24, 3, 13) {real, imag} */,
  {32'hc20fbf48, 32'h4258cd68} /* (24, 3, 12) {real, imag} */,
  {32'hc12a61bc, 32'hc18136d8} /* (24, 3, 11) {real, imag} */,
  {32'h41089b06, 32'hc153c0aa} /* (24, 3, 10) {real, imag} */,
  {32'h412a857a, 32'hbfcd9e60} /* (24, 3, 9) {real, imag} */,
  {32'h422ccf68, 32'h404b73b0} /* (24, 3, 8) {real, imag} */,
  {32'hc24dac52, 32'hc0d447ec} /* (24, 3, 7) {real, imag} */,
  {32'hc252a4b3, 32'h40da3848} /* (24, 3, 6) {real, imag} */,
  {32'h416e6564, 32'hc28fe0a8} /* (24, 3, 5) {real, imag} */,
  {32'h42820570, 32'h4281e138} /* (24, 3, 4) {real, imag} */,
  {32'h42d877de, 32'h42cfc0d9} /* (24, 3, 3) {real, imag} */,
  {32'hc2845e41, 32'h423364bd} /* (24, 3, 2) {real, imag} */,
  {32'hc213488d, 32'hc290a558} /* (24, 3, 1) {real, imag} */,
  {32'h42859d64, 32'hc1f37221} /* (24, 3, 0) {real, imag} */,
  {32'h43888517, 32'h43f40070} /* (24, 2, 31) {real, imag} */,
  {32'hc3823403, 32'hc2b4e650} /* (24, 2, 30) {real, imag} */,
  {32'h42a78328, 32'h42447754} /* (24, 2, 29) {real, imag} */,
  {32'h4242f6b3, 32'hc24e8296} /* (24, 2, 28) {real, imag} */,
  {32'hc32ebb96, 32'hc1b85d9c} /* (24, 2, 27) {real, imag} */,
  {32'h429e9253, 32'h42fb174a} /* (24, 2, 26) {real, imag} */,
  {32'h4196f4a6, 32'h40c22e98} /* (24, 2, 25) {real, imag} */,
  {32'hc330fd1d, 32'hc1d6d748} /* (24, 2, 24) {real, imag} */,
  {32'hc1ec55f2, 32'h41ca82e2} /* (24, 2, 23) {real, imag} */,
  {32'h41c748f4, 32'hc1d59df4} /* (24, 2, 22) {real, imag} */,
  {32'h419a71ab, 32'h4197ed82} /* (24, 2, 21) {real, imag} */,
  {32'hc15ecdf4, 32'hc292de8f} /* (24, 2, 20) {real, imag} */,
  {32'h42285d06, 32'hc1eb853d} /* (24, 2, 19) {real, imag} */,
  {32'h415567b9, 32'hc1d92990} /* (24, 2, 18) {real, imag} */,
  {32'hc0c6966a, 32'hbea6ac00} /* (24, 2, 17) {real, imag} */,
  {32'h416d13b8, 32'h419d37b0} /* (24, 2, 16) {real, imag} */,
  {32'hc12d5d0b, 32'hc0996d00} /* (24, 2, 15) {real, imag} */,
  {32'hc09dee32, 32'h40b49f00} /* (24, 2, 14) {real, imag} */,
  {32'h411d15f0, 32'h3f545020} /* (24, 2, 13) {real, imag} */,
  {32'h423c9939, 32'h423fba0e} /* (24, 2, 12) {real, imag} */,
  {32'h41a6ac77, 32'hc10de65c} /* (24, 2, 11) {real, imag} */,
  {32'hc20dee6e, 32'hc13163d8} /* (24, 2, 10) {real, imag} */,
  {32'hbff704a0, 32'h41bc109e} /* (24, 2, 9) {real, imag} */,
  {32'hc1473310, 32'hc2d1d10c} /* (24, 2, 8) {real, imag} */,
  {32'hc2148475, 32'hc28d4496} /* (24, 2, 7) {real, imag} */,
  {32'h40ad6e90, 32'hc180a6e8} /* (24, 2, 6) {real, imag} */,
  {32'h42832198, 32'hc3416ac8} /* (24, 2, 5) {real, imag} */,
  {32'h42e97562, 32'h4250f012} /* (24, 2, 4) {real, imag} */,
  {32'h42da04f0, 32'hc217dad0} /* (24, 2, 3) {real, imag} */,
  {32'hc39d2d91, 32'hc3c3518d} /* (24, 2, 2) {real, imag} */,
  {32'h439f9f65, 32'h42071f3c} /* (24, 2, 1) {real, imag} */,
  {32'h42fc42b5, 32'h438b19a9} /* (24, 2, 0) {real, imag} */,
  {32'hc38e6341, 32'hc395bcc4} /* (24, 1, 31) {real, imag} */,
  {32'h43561667, 32'h43199e66} /* (24, 1, 30) {real, imag} */,
  {32'h41c0f28c, 32'h41b6a390} /* (24, 1, 29) {real, imag} */,
  {32'h421c0c9e, 32'hc2d48b9a} /* (24, 1, 28) {real, imag} */,
  {32'h428b0384, 32'h4334eb20} /* (24, 1, 27) {real, imag} */,
  {32'hc2799760, 32'h41907299} /* (24, 1, 26) {real, imag} */,
  {32'h42a00209, 32'hc1634290} /* (24, 1, 25) {real, imag} */,
  {32'h4171a1f0, 32'hc2291984} /* (24, 1, 24) {real, imag} */,
  {32'h418970c4, 32'h42c5c97a} /* (24, 1, 23) {real, imag} */,
  {32'hc0ab4ac0, 32'hbffae2b0} /* (24, 1, 22) {real, imag} */,
  {32'hc1a9a0aa, 32'hc1e02abc} /* (24, 1, 21) {real, imag} */,
  {32'h40a61de0, 32'hc1b50eba} /* (24, 1, 20) {real, imag} */,
  {32'h401b2dc0, 32'h41ddd03c} /* (24, 1, 19) {real, imag} */,
  {32'h417eb598, 32'hc27f34c6} /* (24, 1, 18) {real, imag} */,
  {32'hc164f534, 32'h41790630} /* (24, 1, 17) {real, imag} */,
  {32'hc1a37950, 32'hc1a82598} /* (24, 1, 16) {real, imag} */,
  {32'h42a08d6a, 32'h3fbe8880} /* (24, 1, 15) {real, imag} */,
  {32'hc17f9a18, 32'hbe932500} /* (24, 1, 14) {real, imag} */,
  {32'hc05ec7d8, 32'hc1b7875c} /* (24, 1, 13) {real, imag} */,
  {32'hc232ed58, 32'h40893718} /* (24, 1, 12) {real, imag} */,
  {32'h40aa6c6a, 32'h4297607b} /* (24, 1, 11) {real, imag} */,
  {32'h42935904, 32'hc2664dac} /* (24, 1, 10) {real, imag} */,
  {32'hc29b417e, 32'h41c8d134} /* (24, 1, 9) {real, imag} */,
  {32'hc2a5d7a2, 32'h42df64de} /* (24, 1, 8) {real, imag} */,
  {32'hc20b76f8, 32'hc0cbae50} /* (24, 1, 7) {real, imag} */,
  {32'hc145625e, 32'hc0bfcad4} /* (24, 1, 6) {real, imag} */,
  {32'h41c960d2, 32'h43029a02} /* (24, 1, 5) {real, imag} */,
  {32'h42bb06e9, 32'h4293abfe} /* (24, 1, 4) {real, imag} */,
  {32'hc0c97524, 32'hc19c4a48} /* (24, 1, 3) {real, imag} */,
  {32'hc25d46f4, 32'h43f7ccaf} /* (24, 1, 2) {real, imag} */,
  {32'hc31ab97c, 32'hc43b155e} /* (24, 1, 1) {real, imag} */,
  {32'hc36ef09c, 32'hc3e34c68} /* (24, 1, 0) {real, imag} */,
  {32'hc3ad76f9, 32'hc2bc727c} /* (24, 0, 31) {real, imag} */,
  {32'h42ffd7b3, 32'hc2e10236} /* (24, 0, 30) {real, imag} */,
  {32'h41dd4729, 32'h4301f19b} /* (24, 0, 29) {real, imag} */,
  {32'hc12ac770, 32'hc204d0bc} /* (24, 0, 28) {real, imag} */,
  {32'h42e7a1b4, 32'h4279e395} /* (24, 0, 27) {real, imag} */,
  {32'h42c0a852, 32'hc2ab7964} /* (24, 0, 26) {real, imag} */,
  {32'hc300ec64, 32'hc2a60441} /* (24, 0, 25) {real, imag} */,
  {32'h42805624, 32'h42692947} /* (24, 0, 24) {real, imag} */,
  {32'h42046de9, 32'hc20e0e5a} /* (24, 0, 23) {real, imag} */,
  {32'hc2af28b2, 32'h42a4222b} /* (24, 0, 22) {real, imag} */,
  {32'h420e4210, 32'h418675f4} /* (24, 0, 21) {real, imag} */,
  {32'hc19833f9, 32'hc1aa6b21} /* (24, 0, 20) {real, imag} */,
  {32'hc1a367e8, 32'h41f07bd0} /* (24, 0, 19) {real, imag} */,
  {32'h42690062, 32'hc26b3b2c} /* (24, 0, 18) {real, imag} */,
  {32'hc21c4bb3, 32'hc22b2398} /* (24, 0, 17) {real, imag} */,
  {32'hc192a52e, 32'hc0b2b500} /* (24, 0, 16) {real, imag} */,
  {32'hc189014a, 32'hc0966ee0} /* (24, 0, 15) {real, imag} */,
  {32'hc122d0aa, 32'hc11f6fa0} /* (24, 0, 14) {real, imag} */,
  {32'h4022a6d0, 32'h42026a1c} /* (24, 0, 13) {real, imag} */,
  {32'hc1cbcb25, 32'h4004cb18} /* (24, 0, 12) {real, imag} */,
  {32'hc25b28a4, 32'h41677b30} /* (24, 0, 11) {real, imag} */,
  {32'hc0f76560, 32'h414dca08} /* (24, 0, 10) {real, imag} */,
  {32'h41f249ce, 32'hc1d5c42c} /* (24, 0, 9) {real, imag} */,
  {32'hc2d38d82, 32'h418c085a} /* (24, 0, 8) {real, imag} */,
  {32'h42ac9d5c, 32'hc288cbd3} /* (24, 0, 7) {real, imag} */,
  {32'hc228f964, 32'h4294570a} /* (24, 0, 6) {real, imag} */,
  {32'hc0da42e0, 32'h42ec1c16} /* (24, 0, 5) {real, imag} */,
  {32'hc2e37810, 32'h419266bb} /* (24, 0, 4) {real, imag} */,
  {32'h428e316a, 32'hc250b6a8} /* (24, 0, 3) {real, imag} */,
  {32'hc20dcb76, 32'h42b126bc} /* (24, 0, 2) {real, imag} */,
  {32'hc33563f6, 32'hc3ca9af3} /* (24, 0, 1) {real, imag} */,
  {32'hc30d681c, 32'hc348900f} /* (24, 0, 0) {real, imag} */,
  {32'hc320011c, 32'h41373994} /* (23, 31, 31) {real, imag} */,
  {32'h43163f25, 32'h42da83ad} /* (23, 31, 30) {real, imag} */,
  {32'h413a2da7, 32'h437a1e60} /* (23, 31, 29) {real, imag} */,
  {32'hc18780aa, 32'hc283491d} /* (23, 31, 28) {real, imag} */,
  {32'h42905610, 32'h41550ecf} /* (23, 31, 27) {real, imag} */,
  {32'h422ef702, 32'h42248e45} /* (23, 31, 26) {real, imag} */,
  {32'h4242625e, 32'hc224cee5} /* (23, 31, 25) {real, imag} */,
  {32'hc28bba62, 32'hc30a86db} /* (23, 31, 24) {real, imag} */,
  {32'h41e99e8c, 32'hc27af767} /* (23, 31, 23) {real, imag} */,
  {32'hc1f64088, 32'hc20ccac3} /* (23, 31, 22) {real, imag} */,
  {32'hc1cfbe1f, 32'h3f0a3150} /* (23, 31, 21) {real, imag} */,
  {32'hc1995747, 32'hc0eabd6a} /* (23, 31, 20) {real, imag} */,
  {32'hc0ad1ffa, 32'h422957ff} /* (23, 31, 19) {real, imag} */,
  {32'hc1a8b187, 32'h41245951} /* (23, 31, 18) {real, imag} */,
  {32'h411af648, 32'h3fa21940} /* (23, 31, 17) {real, imag} */,
  {32'h41276b58, 32'h41e47d4e} /* (23, 31, 16) {real, imag} */,
  {32'h4111e368, 32'hc19ba860} /* (23, 31, 15) {real, imag} */,
  {32'h4148d9ee, 32'h414d3087} /* (23, 31, 14) {real, imag} */,
  {32'h41b9b3d2, 32'h41ce8b96} /* (23, 31, 13) {real, imag} */,
  {32'hc248cfa4, 32'h4133029d} /* (23, 31, 12) {real, imag} */,
  {32'h41f7736d, 32'hc115ecaf} /* (23, 31, 11) {real, imag} */,
  {32'h423bd214, 32'h41d1b4ae} /* (23, 31, 10) {real, imag} */,
  {32'h40d71210, 32'h420002ef} /* (23, 31, 9) {real, imag} */,
  {32'h418899ba, 32'h41ecde22} /* (23, 31, 8) {real, imag} */,
  {32'hc285fbd1, 32'hc1efd61e} /* (23, 31, 7) {real, imag} */,
  {32'hc2d3856b, 32'hc2988cf0} /* (23, 31, 6) {real, imag} */,
  {32'h41c3cf5a, 32'hc229bd0d} /* (23, 31, 5) {real, imag} */,
  {32'hbf08e4f0, 32'hc21c6b19} /* (23, 31, 4) {real, imag} */,
  {32'h40a75892, 32'h40114c20} /* (23, 31, 3) {real, imag} */,
  {32'h428ed470, 32'h42c1af67} /* (23, 31, 2) {real, imag} */,
  {32'hc202ab66, 32'hc2f0fe5e} /* (23, 31, 1) {real, imag} */,
  {32'hc312e8dc, 32'h42857d40} /* (23, 31, 0) {real, imag} */,
  {32'h42cf3a32, 32'h42e4516d} /* (23, 30, 31) {real, imag} */,
  {32'h4245b65c, 32'hc351139b} /* (23, 30, 30) {real, imag} */,
  {32'hc277e92b, 32'hc2d2c36f} /* (23, 30, 29) {real, imag} */,
  {32'h4250b09a, 32'h42f63806} /* (23, 30, 28) {real, imag} */,
  {32'hc28fd89e, 32'h41f0a673} /* (23, 30, 27) {real, imag} */,
  {32'h42837eb1, 32'hc2017d63} /* (23, 30, 26) {real, imag} */,
  {32'h42d03b41, 32'h41b634c7} /* (23, 30, 25) {real, imag} */,
  {32'hc29cdff0, 32'hc1cce74c} /* (23, 30, 24) {real, imag} */,
  {32'hbfd72d00, 32'h41ff1524} /* (23, 30, 23) {real, imag} */,
  {32'h424d0138, 32'hc2391f38} /* (23, 30, 22) {real, imag} */,
  {32'hc252b3a4, 32'h41cb7fa3} /* (23, 30, 21) {real, imag} */,
  {32'h41915308, 32'h410cacba} /* (23, 30, 20) {real, imag} */,
  {32'hc1427b88, 32'h4181aefa} /* (23, 30, 19) {real, imag} */,
  {32'h4207a9f0, 32'h40e76ed4} /* (23, 30, 18) {real, imag} */,
  {32'h421d294a, 32'hc2013f3c} /* (23, 30, 17) {real, imag} */,
  {32'h419e51ac, 32'h40837470} /* (23, 30, 16) {real, imag} */,
  {32'hc0f4da68, 32'hc08a36b4} /* (23, 30, 15) {real, imag} */,
  {32'h4187c3f5, 32'hc2123996} /* (23, 30, 14) {real, imag} */,
  {32'hc2398898, 32'hc1a3ed42} /* (23, 30, 13) {real, imag} */,
  {32'h40a9e132, 32'h42147660} /* (23, 30, 12) {real, imag} */,
  {32'h41ecb7c8, 32'hc16291ca} /* (23, 30, 11) {real, imag} */,
  {32'h42840df2, 32'hc1c8eb4c} /* (23, 30, 10) {real, imag} */,
  {32'hc1a81616, 32'h419b6ce2} /* (23, 30, 9) {real, imag} */,
  {32'hc1e72e50, 32'h417d52d8} /* (23, 30, 8) {real, imag} */,
  {32'h41847c64, 32'hc253d8ac} /* (23, 30, 7) {real, imag} */,
  {32'h4219d92a, 32'hc29d503c} /* (23, 30, 6) {real, imag} */,
  {32'h3ff65e80, 32'hc1ddc11d} /* (23, 30, 5) {real, imag} */,
  {32'hc29a6a1b, 32'h42e4c362} /* (23, 30, 4) {real, imag} */,
  {32'hc3106e63, 32'hbdd41000} /* (23, 30, 3) {real, imag} */,
  {32'hc221ac6e, 32'hc326f769} /* (23, 30, 2) {real, imag} */,
  {32'h4201eff9, 32'h42c2ab37} /* (23, 30, 1) {real, imag} */,
  {32'h41b9cd2e, 32'h42e7fe0b} /* (23, 30, 0) {real, imag} */,
  {32'hc0f4c30e, 32'h421d79d8} /* (23, 29, 31) {real, imag} */,
  {32'hc2b8755d, 32'h4324cae6} /* (23, 29, 30) {real, imag} */,
  {32'h42aeea0c, 32'h41e610f6} /* (23, 29, 29) {real, imag} */,
  {32'hc13427aa, 32'hc2b784da} /* (23, 29, 28) {real, imag} */,
  {32'h4294295e, 32'hc1092591} /* (23, 29, 27) {real, imag} */,
  {32'h42736f54, 32'h42d8a940} /* (23, 29, 26) {real, imag} */,
  {32'hc247a229, 32'hc23a0ff9} /* (23, 29, 25) {real, imag} */,
  {32'h42301fc2, 32'hc13eadc4} /* (23, 29, 24) {real, imag} */,
  {32'hc16886e2, 32'h3f9ce4a0} /* (23, 29, 23) {real, imag} */,
  {32'hc05ba0a0, 32'hc0affb1c} /* (23, 29, 22) {real, imag} */,
  {32'hc142ba74, 32'hc26ff774} /* (23, 29, 21) {real, imag} */,
  {32'h41e71132, 32'h41984cf4} /* (23, 29, 20) {real, imag} */,
  {32'h41043e4f, 32'h4291026a} /* (23, 29, 19) {real, imag} */,
  {32'hc2145e06, 32'hc14ebcbc} /* (23, 29, 18) {real, imag} */,
  {32'hc115925a, 32'hc1e2d80a} /* (23, 29, 17) {real, imag} */,
  {32'hc0945268, 32'hc130f8ae} /* (23, 29, 16) {real, imag} */,
  {32'h41e61d67, 32'h40ec7df6} /* (23, 29, 15) {real, imag} */,
  {32'hc20108b2, 32'hc00dbbf0} /* (23, 29, 14) {real, imag} */,
  {32'h420c92c4, 32'h403e5fa0} /* (23, 29, 13) {real, imag} */,
  {32'h40174db4, 32'hc19aa43a} /* (23, 29, 12) {real, imag} */,
  {32'h41115f24, 32'h41981598} /* (23, 29, 11) {real, imag} */,
  {32'hc25977b8, 32'hbfcd2790} /* (23, 29, 10) {real, imag} */,
  {32'hc1d9d8df, 32'h42993b7c} /* (23, 29, 9) {real, imag} */,
  {32'hbe220e00, 32'hc1467adc} /* (23, 29, 8) {real, imag} */,
  {32'h422113e7, 32'hc2396f4f} /* (23, 29, 7) {real, imag} */,
  {32'h41d803a4, 32'h4281a2ec} /* (23, 29, 6) {real, imag} */,
  {32'h41ae67b6, 32'hc1d5957c} /* (23, 29, 5) {real, imag} */,
  {32'hc01286a2, 32'hc1d8efc0} /* (23, 29, 4) {real, imag} */,
  {32'h42cd0f2e, 32'hc15bafac} /* (23, 29, 3) {real, imag} */,
  {32'hc1122b38, 32'hc205ae60} /* (23, 29, 2) {real, imag} */,
  {32'hc04cfdc4, 32'hc08dfca0} /* (23, 29, 1) {real, imag} */,
  {32'h42ad374a, 32'h415184b8} /* (23, 29, 0) {real, imag} */,
  {32'hc0a9c914, 32'hc21a78b0} /* (23, 28, 31) {real, imag} */,
  {32'hbfcdf680, 32'hc1c5260c} /* (23, 28, 30) {real, imag} */,
  {32'h42dee63e, 32'hc0b5ecf0} /* (23, 28, 29) {real, imag} */,
  {32'hc1cb5499, 32'hc1e6011d} /* (23, 28, 28) {real, imag} */,
  {32'hc1d27da4, 32'h4195ebce} /* (23, 28, 27) {real, imag} */,
  {32'hc2bf10cc, 32'hc275be8f} /* (23, 28, 26) {real, imag} */,
  {32'h419d9b58, 32'h421441ea} /* (23, 28, 25) {real, imag} */,
  {32'hc1cdab5a, 32'h41c3a06a} /* (23, 28, 24) {real, imag} */,
  {32'h42051adb, 32'hc24e8b9f} /* (23, 28, 23) {real, imag} */,
  {32'h41be7929, 32'h421351d3} /* (23, 28, 22) {real, imag} */,
  {32'h42834e75, 32'h41b86890} /* (23, 28, 21) {real, imag} */,
  {32'hc0d7a2e7, 32'h41d181a2} /* (23, 28, 20) {real, imag} */,
  {32'h4197d4b8, 32'hc1a1aac0} /* (23, 28, 19) {real, imag} */,
  {32'h411c3204, 32'h41454858} /* (23, 28, 18) {real, imag} */,
  {32'hc1f1089d, 32'hc163f134} /* (23, 28, 17) {real, imag} */,
  {32'hc0e879e0, 32'hc1258d76} /* (23, 28, 16) {real, imag} */,
  {32'hc1a176bb, 32'hc10d8e30} /* (23, 28, 15) {real, imag} */,
  {32'h41726760, 32'hc15e4694} /* (23, 28, 14) {real, imag} */,
  {32'h3f73dac0, 32'hc203eb4a} /* (23, 28, 13) {real, imag} */,
  {32'h410fd1fa, 32'hc2044437} /* (23, 28, 12) {real, imag} */,
  {32'h41339f48, 32'h41df8ebc} /* (23, 28, 11) {real, imag} */,
  {32'hc276778a, 32'h421dc06f} /* (23, 28, 10) {real, imag} */,
  {32'hc2129a89, 32'h41ee60f6} /* (23, 28, 9) {real, imag} */,
  {32'hc2470033, 32'hc20af216} /* (23, 28, 8) {real, imag} */,
  {32'h4306161d, 32'hc1ce4a98} /* (23, 28, 7) {real, imag} */,
  {32'h41a10216, 32'hc2846dd7} /* (23, 28, 6) {real, imag} */,
  {32'hc2c3b185, 32'hc2f75bf0} /* (23, 28, 5) {real, imag} */,
  {32'h4255c03e, 32'h414895be} /* (23, 28, 4) {real, imag} */,
  {32'h418a7f98, 32'hc2eba3de} /* (23, 28, 3) {real, imag} */,
  {32'h42398a27, 32'h424d4b3e} /* (23, 28, 2) {real, imag} */,
  {32'h42503bf2, 32'hc1ed99df} /* (23, 28, 1) {real, imag} */,
  {32'h40a4cf58, 32'hc1636e0a} /* (23, 28, 0) {real, imag} */,
  {32'h423bdf40, 32'h419b5898} /* (23, 27, 31) {real, imag} */,
  {32'h42169584, 32'h427fba59} /* (23, 27, 30) {real, imag} */,
  {32'hc2a78a0b, 32'h4126c250} /* (23, 27, 29) {real, imag} */,
  {32'hc21b24a3, 32'hc27a6496} /* (23, 27, 28) {real, imag} */,
  {32'h4266d73b, 32'h4029ae98} /* (23, 27, 27) {real, imag} */,
  {32'hc2ae36c3, 32'h40b8bb49} /* (23, 27, 26) {real, imag} */,
  {32'h42830a6c, 32'h4089b938} /* (23, 27, 25) {real, imag} */,
  {32'h405c6a10, 32'h4196854a} /* (23, 27, 24) {real, imag} */,
  {32'h424d7989, 32'h421c80ee} /* (23, 27, 23) {real, imag} */,
  {32'hc08f75e4, 32'hc0adce07} /* (23, 27, 22) {real, imag} */,
  {32'hc21aeb73, 32'h42a334f4} /* (23, 27, 21) {real, imag} */,
  {32'h41b380b2, 32'hc1224e6e} /* (23, 27, 20) {real, imag} */,
  {32'h41d9f487, 32'h4167a7b0} /* (23, 27, 19) {real, imag} */,
  {32'hc07337e8, 32'hc1167b5f} /* (23, 27, 18) {real, imag} */,
  {32'h4185222a, 32'h42198684} /* (23, 27, 17) {real, imag} */,
  {32'hc085bc28, 32'h407beac0} /* (23, 27, 16) {real, imag} */,
  {32'h40e1b5d2, 32'h4101d7fa} /* (23, 27, 15) {real, imag} */,
  {32'h41bb0d8d, 32'h404c8aa4} /* (23, 27, 14) {real, imag} */,
  {32'h4272e794, 32'h41e34290} /* (23, 27, 13) {real, imag} */,
  {32'hbebce460, 32'hc1bb6d71} /* (23, 27, 12) {real, imag} */,
  {32'hc1c9e2fe, 32'hc12959d4} /* (23, 27, 11) {real, imag} */,
  {32'h41ef8e53, 32'h400e5bc6} /* (23, 27, 10) {real, imag} */,
  {32'hc1e18506, 32'h4258506e} /* (23, 27, 9) {real, imag} */,
  {32'hc2023793, 32'h42cba612} /* (23, 27, 8) {real, imag} */,
  {32'h404a13c8, 32'hc231d87f} /* (23, 27, 7) {real, imag} */,
  {32'h420d033c, 32'h40a68243} /* (23, 27, 6) {real, imag} */,
  {32'h412266ec, 32'hc25104d8} /* (23, 27, 5) {real, imag} */,
  {32'h42417085, 32'h4215df06} /* (23, 27, 4) {real, imag} */,
  {32'hc2729a6a, 32'h42ac6598} /* (23, 27, 3) {real, imag} */,
  {32'hc2ab153c, 32'hc257cf75} /* (23, 27, 2) {real, imag} */,
  {32'hc0caabe4, 32'h425da380} /* (23, 27, 1) {real, imag} */,
  {32'h42902cf0, 32'h42a102b8} /* (23, 27, 0) {real, imag} */,
  {32'h4299f3f3, 32'h41bcd3fb} /* (23, 26, 31) {real, imag} */,
  {32'h41f89cf7, 32'hc3023edf} /* (23, 26, 30) {real, imag} */,
  {32'h4191052b, 32'hc109f474} /* (23, 26, 29) {real, imag} */,
  {32'hc271d11d, 32'h42914f9b} /* (23, 26, 28) {real, imag} */,
  {32'hc2717628, 32'hc162771e} /* (23, 26, 27) {real, imag} */,
  {32'hc201664c, 32'h4262c454} /* (23, 26, 26) {real, imag} */,
  {32'h420bd38f, 32'h41e85520} /* (23, 26, 25) {real, imag} */,
  {32'h4219ff30, 32'h41a777e0} /* (23, 26, 24) {real, imag} */,
  {32'h41450c60, 32'hc0f27dff} /* (23, 26, 23) {real, imag} */,
  {32'h41b1528e, 32'h4111401e} /* (23, 26, 22) {real, imag} */,
  {32'hc11f9217, 32'h424c80e6} /* (23, 26, 21) {real, imag} */,
  {32'h4240a044, 32'hc03615e8} /* (23, 26, 20) {real, imag} */,
  {32'h4191722b, 32'h413d35de} /* (23, 26, 19) {real, imag} */,
  {32'hc17bae0a, 32'hc1b66208} /* (23, 26, 18) {real, imag} */,
  {32'h40c99e11, 32'hc126cce2} /* (23, 26, 17) {real, imag} */,
  {32'h4194424a, 32'h411258a6} /* (23, 26, 16) {real, imag} */,
  {32'hbf529608, 32'h408ef32c} /* (23, 26, 15) {real, imag} */,
  {32'hc1ac4b8f, 32'hc1ab630c} /* (23, 26, 14) {real, imag} */,
  {32'h407f0252, 32'hc0da27bd} /* (23, 26, 13) {real, imag} */,
  {32'hc19fa803, 32'hc210df88} /* (23, 26, 12) {real, imag} */,
  {32'h40b14d3e, 32'h40e0d034} /* (23, 26, 11) {real, imag} */,
  {32'h40ba1b82, 32'h3f7413e0} /* (23, 26, 10) {real, imag} */,
  {32'h4281b360, 32'hc193e66a} /* (23, 26, 9) {real, imag} */,
  {32'h41b2a974, 32'hc1709e50} /* (23, 26, 8) {real, imag} */,
  {32'h4160ac1c, 32'h4114debc} /* (23, 26, 7) {real, imag} */,
  {32'h422021e2, 32'hc2e0b106} /* (23, 26, 6) {real, imag} */,
  {32'h41188700, 32'h418ee2f1} /* (23, 26, 5) {real, imag} */,
  {32'hc211b607, 32'h420b5df0} /* (23, 26, 4) {real, imag} */,
  {32'h40fa7a71, 32'hc1300344} /* (23, 26, 3) {real, imag} */,
  {32'h428e0ca5, 32'hc256e73c} /* (23, 26, 2) {real, imag} */,
  {32'h429a72ed, 32'h41afb3ab} /* (23, 26, 1) {real, imag} */,
  {32'hc2cab314, 32'hc12172e2} /* (23, 26, 0) {real, imag} */,
  {32'hc1b04b9a, 32'h42d833c3} /* (23, 25, 31) {real, imag} */,
  {32'hc2a4e0a9, 32'h41975822} /* (23, 25, 30) {real, imag} */,
  {32'hc1d0761c, 32'hc264a232} /* (23, 25, 29) {real, imag} */,
  {32'hc27e99ba, 32'hc0fd8550} /* (23, 25, 28) {real, imag} */,
  {32'h40ac87b7, 32'h41f50fe6} /* (23, 25, 27) {real, imag} */,
  {32'h418a022a, 32'hc1687698} /* (23, 25, 26) {real, imag} */,
  {32'hc2098c96, 32'hc1979488} /* (23, 25, 25) {real, imag} */,
  {32'hc1faeddc, 32'h42a66952} /* (23, 25, 24) {real, imag} */,
  {32'hc1ffa4e2, 32'hc17d2ad4} /* (23, 25, 23) {real, imag} */,
  {32'hc1cd4f82, 32'h41a03e9c} /* (23, 25, 22) {real, imag} */,
  {32'h4170e8b9, 32'hc106131b} /* (23, 25, 21) {real, imag} */,
  {32'hc1be0d3a, 32'hc1eeb5fd} /* (23, 25, 20) {real, imag} */,
  {32'hc0c33b96, 32'hc24b2a7f} /* (23, 25, 19) {real, imag} */,
  {32'h410b9dc8, 32'hc10c83ed} /* (23, 25, 18) {real, imag} */,
  {32'hc17ed4d7, 32'hc0aa5560} /* (23, 25, 17) {real, imag} */,
  {32'hc17587a4, 32'hc09736d4} /* (23, 25, 16) {real, imag} */,
  {32'hc14dd36f, 32'hc0c2fb90} /* (23, 25, 15) {real, imag} */,
  {32'h417c17b0, 32'h4177bc63} /* (23, 25, 14) {real, imag} */,
  {32'hc17c7e19, 32'hc1bb564a} /* (23, 25, 13) {real, imag} */,
  {32'h41e76c28, 32'h423b5ba2} /* (23, 25, 12) {real, imag} */,
  {32'hc081278e, 32'h413c1f8f} /* (23, 25, 11) {real, imag} */,
  {32'hc1722e64, 32'hc020530c} /* (23, 25, 10) {real, imag} */,
  {32'h41fdbae0, 32'h41301b7c} /* (23, 25, 9) {real, imag} */,
  {32'hc2f0cfab, 32'hbea09b00} /* (23, 25, 8) {real, imag} */,
  {32'hc188038f, 32'h40f3b4c9} /* (23, 25, 7) {real, imag} */,
  {32'hc113b547, 32'h42a44265} /* (23, 25, 6) {real, imag} */,
  {32'h417cc512, 32'h426aae95} /* (23, 25, 5) {real, imag} */,
  {32'h42e4a13f, 32'hc1280b90} /* (23, 25, 4) {real, imag} */,
  {32'hc24ee99a, 32'h420bbb94} /* (23, 25, 3) {real, imag} */,
  {32'h424d8556, 32'hc29d87ce} /* (23, 25, 2) {real, imag} */,
  {32'hc193ed36, 32'hc0d36f80} /* (23, 25, 1) {real, imag} */,
  {32'hc27e05fb, 32'hc25bce54} /* (23, 25, 0) {real, imag} */,
  {32'h429de164, 32'h41dd124c} /* (23, 24, 31) {real, imag} */,
  {32'h404ae808, 32'hc0e88c42} /* (23, 24, 30) {real, imag} */,
  {32'h41948684, 32'h421ed154} /* (23, 24, 29) {real, imag} */,
  {32'h41e2600e, 32'hc2a95e2c} /* (23, 24, 28) {real, imag} */,
  {32'hc2c1353c, 32'hc1f456e9} /* (23, 24, 27) {real, imag} */,
  {32'hc209d310, 32'hc1102125} /* (23, 24, 26) {real, imag} */,
  {32'hc17a6b7c, 32'h41aa3bd1} /* (23, 24, 25) {real, imag} */,
  {32'hc14b69f8, 32'hc1b68da2} /* (23, 24, 24) {real, imag} */,
  {32'hc0b4e4b8, 32'h42741840} /* (23, 24, 23) {real, imag} */,
  {32'h40a55b76, 32'h423bf026} /* (23, 24, 22) {real, imag} */,
  {32'h418d47ec, 32'hc133dd83} /* (23, 24, 21) {real, imag} */,
  {32'hc14bb575, 32'hc1a56bc1} /* (23, 24, 20) {real, imag} */,
  {32'hc181f876, 32'hbf91b2d8} /* (23, 24, 19) {real, imag} */,
  {32'h419c6dba, 32'hc00a1918} /* (23, 24, 18) {real, imag} */,
  {32'hc1010c33, 32'h41886980} /* (23, 24, 17) {real, imag} */,
  {32'hc1045230, 32'h41635639} /* (23, 24, 16) {real, imag} */,
  {32'hc1baa2da, 32'hc01cf920} /* (23, 24, 15) {real, imag} */,
  {32'h40170504, 32'h40cf53f8} /* (23, 24, 14) {real, imag} */,
  {32'hbf3e9da0, 32'hc1e730b6} /* (23, 24, 13) {real, imag} */,
  {32'hc05498ec, 32'hc0a14c34} /* (23, 24, 12) {real, imag} */,
  {32'hc1ec8d94, 32'hc17b3689} /* (23, 24, 11) {real, imag} */,
  {32'h4146654b, 32'h415e97b0} /* (23, 24, 10) {real, imag} */,
  {32'h3f345160, 32'hbf473ca0} /* (23, 24, 9) {real, imag} */,
  {32'hc18e88ac, 32'h4200f046} /* (23, 24, 8) {real, imag} */,
  {32'hc0b52374, 32'h407becf8} /* (23, 24, 7) {real, imag} */,
  {32'h42d15e8a, 32'h414b82e5} /* (23, 24, 6) {real, imag} */,
  {32'h40e6ea08, 32'h415ff55e} /* (23, 24, 5) {real, imag} */,
  {32'hc151e0f4, 32'h423226d0} /* (23, 24, 4) {real, imag} */,
  {32'h417eb1e9, 32'hc20ca02a} /* (23, 24, 3) {real, imag} */,
  {32'hc232c74a, 32'hc210011a} /* (23, 24, 2) {real, imag} */,
  {32'hc2b716bc, 32'h420770be} /* (23, 24, 1) {real, imag} */,
  {32'h431ddfba, 32'h4160e175} /* (23, 24, 0) {real, imag} */,
  {32'hc20871b2, 32'h41f8b241} /* (23, 23, 31) {real, imag} */,
  {32'h4217bdd0, 32'hc1e91f33} /* (23, 23, 30) {real, imag} */,
  {32'h41f2be43, 32'hbfaca280} /* (23, 23, 29) {real, imag} */,
  {32'h41785bb2, 32'h4249d2ab} /* (23, 23, 28) {real, imag} */,
  {32'h421e8482, 32'hc00edee0} /* (23, 23, 27) {real, imag} */,
  {32'h414a57e4, 32'h42187072} /* (23, 23, 26) {real, imag} */,
  {32'hc2573c8a, 32'h41beff37} /* (23, 23, 25) {real, imag} */,
  {32'hc206d01e, 32'h41934fe6} /* (23, 23, 24) {real, imag} */,
  {32'hc1ca8a3c, 32'h41b1570c} /* (23, 23, 23) {real, imag} */,
  {32'h41a9ac44, 32'hc2218165} /* (23, 23, 22) {real, imag} */,
  {32'hc1a92acf, 32'hc1823ad4} /* (23, 23, 21) {real, imag} */,
  {32'hc1aad1ec, 32'h41f9dcee} /* (23, 23, 20) {real, imag} */,
  {32'hc04d18d0, 32'hc0181974} /* (23, 23, 19) {real, imag} */,
  {32'hc0ea2b85, 32'hc1517c68} /* (23, 23, 18) {real, imag} */,
  {32'hc05a929c, 32'h4087934d} /* (23, 23, 17) {real, imag} */,
  {32'h3f849d48, 32'h416688fe} /* (23, 23, 16) {real, imag} */,
  {32'hc0a2cd72, 32'h41353414} /* (23, 23, 15) {real, imag} */,
  {32'h3d322280, 32'hbfc0d980} /* (23, 23, 14) {real, imag} */,
  {32'h41a32468, 32'h41a9c406} /* (23, 23, 13) {real, imag} */,
  {32'h4173ddd4, 32'hc16b2694} /* (23, 23, 12) {real, imag} */,
  {32'h419ba6c3, 32'h40cd347e} /* (23, 23, 11) {real, imag} */,
  {32'h3fc01548, 32'h423a6dff} /* (23, 23, 10) {real, imag} */,
  {32'hbfd9d0a0, 32'hc02ac1e0} /* (23, 23, 9) {real, imag} */,
  {32'h3fc3f610, 32'hc051793c} /* (23, 23, 8) {real, imag} */,
  {32'hc22b0036, 32'hc2024028} /* (23, 23, 7) {real, imag} */,
  {32'hc247a287, 32'h421b5410} /* (23, 23, 6) {real, imag} */,
  {32'hc17b0404, 32'h4106e38e} /* (23, 23, 5) {real, imag} */,
  {32'h41fbca09, 32'hc1e66966} /* (23, 23, 4) {real, imag} */,
  {32'h4163ddae, 32'hc12bd21a} /* (23, 23, 3) {real, imag} */,
  {32'h424a2fb6, 32'h421b5868} /* (23, 23, 2) {real, imag} */,
  {32'hc2595442, 32'hc2100e2c} /* (23, 23, 1) {real, imag} */,
  {32'hc1f6beaa, 32'hc29ae8a4} /* (23, 23, 0) {real, imag} */,
  {32'hc11bc20e, 32'h3ed0a120} /* (23, 22, 31) {real, imag} */,
  {32'h42bb4483, 32'hc0cc5106} /* (23, 22, 30) {real, imag} */,
  {32'hc242e442, 32'hc253824a} /* (23, 22, 29) {real, imag} */,
  {32'h3eeff074, 32'hc19f51e4} /* (23, 22, 28) {real, imag} */,
  {32'h4145da5c, 32'hc1b486d3} /* (23, 22, 27) {real, imag} */,
  {32'hc0640058, 32'h415117ba} /* (23, 22, 26) {real, imag} */,
  {32'hc1d80aac, 32'h4134b619} /* (23, 22, 25) {real, imag} */,
  {32'h411cdf3b, 32'h418583c9} /* (23, 22, 24) {real, imag} */,
  {32'h41220ea7, 32'hc1321c1c} /* (23, 22, 23) {real, imag} */,
  {32'hc0868c7d, 32'h419694b1} /* (23, 22, 22) {real, imag} */,
  {32'h41b2dc4b, 32'hbf0ab918} /* (23, 22, 21) {real, imag} */,
  {32'h412af84d, 32'h412b2208} /* (23, 22, 20) {real, imag} */,
  {32'hc036bd78, 32'h4118bb8c} /* (23, 22, 19) {real, imag} */,
  {32'hbffca890, 32'h41896992} /* (23, 22, 18) {real, imag} */,
  {32'hc143d658, 32'h414920b1} /* (23, 22, 17) {real, imag} */,
  {32'h411864e1, 32'hc17f419b} /* (23, 22, 16) {real, imag} */,
  {32'h4114b340, 32'h406f9bcc} /* (23, 22, 15) {real, imag} */,
  {32'h40ee38ac, 32'h418aee5a} /* (23, 22, 14) {real, imag} */,
  {32'hc1e0fb87, 32'h415fa060} /* (23, 22, 13) {real, imag} */,
  {32'hbfebca48, 32'h4201c921} /* (23, 22, 12) {real, imag} */,
  {32'h41a96541, 32'hc03af756} /* (23, 22, 11) {real, imag} */,
  {32'hc106da6a, 32'hc177ba16} /* (23, 22, 10) {real, imag} */,
  {32'h41e99050, 32'hc1c53006} /* (23, 22, 9) {real, imag} */,
  {32'hc12abe5b, 32'hc1e8165b} /* (23, 22, 8) {real, imag} */,
  {32'h41edeaec, 32'hbc85fc00} /* (23, 22, 7) {real, imag} */,
  {32'h419ea63f, 32'hc2170218} /* (23, 22, 6) {real, imag} */,
  {32'h4257bb85, 32'h41d2625b} /* (23, 22, 5) {real, imag} */,
  {32'h404ab040, 32'hc1229845} /* (23, 22, 4) {real, imag} */,
  {32'h40eeadf4, 32'h419f3464} /* (23, 22, 3) {real, imag} */,
  {32'hc24912a2, 32'h41467b59} /* (23, 22, 2) {real, imag} */,
  {32'h419823eb, 32'h41c43a5a} /* (23, 22, 1) {real, imag} */,
  {32'hc1d5f358, 32'hc197d244} /* (23, 22, 0) {real, imag} */,
  {32'h42313422, 32'hc12e9ae6} /* (23, 21, 31) {real, imag} */,
  {32'hc07f8f63, 32'hc1d69f64} /* (23, 21, 30) {real, imag} */,
  {32'hc1fb5d21, 32'hc285d6b2} /* (23, 21, 29) {real, imag} */,
  {32'h41cb3b3c, 32'h41a24d3a} /* (23, 21, 28) {real, imag} */,
  {32'h4233f14a, 32'hc253038f} /* (23, 21, 27) {real, imag} */,
  {32'h41551cee, 32'hc1f5976b} /* (23, 21, 26) {real, imag} */,
  {32'h41e7625e, 32'hc1a7476b} /* (23, 21, 25) {real, imag} */,
  {32'h41b67d04, 32'hc1907434} /* (23, 21, 24) {real, imag} */,
  {32'h4203871e, 32'h3fb10f86} /* (23, 21, 23) {real, imag} */,
  {32'h416987d8, 32'hc205d35e} /* (23, 21, 22) {real, imag} */,
  {32'hc19cb933, 32'h3fc8cd08} /* (23, 21, 21) {real, imag} */,
  {32'h41124ca1, 32'hc0fd9212} /* (23, 21, 20) {real, imag} */,
  {32'h3f9f4710, 32'hc124f199} /* (23, 21, 19) {real, imag} */,
  {32'h4115d313, 32'hc05b5018} /* (23, 21, 18) {real, imag} */,
  {32'hc110f31a, 32'hc0f0df89} /* (23, 21, 17) {real, imag} */,
  {32'hbfd36880, 32'h40bef81a} /* (23, 21, 16) {real, imag} */,
  {32'h40d26758, 32'h41554398} /* (23, 21, 15) {real, imag} */,
  {32'hbf9ce3d8, 32'hc11b6aae} /* (23, 21, 14) {real, imag} */,
  {32'h412f2fb2, 32'h40bde3be} /* (23, 21, 13) {real, imag} */,
  {32'h40e2302e, 32'h4158cbe3} /* (23, 21, 12) {real, imag} */,
  {32'hc1abfbb3, 32'h41aedbe0} /* (23, 21, 11) {real, imag} */,
  {32'hbf2d2ae0, 32'hc176a6d2} /* (23, 21, 10) {real, imag} */,
  {32'hc21b912e, 32'h4091254a} /* (23, 21, 9) {real, imag} */,
  {32'h4216f8f4, 32'h4028e3e8} /* (23, 21, 8) {real, imag} */,
  {32'h424bc205, 32'hc1e4afcd} /* (23, 21, 7) {real, imag} */,
  {32'h418f9cb6, 32'hc1f41f31} /* (23, 21, 6) {real, imag} */,
  {32'hc2700c7e, 32'hc19a344a} /* (23, 21, 5) {real, imag} */,
  {32'hc1c13bec, 32'h40e7f0cd} /* (23, 21, 4) {real, imag} */,
  {32'hc22d6160, 32'h416f4728} /* (23, 21, 3) {real, imag} */,
  {32'hc0a2a3f6, 32'h4216bb10} /* (23, 21, 2) {real, imag} */,
  {32'hc1440618, 32'h415f7c22} /* (23, 21, 1) {real, imag} */,
  {32'hc23c5390, 32'hc19743ca} /* (23, 21, 0) {real, imag} */,
  {32'h4217adde, 32'h41bc2772} /* (23, 20, 31) {real, imag} */,
  {32'h420dbaee, 32'hc0fe3526} /* (23, 20, 30) {real, imag} */,
  {32'hc1b14f5c, 32'hbf22e2f0} /* (23, 20, 29) {real, imag} */,
  {32'h41083dee, 32'hc0a3f550} /* (23, 20, 28) {real, imag} */,
  {32'h41846d40, 32'h41c75f4f} /* (23, 20, 27) {real, imag} */,
  {32'h41106ce2, 32'hc12d5f7b} /* (23, 20, 26) {real, imag} */,
  {32'h419aa42c, 32'hc07f28e8} /* (23, 20, 25) {real, imag} */,
  {32'hbf0d69d8, 32'hc1a60217} /* (23, 20, 24) {real, imag} */,
  {32'h3db02680, 32'h41aa969b} /* (23, 20, 23) {real, imag} */,
  {32'hc0e273d0, 32'hc15fea1b} /* (23, 20, 22) {real, imag} */,
  {32'h4131ba96, 32'h40b458b2} /* (23, 20, 21) {real, imag} */,
  {32'h40e0c1d1, 32'h3f534880} /* (23, 20, 20) {real, imag} */,
  {32'h4113fa11, 32'hc10c585c} /* (23, 20, 19) {real, imag} */,
  {32'h401a26ac, 32'h408c9aa4} /* (23, 20, 18) {real, imag} */,
  {32'hbfbbefc0, 32'h4080bb8a} /* (23, 20, 17) {real, imag} */,
  {32'hc1312856, 32'h407b9384} /* (23, 20, 16) {real, imag} */,
  {32'h4131fa0c, 32'hc045dfec} /* (23, 20, 15) {real, imag} */,
  {32'h41834268, 32'hc006e8d8} /* (23, 20, 14) {real, imag} */,
  {32'h412d3dbb, 32'h401b01d1} /* (23, 20, 13) {real, imag} */,
  {32'h3ffa95e4, 32'hbefe04e0} /* (23, 20, 12) {real, imag} */,
  {32'h41342bf8, 32'hc1d73cec} /* (23, 20, 11) {real, imag} */,
  {32'hc12f7c48, 32'h411a87f3} /* (23, 20, 10) {real, imag} */,
  {32'hc1258b4f, 32'hc1db2949} /* (23, 20, 9) {real, imag} */,
  {32'h418056c3, 32'hc155b167} /* (23, 20, 8) {real, imag} */,
  {32'hc0eb5d0a, 32'h41ac0d8f} /* (23, 20, 7) {real, imag} */,
  {32'hc2169408, 32'hc2058bed} /* (23, 20, 6) {real, imag} */,
  {32'hc13949e7, 32'h41ee2075} /* (23, 20, 5) {real, imag} */,
  {32'hc0539cf2, 32'hc1cae3ea} /* (23, 20, 4) {real, imag} */,
  {32'hc2150edb, 32'hc0a8368d} /* (23, 20, 3) {real, imag} */,
  {32'hc12a55e6, 32'hc0ce15aa} /* (23, 20, 2) {real, imag} */,
  {32'h41ec5bdb, 32'hc227c8df} /* (23, 20, 1) {real, imag} */,
  {32'hc1cadcf1, 32'hc10ba776} /* (23, 20, 0) {real, imag} */,
  {32'hc2171710, 32'h413a8fc8} /* (23, 19, 31) {real, imag} */,
  {32'hc1456c06, 32'h41bae1ec} /* (23, 19, 30) {real, imag} */,
  {32'hc1198c5d, 32'h420db04c} /* (23, 19, 29) {real, imag} */,
  {32'h4230728b, 32'hc1318b38} /* (23, 19, 28) {real, imag} */,
  {32'hc22202dc, 32'hc190045c} /* (23, 19, 27) {real, imag} */,
  {32'h3f282e20, 32'hc14bcbf1} /* (23, 19, 26) {real, imag} */,
  {32'hbeafd790, 32'h3eb76070} /* (23, 19, 25) {real, imag} */,
  {32'hc16db2e4, 32'h41108002} /* (23, 19, 24) {real, imag} */,
  {32'hc1a9cac2, 32'hc178e696} /* (23, 19, 23) {real, imag} */,
  {32'hc186a16b, 32'hc130c49a} /* (23, 19, 22) {real, imag} */,
  {32'h41af6572, 32'h411cd4f6} /* (23, 19, 21) {real, imag} */,
  {32'hbfeb0b78, 32'hc17ab6a7} /* (23, 19, 20) {real, imag} */,
  {32'h409d8b7a, 32'hc103a3ac} /* (23, 19, 19) {real, imag} */,
  {32'h3f196908, 32'hc0229c3e} /* (23, 19, 18) {real, imag} */,
  {32'hc06e1d4c, 32'h3feecd56} /* (23, 19, 17) {real, imag} */,
  {32'hbf3ecf08, 32'hbee26c10} /* (23, 19, 16) {real, imag} */,
  {32'h40a3ccfa, 32'hc0ac277e} /* (23, 19, 15) {real, imag} */,
  {32'h3fd22d44, 32'h3f14e368} /* (23, 19, 14) {real, imag} */,
  {32'h40292645, 32'hc17010e6} /* (23, 19, 13) {real, imag} */,
  {32'hbf803a58, 32'h414cb6a3} /* (23, 19, 12) {real, imag} */,
  {32'h3fc3eb38, 32'hc06d6e97} /* (23, 19, 11) {real, imag} */,
  {32'h4104aa32, 32'h4123bdc6} /* (23, 19, 10) {real, imag} */,
  {32'h40667184, 32'h410dce4a} /* (23, 19, 9) {real, imag} */,
  {32'h41162a8c, 32'h41d3a725} /* (23, 19, 8) {real, imag} */,
  {32'h409cd22b, 32'hc0d0ef9f} /* (23, 19, 7) {real, imag} */,
  {32'hc193dce3, 32'h4127322f} /* (23, 19, 6) {real, imag} */,
  {32'h40bb7404, 32'h41191e78} /* (23, 19, 5) {real, imag} */,
  {32'h40f6f468, 32'h42273f18} /* (23, 19, 4) {real, imag} */,
  {32'h4001da8c, 32'hc1acc3d4} /* (23, 19, 3) {real, imag} */,
  {32'h42003218, 32'h4094b316} /* (23, 19, 2) {real, imag} */,
  {32'hc0cd3e7c, 32'h41b788c2} /* (23, 19, 1) {real, imag} */,
  {32'hc02af172, 32'h40eb78b1} /* (23, 19, 0) {real, imag} */,
  {32'hc16736bf, 32'hc1d2f166} /* (23, 18, 31) {real, imag} */,
  {32'hc1a227ed, 32'hbfaf4696} /* (23, 18, 30) {real, imag} */,
  {32'h40f74a3c, 32'hc1b8d046} /* (23, 18, 29) {real, imag} */,
  {32'h420c410c, 32'hc224f5c0} /* (23, 18, 28) {real, imag} */,
  {32'h4154b3ba, 32'hc0633ba8} /* (23, 18, 27) {real, imag} */,
  {32'h3f8e5924, 32'hbff0deff} /* (23, 18, 26) {real, imag} */,
  {32'hc22cf9c2, 32'h41374ae5} /* (23, 18, 25) {real, imag} */,
  {32'h415bfce8, 32'h41784d14} /* (23, 18, 24) {real, imag} */,
  {32'hc13218f1, 32'hc1083e06} /* (23, 18, 23) {real, imag} */,
  {32'hc0480049, 32'hc18d597a} /* (23, 18, 22) {real, imag} */,
  {32'h40c3d99e, 32'hc0eefca9} /* (23, 18, 21) {real, imag} */,
  {32'hc069ff0a, 32'h3ea3f178} /* (23, 18, 20) {real, imag} */,
  {32'h3d90ea00, 32'hbfe1d02c} /* (23, 18, 19) {real, imag} */,
  {32'hc01adc54, 32'h404284f9} /* (23, 18, 18) {real, imag} */,
  {32'hc0015a35, 32'h3e847bb0} /* (23, 18, 17) {real, imag} */,
  {32'hc0120ada, 32'hbff708a8} /* (23, 18, 16) {real, imag} */,
  {32'h3fd56ed6, 32'h40ca9dc3} /* (23, 18, 15) {real, imag} */,
  {32'hbce7ea00, 32'hbfb17d56} /* (23, 18, 14) {real, imag} */,
  {32'hc0caec28, 32'h4107d9c8} /* (23, 18, 13) {real, imag} */,
  {32'hc07f9036, 32'hc0d65070} /* (23, 18, 12) {real, imag} */,
  {32'hc0d8314a, 32'h4105c6f4} /* (23, 18, 11) {real, imag} */,
  {32'h3fd85b36, 32'h412babc4} /* (23, 18, 10) {real, imag} */,
  {32'h3f07f510, 32'h414ded48} /* (23, 18, 9) {real, imag} */,
  {32'hc0e9ec70, 32'h3f6855a8} /* (23, 18, 8) {real, imag} */,
  {32'hc1b5fb48, 32'h413fbf87} /* (23, 18, 7) {real, imag} */,
  {32'hc155080e, 32'h4097c568} /* (23, 18, 6) {real, imag} */,
  {32'hbed76030, 32'h41d478c7} /* (23, 18, 5) {real, imag} */,
  {32'h418de397, 32'hc231c378} /* (23, 18, 4) {real, imag} */,
  {32'hc1f1ea8b, 32'hc08f4a16} /* (23, 18, 3) {real, imag} */,
  {32'hc1fad973, 32'h410d8173} /* (23, 18, 2) {real, imag} */,
  {32'h4157a719, 32'hc0f73310} /* (23, 18, 1) {real, imag} */,
  {32'hc0d10f5f, 32'hc1ed053a} /* (23, 18, 0) {real, imag} */,
  {32'hc1ca7449, 32'hc1b32ab2} /* (23, 17, 31) {real, imag} */,
  {32'hbf700fdc, 32'hc1797fb8} /* (23, 17, 30) {real, imag} */,
  {32'h406c1d00, 32'h40f48078} /* (23, 17, 29) {real, imag} */,
  {32'hc1b2cc38, 32'h3fa37e8c} /* (23, 17, 28) {real, imag} */,
  {32'hc138493a, 32'h40a024b6} /* (23, 17, 27) {real, imag} */,
  {32'hc1aef25b, 32'hc0ec4902} /* (23, 17, 26) {real, imag} */,
  {32'h40c1738c, 32'h41171d8c} /* (23, 17, 25) {real, imag} */,
  {32'h41a5af42, 32'h4062ed9e} /* (23, 17, 24) {real, imag} */,
  {32'hc0515f86, 32'h4089b046} /* (23, 17, 23) {real, imag} */,
  {32'h411df8a0, 32'hc1613a76} /* (23, 17, 22) {real, imag} */,
  {32'hc12191fb, 32'hc0a4736b} /* (23, 17, 21) {real, imag} */,
  {32'hc0a836f4, 32'h40d2ff22} /* (23, 17, 20) {real, imag} */,
  {32'h412c18b4, 32'h3fef70b2} /* (23, 17, 19) {real, imag} */,
  {32'h40d89d92, 32'h40c6ca24} /* (23, 17, 18) {real, imag} */,
  {32'h411bea26, 32'hc0835637} /* (23, 17, 17) {real, imag} */,
  {32'hc02038e6, 32'h40401760} /* (23, 17, 16) {real, imag} */,
  {32'h402718a8, 32'h3fd6b254} /* (23, 17, 15) {real, imag} */,
  {32'h3f545c0c, 32'hbfb6de70} /* (23, 17, 14) {real, imag} */,
  {32'h40b0dfa7, 32'hc102a732} /* (23, 17, 13) {real, imag} */,
  {32'hbff5607e, 32'h40f6a562} /* (23, 17, 12) {real, imag} */,
  {32'hbf9a68c0, 32'hc0c56271} /* (23, 17, 11) {real, imag} */,
  {32'hc15b0018, 32'h40cdc635} /* (23, 17, 10) {real, imag} */,
  {32'hc0cd4195, 32'h405194fd} /* (23, 17, 9) {real, imag} */,
  {32'hc0e2ca0c, 32'h40bad4fd} /* (23, 17, 8) {real, imag} */,
  {32'hc17c8e42, 32'h411c7eb6} /* (23, 17, 7) {real, imag} */,
  {32'h40b9609c, 32'hc0219a3f} /* (23, 17, 6) {real, imag} */,
  {32'h40e2181b, 32'hc1ced1ec} /* (23, 17, 5) {real, imag} */,
  {32'hc1513797, 32'h41319bb0} /* (23, 17, 4) {real, imag} */,
  {32'h41c12d6c, 32'hc1ca27d2} /* (23, 17, 3) {real, imag} */,
  {32'h40649497, 32'hc17217a8} /* (23, 17, 2) {real, imag} */,
  {32'hc097d16c, 32'h3ecbd7e0} /* (23, 17, 1) {real, imag} */,
  {32'h413b6ac8, 32'h4100adc6} /* (23, 17, 0) {real, imag} */,
  {32'h4196cd39, 32'hc1a8d8fc} /* (23, 16, 31) {real, imag} */,
  {32'hc0fefcd8, 32'h3ffacce9} /* (23, 16, 30) {real, imag} */,
  {32'hc1057d25, 32'hc104354b} /* (23, 16, 29) {real, imag} */,
  {32'h4107c175, 32'h41c860b3} /* (23, 16, 28) {real, imag} */,
  {32'h41bf7e16, 32'h4180f1b8} /* (23, 16, 27) {real, imag} */,
  {32'h3fce5ed4, 32'hc1a192d8} /* (23, 16, 26) {real, imag} */,
  {32'h410c2962, 32'hc1682875} /* (23, 16, 25) {real, imag} */,
  {32'h40c2212f, 32'hc17446e1} /* (23, 16, 24) {real, imag} */,
  {32'h3e8d6bf0, 32'h40d52ef8} /* (23, 16, 23) {real, imag} */,
  {32'h40168ed6, 32'hc0841896} /* (23, 16, 22) {real, imag} */,
  {32'h403258e0, 32'hc140664a} /* (23, 16, 21) {real, imag} */,
  {32'hc0a7c4b8, 32'h40ef5255} /* (23, 16, 20) {real, imag} */,
  {32'hc124f9e8, 32'h40929f92} /* (23, 16, 19) {real, imag} */,
  {32'hc0e4698a, 32'h3fa19b0e} /* (23, 16, 18) {real, imag} */,
  {32'h40a6099a, 32'h401547c2} /* (23, 16, 17) {real, imag} */,
  {32'hc039e0d6, 32'h4103c884} /* (23, 16, 16) {real, imag} */,
  {32'hc0ab4756, 32'h40dd9e2f} /* (23, 16, 15) {real, imag} */,
  {32'h3fcd9db8, 32'h3f3cf488} /* (23, 16, 14) {real, imag} */,
  {32'h40a07c27, 32'h3f2ba020} /* (23, 16, 13) {real, imag} */,
  {32'hc0e0623a, 32'hc1847305} /* (23, 16, 12) {real, imag} */,
  {32'hbf79fca0, 32'h40ff75fc} /* (23, 16, 11) {real, imag} */,
  {32'h40279a5a, 32'hc1182183} /* (23, 16, 10) {real, imag} */,
  {32'h40ffee8f, 32'hc0f49720} /* (23, 16, 9) {real, imag} */,
  {32'hc0d95689, 32'h40cb59be} /* (23, 16, 8) {real, imag} */,
  {32'hc023aa18, 32'h40e4eaf6} /* (23, 16, 7) {real, imag} */,
  {32'h413e1a8e, 32'hc138b542} /* (23, 16, 6) {real, imag} */,
  {32'h40556538, 32'hc0a0fb20} /* (23, 16, 5) {real, imag} */,
  {32'h4078be28, 32'hc17e524e} /* (23, 16, 4) {real, imag} */,
  {32'h41046913, 32'h413e2021} /* (23, 16, 3) {real, imag} */,
  {32'h4143bd04, 32'h4076585c} /* (23, 16, 2) {real, imag} */,
  {32'hc0f542bb, 32'hc126742d} /* (23, 16, 1) {real, imag} */,
  {32'h41284b8a, 32'h41fac0d2} /* (23, 16, 0) {real, imag} */,
  {32'h41839134, 32'h41229df0} /* (23, 15, 31) {real, imag} */,
  {32'hbd5af2a0, 32'h41cb6e68} /* (23, 15, 30) {real, imag} */,
  {32'hc05b7b12, 32'hc140a84c} /* (23, 15, 29) {real, imag} */,
  {32'h419836a8, 32'h417472fc} /* (23, 15, 28) {real, imag} */,
  {32'hc095ebcd, 32'h3fc53100} /* (23, 15, 27) {real, imag} */,
  {32'hc13d28be, 32'h41cdf444} /* (23, 15, 26) {real, imag} */,
  {32'hc0a78f04, 32'hc119847d} /* (23, 15, 25) {real, imag} */,
  {32'hc0074008, 32'hc110421a} /* (23, 15, 24) {real, imag} */,
  {32'h4197bb61, 32'hc0625e99} /* (23, 15, 23) {real, imag} */,
  {32'h402b5f69, 32'hc124cdd1} /* (23, 15, 22) {real, imag} */,
  {32'hc0cea368, 32'h41960dd8} /* (23, 15, 21) {real, imag} */,
  {32'h407c87d6, 32'hc117c780} /* (23, 15, 20) {real, imag} */,
  {32'hbf3d9bb4, 32'h40e95507} /* (23, 15, 19) {real, imag} */,
  {32'hbfae87e7, 32'h401d7690} /* (23, 15, 18) {real, imag} */,
  {32'hc0452817, 32'hbfed8bb8} /* (23, 15, 17) {real, imag} */,
  {32'hc0d46b38, 32'hbeae3920} /* (23, 15, 16) {real, imag} */,
  {32'hc0892510, 32'h40cfd3d6} /* (23, 15, 15) {real, imag} */,
  {32'h3f8157ad, 32'hc063dbb8} /* (23, 15, 14) {real, imag} */,
  {32'h40a0bda8, 32'hc068411e} /* (23, 15, 13) {real, imag} */,
  {32'h408f59b3, 32'hc09a44f1} /* (23, 15, 12) {real, imag} */,
  {32'hc0ac629e, 32'hbece2e80} /* (23, 15, 11) {real, imag} */,
  {32'h4080174c, 32'hc02cde7c} /* (23, 15, 10) {real, imag} */,
  {32'h41861579, 32'hc0e21e08} /* (23, 15, 9) {real, imag} */,
  {32'h4211e112, 32'hc171b084} /* (23, 15, 8) {real, imag} */,
  {32'h3f7039a4, 32'hc116da39} /* (23, 15, 7) {real, imag} */,
  {32'hc19c3f5f, 32'h419c0084} /* (23, 15, 6) {real, imag} */,
  {32'h40ac099b, 32'hc1dd6b46} /* (23, 15, 5) {real, imag} */,
  {32'hc1a97892, 32'h3fdcfebc} /* (23, 15, 4) {real, imag} */,
  {32'h4182af92, 32'hc11144de} /* (23, 15, 3) {real, imag} */,
  {32'h40315e4c, 32'h41e7c3f8} /* (23, 15, 2) {real, imag} */,
  {32'hc16971e6, 32'hc1852323} /* (23, 15, 1) {real, imag} */,
  {32'h41dfac58, 32'h4026c54c} /* (23, 15, 0) {real, imag} */,
  {32'hc0e5847e, 32'hc14135e5} /* (23, 14, 31) {real, imag} */,
  {32'hc16facf2, 32'h41b96ce5} /* (23, 14, 30) {real, imag} */,
  {32'h419b47aa, 32'hc186fc7a} /* (23, 14, 29) {real, imag} */,
  {32'hc16c2df8, 32'hc16efa04} /* (23, 14, 28) {real, imag} */,
  {32'h4166fcc4, 32'hc20bd2c0} /* (23, 14, 27) {real, imag} */,
  {32'h417e2020, 32'hc0d5ed6c} /* (23, 14, 26) {real, imag} */,
  {32'hc1a46f40, 32'hbf8c3fb8} /* (23, 14, 25) {real, imag} */,
  {32'hc1bbc7a2, 32'h41938e71} /* (23, 14, 24) {real, imag} */,
  {32'hc08e08eb, 32'h4146daeb} /* (23, 14, 23) {real, imag} */,
  {32'h4125b960, 32'h40f8115a} /* (23, 14, 22) {real, imag} */,
  {32'hbf1b933e, 32'h4111ba7a} /* (23, 14, 21) {real, imag} */,
  {32'h40f62384, 32'hbf88a230} /* (23, 14, 20) {real, imag} */,
  {32'h409241d2, 32'h40cda78a} /* (23, 14, 19) {real, imag} */,
  {32'h406386fa, 32'hc079861c} /* (23, 14, 18) {real, imag} */,
  {32'h40391b21, 32'h40a2608c} /* (23, 14, 17) {real, imag} */,
  {32'hc0051ca9, 32'h404778e0} /* (23, 14, 16) {real, imag} */,
  {32'hc0bd8704, 32'hc0572258} /* (23, 14, 15) {real, imag} */,
  {32'h4093a4df, 32'h3f7072b0} /* (23, 14, 14) {real, imag} */,
  {32'hc037c673, 32'h40672014} /* (23, 14, 13) {real, imag} */,
  {32'h412e828c, 32'hc1a2bd85} /* (23, 14, 12) {real, imag} */,
  {32'h3e23b588, 32'h41461d16} /* (23, 14, 11) {real, imag} */,
  {32'h418412c1, 32'hc0955cea} /* (23, 14, 10) {real, imag} */,
  {32'h404c1c62, 32'h3f86bc28} /* (23, 14, 9) {real, imag} */,
  {32'hbfad53c0, 32'hc06ed1c8} /* (23, 14, 8) {real, imag} */,
  {32'h40dbf165, 32'hc0f2fdba} /* (23, 14, 7) {real, imag} */,
  {32'h40a67c2b, 32'h4135aa98} /* (23, 14, 6) {real, imag} */,
  {32'hc1acdd3e, 32'h400ee108} /* (23, 14, 5) {real, imag} */,
  {32'hc140cece, 32'h41867d4e} /* (23, 14, 4) {real, imag} */,
  {32'hc054e1d4, 32'hc13dcbe6} /* (23, 14, 3) {real, imag} */,
  {32'h416f759e, 32'h41f65c51} /* (23, 14, 2) {real, imag} */,
  {32'h40d97d86, 32'hc1b50e72} /* (23, 14, 1) {real, imag} */,
  {32'h4085f174, 32'h4116ce56} /* (23, 14, 0) {real, imag} */,
  {32'h4105f17d, 32'h41e106df} /* (23, 13, 31) {real, imag} */,
  {32'hc06e7828, 32'h414e9b3c} /* (23, 13, 30) {real, imag} */,
  {32'h4155637d, 32'hc1d3f00a} /* (23, 13, 29) {real, imag} */,
  {32'hc184c944, 32'h4238d4ff} /* (23, 13, 28) {real, imag} */,
  {32'hc0b7b98e, 32'hc1963e6b} /* (23, 13, 27) {real, imag} */,
  {32'hc1adc0ad, 32'h403eb268} /* (23, 13, 26) {real, imag} */,
  {32'hc06959c4, 32'hbf9ddb78} /* (23, 13, 25) {real, imag} */,
  {32'hbfdaf060, 32'h40c3ea02} /* (23, 13, 24) {real, imag} */,
  {32'h40d13ee8, 32'h4088dbeb} /* (23, 13, 23) {real, imag} */,
  {32'hc1becc92, 32'hbff3db20} /* (23, 13, 22) {real, imag} */,
  {32'hc08fb16b, 32'h418bd494} /* (23, 13, 21) {real, imag} */,
  {32'hc05df290, 32'hc0502a26} /* (23, 13, 20) {real, imag} */,
  {32'h411c0f39, 32'hbf0ac9c8} /* (23, 13, 19) {real, imag} */,
  {32'h406f6750, 32'hc0d89a3d} /* (23, 13, 18) {real, imag} */,
  {32'h4096895e, 32'hc14b9a81} /* (23, 13, 17) {real, imag} */,
  {32'h3f0784c0, 32'h3f8eca60} /* (23, 13, 16) {real, imag} */,
  {32'hc0f89216, 32'h40d94786} /* (23, 13, 15) {real, imag} */,
  {32'h40edddf4, 32'h40883959} /* (23, 13, 14) {real, imag} */,
  {32'h40a8824a, 32'h410e66a0} /* (23, 13, 13) {real, imag} */,
  {32'h40fcdb4c, 32'h41721faa} /* (23, 13, 12) {real, imag} */,
  {32'hc162e0a8, 32'hc008728c} /* (23, 13, 11) {real, imag} */,
  {32'hc15ddd80, 32'hc02698bc} /* (23, 13, 10) {real, imag} */,
  {32'hc08cdbb0, 32'h4106e4e8} /* (23, 13, 9) {real, imag} */,
  {32'h41db150a, 32'hc15a4897} /* (23, 13, 8) {real, imag} */,
  {32'h416e1213, 32'hc0e69966} /* (23, 13, 7) {real, imag} */,
  {32'hbf3e1da0, 32'hc0f9f576} /* (23, 13, 6) {real, imag} */,
  {32'h413abd99, 32'hc1e534f1} /* (23, 13, 5) {real, imag} */,
  {32'hc1d3d4ac, 32'hc0aff9a0} /* (23, 13, 4) {real, imag} */,
  {32'h41445959, 32'h41696240} /* (23, 13, 3) {real, imag} */,
  {32'hc149f5dc, 32'hc0732ad8} /* (23, 13, 2) {real, imag} */,
  {32'hbe4c3740, 32'h41051722} /* (23, 13, 1) {real, imag} */,
  {32'hc2084ef5, 32'h42822d30} /* (23, 13, 0) {real, imag} */,
  {32'h40b4f889, 32'h41dad4f9} /* (23, 12, 31) {real, imag} */,
  {32'hc1ca7a1a, 32'h415d3e12} /* (23, 12, 30) {real, imag} */,
  {32'hc2047b78, 32'h420b4c65} /* (23, 12, 29) {real, imag} */,
  {32'h4155ee32, 32'hc18c8707} /* (23, 12, 28) {real, imag} */,
  {32'h409fb9f0, 32'hbf588f18} /* (23, 12, 27) {real, imag} */,
  {32'h418315c2, 32'h42020ab3} /* (23, 12, 26) {real, imag} */,
  {32'hc1924782, 32'h40edf8bc} /* (23, 12, 25) {real, imag} */,
  {32'h41988f6c, 32'h414468d4} /* (23, 12, 24) {real, imag} */,
  {32'hc18c83dc, 32'h41495e5e} /* (23, 12, 23) {real, imag} */,
  {32'h41603907, 32'h41292a2c} /* (23, 12, 22) {real, imag} */,
  {32'hc1885942, 32'hc1996d7c} /* (23, 12, 21) {real, imag} */,
  {32'hc058e316, 32'hc0f8a5e8} /* (23, 12, 20) {real, imag} */,
  {32'h410a610e, 32'hbfc9e67c} /* (23, 12, 19) {real, imag} */,
  {32'hc0496668, 32'hc126b08f} /* (23, 12, 18) {real, imag} */,
  {32'hc05b1e5e, 32'hc050d0f8} /* (23, 12, 17) {real, imag} */,
  {32'hbff71d20, 32'hc0b5d6e1} /* (23, 12, 16) {real, imag} */,
  {32'h40210c8a, 32'hc0562028} /* (23, 12, 15) {real, imag} */,
  {32'h409c198c, 32'h410cc531} /* (23, 12, 14) {real, imag} */,
  {32'h40878105, 32'hc170c754} /* (23, 12, 13) {real, imag} */,
  {32'h411beb84, 32'h41e4fc4a} /* (23, 12, 12) {real, imag} */,
  {32'hc13ebf48, 32'h3def7400} /* (23, 12, 11) {real, imag} */,
  {32'hc0aa4182, 32'hc0ade538} /* (23, 12, 10) {real, imag} */,
  {32'hc20cf01f, 32'hc05e95f8} /* (23, 12, 9) {real, imag} */,
  {32'hc18fdac4, 32'h3fef5724} /* (23, 12, 8) {real, imag} */,
  {32'h40e38722, 32'hc22e3f24} /* (23, 12, 7) {real, imag} */,
  {32'h408d628f, 32'h409e3398} /* (23, 12, 6) {real, imag} */,
  {32'hc1e0e352, 32'h406edb0e} /* (23, 12, 5) {real, imag} */,
  {32'h41863268, 32'hc162db8e} /* (23, 12, 4) {real, imag} */,
  {32'h41aca749, 32'h41518e78} /* (23, 12, 3) {real, imag} */,
  {32'h41b5a816, 32'hc141dc0e} /* (23, 12, 2) {real, imag} */,
  {32'h4121a11e, 32'hc0b65b04} /* (23, 12, 1) {real, imag} */,
  {32'h41b4fe36, 32'hc0753882} /* (23, 12, 0) {real, imag} */,
  {32'h4112e78b, 32'h40cf12c7} /* (23, 11, 31) {real, imag} */,
  {32'h419d703b, 32'hc1dc2bee} /* (23, 11, 30) {real, imag} */,
  {32'hbfbf093c, 32'h411339c8} /* (23, 11, 29) {real, imag} */,
  {32'hc22a08a4, 32'h41ff76ea} /* (23, 11, 28) {real, imag} */,
  {32'h424be90d, 32'hc0dc1e9a} /* (23, 11, 27) {real, imag} */,
  {32'h40e1709c, 32'h4236887f} /* (23, 11, 26) {real, imag} */,
  {32'h40f425d6, 32'h41404ebd} /* (23, 11, 25) {real, imag} */,
  {32'h40a00744, 32'hc187408f} /* (23, 11, 24) {real, imag} */,
  {32'hc22edbca, 32'hc01fa617} /* (23, 11, 23) {real, imag} */,
  {32'hc10bb725, 32'hc182b8c6} /* (23, 11, 22) {real, imag} */,
  {32'h41833766, 32'hc13cad23} /* (23, 11, 21) {real, imag} */,
  {32'h41346020, 32'hc0b9ea56} /* (23, 11, 20) {real, imag} */,
  {32'hc057d628, 32'hbf617bf0} /* (23, 11, 19) {real, imag} */,
  {32'hc09b0ceb, 32'h3f874b14} /* (23, 11, 18) {real, imag} */,
  {32'h3de5f160, 32'h4080f0ff} /* (23, 11, 17) {real, imag} */,
  {32'h3e277f80, 32'h401d87f0} /* (23, 11, 16) {real, imag} */,
  {32'h40831dce, 32'hc0d7a449} /* (23, 11, 15) {real, imag} */,
  {32'h4191c61f, 32'h40a299e5} /* (23, 11, 14) {real, imag} */,
  {32'hc0ab96f6, 32'hc181d58c} /* (23, 11, 13) {real, imag} */,
  {32'hc11ff7c8, 32'hc0601f53} /* (23, 11, 12) {real, imag} */,
  {32'hc0f8d2e0, 32'hc0a96b36} /* (23, 11, 11) {real, imag} */,
  {32'hbed7fce0, 32'hc155ec4c} /* (23, 11, 10) {real, imag} */,
  {32'hc0a0b818, 32'h40857528} /* (23, 11, 9) {real, imag} */,
  {32'h3e532050, 32'hc141804a} /* (23, 11, 8) {real, imag} */,
  {32'h4213d34c, 32'hc1745279} /* (23, 11, 7) {real, imag} */,
  {32'h426220fc, 32'h42061bf9} /* (23, 11, 6) {real, imag} */,
  {32'hc137b400, 32'hc1f2b006} /* (23, 11, 5) {real, imag} */,
  {32'hc144e53a, 32'h4232d581} /* (23, 11, 4) {real, imag} */,
  {32'hc12f00b4, 32'hc21b303a} /* (23, 11, 3) {real, imag} */,
  {32'h41a3e4cd, 32'h421f066b} /* (23, 11, 2) {real, imag} */,
  {32'hc1ca62c0, 32'hc177f0b0} /* (23, 11, 1) {real, imag} */,
  {32'h41907abd, 32'hc1c25506} /* (23, 11, 0) {real, imag} */,
  {32'h41fed8c6, 32'h41f68e2c} /* (23, 10, 31) {real, imag} */,
  {32'h40a0648d, 32'hc0aa73d0} /* (23, 10, 30) {real, imag} */,
  {32'h4210f10f, 32'h3f70d560} /* (23, 10, 29) {real, imag} */,
  {32'h410f2024, 32'h429608ca} /* (23, 10, 28) {real, imag} */,
  {32'h40333ece, 32'hc1a67419} /* (23, 10, 27) {real, imag} */,
  {32'h414743ff, 32'hc2473cf0} /* (23, 10, 26) {real, imag} */,
  {32'h417ba254, 32'h408c83f6} /* (23, 10, 25) {real, imag} */,
  {32'hc144da2f, 32'h4095d120} /* (23, 10, 24) {real, imag} */,
  {32'h40cf5e62, 32'hc1e17741} /* (23, 10, 23) {real, imag} */,
  {32'h4097d5dc, 32'h41a67d44} /* (23, 10, 22) {real, imag} */,
  {32'h41af6d94, 32'hc17485d4} /* (23, 10, 21) {real, imag} */,
  {32'h4151e7ae, 32'h4119f0c2} /* (23, 10, 20) {real, imag} */,
  {32'hc0e8db5a, 32'h41d9b0aa} /* (23, 10, 19) {real, imag} */,
  {32'h3f0c7d58, 32'h40e11c30} /* (23, 10, 18) {real, imag} */,
  {32'hc0535690, 32'hc04a9ef2} /* (23, 10, 17) {real, imag} */,
  {32'h3d9e0a80, 32'hc1526b2a} /* (23, 10, 16) {real, imag} */,
  {32'h3dfa3400, 32'h3d7b3380} /* (23, 10, 15) {real, imag} */,
  {32'hc0bd1df5, 32'hc0143d50} /* (23, 10, 14) {real, imag} */,
  {32'hbfcc1528, 32'h417807f5} /* (23, 10, 13) {real, imag} */,
  {32'h41e1d95d, 32'h41638b8e} /* (23, 10, 12) {real, imag} */,
  {32'hc1139b3d, 32'h3f89aa30} /* (23, 10, 11) {real, imag} */,
  {32'h410a8986, 32'h41050fb4} /* (23, 10, 10) {real, imag} */,
  {32'h4100b895, 32'h41b00aef} /* (23, 10, 9) {real, imag} */,
  {32'hc1c93ca8, 32'hc1952110} /* (23, 10, 8) {real, imag} */,
  {32'hc26fc683, 32'hc1da2904} /* (23, 10, 7) {real, imag} */,
  {32'h4215b7fd, 32'h40003790} /* (23, 10, 6) {real, imag} */,
  {32'h411481fe, 32'hc1c02307} /* (23, 10, 5) {real, imag} */,
  {32'h409c52af, 32'hc23dc0b0} /* (23, 10, 4) {real, imag} */,
  {32'hc1b9063e, 32'hc15b38b4} /* (23, 10, 3) {real, imag} */,
  {32'hc0a98903, 32'h429ac105} /* (23, 10, 2) {real, imag} */,
  {32'hc207c805, 32'hc26171aa} /* (23, 10, 1) {real, imag} */,
  {32'h41584c6d, 32'hc0439240} /* (23, 10, 0) {real, imag} */,
  {32'h41896506, 32'hc25ed6c7} /* (23, 9, 31) {real, imag} */,
  {32'hc1804e2e, 32'h4129b279} /* (23, 9, 30) {real, imag} */,
  {32'h40da646c, 32'h419ba2f1} /* (23, 9, 29) {real, imag} */,
  {32'hc1d98cea, 32'hc2a87f9f} /* (23, 9, 28) {real, imag} */,
  {32'h420fa1be, 32'hc1c0e679} /* (23, 9, 27) {real, imag} */,
  {32'h420e8eec, 32'hc14878bd} /* (23, 9, 26) {real, imag} */,
  {32'h401774f8, 32'h416d368f} /* (23, 9, 25) {real, imag} */,
  {32'h42ae1668, 32'h4130215c} /* (23, 9, 24) {real, imag} */,
  {32'hc1e66fbc, 32'hc0b24b42} /* (23, 9, 23) {real, imag} */,
  {32'hc1a035f8, 32'hc1aa2ca9} /* (23, 9, 22) {real, imag} */,
  {32'hc15fabc2, 32'hc125ea26} /* (23, 9, 21) {real, imag} */,
  {32'hc1846c5b, 32'hc0072c30} /* (23, 9, 20) {real, imag} */,
  {32'h418b40fc, 32'h4110d9fd} /* (23, 9, 19) {real, imag} */,
  {32'hc123a95f, 32'hc056159c} /* (23, 9, 18) {real, imag} */,
  {32'hc0c2bd34, 32'h40875402} /* (23, 9, 17) {real, imag} */,
  {32'h40537136, 32'hc0283700} /* (23, 9, 16) {real, imag} */,
  {32'h4168d9b4, 32'h4022f664} /* (23, 9, 15) {real, imag} */,
  {32'hc11e367b, 32'hc05ca37c} /* (23, 9, 14) {real, imag} */,
  {32'hc187e1c0, 32'hc10d92eb} /* (23, 9, 13) {real, imag} */,
  {32'h414f1cb0, 32'h416b9818} /* (23, 9, 12) {real, imag} */,
  {32'hc1b13a2f, 32'hc1064b56} /* (23, 9, 11) {real, imag} */,
  {32'hc140e380, 32'h4149942e} /* (23, 9, 10) {real, imag} */,
  {32'hc18fb27e, 32'hbfae95c8} /* (23, 9, 9) {real, imag} */,
  {32'hc12a89d4, 32'h4117fb64} /* (23, 9, 8) {real, imag} */,
  {32'hc1f57ead, 32'hc1b32fca} /* (23, 9, 7) {real, imag} */,
  {32'h4191aad7, 32'hc22c126c} /* (23, 9, 6) {real, imag} */,
  {32'hc1b79975, 32'h3f002d20} /* (23, 9, 5) {real, imag} */,
  {32'h41ba2ea2, 32'hc1a89343} /* (23, 9, 4) {real, imag} */,
  {32'hc0afcd94, 32'h419c62c7} /* (23, 9, 3) {real, imag} */,
  {32'h41a955e4, 32'h411cbd25} /* (23, 9, 2) {real, imag} */,
  {32'hc2817d8c, 32'h42d67fe4} /* (23, 9, 1) {real, imag} */,
  {32'h41561a1a, 32'hc12896bc} /* (23, 9, 0) {real, imag} */,
  {32'h419f753d, 32'h411ada96} /* (23, 8, 31) {real, imag} */,
  {32'hc127df2d, 32'hc25fd60e} /* (23, 8, 30) {real, imag} */,
  {32'hc1422650, 32'h4176c234} /* (23, 8, 29) {real, imag} */,
  {32'h42944bc0, 32'h418f0918} /* (23, 8, 28) {real, imag} */,
  {32'h40f6cb00, 32'hc274442c} /* (23, 8, 27) {real, imag} */,
  {32'hc0b9a308, 32'hc0959c34} /* (23, 8, 26) {real, imag} */,
  {32'hc0ac1214, 32'hc19dc482} /* (23, 8, 25) {real, imag} */,
  {32'hc1ca3229, 32'hc214720e} /* (23, 8, 24) {real, imag} */,
  {32'h4196581e, 32'hc1be7578} /* (23, 8, 23) {real, imag} */,
  {32'h4217218c, 32'h4097cbc4} /* (23, 8, 22) {real, imag} */,
  {32'hbf01d208, 32'h421a2a87} /* (23, 8, 21) {real, imag} */,
  {32'hbec2fa80, 32'h420186a9} /* (23, 8, 20) {real, imag} */,
  {32'h4173f5d9, 32'hc20dee07} /* (23, 8, 19) {real, imag} */,
  {32'h415d27e3, 32'hc0f0bbe5} /* (23, 8, 18) {real, imag} */,
  {32'hc0c591c4, 32'h419d7acc} /* (23, 8, 17) {real, imag} */,
  {32'hc0a8835a, 32'hc1a308c4} /* (23, 8, 16) {real, imag} */,
  {32'hc0abe648, 32'h3e270140} /* (23, 8, 15) {real, imag} */,
  {32'h41cd3cfc, 32'h4088d2f5} /* (23, 8, 14) {real, imag} */,
  {32'h4117afbf, 32'hc1218854} /* (23, 8, 13) {real, imag} */,
  {32'hc00430d0, 32'hc1e3e972} /* (23, 8, 12) {real, imag} */,
  {32'h3fd46964, 32'h40d906a8} /* (23, 8, 11) {real, imag} */,
  {32'h40a643f4, 32'h41eb8c39} /* (23, 8, 10) {real, imag} */,
  {32'hc16aac29, 32'h413035b3} /* (23, 8, 9) {real, imag} */,
  {32'h42334e18, 32'h411cbf17} /* (23, 8, 8) {real, imag} */,
  {32'hc1e92e5b, 32'hc2269939} /* (23, 8, 7) {real, imag} */,
  {32'hc20ab70c, 32'h4215abe6} /* (23, 8, 6) {real, imag} */,
  {32'h4204a51f, 32'h429c4b86} /* (23, 8, 5) {real, imag} */,
  {32'hc1b2230e, 32'hc21bccf0} /* (23, 8, 4) {real, imag} */,
  {32'hc1b1ee86, 32'h41c9a136} /* (23, 8, 3) {real, imag} */,
  {32'hc222355e, 32'hc1f744f7} /* (23, 8, 2) {real, imag} */,
  {32'h401d9460, 32'hc2774e02} /* (23, 8, 1) {real, imag} */,
  {32'hc1b74118, 32'h428d3099} /* (23, 8, 0) {real, imag} */,
  {32'h420e93eb, 32'hc2fc37da} /* (23, 7, 31) {real, imag} */,
  {32'h4151a897, 32'h420e3306} /* (23, 7, 30) {real, imag} */,
  {32'h4222a6e3, 32'h422e5377} /* (23, 7, 29) {real, imag} */,
  {32'h41e4cb45, 32'h41d3a276} /* (23, 7, 28) {real, imag} */,
  {32'h42c73e97, 32'h43060a73} /* (23, 7, 27) {real, imag} */,
  {32'hc274880a, 32'hc0488638} /* (23, 7, 26) {real, imag} */,
  {32'h417b99c5, 32'hc1e70f30} /* (23, 7, 25) {real, imag} */,
  {32'h42142acb, 32'hc2029231} /* (23, 7, 24) {real, imag} */,
  {32'hc1e263cc, 32'hc1cfab30} /* (23, 7, 23) {real, imag} */,
  {32'hc23d3774, 32'hc1f7bc75} /* (23, 7, 22) {real, imag} */,
  {32'hc1bc3ea0, 32'h40a94338} /* (23, 7, 21) {real, imag} */,
  {32'hc10ec02d, 32'h40e445ce} /* (23, 7, 20) {real, imag} */,
  {32'h4076ff5c, 32'h4179881f} /* (23, 7, 19) {real, imag} */,
  {32'h4091f086, 32'h41527b75} /* (23, 7, 18) {real, imag} */,
  {32'hc11cf8c6, 32'hc0590510} /* (23, 7, 17) {real, imag} */,
  {32'h4115631f, 32'h4156cf10} /* (23, 7, 16) {real, imag} */,
  {32'h419c9b71, 32'hc161d864} /* (23, 7, 15) {real, imag} */,
  {32'h417ad4a5, 32'hc0bd5cea} /* (23, 7, 14) {real, imag} */,
  {32'hc174df8f, 32'h41e34990} /* (23, 7, 13) {real, imag} */,
  {32'hbe430440, 32'hbfa0e1b8} /* (23, 7, 12) {real, imag} */,
  {32'hc1e92366, 32'h4202910d} /* (23, 7, 11) {real, imag} */,
  {32'hc21494bc, 32'hc22e675b} /* (23, 7, 10) {real, imag} */,
  {32'hc1fd45c4, 32'hc0a96c0c} /* (23, 7, 9) {real, imag} */,
  {32'h41f76c67, 32'h415be764} /* (23, 7, 8) {real, imag} */,
  {32'hc1898508, 32'hc1451207} /* (23, 7, 7) {real, imag} */,
  {32'hc27aea9e, 32'hc1d729d5} /* (23, 7, 6) {real, imag} */,
  {32'hc1f17a9c, 32'hc27a9bed} /* (23, 7, 5) {real, imag} */,
  {32'h41b0b21b, 32'hc1c4bdae} /* (23, 7, 4) {real, imag} */,
  {32'hbfe3eca0, 32'hc09f1168} /* (23, 7, 3) {real, imag} */,
  {32'h40b6ee62, 32'h42a65d63} /* (23, 7, 2) {real, imag} */,
  {32'h4238df59, 32'h41f28f0a} /* (23, 7, 1) {real, imag} */,
  {32'h41ba8fbc, 32'h416b8268} /* (23, 7, 0) {real, imag} */,
  {32'h429cd4a9, 32'hc18aa8a5} /* (23, 6, 31) {real, imag} */,
  {32'hc1d49b7a, 32'hc10900cd} /* (23, 6, 30) {real, imag} */,
  {32'hc29d4b2a, 32'h41050ea0} /* (23, 6, 29) {real, imag} */,
  {32'h4244bedd, 32'hc295fc38} /* (23, 6, 28) {real, imag} */,
  {32'hc2acda34, 32'hc167050c} /* (23, 6, 27) {real, imag} */,
  {32'hc2457413, 32'hc24cb13d} /* (23, 6, 26) {real, imag} */,
  {32'h413a48a1, 32'hc23aac26} /* (23, 6, 25) {real, imag} */,
  {32'hc132708e, 32'h42537f5c} /* (23, 6, 24) {real, imag} */,
  {32'h41c3e03c, 32'hbe65cc80} /* (23, 6, 23) {real, imag} */,
  {32'hc261d9f6, 32'h429c26ea} /* (23, 6, 22) {real, imag} */,
  {32'h4121f25b, 32'hc1ef0a9d} /* (23, 6, 21) {real, imag} */,
  {32'h418d2b6c, 32'hc16e98c2} /* (23, 6, 20) {real, imag} */,
  {32'hc0c3dcb1, 32'hc016b080} /* (23, 6, 19) {real, imag} */,
  {32'hc067b2b8, 32'h410f7c81} /* (23, 6, 18) {real, imag} */,
  {32'h42291546, 32'h4190718a} /* (23, 6, 17) {real, imag} */,
  {32'hc14d876c, 32'h4192b09b} /* (23, 6, 16) {real, imag} */,
  {32'hc194cc24, 32'hc008f960} /* (23, 6, 15) {real, imag} */,
  {32'hc1e2b7f6, 32'h41bc3aee} /* (23, 6, 14) {real, imag} */,
  {32'hc10a3200, 32'h4114eaa0} /* (23, 6, 13) {real, imag} */,
  {32'hc1a535cc, 32'h4214447c} /* (23, 6, 12) {real, imag} */,
  {32'h408047da, 32'hc25b990e} /* (23, 6, 11) {real, imag} */,
  {32'hbfedfa40, 32'h4206ee77} /* (23, 6, 10) {real, imag} */,
  {32'h423a447e, 32'hc202dee4} /* (23, 6, 9) {real, imag} */,
  {32'hc0f4738b, 32'hc1dc300c} /* (23, 6, 8) {real, imag} */,
  {32'h41ca9ac0, 32'h3f2f08e0} /* (23, 6, 7) {real, imag} */,
  {32'h413e39fc, 32'h41ca9e8a} /* (23, 6, 6) {real, imag} */,
  {32'hc207552e, 32'hc178966e} /* (23, 6, 5) {real, imag} */,
  {32'h426da83f, 32'hc09fc298} /* (23, 6, 4) {real, imag} */,
  {32'h425fd3d3, 32'h432b0b6c} /* (23, 6, 3) {real, imag} */,
  {32'h4240d117, 32'h41acd8a0} /* (23, 6, 2) {real, imag} */,
  {32'hc28b4a7f, 32'h429ad133} /* (23, 6, 1) {real, imag} */,
  {32'hc2620ed5, 32'h411a268a} /* (23, 6, 0) {real, imag} */,
  {32'hc205c89f, 32'h422553df} /* (23, 5, 31) {real, imag} */,
  {32'h42523c29, 32'hc25cb15e} /* (23, 5, 30) {real, imag} */,
  {32'hc2a61a4c, 32'hc2265f88} /* (23, 5, 29) {real, imag} */,
  {32'hc11acf14, 32'h41a5c4a0} /* (23, 5, 28) {real, imag} */,
  {32'h3f260630, 32'hc271aef8} /* (23, 5, 27) {real, imag} */,
  {32'hc20e5be2, 32'hc290934e} /* (23, 5, 26) {real, imag} */,
  {32'h424d2168, 32'hc074fbc0} /* (23, 5, 25) {real, imag} */,
  {32'h42867532, 32'hc27392d0} /* (23, 5, 24) {real, imag} */,
  {32'h42516011, 32'hc273fa24} /* (23, 5, 23) {real, imag} */,
  {32'h41dc9e16, 32'h4281f12e} /* (23, 5, 22) {real, imag} */,
  {32'hc1de654c, 32'h4102f82a} /* (23, 5, 21) {real, imag} */,
  {32'h416c8cfc, 32'h40b685d0} /* (23, 5, 20) {real, imag} */,
  {32'hc0dc147e, 32'h4166eed8} /* (23, 5, 19) {real, imag} */,
  {32'hc1af1419, 32'h41d3205e} /* (23, 5, 18) {real, imag} */,
  {32'hbf549db0, 32'hc003b604} /* (23, 5, 17) {real, imag} */,
  {32'hc17f35eb, 32'hc17165fe} /* (23, 5, 16) {real, imag} */,
  {32'h413e5e1d, 32'h419bd404} /* (23, 5, 15) {real, imag} */,
  {32'h3fdb8850, 32'h412cdda3} /* (23, 5, 14) {real, imag} */,
  {32'h3f9a2d08, 32'hc144e99c} /* (23, 5, 13) {real, imag} */,
  {32'hc2526363, 32'h3f559440} /* (23, 5, 12) {real, imag} */,
  {32'h408ce71e, 32'hc20f20f2} /* (23, 5, 11) {real, imag} */,
  {32'h3f756680, 32'hc28bef4e} /* (23, 5, 10) {real, imag} */,
  {32'hc1d8141e, 32'hc28ca65a} /* (23, 5, 9) {real, imag} */,
  {32'hc19a9cc2, 32'h42605998} /* (23, 5, 8) {real, imag} */,
  {32'h424375ae, 32'h42b5b906} /* (23, 5, 7) {real, imag} */,
  {32'hc24fd236, 32'hc298151e} /* (23, 5, 6) {real, imag} */,
  {32'h41e1306a, 32'hc0d28e80} /* (23, 5, 5) {real, imag} */,
  {32'h418d1405, 32'h422f6dd0} /* (23, 5, 4) {real, imag} */,
  {32'h428ba640, 32'h41e0bbe1} /* (23, 5, 3) {real, imag} */,
  {32'hc27767c7, 32'hc2510766} /* (23, 5, 2) {real, imag} */,
  {32'h427c5bfb, 32'h42df11c0} /* (23, 5, 1) {real, imag} */,
  {32'h41c49a8a, 32'hc21526b2} /* (23, 5, 0) {real, imag} */,
  {32'h42582a12, 32'hc2bd85e2} /* (23, 4, 31) {real, imag} */,
  {32'hc23844d0, 32'h42ae619e} /* (23, 4, 30) {real, imag} */,
  {32'hc2742c4a, 32'hc27d5122} /* (23, 4, 29) {real, imag} */,
  {32'hc20f1f26, 32'hc1196e5a} /* (23, 4, 28) {real, imag} */,
  {32'hc1fc8599, 32'h424b4a80} /* (23, 4, 27) {real, imag} */,
  {32'h4208835b, 32'hc1b7617a} /* (23, 4, 26) {real, imag} */,
  {32'h41a0c7ae, 32'h420a5c70} /* (23, 4, 25) {real, imag} */,
  {32'hc304deb0, 32'h4218e6e6} /* (23, 4, 24) {real, imag} */,
  {32'hc20ac39b, 32'hc16ad67a} /* (23, 4, 23) {real, imag} */,
  {32'hc19a51f2, 32'h41ffcc8e} /* (23, 4, 22) {real, imag} */,
  {32'hc164e8c8, 32'hc19b3af6} /* (23, 4, 21) {real, imag} */,
  {32'hc0a29bb0, 32'h40f51f9a} /* (23, 4, 20) {real, imag} */,
  {32'hc196aa4f, 32'h41b40a83} /* (23, 4, 19) {real, imag} */,
  {32'h41b1b88f, 32'hc2226179} /* (23, 4, 18) {real, imag} */,
  {32'h40813c8c, 32'h4192ebea} /* (23, 4, 17) {real, imag} */,
  {32'h41991eff, 32'hc1a9d768} /* (23, 4, 16) {real, imag} */,
  {32'hc17fb606, 32'h402386ec} /* (23, 4, 15) {real, imag} */,
  {32'hc13ff77a, 32'hc1d4d552} /* (23, 4, 14) {real, imag} */,
  {32'hc1b527e3, 32'hc1c6e0fd} /* (23, 4, 13) {real, imag} */,
  {32'h42346868, 32'hc2074013} /* (23, 4, 12) {real, imag} */,
  {32'h400708a0, 32'h41b3a2a6} /* (23, 4, 11) {real, imag} */,
  {32'h4203b9d1, 32'hc0fddc6e} /* (23, 4, 10) {real, imag} */,
  {32'h420194c1, 32'hc1ff9d9f} /* (23, 4, 9) {real, imag} */,
  {32'h4292f3e4, 32'h422cfaea} /* (23, 4, 8) {real, imag} */,
  {32'hc18fcb9a, 32'h4236a9d8} /* (23, 4, 7) {real, imag} */,
  {32'h4295df94, 32'h42acf1ce} /* (23, 4, 6) {real, imag} */,
  {32'h42817acf, 32'h427d665e} /* (23, 4, 5) {real, imag} */,
  {32'h42647b98, 32'h40bc3ff1} /* (23, 4, 4) {real, imag} */,
  {32'hc1638728, 32'hc28485cf} /* (23, 4, 3) {real, imag} */,
  {32'hc234dc7c, 32'hc1f2b2f2} /* (23, 4, 2) {real, imag} */,
  {32'h42098e24, 32'h424547c5} /* (23, 4, 1) {real, imag} */,
  {32'h41d3be15, 32'h42bd329e} /* (23, 4, 0) {real, imag} */,
  {32'hbf4a4b60, 32'h4301f7fe} /* (23, 3, 31) {real, imag} */,
  {32'hc30ac511, 32'h42abc953} /* (23, 3, 30) {real, imag} */,
  {32'hc0704160, 32'hc1d15350} /* (23, 3, 29) {real, imag} */,
  {32'hc295da43, 32'hc1cf1944} /* (23, 3, 28) {real, imag} */,
  {32'h42a164ca, 32'hc278c792} /* (23, 3, 27) {real, imag} */,
  {32'h412d0660, 32'hc222108c} /* (23, 3, 26) {real, imag} */,
  {32'hc1950382, 32'hc1c236f0} /* (23, 3, 25) {real, imag} */,
  {32'h42432f63, 32'h4255b97a} /* (23, 3, 24) {real, imag} */,
  {32'hc15276d8, 32'h41aab8d0} /* (23, 3, 23) {real, imag} */,
  {32'h427a3226, 32'hc13ee1d4} /* (23, 3, 22) {real, imag} */,
  {32'hc18f22a8, 32'hc0426710} /* (23, 3, 21) {real, imag} */,
  {32'h41c11508, 32'h41fedbde} /* (23, 3, 20) {real, imag} */,
  {32'h4111c3b8, 32'hc20407f6} /* (23, 3, 19) {real, imag} */,
  {32'h41573b70, 32'hc0c7b9f8} /* (23, 3, 18) {real, imag} */,
  {32'hc1e173a6, 32'h416347eb} /* (23, 3, 17) {real, imag} */,
  {32'hc10dc17e, 32'h404eb928} /* (23, 3, 16) {real, imag} */,
  {32'hc0a12c06, 32'hc11e077d} /* (23, 3, 15) {real, imag} */,
  {32'h4111b210, 32'hc1881cc2} /* (23, 3, 14) {real, imag} */,
  {32'hc1a27a06, 32'h419a514b} /* (23, 3, 13) {real, imag} */,
  {32'hc1fe5622, 32'h426bf5b3} /* (23, 3, 12) {real, imag} */,
  {32'hc1f77378, 32'hc2237a8a} /* (23, 3, 11) {real, imag} */,
  {32'h421dabb0, 32'h42031102} /* (23, 3, 10) {real, imag} */,
  {32'h41c20fe0, 32'hc1f1319c} /* (23, 3, 9) {real, imag} */,
  {32'hbea71100, 32'hc24d8860} /* (23, 3, 8) {real, imag} */,
  {32'h41f9445e, 32'hc1c7b67a} /* (23, 3, 7) {real, imag} */,
  {32'hc1ca6950, 32'hc1d2a9df} /* (23, 3, 6) {real, imag} */,
  {32'h41f901c2, 32'hc28806d3} /* (23, 3, 5) {real, imag} */,
  {32'h4041aee0, 32'hc22d37e0} /* (23, 3, 4) {real, imag} */,
  {32'h42a3012b, 32'hc28e1ba2} /* (23, 3, 3) {real, imag} */,
  {32'hc309f91f, 32'h4308ffa8} /* (23, 3, 2) {real, imag} */,
  {32'hc1298a58, 32'hc2c21fb0} /* (23, 3, 1) {real, imag} */,
  {32'hc01d2918, 32'hc2862053} /* (23, 3, 0) {real, imag} */,
  {32'h42fc1e3c, 32'h42962f98} /* (23, 2, 31) {real, imag} */,
  {32'hc2c55f78, 32'hc2b5bc6b} /* (23, 2, 30) {real, imag} */,
  {32'hc3099638, 32'hc2767b21} /* (23, 2, 29) {real, imag} */,
  {32'h42a41a1d, 32'hbf437b00} /* (23, 2, 28) {real, imag} */,
  {32'hc13eecd8, 32'h4234bad5} /* (23, 2, 27) {real, imag} */,
  {32'hc2f5b0e2, 32'hc266f61e} /* (23, 2, 26) {real, imag} */,
  {32'h40e4e350, 32'h42c26268} /* (23, 2, 25) {real, imag} */,
  {32'hc21cb670, 32'h425f9877} /* (23, 2, 24) {real, imag} */,
  {32'h41388534, 32'hc1ea9f48} /* (23, 2, 23) {real, imag} */,
  {32'h41e8bd14, 32'h42682623} /* (23, 2, 22) {real, imag} */,
  {32'hc127b754, 32'hc28e8c93} /* (23, 2, 21) {real, imag} */,
  {32'hc0302072, 32'hc2277e64} /* (23, 2, 20) {real, imag} */,
  {32'h4206c354, 32'hc029dea0} /* (23, 2, 19) {real, imag} */,
  {32'hc0d3844a, 32'h42039ad6} /* (23, 2, 18) {real, imag} */,
  {32'h404f5e02, 32'h41a9baac} /* (23, 2, 17) {real, imag} */,
  {32'hc152d690, 32'h40272ce0} /* (23, 2, 16) {real, imag} */,
  {32'h414786f0, 32'hc0f5cf9e} /* (23, 2, 15) {real, imag} */,
  {32'hc11342fb, 32'h410bc6aa} /* (23, 2, 14) {real, imag} */,
  {32'hc1cd3cb1, 32'h41f8d4f4} /* (23, 2, 13) {real, imag} */,
  {32'h40439c0e, 32'hc1e76a44} /* (23, 2, 12) {real, imag} */,
  {32'h415266f8, 32'hc24ce4ab} /* (23, 2, 11) {real, imag} */,
  {32'hc20e0b4e, 32'hc2190e6d} /* (23, 2, 10) {real, imag} */,
  {32'h420aeae9, 32'hc1dfe238} /* (23, 2, 9) {real, imag} */,
  {32'h4208df36, 32'hc2df697e} /* (23, 2, 8) {real, imag} */,
  {32'h4284728f, 32'h41e1f310} /* (23, 2, 7) {real, imag} */,
  {32'hc1af9100, 32'h4207bf7a} /* (23, 2, 6) {real, imag} */,
  {32'hc093b398, 32'h42a75582} /* (23, 2, 5) {real, imag} */,
  {32'hc254e96e, 32'h4241d9e8} /* (23, 2, 4) {real, imag} */,
  {32'h42105d86, 32'h42bf6642} /* (23, 2, 3) {real, imag} */,
  {32'hc250f278, 32'hc324d56e} /* (23, 2, 2) {real, imag} */,
  {32'h42f3d57e, 32'hc286c258} /* (23, 2, 1) {real, imag} */,
  {32'hc037fa00, 32'h4281ba82} /* (23, 2, 0) {real, imag} */,
  {32'hc299a83f, 32'hc2d759fd} /* (23, 1, 31) {real, imag} */,
  {32'hc1451a0e, 32'hc1ea00a4} /* (23, 1, 30) {real, imag} */,
  {32'h4296f5ba, 32'hc28661b8} /* (23, 1, 29) {real, imag} */,
  {32'hc2401b68, 32'hc22333b4} /* (23, 1, 28) {real, imag} */,
  {32'h420ffc79, 32'h422be735} /* (23, 1, 27) {real, imag} */,
  {32'h415fa245, 32'h401c27a2} /* (23, 1, 26) {real, imag} */,
  {32'h421c709c, 32'hc22f771b} /* (23, 1, 25) {real, imag} */,
  {32'hc1e558d0, 32'h41fe7ffa} /* (23, 1, 24) {real, imag} */,
  {32'h41ad5490, 32'h422b3e9d} /* (23, 1, 23) {real, imag} */,
  {32'h413dd2f2, 32'hc0968f54} /* (23, 1, 22) {real, imag} */,
  {32'h427244b4, 32'hc1947a1c} /* (23, 1, 21) {real, imag} */,
  {32'h421eb594, 32'hc0ac53c0} /* (23, 1, 20) {real, imag} */,
  {32'hc1c834fa, 32'h41b04af7} /* (23, 1, 19) {real, imag} */,
  {32'h41918874, 32'h415d5948} /* (23, 1, 18) {real, imag} */,
  {32'h41d88b71, 32'h41ecb20c} /* (23, 1, 17) {real, imag} */,
  {32'h4202f15a, 32'hc1b1b744} /* (23, 1, 16) {real, imag} */,
  {32'hbea6cb40, 32'h40dcfdd2} /* (23, 1, 15) {real, imag} */,
  {32'hc218a56d, 32'h41c1dc4c} /* (23, 1, 14) {real, imag} */,
  {32'hc148344c, 32'hc11e3da2} /* (23, 1, 13) {real, imag} */,
  {32'h4128a015, 32'h4200716d} /* (23, 1, 12) {real, imag} */,
  {32'h4224faaa, 32'h42148a3c} /* (23, 1, 11) {real, imag} */,
  {32'hc18f1224, 32'hc210b36e} /* (23, 1, 10) {real, imag} */,
  {32'hc1695080, 32'hc291e97a} /* (23, 1, 9) {real, imag} */,
  {32'hc1d997c0, 32'h42b4196a} /* (23, 1, 8) {real, imag} */,
  {32'h42528544, 32'h41a4c572} /* (23, 1, 7) {real, imag} */,
  {32'hc2010847, 32'hc1837184} /* (23, 1, 6) {real, imag} */,
  {32'h42359c51, 32'hc18d106a} /* (23, 1, 5) {real, imag} */,
  {32'hc1988370, 32'hc296735c} /* (23, 1, 4) {real, imag} */,
  {32'hc224c513, 32'hc1111df0} /* (23, 1, 3) {real, imag} */,
  {32'hc1b55b5d, 32'h42f72f4d} /* (23, 1, 2) {real, imag} */,
  {32'hc2b98911, 32'hc338a2fc} /* (23, 1, 1) {real, imag} */,
  {32'hc3016198, 32'hc3068ac2} /* (23, 1, 0) {real, imag} */,
  {32'hc307a91e, 32'h4283d1b6} /* (23, 0, 31) {real, imag} */,
  {32'hc26499ea, 32'h4167d9aa} /* (23, 0, 30) {real, imag} */,
  {32'h4319e11e, 32'h416bf247} /* (23, 0, 29) {real, imag} */,
  {32'hc2958a7d, 32'hc2815db2} /* (23, 0, 28) {real, imag} */,
  {32'h4284656e, 32'h422cb3f0} /* (23, 0, 27) {real, imag} */,
  {32'hc17ece3e, 32'h428f13c2} /* (23, 0, 26) {real, imag} */,
  {32'hc2345e58, 32'hc24c003a} /* (23, 0, 25) {real, imag} */,
  {32'h42a7e8cd, 32'hc30b6576} /* (23, 0, 24) {real, imag} */,
  {32'h41eadff5, 32'h40c4b7e8} /* (23, 0, 23) {real, imag} */,
  {32'hc1f0ff1a, 32'hc225af46} /* (23, 0, 22) {real, imag} */,
  {32'hc16be6fc, 32'h422f80c8} /* (23, 0, 21) {real, imag} */,
  {32'h40c1776f, 32'hc18c4a10} /* (23, 0, 20) {real, imag} */,
  {32'hc1e9a5e6, 32'hc123d985} /* (23, 0, 19) {real, imag} */,
  {32'h419b6748, 32'hc1d51116} /* (23, 0, 18) {real, imag} */,
  {32'hc0702b48, 32'h41252876} /* (23, 0, 17) {real, imag} */,
  {32'h40f3aeca, 32'h41c0dff0} /* (23, 0, 16) {real, imag} */,
  {32'hc104a436, 32'hc102a1ea} /* (23, 0, 15) {real, imag} */,
  {32'hc19f61b8, 32'h416cabd1} /* (23, 0, 14) {real, imag} */,
  {32'h421a8a1d, 32'h411a283b} /* (23, 0, 13) {real, imag} */,
  {32'h402ca36e, 32'h3f308b70} /* (23, 0, 12) {real, imag} */,
  {32'hc19f471a, 32'hc03dedf8} /* (23, 0, 11) {real, imag} */,
  {32'h42bb3720, 32'h418d606c} /* (23, 0, 10) {real, imag} */,
  {32'h41a55593, 32'h427ca8b9} /* (23, 0, 9) {real, imag} */,
  {32'hc298721b, 32'h42aa85a8} /* (23, 0, 8) {real, imag} */,
  {32'h4178c072, 32'hc203b7f8} /* (23, 0, 7) {real, imag} */,
  {32'hc28c67e7, 32'hc181a3d8} /* (23, 0, 6) {real, imag} */,
  {32'h424a25c1, 32'h4106bafe} /* (23, 0, 5) {real, imag} */,
  {32'h424e5482, 32'hc11d796c} /* (23, 0, 4) {real, imag} */,
  {32'hc29bfccc, 32'hc18a9164} /* (23, 0, 3) {real, imag} */,
  {32'h41fae6d4, 32'h41d20c4b} /* (23, 0, 2) {real, imag} */,
  {32'hc27b2318, 32'hc2e71cb2} /* (23, 0, 1) {real, imag} */,
  {32'hc1a5d9aa, 32'hc3401eb6} /* (23, 0, 0) {real, imag} */,
  {32'hc32ee7ef, 32'h425cd792} /* (22, 31, 31) {real, imag} */,
  {32'h42063bea, 32'h42845d5a} /* (22, 31, 30) {real, imag} */,
  {32'h425bbeb0, 32'hc2a0d075} /* (22, 31, 29) {real, imag} */,
  {32'hc20cb128, 32'hc21011a8} /* (22, 31, 28) {real, imag} */,
  {32'h41292ca4, 32'h419961af} /* (22, 31, 27) {real, imag} */,
  {32'h4202f16f, 32'hc22a7e2a} /* (22, 31, 26) {real, imag} */,
  {32'h41fb7ca8, 32'hc1a43b1d} /* (22, 31, 25) {real, imag} */,
  {32'hc212ba7a, 32'hc07286e8} /* (22, 31, 24) {real, imag} */,
  {32'h42272078, 32'hc19bdeed} /* (22, 31, 23) {real, imag} */,
  {32'h3f630180, 32'hc0d64d64} /* (22, 31, 22) {real, imag} */,
  {32'h41dfce59, 32'hc248a61c} /* (22, 31, 21) {real, imag} */,
  {32'hc1952741, 32'hc02faa60} /* (22, 31, 20) {real, imag} */,
  {32'hc120e439, 32'hbe77fe00} /* (22, 31, 19) {real, imag} */,
  {32'h40945a9c, 32'hc2369011} /* (22, 31, 18) {real, imag} */,
  {32'h3f0443e0, 32'h41dbb071} /* (22, 31, 17) {real, imag} */,
  {32'hc1ac4fe1, 32'hc1c6cf6f} /* (22, 31, 16) {real, imag} */,
  {32'hc1c98537, 32'h403372d8} /* (22, 31, 15) {real, imag} */,
  {32'hc00ba8f8, 32'h40a37fa0} /* (22, 31, 14) {real, imag} */,
  {32'h4187be62, 32'h3fb1ab40} /* (22, 31, 13) {real, imag} */,
  {32'h41870ba9, 32'hc19b1774} /* (22, 31, 12) {real, imag} */,
  {32'h42453da6, 32'h412022c2} /* (22, 31, 11) {real, imag} */,
  {32'hc245066e, 32'hc1c11247} /* (22, 31, 10) {real, imag} */,
  {32'hc0bbaa04, 32'hc2049170} /* (22, 31, 9) {real, imag} */,
  {32'h404d7658, 32'h40fb3b14} /* (22, 31, 8) {real, imag} */,
  {32'h4142e145, 32'h4199d975} /* (22, 31, 7) {real, imag} */,
  {32'h42cda2d8, 32'hc2c31b7f} /* (22, 31, 6) {real, imag} */,
  {32'h42afb88a, 32'h424c9250} /* (22, 31, 5) {real, imag} */,
  {32'hc1e5c135, 32'hc2f88542} /* (22, 31, 4) {real, imag} */,
  {32'h41ded948, 32'h4251b74e} /* (22, 31, 3) {real, imag} */,
  {32'h42a62adb, 32'hc1a17841} /* (22, 31, 2) {real, imag} */,
  {32'hc2e15702, 32'hc28210a5} /* (22, 31, 1) {real, imag} */,
  {32'hc27fd99a, 32'hc241afb0} /* (22, 31, 0) {real, imag} */,
  {32'h429dd48d, 32'h40a49e18} /* (22, 30, 31) {real, imag} */,
  {32'hc2d83d7a, 32'h3fe02674} /* (22, 30, 30) {real, imag} */,
  {32'hc22eee2d, 32'hc25692bc} /* (22, 30, 29) {real, imag} */,
  {32'h402d23c0, 32'h429c11ae} /* (22, 30, 28) {real, imag} */,
  {32'hc287ec26, 32'hc12e52a3} /* (22, 30, 27) {real, imag} */,
  {32'h42595da2, 32'h414cfa2a} /* (22, 30, 26) {real, imag} */,
  {32'h426c5f0a, 32'h421c05dc} /* (22, 30, 25) {real, imag} */,
  {32'hc227cde4, 32'hc2853e60} /* (22, 30, 24) {real, imag} */,
  {32'hc1ec1908, 32'h41b6d9f9} /* (22, 30, 23) {real, imag} */,
  {32'h418a5051, 32'hc17179ce} /* (22, 30, 22) {real, imag} */,
  {32'h4203aa3c, 32'h42240c60} /* (22, 30, 21) {real, imag} */,
  {32'hc1470be1, 32'h40e097f8} /* (22, 30, 20) {real, imag} */,
  {32'hc0f42418, 32'hc232cb68} /* (22, 30, 19) {real, imag} */,
  {32'hc2164c59, 32'hc18250a2} /* (22, 30, 18) {real, imag} */,
  {32'h420d6406, 32'h41d4abd3} /* (22, 30, 17) {real, imag} */,
  {32'h41c45ad0, 32'h4012a208} /* (22, 30, 16) {real, imag} */,
  {32'hc2135aae, 32'h4053abb8} /* (22, 30, 15) {real, imag} */,
  {32'h419228b6, 32'h41695271} /* (22, 30, 14) {real, imag} */,
  {32'hc1f3e268, 32'hc1ea23e8} /* (22, 30, 13) {real, imag} */,
  {32'hc1dc270c, 32'hc17b77b4} /* (22, 30, 12) {real, imag} */,
  {32'hbf3bf1a0, 32'h40fcda50} /* (22, 30, 11) {real, imag} */,
  {32'h428be256, 32'hc22744c2} /* (22, 30, 10) {real, imag} */,
  {32'hc21b9f4a, 32'h4140a062} /* (22, 30, 9) {real, imag} */,
  {32'h42f50c06, 32'h423b3410} /* (22, 30, 8) {real, imag} */,
  {32'hc0a0d680, 32'h40c991bc} /* (22, 30, 7) {real, imag} */,
  {32'hc1815051, 32'h422b53b0} /* (22, 30, 6) {real, imag} */,
  {32'hc1c36802, 32'hbf025230} /* (22, 30, 5) {real, imag} */,
  {32'h4260ba18, 32'h4250b834} /* (22, 30, 4) {real, imag} */,
  {32'hc2880bba, 32'h42b8b4a8} /* (22, 30, 3) {real, imag} */,
  {32'hc31c4acf, 32'h410cc4e2} /* (22, 30, 2) {real, imag} */,
  {32'h42fdb085, 32'hc156b2fc} /* (22, 30, 1) {real, imag} */,
  {32'h42306348, 32'h41519b82} /* (22, 30, 0) {real, imag} */,
  {32'h41766df0, 32'hc26fb12a} /* (22, 29, 31) {real, imag} */,
  {32'h42cf8d48, 32'hc273ff24} /* (22, 29, 30) {real, imag} */,
  {32'hc20df0be, 32'h4291166f} /* (22, 29, 29) {real, imag} */,
  {32'h41daf23d, 32'h4229383d} /* (22, 29, 28) {real, imag} */,
  {32'h4132e140, 32'hbe056e00} /* (22, 29, 27) {real, imag} */,
  {32'h40eaaf6c, 32'h422adc72} /* (22, 29, 26) {real, imag} */,
  {32'hc07a1098, 32'h4169a76b} /* (22, 29, 25) {real, imag} */,
  {32'h41a9bc7a, 32'h4203e0e4} /* (22, 29, 24) {real, imag} */,
  {32'hc18851f7, 32'h420ff0c3} /* (22, 29, 23) {real, imag} */,
  {32'hc1c328ce, 32'hc1214275} /* (22, 29, 22) {real, imag} */,
  {32'h4186aeaa, 32'h421a3a9c} /* (22, 29, 21) {real, imag} */,
  {32'h40bf46bc, 32'h41226dee} /* (22, 29, 20) {real, imag} */,
  {32'hc16ef024, 32'h41643f9e} /* (22, 29, 19) {real, imag} */,
  {32'hc031f438, 32'hc0d0cf70} /* (22, 29, 18) {real, imag} */,
  {32'h3ff69a60, 32'h410429f8} /* (22, 29, 17) {real, imag} */,
  {32'hc05ce8c8, 32'h41483e6e} /* (22, 29, 16) {real, imag} */,
  {32'hc0bf3e58, 32'hbfd9d1c0} /* (22, 29, 15) {real, imag} */,
  {32'h4102062e, 32'hc1d8a266} /* (22, 29, 14) {real, imag} */,
  {32'h416d8584, 32'hc206ef56} /* (22, 29, 13) {real, imag} */,
  {32'hc22e5db8, 32'hc120ee5a} /* (22, 29, 12) {real, imag} */,
  {32'h40f676fa, 32'hc00f1e20} /* (22, 29, 11) {real, imag} */,
  {32'hc1ce76e4, 32'h41095ebf} /* (22, 29, 10) {real, imag} */,
  {32'hc1b290a9, 32'hc2509d61} /* (22, 29, 9) {real, imag} */,
  {32'h425089a7, 32'hc2a0d266} /* (22, 29, 8) {real, imag} */,
  {32'h4181a697, 32'h408b134e} /* (22, 29, 7) {real, imag} */,
  {32'hc2192c0e, 32'hc280a9d5} /* (22, 29, 6) {real, imag} */,
  {32'h42846ba4, 32'h426412c0} /* (22, 29, 5) {real, imag} */,
  {32'h4021b528, 32'hc210885d} /* (22, 29, 4) {real, imag} */,
  {32'h418168e1, 32'h42a135f5} /* (22, 29, 3) {real, imag} */,
  {32'h4315aa3e, 32'h3f00c4c0} /* (22, 29, 2) {real, imag} */,
  {32'h425c489a, 32'hc274f3e6} /* (22, 29, 1) {real, imag} */,
  {32'hc1cf0577, 32'h411a2d76} /* (22, 29, 0) {real, imag} */,
  {32'hc1f02df7, 32'h4302a482} /* (22, 28, 31) {real, imag} */,
  {32'h42a52cbe, 32'hc2331ebc} /* (22, 28, 30) {real, imag} */,
  {32'hc28a5d15, 32'hc28f5e12} /* (22, 28, 29) {real, imag} */,
  {32'hbfcbe620, 32'h4283a8aa} /* (22, 28, 28) {real, imag} */,
  {32'hc11dce5a, 32'h42233435} /* (22, 28, 27) {real, imag} */,
  {32'hc212f594, 32'hc0bf120c} /* (22, 28, 26) {real, imag} */,
  {32'hc2b29ffe, 32'h422a6db2} /* (22, 28, 25) {real, imag} */,
  {32'hc1af23b5, 32'h41b6c24c} /* (22, 28, 24) {real, imag} */,
  {32'hc07567b8, 32'h425ee684} /* (22, 28, 23) {real, imag} */,
  {32'h415c9dd7, 32'hc19c435b} /* (22, 28, 22) {real, imag} */,
  {32'hc1e66906, 32'hc0c0a350} /* (22, 28, 21) {real, imag} */,
  {32'hc09038dc, 32'hc19a443f} /* (22, 28, 20) {real, imag} */,
  {32'h4162ec06, 32'h4023ece0} /* (22, 28, 19) {real, imag} */,
  {32'h3f87b57c, 32'hc1dad4a3} /* (22, 28, 18) {real, imag} */,
  {32'hc1cf5c5b, 32'hc10a856e} /* (22, 28, 17) {real, imag} */,
  {32'h400677c0, 32'h406d4918} /* (22, 28, 16) {real, imag} */,
  {32'h404a3ba8, 32'h40145cf8} /* (22, 28, 15) {real, imag} */,
  {32'h41377230, 32'hc1d0d431} /* (22, 28, 14) {real, imag} */,
  {32'h4106f94a, 32'h4278084c} /* (22, 28, 13) {real, imag} */,
  {32'hc14dc63a, 32'hc1c8881f} /* (22, 28, 12) {real, imag} */,
  {32'hc007c5b4, 32'h411fc844} /* (22, 28, 11) {real, imag} */,
  {32'hc1d780ca, 32'h426d0258} /* (22, 28, 10) {real, imag} */,
  {32'hc205f828, 32'h422f2b8c} /* (22, 28, 9) {real, imag} */,
  {32'hc1559636, 32'h42b44b79} /* (22, 28, 8) {real, imag} */,
  {32'h41e33702, 32'hc1945709} /* (22, 28, 7) {real, imag} */,
  {32'hc21d7e48, 32'hc239d4a8} /* (22, 28, 6) {real, imag} */,
  {32'h41b9b61d, 32'hc2052c3b} /* (22, 28, 5) {real, imag} */,
  {32'h42e15052, 32'hc18f24e7} /* (22, 28, 4) {real, imag} */,
  {32'hc2b2c24d, 32'hc2b1ba92} /* (22, 28, 3) {real, imag} */,
  {32'h42b6b48c, 32'h40336480} /* (22, 28, 2) {real, imag} */,
  {32'h41454bb2, 32'h40a29f20} /* (22, 28, 1) {real, imag} */,
  {32'hc2b27f32, 32'h41cdc3bd} /* (22, 28, 0) {real, imag} */,
  {32'h42613350, 32'hc2b158f0} /* (22, 27, 31) {real, imag} */,
  {32'h4034d640, 32'h41eeb75a} /* (22, 27, 30) {real, imag} */,
  {32'h418dc034, 32'h41ae18aa} /* (22, 27, 29) {real, imag} */,
  {32'h42278745, 32'h422278bc} /* (22, 27, 28) {real, imag} */,
  {32'hc282dcf7, 32'hc2293198} /* (22, 27, 27) {real, imag} */,
  {32'hc22a8ed5, 32'hc2615dcc} /* (22, 27, 26) {real, imag} */,
  {32'h429a1a78, 32'hc0974130} /* (22, 27, 25) {real, imag} */,
  {32'hc09616fc, 32'h41e5afb7} /* (22, 27, 24) {real, imag} */,
  {32'h41c14280, 32'h3f68b0d0} /* (22, 27, 23) {real, imag} */,
  {32'hc1bd15f4, 32'h4208eb68} /* (22, 27, 22) {real, imag} */,
  {32'hc129e554, 32'hc2080e07} /* (22, 27, 21) {real, imag} */,
  {32'h4125ef1c, 32'hbf0d0ec0} /* (22, 27, 20) {real, imag} */,
  {32'hc1b261f0, 32'h41bc88f6} /* (22, 27, 19) {real, imag} */,
  {32'h41cf8022, 32'h41537bdb} /* (22, 27, 18) {real, imag} */,
  {32'hc1764771, 32'hc11bab2a} /* (22, 27, 17) {real, imag} */,
  {32'hc1445150, 32'h4037fe40} /* (22, 27, 16) {real, imag} */,
  {32'h419371cb, 32'h4019a098} /* (22, 27, 15) {real, imag} */,
  {32'hc0992c3c, 32'h4185e202} /* (22, 27, 14) {real, imag} */,
  {32'hc0a1ddd8, 32'h41855056} /* (22, 27, 13) {real, imag} */,
  {32'hbdf5e500, 32'hc1620f92} /* (22, 27, 12) {real, imag} */,
  {32'h4188cdd2, 32'h414c2593} /* (22, 27, 11) {real, imag} */,
  {32'hc1b926d4, 32'hc29e68fe} /* (22, 27, 10) {real, imag} */,
  {32'h3dc35480, 32'hc1c065cc} /* (22, 27, 9) {real, imag} */,
  {32'hc1e898e5, 32'h41e068e9} /* (22, 27, 8) {real, imag} */,
  {32'hbfdaf4a0, 32'h412a619a} /* (22, 27, 7) {real, imag} */,
  {32'h422b2aaf, 32'hc24e778c} /* (22, 27, 6) {real, imag} */,
  {32'hc281b62b, 32'h41583bd9} /* (22, 27, 5) {real, imag} */,
  {32'hc17479dd, 32'h41eadf90} /* (22, 27, 4) {real, imag} */,
  {32'h4245214a, 32'hbf7a0440} /* (22, 27, 3) {real, imag} */,
  {32'hc1882f77, 32'hc26b7bf1} /* (22, 27, 2) {real, imag} */,
  {32'hc2550e3e, 32'h43087741} /* (22, 27, 1) {real, imag} */,
  {32'h42758348, 32'h42a69388} /* (22, 27, 0) {real, imag} */,
  {32'h419ef180, 32'hc2a3a889} /* (22, 26, 31) {real, imag} */,
  {32'hc2b6fe4c, 32'h421750fc} /* (22, 26, 30) {real, imag} */,
  {32'h42429491, 32'hc1f31ba6} /* (22, 26, 29) {real, imag} */,
  {32'h40177be0, 32'hc19297f0} /* (22, 26, 28) {real, imag} */,
  {32'hc1c011b6, 32'h41d3b400} /* (22, 26, 27) {real, imag} */,
  {32'h40e5309a, 32'hc2103e16} /* (22, 26, 26) {real, imag} */,
  {32'h419b52cc, 32'h425bf80d} /* (22, 26, 25) {real, imag} */,
  {32'h4293983f, 32'hc1e4525a} /* (22, 26, 24) {real, imag} */,
  {32'hc1b42806, 32'hbfc8ee20} /* (22, 26, 23) {real, imag} */,
  {32'hc242fcb0, 32'h41d18f4d} /* (22, 26, 22) {real, imag} */,
  {32'hbf1a2058, 32'hc231cbbe} /* (22, 26, 21) {real, imag} */,
  {32'hbfe374f8, 32'hc1944e68} /* (22, 26, 20) {real, imag} */,
  {32'h40e4da32, 32'h41b20aac} /* (22, 26, 19) {real, imag} */,
  {32'h3faa1110, 32'hc179907d} /* (22, 26, 18) {real, imag} */,
  {32'hc1b07f57, 32'hc197784c} /* (22, 26, 17) {real, imag} */,
  {32'hc15ca9e6, 32'hc02df9d0} /* (22, 26, 16) {real, imag} */,
  {32'hc0f05b14, 32'hc096e298} /* (22, 26, 15) {real, imag} */,
  {32'h3eb9b8c0, 32'h41e5fcfa} /* (22, 26, 14) {real, imag} */,
  {32'hbfb538f8, 32'hc19f7554} /* (22, 26, 13) {real, imag} */,
  {32'h41a15f80, 32'h3f8d39c8} /* (22, 26, 12) {real, imag} */,
  {32'hbf91f4cc, 32'h40c175e0} /* (22, 26, 11) {real, imag} */,
  {32'hc13ee720, 32'hc27c5714} /* (22, 26, 10) {real, imag} */,
  {32'h42370863, 32'h4212cd91} /* (22, 26, 9) {real, imag} */,
  {32'h40b13e00, 32'hc17d5120} /* (22, 26, 8) {real, imag} */,
  {32'h4092f6de, 32'h411de7a4} /* (22, 26, 7) {real, imag} */,
  {32'hc04cdb34, 32'h410f85a2} /* (22, 26, 6) {real, imag} */,
  {32'hc0fbcaa0, 32'h4287a447} /* (22, 26, 5) {real, imag} */,
  {32'h429ad39d, 32'hc0537b5c} /* (22, 26, 4) {real, imag} */,
  {32'hc2d90730, 32'h3f676b30} /* (22, 26, 3) {real, imag} */,
  {32'h406b8e70, 32'hc1f42eb8} /* (22, 26, 2) {real, imag} */,
  {32'h42239bde, 32'h41fa9943} /* (22, 26, 1) {real, imag} */,
  {32'hc28378f4, 32'h42155d2e} /* (22, 26, 0) {real, imag} */,
  {32'h410ecfe2, 32'h429559f6} /* (22, 25, 31) {real, imag} */,
  {32'hc20fba36, 32'h42a3d6ab} /* (22, 25, 30) {real, imag} */,
  {32'hc15621a4, 32'hc1f1f0d9} /* (22, 25, 29) {real, imag} */,
  {32'h40f3f2f8, 32'h41df32e5} /* (22, 25, 28) {real, imag} */,
  {32'h41821a78, 32'h422367d3} /* (22, 25, 27) {real, imag} */,
  {32'h4192fa23, 32'h4250053a} /* (22, 25, 26) {real, imag} */,
  {32'hc1637b72, 32'hc0ec7eda} /* (22, 25, 25) {real, imag} */,
  {32'hc188dd6a, 32'h410a6770} /* (22, 25, 24) {real, imag} */,
  {32'h41db64c7, 32'h4214caa3} /* (22, 25, 23) {real, imag} */,
  {32'hc1d514c0, 32'h4247bc18} /* (22, 25, 22) {real, imag} */,
  {32'h4165d371, 32'hc12a6826} /* (22, 25, 21) {real, imag} */,
  {32'hc14bf5be, 32'hc11365b4} /* (22, 25, 20) {real, imag} */,
  {32'h41d1deae, 32'h3dc70300} /* (22, 25, 19) {real, imag} */,
  {32'h40436197, 32'h41054784} /* (22, 25, 18) {real, imag} */,
  {32'hc180f9ba, 32'hc1095d58} /* (22, 25, 17) {real, imag} */,
  {32'hc0545080, 32'h41d8c94f} /* (22, 25, 16) {real, imag} */,
  {32'hc0a70490, 32'hc1c02988} /* (22, 25, 15) {real, imag} */,
  {32'h40917570, 32'h40145990} /* (22, 25, 14) {real, imag} */,
  {32'hc0de0e68, 32'h41c0e399} /* (22, 25, 13) {real, imag} */,
  {32'hc09f8a0c, 32'h40f01ee5} /* (22, 25, 12) {real, imag} */,
  {32'hc0932dba, 32'h41ba79ad} /* (22, 25, 11) {real, imag} */,
  {32'h4003aaf4, 32'h419fd4e8} /* (22, 25, 10) {real, imag} */,
  {32'h41ab3bf7, 32'h41f54726} /* (22, 25, 9) {real, imag} */,
  {32'h415addd7, 32'h4282ab1a} /* (22, 25, 8) {real, imag} */,
  {32'h42382fc4, 32'h41c85fd2} /* (22, 25, 7) {real, imag} */,
  {32'h41615a82, 32'h414a9b28} /* (22, 25, 6) {real, imag} */,
  {32'h421a6423, 32'hc2484af1} /* (22, 25, 5) {real, imag} */,
  {32'h426e8b15, 32'hc23a66e8} /* (22, 25, 4) {real, imag} */,
  {32'hc20971e1, 32'hc13f6956} /* (22, 25, 3) {real, imag} */,
  {32'h41536437, 32'hc2870005} /* (22, 25, 2) {real, imag} */,
  {32'hc22280a4, 32'hc2691d85} /* (22, 25, 1) {real, imag} */,
  {32'h422760ae, 32'h423bd8f8} /* (22, 25, 0) {real, imag} */,
  {32'hc1977d43, 32'hc1d895ce} /* (22, 24, 31) {real, imag} */,
  {32'hc267cf06, 32'h421714be} /* (22, 24, 30) {real, imag} */,
  {32'h427c06a7, 32'h41c3508b} /* (22, 24, 29) {real, imag} */,
  {32'h415ced36, 32'hc250f258} /* (22, 24, 28) {real, imag} */,
  {32'h41c447ee, 32'h421426a3} /* (22, 24, 27) {real, imag} */,
  {32'h425d6051, 32'hc1ccdb47} /* (22, 24, 26) {real, imag} */,
  {32'h4287c4dc, 32'h4067d53a} /* (22, 24, 25) {real, imag} */,
  {32'hc0bc1fc8, 32'hc23eec0c} /* (22, 24, 24) {real, imag} */,
  {32'hc1f41b83, 32'h4184a1b3} /* (22, 24, 23) {real, imag} */,
  {32'hbf88a95c, 32'h408f9ed6} /* (22, 24, 22) {real, imag} */,
  {32'h41e9962c, 32'h404edc84} /* (22, 24, 21) {real, imag} */,
  {32'hc1e4c20d, 32'hc15613ce} /* (22, 24, 20) {real, imag} */,
  {32'h4120d64e, 32'hc122e34f} /* (22, 24, 19) {real, imag} */,
  {32'h41633baa, 32'h418465c7} /* (22, 24, 18) {real, imag} */,
  {32'h3fa93840, 32'hc1049548} /* (22, 24, 17) {real, imag} */,
  {32'h4145fd20, 32'hc12cb7c2} /* (22, 24, 16) {real, imag} */,
  {32'h3f8a79c0, 32'h414a68ee} /* (22, 24, 15) {real, imag} */,
  {32'h4129d326, 32'h40a4edfc} /* (22, 24, 14) {real, imag} */,
  {32'h3fadcf50, 32'h41228071} /* (22, 24, 13) {real, imag} */,
  {32'hc1aafd3f, 32'hc1819ec1} /* (22, 24, 12) {real, imag} */,
  {32'h3f617b20, 32'hc14759a1} /* (22, 24, 11) {real, imag} */,
  {32'hc14caf3c, 32'h40b816e6} /* (22, 24, 10) {real, imag} */,
  {32'hc00e2b98, 32'hc110ff38} /* (22, 24, 9) {real, imag} */,
  {32'h41a2fa64, 32'hc0565848} /* (22, 24, 8) {real, imag} */,
  {32'hc2349aa7, 32'hc0c9f7df} /* (22, 24, 7) {real, imag} */,
  {32'hc26635fb, 32'h4191b4b9} /* (22, 24, 6) {real, imag} */,
  {32'h4213f105, 32'h4100a5bb} /* (22, 24, 5) {real, imag} */,
  {32'hc1fa7a53, 32'h42236ca0} /* (22, 24, 4) {real, imag} */,
  {32'hc228e4a5, 32'hc1a116b5} /* (22, 24, 3) {real, imag} */,
  {32'hc19d7a30, 32'hc203ec00} /* (22, 24, 2) {real, imag} */,
  {32'hc106b42e, 32'hc1558cdd} /* (22, 24, 1) {real, imag} */,
  {32'h42aa4656, 32'h41fb0e75} /* (22, 24, 0) {real, imag} */,
  {32'hc2116038, 32'hc227f491} /* (22, 23, 31) {real, imag} */,
  {32'hc09b86f4, 32'hc2b132d8} /* (22, 23, 30) {real, imag} */,
  {32'h422ec116, 32'hc1f3f9b1} /* (22, 23, 29) {real, imag} */,
  {32'h41c31cd7, 32'hc1ad2412} /* (22, 23, 28) {real, imag} */,
  {32'hc0f70274, 32'hc1385918} /* (22, 23, 27) {real, imag} */,
  {32'h411af21a, 32'h41855096} /* (22, 23, 26) {real, imag} */,
  {32'h4223e2df, 32'hc244e624} /* (22, 23, 25) {real, imag} */,
  {32'h424f4704, 32'hbfbdc564} /* (22, 23, 24) {real, imag} */,
  {32'h40280ea0, 32'hc1f3e8a2} /* (22, 23, 23) {real, imag} */,
  {32'h4136db93, 32'h41e3bee8} /* (22, 23, 22) {real, imag} */,
  {32'h41030039, 32'h416eac3e} /* (22, 23, 21) {real, imag} */,
  {32'h4100f576, 32'hbf5c8dd8} /* (22, 23, 20) {real, imag} */,
  {32'hc1a8563d, 32'hc039f302} /* (22, 23, 19) {real, imag} */,
  {32'hc0887236, 32'hbf8c3be0} /* (22, 23, 18) {real, imag} */,
  {32'h40c4e116, 32'h3f1f86a0} /* (22, 23, 17) {real, imag} */,
  {32'hbf742bc8, 32'hc12bf1ec} /* (22, 23, 16) {real, imag} */,
  {32'hbf2c9590, 32'hc110eadc} /* (22, 23, 15) {real, imag} */,
  {32'hc11e2a0f, 32'hc04f8d90} /* (22, 23, 14) {real, imag} */,
  {32'hc0ecd0a3, 32'hbfe4f91c} /* (22, 23, 13) {real, imag} */,
  {32'hc1aa4c4f, 32'h40fbe977} /* (22, 23, 12) {real, imag} */,
  {32'hc1856360, 32'h40f953fb} /* (22, 23, 11) {real, imag} */,
  {32'hc1618dbb, 32'hc20bbdd6} /* (22, 23, 10) {real, imag} */,
  {32'hc139f31a, 32'hc1d448e0} /* (22, 23, 9) {real, imag} */,
  {32'h412644c6, 32'h3e53fc20} /* (22, 23, 8) {real, imag} */,
  {32'h40d02508, 32'h40eb8fa8} /* (22, 23, 7) {real, imag} */,
  {32'hbf9c4840, 32'h42053043} /* (22, 23, 6) {real, imag} */,
  {32'h41f343ab, 32'hc217cacf} /* (22, 23, 5) {real, imag} */,
  {32'hc12b9c7e, 32'hc1525dcc} /* (22, 23, 4) {real, imag} */,
  {32'h41119fda, 32'hc219c85b} /* (22, 23, 3) {real, imag} */,
  {32'hc211747e, 32'hc1bcba78} /* (22, 23, 2) {real, imag} */,
  {32'h4181205b, 32'hc18c57de} /* (22, 23, 1) {real, imag} */,
  {32'h3fee1034, 32'h42429bde} /* (22, 23, 0) {real, imag} */,
  {32'h4249f9b7, 32'h41f54a88} /* (22, 22, 31) {real, imag} */,
  {32'h41a9aea2, 32'h41c20540} /* (22, 22, 30) {real, imag} */,
  {32'h41d99759, 32'hc0798e54} /* (22, 22, 29) {real, imag} */,
  {32'hc20f7d19, 32'h4266bfa6} /* (22, 22, 28) {real, imag} */,
  {32'hc0aee83c, 32'h40f7817e} /* (22, 22, 27) {real, imag} */,
  {32'h41c3dc9a, 32'hc22fd7ae} /* (22, 22, 26) {real, imag} */,
  {32'hc18f07e0, 32'h41401637} /* (22, 22, 25) {real, imag} */,
  {32'hc02c20f0, 32'hc1a8bc52} /* (22, 22, 24) {real, imag} */,
  {32'hc1ca0c29, 32'h415c6e19} /* (22, 22, 23) {real, imag} */,
  {32'hc1dc55d4, 32'h40b19d4a} /* (22, 22, 22) {real, imag} */,
  {32'h41c0c745, 32'h416ec637} /* (22, 22, 21) {real, imag} */,
  {32'h3f25f4fc, 32'h4126b9ed} /* (22, 22, 20) {real, imag} */,
  {32'h3f694830, 32'h4106cd80} /* (22, 22, 19) {real, imag} */,
  {32'h3fbc4e9c, 32'hc16a0c9a} /* (22, 22, 18) {real, imag} */,
  {32'h415dc0d2, 32'h403b64d4} /* (22, 22, 17) {real, imag} */,
  {32'hc100e639, 32'h3f9672e0} /* (22, 22, 16) {real, imag} */,
  {32'h402630a6, 32'h40d2848a} /* (22, 22, 15) {real, imag} */,
  {32'hc05a109e, 32'hc1628796} /* (22, 22, 14) {real, imag} */,
  {32'h417cdb43, 32'hc0f335f3} /* (22, 22, 13) {real, imag} */,
  {32'h4109c5f4, 32'h413c7d89} /* (22, 22, 12) {real, imag} */,
  {32'h41c4a43b, 32'hbef90560} /* (22, 22, 11) {real, imag} */,
  {32'h40439db4, 32'hc202d5e0} /* (22, 22, 10) {real, imag} */,
  {32'h41e0e91b, 32'h41eef1d6} /* (22, 22, 9) {real, imag} */,
  {32'h41d6bf6c, 32'h40a5bbce} /* (22, 22, 8) {real, imag} */,
  {32'h40b03890, 32'hc0cd81b6} /* (22, 22, 7) {real, imag} */,
  {32'hc16b6f47, 32'h41050dc2} /* (22, 22, 6) {real, imag} */,
  {32'h413012b8, 32'h41eb84be} /* (22, 22, 5) {real, imag} */,
  {32'hc1b87ea4, 32'hc1eb281c} /* (22, 22, 4) {real, imag} */,
  {32'h41ac73fb, 32'hc18a376e} /* (22, 22, 3) {real, imag} */,
  {32'h418e0c9a, 32'h4078dec0} /* (22, 22, 2) {real, imag} */,
  {32'h420427e9, 32'hc1b81e56} /* (22, 22, 1) {real, imag} */,
  {32'hc174ec43, 32'hbf42f280} /* (22, 22, 0) {real, imag} */,
  {32'hc007c589, 32'h42121dad} /* (22, 21, 31) {real, imag} */,
  {32'h3faed53b, 32'hbffdf630} /* (22, 21, 30) {real, imag} */,
  {32'hc252a1e0, 32'hc0a3fa7e} /* (22, 21, 29) {real, imag} */,
  {32'hc2848b18, 32'h40303238} /* (22, 21, 28) {real, imag} */,
  {32'hc00f8d2c, 32'hc231e0a4} /* (22, 21, 27) {real, imag} */,
  {32'h403c5c7c, 32'h41d26c8b} /* (22, 21, 26) {real, imag} */,
  {32'hc0853b66, 32'h420c39f7} /* (22, 21, 25) {real, imag} */,
  {32'hc0a452f2, 32'hc275ec9e} /* (22, 21, 24) {real, imag} */,
  {32'hc179d600, 32'hc12effbb} /* (22, 21, 23) {real, imag} */,
  {32'hc128367b, 32'hc0762538} /* (22, 21, 22) {real, imag} */,
  {32'hc17ea705, 32'hc1736052} /* (22, 21, 21) {real, imag} */,
  {32'h4055f040, 32'hc047a3d8} /* (22, 21, 20) {real, imag} */,
  {32'h41334d0d, 32'h3f8e9cb6} /* (22, 21, 19) {real, imag} */,
  {32'hc0c3a4d6, 32'hbd28d600} /* (22, 21, 18) {real, imag} */,
  {32'h4008e2e0, 32'h3fcb1724} /* (22, 21, 17) {real, imag} */,
  {32'hc09bfff8, 32'h4124bf01} /* (22, 21, 16) {real, imag} */,
  {32'h40c50c58, 32'hc08ad431} /* (22, 21, 15) {real, imag} */,
  {32'hc0c5f3ae, 32'hc13aaf0e} /* (22, 21, 14) {real, imag} */,
  {32'h40f0928a, 32'h408a5d80} /* (22, 21, 13) {real, imag} */,
  {32'h40031ba0, 32'h41886313} /* (22, 21, 12) {real, imag} */,
  {32'hc1ad1b2e, 32'h418ddfed} /* (22, 21, 11) {real, imag} */,
  {32'hc1f9a7e4, 32'hc1c9b3f3} /* (22, 21, 10) {real, imag} */,
  {32'hc1a1e13c, 32'hc14e305f} /* (22, 21, 9) {real, imag} */,
  {32'hc19166ba, 32'hc22c6176} /* (22, 21, 8) {real, imag} */,
  {32'h4146973d, 32'hc099b56e} /* (22, 21, 7) {real, imag} */,
  {32'hc10b1c53, 32'hc1fccad5} /* (22, 21, 6) {real, imag} */,
  {32'hc19c4626, 32'h4166a026} /* (22, 21, 5) {real, imag} */,
  {32'h400b6950, 32'h425f0bf6} /* (22, 21, 4) {real, imag} */,
  {32'h42480be6, 32'hc18f32e0} /* (22, 21, 3) {real, imag} */,
  {32'h3fe1e7f5, 32'h426d233a} /* (22, 21, 2) {real, imag} */,
  {32'hbcff0080, 32'h421d97e7} /* (22, 21, 1) {real, imag} */,
  {32'hc1ebb2a8, 32'hc11b2c15} /* (22, 21, 0) {real, imag} */,
  {32'h402d642b, 32'h42108dc7} /* (22, 20, 31) {real, imag} */,
  {32'h4202844e, 32'h41223a8c} /* (22, 20, 30) {real, imag} */,
  {32'hc0904876, 32'hc108d8f0} /* (22, 20, 29) {real, imag} */,
  {32'hc130d02d, 32'h3ca85b80} /* (22, 20, 28) {real, imag} */,
  {32'hc263da6a, 32'hc1bda6a2} /* (22, 20, 27) {real, imag} */,
  {32'hc163add6, 32'hc0c40ee2} /* (22, 20, 26) {real, imag} */,
  {32'h41d87586, 32'h41ca890d} /* (22, 20, 25) {real, imag} */,
  {32'h41170e2c, 32'h4204c510} /* (22, 20, 24) {real, imag} */,
  {32'h416023d3, 32'hc1b5f409} /* (22, 20, 23) {real, imag} */,
  {32'h405a0180, 32'hc1acbf78} /* (22, 20, 22) {real, imag} */,
  {32'h411af365, 32'h406eaed2} /* (22, 20, 21) {real, imag} */,
  {32'h40c30aec, 32'hbf3dee0c} /* (22, 20, 20) {real, imag} */,
  {32'h412e09bb, 32'h40cb0aaf} /* (22, 20, 19) {real, imag} */,
  {32'h4145bb6e, 32'h3fdb3db4} /* (22, 20, 18) {real, imag} */,
  {32'h3f177da4, 32'hc14de58a} /* (22, 20, 17) {real, imag} */,
  {32'hc11848ee, 32'h3eb18c40} /* (22, 20, 16) {real, imag} */,
  {32'h3ef25de8, 32'h409e926b} /* (22, 20, 15) {real, imag} */,
  {32'h40996f1c, 32'hbdab5ac0} /* (22, 20, 14) {real, imag} */,
  {32'h41481d85, 32'h411e7d7a} /* (22, 20, 13) {real, imag} */,
  {32'hbe9c2e00, 32'hc0cb52da} /* (22, 20, 12) {real, imag} */,
  {32'hc1646191, 32'hc0ead5f1} /* (22, 20, 11) {real, imag} */,
  {32'hc18335e7, 32'h3f57b110} /* (22, 20, 10) {real, imag} */,
  {32'h4124f23d, 32'hc0b3e984} /* (22, 20, 9) {real, imag} */,
  {32'hc1c22ed4, 32'h4202c722} /* (22, 20, 8) {real, imag} */,
  {32'hc19ad65a, 32'hbda52700} /* (22, 20, 7) {real, imag} */,
  {32'h414ae0e4, 32'h4122bd97} /* (22, 20, 6) {real, imag} */,
  {32'hc192c47b, 32'hc2376687} /* (22, 20, 5) {real, imag} */,
  {32'h4214a041, 32'h40073d6f} /* (22, 20, 4) {real, imag} */,
  {32'h41ca170c, 32'hc129d38a} /* (22, 20, 3) {real, imag} */,
  {32'h420da722, 32'hc121d03c} /* (22, 20, 2) {real, imag} */,
  {32'h408662b8, 32'hc20c5c7f} /* (22, 20, 1) {real, imag} */,
  {32'hc23049f2, 32'hbe547e80} /* (22, 20, 0) {real, imag} */,
  {32'hc11ebe8e, 32'h41a5efdd} /* (22, 19, 31) {real, imag} */,
  {32'h41426cc7, 32'h4056c966} /* (22, 19, 30) {real, imag} */,
  {32'h40e3026c, 32'hc0fb14ef} /* (22, 19, 29) {real, imag} */,
  {32'hc131a4a6, 32'hc0700b64} /* (22, 19, 28) {real, imag} */,
  {32'h41960cc5, 32'hc16c1365} /* (22, 19, 27) {real, imag} */,
  {32'h4036cb72, 32'h3ef69100} /* (22, 19, 26) {real, imag} */,
  {32'h4149c79e, 32'hbffeacc0} /* (22, 19, 25) {real, imag} */,
  {32'h40e79280, 32'h4086c6d7} /* (22, 19, 24) {real, imag} */,
  {32'h3fd598a4, 32'hc18578da} /* (22, 19, 23) {real, imag} */,
  {32'h418ce544, 32'h3f041d60} /* (22, 19, 22) {real, imag} */,
  {32'hc0ae4250, 32'hc0e979a2} /* (22, 19, 21) {real, imag} */,
  {32'h411d33de, 32'h3fa7e6a8} /* (22, 19, 20) {real, imag} */,
  {32'hc0e88c77, 32'h40e1530f} /* (22, 19, 19) {real, imag} */,
  {32'hc098c716, 32'h407b2e4e} /* (22, 19, 18) {real, imag} */,
  {32'h3ea7bcf0, 32'hc111d212} /* (22, 19, 17) {real, imag} */,
  {32'hc0746cb5, 32'h4158795e} /* (22, 19, 16) {real, imag} */,
  {32'hbff0c7c4, 32'hc00d9460} /* (22, 19, 15) {real, imag} */,
  {32'hc0e14a0c, 32'hc15d7542} /* (22, 19, 14) {real, imag} */,
  {32'h40ef03f9, 32'hc0f90839} /* (22, 19, 13) {real, imag} */,
  {32'hc140e8fe, 32'hc18ee74a} /* (22, 19, 12) {real, imag} */,
  {32'hbe493690, 32'h3fa5abfa} /* (22, 19, 11) {real, imag} */,
  {32'h3fba60c0, 32'hc079ce0c} /* (22, 19, 10) {real, imag} */,
  {32'h413eadde, 32'h40a7c397} /* (22, 19, 9) {real, imag} */,
  {32'hc14cbcf0, 32'h3cfa1100} /* (22, 19, 8) {real, imag} */,
  {32'h412cabf8, 32'h406aa304} /* (22, 19, 7) {real, imag} */,
  {32'h41113c64, 32'hc15be47d} /* (22, 19, 6) {real, imag} */,
  {32'h41a89abf, 32'hc0210344} /* (22, 19, 5) {real, imag} */,
  {32'hc18dd90b, 32'h41a354ec} /* (22, 19, 4) {real, imag} */,
  {32'hc202a046, 32'h4132f8b8} /* (22, 19, 3) {real, imag} */,
  {32'h41a6b498, 32'h40c74c0f} /* (22, 19, 2) {real, imag} */,
  {32'h41d65675, 32'h411ac424} /* (22, 19, 1) {real, imag} */,
  {32'h4124906a, 32'hc21b7734} /* (22, 19, 0) {real, imag} */,
  {32'hc2093744, 32'hc227b199} /* (22, 18, 31) {real, imag} */,
  {32'hc16c0720, 32'h3ecea490} /* (22, 18, 30) {real, imag} */,
  {32'h4197711e, 32'h3fb611d8} /* (22, 18, 29) {real, imag} */,
  {32'h4009a3fc, 32'hc1eb1616} /* (22, 18, 28) {real, imag} */,
  {32'hc163cbfe, 32'h4167633b} /* (22, 18, 27) {real, imag} */,
  {32'hc09ca25b, 32'h41b16a7c} /* (22, 18, 26) {real, imag} */,
  {32'h40935c66, 32'h4182a402} /* (22, 18, 25) {real, imag} */,
  {32'hbfb783ec, 32'h40d2353c} /* (22, 18, 24) {real, imag} */,
  {32'hc1902a6c, 32'h40c6d2fc} /* (22, 18, 23) {real, imag} */,
  {32'h40123320, 32'h41aea1db} /* (22, 18, 22) {real, imag} */,
  {32'hc12fe7a9, 32'h406d8158} /* (22, 18, 21) {real, imag} */,
  {32'h40f2705c, 32'hc0cde891} /* (22, 18, 20) {real, imag} */,
  {32'hbebceaf8, 32'hbf640348} /* (22, 18, 19) {real, imag} */,
  {32'hbfa4ae10, 32'hc0ff98cd} /* (22, 18, 18) {real, imag} */,
  {32'hc083bc66, 32'hc0d80182} /* (22, 18, 17) {real, imag} */,
  {32'h404a3f58, 32'h3f2ac338} /* (22, 18, 16) {real, imag} */,
  {32'hc05e035c, 32'h414756af} /* (22, 18, 15) {real, imag} */,
  {32'hc0d49248, 32'h3f184d68} /* (22, 18, 14) {real, imag} */,
  {32'hc0ea1976, 32'h3f5e2760} /* (22, 18, 13) {real, imag} */,
  {32'h415a9fee, 32'hc0881e53} /* (22, 18, 12) {real, imag} */,
  {32'h412ac02f, 32'hc0b6391c} /* (22, 18, 11) {real, imag} */,
  {32'h4166b0e8, 32'hc00cae50} /* (22, 18, 10) {real, imag} */,
  {32'h41144ff9, 32'h417a80d2} /* (22, 18, 9) {real, imag} */,
  {32'h40701696, 32'h409949da} /* (22, 18, 8) {real, imag} */,
  {32'hc10d0705, 32'h414068a0} /* (22, 18, 7) {real, imag} */,
  {32'h41205ea8, 32'h4184ace0} /* (22, 18, 6) {real, imag} */,
  {32'h3f0695b8, 32'hc1aba2dc} /* (22, 18, 5) {real, imag} */,
  {32'h419385ba, 32'hc004878c} /* (22, 18, 4) {real, imag} */,
  {32'hc18ef8dc, 32'h413987fd} /* (22, 18, 3) {real, imag} */,
  {32'h41b5fe9c, 32'hc029252a} /* (22, 18, 2) {real, imag} */,
  {32'h3ffa3d90, 32'hc0749eb0} /* (22, 18, 1) {real, imag} */,
  {32'hc16b68a6, 32'hc184c91a} /* (22, 18, 0) {real, imag} */,
  {32'hc04ab125, 32'h40d41336} /* (22, 17, 31) {real, imag} */,
  {32'h4036af38, 32'hc0a3d715} /* (22, 17, 30) {real, imag} */,
  {32'h4059981a, 32'h406ca6ee} /* (22, 17, 29) {real, imag} */,
  {32'h41137b40, 32'hbf77da05} /* (22, 17, 28) {real, imag} */,
  {32'h41e24eb2, 32'hbfe2b648} /* (22, 17, 27) {real, imag} */,
  {32'hc03f1122, 32'hc024f1dd} /* (22, 17, 26) {real, imag} */,
  {32'h40f2a822, 32'hc19c5f3f} /* (22, 17, 25) {real, imag} */,
  {32'h40110e48, 32'hbf58e410} /* (22, 17, 24) {real, imag} */,
  {32'h4021c81c, 32'h41857ff6} /* (22, 17, 23) {real, imag} */,
  {32'hc07b304c, 32'hc0bf2ce8} /* (22, 17, 22) {real, imag} */,
  {32'h40c347e0, 32'h414a6ca6} /* (22, 17, 21) {real, imag} */,
  {32'hbfe80294, 32'hc0a9e474} /* (22, 17, 20) {real, imag} */,
  {32'hbfd67044, 32'h41347b6a} /* (22, 17, 19) {real, imag} */,
  {32'hc0ad7c66, 32'hc13726a6} /* (22, 17, 18) {real, imag} */,
  {32'hbf991cbe, 32'h4040acf7} /* (22, 17, 17) {real, imag} */,
  {32'h40310854, 32'hbfcabd30} /* (22, 17, 16) {real, imag} */,
  {32'hbf70398c, 32'h3ffeba7e} /* (22, 17, 15) {real, imag} */,
  {32'h4035ade4, 32'h408cda2f} /* (22, 17, 14) {real, imag} */,
  {32'h40901349, 32'hc179d812} /* (22, 17, 13) {real, imag} */,
  {32'hbe91f6a0, 32'h410db16a} /* (22, 17, 12) {real, imag} */,
  {32'hc01da660, 32'hc0b5e924} /* (22, 17, 11) {real, imag} */,
  {32'h417d2cf1, 32'hc0084da1} /* (22, 17, 10) {real, imag} */,
  {32'hc19702d2, 32'hc1278fd5} /* (22, 17, 9) {real, imag} */,
  {32'hbf3b6d40, 32'hc19dd63a} /* (22, 17, 8) {real, imag} */,
  {32'h41c6e286, 32'h420f1630} /* (22, 17, 7) {real, imag} */,
  {32'hc0d67327, 32'h40926406} /* (22, 17, 6) {real, imag} */,
  {32'hc1656444, 32'h3d689500} /* (22, 17, 5) {real, imag} */,
  {32'hc0f3cc35, 32'h40089e8f} /* (22, 17, 4) {real, imag} */,
  {32'h415b2a12, 32'hc19a80e8} /* (22, 17, 3) {real, imag} */,
  {32'h416a758c, 32'hc122d10a} /* (22, 17, 2) {real, imag} */,
  {32'hc0337599, 32'hc133453f} /* (22, 17, 1) {real, imag} */,
  {32'h3fa88f88, 32'hc1dd0e40} /* (22, 17, 0) {real, imag} */,
  {32'h41beff5f, 32'hc1013de2} /* (22, 16, 31) {real, imag} */,
  {32'h41907af6, 32'h410ec676} /* (22, 16, 30) {real, imag} */,
  {32'h41c75f52, 32'hc18248b8} /* (22, 16, 29) {real, imag} */,
  {32'h41b357e2, 32'hc12071cc} /* (22, 16, 28) {real, imag} */,
  {32'h40c17c99, 32'h4157a39e} /* (22, 16, 27) {real, imag} */,
  {32'hc0bc3174, 32'hc0f54e17} /* (22, 16, 26) {real, imag} */,
  {32'hbe8ea178, 32'h3fdf18a8} /* (22, 16, 25) {real, imag} */,
  {32'hc12fa148, 32'hc11e0ac6} /* (22, 16, 24) {real, imag} */,
  {32'h407c2e1c, 32'h409838e8} /* (22, 16, 23) {real, imag} */,
  {32'h40003e33, 32'hbd0a94e0} /* (22, 16, 22) {real, imag} */,
  {32'h3f09c568, 32'hc0f117d1} /* (22, 16, 21) {real, imag} */,
  {32'h3ee9eea0, 32'hc0704145} /* (22, 16, 20) {real, imag} */,
  {32'hc0c77be6, 32'hbfd3d458} /* (22, 16, 19) {real, imag} */,
  {32'h40a00482, 32'hc0a8780e} /* (22, 16, 18) {real, imag} */,
  {32'h4040d3ab, 32'h409d9b57} /* (22, 16, 17) {real, imag} */,
  {32'hbfce95ec, 32'h3f9f1da4} /* (22, 16, 16) {real, imag} */,
  {32'h403b3693, 32'hc0a38305} /* (22, 16, 15) {real, imag} */,
  {32'h4067fb03, 32'h4085d71e} /* (22, 16, 14) {real, imag} */,
  {32'h4048f4d5, 32'hc08eaeee} /* (22, 16, 13) {real, imag} */,
  {32'hc11d1821, 32'hc0b98ca4} /* (22, 16, 12) {real, imag} */,
  {32'hc10ef656, 32'h3e3320e0} /* (22, 16, 11) {real, imag} */,
  {32'hc09053fc, 32'hbe4510b8} /* (22, 16, 10) {real, imag} */,
  {32'h4179b185, 32'h4106ae3e} /* (22, 16, 9) {real, imag} */,
  {32'hc0cebfc1, 32'h401c4ee0} /* (22, 16, 8) {real, imag} */,
  {32'h405816f7, 32'hc2067e7f} /* (22, 16, 7) {real, imag} */,
  {32'h412b71b6, 32'h410bbc37} /* (22, 16, 6) {real, imag} */,
  {32'hc1125f06, 32'hc164976e} /* (22, 16, 5) {real, imag} */,
  {32'hc1dbafb6, 32'h40bf50d1} /* (22, 16, 4) {real, imag} */,
  {32'hc1aeefda, 32'h40aaa78e} /* (22, 16, 3) {real, imag} */,
  {32'h4009e580, 32'h40aa6600} /* (22, 16, 2) {real, imag} */,
  {32'hc1a5453d, 32'h40ac8c80} /* (22, 16, 1) {real, imag} */,
  {32'h418bcb55, 32'hc0562c5a} /* (22, 16, 0) {real, imag} */,
  {32'h40032fc3, 32'h3f93cbf2} /* (22, 15, 31) {real, imag} */,
  {32'h3f5c3630, 32'h41b93993} /* (22, 15, 30) {real, imag} */,
  {32'h4090e7a6, 32'hc12e43ae} /* (22, 15, 29) {real, imag} */,
  {32'hc1b5a99e, 32'hc1fcaf22} /* (22, 15, 28) {real, imag} */,
  {32'h403657c2, 32'h4115c76d} /* (22, 15, 27) {real, imag} */,
  {32'hc089c5e8, 32'h4175cdd3} /* (22, 15, 26) {real, imag} */,
  {32'h402393b0, 32'h4095ad3c} /* (22, 15, 25) {real, imag} */,
  {32'hbf997938, 32'h418505fb} /* (22, 15, 24) {real, imag} */,
  {32'h3fc1f130, 32'hc0f96428} /* (22, 15, 23) {real, imag} */,
  {32'hc134e49a, 32'hc0be73d4} /* (22, 15, 22) {real, imag} */,
  {32'h40589c46, 32'hc0cc273f} /* (22, 15, 21) {real, imag} */,
  {32'hc095e1aa, 32'h3fcdc874} /* (22, 15, 20) {real, imag} */,
  {32'h4012c526, 32'hc0997cb2} /* (22, 15, 19) {real, imag} */,
  {32'h410a3788, 32'h3fa51ab0} /* (22, 15, 18) {real, imag} */,
  {32'h408f3c18, 32'hbcbab580} /* (22, 15, 17) {real, imag} */,
  {32'hbf0fc3f8, 32'h3e3d7080} /* (22, 15, 16) {real, imag} */,
  {32'hbc09d700, 32'hbed073d8} /* (22, 15, 15) {real, imag} */,
  {32'h402850f6, 32'h40ac2784} /* (22, 15, 14) {real, imag} */,
  {32'h409d8868, 32'h40eb0fa0} /* (22, 15, 13) {real, imag} */,
  {32'h3e9c4c20, 32'hc12341dc} /* (22, 15, 12) {real, imag} */,
  {32'hbfb72755, 32'hbf89c330} /* (22, 15, 11) {real, imag} */,
  {32'hc143e8e6, 32'h40669f10} /* (22, 15, 10) {real, imag} */,
  {32'h41c3a501, 32'hba496000} /* (22, 15, 9) {real, imag} */,
  {32'h410b9965, 32'hc1219c96} /* (22, 15, 8) {real, imag} */,
  {32'h4097a21a, 32'hc13be796} /* (22, 15, 7) {real, imag} */,
  {32'h407d34c0, 32'hc0f23a7e} /* (22, 15, 6) {real, imag} */,
  {32'hc1283058, 32'h410cb17d} /* (22, 15, 5) {real, imag} */,
  {32'h4097fd34, 32'hc087a3de} /* (22, 15, 4) {real, imag} */,
  {32'hc04d92b2, 32'h4143598a} /* (22, 15, 3) {real, imag} */,
  {32'h40e7f0f0, 32'h41f28f61} /* (22, 15, 2) {real, imag} */,
  {32'hc110bc4d, 32'hc10ab0c4} /* (22, 15, 1) {real, imag} */,
  {32'h413de90c, 32'h4040fe68} /* (22, 15, 0) {real, imag} */,
  {32'h421b2446, 32'hc03904d6} /* (22, 14, 31) {real, imag} */,
  {32'h3ee48c4c, 32'hc1a77b49} /* (22, 14, 30) {real, imag} */,
  {32'h40f264c9, 32'h418395c5} /* (22, 14, 29) {real, imag} */,
  {32'h40c7e722, 32'hc12408ab} /* (22, 14, 28) {real, imag} */,
  {32'h41eaa661, 32'h4142d186} /* (22, 14, 27) {real, imag} */,
  {32'hc1018001, 32'hc11f34a8} /* (22, 14, 26) {real, imag} */,
  {32'h3fd97cb4, 32'h40f81dc6} /* (22, 14, 25) {real, imag} */,
  {32'h4103e098, 32'h40af2957} /* (22, 14, 24) {real, imag} */,
  {32'hc11f0cd1, 32'h40e449fb} /* (22, 14, 23) {real, imag} */,
  {32'h40f04623, 32'hc178027a} /* (22, 14, 22) {real, imag} */,
  {32'hbf4aa6a0, 32'h40bebfa6} /* (22, 14, 21) {real, imag} */,
  {32'h41493826, 32'h41d48af2} /* (22, 14, 20) {real, imag} */,
  {32'hc0c8b249, 32'hc08d834c} /* (22, 14, 19) {real, imag} */,
  {32'h4052a716, 32'hc08e57c6} /* (22, 14, 18) {real, imag} */,
  {32'hc05b1958, 32'h401c9d93} /* (22, 14, 17) {real, imag} */,
  {32'hbfa18bd8, 32'hc001b17c} /* (22, 14, 16) {real, imag} */,
  {32'h40242090, 32'hc052b737} /* (22, 14, 15) {real, imag} */,
  {32'hc11ec414, 32'hbff55e76} /* (22, 14, 14) {real, imag} */,
  {32'h3f9258e4, 32'hc0607f4f} /* (22, 14, 13) {real, imag} */,
  {32'hc11df454, 32'hc0eab77e} /* (22, 14, 12) {real, imag} */,
  {32'hc0e07a54, 32'h405d8870} /* (22, 14, 11) {real, imag} */,
  {32'h4117150f, 32'hc1843ed9} /* (22, 14, 10) {real, imag} */,
  {32'h41861549, 32'hc0f1ac85} /* (22, 14, 9) {real, imag} */,
  {32'hbf08d8dc, 32'hc0d2aca1} /* (22, 14, 8) {real, imag} */,
  {32'h411fadb0, 32'hc0d4a2e6} /* (22, 14, 7) {real, imag} */,
  {32'hc1145ed7, 32'h4082ae28} /* (22, 14, 6) {real, imag} */,
  {32'h413bb12a, 32'hc147d1b2} /* (22, 14, 5) {real, imag} */,
  {32'h41aaa660, 32'h412cc4f1} /* (22, 14, 4) {real, imag} */,
  {32'h3e9a26b0, 32'h40f36b50} /* (22, 14, 3) {real, imag} */,
  {32'h4056982e, 32'hc1efe047} /* (22, 14, 2) {real, imag} */,
  {32'hbeb84500, 32'h40e5ed09} /* (22, 14, 1) {real, imag} */,
  {32'hc12785c3, 32'h41c5edd4} /* (22, 14, 0) {real, imag} */,
  {32'h41a961be, 32'h3d8bf640} /* (22, 13, 31) {real, imag} */,
  {32'h41d104d4, 32'hc15d76c5} /* (22, 13, 30) {real, imag} */,
  {32'hc1e3263e, 32'hbf4a6560} /* (22, 13, 29) {real, imag} */,
  {32'hc18128f0, 32'h41334de6} /* (22, 13, 28) {real, imag} */,
  {32'h406fb538, 32'hbdd8c780} /* (22, 13, 27) {real, imag} */,
  {32'h426f25ca, 32'h41b59b84} /* (22, 13, 26) {real, imag} */,
  {32'h413543ae, 32'h414f8bfc} /* (22, 13, 25) {real, imag} */,
  {32'hc0eff44f, 32'hc0331848} /* (22, 13, 24) {real, imag} */,
  {32'hc19632c9, 32'h40b4675e} /* (22, 13, 23) {real, imag} */,
  {32'h40d324b4, 32'hc18748e5} /* (22, 13, 22) {real, imag} */,
  {32'hc0ec1614, 32'h40b84dce} /* (22, 13, 21) {real, imag} */,
  {32'hc0cd0002, 32'h40eff78f} /* (22, 13, 20) {real, imag} */,
  {32'h40edfbe0, 32'hc11d2883} /* (22, 13, 19) {real, imag} */,
  {32'h3f8566a0, 32'hc1798f22} /* (22, 13, 18) {real, imag} */,
  {32'h404dbcf0, 32'hc0925c23} /* (22, 13, 17) {real, imag} */,
  {32'h410e8131, 32'h40b321e0} /* (22, 13, 16) {real, imag} */,
  {32'h41114d60, 32'h411b1d2c} /* (22, 13, 15) {real, imag} */,
  {32'h403fe470, 32'hc100ea52} /* (22, 13, 14) {real, imag} */,
  {32'hc0f64e1a, 32'hc0a89cbe} /* (22, 13, 13) {real, imag} */,
  {32'h400c8ddc, 32'hc053abee} /* (22, 13, 12) {real, imag} */,
  {32'h3ec9a9e0, 32'h418821e2} /* (22, 13, 11) {real, imag} */,
  {32'h4139a1e6, 32'h417dc02a} /* (22, 13, 10) {real, imag} */,
  {32'hc169bbf2, 32'h41a52612} /* (22, 13, 9) {real, imag} */,
  {32'h40467a62, 32'hc1310aba} /* (22, 13, 8) {real, imag} */,
  {32'hc18ed20f, 32'hc15b4586} /* (22, 13, 7) {real, imag} */,
  {32'h4166bcea, 32'hc0987b26} /* (22, 13, 6) {real, imag} */,
  {32'hc1dc66fb, 32'hc1bcb944} /* (22, 13, 5) {real, imag} */,
  {32'h421dc56e, 32'h3fec2024} /* (22, 13, 4) {real, imag} */,
  {32'h417e5123, 32'h413158da} /* (22, 13, 3) {real, imag} */,
  {32'hc1ba7294, 32'hc19921cc} /* (22, 13, 2) {real, imag} */,
  {32'hc0b63828, 32'hc10de5de} /* (22, 13, 1) {real, imag} */,
  {32'hc11dec5f, 32'h4091670c} /* (22, 13, 0) {real, imag} */,
  {32'hc09cadbc, 32'hc2046c55} /* (22, 12, 31) {real, imag} */,
  {32'h41417b96, 32'hc0408922} /* (22, 12, 30) {real, imag} */,
  {32'hc20298e4, 32'h4042bcd8} /* (22, 12, 29) {real, imag} */,
  {32'hc1bcd3f0, 32'h41eeddc0} /* (22, 12, 28) {real, imag} */,
  {32'h3ff8c5c2, 32'h3e9356bc} /* (22, 12, 27) {real, imag} */,
  {32'h41fee736, 32'h42050f00} /* (22, 12, 26) {real, imag} */,
  {32'hc1896182, 32'hc1bce8af} /* (22, 12, 25) {real, imag} */,
  {32'hc088ef0d, 32'hc17f0422} /* (22, 12, 24) {real, imag} */,
  {32'hc167709c, 32'hc139d1d6} /* (22, 12, 23) {real, imag} */,
  {32'hc1923d74, 32'hbd8ec740} /* (22, 12, 22) {real, imag} */,
  {32'hc1225188, 32'h3f542a58} /* (22, 12, 21) {real, imag} */,
  {32'hc153377e, 32'hc13bd60e} /* (22, 12, 20) {real, imag} */,
  {32'h40cc3fb8, 32'h3f756bf0} /* (22, 12, 19) {real, imag} */,
  {32'h414e5b8e, 32'h4147c4b8} /* (22, 12, 18) {real, imag} */,
  {32'hc058a193, 32'hc0ee06e8} /* (22, 12, 17) {real, imag} */,
  {32'h4181d1da, 32'hbf8ffef8} /* (22, 12, 16) {real, imag} */,
  {32'hbfc0bd0e, 32'hbedaec00} /* (22, 12, 15) {real, imag} */,
  {32'hc0ad1a2c, 32'h40004bda} /* (22, 12, 14) {real, imag} */,
  {32'h3f3f559c, 32'hc0db704f} /* (22, 12, 13) {real, imag} */,
  {32'hc11357b2, 32'hc0f855cc} /* (22, 12, 12) {real, imag} */,
  {32'h40bba370, 32'h40e759f5} /* (22, 12, 11) {real, imag} */,
  {32'h4090eb62, 32'h40ee7821} /* (22, 12, 10) {real, imag} */,
  {32'h4094bcf0, 32'hc11d2172} /* (22, 12, 9) {real, imag} */,
  {32'h41081732, 32'h40e96110} /* (22, 12, 8) {real, imag} */,
  {32'h418a1e34, 32'h41dbaf9b} /* (22, 12, 7) {real, imag} */,
  {32'hc1a5b2a6, 32'h418536c7} /* (22, 12, 6) {real, imag} */,
  {32'hbfd6db66, 32'h4000ba04} /* (22, 12, 5) {real, imag} */,
  {32'h41e2f5f4, 32'h408c6bc2} /* (22, 12, 4) {real, imag} */,
  {32'hc20fbef4, 32'h418f35f8} /* (22, 12, 3) {real, imag} */,
  {32'h3febff34, 32'h41958b6b} /* (22, 12, 2) {real, imag} */,
  {32'h41a40079, 32'hc0b358f0} /* (22, 12, 1) {real, imag} */,
  {32'h411ba083, 32'hc1e59cc4} /* (22, 12, 0) {real, imag} */,
  {32'hc228fb60, 32'hc1a8bff3} /* (22, 11, 31) {real, imag} */,
  {32'h417f68c4, 32'h4164c3b5} /* (22, 11, 30) {real, imag} */,
  {32'h413bf346, 32'h3fa36810} /* (22, 11, 29) {real, imag} */,
  {32'hc0b7cd2a, 32'hc123cd8b} /* (22, 11, 28) {real, imag} */,
  {32'hc1a61fa1, 32'hc1c05656} /* (22, 11, 27) {real, imag} */,
  {32'h420286c5, 32'hc2308b47} /* (22, 11, 26) {real, imag} */,
  {32'h3fcc0af0, 32'h4110589e} /* (22, 11, 25) {real, imag} */,
  {32'hc0eaf78b, 32'hc20fd5e3} /* (22, 11, 24) {real, imag} */,
  {32'h4200932a, 32'h41ca829d} /* (22, 11, 23) {real, imag} */,
  {32'hc0b1ec64, 32'hbebae660} /* (22, 11, 22) {real, imag} */,
  {32'h419b02a0, 32'hc1753160} /* (22, 11, 21) {real, imag} */,
  {32'hc137a913, 32'hc085ec66} /* (22, 11, 20) {real, imag} */,
  {32'hbea5d608, 32'hc185c4cc} /* (22, 11, 19) {real, imag} */,
  {32'hc1659e50, 32'h4019fef8} /* (22, 11, 18) {real, imag} */,
  {32'h40759a30, 32'hbf172b08} /* (22, 11, 17) {real, imag} */,
  {32'h41179b6c, 32'hc100a64b} /* (22, 11, 16) {real, imag} */,
  {32'hbf4558c0, 32'h40e3815d} /* (22, 11, 15) {real, imag} */,
  {32'hc0f6d778, 32'hc0c31b80} /* (22, 11, 14) {real, imag} */,
  {32'h4103a818, 32'h410ca713} /* (22, 11, 13) {real, imag} */,
  {32'h410a420d, 32'h40b02b94} /* (22, 11, 12) {real, imag} */,
  {32'h410bfd20, 32'hbfe39580} /* (22, 11, 11) {real, imag} */,
  {32'hc0e03904, 32'hc188d374} /* (22, 11, 10) {real, imag} */,
  {32'hc0e4bf68, 32'h4093fa9c} /* (22, 11, 9) {real, imag} */,
  {32'hc0c6b70d, 32'h40fe6d1e} /* (22, 11, 8) {real, imag} */,
  {32'hc1e932df, 32'h41b870d1} /* (22, 11, 7) {real, imag} */,
  {32'hc216e617, 32'h41830648} /* (22, 11, 6) {real, imag} */,
  {32'h414aaec6, 32'hc24c3815} /* (22, 11, 5) {real, imag} */,
  {32'h40ea5390, 32'h4154d069} /* (22, 11, 4) {real, imag} */,
  {32'h41116f16, 32'hc23c75d2} /* (22, 11, 3) {real, imag} */,
  {32'hc1efbda2, 32'h4012548c} /* (22, 11, 2) {real, imag} */,
  {32'h40253cc0, 32'h4178a03e} /* (22, 11, 1) {real, imag} */,
  {32'h4226379a, 32'h4198abee} /* (22, 11, 0) {real, imag} */,
  {32'h41227ac4, 32'hc083080f} /* (22, 10, 31) {real, imag} */,
  {32'hc1ca27ca, 32'hc20a6b11} /* (22, 10, 30) {real, imag} */,
  {32'hc1d6a3d2, 32'hc1ad0527} /* (22, 10, 29) {real, imag} */,
  {32'h419b38c0, 32'hc04a2610} /* (22, 10, 28) {real, imag} */,
  {32'h41a88a70, 32'h3f3c0e40} /* (22, 10, 27) {real, imag} */,
  {32'hc0fbd1f2, 32'h40960560} /* (22, 10, 26) {real, imag} */,
  {32'h407251a8, 32'hc0821f60} /* (22, 10, 25) {real, imag} */,
  {32'h404050fa, 32'h4179c9be} /* (22, 10, 24) {real, imag} */,
  {32'h4100e9fa, 32'h3f84b2c8} /* (22, 10, 23) {real, imag} */,
  {32'h4135e294, 32'h40bd1c6e} /* (22, 10, 22) {real, imag} */,
  {32'hc1a0aec6, 32'h3fed6c10} /* (22, 10, 21) {real, imag} */,
  {32'h4037d92c, 32'h3fb82084} /* (22, 10, 20) {real, imag} */,
  {32'hc1549d3e, 32'h41b858fa} /* (22, 10, 19) {real, imag} */,
  {32'hc0e0668e, 32'h4077f234} /* (22, 10, 18) {real, imag} */,
  {32'hc089b2ad, 32'h40bc4cc4} /* (22, 10, 17) {real, imag} */,
  {32'hc010e1b2, 32'h40a0f098} /* (22, 10, 16) {real, imag} */,
  {32'h3f9c8f74, 32'hc12ea8a6} /* (22, 10, 15) {real, imag} */,
  {32'h412230b9, 32'h408f74ea} /* (22, 10, 14) {real, imag} */,
  {32'hc196542d, 32'hc04dce80} /* (22, 10, 13) {real, imag} */,
  {32'hc1837b70, 32'h3fdd15d4} /* (22, 10, 12) {real, imag} */,
  {32'h3fd1cc18, 32'h4086c524} /* (22, 10, 11) {real, imag} */,
  {32'h40f51834, 32'h41c9d1b4} /* (22, 10, 10) {real, imag} */,
  {32'hc17efbb8, 32'hbf9f8580} /* (22, 10, 9) {real, imag} */,
  {32'hc17861a6, 32'h41da4eef} /* (22, 10, 8) {real, imag} */,
  {32'h412f00f0, 32'hc1e0ba68} /* (22, 10, 7) {real, imag} */,
  {32'hc1d79f00, 32'h424b9820} /* (22, 10, 6) {real, imag} */,
  {32'h40ba0b82, 32'h426301aa} /* (22, 10, 5) {real, imag} */,
  {32'h4124be8e, 32'hc1f03832} /* (22, 10, 4) {real, imag} */,
  {32'hc1d58716, 32'hc03a2c98} /* (22, 10, 3) {real, imag} */,
  {32'h4188fc70, 32'h41baf11e} /* (22, 10, 2) {real, imag} */,
  {32'hc1aa401c, 32'hc1923bb8} /* (22, 10, 1) {real, imag} */,
  {32'h417b6afc, 32'h422e48de} /* (22, 10, 0) {real, imag} */,
  {32'h41e58b09, 32'h4169b678} /* (22, 9, 31) {real, imag} */,
  {32'h421e6e61, 32'h4248d728} /* (22, 9, 30) {real, imag} */,
  {32'h408a22da, 32'hc21a295d} /* (22, 9, 29) {real, imag} */,
  {32'h4244af63, 32'h404d91dc} /* (22, 9, 28) {real, imag} */,
  {32'hc154e379, 32'hc1e5e518} /* (22, 9, 27) {real, imag} */,
  {32'hc1cf7588, 32'h4219b4cf} /* (22, 9, 26) {real, imag} */,
  {32'hc21fd758, 32'hc1a76bf2} /* (22, 9, 25) {real, imag} */,
  {32'h4099ca31, 32'h41b2b346} /* (22, 9, 24) {real, imag} */,
  {32'h41d706c9, 32'h410ab334} /* (22, 9, 23) {real, imag} */,
  {32'hc1cc9cf4, 32'h40e101b4} /* (22, 9, 22) {real, imag} */,
  {32'hc19390bf, 32'hc197d3d6} /* (22, 9, 21) {real, imag} */,
  {32'h41cdac43, 32'h40759b54} /* (22, 9, 20) {real, imag} */,
  {32'h413e552e, 32'h41be84cb} /* (22, 9, 19) {real, imag} */,
  {32'hc0cc26b8, 32'h4090dd18} /* (22, 9, 18) {real, imag} */,
  {32'h40b4c529, 32'h40e8bb28} /* (22, 9, 17) {real, imag} */,
  {32'h40e52336, 32'hc10cafe9} /* (22, 9, 16) {real, imag} */,
  {32'h41266638, 32'hc0e745e4} /* (22, 9, 15) {real, imag} */,
  {32'h419f8373, 32'h3f0ca400} /* (22, 9, 14) {real, imag} */,
  {32'hc06eda32, 32'hbf81d470} /* (22, 9, 13) {real, imag} */,
  {32'h411212c2, 32'h420b7dc5} /* (22, 9, 12) {real, imag} */,
  {32'h41eb6f85, 32'h3fbfac68} /* (22, 9, 11) {real, imag} */,
  {32'h414c4127, 32'hc1d640dd} /* (22, 9, 10) {real, imag} */,
  {32'hc25090f2, 32'hbe4fa5a0} /* (22, 9, 9) {real, imag} */,
  {32'hc0a4e08f, 32'hc1163a39} /* (22, 9, 8) {real, imag} */,
  {32'h414ecb8c, 32'h41d8d31a} /* (22, 9, 7) {real, imag} */,
  {32'h4235a9b0, 32'h4098b3a0} /* (22, 9, 6) {real, imag} */,
  {32'hc1bd633c, 32'h4209aa56} /* (22, 9, 5) {real, imag} */,
  {32'hc1edda62, 32'h41d8ab08} /* (22, 9, 4) {real, imag} */,
  {32'h41a52384, 32'hc1b8906a} /* (22, 9, 3) {real, imag} */,
  {32'hc227b23f, 32'hc17f4592} /* (22, 9, 2) {real, imag} */,
  {32'h40ac9fb4, 32'hc253d168} /* (22, 9, 1) {real, imag} */,
  {32'hbff2be90, 32'h41468033} /* (22, 9, 0) {real, imag} */,
  {32'hbfebf4a0, 32'h421143e8} /* (22, 8, 31) {real, imag} */,
  {32'h41266b40, 32'hc1d27dae} /* (22, 8, 30) {real, imag} */,
  {32'h418a8b56, 32'hc280052c} /* (22, 8, 29) {real, imag} */,
  {32'h40f3133c, 32'h422d2c96} /* (22, 8, 28) {real, imag} */,
  {32'hc18f2a20, 32'h422bc408} /* (22, 8, 27) {real, imag} */,
  {32'hc2536134, 32'hc216b73a} /* (22, 8, 26) {real, imag} */,
  {32'h3e5e3400, 32'hc121a660} /* (22, 8, 25) {real, imag} */,
  {32'h4117813c, 32'h403ccafb} /* (22, 8, 24) {real, imag} */,
  {32'h40bc943a, 32'hc14ceed8} /* (22, 8, 23) {real, imag} */,
  {32'hc0ea010a, 32'h41101bff} /* (22, 8, 22) {real, imag} */,
  {32'h403c88c4, 32'hc00c8cb4} /* (22, 8, 21) {real, imag} */,
  {32'hc2165568, 32'hc1105d17} /* (22, 8, 20) {real, imag} */,
  {32'hc12d6e2a, 32'hc0807172} /* (22, 8, 19) {real, imag} */,
  {32'h41017004, 32'hbff0cb60} /* (22, 8, 18) {real, imag} */,
  {32'hc1eb0244, 32'h3e3ab2e0} /* (22, 8, 17) {real, imag} */,
  {32'h401ed296, 32'hbf862108} /* (22, 8, 16) {real, imag} */,
  {32'h4207ddd4, 32'hc0c8622d} /* (22, 8, 15) {real, imag} */,
  {32'h410913e0, 32'h40a108b4} /* (22, 8, 14) {real, imag} */,
  {32'hc078ccaf, 32'h4135d143} /* (22, 8, 13) {real, imag} */,
  {32'h4184fdba, 32'h41cd0b68} /* (22, 8, 12) {real, imag} */,
  {32'hc09d6abe, 32'h4171ab8b} /* (22, 8, 11) {real, imag} */,
  {32'hc166f717, 32'hc1d52a12} /* (22, 8, 10) {real, imag} */,
  {32'h410e9d32, 32'hc1827a0d} /* (22, 8, 9) {real, imag} */,
  {32'hc135d876, 32'hbf24e194} /* (22, 8, 8) {real, imag} */,
  {32'hc2069d96, 32'h4237e284} /* (22, 8, 7) {real, imag} */,
  {32'hc2a7bb70, 32'h4058eec8} /* (22, 8, 6) {real, imag} */,
  {32'h4293e828, 32'hc2705e24} /* (22, 8, 5) {real, imag} */,
  {32'hc129b966, 32'hc221b7f8} /* (22, 8, 4) {real, imag} */,
  {32'h419c2d02, 32'h428a0e88} /* (22, 8, 3) {real, imag} */,
  {32'hc1f399ba, 32'hc220904d} /* (22, 8, 2) {real, imag} */,
  {32'h4234157d, 32'hc16fd780} /* (22, 8, 1) {real, imag} */,
  {32'hc08aa7dd, 32'hc1495477} /* (22, 8, 0) {real, imag} */,
  {32'hc1c8a368, 32'hc1bbfad2} /* (22, 7, 31) {real, imag} */,
  {32'hc1fd016d, 32'h428808d9} /* (22, 7, 30) {real, imag} */,
  {32'hc27be6ed, 32'h426c2633} /* (22, 7, 29) {real, imag} */,
  {32'h41cf448f, 32'h400d63a8} /* (22, 7, 28) {real, imag} */,
  {32'h4250c816, 32'h428113f2} /* (22, 7, 27) {real, imag} */,
  {32'hc280e30f, 32'h416ccac8} /* (22, 7, 26) {real, imag} */,
  {32'hc1a9c7a2, 32'hc23759ce} /* (22, 7, 25) {real, imag} */,
  {32'h41663495, 32'h410b15b4} /* (22, 7, 24) {real, imag} */,
  {32'hc0955cd2, 32'hc1271a96} /* (22, 7, 23) {real, imag} */,
  {32'h41484413, 32'h420c0556} /* (22, 7, 22) {real, imag} */,
  {32'hc1332e9f, 32'hc1b2af5c} /* (22, 7, 21) {real, imag} */,
  {32'hc159ab76, 32'h406916a2} /* (22, 7, 20) {real, imag} */,
  {32'hc1e8ef78, 32'h40a66aa2} /* (22, 7, 19) {real, imag} */,
  {32'h40b925ac, 32'hc03d1798} /* (22, 7, 18) {real, imag} */,
  {32'hc0220b74, 32'hbecfe2c0} /* (22, 7, 17) {real, imag} */,
  {32'hc11f2129, 32'h40d1f640} /* (22, 7, 16) {real, imag} */,
  {32'h4088ca16, 32'h419607ab} /* (22, 7, 15) {real, imag} */,
  {32'h3feb06d0, 32'hc1943d1b} /* (22, 7, 14) {real, imag} */,
  {32'hc13aade8, 32'hc13123f9} /* (22, 7, 13) {real, imag} */,
  {32'h411a7ab6, 32'hc137e46c} /* (22, 7, 12) {real, imag} */,
  {32'hc17b46f9, 32'hc17119fc} /* (22, 7, 11) {real, imag} */,
  {32'hc205753b, 32'hc2009b0c} /* (22, 7, 10) {real, imag} */,
  {32'hbf19e270, 32'h423410f4} /* (22, 7, 9) {real, imag} */,
  {32'hc1bab13e, 32'h40f8c448} /* (22, 7, 8) {real, imag} */,
  {32'h401274dc, 32'hc25a80bc} /* (22, 7, 7) {real, imag} */,
  {32'h4274b02a, 32'h42688172} /* (22, 7, 6) {real, imag} */,
  {32'h4280e2c2, 32'hc1c1fb37} /* (22, 7, 5) {real, imag} */,
  {32'h40cdf324, 32'hc1dd2a7f} /* (22, 7, 4) {real, imag} */,
  {32'h427011d1, 32'h41917bb6} /* (22, 7, 3) {real, imag} */,
  {32'h41c91b39, 32'hc18ff699} /* (22, 7, 2) {real, imag} */,
  {32'h42818608, 32'h427eb097} /* (22, 7, 1) {real, imag} */,
  {32'hc1cdfe28, 32'hc20326d4} /* (22, 7, 0) {real, imag} */,
  {32'h418f8319, 32'h410b5302} /* (22, 6, 31) {real, imag} */,
  {32'h414e1008, 32'h407c9ed8} /* (22, 6, 30) {real, imag} */,
  {32'h42ad9b34, 32'hc150e2ba} /* (22, 6, 29) {real, imag} */,
  {32'hc2ab636c, 32'hc18140a2} /* (22, 6, 28) {real, imag} */,
  {32'hc25e5a24, 32'h42993b8c} /* (22, 6, 27) {real, imag} */,
  {32'h40320b88, 32'hbfae6fc0} /* (22, 6, 26) {real, imag} */,
  {32'h428cb446, 32'h4219968e} /* (22, 6, 25) {real, imag} */,
  {32'hc127e4bb, 32'hc17d9855} /* (22, 6, 24) {real, imag} */,
  {32'hc047b83c, 32'hc095e557} /* (22, 6, 23) {real, imag} */,
  {32'h413c70d9, 32'hc1b8d3f1} /* (22, 6, 22) {real, imag} */,
  {32'hbfb8a3b8, 32'hc2069e3e} /* (22, 6, 21) {real, imag} */,
  {32'h41a40041, 32'hc05a6e90} /* (22, 6, 20) {real, imag} */,
  {32'h41319e68, 32'hc06b8800} /* (22, 6, 19) {real, imag} */,
  {32'hc0819dce, 32'h41588b88} /* (22, 6, 18) {real, imag} */,
  {32'hc12b4642, 32'h3f3edc58} /* (22, 6, 17) {real, imag} */,
  {32'hc055a100, 32'h402635c0} /* (22, 6, 16) {real, imag} */,
  {32'h4180adb7, 32'hc07cc022} /* (22, 6, 15) {real, imag} */,
  {32'hc12be22f, 32'hc0a89990} /* (22, 6, 14) {real, imag} */,
  {32'h4222c31a, 32'h41819602} /* (22, 6, 13) {real, imag} */,
  {32'h411c6ce2, 32'h422e1455} /* (22, 6, 12) {real, imag} */,
  {32'h40e58646, 32'h42031486} /* (22, 6, 11) {real, imag} */,
  {32'h4195909e, 32'hc1b640c7} /* (22, 6, 10) {real, imag} */,
  {32'hc097512a, 32'h40ee94af} /* (22, 6, 9) {real, imag} */,
  {32'h4228b453, 32'hc0774134} /* (22, 6, 8) {real, imag} */,
  {32'h415b27b0, 32'h40efcf9c} /* (22, 6, 7) {real, imag} */,
  {32'h422436d6, 32'hc203405a} /* (22, 6, 6) {real, imag} */,
  {32'hc29bb504, 32'h40b5aec8} /* (22, 6, 5) {real, imag} */,
  {32'hc1036a54, 32'hc1a0c17a} /* (22, 6, 4) {real, imag} */,
  {32'hc0d54788, 32'hc26c1de2} /* (22, 6, 3) {real, imag} */,
  {32'hc29951e6, 32'h422b3936} /* (22, 6, 2) {real, imag} */,
  {32'h4024a368, 32'hc1adbfa8} /* (22, 6, 1) {real, imag} */,
  {32'h426622be, 32'h42549026} /* (22, 6, 0) {real, imag} */,
  {32'h41bf4150, 32'hc27353e0} /* (22, 5, 31) {real, imag} */,
  {32'h3fc69f80, 32'h41cd49c1} /* (22, 5, 30) {real, imag} */,
  {32'h41975872, 32'h426c5661} /* (22, 5, 29) {real, imag} */,
  {32'hc2cf66b6, 32'h4165a3f2} /* (22, 5, 28) {real, imag} */,
  {32'h429e3c7a, 32'h41babc1a} /* (22, 5, 27) {real, imag} */,
  {32'h42016403, 32'hc2820b25} /* (22, 5, 26) {real, imag} */,
  {32'h4172ac28, 32'hc1c6759b} /* (22, 5, 25) {real, imag} */,
  {32'hc200d7e2, 32'hc13ba771} /* (22, 5, 24) {real, imag} */,
  {32'hc062b688, 32'hc1a34629} /* (22, 5, 23) {real, imag} */,
  {32'h414d6c8c, 32'h424df6dc} /* (22, 5, 22) {real, imag} */,
  {32'h412179de, 32'h41919650} /* (22, 5, 21) {real, imag} */,
  {32'hc0bf2380, 32'h41ad2a5c} /* (22, 5, 20) {real, imag} */,
  {32'h40a3c98e, 32'hc05bd284} /* (22, 5, 19) {real, imag} */,
  {32'h41d98920, 32'h3ffd8f84} /* (22, 5, 18) {real, imag} */,
  {32'h40948c55, 32'h3e12c800} /* (22, 5, 17) {real, imag} */,
  {32'hc1c94a8b, 32'hc0eabda8} /* (22, 5, 16) {real, imag} */,
  {32'hbffb8d8c, 32'hc0ac3908} /* (22, 5, 15) {real, imag} */,
  {32'h410992b8, 32'hc130bff0} /* (22, 5, 14) {real, imag} */,
  {32'hc0153414, 32'hc0e5d4f6} /* (22, 5, 13) {real, imag} */,
  {32'h40aaeef0, 32'hc134a39c} /* (22, 5, 12) {real, imag} */,
  {32'h41e13377, 32'h412f26bb} /* (22, 5, 11) {real, imag} */,
  {32'hc221da78, 32'hc09fb594} /* (22, 5, 10) {real, imag} */,
  {32'h41ae0453, 32'h41dc963b} /* (22, 5, 9) {real, imag} */,
  {32'hbfd0f010, 32'h40e883e6} /* (22, 5, 8) {real, imag} */,
  {32'hc10121ec, 32'hc20419a2} /* (22, 5, 7) {real, imag} */,
  {32'hc1fbc0e4, 32'h42311268} /* (22, 5, 6) {real, imag} */,
  {32'h4121c9e4, 32'hc24e569f} /* (22, 5, 5) {real, imag} */,
  {32'h42563ccc, 32'h427c0e48} /* (22, 5, 4) {real, imag} */,
  {32'hc28818f6, 32'h42370d73} /* (22, 5, 3) {real, imag} */,
  {32'hc21a64be, 32'hc1123346} /* (22, 5, 2) {real, imag} */,
  {32'hc24cc130, 32'h410ce612} /* (22, 5, 1) {real, imag} */,
  {32'h4240eb7e, 32'hc22b54a1} /* (22, 5, 0) {real, imag} */,
  {32'h421bb8d1, 32'h41bb132e} /* (22, 4, 31) {real, imag} */,
  {32'h40cfffe8, 32'h42815614} /* (22, 4, 30) {real, imag} */,
  {32'hc26abdc2, 32'h4287f844} /* (22, 4, 29) {real, imag} */,
  {32'h40786880, 32'hc2a18ca5} /* (22, 4, 28) {real, imag} */,
  {32'hc1f209fd, 32'h4191dc07} /* (22, 4, 27) {real, imag} */,
  {32'hc2a03e08, 32'hc2b008b6} /* (22, 4, 26) {real, imag} */,
  {32'h4201a66b, 32'hc1fb6d24} /* (22, 4, 25) {real, imag} */,
  {32'h41ced19a, 32'h40598094} /* (22, 4, 24) {real, imag} */,
  {32'hc2260ca4, 32'h414620e5} /* (22, 4, 23) {real, imag} */,
  {32'hc04a7460, 32'h422a15e2} /* (22, 4, 22) {real, imag} */,
  {32'h42690be6, 32'h408dc4b2} /* (22, 4, 21) {real, imag} */,
  {32'hc28f32ac, 32'hc217e472} /* (22, 4, 20) {real, imag} */,
  {32'h418153a6, 32'hc0286184} /* (22, 4, 19) {real, imag} */,
  {32'hc180da32, 32'hc1383dd8} /* (22, 4, 18) {real, imag} */,
  {32'h4132ef93, 32'hc183f170} /* (22, 4, 17) {real, imag} */,
  {32'hc12d8ecd, 32'h40ccdb78} /* (22, 4, 16) {real, imag} */,
  {32'h4111c835, 32'h4073593e} /* (22, 4, 15) {real, imag} */,
  {32'hc19af0fe, 32'hc147c150} /* (22, 4, 14) {real, imag} */,
  {32'h4130b353, 32'hc10d9925} /* (22, 4, 13) {real, imag} */,
  {32'hc1892b08, 32'h4136c00e} /* (22, 4, 12) {real, imag} */,
  {32'h40b9f5f4, 32'hc16d19c7} /* (22, 4, 11) {real, imag} */,
  {32'h3eadaf80, 32'h41fdbf71} /* (22, 4, 10) {real, imag} */,
  {32'h3fa8ab90, 32'h4200aa9f} /* (22, 4, 9) {real, imag} */,
  {32'h42267643, 32'hc1c1a2aa} /* (22, 4, 8) {real, imag} */,
  {32'h422181dd, 32'hc22dfb74} /* (22, 4, 7) {real, imag} */,
  {32'hbf782b00, 32'h4021a7f0} /* (22, 4, 6) {real, imag} */,
  {32'h40aa4924, 32'h42487ac2} /* (22, 4, 5) {real, imag} */,
  {32'hc3229947, 32'hc01dc0e0} /* (22, 4, 4) {real, imag} */,
  {32'h3f95b9c0, 32'hc1c25e72} /* (22, 4, 3) {real, imag} */,
  {32'hc247f9a3, 32'h429742a8} /* (22, 4, 2) {real, imag} */,
  {32'h41bed296, 32'hc25a4c6d} /* (22, 4, 1) {real, imag} */,
  {32'hc15a6e33, 32'hc22fd733} /* (22, 4, 0) {real, imag} */,
  {32'hc2d17e2b, 32'h426a49c3} /* (22, 3, 31) {real, imag} */,
  {32'hc205a4fb, 32'h42c87cef} /* (22, 3, 30) {real, imag} */,
  {32'hc0dee60c, 32'hc1b27a50} /* (22, 3, 29) {real, imag} */,
  {32'h42216f78, 32'h41d107bc} /* (22, 3, 28) {real, imag} */,
  {32'h420b3df4, 32'h42465ae2} /* (22, 3, 27) {real, imag} */,
  {32'h40da5dfa, 32'hc1c9d220} /* (22, 3, 26) {real, imag} */,
  {32'hc10c9c33, 32'hc19c701a} /* (22, 3, 25) {real, imag} */,
  {32'h40e69854, 32'hc2bcca7c} /* (22, 3, 24) {real, imag} */,
  {32'h41d70ba4, 32'hc06f6330} /* (22, 3, 23) {real, imag} */,
  {32'hc27f76ff, 32'hc1cdf09f} /* (22, 3, 22) {real, imag} */,
  {32'hc1a1ec9e, 32'hc1164dd2} /* (22, 3, 21) {real, imag} */,
  {32'h410aa546, 32'hc21268a5} /* (22, 3, 20) {real, imag} */,
  {32'hc0f04eee, 32'hc165f3eb} /* (22, 3, 19) {real, imag} */,
  {32'hc126e4c9, 32'hc20b50fe} /* (22, 3, 18) {real, imag} */,
  {32'h3e8f32a0, 32'h41405c78} /* (22, 3, 17) {real, imag} */,
  {32'h419f3a50, 32'h418687ae} /* (22, 3, 16) {real, imag} */,
  {32'h4110bb2b, 32'hc0c980e0} /* (22, 3, 15) {real, imag} */,
  {32'hc13b48bf, 32'h41ecd170} /* (22, 3, 14) {real, imag} */,
  {32'hc181bb5a, 32'h40ee7bda} /* (22, 3, 13) {real, imag} */,
  {32'h4226126a, 32'h40a6b94a} /* (22, 3, 12) {real, imag} */,
  {32'hc1a9b5ee, 32'h410841ae} /* (22, 3, 11) {real, imag} */,
  {32'hc0398b10, 32'h417bff1a} /* (22, 3, 10) {real, imag} */,
  {32'h41d6f078, 32'hc1c0e668} /* (22, 3, 9) {real, imag} */,
  {32'hc1a6dbd1, 32'h412751c4} /* (22, 3, 8) {real, imag} */,
  {32'hc2053ce7, 32'h418b72f0} /* (22, 3, 7) {real, imag} */,
  {32'h418b71c2, 32'hc2bbf80a} /* (22, 3, 6) {real, imag} */,
  {32'hc20c7488, 32'hc2b0def3} /* (22, 3, 5) {real, imag} */,
  {32'hc1ad4735, 32'hc119f237} /* (22, 3, 4) {real, imag} */,
  {32'hc257537a, 32'h4094999e} /* (22, 3, 3) {real, imag} */,
  {32'hc1a002b6, 32'h4256a662} /* (22, 3, 2) {real, imag} */,
  {32'hc28f24e1, 32'h4277d3e3} /* (22, 3, 1) {real, imag} */,
  {32'hc28a40c4, 32'h42c3f51c} /* (22, 3, 0) {real, imag} */,
  {32'h4285900f, 32'h42b98747} /* (22, 2, 31) {real, imag} */,
  {32'hc11a1328, 32'h41616339} /* (22, 2, 30) {real, imag} */,
  {32'h42da1d30, 32'h40c68f20} /* (22, 2, 29) {real, imag} */,
  {32'h418a9b63, 32'hc33cd1b3} /* (22, 2, 28) {real, imag} */,
  {32'hc0a96db8, 32'hc27bef32} /* (22, 2, 27) {real, imag} */,
  {32'h4205d68e, 32'h42286cb6} /* (22, 2, 26) {real, imag} */,
  {32'hc11aaffe, 32'hc2286028} /* (22, 2, 25) {real, imag} */,
  {32'hc27acf2e, 32'hc1e52baa} /* (22, 2, 24) {real, imag} */,
  {32'hc207b34b, 32'h40298230} /* (22, 2, 23) {real, imag} */,
  {32'h40966752, 32'hc0f9ca18} /* (22, 2, 22) {real, imag} */,
  {32'hc0dc41ec, 32'h4068b10e} /* (22, 2, 21) {real, imag} */,
  {32'hc1b5faf1, 32'h42157f50} /* (22, 2, 20) {real, imag} */,
  {32'h410b5a02, 32'h416836b6} /* (22, 2, 19) {real, imag} */,
  {32'h416aa472, 32'h41f2a8be} /* (22, 2, 18) {real, imag} */,
  {32'hc1369048, 32'h40b380ae} /* (22, 2, 17) {real, imag} */,
  {32'h40b1be10, 32'hbe816c40} /* (22, 2, 16) {real, imag} */,
  {32'h40699422, 32'h41017a3f} /* (22, 2, 15) {real, imag} */,
  {32'h42084250, 32'hc1d1461e} /* (22, 2, 14) {real, imag} */,
  {32'h40f556f4, 32'hc1ed3bb7} /* (22, 2, 13) {real, imag} */,
  {32'hc1a983d5, 32'hc1d241f5} /* (22, 2, 12) {real, imag} */,
  {32'hc001d6a8, 32'h4182f820} /* (22, 2, 11) {real, imag} */,
  {32'hc182ab2e, 32'h422285d2} /* (22, 2, 10) {real, imag} */,
  {32'hc1d77a06, 32'hc19f8722} /* (22, 2, 9) {real, imag} */,
  {32'hc232472e, 32'hc2b6dbda} /* (22, 2, 8) {real, imag} */,
  {32'h40ea310c, 32'h42847d0a} /* (22, 2, 7) {real, imag} */,
  {32'h40f5ad84, 32'hc1c53d9c} /* (22, 2, 6) {real, imag} */,
  {32'hc2a2d138, 32'hc22ffe4e} /* (22, 2, 5) {real, imag} */,
  {32'h41189127, 32'h4271f38c} /* (22, 2, 4) {real, imag} */,
  {32'hc157b53c, 32'h42b74786} /* (22, 2, 3) {real, imag} */,
  {32'hc3260cb8, 32'h40e2e706} /* (22, 2, 2) {real, imag} */,
  {32'h42072cea, 32'hc29b8ce5} /* (22, 2, 1) {real, imag} */,
  {32'h431715d0, 32'h41fb8353} /* (22, 2, 0) {real, imag} */,
  {32'hc2be1d16, 32'hc22c2e28} /* (22, 1, 31) {real, imag} */,
  {32'h42926038, 32'h42d43dec} /* (22, 1, 30) {real, imag} */,
  {32'h41e55c78, 32'hc2c69876} /* (22, 1, 29) {real, imag} */,
  {32'hc222c9c2, 32'hbf37d198} /* (22, 1, 28) {real, imag} */,
  {32'hc1c2b6cc, 32'h4322a7d2} /* (22, 1, 27) {real, imag} */,
  {32'hc1afd438, 32'h424011cf} /* (22, 1, 26) {real, imag} */,
  {32'hc1ce67d0, 32'hc21863fd} /* (22, 1, 25) {real, imag} */,
  {32'hc104b678, 32'h426b227a} /* (22, 1, 24) {real, imag} */,
  {32'h417bf7f6, 32'hc0eca9d6} /* (22, 1, 23) {real, imag} */,
  {32'h41e28d7c, 32'h41b8c6da} /* (22, 1, 22) {real, imag} */,
  {32'h4115c1c2, 32'hc10a3ecc} /* (22, 1, 21) {real, imag} */,
  {32'h3feb7df8, 32'h40f53a61} /* (22, 1, 20) {real, imag} */,
  {32'h41ed6f72, 32'h421eb2ec} /* (22, 1, 19) {real, imag} */,
  {32'hc0e4c852, 32'hc10586bc} /* (22, 1, 18) {real, imag} */,
  {32'hc1334ea9, 32'hc1ac96c4} /* (22, 1, 17) {real, imag} */,
  {32'h40f7de74, 32'h4000c740} /* (22, 1, 16) {real, imag} */,
  {32'h41563381, 32'h412da518} /* (22, 1, 15) {real, imag} */,
  {32'hc16f7e37, 32'hc129fa84} /* (22, 1, 14) {real, imag} */,
  {32'hc10df20c, 32'hc0b2cb4c} /* (22, 1, 13) {real, imag} */,
  {32'hc195b554, 32'hbfc3f204} /* (22, 1, 12) {real, imag} */,
  {32'h4102383a, 32'hc1e15c8e} /* (22, 1, 11) {real, imag} */,
  {32'h4107f248, 32'h41ee0a9a} /* (22, 1, 10) {real, imag} */,
  {32'hc288d1cb, 32'hc1c0117e} /* (22, 1, 9) {real, imag} */,
  {32'hc19d3590, 32'hc1f143c3} /* (22, 1, 8) {real, imag} */,
  {32'h40f7a0c8, 32'hc2cc1d16} /* (22, 1, 7) {real, imag} */,
  {32'h42209580, 32'h4201f27f} /* (22, 1, 6) {real, imag} */,
  {32'h430e4902, 32'h4233531a} /* (22, 1, 5) {real, imag} */,
  {32'hc22c0f48, 32'hc183e2a7} /* (22, 1, 4) {real, imag} */,
  {32'h430b1f1f, 32'h3ed19380} /* (22, 1, 3) {real, imag} */,
  {32'h41fbf3a8, 32'h42bb3bc0} /* (22, 1, 2) {real, imag} */,
  {32'hc28184be, 32'hc30a33cf} /* (22, 1, 1) {real, imag} */,
  {32'h428004c0, 32'hc31b0ef1} /* (22, 1, 0) {real, imag} */,
  {32'hc2d0398b, 32'h42cd5d5d} /* (22, 0, 31) {real, imag} */,
  {32'h4245643a, 32'h42a97762} /* (22, 0, 30) {real, imag} */,
  {32'hc30bdca4, 32'h410150be} /* (22, 0, 29) {real, imag} */,
  {32'hc124af6c, 32'hbf3be1c0} /* (22, 0, 28) {real, imag} */,
  {32'hc1c942b4, 32'hc2848356} /* (22, 0, 27) {real, imag} */,
  {32'h4136cb56, 32'hc0892ba0} /* (22, 0, 26) {real, imag} */,
  {32'hc23dd76f, 32'hc2a52804} /* (22, 0, 25) {real, imag} */,
  {32'hc2a0d834, 32'hc22a0aea} /* (22, 0, 24) {real, imag} */,
  {32'h4276b903, 32'hc268c0b0} /* (22, 0, 23) {real, imag} */,
  {32'hc0baed68, 32'hc0f1fe00} /* (22, 0, 22) {real, imag} */,
  {32'hc03e5118, 32'h4238861b} /* (22, 0, 21) {real, imag} */,
  {32'h408af9cc, 32'h419ba2e5} /* (22, 0, 20) {real, imag} */,
  {32'h408df0e6, 32'hc204f45e} /* (22, 0, 19) {real, imag} */,
  {32'hc0ea7b9c, 32'h419316d9} /* (22, 0, 18) {real, imag} */,
  {32'h413484f6, 32'hc12d7a99} /* (22, 0, 17) {real, imag} */,
  {32'h41a17744, 32'hc2255080} /* (22, 0, 16) {real, imag} */,
  {32'h40d307f4, 32'h41b31c8c} /* (22, 0, 15) {real, imag} */,
  {32'hc10b6aa6, 32'h40826d8c} /* (22, 0, 14) {real, imag} */,
  {32'hc1af0d72, 32'h41e22765} /* (22, 0, 13) {real, imag} */,
  {32'h420a140a, 32'hc0d3bc64} /* (22, 0, 12) {real, imag} */,
  {32'h42036ea2, 32'h41b2d6fa} /* (22, 0, 11) {real, imag} */,
  {32'hc16dab10, 32'hc1ebb2a8} /* (22, 0, 10) {real, imag} */,
  {32'h42bc53c4, 32'h413c7650} /* (22, 0, 9) {real, imag} */,
  {32'hc17ffca0, 32'hc1a35fee} /* (22, 0, 8) {real, imag} */,
  {32'h41d0ade6, 32'h4197bf08} /* (22, 0, 7) {real, imag} */,
  {32'hc2671a2e, 32'h42f255a4} /* (22, 0, 6) {real, imag} */,
  {32'h432d08a2, 32'h428add02} /* (22, 0, 5) {real, imag} */,
  {32'h42c040b0, 32'h42e1f3ea} /* (22, 0, 4) {real, imag} */,
  {32'hc29b8a06, 32'h42521834} /* (22, 0, 3) {real, imag} */,
  {32'hc0c18e54, 32'h41d2c85d} /* (22, 0, 2) {real, imag} */,
  {32'hc2264fce, 32'hc1e251b4} /* (22, 0, 1) {real, imag} */,
  {32'hc214a857, 32'h4212cb0c} /* (22, 0, 0) {real, imag} */,
  {32'h4389bb5d, 32'hc1e41548} /* (21, 31, 31) {real, imag} */,
  {32'hc34201bd, 32'h426675ab} /* (21, 31, 30) {real, imag} */,
  {32'h427c7ae7, 32'hc1afc416} /* (21, 31, 29) {real, imag} */,
  {32'h420b311e, 32'hc22c1d86} /* (21, 31, 28) {real, imag} */,
  {32'hc28da48c, 32'hc1fb3658} /* (21, 31, 27) {real, imag} */,
  {32'h42871bb1, 32'h41802080} /* (21, 31, 26) {real, imag} */,
  {32'hc2082297, 32'h41d363dd} /* (21, 31, 25) {real, imag} */,
  {32'hc29fe38e, 32'hc21ae5f3} /* (21, 31, 24) {real, imag} */,
  {32'h42399589, 32'h41afd4ff} /* (21, 31, 23) {real, imag} */,
  {32'hbf7d0720, 32'hc1325f2e} /* (21, 31, 22) {real, imag} */,
  {32'hc1ac187a, 32'h40301426} /* (21, 31, 21) {real, imag} */,
  {32'hc062a4f2, 32'hc1961b9e} /* (21, 31, 20) {real, imag} */,
  {32'h41859e02, 32'h41030fb2} /* (21, 31, 19) {real, imag} */,
  {32'h42368971, 32'h419a161d} /* (21, 31, 18) {real, imag} */,
  {32'hc0109d80, 32'hc1a39d51} /* (21, 31, 17) {real, imag} */,
  {32'hc0a58fc0, 32'h413d3a0c} /* (21, 31, 16) {real, imag} */,
  {32'h41f35378, 32'h41b4b4e9} /* (21, 31, 15) {real, imag} */,
  {32'hbff87520, 32'h401077d0} /* (21, 31, 14) {real, imag} */,
  {32'h40eed132, 32'h41ee6321} /* (21, 31, 13) {real, imag} */,
  {32'h41249b5c, 32'hc223fddc} /* (21, 31, 12) {real, imag} */,
  {32'hc0d453d8, 32'h40fa42dd} /* (21, 31, 11) {real, imag} */,
  {32'hc1016f1a, 32'h41f89d11} /* (21, 31, 10) {real, imag} */,
  {32'hc09839b0, 32'h41711b6a} /* (21, 31, 9) {real, imag} */,
  {32'h41d3ef76, 32'h42b8ce42} /* (21, 31, 8) {real, imag} */,
  {32'hc18e04c8, 32'h424927b0} /* (21, 31, 7) {real, imag} */,
  {32'hc25c4764, 32'hc15d06a0} /* (21, 31, 6) {real, imag} */,
  {32'hc2f962e4, 32'hc26499ec} /* (21, 31, 5) {real, imag} */,
  {32'h424e8862, 32'hc2fab04b} /* (21, 31, 4) {real, imag} */,
  {32'hc121a5a4, 32'hc23bdbe9} /* (21, 31, 3) {real, imag} */,
  {32'hc2e804b2, 32'h413335a4} /* (21, 31, 2) {real, imag} */,
  {32'h4212ec4a, 32'h42b65580} /* (21, 31, 1) {real, imag} */,
  {32'h432ee17c, 32'h420d67ab} /* (21, 31, 0) {real, imag} */,
  {32'hc231cdd4, 32'hc1fb0054} /* (21, 30, 31) {real, imag} */,
  {32'h41935ba4, 32'h430d5ed0} /* (21, 30, 30) {real, imag} */,
  {32'hc1d02ca9, 32'h3f9f7e3c} /* (21, 30, 29) {real, imag} */,
  {32'hc24dcc10, 32'h4213aef0} /* (21, 30, 28) {real, imag} */,
  {32'h425cdd95, 32'hc14addb5} /* (21, 30, 27) {real, imag} */,
  {32'h41a9a00f, 32'h4235bbba} /* (21, 30, 26) {real, imag} */,
  {32'h41dc593f, 32'hc1dd1c48} /* (21, 30, 25) {real, imag} */,
  {32'hc1b62dc8, 32'hc28a358c} /* (21, 30, 24) {real, imag} */,
  {32'hc210f68e, 32'h423614c6} /* (21, 30, 23) {real, imag} */,
  {32'hc298d298, 32'h40fb2f20} /* (21, 30, 22) {real, imag} */,
  {32'h41da163a, 32'hc2274829} /* (21, 30, 21) {real, imag} */,
  {32'h425e4fb8, 32'hc01d8eb8} /* (21, 30, 20) {real, imag} */,
  {32'hc198eb9e, 32'h40d3e1b7} /* (21, 30, 19) {real, imag} */,
  {32'hc1a0dfcc, 32'h406b7b08} /* (21, 30, 18) {real, imag} */,
  {32'h410c3aec, 32'h41f07907} /* (21, 30, 17) {real, imag} */,
  {32'h3cfc7000, 32'hc110b940} /* (21, 30, 16) {real, imag} */,
  {32'hc07a2250, 32'hc1bfc457} /* (21, 30, 15) {real, imag} */,
  {32'hc1164ff8, 32'hc0205408} /* (21, 30, 14) {real, imag} */,
  {32'h419c9836, 32'hc0a8b91f} /* (21, 30, 13) {real, imag} */,
  {32'hc16f5f7e, 32'hc1ccaec0} /* (21, 30, 12) {real, imag} */,
  {32'h405df680, 32'h4164617d} /* (21, 30, 11) {real, imag} */,
  {32'h40cd9ce0, 32'hc195fafc} /* (21, 30, 10) {real, imag} */,
  {32'h424b74f4, 32'hc064d758} /* (21, 30, 9) {real, imag} */,
  {32'h41230510, 32'h428b3c92} /* (21, 30, 8) {real, imag} */,
  {32'hc268fc3e, 32'hc2c469b6} /* (21, 30, 7) {real, imag} */,
  {32'h41809e13, 32'hc23d9c0a} /* (21, 30, 6) {real, imag} */,
  {32'hc08da410, 32'hc18e3108} /* (21, 30, 5) {real, imag} */,
  {32'h4167d2fe, 32'h40a60dde} /* (21, 30, 4) {real, imag} */,
  {32'h40e7fe3c, 32'h3f710e08} /* (21, 30, 3) {real, imag} */,
  {32'h432e0860, 32'h411b6c78} /* (21, 30, 2) {real, imag} */,
  {32'hc33c3263, 32'hc2d1bb7f} /* (21, 30, 1) {real, imag} */,
  {32'hc2c2e52d, 32'hc0bf8a2d} /* (21, 30, 0) {real, imag} */,
  {32'hc1d1ad44, 32'hc23b4e40} /* (21, 29, 31) {real, imag} */,
  {32'hc2cf1c44, 32'h405ad770} /* (21, 29, 30) {real, imag} */,
  {32'hc2a4247b, 32'h422d38b8} /* (21, 29, 29) {real, imag} */,
  {32'hc1def8d5, 32'hc1ca4bc5} /* (21, 29, 28) {real, imag} */,
  {32'hc1855296, 32'h41a6675e} /* (21, 29, 27) {real, imag} */,
  {32'h41a3589c, 32'h41c78f07} /* (21, 29, 26) {real, imag} */,
  {32'h41b7b6b3, 32'hc03d0ca0} /* (21, 29, 25) {real, imag} */,
  {32'hc1a04f96, 32'hc2465aa8} /* (21, 29, 24) {real, imag} */,
  {32'h426977fc, 32'h41455ba2} /* (21, 29, 23) {real, imag} */,
  {32'hc1e11319, 32'h408242f8} /* (21, 29, 22) {real, imag} */,
  {32'h41c54f95, 32'hc1ef5d21} /* (21, 29, 21) {real, imag} */,
  {32'hc17ac052, 32'hc1d76bfc} /* (21, 29, 20) {real, imag} */,
  {32'h4153d8ca, 32'h41037f39} /* (21, 29, 19) {real, imag} */,
  {32'h41991320, 32'hc15a5932} /* (21, 29, 18) {real, imag} */,
  {32'hc116b1eb, 32'h4126c17c} /* (21, 29, 17) {real, imag} */,
  {32'hc1c0b7ca, 32'h40bc4d74} /* (21, 29, 16) {real, imag} */,
  {32'h40a99eea, 32'hc153fce4} /* (21, 29, 15) {real, imag} */,
  {32'hc1575624, 32'hc136da06} /* (21, 29, 14) {real, imag} */,
  {32'hc156fe3e, 32'h407c5114} /* (21, 29, 13) {real, imag} */,
  {32'hc1684522, 32'hc24161fe} /* (21, 29, 12) {real, imag} */,
  {32'hc2193792, 32'h411ec22a} /* (21, 29, 11) {real, imag} */,
  {32'hc1f15ffb, 32'h4151bf00} /* (21, 29, 10) {real, imag} */,
  {32'h423731ec, 32'h41d3a409} /* (21, 29, 9) {real, imag} */,
  {32'hc0a539ca, 32'h4213462c} /* (21, 29, 8) {real, imag} */,
  {32'hc2177fbe, 32'h428bf6af} /* (21, 29, 7) {real, imag} */,
  {32'hc2362572, 32'hc24bb2fc} /* (21, 29, 6) {real, imag} */,
  {32'h41e9d9be, 32'h42d46574} /* (21, 29, 5) {real, imag} */,
  {32'h423e2f16, 32'h41fef287} /* (21, 29, 4) {real, imag} */,
  {32'h425d3192, 32'hc21e8724} /* (21, 29, 3) {real, imag} */,
  {32'hc1aecd40, 32'h42ec4e8c} /* (21, 29, 2) {real, imag} */,
  {32'h421670dc, 32'hc2d18c2c} /* (21, 29, 1) {real, imag} */,
  {32'h42ba135a, 32'hc2278902} /* (21, 29, 0) {real, imag} */,
  {32'h42f582cc, 32'hbfe1f2c8} /* (21, 28, 31) {real, imag} */,
  {32'hc2b50fb4, 32'h42ef4639} /* (21, 28, 30) {real, imag} */,
  {32'h42a8b297, 32'h41f479b8} /* (21, 28, 29) {real, imag} */,
  {32'h4191779c, 32'hc235043c} /* (21, 28, 28) {real, imag} */,
  {32'hc25f96ba, 32'hc1ec30ec} /* (21, 28, 27) {real, imag} */,
  {32'hc2986c66, 32'hc2484eef} /* (21, 28, 26) {real, imag} */,
  {32'h42a31da5, 32'h423af418} /* (21, 28, 25) {real, imag} */,
  {32'hc0b12c7c, 32'h4195c978} /* (21, 28, 24) {real, imag} */,
  {32'hc012e9bc, 32'h42621e07} /* (21, 28, 23) {real, imag} */,
  {32'h4012beb0, 32'h41f599f7} /* (21, 28, 22) {real, imag} */,
  {32'hc1f6ada2, 32'hc0bfea69} /* (21, 28, 21) {real, imag} */,
  {32'hc1ee18f2, 32'hc1c2f77a} /* (21, 28, 20) {real, imag} */,
  {32'hc1ea1551, 32'h4092dab2} /* (21, 28, 19) {real, imag} */,
  {32'hbfef0e50, 32'hc156cf6e} /* (21, 28, 18) {real, imag} */,
  {32'h418ae73a, 32'hc00262b4} /* (21, 28, 17) {real, imag} */,
  {32'hc036c8e0, 32'hc1934738} /* (21, 28, 16) {real, imag} */,
  {32'hbddfe200, 32'h41b27574} /* (21, 28, 15) {real, imag} */,
  {32'h3fc71a30, 32'h4188727b} /* (21, 28, 14) {real, imag} */,
  {32'h41865d81, 32'h4124f8d9} /* (21, 28, 13) {real, imag} */,
  {32'h418fe336, 32'hc1a89796} /* (21, 28, 12) {real, imag} */,
  {32'hbf69e2b0, 32'hc16d7c78} /* (21, 28, 11) {real, imag} */,
  {32'hc23900a9, 32'hc02fd0d8} /* (21, 28, 10) {real, imag} */,
  {32'hc1d03338, 32'h4173fe6c} /* (21, 28, 9) {real, imag} */,
  {32'h40ef22ec, 32'hc121b6a3} /* (21, 28, 8) {real, imag} */,
  {32'hc134f928, 32'hc2ae5f8e} /* (21, 28, 7) {real, imag} */,
  {32'h422f2550, 32'h41f67002} /* (21, 28, 6) {real, imag} */,
  {32'hc2cae5d3, 32'hc24729ce} /* (21, 28, 5) {real, imag} */,
  {32'h414260b3, 32'h4232b71a} /* (21, 28, 4) {real, imag} */,
  {32'hc0c8a510, 32'hc231dba8} /* (21, 28, 3) {real, imag} */,
  {32'h40040bc0, 32'h42988b0b} /* (21, 28, 2) {real, imag} */,
  {32'h41432874, 32'hc1b5a6c0} /* (21, 28, 1) {real, imag} */,
  {32'h4218446d, 32'h417c5c5b} /* (21, 28, 0) {real, imag} */,
  {32'hc31f86ac, 32'h425b224e} /* (21, 27, 31) {real, imag} */,
  {32'h425776ec, 32'h41c023bc} /* (21, 27, 30) {real, imag} */,
  {32'hc03f0482, 32'h425565ba} /* (21, 27, 29) {real, imag} */,
  {32'hc147e23a, 32'h427ac2eb} /* (21, 27, 28) {real, imag} */,
  {32'h418b2413, 32'hc27cee78} /* (21, 27, 27) {real, imag} */,
  {32'hc190b870, 32'h41807ca4} /* (21, 27, 26) {real, imag} */,
  {32'hc22786e4, 32'h420ff730} /* (21, 27, 25) {real, imag} */,
  {32'h4236d746, 32'hc1818c00} /* (21, 27, 24) {real, imag} */,
  {32'h41a090fe, 32'h422c9ffc} /* (21, 27, 23) {real, imag} */,
  {32'hc0901cb4, 32'hc1c3e162} /* (21, 27, 22) {real, imag} */,
  {32'h41ae3677, 32'hc2034152} /* (21, 27, 21) {real, imag} */,
  {32'hc2096f3c, 32'h40408c14} /* (21, 27, 20) {real, imag} */,
  {32'hc1ad1de9, 32'hc13533c4} /* (21, 27, 19) {real, imag} */,
  {32'hc1639f9e, 32'hc04e1174} /* (21, 27, 18) {real, imag} */,
  {32'h41a08d79, 32'h40e05b2c} /* (21, 27, 17) {real, imag} */,
  {32'h41852eaf, 32'h3f44f470} /* (21, 27, 16) {real, imag} */,
  {32'hbfc9df90, 32'hc0334648} /* (21, 27, 15) {real, imag} */,
  {32'hc10d12e2, 32'h40dc80b6} /* (21, 27, 14) {real, imag} */,
  {32'hc0cc3ff5, 32'hc1e87142} /* (21, 27, 13) {real, imag} */,
  {32'h41254564, 32'hc1376e85} /* (21, 27, 12) {real, imag} */,
  {32'h4168662a, 32'h41adbae8} /* (21, 27, 11) {real, imag} */,
  {32'hc2043bfe, 32'hc0b00560} /* (21, 27, 10) {real, imag} */,
  {32'h3f8bb1a8, 32'h41d2a379} /* (21, 27, 9) {real, imag} */,
  {32'h40f68bec, 32'hc0de6c38} /* (21, 27, 8) {real, imag} */,
  {32'hc1bae1f4, 32'hc21f0f18} /* (21, 27, 7) {real, imag} */,
  {32'hc1430dab, 32'hc1333dd4} /* (21, 27, 6) {real, imag} */,
  {32'h421dc434, 32'h41c85b74} /* (21, 27, 5) {real, imag} */,
  {32'h41baaa71, 32'h428305c6} /* (21, 27, 4) {real, imag} */,
  {32'h40e54b19, 32'hbf818d40} /* (21, 27, 3) {real, imag} */,
  {32'h42247aaa, 32'hc25b099c} /* (21, 27, 2) {real, imag} */,
  {32'hc275a018, 32'hc2aaa6d1} /* (21, 27, 1) {real, imag} */,
  {32'hc264a594, 32'hc1b3e218} /* (21, 27, 0) {real, imag} */,
  {32'h423bdffe, 32'hc198627c} /* (21, 26, 31) {real, imag} */,
  {32'hc0de3ab1, 32'hc21ede22} /* (21, 26, 30) {real, imag} */,
  {32'h42159dfb, 32'hc108d300} /* (21, 26, 29) {real, imag} */,
  {32'h42515386, 32'h42236d02} /* (21, 26, 28) {real, imag} */,
  {32'h420ce183, 32'h41860b6e} /* (21, 26, 27) {real, imag} */,
  {32'hc20b940b, 32'hc23586f2} /* (21, 26, 26) {real, imag} */,
  {32'hc201cb5a, 32'h4188cfb0} /* (21, 26, 25) {real, imag} */,
  {32'hc217cde2, 32'h409b5ab0} /* (21, 26, 24) {real, imag} */,
  {32'h421d3227, 32'hc1e1b873} /* (21, 26, 23) {real, imag} */,
  {32'hbfe84b10, 32'hc26821f2} /* (21, 26, 22) {real, imag} */,
  {32'h40f93b92, 32'hc1cf3e61} /* (21, 26, 21) {real, imag} */,
  {32'hbf586ac0, 32'hc1aa7f3f} /* (21, 26, 20) {real, imag} */,
  {32'hc0ef6664, 32'hc0832d4a} /* (21, 26, 19) {real, imag} */,
  {32'hc0afad8e, 32'hc0ee33ac} /* (21, 26, 18) {real, imag} */,
  {32'h40875fdc, 32'h40de9bde} /* (21, 26, 17) {real, imag} */,
  {32'h414cc1c0, 32'hc1631c5b} /* (21, 26, 16) {real, imag} */,
  {32'h41111bc2, 32'h416b9b59} /* (21, 26, 15) {real, imag} */,
  {32'h41743b85, 32'hc14c541a} /* (21, 26, 14) {real, imag} */,
  {32'hc17016ce, 32'h4180c6c6} /* (21, 26, 13) {real, imag} */,
  {32'h418b7374, 32'hc1e94fad} /* (21, 26, 12) {real, imag} */,
  {32'hc1068937, 32'hc1715a56} /* (21, 26, 11) {real, imag} */,
  {32'h402537a8, 32'h41fe6acb} /* (21, 26, 10) {real, imag} */,
  {32'h4136a360, 32'h40beb5c4} /* (21, 26, 9) {real, imag} */,
  {32'hc25ac73c, 32'hc218c834} /* (21, 26, 8) {real, imag} */,
  {32'hc0f35ee8, 32'h41a33882} /* (21, 26, 7) {real, imag} */,
  {32'hc213d7e7, 32'h419b360c} /* (21, 26, 6) {real, imag} */,
  {32'hc240c1b7, 32'hc1a57ab8} /* (21, 26, 5) {real, imag} */,
  {32'h420f113a, 32'h418bdce9} /* (21, 26, 4) {real, imag} */,
  {32'hc26b2781, 32'h42476f6c} /* (21, 26, 3) {real, imag} */,
  {32'hc0b11703, 32'hc1ff6ce5} /* (21, 26, 2) {real, imag} */,
  {32'h4304ab5e, 32'hc232539e} /* (21, 26, 1) {real, imag} */,
  {32'hc2af1353, 32'h4179ab3d} /* (21, 26, 0) {real, imag} */,
  {32'h42b82c73, 32'h41bc394c} /* (21, 25, 31) {real, imag} */,
  {32'hbf11ad60, 32'hc0bfe878} /* (21, 25, 30) {real, imag} */,
  {32'hc1cef6be, 32'h4297b1fe} /* (21, 25, 29) {real, imag} */,
  {32'h420cbf1c, 32'hc196921d} /* (21, 25, 28) {real, imag} */,
  {32'hc2152033, 32'h42a3ee94} /* (21, 25, 27) {real, imag} */,
  {32'h428d23f2, 32'h3ffcae28} /* (21, 25, 26) {real, imag} */,
  {32'h41aa09e0, 32'hc2366414} /* (21, 25, 25) {real, imag} */,
  {32'h4219ccc0, 32'hc128c78d} /* (21, 25, 24) {real, imag} */,
  {32'h413702c0, 32'h3b428000} /* (21, 25, 23) {real, imag} */,
  {32'hc0db4f9c, 32'h41422949} /* (21, 25, 22) {real, imag} */,
  {32'h41d96dad, 32'hc19ff09b} /* (21, 25, 21) {real, imag} */,
  {32'hbffd58b0, 32'h3f1109d0} /* (21, 25, 20) {real, imag} */,
  {32'hc16f1ffc, 32'h419f928f} /* (21, 25, 19) {real, imag} */,
  {32'h40aac27c, 32'h4120d204} /* (21, 25, 18) {real, imag} */,
  {32'hc11aae47, 32'hc162aec2} /* (21, 25, 17) {real, imag} */,
  {32'hc16ab8ea, 32'h3fb349a8} /* (21, 25, 16) {real, imag} */,
  {32'h4089d22e, 32'hc05c8c70} /* (21, 25, 15) {real, imag} */,
  {32'hc026d988, 32'h40df8708} /* (21, 25, 14) {real, imag} */,
  {32'hc0fcce48, 32'hc1cee1a9} /* (21, 25, 13) {real, imag} */,
  {32'h421af264, 32'hc15a7460} /* (21, 25, 12) {real, imag} */,
  {32'hc1cbe38b, 32'h400590d8} /* (21, 25, 11) {real, imag} */,
  {32'h4026f268, 32'hc229cd6b} /* (21, 25, 10) {real, imag} */,
  {32'hc20d35f2, 32'h416b32ec} /* (21, 25, 9) {real, imag} */,
  {32'h41f58f4d, 32'h40b3c5de} /* (21, 25, 8) {real, imag} */,
  {32'hc0d793f2, 32'h41686abe} /* (21, 25, 7) {real, imag} */,
  {32'hc1bd4545, 32'h41a1f724} /* (21, 25, 6) {real, imag} */,
  {32'hc2693ebd, 32'hc15a3f74} /* (21, 25, 5) {real, imag} */,
  {32'h3f858b90, 32'h41be81e5} /* (21, 25, 4) {real, imag} */,
  {32'h425acc6d, 32'hc29b9474} /* (21, 25, 3) {real, imag} */,
  {32'hc23086ba, 32'h4085a918} /* (21, 25, 2) {real, imag} */,
  {32'h42a40da7, 32'h41aa4c24} /* (21, 25, 1) {real, imag} */,
  {32'hc28dc3a4, 32'hc1e56038} /* (21, 25, 0) {real, imag} */,
  {32'h3fb5bdb4, 32'h41a8b976} /* (21, 24, 31) {real, imag} */,
  {32'hc1ddfc02, 32'hbe8323e0} /* (21, 24, 30) {real, imag} */,
  {32'h41abb176, 32'hbf417310} /* (21, 24, 29) {real, imag} */,
  {32'hc2188158, 32'hc2018e71} /* (21, 24, 28) {real, imag} */,
  {32'hc1af5c64, 32'hc217a92d} /* (21, 24, 27) {real, imag} */,
  {32'hc256e56c, 32'hc1d481d4} /* (21, 24, 26) {real, imag} */,
  {32'h4228c906, 32'hc01ca0f4} /* (21, 24, 25) {real, imag} */,
  {32'h4221fe79, 32'h4043c548} /* (21, 24, 24) {real, imag} */,
  {32'hc187f1f8, 32'h40ef1886} /* (21, 24, 23) {real, imag} */,
  {32'hc19739e6, 32'h4162f253} /* (21, 24, 22) {real, imag} */,
  {32'hc05e6608, 32'h41831428} /* (21, 24, 21) {real, imag} */,
  {32'hc047c34b, 32'hc12f483f} /* (21, 24, 20) {real, imag} */,
  {32'h4122bb5a, 32'hc201e31a} /* (21, 24, 19) {real, imag} */,
  {32'hc0dd4c60, 32'hc0662dc5} /* (21, 24, 18) {real, imag} */,
  {32'hc0f8c7f2, 32'hc07fd7a0} /* (21, 24, 17) {real, imag} */,
  {32'h40b2782d, 32'h3e6f9600} /* (21, 24, 16) {real, imag} */,
  {32'hc0f896a8, 32'h40e7941c} /* (21, 24, 15) {real, imag} */,
  {32'h4155d046, 32'h4134d61c} /* (21, 24, 14) {real, imag} */,
  {32'hbf529f18, 32'hc05a31c8} /* (21, 24, 13) {real, imag} */,
  {32'hbff5bad6, 32'h41368e69} /* (21, 24, 12) {real, imag} */,
  {32'h42174cb0, 32'hbf8b287c} /* (21, 24, 11) {real, imag} */,
  {32'h421e2de9, 32'hc19fb6ca} /* (21, 24, 10) {real, imag} */,
  {32'hc0a41e9e, 32'hc1bbdbc0} /* (21, 24, 9) {real, imag} */,
  {32'hc1a1e6b2, 32'h41b81ecf} /* (21, 24, 8) {real, imag} */,
  {32'hc27fa21e, 32'h41a8d3bc} /* (21, 24, 7) {real, imag} */,
  {32'h41071a98, 32'h40f6709e} /* (21, 24, 6) {real, imag} */,
  {32'h402d7894, 32'h4202be21} /* (21, 24, 5) {real, imag} */,
  {32'h42046e3e, 32'h4211a32f} /* (21, 24, 4) {real, imag} */,
  {32'hc1a4fa56, 32'hc17e8fb5} /* (21, 24, 3) {real, imag} */,
  {32'hc1ea198a, 32'hc185e530} /* (21, 24, 2) {real, imag} */,
  {32'hc1006968, 32'h41f117ee} /* (21, 24, 1) {real, imag} */,
  {32'h418217e1, 32'hc1979cdc} /* (21, 24, 0) {real, imag} */,
  {32'h42af45ac, 32'hc0d7b8b5} /* (21, 23, 31) {real, imag} */,
  {32'hbfc74650, 32'h4221ac62} /* (21, 23, 30) {real, imag} */,
  {32'h409c14ae, 32'h422e87a6} /* (21, 23, 29) {real, imag} */,
  {32'hbf8a6940, 32'hc1aed19c} /* (21, 23, 28) {real, imag} */,
  {32'h41d87a97, 32'h415d5d49} /* (21, 23, 27) {real, imag} */,
  {32'h41052bb9, 32'hc1ea3038} /* (21, 23, 26) {real, imag} */,
  {32'hc01dc0f0, 32'hc103c63c} /* (21, 23, 25) {real, imag} */,
  {32'h41d2f45f, 32'hc0b19656} /* (21, 23, 24) {real, imag} */,
  {32'hc1a132d8, 32'h401b0978} /* (21, 23, 23) {real, imag} */,
  {32'hc181cb4b, 32'h3f8b9448} /* (21, 23, 22) {real, imag} */,
  {32'hc18ec6f6, 32'hc096d102} /* (21, 23, 21) {real, imag} */,
  {32'h4114a55e, 32'hc17df5fe} /* (21, 23, 20) {real, imag} */,
  {32'h40874724, 32'hc13df535} /* (21, 23, 19) {real, imag} */,
  {32'hc118af88, 32'hc05e0d89} /* (21, 23, 18) {real, imag} */,
  {32'hc0f37ff2, 32'h4003b3b4} /* (21, 23, 17) {real, imag} */,
  {32'h409b815c, 32'h41122f52} /* (21, 23, 16) {real, imag} */,
  {32'hc0b03b6a, 32'h41accc32} /* (21, 23, 15) {real, imag} */,
  {32'hc08a5c45, 32'hbfabfd52} /* (21, 23, 14) {real, imag} */,
  {32'h40be6e30, 32'hc0d35b42} /* (21, 23, 13) {real, imag} */,
  {32'hc09bb684, 32'h40dfd809} /* (21, 23, 12) {real, imag} */,
  {32'h411172ff, 32'h4105e283} /* (21, 23, 11) {real, imag} */,
  {32'hc1ff6f39, 32'h41c72342} /* (21, 23, 10) {real, imag} */,
  {32'hc1befc44, 32'hc1864761} /* (21, 23, 9) {real, imag} */,
  {32'hc1fa1077, 32'hc1d373da} /* (21, 23, 8) {real, imag} */,
  {32'h41c246c5, 32'hc2037e88} /* (21, 23, 7) {real, imag} */,
  {32'hbfa9d7f8, 32'h40e895da} /* (21, 23, 6) {real, imag} */,
  {32'hc1cdff6b, 32'hc1ed9620} /* (21, 23, 5) {real, imag} */,
  {32'hc24c0964, 32'hc0fd98a6} /* (21, 23, 4) {real, imag} */,
  {32'hc2079940, 32'hc068c1e0} /* (21, 23, 3) {real, imag} */,
  {32'h42140f38, 32'hc20ce794} /* (21, 23, 2) {real, imag} */,
  {32'hc2186deb, 32'h41032d98} /* (21, 23, 1) {real, imag} */,
  {32'h4245c822, 32'h4258ca22} /* (21, 23, 0) {real, imag} */,
  {32'hc26343a7, 32'hc211863f} /* (21, 22, 31) {real, imag} */,
  {32'hc1dc5184, 32'h4136f4b1} /* (21, 22, 30) {real, imag} */,
  {32'hc145f5e8, 32'hc1fd2417} /* (21, 22, 29) {real, imag} */,
  {32'hc1878d5c, 32'hc1961620} /* (21, 22, 28) {real, imag} */,
  {32'hc1674d95, 32'h419242f2} /* (21, 22, 27) {real, imag} */,
  {32'h4121e4ee, 32'h4120e135} /* (21, 22, 26) {real, imag} */,
  {32'h40f94dbd, 32'h3f87a480} /* (21, 22, 25) {real, imag} */,
  {32'h416151bc, 32'h41d7f7be} /* (21, 22, 24) {real, imag} */,
  {32'hc1b49ab5, 32'h4220f379} /* (21, 22, 23) {real, imag} */,
  {32'h4139e55a, 32'hc1af9005} /* (21, 22, 22) {real, imag} */,
  {32'h4088c586, 32'h4000a277} /* (21, 22, 21) {real, imag} */,
  {32'h418f3e36, 32'hc0665739} /* (21, 22, 20) {real, imag} */,
  {32'hc17ef62e, 32'h40e0cfb6} /* (21, 22, 19) {real, imag} */,
  {32'h417482a3, 32'hc0bf1ca4} /* (21, 22, 18) {real, imag} */,
  {32'hbf193ec0, 32'hc002aefe} /* (21, 22, 17) {real, imag} */,
  {32'hbf3c4c78, 32'h40bdb918} /* (21, 22, 16) {real, imag} */,
  {32'h40c51850, 32'h3f6358b8} /* (21, 22, 15) {real, imag} */,
  {32'hc117e1c5, 32'hc11b8bae} /* (21, 22, 14) {real, imag} */,
  {32'h405d9266, 32'h409311da} /* (21, 22, 13) {real, imag} */,
  {32'hc1611595, 32'hc0b28a90} /* (21, 22, 12) {real, imag} */,
  {32'h40eb417a, 32'hc0575a67} /* (21, 22, 11) {real, imag} */,
  {32'hc13b4282, 32'h3eb72c80} /* (21, 22, 10) {real, imag} */,
  {32'hc21c60c6, 32'hc1a540f6} /* (21, 22, 9) {real, imag} */,
  {32'h4261726b, 32'h4239743b} /* (21, 22, 8) {real, imag} */,
  {32'hbfdec9b4, 32'hc2537fda} /* (21, 22, 7) {real, imag} */,
  {32'hc1162522, 32'h41e8c106} /* (21, 22, 6) {real, imag} */,
  {32'h41e3a6be, 32'h414a8cd0} /* (21, 22, 5) {real, imag} */,
  {32'h40d2f94e, 32'hc1f01014} /* (21, 22, 4) {real, imag} */,
  {32'h4206a8ec, 32'h41adadb9} /* (21, 22, 3) {real, imag} */,
  {32'hc14c4e18, 32'h410effc3} /* (21, 22, 2) {real, imag} */,
  {32'hc0e140c0, 32'hc00fb470} /* (21, 22, 1) {real, imag} */,
  {32'hc15440fe, 32'hc2886924} /* (21, 22, 0) {real, imag} */,
  {32'hbf9183b0, 32'h41379aa9} /* (21, 21, 31) {real, imag} */,
  {32'hc15926f6, 32'hbfc2df80} /* (21, 21, 30) {real, imag} */,
  {32'hc2200a65, 32'hc0d41a0b} /* (21, 21, 29) {real, imag} */,
  {32'hc236f08a, 32'hc23baf8d} /* (21, 21, 28) {real, imag} */,
  {32'hc0929900, 32'h40adf753} /* (21, 21, 27) {real, imag} */,
  {32'hc0d73f7a, 32'h419bb105} /* (21, 21, 26) {real, imag} */,
  {32'hbf686fa0, 32'h40545900} /* (21, 21, 25) {real, imag} */,
  {32'h40760da8, 32'hc1039cc8} /* (21, 21, 24) {real, imag} */,
  {32'hc144e6c5, 32'h40f28020} /* (21, 21, 23) {real, imag} */,
  {32'h40658cac, 32'h411e19ed} /* (21, 21, 22) {real, imag} */,
  {32'hbf1f04bc, 32'hc19e40c1} /* (21, 21, 21) {real, imag} */,
  {32'h411387b0, 32'hc0844574} /* (21, 21, 20) {real, imag} */,
  {32'hc074d7b8, 32'h404cbfb6} /* (21, 21, 19) {real, imag} */,
  {32'hc0635714, 32'h410fc016} /* (21, 21, 18) {real, imag} */,
  {32'h3faaaee8, 32'hc0848314} /* (21, 21, 17) {real, imag} */,
  {32'hc0482860, 32'h4071dd88} /* (21, 21, 16) {real, imag} */,
  {32'hbffcb548, 32'hc11e088a} /* (21, 21, 15) {real, imag} */,
  {32'hc15851dd, 32'h411fd398} /* (21, 21, 14) {real, imag} */,
  {32'hc0c2e03c, 32'h40964b63} /* (21, 21, 13) {real, imag} */,
  {32'hc0ca156c, 32'h41a1f990} /* (21, 21, 12) {real, imag} */,
  {32'h409389d6, 32'h40efe075} /* (21, 21, 11) {real, imag} */,
  {32'h414e2a5f, 32'h4101b3f7} /* (21, 21, 10) {real, imag} */,
  {32'hc09fb686, 32'h3fa88f48} /* (21, 21, 9) {real, imag} */,
  {32'h418bc169, 32'h417a9df0} /* (21, 21, 8) {real, imag} */,
  {32'hc1b173f7, 32'h413b9ad5} /* (21, 21, 7) {real, imag} */,
  {32'h416f1dc9, 32'h41cc3af3} /* (21, 21, 6) {real, imag} */,
  {32'hc10512db, 32'h4199862b} /* (21, 21, 5) {real, imag} */,
  {32'hc0afa5e0, 32'h40bcfe08} /* (21, 21, 4) {real, imag} */,
  {32'hc1e384b6, 32'hc112c29c} /* (21, 21, 3) {real, imag} */,
  {32'hc1cb08c5, 32'hc258e962} /* (21, 21, 2) {real, imag} */,
  {32'hc26e1b02, 32'hc15d07af} /* (21, 21, 1) {real, imag} */,
  {32'hc1801f6c, 32'h42030c34} /* (21, 21, 0) {real, imag} */,
  {32'hc1e352b8, 32'h41c79682} /* (21, 20, 31) {real, imag} */,
  {32'hc1cf5b7e, 32'hc1eb9ed2} /* (21, 20, 30) {real, imag} */,
  {32'hc1711350, 32'hc0ed6226} /* (21, 20, 29) {real, imag} */,
  {32'h40b6227a, 32'hc01de9f0} /* (21, 20, 28) {real, imag} */,
  {32'hc12c3b6c, 32'h41a9df1e} /* (21, 20, 27) {real, imag} */,
  {32'h40bdd0b3, 32'h40070c40} /* (21, 20, 26) {real, imag} */,
  {32'h41b82fea, 32'h40705898} /* (21, 20, 25) {real, imag} */,
  {32'hc1465158, 32'h412f6e2c} /* (21, 20, 24) {real, imag} */,
  {32'h40547982, 32'hc08506f4} /* (21, 20, 23) {real, imag} */,
  {32'h4094553f, 32'hbeaf81d0} /* (21, 20, 22) {real, imag} */,
  {32'hc09b8ade, 32'h407a1b20} /* (21, 20, 21) {real, imag} */,
  {32'hbe16cea0, 32'h40655152} /* (21, 20, 20) {real, imag} */,
  {32'h406f9a17, 32'h414d5d62} /* (21, 20, 19) {real, imag} */,
  {32'h3ef6b490, 32'hc095b15b} /* (21, 20, 18) {real, imag} */,
  {32'hc031940a, 32'h40f36d5c} /* (21, 20, 17) {real, imag} */,
  {32'hbfc90b2c, 32'h3eb47e80} /* (21, 20, 16) {real, imag} */,
  {32'hc07b767a, 32'h41081dfe} /* (21, 20, 15) {real, imag} */,
  {32'h41143300, 32'h414c125e} /* (21, 20, 14) {real, imag} */,
  {32'hc1012023, 32'hc11d92aa} /* (21, 20, 13) {real, imag} */,
  {32'hbfec99d4, 32'h416e7af4} /* (21, 20, 12) {real, imag} */,
  {32'h3fe52628, 32'h41738bee} /* (21, 20, 11) {real, imag} */,
  {32'hc13652ac, 32'h41703060} /* (21, 20, 10) {real, imag} */,
  {32'hc0c9fe91, 32'h40ca5012} /* (21, 20, 9) {real, imag} */,
  {32'h405dbc4e, 32'hc1afd2a6} /* (21, 20, 8) {real, imag} */,
  {32'hc1734bcc, 32'hc15b8c38} /* (21, 20, 7) {real, imag} */,
  {32'hc193b0b7, 32'hc1f01924} /* (21, 20, 6) {real, imag} */,
  {32'h415deb08, 32'h416587f5} /* (21, 20, 5) {real, imag} */,
  {32'h4196240a, 32'hc0827be2} /* (21, 20, 4) {real, imag} */,
  {32'hbeccf630, 32'hbff00f98} /* (21, 20, 3) {real, imag} */,
  {32'hc2060716, 32'h402dbaa0} /* (21, 20, 2) {real, imag} */,
  {32'h4199a112, 32'hc1d3436e} /* (21, 20, 1) {real, imag} */,
  {32'h403ad12a, 32'h419dfbea} /* (21, 20, 0) {real, imag} */,
  {32'hc137c814, 32'hc081df8a} /* (21, 19, 31) {real, imag} */,
  {32'hc112da72, 32'hc181f162} /* (21, 19, 30) {real, imag} */,
  {32'hc1a8a4c5, 32'h3fe9e488} /* (21, 19, 29) {real, imag} */,
  {32'h41299059, 32'hc1233ece} /* (21, 19, 28) {real, imag} */,
  {32'h405a364a, 32'h41ada590} /* (21, 19, 27) {real, imag} */,
  {32'h417dd471, 32'hbe9d5600} /* (21, 19, 26) {real, imag} */,
  {32'hbfb49970, 32'hc08de706} /* (21, 19, 25) {real, imag} */,
  {32'h41167e56, 32'h40a04b60} /* (21, 19, 24) {real, imag} */,
  {32'hc08cd97b, 32'h411da0a0} /* (21, 19, 23) {real, imag} */,
  {32'h4024010b, 32'hc07d64ba} /* (21, 19, 22) {real, imag} */,
  {32'h40a84d23, 32'h4123d8f8} /* (21, 19, 21) {real, imag} */,
  {32'h40a46724, 32'h409b0c20} /* (21, 19, 20) {real, imag} */,
  {32'hbf931034, 32'h40976798} /* (21, 19, 19) {real, imag} */,
  {32'h3ff44023, 32'h3ffa771c} /* (21, 19, 18) {real, imag} */,
  {32'hc012bbf0, 32'h404e8cea} /* (21, 19, 17) {real, imag} */,
  {32'hc01080bc, 32'h3ffd381c} /* (21, 19, 16) {real, imag} */,
  {32'hc09d3cd6, 32'hbfa671c4} /* (21, 19, 15) {real, imag} */,
  {32'h3dd33eb0, 32'hc11883fa} /* (21, 19, 14) {real, imag} */,
  {32'hbfe37404, 32'h409490f4} /* (21, 19, 13) {real, imag} */,
  {32'h405abd53, 32'hc0f383b8} /* (21, 19, 12) {real, imag} */,
  {32'hbf07e278, 32'h3fd79df4} /* (21, 19, 11) {real, imag} */,
  {32'h4119a15b, 32'h416f5bf6} /* (21, 19, 10) {real, imag} */,
  {32'h4173abee, 32'hc135fa88} /* (21, 19, 9) {real, imag} */,
  {32'h4087ed93, 32'hbf9a9472} /* (21, 19, 8) {real, imag} */,
  {32'h4198d9d1, 32'h40f4b6f8} /* (21, 19, 7) {real, imag} */,
  {32'h4125c261, 32'hc085b40e} /* (21, 19, 6) {real, imag} */,
  {32'hc12a86c6, 32'hc163f670} /* (21, 19, 5) {real, imag} */,
  {32'hc0ae8966, 32'h3ee9c6c0} /* (21, 19, 4) {real, imag} */,
  {32'h40dd832f, 32'hc18d89dc} /* (21, 19, 3) {real, imag} */,
  {32'h4100580e, 32'hc1c3c4f2} /* (21, 19, 2) {real, imag} */,
  {32'h411793d8, 32'h418afc30} /* (21, 19, 1) {real, imag} */,
  {32'h41a97eaa, 32'hc14cad16} /* (21, 19, 0) {real, imag} */,
  {32'hc1925b52, 32'hc1cd5faf} /* (21, 18, 31) {real, imag} */,
  {32'h413416b8, 32'hc087aeda} /* (21, 18, 30) {real, imag} */,
  {32'h3fb1e486, 32'h417c81dd} /* (21, 18, 29) {real, imag} */,
  {32'h3f897b2c, 32'h403c6dd6} /* (21, 18, 28) {real, imag} */,
  {32'h3fcb1a33, 32'hc1999508} /* (21, 18, 27) {real, imag} */,
  {32'hbe82fdc0, 32'h40d2c890} /* (21, 18, 26) {real, imag} */,
  {32'hc1302766, 32'h3fd68fb6} /* (21, 18, 25) {real, imag} */,
  {32'h3f5f6558, 32'h40a199ac} /* (21, 18, 24) {real, imag} */,
  {32'hc098407b, 32'h4018e8ac} /* (21, 18, 23) {real, imag} */,
  {32'hc0c7885d, 32'hbfba4152} /* (21, 18, 22) {real, imag} */,
  {32'hbf3f6238, 32'hc0ff275c} /* (21, 18, 21) {real, imag} */,
  {32'h3f1a0600, 32'h4062efff} /* (21, 18, 20) {real, imag} */,
  {32'h40cc4440, 32'hc046ae80} /* (21, 18, 19) {real, imag} */,
  {32'h400128be, 32'h4009a94f} /* (21, 18, 18) {real, imag} */,
  {32'hc01d8454, 32'hc03f09f4} /* (21, 18, 17) {real, imag} */,
  {32'h40ae5c06, 32'h40ec268f} /* (21, 18, 16) {real, imag} */,
  {32'h3f9e7908, 32'hc00565ec} /* (21, 18, 15) {real, imag} */,
  {32'h410695bc, 32'hc08d2934} /* (21, 18, 14) {real, imag} */,
  {32'h405f3f39, 32'h409c6474} /* (21, 18, 13) {real, imag} */,
  {32'hbf4bae6c, 32'h3e9d2928} /* (21, 18, 12) {real, imag} */,
  {32'hbf1ee46c, 32'hbf40bf80} /* (21, 18, 11) {real, imag} */,
  {32'hc1a09585, 32'hbefe9348} /* (21, 18, 10) {real, imag} */,
  {32'h41219a8e, 32'hc0c7afca} /* (21, 18, 9) {real, imag} */,
  {32'hc1206836, 32'h41734532} /* (21, 18, 8) {real, imag} */,
  {32'hbecced50, 32'hbf4859cc} /* (21, 18, 7) {real, imag} */,
  {32'hc0d3aca6, 32'hbf9bc8aa} /* (21, 18, 6) {real, imag} */,
  {32'h407e1336, 32'h3ea481a0} /* (21, 18, 5) {real, imag} */,
  {32'hc0fe1ef7, 32'hc10e5f8e} /* (21, 18, 4) {real, imag} */,
  {32'h411205a3, 32'h418ea8be} /* (21, 18, 3) {real, imag} */,
  {32'hc1558cac, 32'hc161794d} /* (21, 18, 2) {real, imag} */,
  {32'hc012086c, 32'h419e9a11} /* (21, 18, 1) {real, imag} */,
  {32'hc09ef432, 32'h41969bf8} /* (21, 18, 0) {real, imag} */,
  {32'h411bf155, 32'hc0f32162} /* (21, 17, 31) {real, imag} */,
  {32'h3fe00b10, 32'h3e83f764} /* (21, 17, 30) {real, imag} */,
  {32'hbea8d7a0, 32'hc190092a} /* (21, 17, 29) {real, imag} */,
  {32'h401b3046, 32'h417ac85c} /* (21, 17, 28) {real, imag} */,
  {32'h414dd694, 32'hc128419e} /* (21, 17, 27) {real, imag} */,
  {32'hc0ca5a66, 32'hc11e1301} /* (21, 17, 26) {real, imag} */,
  {32'h40e03618, 32'h40b9e03f} /* (21, 17, 25) {real, imag} */,
  {32'hbf4f1e80, 32'hc12f0555} /* (21, 17, 24) {real, imag} */,
  {32'hc0aca517, 32'hbf28b254} /* (21, 17, 23) {real, imag} */,
  {32'h408bfcee, 32'h4091c0d0} /* (21, 17, 22) {real, imag} */,
  {32'h412971cc, 32'h4128a20f} /* (21, 17, 21) {real, imag} */,
  {32'h4006b81b, 32'h3f9c7be0} /* (21, 17, 20) {real, imag} */,
  {32'hc0e830ba, 32'h3fd22b74} /* (21, 17, 19) {real, imag} */,
  {32'h3f7d8b60, 32'hc0182108} /* (21, 17, 18) {real, imag} */,
  {32'hc00d114a, 32'h3f757828} /* (21, 17, 17) {real, imag} */,
  {32'hc06867ae, 32'hbfaa93a4} /* (21, 17, 16) {real, imag} */,
  {32'h3e81f770, 32'h3f951334} /* (21, 17, 15) {real, imag} */,
  {32'h3fa8fd50, 32'h4098afbb} /* (21, 17, 14) {real, imag} */,
  {32'h3fd436a0, 32'h40d44423} /* (21, 17, 13) {real, imag} */,
  {32'hc09578a2, 32'h40418f44} /* (21, 17, 12) {real, imag} */,
  {32'h40c72339, 32'hc0f9ddd2} /* (21, 17, 11) {real, imag} */,
  {32'h3f911922, 32'hc034a438} /* (21, 17, 10) {real, imag} */,
  {32'hc0e59cf9, 32'h401f7d77} /* (21, 17, 9) {real, imag} */,
  {32'hc19004b6, 32'hc15775bd} /* (21, 17, 8) {real, imag} */,
  {32'h4036fa50, 32'h4098e85d} /* (21, 17, 7) {real, imag} */,
  {32'h3f85a1b2, 32'h4088e732} /* (21, 17, 6) {real, imag} */,
  {32'hc021c112, 32'hc18e0fa4} /* (21, 17, 5) {real, imag} */,
  {32'hc05b131a, 32'h3f8c5964} /* (21, 17, 4) {real, imag} */,
  {32'hc14f3f4e, 32'hc13ffa2c} /* (21, 17, 3) {real, imag} */,
  {32'hc15f2752, 32'hc0172b16} /* (21, 17, 2) {real, imag} */,
  {32'h4194e408, 32'h411ec813} /* (21, 17, 1) {real, imag} */,
  {32'h41021168, 32'h3fbae174} /* (21, 17, 0) {real, imag} */,
  {32'hc0f6c0c8, 32'h40e47a25} /* (21, 16, 31) {real, imag} */,
  {32'h40a5a11d, 32'hc116f355} /* (21, 16, 30) {real, imag} */,
  {32'h41501995, 32'h3f811aac} /* (21, 16, 29) {real, imag} */,
  {32'h410c168c, 32'h3f82c916} /* (21, 16, 28) {real, imag} */,
  {32'hc15f1a57, 32'hc0b3b07e} /* (21, 16, 27) {real, imag} */,
  {32'h3fa9a860, 32'hc14d660f} /* (21, 16, 26) {real, imag} */,
  {32'h41113664, 32'h41831e6b} /* (21, 16, 25) {real, imag} */,
  {32'h40da1e12, 32'h413d4982} /* (21, 16, 24) {real, imag} */,
  {32'hbe82c040, 32'h417d325e} /* (21, 16, 23) {real, imag} */,
  {32'hc0596a01, 32'h40918e00} /* (21, 16, 22) {real, imag} */,
  {32'h4048eeb8, 32'h40c5107e} /* (21, 16, 21) {real, imag} */,
  {32'h4008f120, 32'hc0877be8} /* (21, 16, 20) {real, imag} */,
  {32'h4104780a, 32'h40414e58} /* (21, 16, 19) {real, imag} */,
  {32'h3d994850, 32'h3f81fe10} /* (21, 16, 18) {real, imag} */,
  {32'hc016980b, 32'h404702e4} /* (21, 16, 17) {real, imag} */,
  {32'h3f87f9d0, 32'hbe550860} /* (21, 16, 16) {real, imag} */,
  {32'h404390af, 32'h3ec55a04} /* (21, 16, 15) {real, imag} */,
  {32'h3fab025d, 32'hbfa03ffc} /* (21, 16, 14) {real, imag} */,
  {32'hc04706f7, 32'hc05b7d1c} /* (21, 16, 13) {real, imag} */,
  {32'hc08170e5, 32'h406cbd0d} /* (21, 16, 12) {real, imag} */,
  {32'hc0860c07, 32'hc0e50f32} /* (21, 16, 11) {real, imag} */,
  {32'hbfedd836, 32'hbffd8946} /* (21, 16, 10) {real, imag} */,
  {32'h41ba4087, 32'hc0262b28} /* (21, 16, 9) {real, imag} */,
  {32'h40ec2580, 32'h4066c148} /* (21, 16, 8) {real, imag} */,
  {32'hc0565d8e, 32'hbfde5e90} /* (21, 16, 7) {real, imag} */,
  {32'hc1156a8a, 32'h40cc855a} /* (21, 16, 6) {real, imag} */,
  {32'h3ecb6ee0, 32'hc1986702} /* (21, 16, 5) {real, imag} */,
  {32'hc106645e, 32'hbf90a2b4} /* (21, 16, 4) {real, imag} */,
  {32'hc108c33f, 32'h409f1879} /* (21, 16, 3) {real, imag} */,
  {32'hbee1d2b0, 32'hbf812298} /* (21, 16, 2) {real, imag} */,
  {32'hbf682f74, 32'hc10c0ce1} /* (21, 16, 1) {real, imag} */,
  {32'h41afffc1, 32'hc093100d} /* (21, 16, 0) {real, imag} */,
  {32'hc12b4951, 32'hbf740dd8} /* (21, 15, 31) {real, imag} */,
  {32'h42330ab0, 32'hc01f8278} /* (21, 15, 30) {real, imag} */,
  {32'h4101a71c, 32'h4149ecd6} /* (21, 15, 29) {real, imag} */,
  {32'h4009089b, 32'h41220a7e} /* (21, 15, 28) {real, imag} */,
  {32'h411d743b, 32'h41136edc} /* (21, 15, 27) {real, imag} */,
  {32'hc1665f34, 32'hc1516369} /* (21, 15, 26) {real, imag} */,
  {32'hc18d3db1, 32'h402cd390} /* (21, 15, 25) {real, imag} */,
  {32'hbed26b50, 32'hbfc7c3f0} /* (21, 15, 24) {real, imag} */,
  {32'hc11d0638, 32'h40f5c0b8} /* (21, 15, 23) {real, imag} */,
  {32'h400f1848, 32'h407b34f6} /* (21, 15, 22) {real, imag} */,
  {32'hc1031d84, 32'hc1149b54} /* (21, 15, 21) {real, imag} */,
  {32'h3f276afc, 32'hc08c62cf} /* (21, 15, 20) {real, imag} */,
  {32'hc0e7738f, 32'h40445273} /* (21, 15, 19) {real, imag} */,
  {32'h3ef056e0, 32'hc0508806} /* (21, 15, 18) {real, imag} */,
  {32'hc0921379, 32'hbfefada4} /* (21, 15, 17) {real, imag} */,
  {32'hc0636ad5, 32'hc07ada39} /* (21, 15, 16) {real, imag} */,
  {32'hc092fedf, 32'h3e789620} /* (21, 15, 15) {real, imag} */,
  {32'h4063bbf4, 32'hbe6f4148} /* (21, 15, 14) {real, imag} */,
  {32'h3e1a82e0, 32'h3f16d48c} /* (21, 15, 13) {real, imag} */,
  {32'hbfc2c04e, 32'h4044d05a} /* (21, 15, 12) {real, imag} */,
  {32'hc11d10da, 32'h415a7120} /* (21, 15, 11) {real, imag} */,
  {32'h4039cb8c, 32'h3d4f5780} /* (21, 15, 10) {real, imag} */,
  {32'hc0bde303, 32'h411b633c} /* (21, 15, 9) {real, imag} */,
  {32'hc135e466, 32'hc0002502} /* (21, 15, 8) {real, imag} */,
  {32'h40bae8c9, 32'hc1108f66} /* (21, 15, 7) {real, imag} */,
  {32'h4023a5be, 32'h4101381d} /* (21, 15, 6) {real, imag} */,
  {32'hc1242da1, 32'h40dbd6f7} /* (21, 15, 5) {real, imag} */,
  {32'hbfb5b466, 32'h413bb9c6} /* (21, 15, 4) {real, imag} */,
  {32'hc00114ec, 32'hc1d7ee0b} /* (21, 15, 3) {real, imag} */,
  {32'h413a262a, 32'hc0f7b9dc} /* (21, 15, 2) {real, imag} */,
  {32'h41343e73, 32'h40a059f3} /* (21, 15, 1) {real, imag} */,
  {32'hc0ec6194, 32'h413abec6} /* (21, 15, 0) {real, imag} */,
  {32'h40e848c3, 32'h40167220} /* (21, 14, 31) {real, imag} */,
  {32'hc031da28, 32'hc110c175} /* (21, 14, 30) {real, imag} */,
  {32'h40528106, 32'h4194c968} /* (21, 14, 29) {real, imag} */,
  {32'h3f840a18, 32'hc08642f6} /* (21, 14, 28) {real, imag} */,
  {32'hc1662c31, 32'hbf919354} /* (21, 14, 27) {real, imag} */,
  {32'hc0d1bbac, 32'hbebb5a68} /* (21, 14, 26) {real, imag} */,
  {32'hc0d3383e, 32'h411a77b4} /* (21, 14, 25) {real, imag} */,
  {32'h40a2ec5e, 32'h40cba430} /* (21, 14, 24) {real, imag} */,
  {32'h41675310, 32'h4109e770} /* (21, 14, 23) {real, imag} */,
  {32'h3fe53542, 32'hc103e01d} /* (21, 14, 22) {real, imag} */,
  {32'hbfcfaf4e, 32'hc15321ea} /* (21, 14, 21) {real, imag} */,
  {32'h40bc3dff, 32'h4102c698} /* (21, 14, 20) {real, imag} */,
  {32'hc085d857, 32'h40225190} /* (21, 14, 19) {real, imag} */,
  {32'h41161200, 32'hbf9329a8} /* (21, 14, 18) {real, imag} */,
  {32'h40a72a7d, 32'hc0ae96d4} /* (21, 14, 17) {real, imag} */,
  {32'h40c91bbf, 32'h40008d99} /* (21, 14, 16) {real, imag} */,
  {32'hbee32b10, 32'hbf403184} /* (21, 14, 15) {real, imag} */,
  {32'h4016c336, 32'hc0d2912a} /* (21, 14, 14) {real, imag} */,
  {32'h40511fb8, 32'hc101c46a} /* (21, 14, 13) {real, imag} */,
  {32'hc0aa9ec9, 32'h40127052} /* (21, 14, 12) {real, imag} */,
  {32'hc096172e, 32'h3f7a0ce8} /* (21, 14, 11) {real, imag} */,
  {32'h4077e4cb, 32'hc16ec771} /* (21, 14, 10) {real, imag} */,
  {32'h3f1e89a0, 32'hc197bc89} /* (21, 14, 9) {real, imag} */,
  {32'hc13f1745, 32'hc0ceb832} /* (21, 14, 8) {real, imag} */,
  {32'h417128df, 32'h3fe98b6c} /* (21, 14, 7) {real, imag} */,
  {32'h3f4e51f4, 32'h40e5c16e} /* (21, 14, 6) {real, imag} */,
  {32'hc1164c67, 32'hc1797052} /* (21, 14, 5) {real, imag} */,
  {32'h4008aefe, 32'h40d9b87a} /* (21, 14, 4) {real, imag} */,
  {32'hc0949984, 32'h40ac60fc} /* (21, 14, 3) {real, imag} */,
  {32'h419f5c11, 32'hc1e38ce6} /* (21, 14, 2) {real, imag} */,
  {32'h4156df6e, 32'hc19ea27f} /* (21, 14, 1) {real, imag} */,
  {32'h41514afe, 32'h405587a1} /* (21, 14, 0) {real, imag} */,
  {32'hc11d1837, 32'h40bc1e38} /* (21, 13, 31) {real, imag} */,
  {32'hbea0dee0, 32'h410f43ad} /* (21, 13, 30) {real, imag} */,
  {32'hc0925fee, 32'h4197f368} /* (21, 13, 29) {real, imag} */,
  {32'h4115afc4, 32'hc117ab7f} /* (21, 13, 28) {real, imag} */,
  {32'h4023ad27, 32'hc154e6a8} /* (21, 13, 27) {real, imag} */,
  {32'h412f52eb, 32'hc156625c} /* (21, 13, 26) {real, imag} */,
  {32'hc0dfc442, 32'hc1960771} /* (21, 13, 25) {real, imag} */,
  {32'hc056e3d8, 32'h4119afae} /* (21, 13, 24) {real, imag} */,
  {32'h419116a0, 32'h4137c34c} /* (21, 13, 23) {real, imag} */,
  {32'hc08936f8, 32'h40b9f9dc} /* (21, 13, 22) {real, imag} */,
  {32'hc080f8c0, 32'hbf93bf28} /* (21, 13, 21) {real, imag} */,
  {32'hbda015c0, 32'hbff53af0} /* (21, 13, 20) {real, imag} */,
  {32'h3fbf2d80, 32'h4095f447} /* (21, 13, 19) {real, imag} */,
  {32'hc0bc5070, 32'h3fa056c4} /* (21, 13, 18) {real, imag} */,
  {32'h40b769aa, 32'h40680468} /* (21, 13, 17) {real, imag} */,
  {32'h3f6c8304, 32'h409f61e2} /* (21, 13, 16) {real, imag} */,
  {32'hbfdbb158, 32'h40ea7988} /* (21, 13, 15) {real, imag} */,
  {32'h4089797c, 32'hbfc8d9bc} /* (21, 13, 14) {real, imag} */,
  {32'h3f82a570, 32'h3f8f917c} /* (21, 13, 13) {real, imag} */,
  {32'hbe4648a0, 32'hc120fa0c} /* (21, 13, 12) {real, imag} */,
  {32'hc17d69f4, 32'h40b0b02e} /* (21, 13, 11) {real, imag} */,
  {32'h407d8548, 32'hc15fe86a} /* (21, 13, 10) {real, imag} */,
  {32'hc1c9ed0c, 32'hc1164f74} /* (21, 13, 9) {real, imag} */,
  {32'h4114b044, 32'h4082d394} /* (21, 13, 8) {real, imag} */,
  {32'hbb599400, 32'h41202f0a} /* (21, 13, 7) {real, imag} */,
  {32'hc0e7b45d, 32'hc1dd7822} /* (21, 13, 6) {real, imag} */,
  {32'h410550aa, 32'h4184f58a} /* (21, 13, 5) {real, imag} */,
  {32'h42006e3d, 32'h418c646e} /* (21, 13, 4) {real, imag} */,
  {32'h41b3df28, 32'hc1e1d8ea} /* (21, 13, 3) {real, imag} */,
  {32'h41a02180, 32'hc01ced28} /* (21, 13, 2) {real, imag} */,
  {32'h420061b8, 32'h419b7b61} /* (21, 13, 1) {real, imag} */,
  {32'hbf6157a4, 32'h41290c3f} /* (21, 13, 0) {real, imag} */,
  {32'hc0bf7c30, 32'h4171cc78} /* (21, 12, 31) {real, imag} */,
  {32'hc1768ade, 32'hc16f62b8} /* (21, 12, 30) {real, imag} */,
  {32'h41e28f0b, 32'h3fdc470c} /* (21, 12, 29) {real, imag} */,
  {32'hbf8bdfb0, 32'hc10c15ec} /* (21, 12, 28) {real, imag} */,
  {32'hc1465fc9, 32'hc2004b7b} /* (21, 12, 27) {real, imag} */,
  {32'h40ad8990, 32'hc122fad7} /* (21, 12, 26) {real, imag} */,
  {32'h4139c645, 32'h417fe1be} /* (21, 12, 25) {real, imag} */,
  {32'hc1804592, 32'hc12bcc23} /* (21, 12, 24) {real, imag} */,
  {32'hbe5cecc0, 32'hc09ec43c} /* (21, 12, 23) {real, imag} */,
  {32'hc09e478c, 32'hc1def39a} /* (21, 12, 22) {real, imag} */,
  {32'hc0c99786, 32'h401931b4} /* (21, 12, 21) {real, imag} */,
  {32'h411679ce, 32'h4102d17e} /* (21, 12, 20) {real, imag} */,
  {32'h40a8efdd, 32'h4124cd00} /* (21, 12, 19) {real, imag} */,
  {32'h410c0cee, 32'h410384f6} /* (21, 12, 18) {real, imag} */,
  {32'hc0a5c895, 32'h40dd82d0} /* (21, 12, 17) {real, imag} */,
  {32'hc09a0e62, 32'h4040c5c4} /* (21, 12, 16) {real, imag} */,
  {32'h4065686e, 32'hc09c107c} /* (21, 12, 15) {real, imag} */,
  {32'hc0c3d695, 32'hbf15e018} /* (21, 12, 14) {real, imag} */,
  {32'h4107a436, 32'hc0a34755} /* (21, 12, 13) {real, imag} */,
  {32'hc09ab1da, 32'h413cee3e} /* (21, 12, 12) {real, imag} */,
  {32'h40d3998e, 32'hbf906f78} /* (21, 12, 11) {real, imag} */,
  {32'hc1c458c7, 32'hc1544aac} /* (21, 12, 10) {real, imag} */,
  {32'hc1c34c36, 32'h40dfc2a0} /* (21, 12, 9) {real, imag} */,
  {32'h40732566, 32'hc158c08d} /* (21, 12, 8) {real, imag} */,
  {32'h407249f4, 32'hc0684dd0} /* (21, 12, 7) {real, imag} */,
  {32'hc1e9a75e, 32'h414e3ee1} /* (21, 12, 6) {real, imag} */,
  {32'h41bf2650, 32'h41018c28} /* (21, 12, 5) {real, imag} */,
  {32'hc15f6597, 32'h41005cc2} /* (21, 12, 4) {real, imag} */,
  {32'hbf9fadd0, 32'hc16a91f0} /* (21, 12, 3) {real, imag} */,
  {32'h4184859d, 32'hc07c7b22} /* (21, 12, 2) {real, imag} */,
  {32'h3fb47ff2, 32'hc0a7e1b4} /* (21, 12, 1) {real, imag} */,
  {32'hc1d45020, 32'h4194377c} /* (21, 12, 0) {real, imag} */,
  {32'h41c00fbd, 32'hc20bf7ea} /* (21, 11, 31) {real, imag} */,
  {32'h41ba0e2e, 32'h412d9754} /* (21, 11, 30) {real, imag} */,
  {32'hc2110034, 32'h418cd817} /* (21, 11, 29) {real, imag} */,
  {32'h417e0296, 32'hc1b26d3e} /* (21, 11, 28) {real, imag} */,
  {32'h40cd5472, 32'hc199b16e} /* (21, 11, 27) {real, imag} */,
  {32'hc194e0fd, 32'h4186c57c} /* (21, 11, 26) {real, imag} */,
  {32'h41a10039, 32'h3f062260} /* (21, 11, 25) {real, imag} */,
  {32'hc0e06018, 32'h3f170580} /* (21, 11, 24) {real, imag} */,
  {32'h4168bc44, 32'h3d168c00} /* (21, 11, 23) {real, imag} */,
  {32'hc0f53d72, 32'h40d56dff} /* (21, 11, 22) {real, imag} */,
  {32'hc1090e1f, 32'h4062ba88} /* (21, 11, 21) {real, imag} */,
  {32'hc07e8479, 32'hc175e860} /* (21, 11, 20) {real, imag} */,
  {32'h409be090, 32'h40903dc4} /* (21, 11, 19) {real, imag} */,
  {32'hc03f1ca6, 32'h3f776760} /* (21, 11, 18) {real, imag} */,
  {32'h4085bb76, 32'h409c38b0} /* (21, 11, 17) {real, imag} */,
  {32'hc132d93a, 32'hc0257db6} /* (21, 11, 16) {real, imag} */,
  {32'hc09e2f3a, 32'h3f7bfa80} /* (21, 11, 15) {real, imag} */,
  {32'h4019c172, 32'hc1358f81} /* (21, 11, 14) {real, imag} */,
  {32'h40982b64, 32'h4082a33c} /* (21, 11, 13) {real, imag} */,
  {32'h3fb898ce, 32'hc0930e81} /* (21, 11, 12) {real, imag} */,
  {32'h40788245, 32'hbe0d7d80} /* (21, 11, 11) {real, imag} */,
  {32'h3d978360, 32'hc0a531c7} /* (21, 11, 10) {real, imag} */,
  {32'h40bce661, 32'hc1adf12a} /* (21, 11, 9) {real, imag} */,
  {32'hc2062f36, 32'h416302e8} /* (21, 11, 8) {real, imag} */,
  {32'h417eb9da, 32'h42239c34} /* (21, 11, 7) {real, imag} */,
  {32'h41c84b37, 32'hc11a76a3} /* (21, 11, 6) {real, imag} */,
  {32'hc0e91212, 32'hc11d86eb} /* (21, 11, 5) {real, imag} */,
  {32'hc1dd5bf5, 32'hbfc66b60} /* (21, 11, 4) {real, imag} */,
  {32'h416bfbee, 32'h4254d5e8} /* (21, 11, 3) {real, imag} */,
  {32'h406aae7c, 32'h41182140} /* (21, 11, 2) {real, imag} */,
  {32'hc1ceacf7, 32'hc2531e3e} /* (21, 11, 1) {real, imag} */,
  {32'hc239f3d6, 32'hbfbcd2e4} /* (21, 11, 0) {real, imag} */,
  {32'hbfc12aa9, 32'h411ab53a} /* (21, 10, 31) {real, imag} */,
  {32'hc03a644e, 32'h40d5a9ae} /* (21, 10, 30) {real, imag} */,
  {32'h414434a6, 32'h3f3e1c08} /* (21, 10, 29) {real, imag} */,
  {32'hc18a684e, 32'h3fcb47f0} /* (21, 10, 28) {real, imag} */,
  {32'hc1f32f7c, 32'h4140f8ae} /* (21, 10, 27) {real, imag} */,
  {32'h41e4c802, 32'hc18c10d6} /* (21, 10, 26) {real, imag} */,
  {32'h418524bc, 32'h3fd93bf0} /* (21, 10, 25) {real, imag} */,
  {32'h41c4d3a0, 32'hc1b51c80} /* (21, 10, 24) {real, imag} */,
  {32'hc1443090, 32'h420a025d} /* (21, 10, 23) {real, imag} */,
  {32'h4180d530, 32'hbcb6e100} /* (21, 10, 22) {real, imag} */,
  {32'h41a22179, 32'h3f2ee670} /* (21, 10, 21) {real, imag} */,
  {32'hc14de526, 32'h3ec59a88} /* (21, 10, 20) {real, imag} */,
  {32'h3d0d1400, 32'hc16de2b5} /* (21, 10, 19) {real, imag} */,
  {32'hc0e7eecc, 32'hc189c7a1} /* (21, 10, 18) {real, imag} */,
  {32'hbefe4f58, 32'hc147a950} /* (21, 10, 17) {real, imag} */,
  {32'hc0f4a720, 32'h3fa52f34} /* (21, 10, 16) {real, imag} */,
  {32'hc09afef4, 32'hbd3b9780} /* (21, 10, 15) {real, imag} */,
  {32'h41ee7dd1, 32'h411b8c20} /* (21, 10, 14) {real, imag} */,
  {32'hc0ecfb42, 32'hc05d419c} /* (21, 10, 13) {real, imag} */,
  {32'hc10d758c, 32'h408cc6b0} /* (21, 10, 12) {real, imag} */,
  {32'hbffecff0, 32'h41b391b6} /* (21, 10, 11) {real, imag} */,
  {32'hc182a792, 32'h40158642} /* (21, 10, 10) {real, imag} */,
  {32'hc116cfd8, 32'hc22c84c5} /* (21, 10, 9) {real, imag} */,
  {32'h420c3be8, 32'hc090fa8c} /* (21, 10, 8) {real, imag} */,
  {32'h41c3c21a, 32'hc03a21e8} /* (21, 10, 7) {real, imag} */,
  {32'h41c0743e, 32'hc1a58562} /* (21, 10, 6) {real, imag} */,
  {32'h41f4027c, 32'hc1e3d9d9} /* (21, 10, 5) {real, imag} */,
  {32'hc241173b, 32'hc16ead7a} /* (21, 10, 4) {real, imag} */,
  {32'hc12d0ac2, 32'hc170e4ac} /* (21, 10, 3) {real, imag} */,
  {32'h405d647a, 32'h419ae988} /* (21, 10, 2) {real, imag} */,
  {32'h4000e0c2, 32'h424c660a} /* (21, 10, 1) {real, imag} */,
  {32'h406ae998, 32'hc1487578} /* (21, 10, 0) {real, imag} */,
  {32'hc1d527e4, 32'hc1aa1af6} /* (21, 9, 31) {real, imag} */,
  {32'hc1e6b4f1, 32'hc0e85f70} /* (21, 9, 30) {real, imag} */,
  {32'hc1060800, 32'hc23167b7} /* (21, 9, 29) {real, imag} */,
  {32'hc11a9b86, 32'h418ab6f8} /* (21, 9, 28) {real, imag} */,
  {32'hc1fa393c, 32'h42179d93} /* (21, 9, 27) {real, imag} */,
  {32'h419c29a4, 32'hc150e76e} /* (21, 9, 26) {real, imag} */,
  {32'h4127f644, 32'hc17007d4} /* (21, 9, 25) {real, imag} */,
  {32'h41e809a7, 32'hc1bf3866} /* (21, 9, 24) {real, imag} */,
  {32'h41d4a82e, 32'hbf26ef88} /* (21, 9, 23) {real, imag} */,
  {32'h4024f070, 32'hc14c64c4} /* (21, 9, 22) {real, imag} */,
  {32'h40ae5b1e, 32'h41855748} /* (21, 9, 21) {real, imag} */,
  {32'hbf9cfa74, 32'h40d772a1} /* (21, 9, 20) {real, imag} */,
  {32'h3fc145a4, 32'hc01be8fc} /* (21, 9, 19) {real, imag} */,
  {32'h400b05b2, 32'hbfb17530} /* (21, 9, 18) {real, imag} */,
  {32'hc0ccb020, 32'hc0b1947d} /* (21, 9, 17) {real, imag} */,
  {32'h40d6b485, 32'hc0bac172} /* (21, 9, 16) {real, imag} */,
  {32'h4075afb4, 32'h4055dd0a} /* (21, 9, 15) {real, imag} */,
  {32'hc1449150, 32'hbfa06b40} /* (21, 9, 14) {real, imag} */,
  {32'hc12d6180, 32'h40a4461a} /* (21, 9, 13) {real, imag} */,
  {32'h4089abdd, 32'hc038edbe} /* (21, 9, 12) {real, imag} */,
  {32'hc1802b26, 32'hc14b884b} /* (21, 9, 11) {real, imag} */,
  {32'h41eff376, 32'h414157a8} /* (21, 9, 10) {real, imag} */,
  {32'h4190c7ee, 32'h4132a712} /* (21, 9, 9) {real, imag} */,
  {32'h4170bf8a, 32'hc15285f4} /* (21, 9, 8) {real, imag} */,
  {32'hc2137219, 32'hc17f32c6} /* (21, 9, 7) {real, imag} */,
  {32'h41f87a04, 32'h41ec6153} /* (21, 9, 6) {real, imag} */,
  {32'hc1eb4770, 32'h413f9a3c} /* (21, 9, 5) {real, imag} */,
  {32'hc1ab045d, 32'h41497743} /* (21, 9, 4) {real, imag} */,
  {32'h4201c438, 32'h4158ca97} /* (21, 9, 3) {real, imag} */,
  {32'hc29449a8, 32'hc2472b46} /* (21, 9, 2) {real, imag} */,
  {32'hc0b1d9d0, 32'hc14d79f0} /* (21, 9, 1) {real, imag} */,
  {32'h4166de3e, 32'h417134df} /* (21, 9, 0) {real, imag} */,
  {32'hc20d9900, 32'hc258d795} /* (21, 8, 31) {real, imag} */,
  {32'h425ef466, 32'hc233c9a3} /* (21, 8, 30) {real, imag} */,
  {32'h4143f98c, 32'h400e95b8} /* (21, 8, 29) {real, imag} */,
  {32'h4201e131, 32'h419028e8} /* (21, 8, 28) {real, imag} */,
  {32'hbfa40a40, 32'hc1138048} /* (21, 8, 27) {real, imag} */,
  {32'h428bbc57, 32'h41218d29} /* (21, 8, 26) {real, imag} */,
  {32'h41ca8d28, 32'hc221d34c} /* (21, 8, 25) {real, imag} */,
  {32'h4129f5f6, 32'h41b181ff} /* (21, 8, 24) {real, imag} */,
  {32'hc2244e90, 32'hc18a12c1} /* (21, 8, 23) {real, imag} */,
  {32'hc12632d2, 32'hc1bb1ca2} /* (21, 8, 22) {real, imag} */,
  {32'hc18a7adb, 32'h406d1144} /* (21, 8, 21) {real, imag} */,
  {32'hc08824c2, 32'h41108fb8} /* (21, 8, 20) {real, imag} */,
  {32'h41653eb9, 32'h40866811} /* (21, 8, 19) {real, imag} */,
  {32'hbdb6cb80, 32'h3ec083a0} /* (21, 8, 18) {real, imag} */,
  {32'h40bd637b, 32'h402f4e0c} /* (21, 8, 17) {real, imag} */,
  {32'h4145b57c, 32'hc14e7ab6} /* (21, 8, 16) {real, imag} */,
  {32'hc036f746, 32'h3ff916d8} /* (21, 8, 15) {real, imag} */,
  {32'hc1163667, 32'h40ffa5ce} /* (21, 8, 14) {real, imag} */,
  {32'h40fe12d6, 32'h41921d7c} /* (21, 8, 13) {real, imag} */,
  {32'hc1411c0f, 32'h40436292} /* (21, 8, 12) {real, imag} */,
  {32'hc0aca659, 32'hc04739ac} /* (21, 8, 11) {real, imag} */,
  {32'h41864f6b, 32'hc1140210} /* (21, 8, 10) {real, imag} */,
  {32'hc0e5ed30, 32'hc0fe76f4} /* (21, 8, 9) {real, imag} */,
  {32'hc20654dc, 32'h415a359e} /* (21, 8, 8) {real, imag} */,
  {32'hc1cded48, 32'h422e9366} /* (21, 8, 7) {real, imag} */,
  {32'hc217da00, 32'h4027f260} /* (21, 8, 6) {real, imag} */,
  {32'h42261b36, 32'h420a68c3} /* (21, 8, 5) {real, imag} */,
  {32'h40d5acb6, 32'hc237095b} /* (21, 8, 4) {real, imag} */,
  {32'h420949d2, 32'h420615c6} /* (21, 8, 3) {real, imag} */,
  {32'hc25935be, 32'hc1a99542} /* (21, 8, 2) {real, imag} */,
  {32'hc1a93e84, 32'h40aa7c48} /* (21, 8, 1) {real, imag} */,
  {32'hc24ffd39, 32'hc298cf35} /* (21, 8, 0) {real, imag} */,
  {32'hc20ad1ca, 32'hc07d37ae} /* (21, 7, 31) {real, imag} */,
  {32'h40f9421a, 32'h4239d33e} /* (21, 7, 30) {real, imag} */,
  {32'hc0e170b6, 32'hc12a76db} /* (21, 7, 29) {real, imag} */,
  {32'h41e4aae4, 32'hc198b6c5} /* (21, 7, 28) {real, imag} */,
  {32'h41c26285, 32'h426e96ba} /* (21, 7, 27) {real, imag} */,
  {32'hc201cd27, 32'h426d8d9c} /* (21, 7, 26) {real, imag} */,
  {32'h3e6eed80, 32'hc1b3edf9} /* (21, 7, 25) {real, imag} */,
  {32'h41ed3a45, 32'h418d0b4d} /* (21, 7, 24) {real, imag} */,
  {32'hc19ab7a5, 32'h413765de} /* (21, 7, 23) {real, imag} */,
  {32'h41ba7b48, 32'h41c1ac10} /* (21, 7, 22) {real, imag} */,
  {32'h402cd07a, 32'hc12b2521} /* (21, 7, 21) {real, imag} */,
  {32'hbdc55280, 32'hc1988af7} /* (21, 7, 20) {real, imag} */,
  {32'hbfa2a45c, 32'h409b4430} /* (21, 7, 19) {real, imag} */,
  {32'hc0b6b6c8, 32'hbfe35dc8} /* (21, 7, 18) {real, imag} */,
  {32'hc10f7018, 32'hc1ba790c} /* (21, 7, 17) {real, imag} */,
  {32'h3d8c6d00, 32'hbf9d8c30} /* (21, 7, 16) {real, imag} */,
  {32'h41275060, 32'hc131d287} /* (21, 7, 15) {real, imag} */,
  {32'hc1909170, 32'h4147f7c5} /* (21, 7, 14) {real, imag} */,
  {32'h41359a02, 32'hc00b3b80} /* (21, 7, 13) {real, imag} */,
  {32'h41805aba, 32'h41b9158d} /* (21, 7, 12) {real, imag} */,
  {32'hc0307bb6, 32'h41068599} /* (21, 7, 11) {real, imag} */,
  {32'hc13db709, 32'hc187b74e} /* (21, 7, 10) {real, imag} */,
  {32'hc1511aca, 32'h41a5c251} /* (21, 7, 9) {real, imag} */,
  {32'h41438c02, 32'hc1b81b47} /* (21, 7, 8) {real, imag} */,
  {32'hc176e71a, 32'hc1870b93} /* (21, 7, 7) {real, imag} */,
  {32'hc222b267, 32'hc18a9b8f} /* (21, 7, 6) {real, imag} */,
  {32'hc1854235, 32'h41ab69e4} /* (21, 7, 5) {real, imag} */,
  {32'hc03a133c, 32'h4140280e} /* (21, 7, 4) {real, imag} */,
  {32'hc1a14948, 32'hc20bb1f7} /* (21, 7, 3) {real, imag} */,
  {32'hbf8de828, 32'h4179348d} /* (21, 7, 2) {real, imag} */,
  {32'h41ea7214, 32'hc0e5e9e9} /* (21, 7, 1) {real, imag} */,
  {32'h426a3984, 32'hc1d3deef} /* (21, 7, 0) {real, imag} */,
  {32'hc1958bb8, 32'hc1be6579} /* (21, 6, 31) {real, imag} */,
  {32'hc183f9be, 32'h4208374d} /* (21, 6, 30) {real, imag} */,
  {32'hc205ae7b, 32'hc1a82389} /* (21, 6, 29) {real, imag} */,
  {32'hc18458dc, 32'h41b82548} /* (21, 6, 28) {real, imag} */,
  {32'hc247138e, 32'h420bbf44} /* (21, 6, 27) {real, imag} */,
  {32'h420d0bd7, 32'h418a9c4a} /* (21, 6, 26) {real, imag} */,
  {32'hc0916fa8, 32'hc05432e8} /* (21, 6, 25) {real, imag} */,
  {32'h41c67344, 32'h421db5ab} /* (21, 6, 24) {real, imag} */,
  {32'h4270e7d0, 32'hc1ff895c} /* (21, 6, 23) {real, imag} */,
  {32'hc043c252, 32'hc1bd28da} /* (21, 6, 22) {real, imag} */,
  {32'hc150d5a8, 32'hc138563c} /* (21, 6, 21) {real, imag} */,
  {32'h414395f7, 32'h40a2916b} /* (21, 6, 20) {real, imag} */,
  {32'h411ca126, 32'hc14ddaa4} /* (21, 6, 19) {real, imag} */,
  {32'h40eafa18, 32'h41ae30f6} /* (21, 6, 18) {real, imag} */,
  {32'hc18ab08c, 32'h3f64c758} /* (21, 6, 17) {real, imag} */,
  {32'hc106efa0, 32'hc09e4400} /* (21, 6, 16) {real, imag} */,
  {32'h41463c53, 32'hc1306b92} /* (21, 6, 15) {real, imag} */,
  {32'hc151119c, 32'h41be564e} /* (21, 6, 14) {real, imag} */,
  {32'hc13cb9ca, 32'hc128edc8} /* (21, 6, 13) {real, imag} */,
  {32'hc18660d4, 32'hc1138002} /* (21, 6, 12) {real, imag} */,
  {32'h41d045e0, 32'hc1db22aa} /* (21, 6, 11) {real, imag} */,
  {32'h408a370d, 32'h404c2974} /* (21, 6, 10) {real, imag} */,
  {32'hc0b39920, 32'h41ab9bfe} /* (21, 6, 9) {real, imag} */,
  {32'hc1296658, 32'hc0fe0046} /* (21, 6, 8) {real, imag} */,
  {32'h42277ea5, 32'h41ff8399} /* (21, 6, 7) {real, imag} */,
  {32'h41a1969a, 32'h41582df1} /* (21, 6, 6) {real, imag} */,
  {32'h419e81d4, 32'h40235c08} /* (21, 6, 5) {real, imag} */,
  {32'h42515cbe, 32'hc248e2d8} /* (21, 6, 4) {real, imag} */,
  {32'hc2073a15, 32'hc25e2b1c} /* (21, 6, 3) {real, imag} */,
  {32'hc289fc6e, 32'h42b7a09a} /* (21, 6, 2) {real, imag} */,
  {32'h4155eff0, 32'h425212c8} /* (21, 6, 1) {real, imag} */,
  {32'h42291b32, 32'hc238cd32} /* (21, 6, 0) {real, imag} */,
  {32'hc1f9600c, 32'hc0b73e48} /* (21, 5, 31) {real, imag} */,
  {32'h41a61e76, 32'h431715bf} /* (21, 5, 30) {real, imag} */,
  {32'h4114d3bc, 32'hc17563fd} /* (21, 5, 29) {real, imag} */,
  {32'hc1da71c3, 32'h41c0ead3} /* (21, 5, 28) {real, imag} */,
  {32'hc1678428, 32'h425e6348} /* (21, 5, 27) {real, imag} */,
  {32'hc0f2b058, 32'hc265d54c} /* (21, 5, 26) {real, imag} */,
  {32'hc1937e91, 32'hc2185611} /* (21, 5, 25) {real, imag} */,
  {32'h42157e7d, 32'h417a71d6} /* (21, 5, 24) {real, imag} */,
  {32'h41a31bd0, 32'hc0e8a2a2} /* (21, 5, 23) {real, imag} */,
  {32'hc1a339e6, 32'h419b1f30} /* (21, 5, 22) {real, imag} */,
  {32'hc1149908, 32'hc14ae0dd} /* (21, 5, 21) {real, imag} */,
  {32'h412d9572, 32'h3ffe4e90} /* (21, 5, 20) {real, imag} */,
  {32'h413f8c51, 32'h40bdd6de} /* (21, 5, 19) {real, imag} */,
  {32'hc0414ab0, 32'h3ebb7680} /* (21, 5, 18) {real, imag} */,
  {32'hc10a08dd, 32'hbf538650} /* (21, 5, 17) {real, imag} */,
  {32'h41213b06, 32'hbfc92160} /* (21, 5, 16) {real, imag} */,
  {32'h41ad5810, 32'hc1be5300} /* (21, 5, 15) {real, imag} */,
  {32'h40919668, 32'hc1342a24} /* (21, 5, 14) {real, imag} */,
  {32'h409cf91e, 32'h410ba4db} /* (21, 5, 13) {real, imag} */,
  {32'hc117868e, 32'hc1341fde} /* (21, 5, 12) {real, imag} */,
  {32'h3fe8b840, 32'hc193f00e} /* (21, 5, 11) {real, imag} */,
  {32'h40eeb320, 32'h420a779c} /* (21, 5, 10) {real, imag} */,
  {32'h41b24884, 32'hc11023e9} /* (21, 5, 9) {real, imag} */,
  {32'h4242c687, 32'hc2104904} /* (21, 5, 8) {real, imag} */,
  {32'hc18a63b3, 32'h428b4743} /* (21, 5, 7) {real, imag} */,
  {32'hc22bb07a, 32'hc1796038} /* (21, 5, 6) {real, imag} */,
  {32'h42d37433, 32'hbf05fc80} /* (21, 5, 5) {real, imag} */,
  {32'h418c2d41, 32'h3d747600} /* (21, 5, 4) {real, imag} */,
  {32'hc1c0c492, 32'h422b1cfe} /* (21, 5, 3) {real, imag} */,
  {32'hc2722a9f, 32'h41d8b8a2} /* (21, 5, 2) {real, imag} */,
  {32'hc1befc9c, 32'hc2aa75e4} /* (21, 5, 1) {real, imag} */,
  {32'hc257f2c6, 32'hc2c22abe} /* (21, 5, 0) {real, imag} */,
  {32'hc1091692, 32'hc1e1613c} /* (21, 4, 31) {real, imag} */,
  {32'hc292191a, 32'hc213bc2e} /* (21, 4, 30) {real, imag} */,
  {32'h4278e642, 32'h431af20a} /* (21, 4, 29) {real, imag} */,
  {32'hc0d9dfdb, 32'h41041722} /* (21, 4, 28) {real, imag} */,
  {32'h418cccf6, 32'hc1b9b2ea} /* (21, 4, 27) {real, imag} */,
  {32'hc12075e8, 32'h41e891a4} /* (21, 4, 26) {real, imag} */,
  {32'h41b365e9, 32'h42481fc9} /* (21, 4, 25) {real, imag} */,
  {32'hc217217a, 32'hc153dfa0} /* (21, 4, 24) {real, imag} */,
  {32'hc235742b, 32'h3f984040} /* (21, 4, 23) {real, imag} */,
  {32'hc107a22d, 32'h4098c42a} /* (21, 4, 22) {real, imag} */,
  {32'h41656e4c, 32'h40f8da08} /* (21, 4, 21) {real, imag} */,
  {32'h41550b62, 32'h3e9485b4} /* (21, 4, 20) {real, imag} */,
  {32'hc199fa6b, 32'hc1af7451} /* (21, 4, 19) {real, imag} */,
  {32'hc18e983c, 32'h408dbdae} /* (21, 4, 18) {real, imag} */,
  {32'hbf532120, 32'h40b45ad4} /* (21, 4, 17) {real, imag} */,
  {32'h417597ca, 32'hc1c293e5} /* (21, 4, 16) {real, imag} */,
  {32'hc14fa39a, 32'h4106753c} /* (21, 4, 15) {real, imag} */,
  {32'h4009709e, 32'hc1acfb1c} /* (21, 4, 14) {real, imag} */,
  {32'h4173d2f2, 32'h402819c8} /* (21, 4, 13) {real, imag} */,
  {32'hc12bfeca, 32'hbf003d7a} /* (21, 4, 12) {real, imag} */,
  {32'hbff88d10, 32'h409eb260} /* (21, 4, 11) {real, imag} */,
  {32'h41c08c6e, 32'h4201a738} /* (21, 4, 10) {real, imag} */,
  {32'h417140f8, 32'h41c6dffc} /* (21, 4, 9) {real, imag} */,
  {32'hc23b89de, 32'hc21fd586} /* (21, 4, 8) {real, imag} */,
  {32'hc0ce6f33, 32'h40e67b98} /* (21, 4, 7) {real, imag} */,
  {32'h4269aa88, 32'h4220d592} /* (21, 4, 6) {real, imag} */,
  {32'h4155d43a, 32'h422199c0} /* (21, 4, 5) {real, imag} */,
  {32'hc1b12839, 32'h4161a820} /* (21, 4, 4) {real, imag} */,
  {32'hc168265e, 32'h425b00d2} /* (21, 4, 3) {real, imag} */,
  {32'h42cbb9c2, 32'h4200d026} /* (21, 4, 2) {real, imag} */,
  {32'h428494e3, 32'hc0dd209e} /* (21, 4, 1) {real, imag} */,
  {32'h4029384a, 32'h3f3632a0} /* (21, 4, 0) {real, imag} */,
  {32'hc209c4f8, 32'h420e8660} /* (21, 3, 31) {real, imag} */,
  {32'hc1778c28, 32'hc30501ca} /* (21, 3, 30) {real, imag} */,
  {32'h41d250d0, 32'hc18821d1} /* (21, 3, 29) {real, imag} */,
  {32'h41469f1e, 32'h41d09cec} /* (21, 3, 28) {real, imag} */,
  {32'h41f74d38, 32'h420ba125} /* (21, 3, 27) {real, imag} */,
  {32'hc1efaed4, 32'h42273786} /* (21, 3, 26) {real, imag} */,
  {32'h4120ee15, 32'hc2a325d8} /* (21, 3, 25) {real, imag} */,
  {32'hc1b61d0f, 32'hc19e34b1} /* (21, 3, 24) {real, imag} */,
  {32'hc242363e, 32'hc1221d58} /* (21, 3, 23) {real, imag} */,
  {32'h424354a6, 32'hc02cc80c} /* (21, 3, 22) {real, imag} */,
  {32'hc0e02ae2, 32'h40fe7556} /* (21, 3, 21) {real, imag} */,
  {32'h406a91e0, 32'h40812f46} /* (21, 3, 20) {real, imag} */,
  {32'h4204566e, 32'h410b65f0} /* (21, 3, 19) {real, imag} */,
  {32'hc1c31ebc, 32'hc0985e28} /* (21, 3, 18) {real, imag} */,
  {32'h410b1071, 32'h409ca81c} /* (21, 3, 17) {real, imag} */,
  {32'h41b62bef, 32'h4219b96c} /* (21, 3, 16) {real, imag} */,
  {32'hc1877264, 32'h41878241} /* (21, 3, 15) {real, imag} */,
  {32'h40a1317a, 32'h3f8f0860} /* (21, 3, 14) {real, imag} */,
  {32'h41144b29, 32'hc12725a2} /* (21, 3, 13) {real, imag} */,
  {32'hc1ad45d0, 32'h41e9c514} /* (21, 3, 12) {real, imag} */,
  {32'hc1867d40, 32'h406e61e4} /* (21, 3, 11) {real, imag} */,
  {32'h41a72fb4, 32'hbf01a550} /* (21, 3, 10) {real, imag} */,
  {32'hc0331c68, 32'h41d48e92} /* (21, 3, 9) {real, imag} */,
  {32'hc19ccc8b, 32'hc259d41a} /* (21, 3, 8) {real, imag} */,
  {32'hc06f3524, 32'hc1d1bff7} /* (21, 3, 7) {real, imag} */,
  {32'h41e08b3c, 32'h410cbc80} /* (21, 3, 6) {real, imag} */,
  {32'h4299076e, 32'h423ead4f} /* (21, 3, 5) {real, imag} */,
  {32'h40fe284c, 32'h423b74ae} /* (21, 3, 4) {real, imag} */,
  {32'hc1c972a4, 32'h4131a814} /* (21, 3, 3) {real, imag} */,
  {32'h425c8434, 32'hc2d60e7f} /* (21, 3, 2) {real, imag} */,
  {32'h4187a394, 32'h42bf0c42} /* (21, 3, 1) {real, imag} */,
  {32'h41a25bbb, 32'hc2329aaa} /* (21, 3, 0) {real, imag} */,
  {32'hc342f9f4, 32'hc29c5ac1} /* (21, 2, 31) {real, imag} */,
  {32'h432cbf0b, 32'h42b403f1} /* (21, 2, 30) {real, imag} */,
  {32'hc2acd15c, 32'hc1e1c09c} /* (21, 2, 29) {real, imag} */,
  {32'hc22aa37e, 32'h423a763f} /* (21, 2, 28) {real, imag} */,
  {32'h3ef690a0, 32'h416465dc} /* (21, 2, 27) {real, imag} */,
  {32'hc222ce93, 32'hc0fdd178} /* (21, 2, 26) {real, imag} */,
  {32'h42509d80, 32'hc0c90990} /* (21, 2, 25) {real, imag} */,
  {32'h42106616, 32'h415a49dc} /* (21, 2, 24) {real, imag} */,
  {32'hc2134392, 32'hc0781610} /* (21, 2, 23) {real, imag} */,
  {32'h400d8d50, 32'h41574148} /* (21, 2, 22) {real, imag} */,
  {32'hc10f7f75, 32'h41ad5d8e} /* (21, 2, 21) {real, imag} */,
  {32'hc23d0e29, 32'hc1118dde} /* (21, 2, 20) {real, imag} */,
  {32'h41a049a5, 32'hc0cf7880} /* (21, 2, 19) {real, imag} */,
  {32'h4000a638, 32'hc0c77314} /* (21, 2, 18) {real, imag} */,
  {32'h3fa37f50, 32'h417cf38c} /* (21, 2, 17) {real, imag} */,
  {32'h4000b478, 32'hc11af9d4} /* (21, 2, 16) {real, imag} */,
  {32'h41a4b153, 32'hc182b872} /* (21, 2, 15) {real, imag} */,
  {32'h4133eb32, 32'h41b6815b} /* (21, 2, 14) {real, imag} */,
  {32'h415358b2, 32'hc1c1dbec} /* (21, 2, 13) {real, imag} */,
  {32'h410dfc94, 32'h413959ea} /* (21, 2, 12) {real, imag} */,
  {32'hc0db6ad2, 32'h41fb6fc6} /* (21, 2, 11) {real, imag} */,
  {32'h425decc9, 32'hc1ce6620} /* (21, 2, 10) {real, imag} */,
  {32'h4209f95e, 32'h4163660c} /* (21, 2, 9) {real, imag} */,
  {32'h41db79fb, 32'h41ff6c82} /* (21, 2, 8) {real, imag} */,
  {32'h417297c2, 32'h42205430} /* (21, 2, 7) {real, imag} */,
  {32'h41c051ba, 32'h42dbbbd6} /* (21, 2, 6) {real, imag} */,
  {32'hc1d462d0, 32'h41c3a18e} /* (21, 2, 5) {real, imag} */,
  {32'h42ae31b9, 32'hc238a279} /* (21, 2, 4) {real, imag} */,
  {32'hc20e2f6b, 32'h42732c48} /* (21, 2, 3) {real, imag} */,
  {32'h42eba64d, 32'h40ce61f0} /* (21, 2, 2) {real, imag} */,
  {32'hc280c310, 32'hc294891f} /* (21, 2, 1) {real, imag} */,
  {32'hc203b0f6, 32'hc2dd8ec8} /* (21, 2, 0) {real, imag} */,
  {32'h429548dc, 32'h42072222} /* (21, 1, 31) {real, imag} */,
  {32'h4215ff2b, 32'hc30131f6} /* (21, 1, 30) {real, imag} */,
  {32'h425760d4, 32'h42775eac} /* (21, 1, 29) {real, imag} */,
  {32'h3c5b7000, 32'h42a6146b} /* (21, 1, 28) {real, imag} */,
  {32'hc17f8794, 32'hc2caf0b9} /* (21, 1, 27) {real, imag} */,
  {32'h426435b3, 32'hc2124966} /* (21, 1, 26) {real, imag} */,
  {32'h416418b8, 32'h41fef04f} /* (21, 1, 25) {real, imag} */,
  {32'hc2096141, 32'h3f546ac0} /* (21, 1, 24) {real, imag} */,
  {32'h4246a48c, 32'hc25289b2} /* (21, 1, 23) {real, imag} */,
  {32'h4191dfb8, 32'h42297f7f} /* (21, 1, 22) {real, imag} */,
  {32'hc20b16b5, 32'h41b81a17} /* (21, 1, 21) {real, imag} */,
  {32'hc1fb9914, 32'hc0cd5031} /* (21, 1, 20) {real, imag} */,
  {32'h4143dfd2, 32'h41df5954} /* (21, 1, 19) {real, imag} */,
  {32'hc1e3a3e4, 32'hbef21840} /* (21, 1, 18) {real, imag} */,
  {32'h4189a693, 32'h4163f0a4} /* (21, 1, 17) {real, imag} */,
  {32'h40e2bd40, 32'hc0fc2c00} /* (21, 1, 16) {real, imag} */,
  {32'h4112317a, 32'hc196721e} /* (21, 1, 15) {real, imag} */,
  {32'hc0a76b00, 32'hc20280e0} /* (21, 1, 14) {real, imag} */,
  {32'h41d8a5d1, 32'hc15ccc25} /* (21, 1, 13) {real, imag} */,
  {32'hbf5dc880, 32'hc0cf60df} /* (21, 1, 12) {real, imag} */,
  {32'h41067405, 32'hc23658d0} /* (21, 1, 11) {real, imag} */,
  {32'hc22c252e, 32'hc1ef137a} /* (21, 1, 10) {real, imag} */,
  {32'hc2243c4c, 32'h41cae4a5} /* (21, 1, 9) {real, imag} */,
  {32'h41daf502, 32'hc142eb14} /* (21, 1, 8) {real, imag} */,
  {32'h4285bdf5, 32'h422f07c0} /* (21, 1, 7) {real, imag} */,
  {32'h42389141, 32'hc1a22481} /* (21, 1, 6) {real, imag} */,
  {32'hc1ef38fe, 32'h41a165d4} /* (21, 1, 5) {real, imag} */,
  {32'hc2bebe7a, 32'h42d7c4ad} /* (21, 1, 4) {real, imag} */,
  {32'hc0991804, 32'hc20d4bd0} /* (21, 1, 3) {real, imag} */,
  {32'hc289a43c, 32'hc3764092} /* (21, 1, 2) {real, imag} */,
  {32'h430d4776, 32'h4320538a} /* (21, 1, 1) {real, imag} */,
  {32'h4306ff40, 32'h4358d560} /* (21, 1, 0) {real, imag} */,
  {32'h430c8344, 32'h4296a9aa} /* (21, 0, 31) {real, imag} */,
  {32'hc1f89900, 32'h43049586} /* (21, 0, 30) {real, imag} */,
  {32'h420d6d40, 32'h400c4090} /* (21, 0, 29) {real, imag} */,
  {32'h42955309, 32'h415215ed} /* (21, 0, 28) {real, imag} */,
  {32'h4202091e, 32'hc228a50e} /* (21, 0, 27) {real, imag} */,
  {32'hc1da6568, 32'h40fd54cc} /* (21, 0, 26) {real, imag} */,
  {32'h420798e9, 32'h4260cba6} /* (21, 0, 25) {real, imag} */,
  {32'hc1dbc6f8, 32'hc18c5472} /* (21, 0, 24) {real, imag} */,
  {32'hc1de587b, 32'h41f82914} /* (21, 0, 23) {real, imag} */,
  {32'hc16a44b1, 32'h4108f04e} /* (21, 0, 22) {real, imag} */,
  {32'hc0c4be84, 32'h416c669b} /* (21, 0, 21) {real, imag} */,
  {32'h40e07e9e, 32'h4196b4f6} /* (21, 0, 20) {real, imag} */,
  {32'hc1d44cb6, 32'h41b1118d} /* (21, 0, 19) {real, imag} */,
  {32'h3f3eb4a0, 32'h421e6d29} /* (21, 0, 18) {real, imag} */,
  {32'hc1184d5c, 32'hc0d4afda} /* (21, 0, 17) {real, imag} */,
  {32'h411fbf1c, 32'h415a0d68} /* (21, 0, 16) {real, imag} */,
  {32'hc11270e4, 32'h41936a36} /* (21, 0, 15) {real, imag} */,
  {32'h4112c02a, 32'h40805108} /* (21, 0, 14) {real, imag} */,
  {32'hc12e1a53, 32'h408b0c24} /* (21, 0, 13) {real, imag} */,
  {32'h4137fa45, 32'h40dd1d5e} /* (21, 0, 12) {real, imag} */,
  {32'h413cc302, 32'hc1d0577e} /* (21, 0, 11) {real, imag} */,
  {32'hc151326d, 32'hc1dbb43f} /* (21, 0, 10) {real, imag} */,
  {32'hc24b90e2, 32'hc2883254} /* (21, 0, 9) {real, imag} */,
  {32'h42add182, 32'hc304da6b} /* (21, 0, 8) {real, imag} */,
  {32'hc1456aa0, 32'hc10d1200} /* (21, 0, 7) {real, imag} */,
  {32'h41ccfd96, 32'h4113d1da} /* (21, 0, 6) {real, imag} */,
  {32'hc28d778b, 32'h4259270c} /* (21, 0, 5) {real, imag} */,
  {32'h41884cec, 32'h41822081} /* (21, 0, 4) {real, imag} */,
  {32'h4213ceb4, 32'hc2e2f660} /* (21, 0, 3) {real, imag} */,
  {32'h42f23554, 32'hc1367684} /* (21, 0, 2) {real, imag} */,
  {32'h42a158cc, 32'h430f8097} /* (21, 0, 1) {real, imag} */,
  {32'h430043e7, 32'h429469d9} /* (21, 0, 0) {real, imag} */,
  {32'h41e34ff2, 32'hbed40fe8} /* (20, 31, 31) {real, imag} */,
  {32'h4266efe8, 32'h4226b880} /* (20, 31, 30) {real, imag} */,
  {32'h421f8336, 32'hc20d662b} /* (20, 31, 29) {real, imag} */,
  {32'hc2b2205a, 32'hc1830164} /* (20, 31, 28) {real, imag} */,
  {32'hc0fedd18, 32'hc2731924} /* (20, 31, 27) {real, imag} */,
  {32'hc0d1a6f0, 32'hc250536e} /* (20, 31, 26) {real, imag} */,
  {32'hc13f3a64, 32'hc1f523f8} /* (20, 31, 25) {real, imag} */,
  {32'h424551e5, 32'hc1df6e2a} /* (20, 31, 24) {real, imag} */,
  {32'hc19e981d, 32'hc1819cb2} /* (20, 31, 23) {real, imag} */,
  {32'hc11d4877, 32'h41ab14b2} /* (20, 31, 22) {real, imag} */,
  {32'h4198a855, 32'h41d99ad9} /* (20, 31, 21) {real, imag} */,
  {32'hc199d2c1, 32'hc18771ef} /* (20, 31, 20) {real, imag} */,
  {32'h418604e7, 32'h40db34d2} /* (20, 31, 19) {real, imag} */,
  {32'h3fa86e90, 32'h4011223e} /* (20, 31, 18) {real, imag} */,
  {32'h406580f0, 32'hc100be9a} /* (20, 31, 17) {real, imag} */,
  {32'h4151707c, 32'hc07cb834} /* (20, 31, 16) {real, imag} */,
  {32'h4146a46c, 32'h40974420} /* (20, 31, 15) {real, imag} */,
  {32'hc0eec0fc, 32'h40313dd2} /* (20, 31, 14) {real, imag} */,
  {32'h3f2bb800, 32'h41786197} /* (20, 31, 13) {real, imag} */,
  {32'hc1b2888b, 32'h41b86831} /* (20, 31, 12) {real, imag} */,
  {32'h4111e588, 32'hc13a6dce} /* (20, 31, 11) {real, imag} */,
  {32'hc137ed79, 32'hc1e0469c} /* (20, 31, 10) {real, imag} */,
  {32'h41494cee, 32'h411c767b} /* (20, 31, 9) {real, imag} */,
  {32'hc180c506, 32'hc1d502be} /* (20, 31, 8) {real, imag} */,
  {32'h417f75ca, 32'hc1126538} /* (20, 31, 7) {real, imag} */,
  {32'hc2270170, 32'h41e1e575} /* (20, 31, 6) {real, imag} */,
  {32'hc28d3774, 32'h41853187} /* (20, 31, 5) {real, imag} */,
  {32'hc2a43802, 32'hc2238ab3} /* (20, 31, 4) {real, imag} */,
  {32'h40f8a730, 32'hbf99aee0} /* (20, 31, 3) {real, imag} */,
  {32'h428b096e, 32'h41774362} /* (20, 31, 2) {real, imag} */,
  {32'hc20e69fb, 32'h3e98e8a8} /* (20, 31, 1) {real, imag} */,
  {32'h426444cd, 32'hc06c96b4} /* (20, 31, 0) {real, imag} */,
  {32'h422892a8, 32'hc2975bb0} /* (20, 30, 31) {real, imag} */,
  {32'hc1c7d76a, 32'hc27ed7d3} /* (20, 30, 30) {real, imag} */,
  {32'h41c3fc98, 32'h4232af90} /* (20, 30, 29) {real, imag} */,
  {32'hc09b192c, 32'h425f0f8b} /* (20, 30, 28) {real, imag} */,
  {32'hc1b12a42, 32'hc1cf2c1b} /* (20, 30, 27) {real, imag} */,
  {32'h427a63da, 32'hc244f425} /* (20, 30, 26) {real, imag} */,
  {32'h41173ada, 32'h42942507} /* (20, 30, 25) {real, imag} */,
  {32'hc210030d, 32'h425411ea} /* (20, 30, 24) {real, imag} */,
  {32'h3fdd9f78, 32'h42077f3a} /* (20, 30, 23) {real, imag} */,
  {32'hc1acded5, 32'h418ed25b} /* (20, 30, 22) {real, imag} */,
  {32'h41032a10, 32'h411a0bea} /* (20, 30, 21) {real, imag} */,
  {32'hc1f12470, 32'hc15e3cc2} /* (20, 30, 20) {real, imag} */,
  {32'h4159ea97, 32'h403f81fa} /* (20, 30, 19) {real, imag} */,
  {32'h4108958a, 32'h41d9faff} /* (20, 30, 18) {real, imag} */,
  {32'hc0b6c37c, 32'h40bbe1ea} /* (20, 30, 17) {real, imag} */,
  {32'h404b05d0, 32'h400f7028} /* (20, 30, 16) {real, imag} */,
  {32'h41b36c11, 32'hc127a75b} /* (20, 30, 15) {real, imag} */,
  {32'hc19de40b, 32'hc1a37c7d} /* (20, 30, 14) {real, imag} */,
  {32'hc11a1a77, 32'h41357e52} /* (20, 30, 13) {real, imag} */,
  {32'h3f3a0a00, 32'h41907c3f} /* (20, 30, 12) {real, imag} */,
  {32'h40990390, 32'hc235c908} /* (20, 30, 11) {real, imag} */,
  {32'hc1e94135, 32'h41eea461} /* (20, 30, 10) {real, imag} */,
  {32'hc1f92078, 32'h406b22b8} /* (20, 30, 9) {real, imag} */,
  {32'h41873e3a, 32'hc21b7c50} /* (20, 30, 8) {real, imag} */,
  {32'h40a84640, 32'h41259fee} /* (20, 30, 7) {real, imag} */,
  {32'hc2b2e8c9, 32'h41ac2086} /* (20, 30, 6) {real, imag} */,
  {32'h423a4e15, 32'hc103b742} /* (20, 30, 5) {real, imag} */,
  {32'h420fba02, 32'h41db6e9a} /* (20, 30, 4) {real, imag} */,
  {32'hc221c840, 32'hc232f214} /* (20, 30, 3) {real, imag} */,
  {32'hc1b59e44, 32'hc1ca6282} /* (20, 30, 2) {real, imag} */,
  {32'h400cbff8, 32'h428cfc5c} /* (20, 30, 1) {real, imag} */,
  {32'hc19f942a, 32'hc174a20e} /* (20, 30, 0) {real, imag} */,
  {32'hc1c08d70, 32'h42071902} /* (20, 29, 31) {real, imag} */,
  {32'h4285df3d, 32'h415bb1c7} /* (20, 29, 30) {real, imag} */,
  {32'hc2ab519a, 32'hc2333e0f} /* (20, 29, 29) {real, imag} */,
  {32'h417bde26, 32'h409ce198} /* (20, 29, 28) {real, imag} */,
  {32'h40b2572a, 32'hc235840f} /* (20, 29, 27) {real, imag} */,
  {32'hc14b6d7d, 32'h4280eeb7} /* (20, 29, 26) {real, imag} */,
  {32'hc1ce4934, 32'h41b20da8} /* (20, 29, 25) {real, imag} */,
  {32'h41a66de0, 32'hc082f797} /* (20, 29, 24) {real, imag} */,
  {32'hbf3eb990, 32'h422cef0a} /* (20, 29, 23) {real, imag} */,
  {32'h3f9e94e0, 32'hc18d088e} /* (20, 29, 22) {real, imag} */,
  {32'h42041b44, 32'h3e7c0900} /* (20, 29, 21) {real, imag} */,
  {32'hbfa7684c, 32'h409139b8} /* (20, 29, 20) {real, imag} */,
  {32'h3feea7c8, 32'hbfac148c} /* (20, 29, 19) {real, imag} */,
  {32'hc16cf65c, 32'h3f66f360} /* (20, 29, 18) {real, imag} */,
  {32'h41874b94, 32'hc1b61132} /* (20, 29, 17) {real, imag} */,
  {32'h3f26e920, 32'hc166657c} /* (20, 29, 16) {real, imag} */,
  {32'hc1081c51, 32'hc1473904} /* (20, 29, 15) {real, imag} */,
  {32'h4163de78, 32'hc02d9658} /* (20, 29, 14) {real, imag} */,
  {32'h4156f3c1, 32'hc0b2843b} /* (20, 29, 13) {real, imag} */,
  {32'h410bc5f8, 32'h411799ec} /* (20, 29, 12) {real, imag} */,
  {32'h42185788, 32'hc1dbd1e6} /* (20, 29, 11) {real, imag} */,
  {32'h4174ac5a, 32'h40503024} /* (20, 29, 10) {real, imag} */,
  {32'h40362a04, 32'hc0d731fc} /* (20, 29, 9) {real, imag} */,
  {32'h414b7880, 32'h410a9a58} /* (20, 29, 8) {real, imag} */,
  {32'hc108c1a1, 32'h41b164a6} /* (20, 29, 7) {real, imag} */,
  {32'h41a60446, 32'h410d2608} /* (20, 29, 6) {real, imag} */,
  {32'hc1eee0e6, 32'h416ad374} /* (20, 29, 5) {real, imag} */,
  {32'hc2012ba2, 32'hc28c25a4} /* (20, 29, 4) {real, imag} */,
  {32'h420c9093, 32'h41dba062} /* (20, 29, 3) {real, imag} */,
  {32'hc230436e, 32'hc134fe0d} /* (20, 29, 2) {real, imag} */,
  {32'h42a0e563, 32'h41cef548} /* (20, 29, 1) {real, imag} */,
  {32'h42209e94, 32'hbf307e78} /* (20, 29, 0) {real, imag} */,
  {32'h42214158, 32'hbf2e5918} /* (20, 28, 31) {real, imag} */,
  {32'h40bd6522, 32'hc26bc412} /* (20, 28, 30) {real, imag} */,
  {32'h4229634e, 32'hc1c0f310} /* (20, 28, 29) {real, imag} */,
  {32'hc1c941e8, 32'h41368c40} /* (20, 28, 28) {real, imag} */,
  {32'hc176bf74, 32'hc28acbb7} /* (20, 28, 27) {real, imag} */,
  {32'h418ca34f, 32'h41b11b90} /* (20, 28, 26) {real, imag} */,
  {32'hbff15a40, 32'h41b20e56} /* (20, 28, 25) {real, imag} */,
  {32'h424c3427, 32'hc1431b94} /* (20, 28, 24) {real, imag} */,
  {32'h41909512, 32'h4189028a} /* (20, 28, 23) {real, imag} */,
  {32'h419709ec, 32'hc160395e} /* (20, 28, 22) {real, imag} */,
  {32'h40c4daa4, 32'hc20aa82b} /* (20, 28, 21) {real, imag} */,
  {32'h3f5f2c60, 32'hc0964cb4} /* (20, 28, 20) {real, imag} */,
  {32'h3e18b540, 32'h40584ab4} /* (20, 28, 19) {real, imag} */,
  {32'h3f6c46c0, 32'hc00cdca0} /* (20, 28, 18) {real, imag} */,
  {32'h4019012a, 32'h4181d299} /* (20, 28, 17) {real, imag} */,
  {32'h3fb5c180, 32'h40d51cf8} /* (20, 28, 16) {real, imag} */,
  {32'hbd556880, 32'hbf7887a8} /* (20, 28, 15) {real, imag} */,
  {32'hc072f778, 32'h41f502a0} /* (20, 28, 14) {real, imag} */,
  {32'hc19db474, 32'hc10a5643} /* (20, 28, 13) {real, imag} */,
  {32'hc1ca9093, 32'hc142deea} /* (20, 28, 12) {real, imag} */,
  {32'h4219e7ae, 32'h40730d04} /* (20, 28, 11) {real, imag} */,
  {32'hc15692bc, 32'hc15e2ca0} /* (20, 28, 10) {real, imag} */,
  {32'h4206c0aa, 32'h411e2e43} /* (20, 28, 9) {real, imag} */,
  {32'h414db74c, 32'hc167650e} /* (20, 28, 8) {real, imag} */,
  {32'hc151e9d4, 32'hc0587f34} /* (20, 28, 7) {real, imag} */,
  {32'h41715a7e, 32'h4129aa11} /* (20, 28, 6) {real, imag} */,
  {32'h41efdf3c, 32'h418e8a0c} /* (20, 28, 5) {real, imag} */,
  {32'hc253e5dc, 32'hc2a14448} /* (20, 28, 4) {real, imag} */,
  {32'hc2873935, 32'hc22b9600} /* (20, 28, 3) {real, imag} */,
  {32'h419042de, 32'h4280179a} /* (20, 28, 2) {real, imag} */,
  {32'h40e90000, 32'h415b220a} /* (20, 28, 1) {real, imag} */,
  {32'hc279c51a, 32'h41fba41a} /* (20, 28, 0) {real, imag} */,
  {32'h420e17f6, 32'h42815510} /* (20, 27, 31) {real, imag} */,
  {32'hc2a26202, 32'h429ae8d3} /* (20, 27, 30) {real, imag} */,
  {32'hc14f0e77, 32'hc2a6abdb} /* (20, 27, 29) {real, imag} */,
  {32'hc15a62b2, 32'h4153a6c4} /* (20, 27, 28) {real, imag} */,
  {32'hc20b0521, 32'hc191010b} /* (20, 27, 27) {real, imag} */,
  {32'hc2b2b2dc, 32'h40e76c58} /* (20, 27, 26) {real, imag} */,
  {32'h42419fd8, 32'hc10e9b36} /* (20, 27, 25) {real, imag} */,
  {32'hc17fe42f, 32'hc21187ae} /* (20, 27, 24) {real, imag} */,
  {32'hc1422232, 32'hc1710537} /* (20, 27, 23) {real, imag} */,
  {32'h40dd90da, 32'h40260348} /* (20, 27, 22) {real, imag} */,
  {32'h41c5200a, 32'h40e0f3c5} /* (20, 27, 21) {real, imag} */,
  {32'h41c9f122, 32'hc185ec98} /* (20, 27, 20) {real, imag} */,
  {32'hc050f6bc, 32'h418e712a} /* (20, 27, 19) {real, imag} */,
  {32'h412ace6a, 32'h4148905c} /* (20, 27, 18) {real, imag} */,
  {32'hc15f7a22, 32'h41672171} /* (20, 27, 17) {real, imag} */,
  {32'h3fdaf0b8, 32'hc0721100} /* (20, 27, 16) {real, imag} */,
  {32'h4191a691, 32'hc104b59d} /* (20, 27, 15) {real, imag} */,
  {32'hbfcd1410, 32'h418855ee} /* (20, 27, 14) {real, imag} */,
  {32'h3fbc0b78, 32'h40ebd217} /* (20, 27, 13) {real, imag} */,
  {32'hc2077136, 32'h40bba444} /* (20, 27, 12) {real, imag} */,
  {32'hc165daa8, 32'h416023ea} /* (20, 27, 11) {real, imag} */,
  {32'h41b22fb8, 32'hc27d8888} /* (20, 27, 10) {real, imag} */,
  {32'hc2720b44, 32'hc1c33cce} /* (20, 27, 9) {real, imag} */,
  {32'hc089e0de, 32'h422e4d36} /* (20, 27, 8) {real, imag} */,
  {32'h40f7039c, 32'h421b9558} /* (20, 27, 7) {real, imag} */,
  {32'h42255d77, 32'hc1b86100} /* (20, 27, 6) {real, imag} */,
  {32'hc1c8daa0, 32'h418245e1} /* (20, 27, 5) {real, imag} */,
  {32'h41bd929d, 32'hc2351a83} /* (20, 27, 4) {real, imag} */,
  {32'h41121b15, 32'hc2a357ed} /* (20, 27, 3) {real, imag} */,
  {32'h42110c77, 32'hc1043060} /* (20, 27, 2) {real, imag} */,
  {32'h4239df72, 32'h425e4e63} /* (20, 27, 1) {real, imag} */,
  {32'hc1ac6c2c, 32'h41bdbc9a} /* (20, 27, 0) {real, imag} */,
  {32'hc22e0eca, 32'h422a172e} /* (20, 26, 31) {real, imag} */,
  {32'h421c511a, 32'hc226eb6c} /* (20, 26, 30) {real, imag} */,
  {32'h410e339c, 32'hc0bd9359} /* (20, 26, 29) {real, imag} */,
  {32'h413568cc, 32'h3fee76c0} /* (20, 26, 28) {real, imag} */,
  {32'hc280f6f0, 32'h4117dc60} /* (20, 26, 27) {real, imag} */,
  {32'h4220c28a, 32'h411ee3f0} /* (20, 26, 26) {real, imag} */,
  {32'hc21607ae, 32'hc1182cc6} /* (20, 26, 25) {real, imag} */,
  {32'h40f789cc, 32'hc185a4ed} /* (20, 26, 24) {real, imag} */,
  {32'h40fbbe28, 32'hc1412706} /* (20, 26, 23) {real, imag} */,
  {32'h41681896, 32'hc00a1f58} /* (20, 26, 22) {real, imag} */,
  {32'hc1d6225c, 32'h3ea74fa0} /* (20, 26, 21) {real, imag} */,
  {32'hc0b01d7d, 32'h40f0dc19} /* (20, 26, 20) {real, imag} */,
  {32'h410a029f, 32'hbfb6b5e4} /* (20, 26, 19) {real, imag} */,
  {32'h4088a311, 32'hc198e49a} /* (20, 26, 18) {real, imag} */,
  {32'h4042b678, 32'h3f68ade0} /* (20, 26, 17) {real, imag} */,
  {32'hc089dc34, 32'hc062eb08} /* (20, 26, 16) {real, imag} */,
  {32'hc13b0966, 32'hbf98bdd0} /* (20, 26, 15) {real, imag} */,
  {32'h40b75c67, 32'h40f8f8a8} /* (20, 26, 14) {real, imag} */,
  {32'h41050d29, 32'hc1677f9e} /* (20, 26, 13) {real, imag} */,
  {32'hc0ed0121, 32'h415b0fb8} /* (20, 26, 12) {real, imag} */,
  {32'h4110bdb8, 32'hc17759a6} /* (20, 26, 11) {real, imag} */,
  {32'h4188b800, 32'hbfd28620} /* (20, 26, 10) {real, imag} */,
  {32'h40fab388, 32'hc19b2e65} /* (20, 26, 9) {real, imag} */,
  {32'hc221bbf0, 32'h42025e08} /* (20, 26, 8) {real, imag} */,
  {32'h3f0cad60, 32'hc1dd9b29} /* (20, 26, 7) {real, imag} */,
  {32'h41ca7da4, 32'h423f8fca} /* (20, 26, 6) {real, imag} */,
  {32'h4195fbe0, 32'h41f02df8} /* (20, 26, 5) {real, imag} */,
  {32'hc18dd3dc, 32'h41a463f8} /* (20, 26, 4) {real, imag} */,
  {32'hc22f59e5, 32'h41178ad6} /* (20, 26, 3) {real, imag} */,
  {32'h41996a8a, 32'hc2242be8} /* (20, 26, 2) {real, imag} */,
  {32'h41da360c, 32'h425445b6} /* (20, 26, 1) {real, imag} */,
  {32'hc216b1d2, 32'hc2282da2} /* (20, 26, 0) {real, imag} */,
  {32'hc22ebef6, 32'hc21c4eca} /* (20, 25, 31) {real, imag} */,
  {32'hc224bed3, 32'hc2308b74} /* (20, 25, 30) {real, imag} */,
  {32'h41f9d726, 32'h420ec3ea} /* (20, 25, 29) {real, imag} */,
  {32'h40efc54e, 32'h4204ac6e} /* (20, 25, 28) {real, imag} */,
  {32'h4165b99c, 32'h405414c0} /* (20, 25, 27) {real, imag} */,
  {32'hc1da78b3, 32'hc164cfaf} /* (20, 25, 26) {real, imag} */,
  {32'hc17fbbbb, 32'h41875cd6} /* (20, 25, 25) {real, imag} */,
  {32'h41f708e6, 32'h40ed0f32} /* (20, 25, 24) {real, imag} */,
  {32'hc1820ddb, 32'h3ff7f739} /* (20, 25, 23) {real, imag} */,
  {32'hc16436e7, 32'hc13a7a9e} /* (20, 25, 22) {real, imag} */,
  {32'hc1a560ce, 32'hc01e3f40} /* (20, 25, 21) {real, imag} */,
  {32'h41bd04ac, 32'hc0c6f1e8} /* (20, 25, 20) {real, imag} */,
  {32'hbf917740, 32'h413c3252} /* (20, 25, 19) {real, imag} */,
  {32'h411e0a6f, 32'h4115470e} /* (20, 25, 18) {real, imag} */,
  {32'h40e3ef11, 32'hc10f2618} /* (20, 25, 17) {real, imag} */,
  {32'h414fdfad, 32'h41942e00} /* (20, 25, 16) {real, imag} */,
  {32'hc03e276e, 32'h410ca5dc} /* (20, 25, 15) {real, imag} */,
  {32'hc1ae0dc4, 32'h4013d638} /* (20, 25, 14) {real, imag} */,
  {32'h40b56904, 32'hbe5d1500} /* (20, 25, 13) {real, imag} */,
  {32'hc0c3d19a, 32'hc1263408} /* (20, 25, 12) {real, imag} */,
  {32'h40a64bae, 32'h418a7334} /* (20, 25, 11) {real, imag} */,
  {32'h40cb09a6, 32'h413a61fa} /* (20, 25, 10) {real, imag} */,
  {32'h4233a1f4, 32'hbfe66be9} /* (20, 25, 9) {real, imag} */,
  {32'hc1c1807e, 32'hc218e714} /* (20, 25, 8) {real, imag} */,
  {32'hc1a9d244, 32'h41d6ac42} /* (20, 25, 7) {real, imag} */,
  {32'hc20d357d, 32'h4135cf71} /* (20, 25, 6) {real, imag} */,
  {32'h41b8149a, 32'hc241e9ea} /* (20, 25, 5) {real, imag} */,
  {32'h41a4ac36, 32'hc1b6cb17} /* (20, 25, 4) {real, imag} */,
  {32'h41428a6b, 32'h41db7a2c} /* (20, 25, 3) {real, imag} */,
  {32'hc040b2d0, 32'h41640886} /* (20, 25, 2) {real, imag} */,
  {32'h41e1f404, 32'hc1985fcc} /* (20, 25, 1) {real, imag} */,
  {32'h42075487, 32'h4281af11} /* (20, 25, 0) {real, imag} */,
  {32'h402466a0, 32'h412f1978} /* (20, 24, 31) {real, imag} */,
  {32'h4272d849, 32'h421bf6fe} /* (20, 24, 30) {real, imag} */,
  {32'h423fd6ea, 32'hc1aca789} /* (20, 24, 29) {real, imag} */,
  {32'h422a7147, 32'h418b2fce} /* (20, 24, 28) {real, imag} */,
  {32'h412b632c, 32'hc1a8c4c2} /* (20, 24, 27) {real, imag} */,
  {32'h41e69a67, 32'hc0540888} /* (20, 24, 26) {real, imag} */,
  {32'h41dbd110, 32'hc141dd06} /* (20, 24, 25) {real, imag} */,
  {32'hc08d27be, 32'hc178dd95} /* (20, 24, 24) {real, imag} */,
  {32'hc1cf64e2, 32'h413adff0} /* (20, 24, 23) {real, imag} */,
  {32'hc12eb3c9, 32'h40983ae1} /* (20, 24, 22) {real, imag} */,
  {32'h40936dd2, 32'hbf447118} /* (20, 24, 21) {real, imag} */,
  {32'h4182febc, 32'h40c702b5} /* (20, 24, 20) {real, imag} */,
  {32'h40f3c764, 32'h407c1149} /* (20, 24, 19) {real, imag} */,
  {32'hc0cc9782, 32'hc13cce85} /* (20, 24, 18) {real, imag} */,
  {32'hbfeacf7e, 32'hc0d6ab82} /* (20, 24, 17) {real, imag} */,
  {32'hc0889239, 32'hc1444d9f} /* (20, 24, 16) {real, imag} */,
  {32'h40985358, 32'hc0a81376} /* (20, 24, 15) {real, imag} */,
  {32'h404e792c, 32'h4033dc94} /* (20, 24, 14) {real, imag} */,
  {32'hc0b0233c, 32'h400f67ff} /* (20, 24, 13) {real, imag} */,
  {32'h3fbe9a08, 32'hbf411b68} /* (20, 24, 12) {real, imag} */,
  {32'h3f82461a, 32'hbf626e38} /* (20, 24, 11) {real, imag} */,
  {32'hc1824fc0, 32'h407f482e} /* (20, 24, 10) {real, imag} */,
  {32'h3f6bbb70, 32'hc13173c0} /* (20, 24, 9) {real, imag} */,
  {32'hc0a5acc4, 32'hc1e19d64} /* (20, 24, 8) {real, imag} */,
  {32'h418411a2, 32'h409a69b4} /* (20, 24, 7) {real, imag} */,
  {32'h40c81c8c, 32'hc1c6ea6d} /* (20, 24, 6) {real, imag} */,
  {32'hc2014631, 32'hc07ac144} /* (20, 24, 5) {real, imag} */,
  {32'h41aaa77e, 32'hc158b364} /* (20, 24, 4) {real, imag} */,
  {32'hc1960543, 32'hc185df73} /* (20, 24, 3) {real, imag} */,
  {32'hc203b15f, 32'h42116f36} /* (20, 24, 2) {real, imag} */,
  {32'hc1744732, 32'hc2038520} /* (20, 24, 1) {real, imag} */,
  {32'h411412fa, 32'h3fa10db8} /* (20, 24, 0) {real, imag} */,
  {32'hc27032d6, 32'h41d14cea} /* (20, 23, 31) {real, imag} */,
  {32'hc106f09b, 32'h40debbb0} /* (20, 23, 30) {real, imag} */,
  {32'hc1a07ca7, 32'h4241984b} /* (20, 23, 29) {real, imag} */,
  {32'hc1b91335, 32'hc164f0b0} /* (20, 23, 28) {real, imag} */,
  {32'h42329ffe, 32'h41b15226} /* (20, 23, 27) {real, imag} */,
  {32'h41a5a5fe, 32'h40e2b95a} /* (20, 23, 26) {real, imag} */,
  {32'hc18740c1, 32'h40872f38} /* (20, 23, 25) {real, imag} */,
  {32'hc15fd592, 32'h4031beb8} /* (20, 23, 24) {real, imag} */,
  {32'hc139cff2, 32'h410397c1} /* (20, 23, 23) {real, imag} */,
  {32'hc18b6ec5, 32'hc1404f03} /* (20, 23, 22) {real, imag} */,
  {32'h40ad698c, 32'hc1af96fc} /* (20, 23, 21) {real, imag} */,
  {32'hc0fed9c4, 32'h40591abf} /* (20, 23, 20) {real, imag} */,
  {32'hc1378402, 32'hc0e2161c} /* (20, 23, 19) {real, imag} */,
  {32'hc0acbbc4, 32'hc15ff24d} /* (20, 23, 18) {real, imag} */,
  {32'hc09dea4b, 32'hc02da198} /* (20, 23, 17) {real, imag} */,
  {32'h3fe45a90, 32'hc0786a4c} /* (20, 23, 16) {real, imag} */,
  {32'h3f454218, 32'h4108203e} /* (20, 23, 15) {real, imag} */,
  {32'h3fac4bda, 32'h4010cbd4} /* (20, 23, 14) {real, imag} */,
  {32'h415c8446, 32'h40abf698} /* (20, 23, 13) {real, imag} */,
  {32'hc071bcb0, 32'h4101b488} /* (20, 23, 12) {real, imag} */,
  {32'hbf8fe8c0, 32'h3fffc408} /* (20, 23, 11) {real, imag} */,
  {32'hc05c84ce, 32'h404934f4} /* (20, 23, 10) {real, imag} */,
  {32'hc20bc180, 32'hc1886a4c} /* (20, 23, 9) {real, imag} */,
  {32'h41501556, 32'hc0fcfd58} /* (20, 23, 8) {real, imag} */,
  {32'hc0d73cfd, 32'h4201e97d} /* (20, 23, 7) {real, imag} */,
  {32'hc0155034, 32'hbfbb2778} /* (20, 23, 6) {real, imag} */,
  {32'hc002d600, 32'hc167b4b3} /* (20, 23, 5) {real, imag} */,
  {32'h3fcf32e0, 32'hc14322f0} /* (20, 23, 4) {real, imag} */,
  {32'h41472062, 32'hc1abda62} /* (20, 23, 3) {real, imag} */,
  {32'h3ffb895e, 32'hc28aa931} /* (20, 23, 2) {real, imag} */,
  {32'hc1b634fb, 32'hc19457e4} /* (20, 23, 1) {real, imag} */,
  {32'h40f5385c, 32'h41dd4998} /* (20, 23, 0) {real, imag} */,
  {32'hc191a8ba, 32'h420b2100} /* (20, 22, 31) {real, imag} */,
  {32'h41a5a12e, 32'hc1528338} /* (20, 22, 30) {real, imag} */,
  {32'hc21a9c43, 32'h416fa0f6} /* (20, 22, 29) {real, imag} */,
  {32'h41f14393, 32'h41166c9a} /* (20, 22, 28) {real, imag} */,
  {32'hc18e7218, 32'hc18b040e} /* (20, 22, 27) {real, imag} */,
  {32'hc22a6301, 32'h410bf51a} /* (20, 22, 26) {real, imag} */,
  {32'hc1145f90, 32'h4145e860} /* (20, 22, 25) {real, imag} */,
  {32'hc008d782, 32'h41146cc4} /* (20, 22, 24) {real, imag} */,
  {32'hc18783db, 32'h3f98dd24} /* (20, 22, 23) {real, imag} */,
  {32'hc02ed7c0, 32'hc07e39b6} /* (20, 22, 22) {real, imag} */,
  {32'hc060d666, 32'h3e759ea0} /* (20, 22, 21) {real, imag} */,
  {32'hc13965c2, 32'hc1765e49} /* (20, 22, 20) {real, imag} */,
  {32'hc0b55fba, 32'hbe4bbd00} /* (20, 22, 19) {real, imag} */,
  {32'h419ef5c4, 32'h40aceb1a} /* (20, 22, 18) {real, imag} */,
  {32'h413b1d7e, 32'hc140d8b9} /* (20, 22, 17) {real, imag} */,
  {32'hc0ac262b, 32'hbf32db28} /* (20, 22, 16) {real, imag} */,
  {32'hbfcd0480, 32'h3ca2aa00} /* (20, 22, 15) {real, imag} */,
  {32'hc11c0962, 32'h40ca9830} /* (20, 22, 14) {real, imag} */,
  {32'h41135e4d, 32'hc0cb605e} /* (20, 22, 13) {real, imag} */,
  {32'h404d9916, 32'h408314ee} /* (20, 22, 12) {real, imag} */,
  {32'h410bf6e2, 32'hbf0a06a8} /* (20, 22, 11) {real, imag} */,
  {32'h40c3aa6c, 32'h3fbb240c} /* (20, 22, 10) {real, imag} */,
  {32'h3fe7ded0, 32'h413b98ec} /* (20, 22, 9) {real, imag} */,
  {32'hc132e70e, 32'h418e60f1} /* (20, 22, 8) {real, imag} */,
  {32'h3fffde80, 32'h410e9424} /* (20, 22, 7) {real, imag} */,
  {32'hc1c497aa, 32'h401b359a} /* (20, 22, 6) {real, imag} */,
  {32'hc1018bcc, 32'hc23517fb} /* (20, 22, 5) {real, imag} */,
  {32'h40eb5c14, 32'h40bd88bd} /* (20, 22, 4) {real, imag} */,
  {32'hc09c46b8, 32'h417d4672} /* (20, 22, 3) {real, imag} */,
  {32'hc0bfa26c, 32'hc137ba58} /* (20, 22, 2) {real, imag} */,
  {32'hc1e53ee2, 32'hc0b135e4} /* (20, 22, 1) {real, imag} */,
  {32'hc11d75f2, 32'h410646a4} /* (20, 22, 0) {real, imag} */,
  {32'hc02a29b8, 32'h410edc41} /* (20, 21, 31) {real, imag} */,
  {32'h41e94bfb, 32'hc194b878} /* (20, 21, 30) {real, imag} */,
  {32'h420704c0, 32'hc193240c} /* (20, 21, 29) {real, imag} */,
  {32'h3fc7bf28, 32'h411f73ca} /* (20, 21, 28) {real, imag} */,
  {32'h409c1d24, 32'hc13843f3} /* (20, 21, 27) {real, imag} */,
  {32'hc204c18e, 32'hbf8f3c74} /* (20, 21, 26) {real, imag} */,
  {32'hc1879d9a, 32'hc15bfce9} /* (20, 21, 25) {real, imag} */,
  {32'h41913d31, 32'hc1282234} /* (20, 21, 24) {real, imag} */,
  {32'h41eaa445, 32'hc1d280e2} /* (20, 21, 23) {real, imag} */,
  {32'hc17b726e, 32'h407bc8f3} /* (20, 21, 22) {real, imag} */,
  {32'h403b2d98, 32'hc0aaffa7} /* (20, 21, 21) {real, imag} */,
  {32'h412c88d3, 32'h402626a2} /* (20, 21, 20) {real, imag} */,
  {32'hc0aca3a0, 32'h3f70f618} /* (20, 21, 19) {real, imag} */,
  {32'h40927680, 32'hc0a3a236} /* (20, 21, 18) {real, imag} */,
  {32'hc03ce3c8, 32'h40de5ed9} /* (20, 21, 17) {real, imag} */,
  {32'h3f735d58, 32'hc09de0ea} /* (20, 21, 16) {real, imag} */,
  {32'hbf211cc0, 32'h404e9432} /* (20, 21, 15) {real, imag} */,
  {32'h40b2af60, 32'h3fbf6286} /* (20, 21, 14) {real, imag} */,
  {32'hbf641d60, 32'hc143aaee} /* (20, 21, 13) {real, imag} */,
  {32'h416f2ac7, 32'hc13837b0} /* (20, 21, 12) {real, imag} */,
  {32'h4125a146, 32'h412168a6} /* (20, 21, 11) {real, imag} */,
  {32'h418574e5, 32'hc0c4aa36} /* (20, 21, 10) {real, imag} */,
  {32'hc0cb4fec, 32'hc0402e0c} /* (20, 21, 9) {real, imag} */,
  {32'h40843304, 32'h418b62ef} /* (20, 21, 8) {real, imag} */,
  {32'h4204848b, 32'h4027242c} /* (20, 21, 7) {real, imag} */,
  {32'h410ea860, 32'h3fcbccd0} /* (20, 21, 6) {real, imag} */,
  {32'h40ad7d5c, 32'hc180b84e} /* (20, 21, 5) {real, imag} */,
  {32'hc1a363e2, 32'hc0b1bfe7} /* (20, 21, 4) {real, imag} */,
  {32'h419b6768, 32'h41334f3c} /* (20, 21, 3) {real, imag} */,
  {32'hc200b2a6, 32'h4168972d} /* (20, 21, 2) {real, imag} */,
  {32'h40d49e78, 32'h41d62fea} /* (20, 21, 1) {real, imag} */,
  {32'hc0d907a1, 32'h420ba483} /* (20, 21, 0) {real, imag} */,
  {32'hc0fb4bbb, 32'h41216ef7} /* (20, 20, 31) {real, imag} */,
  {32'hc086239a, 32'h4196737e} /* (20, 20, 30) {real, imag} */,
  {32'h41f80373, 32'hc1c3d520} /* (20, 20, 29) {real, imag} */,
  {32'hc0dae6a5, 32'h40378756} /* (20, 20, 28) {real, imag} */,
  {32'h4194e234, 32'h41355264} /* (20, 20, 27) {real, imag} */,
  {32'hc041c6ae, 32'h41f87afe} /* (20, 20, 26) {real, imag} */,
  {32'hc0494dbc, 32'hc06f3602} /* (20, 20, 25) {real, imag} */,
  {32'hc0c0d11c, 32'hbfa798d4} /* (20, 20, 24) {real, imag} */,
  {32'h41d65059, 32'h417d7f44} /* (20, 20, 23) {real, imag} */,
  {32'hc126921a, 32'hc17ff454} /* (20, 20, 22) {real, imag} */,
  {32'hbec26fd8, 32'h40f02378} /* (20, 20, 21) {real, imag} */,
  {32'hc14c25e3, 32'h40a95589} /* (20, 20, 20) {real, imag} */,
  {32'hc0ec3612, 32'h3ee831f8} /* (20, 20, 19) {real, imag} */,
  {32'hc0b2b718, 32'h40c10b81} /* (20, 20, 18) {real, imag} */,
  {32'h405d53d8, 32'h4064679c} /* (20, 20, 17) {real, imag} */,
  {32'h40db0d64, 32'hc04c3330} /* (20, 20, 16) {real, imag} */,
  {32'hc07f106c, 32'h3f0708f0} /* (20, 20, 15) {real, imag} */,
  {32'hc0f403d4, 32'hbfd070f4} /* (20, 20, 14) {real, imag} */,
  {32'hc08cb60e, 32'h40cbf284} /* (20, 20, 13) {real, imag} */,
  {32'h3f978280, 32'hc0c43777} /* (20, 20, 12) {real, imag} */,
  {32'h3db311a0, 32'hbdf0b8e0} /* (20, 20, 11) {real, imag} */,
  {32'h40ce2f8b, 32'h4114e336} /* (20, 20, 10) {real, imag} */,
  {32'hc105f4aa, 32'h4117ca08} /* (20, 20, 9) {real, imag} */,
  {32'h40a0e3e0, 32'h411b3b90} /* (20, 20, 8) {real, imag} */,
  {32'hc019458c, 32'h41572e54} /* (20, 20, 7) {real, imag} */,
  {32'h408293a1, 32'h4155ae55} /* (20, 20, 6) {real, imag} */,
  {32'hc0ac0c2e, 32'h41217b64} /* (20, 20, 5) {real, imag} */,
  {32'hc1a94045, 32'hc0f8df4d} /* (20, 20, 4) {real, imag} */,
  {32'h41aa0659, 32'hc1aa9620} /* (20, 20, 3) {real, imag} */,
  {32'h402bf773, 32'h4120fe22} /* (20, 20, 2) {real, imag} */,
  {32'hc1574306, 32'hc1b80d84} /* (20, 20, 1) {real, imag} */,
  {32'h41ea46bf, 32'hc23afaa9} /* (20, 20, 0) {real, imag} */,
  {32'hc139e6ee, 32'hc1b1a902} /* (20, 19, 31) {real, imag} */,
  {32'hc089be04, 32'h40b0506d} /* (20, 19, 30) {real, imag} */,
  {32'h402b13e4, 32'h4190bc7d} /* (20, 19, 29) {real, imag} */,
  {32'hc12d49a9, 32'h41d45765} /* (20, 19, 28) {real, imag} */,
  {32'h4216a146, 32'h409693a0} /* (20, 19, 27) {real, imag} */,
  {32'h3ff6b72e, 32'hc016cf08} /* (20, 19, 26) {real, imag} */,
  {32'h4110e149, 32'h40cfda0c} /* (20, 19, 25) {real, imag} */,
  {32'h413f720c, 32'h3ec05e78} /* (20, 19, 24) {real, imag} */,
  {32'h413f1640, 32'hbf4e4d66} /* (20, 19, 23) {real, imag} */,
  {32'h40290712, 32'h40dab8f5} /* (20, 19, 22) {real, imag} */,
  {32'h4110f1cd, 32'hc0eb4d13} /* (20, 19, 21) {real, imag} */,
  {32'hbf4786a8, 32'h40a8ab70} /* (20, 19, 20) {real, imag} */,
  {32'hbf22e850, 32'hbf7e1a08} /* (20, 19, 19) {real, imag} */,
  {32'hc015064c, 32'h3f5e8004} /* (20, 19, 18) {real, imag} */,
  {32'hc02cfc66, 32'hc030a53c} /* (20, 19, 17) {real, imag} */,
  {32'hc0cec988, 32'hbfa7f470} /* (20, 19, 16) {real, imag} */,
  {32'hc020f1a2, 32'h404b6efc} /* (20, 19, 15) {real, imag} */,
  {32'hc0c02a7a, 32'hc0b78334} /* (20, 19, 14) {real, imag} */,
  {32'hc0936b26, 32'hc0246dba} /* (20, 19, 13) {real, imag} */,
  {32'hbf901140, 32'hc1158dba} /* (20, 19, 12) {real, imag} */,
  {32'h41502447, 32'hbf627518} /* (20, 19, 11) {real, imag} */,
  {32'h3f6b3010, 32'hbfc294ec} /* (20, 19, 10) {real, imag} */,
  {32'h40d3e8d5, 32'h4088deec} /* (20, 19, 9) {real, imag} */,
  {32'h410b329c, 32'hbed43548} /* (20, 19, 8) {real, imag} */,
  {32'h3fcb2828, 32'hc03f5e78} /* (20, 19, 7) {real, imag} */,
  {32'hc10864e4, 32'hc1b135ff} /* (20, 19, 6) {real, imag} */,
  {32'hc195b5d3, 32'hc1b2fd36} /* (20, 19, 5) {real, imag} */,
  {32'hc0d1dc3e, 32'h3fb36e00} /* (20, 19, 4) {real, imag} */,
  {32'hc1db71f4, 32'hc1e05ec7} /* (20, 19, 3) {real, imag} */,
  {32'h4181ce87, 32'hc0fc9437} /* (20, 19, 2) {real, imag} */,
  {32'hc1d5343d, 32'h40cd8f66} /* (20, 19, 1) {real, imag} */,
  {32'h41b03ace, 32'hc0022cee} /* (20, 19, 0) {real, imag} */,
  {32'h406bc838, 32'h4021daf8} /* (20, 18, 31) {real, imag} */,
  {32'h4140ed78, 32'h410ed85c} /* (20, 18, 30) {real, imag} */,
  {32'hc14a23aa, 32'h3f3bbedc} /* (20, 18, 29) {real, imag} */,
  {32'hc19f6fd0, 32'hc16a7e5f} /* (20, 18, 28) {real, imag} */,
  {32'hc10ce8dd, 32'h42094244} /* (20, 18, 27) {real, imag} */,
  {32'hc0e489ce, 32'h415bc78a} /* (20, 18, 26) {real, imag} */,
  {32'hc1c277dc, 32'h3f2b3f3c} /* (20, 18, 25) {real, imag} */,
  {32'h40910df6, 32'hbf2485f6} /* (20, 18, 24) {real, imag} */,
  {32'hc13df208, 32'hc0cea4a6} /* (20, 18, 23) {real, imag} */,
  {32'hc0760eec, 32'hc088740b} /* (20, 18, 22) {real, imag} */,
  {32'h40950514, 32'hc074ef44} /* (20, 18, 21) {real, imag} */,
  {32'h3f272dac, 32'hc04ed4d8} /* (20, 18, 20) {real, imag} */,
  {32'h408cf067, 32'hc08e428e} /* (20, 18, 19) {real, imag} */,
  {32'h406e5c62, 32'h410318f3} /* (20, 18, 18) {real, imag} */,
  {32'h411aa41a, 32'h40cd39f2} /* (20, 18, 17) {real, imag} */,
  {32'hbfa05722, 32'h40a02f22} /* (20, 18, 16) {real, imag} */,
  {32'hbfbb31cc, 32'hbfe79b9e} /* (20, 18, 15) {real, imag} */,
  {32'h3f1095e8, 32'hbeca6ce0} /* (20, 18, 14) {real, imag} */,
  {32'h40b37bd5, 32'h409af46a} /* (20, 18, 13) {real, imag} */,
  {32'h40e57e86, 32'h4035d5b8} /* (20, 18, 12) {real, imag} */,
  {32'h412f589e, 32'h40c0d286} /* (20, 18, 11) {real, imag} */,
  {32'hc1773355, 32'hbf0e94a8} /* (20, 18, 10) {real, imag} */,
  {32'hc12cded6, 32'hc08d6b78} /* (20, 18, 9) {real, imag} */,
  {32'hbf76663e, 32'hc0813107} /* (20, 18, 8) {real, imag} */,
  {32'hc0f0bd42, 32'hc00b244b} /* (20, 18, 7) {real, imag} */,
  {32'hc1a17106, 32'hc100ceaa} /* (20, 18, 6) {real, imag} */,
  {32'h3f2dec10, 32'h416b322a} /* (20, 18, 5) {real, imag} */,
  {32'h41caed7a, 32'h3ede9060} /* (20, 18, 4) {real, imag} */,
  {32'h4029d2ae, 32'hc0164385} /* (20, 18, 3) {real, imag} */,
  {32'hc15892da, 32'hc159f916} /* (20, 18, 2) {real, imag} */,
  {32'hc16be35a, 32'h411c3f66} /* (20, 18, 1) {real, imag} */,
  {32'hc01e86bc, 32'hc12751c8} /* (20, 18, 0) {real, imag} */,
  {32'h4026438c, 32'hc0f5a4bb} /* (20, 17, 31) {real, imag} */,
  {32'h3f8032be, 32'hc026d445} /* (20, 17, 30) {real, imag} */,
  {32'hc0d0c5f8, 32'hbf0aa09e} /* (20, 17, 29) {real, imag} */,
  {32'hc17722c9, 32'h418c301a} /* (20, 17, 28) {real, imag} */,
  {32'hc0e9bf5a, 32'hc1324799} /* (20, 17, 27) {real, imag} */,
  {32'h3ffcc148, 32'h41a95370} /* (20, 17, 26) {real, imag} */,
  {32'h3fdd8a9c, 32'hc105024e} /* (20, 17, 25) {real, imag} */,
  {32'h404705aa, 32'h41485852} /* (20, 17, 24) {real, imag} */,
  {32'hbf3143b0, 32'hc023f2bc} /* (20, 17, 23) {real, imag} */,
  {32'hc1129ab0, 32'h3f60f0c2} /* (20, 17, 22) {real, imag} */,
  {32'h3fe6c938, 32'hc0de610d} /* (20, 17, 21) {real, imag} */,
  {32'h4015a60c, 32'h4123f276} /* (20, 17, 20) {real, imag} */,
  {32'h40bde2b6, 32'h408798bd} /* (20, 17, 19) {real, imag} */,
  {32'hbfa09466, 32'hbf42ccb4} /* (20, 17, 18) {real, imag} */,
  {32'hbf87583c, 32'h4023ec44} /* (20, 17, 17) {real, imag} */,
  {32'hbee378f0, 32'hbfde9b48} /* (20, 17, 16) {real, imag} */,
  {32'h40655b7a, 32'hc0bb8752} /* (20, 17, 15) {real, imag} */,
  {32'h40182d1b, 32'h3fec4f82} /* (20, 17, 14) {real, imag} */,
  {32'h3f73bbc0, 32'hbf3c8618} /* (20, 17, 13) {real, imag} */,
  {32'hc16c3e57, 32'hbf97752c} /* (20, 17, 12) {real, imag} */,
  {32'hc0adcbee, 32'hc05c70d2} /* (20, 17, 11) {real, imag} */,
  {32'h3ec66570, 32'h40365d30} /* (20, 17, 10) {real, imag} */,
  {32'h418ab7ae, 32'h3f5d3be8} /* (20, 17, 9) {real, imag} */,
  {32'h41439faa, 32'hc09c41e8} /* (20, 17, 8) {real, imag} */,
  {32'hc09f7b93, 32'hc0e3e544} /* (20, 17, 7) {real, imag} */,
  {32'hc08b48fa, 32'hc1388211} /* (20, 17, 6) {real, imag} */,
  {32'hc0c3f34e, 32'hc04747a0} /* (20, 17, 5) {real, imag} */,
  {32'h40e882ea, 32'hc03218b6} /* (20, 17, 4) {real, imag} */,
  {32'h41467e48, 32'h4034a0c0} /* (20, 17, 3) {real, imag} */,
  {32'h40e800a4, 32'hc1107f54} /* (20, 17, 2) {real, imag} */,
  {32'h41174200, 32'h40c9a78d} /* (20, 17, 1) {real, imag} */,
  {32'h4183044d, 32'hbeb41620} /* (20, 17, 0) {real, imag} */,
  {32'h40cbe33a, 32'h3e9f1770} /* (20, 16, 31) {real, imag} */,
  {32'hc02720cc, 32'hc0e3aafc} /* (20, 16, 30) {real, imag} */,
  {32'hc17cfb4d, 32'h403af46a} /* (20, 16, 29) {real, imag} */,
  {32'hbe74f780, 32'hc11ef7f5} /* (20, 16, 28) {real, imag} */,
  {32'h3dacb6e0, 32'hc0e321ed} /* (20, 16, 27) {real, imag} */,
  {32'hc17b1cc5, 32'h4121137c} /* (20, 16, 26) {real, imag} */,
  {32'h400328c6, 32'h412e6f63} /* (20, 16, 25) {real, imag} */,
  {32'hbf8cd5b8, 32'h411e23a0} /* (20, 16, 24) {real, imag} */,
  {32'h40df778a, 32'hc10c40dd} /* (20, 16, 23) {real, imag} */,
  {32'hc07d8e1e, 32'hbfd07cda} /* (20, 16, 22) {real, imag} */,
  {32'h3f1ce440, 32'hbd6e5120} /* (20, 16, 21) {real, imag} */,
  {32'hc0a72e31, 32'h3fdb3ccf} /* (20, 16, 20) {real, imag} */,
  {32'hc0d0f7d6, 32'hc0a0b47f} /* (20, 16, 19) {real, imag} */,
  {32'hc059288d, 32'hbfcd9280} /* (20, 16, 18) {real, imag} */,
  {32'hc070e13f, 32'hc0914b38} /* (20, 16, 17) {real, imag} */,
  {32'hc053f5fb, 32'hbedfb3dc} /* (20, 16, 16) {real, imag} */,
  {32'h40089025, 32'hc07d4e58} /* (20, 16, 15) {real, imag} */,
  {32'h3fe743c6, 32'h3fe0cdf0} /* (20, 16, 14) {real, imag} */,
  {32'hc0e90788, 32'hc0c34cab} /* (20, 16, 13) {real, imag} */,
  {32'h40f91ba7, 32'h3e5c7178} /* (20, 16, 12) {real, imag} */,
  {32'h410d164e, 32'h403717f0} /* (20, 16, 11) {real, imag} */,
  {32'hbf4a9f18, 32'h40ab3862} /* (20, 16, 10) {real, imag} */,
  {32'h4096c746, 32'hbfdf010a} /* (20, 16, 9) {real, imag} */,
  {32'hc11c97b7, 32'h40ace780} /* (20, 16, 8) {real, imag} */,
  {32'h4054a818, 32'hc0b24df2} /* (20, 16, 7) {real, imag} */,
  {32'hc0840686, 32'h40de0f44} /* (20, 16, 6) {real, imag} */,
  {32'h3fbfabae, 32'hc18315a3} /* (20, 16, 5) {real, imag} */,
  {32'hc18d5939, 32'h40e0fcbe} /* (20, 16, 4) {real, imag} */,
  {32'hc12049ff, 32'hc13ab6b4} /* (20, 16, 3) {real, imag} */,
  {32'h41918076, 32'hc1b1e0c8} /* (20, 16, 2) {real, imag} */,
  {32'h40d41f96, 32'h4173378c} /* (20, 16, 1) {real, imag} */,
  {32'h40aceeae, 32'h3fee944b} /* (20, 16, 0) {real, imag} */,
  {32'hc0c078f0, 32'h41dab440} /* (20, 15, 31) {real, imag} */,
  {32'h409cdcfe, 32'hc09b00c5} /* (20, 15, 30) {real, imag} */,
  {32'h4116ebfd, 32'h41015206} /* (20, 15, 29) {real, imag} */,
  {32'hc0524536, 32'hbdd1df00} /* (20, 15, 28) {real, imag} */,
  {32'hc1223afa, 32'hc17d8036} /* (20, 15, 27) {real, imag} */,
  {32'h41fe9ef9, 32'h40d92ba7} /* (20, 15, 26) {real, imag} */,
  {32'h415a8524, 32'h404fbefe} /* (20, 15, 25) {real, imag} */,
  {32'h3dc50a80, 32'h418a3661} /* (20, 15, 24) {real, imag} */,
  {32'hc0a83079, 32'hc122e65b} /* (20, 15, 23) {real, imag} */,
  {32'hc06bfdb2, 32'hc03a4d26} /* (20, 15, 22) {real, imag} */,
  {32'hc0045712, 32'hc003d67e} /* (20, 15, 21) {real, imag} */,
  {32'hbf03e524, 32'hc00a23e2} /* (20, 15, 20) {real, imag} */,
  {32'hc00c12c6, 32'hc0430bb8} /* (20, 15, 19) {real, imag} */,
  {32'h40c941ba, 32'hc02f32c2} /* (20, 15, 18) {real, imag} */,
  {32'h4047b71d, 32'h3fed0f38} /* (20, 15, 17) {real, imag} */,
  {32'hbebe0630, 32'hbe2924c0} /* (20, 15, 16) {real, imag} */,
  {32'hbea94280, 32'h3f3cbe30} /* (20, 15, 15) {real, imag} */,
  {32'hbf8cc5a6, 32'hbfb5508c} /* (20, 15, 14) {real, imag} */,
  {32'h401ae5fe, 32'hbf7fb7f2} /* (20, 15, 13) {real, imag} */,
  {32'h405bc753, 32'hc033c78e} /* (20, 15, 12) {real, imag} */,
  {32'h401f7d72, 32'h4067c192} /* (20, 15, 11) {real, imag} */,
  {32'h410cbb1a, 32'hc1209896} /* (20, 15, 10) {real, imag} */,
  {32'hc15dacec, 32'h41192bcd} /* (20, 15, 9) {real, imag} */,
  {32'hc0353934, 32'hc0560e1a} /* (20, 15, 8) {real, imag} */,
  {32'hc11a6580, 32'h41509138} /* (20, 15, 7) {real, imag} */,
  {32'h3f909230, 32'hc1ad1704} /* (20, 15, 6) {real, imag} */,
  {32'h40851e0f, 32'hc08eab44} /* (20, 15, 5) {real, imag} */,
  {32'h413b0ba4, 32'hc1b7cdbb} /* (20, 15, 4) {real, imag} */,
  {32'hc11cc9e7, 32'h3fada294} /* (20, 15, 3) {real, imag} */,
  {32'h41a2273c, 32'h409c090b} /* (20, 15, 2) {real, imag} */,
  {32'hbf7a1cf0, 32'h4043f46c} /* (20, 15, 1) {real, imag} */,
  {32'hc0328d56, 32'h4182c33c} /* (20, 15, 0) {real, imag} */,
  {32'h41974a42, 32'h3fb2c6f4} /* (20, 14, 31) {real, imag} */,
  {32'hc103b7fe, 32'hc1cfad36} /* (20, 14, 30) {real, imag} */,
  {32'hc0f58e42, 32'hc0b21a10} /* (20, 14, 29) {real, imag} */,
  {32'h3f666bc4, 32'h41668f84} /* (20, 14, 28) {real, imag} */,
  {32'h40f81fac, 32'hc1069888} /* (20, 14, 27) {real, imag} */,
  {32'hc0379509, 32'h41c7083a} /* (20, 14, 26) {real, imag} */,
  {32'h40e76672, 32'hc06dea72} /* (20, 14, 25) {real, imag} */,
  {32'hc03ef36d, 32'h40d0be37} /* (20, 14, 24) {real, imag} */,
  {32'h41780dc0, 32'h405f7101} /* (20, 14, 23) {real, imag} */,
  {32'h4135e014, 32'hc15174e6} /* (20, 14, 22) {real, imag} */,
  {32'hc0f0fc12, 32'h40a81298} /* (20, 14, 21) {real, imag} */,
  {32'hc105c04b, 32'hbfaebf67} /* (20, 14, 20) {real, imag} */,
  {32'h40cb8df6, 32'hc0e9d0f0} /* (20, 14, 19) {real, imag} */,
  {32'hbfe9e250, 32'h4118555c} /* (20, 14, 18) {real, imag} */,
  {32'hc0d4d876, 32'h400278ec} /* (20, 14, 17) {real, imag} */,
  {32'hc0b92418, 32'h3f8da028} /* (20, 14, 16) {real, imag} */,
  {32'hbe948658, 32'h40369d58} /* (20, 14, 15) {real, imag} */,
  {32'hc0693ed0, 32'h41155c32} /* (20, 14, 14) {real, imag} */,
  {32'h3fbcd8ba, 32'hc09f0874} /* (20, 14, 13) {real, imag} */,
  {32'hc0a3e476, 32'h3f4d465e} /* (20, 14, 12) {real, imag} */,
  {32'h40ca028e, 32'hc0ca765a} /* (20, 14, 11) {real, imag} */,
  {32'hc155f348, 32'h41209e1c} /* (20, 14, 10) {real, imag} */,
  {32'h40312828, 32'hc12b0986} /* (20, 14, 9) {real, imag} */,
  {32'hbf8638ba, 32'h402814aa} /* (20, 14, 8) {real, imag} */,
  {32'h40afdcca, 32'h400874b0} /* (20, 14, 7) {real, imag} */,
  {32'h3ebd1638, 32'hc000e68c} /* (20, 14, 6) {real, imag} */,
  {32'hc0beabd0, 32'hc14859d4} /* (20, 14, 5) {real, imag} */,
  {32'h4101f86a, 32'h410dc740} /* (20, 14, 4) {real, imag} */,
  {32'h41cf95c4, 32'h4119a6de} /* (20, 14, 3) {real, imag} */,
  {32'hc1486bd4, 32'h3db75180} /* (20, 14, 2) {real, imag} */,
  {32'h40bdb12e, 32'hc1096808} /* (20, 14, 1) {real, imag} */,
  {32'h4125a86c, 32'hc18b173e} /* (20, 14, 0) {real, imag} */,
  {32'h41591e36, 32'hc19f5314} /* (20, 13, 31) {real, imag} */,
  {32'h41c3da38, 32'hc17687bb} /* (20, 13, 30) {real, imag} */,
  {32'hbea13640, 32'h418f51d2} /* (20, 13, 29) {real, imag} */,
  {32'h4087f13c, 32'h40494bfc} /* (20, 13, 28) {real, imag} */,
  {32'hc107de0c, 32'h41431999} /* (20, 13, 27) {real, imag} */,
  {32'hc178f4b4, 32'h41a8fd5e} /* (20, 13, 26) {real, imag} */,
  {32'hc0161cd2, 32'h40114780} /* (20, 13, 25) {real, imag} */,
  {32'hc1601d0a, 32'hc19599ca} /* (20, 13, 24) {real, imag} */,
  {32'hc0af24d4, 32'hbf617b40} /* (20, 13, 23) {real, imag} */,
  {32'hbe8b1080, 32'hbfdc9128} /* (20, 13, 22) {real, imag} */,
  {32'hc0ba4cd2, 32'h400fe32c} /* (20, 13, 21) {real, imag} */,
  {32'h411f5390, 32'hc05e9ad4} /* (20, 13, 20) {real, imag} */,
  {32'h40873378, 32'h3ea42f30} /* (20, 13, 19) {real, imag} */,
  {32'h4000146c, 32'hc055d09f} /* (20, 13, 18) {real, imag} */,
  {32'hc06d628e, 32'h3f98831e} /* (20, 13, 17) {real, imag} */,
  {32'hc013582e, 32'h3f9e57c8} /* (20, 13, 16) {real, imag} */,
  {32'h408b8e5d, 32'h3f21270c} /* (20, 13, 15) {real, imag} */,
  {32'h401eb748, 32'hbff4e0a2} /* (20, 13, 14) {real, imag} */,
  {32'h3df06500, 32'hc0d62e97} /* (20, 13, 13) {real, imag} */,
  {32'h3ff7d380, 32'h407d05ac} /* (20, 13, 12) {real, imag} */,
  {32'h3f3b9a34, 32'hc0e0bbf2} /* (20, 13, 11) {real, imag} */,
  {32'h41a9986a, 32'h41737b6d} /* (20, 13, 10) {real, imag} */,
  {32'hc16fa3ca, 32'hbe3efaa0} /* (20, 13, 9) {real, imag} */,
  {32'hc0607e0e, 32'h3dde2780} /* (20, 13, 8) {real, imag} */,
  {32'hc08e2fb1, 32'h412a766c} /* (20, 13, 7) {real, imag} */,
  {32'h4103fe2c, 32'h41fd1f16} /* (20, 13, 6) {real, imag} */,
  {32'h3ebb2f30, 32'hc1ecd3f4} /* (20, 13, 5) {real, imag} */,
  {32'h417b3f82, 32'hc1c6258e} /* (20, 13, 4) {real, imag} */,
  {32'h41654690, 32'h418d261e} /* (20, 13, 3) {real, imag} */,
  {32'hc039f7a0, 32'hc1b2e285} /* (20, 13, 2) {real, imag} */,
  {32'h40b4d36c, 32'h409ad268} /* (20, 13, 1) {real, imag} */,
  {32'hbfa227f4, 32'h41deb92a} /* (20, 13, 0) {real, imag} */,
  {32'h41a2e12e, 32'h412f0b79} /* (20, 12, 31) {real, imag} */,
  {32'h40881d74, 32'hc053d560} /* (20, 12, 30) {real, imag} */,
  {32'h41884cb3, 32'hc1144614} /* (20, 12, 29) {real, imag} */,
  {32'h41400862, 32'hc1e2dd6e} /* (20, 12, 28) {real, imag} */,
  {32'hc2345176, 32'hbfbc6354} /* (20, 12, 27) {real, imag} */,
  {32'hc0cab6e4, 32'hbfe90800} /* (20, 12, 26) {real, imag} */,
  {32'h4112cf0e, 32'hc1bbdcd6} /* (20, 12, 25) {real, imag} */,
  {32'hc0e44b30, 32'h4185ee32} /* (20, 12, 24) {real, imag} */,
  {32'hc16bc602, 32'h3ff5bd94} /* (20, 12, 23) {real, imag} */,
  {32'hc0dee22c, 32'h41fce9de} /* (20, 12, 22) {real, imag} */,
  {32'h4123613a, 32'hbec55ae0} /* (20, 12, 21) {real, imag} */,
  {32'h4017a438, 32'hc18747ac} /* (20, 12, 20) {real, imag} */,
  {32'h40c0c23e, 32'hbfc9b8ac} /* (20, 12, 19) {real, imag} */,
  {32'h3e812e28, 32'hc09334a8} /* (20, 12, 18) {real, imag} */,
  {32'hc0607b8e, 32'h3fef1afc} /* (20, 12, 17) {real, imag} */,
  {32'hc00a4e8a, 32'hbf873248} /* (20, 12, 16) {real, imag} */,
  {32'h406f5956, 32'hc0b1adaf} /* (20, 12, 15) {real, imag} */,
  {32'hc09fa490, 32'hc09ec4d8} /* (20, 12, 14) {real, imag} */,
  {32'h40a8f5ca, 32'hc03c982e} /* (20, 12, 13) {real, imag} */,
  {32'h41308152, 32'hc08c9e36} /* (20, 12, 12) {real, imag} */,
  {32'hc141b562, 32'hc0b33d39} /* (20, 12, 11) {real, imag} */,
  {32'h3f839d9e, 32'h3fea79e0} /* (20, 12, 10) {real, imag} */,
  {32'h410b20be, 32'hc0afd5bf} /* (20, 12, 9) {real, imag} */,
  {32'hc1cb1bd0, 32'hbf73c288} /* (20, 12, 8) {real, imag} */,
  {32'hc036d9cc, 32'h4136cc04} /* (20, 12, 7) {real, imag} */,
  {32'h414a230a, 32'h40430740} /* (20, 12, 6) {real, imag} */,
  {32'h4164b39e, 32'hc0ac9d94} /* (20, 12, 5) {real, imag} */,
  {32'hc181ec95, 32'hbf9f3438} /* (20, 12, 4) {real, imag} */,
  {32'h4181fe97, 32'h41a9807c} /* (20, 12, 3) {real, imag} */,
  {32'hc0c898e4, 32'h42411f46} /* (20, 12, 2) {real, imag} */,
  {32'h4181a10e, 32'h41632c59} /* (20, 12, 1) {real, imag} */,
  {32'hbfcaaf8c, 32'hc116774c} /* (20, 12, 0) {real, imag} */,
  {32'h4182702e, 32'hc19aab81} /* (20, 11, 31) {real, imag} */,
  {32'h419fcb69, 32'h41de5477} /* (20, 11, 30) {real, imag} */,
  {32'hbe829310, 32'hc1b1e1bc} /* (20, 11, 29) {real, imag} */,
  {32'h412fb044, 32'h4213ccb1} /* (20, 11, 28) {real, imag} */,
  {32'h41e363a3, 32'h41548f22} /* (20, 11, 27) {real, imag} */,
  {32'hc1aea442, 32'hc15d025f} /* (20, 11, 26) {real, imag} */,
  {32'h41cb0b52, 32'h416c28ae} /* (20, 11, 25) {real, imag} */,
  {32'hc150f038, 32'hc057663b} /* (20, 11, 24) {real, imag} */,
  {32'h40e28fba, 32'h4129fad4} /* (20, 11, 23) {real, imag} */,
  {32'hc18193a6, 32'hc1a7e9c3} /* (20, 11, 22) {real, imag} */,
  {32'hc0f7a767, 32'h404b1168} /* (20, 11, 21) {real, imag} */,
  {32'h40c49534, 32'h40c61bc7} /* (20, 11, 20) {real, imag} */,
  {32'h40b5ae55, 32'hc03b1368} /* (20, 11, 19) {real, imag} */,
  {32'hbea7a4c4, 32'hc0613ec2} /* (20, 11, 18) {real, imag} */,
  {32'h3fdf7880, 32'hc02fc419} /* (20, 11, 17) {real, imag} */,
  {32'h3e2dd810, 32'h3ff6a310} /* (20, 11, 16) {real, imag} */,
  {32'hc098c970, 32'h3e35a510} /* (20, 11, 15) {real, imag} */,
  {32'h3f27b822, 32'h40d130df} /* (20, 11, 14) {real, imag} */,
  {32'hc1237dfa, 32'h412fc60f} /* (20, 11, 13) {real, imag} */,
  {32'hc12d0314, 32'h411c2962} /* (20, 11, 12) {real, imag} */,
  {32'h4121dde0, 32'hc18ac722} /* (20, 11, 11) {real, imag} */,
  {32'hbf1076f0, 32'hc1195dcc} /* (20, 11, 10) {real, imag} */,
  {32'h4186d9ca, 32'hc16a7714} /* (20, 11, 9) {real, imag} */,
  {32'h4181ff48, 32'hc12c6ca9} /* (20, 11, 8) {real, imag} */,
  {32'hc1c1452a, 32'h40d662f4} /* (20, 11, 7) {real, imag} */,
  {32'hbf9c4878, 32'h40a3031a} /* (20, 11, 6) {real, imag} */,
  {32'hc1c188d3, 32'hc14bbb88} /* (20, 11, 5) {real, imag} */,
  {32'h419f4193, 32'h40c1bdd6} /* (20, 11, 4) {real, imag} */,
  {32'hc166e368, 32'h418b82d8} /* (20, 11, 3) {real, imag} */,
  {32'h4175d8f6, 32'h40bbbdcc} /* (20, 11, 2) {real, imag} */,
  {32'h40eeddfe, 32'hc1800077} /* (20, 11, 1) {real, imag} */,
  {32'h40b43ba4, 32'h40e0c874} /* (20, 11, 0) {real, imag} */,
  {32'hc09affa0, 32'hc238a1bf} /* (20, 10, 31) {real, imag} */,
  {32'h4218aa19, 32'hc021c590} /* (20, 10, 30) {real, imag} */,
  {32'h42249596, 32'h4188a290} /* (20, 10, 29) {real, imag} */,
  {32'hbfe1f5d0, 32'h41aab24d} /* (20, 10, 28) {real, imag} */,
  {32'h41a6f207, 32'hc0d1f550} /* (20, 10, 27) {real, imag} */,
  {32'h418b7986, 32'h4210d66c} /* (20, 10, 26) {real, imag} */,
  {32'hc1229a96, 32'h41441cc6} /* (20, 10, 25) {real, imag} */,
  {32'hc18d17e8, 32'h40479a2e} /* (20, 10, 24) {real, imag} */,
  {32'h40b34be7, 32'hbf583920} /* (20, 10, 23) {real, imag} */,
  {32'hc11a7bf8, 32'hc08c8902} /* (20, 10, 22) {real, imag} */,
  {32'hc0fcaede, 32'hc13e21e2} /* (20, 10, 21) {real, imag} */,
  {32'hc13f07ba, 32'h40866c2e} /* (20, 10, 20) {real, imag} */,
  {32'hc0491438, 32'hbfe03688} /* (20, 10, 19) {real, imag} */,
  {32'h3f3941b0, 32'hc085b82a} /* (20, 10, 18) {real, imag} */,
  {32'h4097a9c8, 32'h40e86be2} /* (20, 10, 17) {real, imag} */,
  {32'h40ef283c, 32'hc15b0e8d} /* (20, 10, 16) {real, imag} */,
  {32'hc00eae98, 32'h3f0e5690} /* (20, 10, 15) {real, imag} */,
  {32'hc0fb242e, 32'hc0550cbd} /* (20, 10, 14) {real, imag} */,
  {32'hbfcbb170, 32'h4027c3d0} /* (20, 10, 13) {real, imag} */,
  {32'h4019ef40, 32'hc0257d74} /* (20, 10, 12) {real, imag} */,
  {32'h412818f9, 32'h3e9021c0} /* (20, 10, 11) {real, imag} */,
  {32'h4180a38b, 32'hc1b62534} /* (20, 10, 10) {real, imag} */,
  {32'hbd8c4640, 32'h40838368} /* (20, 10, 9) {real, imag} */,
  {32'h415d7b9f, 32'h412c87f4} /* (20, 10, 8) {real, imag} */,
  {32'h41a373bf, 32'hc1adc391} /* (20, 10, 7) {real, imag} */,
  {32'hbff4a1d8, 32'hc1356360} /* (20, 10, 6) {real, imag} */,
  {32'h4122295c, 32'h421fe7e5} /* (20, 10, 5) {real, imag} */,
  {32'h41a1d108, 32'h41763a06} /* (20, 10, 4) {real, imag} */,
  {32'hc28b8791, 32'h410a4d59} /* (20, 10, 3) {real, imag} */,
  {32'h4207b5e7, 32'h3e9185ec} /* (20, 10, 2) {real, imag} */,
  {32'hc218aa08, 32'hbfc5b5e0} /* (20, 10, 1) {real, imag} */,
  {32'hc02ab4e3, 32'hc213de51} /* (20, 10, 0) {real, imag} */,
  {32'hc1fc0fa5, 32'hc129791e} /* (20, 9, 31) {real, imag} */,
  {32'h41caec94, 32'h416aa152} /* (20, 9, 30) {real, imag} */,
  {32'hc0664f34, 32'hc09cc624} /* (20, 9, 29) {real, imag} */,
  {32'hc15350e8, 32'hc203f8e5} /* (20, 9, 28) {real, imag} */,
  {32'hbf6df7c0, 32'hc2036df9} /* (20, 9, 27) {real, imag} */,
  {32'hc0e1f5c9, 32'hc1d33324} /* (20, 9, 26) {real, imag} */,
  {32'h416d0f0c, 32'h40e18b46} /* (20, 9, 25) {real, imag} */,
  {32'hbfc07dc0, 32'hc0a32db9} /* (20, 9, 24) {real, imag} */,
  {32'h40b08460, 32'h4101f6f4} /* (20, 9, 23) {real, imag} */,
  {32'h403ded6a, 32'hbdabebc0} /* (20, 9, 22) {real, imag} */,
  {32'hc0832316, 32'h40cf9aba} /* (20, 9, 21) {real, imag} */,
  {32'hc088bf00, 32'h41adc85e} /* (20, 9, 20) {real, imag} */,
  {32'h415e2e03, 32'hc13000d6} /* (20, 9, 19) {real, imag} */,
  {32'h40333d8d, 32'h4103549e} /* (20, 9, 18) {real, imag} */,
  {32'hc03119fa, 32'h3fbc53b0} /* (20, 9, 17) {real, imag} */,
  {32'h3f87cc40, 32'hc0dbae64} /* (20, 9, 16) {real, imag} */,
  {32'hc00f4cb6, 32'h40c61e9c} /* (20, 9, 15) {real, imag} */,
  {32'h409d1012, 32'h4156fb52} /* (20, 9, 14) {real, imag} */,
  {32'hc00d84bc, 32'hc19d6f50} /* (20, 9, 13) {real, imag} */,
  {32'h419dc3e0, 32'h410c7a29} /* (20, 9, 12) {real, imag} */,
  {32'h415a4c7f, 32'h40de600a} /* (20, 9, 11) {real, imag} */,
  {32'hc0ea70dd, 32'h4135d9a6} /* (20, 9, 10) {real, imag} */,
  {32'hc16b1e28, 32'h4123a358} /* (20, 9, 9) {real, imag} */,
  {32'hc192249e, 32'h416ca85e} /* (20, 9, 8) {real, imag} */,
  {32'h40d3b699, 32'hc0f64a0c} /* (20, 9, 7) {real, imag} */,
  {32'h4046e90a, 32'hc2129732} /* (20, 9, 6) {real, imag} */,
  {32'h424afb41, 32'h41a0d256} /* (20, 9, 5) {real, imag} */,
  {32'hc1ff466a, 32'h4192e2c5} /* (20, 9, 4) {real, imag} */,
  {32'h419d46c6, 32'hc1d3f7b6} /* (20, 9, 3) {real, imag} */,
  {32'hc1759f0f, 32'h3f965e54} /* (20, 9, 2) {real, imag} */,
  {32'hc112abd2, 32'h428072bb} /* (20, 9, 1) {real, imag} */,
  {32'hc20314a6, 32'hc2026f76} /* (20, 9, 0) {real, imag} */,
  {32'hc19f9f86, 32'hc02e17d4} /* (20, 8, 31) {real, imag} */,
  {32'hc1c6da12, 32'hc1e5819a} /* (20, 8, 30) {real, imag} */,
  {32'hc228f174, 32'h40a07a30} /* (20, 8, 29) {real, imag} */,
  {32'h41bf5e48, 32'hc143bc3f} /* (20, 8, 28) {real, imag} */,
  {32'h41100e63, 32'hc13a8824} /* (20, 8, 27) {real, imag} */,
  {32'h3fa84684, 32'h40a3ca4c} /* (20, 8, 26) {real, imag} */,
  {32'hc13de882, 32'h415235f2} /* (20, 8, 25) {real, imag} */,
  {32'hc0beeda5, 32'hc2174867} /* (20, 8, 24) {real, imag} */,
  {32'h414f847a, 32'h4162c1da} /* (20, 8, 23) {real, imag} */,
  {32'h40787c00, 32'hc1bd8e1f} /* (20, 8, 22) {real, imag} */,
  {32'h40b98470, 32'h41a0ba5f} /* (20, 8, 21) {real, imag} */,
  {32'h3fb58fb0, 32'hc0eb77a2} /* (20, 8, 20) {real, imag} */,
  {32'h4021ad68, 32'hbfd2f860} /* (20, 8, 19) {real, imag} */,
  {32'h3f850500, 32'hc1031b30} /* (20, 8, 18) {real, imag} */,
  {32'hc023b3df, 32'h400505e9} /* (20, 8, 17) {real, imag} */,
  {32'h407d2040, 32'h407063f2} /* (20, 8, 16) {real, imag} */,
  {32'h404707ed, 32'hc0786f9f} /* (20, 8, 15) {real, imag} */,
  {32'hc145a982, 32'h414673f6} /* (20, 8, 14) {real, imag} */,
  {32'h41d2889f, 32'hc04001e0} /* (20, 8, 13) {real, imag} */,
  {32'h41a7fcef, 32'hc1cb9bd0} /* (20, 8, 12) {real, imag} */,
  {32'hc09b6590, 32'h415eb99a} /* (20, 8, 11) {real, imag} */,
  {32'hc216c919, 32'hc1ef0839} /* (20, 8, 10) {real, imag} */,
  {32'hbe5c9860, 32'hc14e5394} /* (20, 8, 9) {real, imag} */,
  {32'hbd217d80, 32'hc1e02992} /* (20, 8, 8) {real, imag} */,
  {32'hc2237882, 32'h3fe803a0} /* (20, 8, 7) {real, imag} */,
  {32'h4153dcc0, 32'hc250d282} /* (20, 8, 6) {real, imag} */,
  {32'hc12f9b23, 32'h425fb01f} /* (20, 8, 5) {real, imag} */,
  {32'hc2030678, 32'hc1cdd7c0} /* (20, 8, 4) {real, imag} */,
  {32'h41963555, 32'hc28e8f79} /* (20, 8, 3) {real, imag} */,
  {32'hc19b58fe, 32'hc155917d} /* (20, 8, 2) {real, imag} */,
  {32'h412df679, 32'h418fb370} /* (20, 8, 1) {real, imag} */,
  {32'h4286ab94, 32'hc03ae1a2} /* (20, 8, 0) {real, imag} */,
  {32'h412bab34, 32'h426ae9f5} /* (20, 7, 31) {real, imag} */,
  {32'hc1471d4c, 32'hc0a237b9} /* (20, 7, 30) {real, imag} */,
  {32'hc2165862, 32'h428c71ce} /* (20, 7, 29) {real, imag} */,
  {32'hc08888c8, 32'hc1ae0ffd} /* (20, 7, 28) {real, imag} */,
  {32'h3f9075b0, 32'h4188f546} /* (20, 7, 27) {real, imag} */,
  {32'h41e08ce6, 32'hc2647b68} /* (20, 7, 26) {real, imag} */,
  {32'h4171add5, 32'h41c20f62} /* (20, 7, 25) {real, imag} */,
  {32'h40d72718, 32'h411563c2} /* (20, 7, 24) {real, imag} */,
  {32'hc196adbe, 32'h41250b5a} /* (20, 7, 23) {real, imag} */,
  {32'h417c08cc, 32'h4192367a} /* (20, 7, 22) {real, imag} */,
  {32'h400385ec, 32'h414d2a21} /* (20, 7, 21) {real, imag} */,
  {32'h40579294, 32'hc08c468d} /* (20, 7, 20) {real, imag} */,
  {32'hc00df9a4, 32'hbfa59460} /* (20, 7, 19) {real, imag} */,
  {32'h415491ed, 32'h3fb5aeb4} /* (20, 7, 18) {real, imag} */,
  {32'hc1022b5c, 32'hc01d1730} /* (20, 7, 17) {real, imag} */,
  {32'hc16b9cd4, 32'h3f3ef690} /* (20, 7, 16) {real, imag} */,
  {32'hc0d06829, 32'h40fbf758} /* (20, 7, 15) {real, imag} */,
  {32'h416aa681, 32'h40beb8e3} /* (20, 7, 14) {real, imag} */,
  {32'hbfe9ed18, 32'h41846bdc} /* (20, 7, 13) {real, imag} */,
  {32'hc11af35e, 32'hc0a526b7} /* (20, 7, 12) {real, imag} */,
  {32'h40497fbc, 32'h409b75b6} /* (20, 7, 11) {real, imag} */,
  {32'hc18bf606, 32'h419f608e} /* (20, 7, 10) {real, imag} */,
  {32'h41d6d79e, 32'h4172a30c} /* (20, 7, 9) {real, imag} */,
  {32'hc1aed59c, 32'h423b12b8} /* (20, 7, 8) {real, imag} */,
  {32'h4107836b, 32'hc11087a3} /* (20, 7, 7) {real, imag} */,
  {32'h42208469, 32'hc1c85f5f} /* (20, 7, 6) {real, imag} */,
  {32'hc22a5d1e, 32'hc1e7fb16} /* (20, 7, 5) {real, imag} */,
  {32'hc1a8c626, 32'hc1998fc7} /* (20, 7, 4) {real, imag} */,
  {32'hc0ed0a68, 32'hc1704a0e} /* (20, 7, 3) {real, imag} */,
  {32'h42477d48, 32'hc1266738} /* (20, 7, 2) {real, imag} */,
  {32'h41ca2416, 32'hc2082c49} /* (20, 7, 1) {real, imag} */,
  {32'hc205301e, 32'hc1e2fc64} /* (20, 7, 0) {real, imag} */,
  {32'hc1e564ba, 32'h41388bc6} /* (20, 6, 31) {real, imag} */,
  {32'hc2a2441a, 32'hc1c45bfc} /* (20, 6, 30) {real, imag} */,
  {32'h41b635bc, 32'hc24d3070} /* (20, 6, 29) {real, imag} */,
  {32'h41f494a5, 32'h41184e48} /* (20, 6, 28) {real, imag} */,
  {32'h4233d40c, 32'h414ad727} /* (20, 6, 27) {real, imag} */,
  {32'hc28b7e81, 32'h41628d0e} /* (20, 6, 26) {real, imag} */,
  {32'h41474256, 32'h414e1a5d} /* (20, 6, 25) {real, imag} */,
  {32'h42186740, 32'hc16ef5fc} /* (20, 6, 24) {real, imag} */,
  {32'hc17aca42, 32'hc14e4614} /* (20, 6, 23) {real, imag} */,
  {32'h4098d558, 32'h41a8abaf} /* (20, 6, 22) {real, imag} */,
  {32'hc0d8ac84, 32'h414100ea} /* (20, 6, 21) {real, imag} */,
  {32'hc0f2271d, 32'hc1a60ec4} /* (20, 6, 20) {real, imag} */,
  {32'h41a176b8, 32'h3f86c224} /* (20, 6, 19) {real, imag} */,
  {32'h40409d40, 32'hc17729ae} /* (20, 6, 18) {real, imag} */,
  {32'h412203e5, 32'h40cea330} /* (20, 6, 17) {real, imag} */,
  {32'hbef56060, 32'h40bf9368} /* (20, 6, 16) {real, imag} */,
  {32'hc11dcef3, 32'hc12df1fc} /* (20, 6, 15) {real, imag} */,
  {32'h4149c174, 32'hbeec4290} /* (20, 6, 14) {real, imag} */,
  {32'h40be275a, 32'h40cf61df} /* (20, 6, 13) {real, imag} */,
  {32'h4165d1ca, 32'hc11cca43} /* (20, 6, 12) {real, imag} */,
  {32'hc101ab82, 32'h40159e62} /* (20, 6, 11) {real, imag} */,
  {32'h40cbe890, 32'h408bd5ec} /* (20, 6, 10) {real, imag} */,
  {32'hc1aa1f53, 32'hc165c14c} /* (20, 6, 9) {real, imag} */,
  {32'hc1c2fe88, 32'hc17b798c} /* (20, 6, 8) {real, imag} */,
  {32'h425192de, 32'h3fb41970} /* (20, 6, 7) {real, imag} */,
  {32'h40457a20, 32'h41a0f5df} /* (20, 6, 6) {real, imag} */,
  {32'h408d6e9c, 32'hc19ae324} /* (20, 6, 5) {real, imag} */,
  {32'hc1524626, 32'h4294095b} /* (20, 6, 4) {real, imag} */,
  {32'h42645546, 32'hc1b97037} /* (20, 6, 3) {real, imag} */,
  {32'h41cfb551, 32'hbf5f2170} /* (20, 6, 2) {real, imag} */,
  {32'hc1e8409a, 32'hc26c382e} /* (20, 6, 1) {real, imag} */,
  {32'hc106854b, 32'hc0cb1c98} /* (20, 6, 0) {real, imag} */,
  {32'h41d2775d, 32'hbfa0cfe0} /* (20, 5, 31) {real, imag} */,
  {32'h403e7b3c, 32'hc14c9a02} /* (20, 5, 30) {real, imag} */,
  {32'hc2771111, 32'hc2197907} /* (20, 5, 29) {real, imag} */,
  {32'hc1a9373b, 32'h407382e8} /* (20, 5, 28) {real, imag} */,
  {32'h4189fd8f, 32'h4200789d} /* (20, 5, 27) {real, imag} */,
  {32'hc129a11d, 32'h424e09b0} /* (20, 5, 26) {real, imag} */,
  {32'hc16c9ba5, 32'h40f0c6f4} /* (20, 5, 25) {real, imag} */,
  {32'hc248a42e, 32'hc1688a0e} /* (20, 5, 24) {real, imag} */,
  {32'h41dfd95f, 32'h422e80a0} /* (20, 5, 23) {real, imag} */,
  {32'hc12af941, 32'hc0874a7b} /* (20, 5, 22) {real, imag} */,
  {32'hc1a7cffa, 32'hc21a1cb0} /* (20, 5, 21) {real, imag} */,
  {32'hc04c7ce2, 32'h41940849} /* (20, 5, 20) {real, imag} */,
  {32'h40bb018c, 32'hc0bc9f60} /* (20, 5, 19) {real, imag} */,
  {32'hc1270463, 32'h4090c23f} /* (20, 5, 18) {real, imag} */,
  {32'h40a6a39a, 32'h3f5216b0} /* (20, 5, 17) {real, imag} */,
  {32'hc15898c2, 32'h40293b64} /* (20, 5, 16) {real, imag} */,
  {32'hbfd3df18, 32'h4132d18d} /* (20, 5, 15) {real, imag} */,
  {32'h3f7b8710, 32'h40c48a45} /* (20, 5, 14) {real, imag} */,
  {32'h3fdd78f0, 32'h4130b69a} /* (20, 5, 13) {real, imag} */,
  {32'hbfaa7fcc, 32'hc11117ba} /* (20, 5, 12) {real, imag} */,
  {32'h41bca24e, 32'h40a599f0} /* (20, 5, 11) {real, imag} */,
  {32'hc185d7e2, 32'hc0b9220d} /* (20, 5, 10) {real, imag} */,
  {32'hc1dee443, 32'h41a5a288} /* (20, 5, 9) {real, imag} */,
  {32'hc01e3080, 32'hc24965a0} /* (20, 5, 8) {real, imag} */,
  {32'h421579d2, 32'hc2051716} /* (20, 5, 7) {real, imag} */,
  {32'hc2058488, 32'h41c6b86f} /* (20, 5, 6) {real, imag} */,
  {32'hc20bf0d0, 32'h42438245} /* (20, 5, 5) {real, imag} */,
  {32'hc12a8280, 32'h423e9fb0} /* (20, 5, 4) {real, imag} */,
  {32'hc1b227ce, 32'hc1241475} /* (20, 5, 3) {real, imag} */,
  {32'hc20745ad, 32'hbdecc440} /* (20, 5, 2) {real, imag} */,
  {32'h41d5978b, 32'h424f8085} /* (20, 5, 1) {real, imag} */,
  {32'h41e65c8d, 32'h4177df6f} /* (20, 5, 0) {real, imag} */,
  {32'h41b283a3, 32'hc102ed61} /* (20, 4, 31) {real, imag} */,
  {32'h4210b3cb, 32'hc1f97558} /* (20, 4, 30) {real, imag} */,
  {32'hc26297c0, 32'h40995458} /* (20, 4, 29) {real, imag} */,
  {32'hc195de12, 32'hc1232a70} /* (20, 4, 28) {real, imag} */,
  {32'h3f0a0600, 32'h4290595e} /* (20, 4, 27) {real, imag} */,
  {32'h42369c14, 32'h41b652ae} /* (20, 4, 26) {real, imag} */,
  {32'h413096c1, 32'h40a9b1e8} /* (20, 4, 25) {real, imag} */,
  {32'hc2241a4c, 32'hc224f2cc} /* (20, 4, 24) {real, imag} */,
  {32'h42001a50, 32'hc1722d48} /* (20, 4, 23) {real, imag} */,
  {32'h41957581, 32'hc1b92c28} /* (20, 4, 22) {real, imag} */,
  {32'hc21d9fe8, 32'hc12497a4} /* (20, 4, 21) {real, imag} */,
  {32'hc1667447, 32'h40b00097} /* (20, 4, 20) {real, imag} */,
  {32'h40ba77c2, 32'hbfbd4920} /* (20, 4, 19) {real, imag} */,
  {32'h40a127ce, 32'h41b2c29c} /* (20, 4, 18) {real, imag} */,
  {32'h40d81a03, 32'hc12b5204} /* (20, 4, 17) {real, imag} */,
  {32'hc04ed36c, 32'h4082df00} /* (20, 4, 16) {real, imag} */,
  {32'h40e88ac7, 32'hc0abfec0} /* (20, 4, 15) {real, imag} */,
  {32'h41262f0b, 32'hc01ce264} /* (20, 4, 14) {real, imag} */,
  {32'hc1685fb9, 32'hc1596314} /* (20, 4, 13) {real, imag} */,
  {32'h414602f3, 32'h3ffcc3d4} /* (20, 4, 12) {real, imag} */,
  {32'hc049d940, 32'hc10aad3c} /* (20, 4, 11) {real, imag} */,
  {32'hc238aa86, 32'hc1c104f8} /* (20, 4, 10) {real, imag} */,
  {32'h40d52c82, 32'h424140e8} /* (20, 4, 9) {real, imag} */,
  {32'hc1bfb2f0, 32'h416cff80} /* (20, 4, 8) {real, imag} */,
  {32'h40fb45ee, 32'h420e7933} /* (20, 4, 7) {real, imag} */,
  {32'hc018ab98, 32'hc191cc2a} /* (20, 4, 6) {real, imag} */,
  {32'hc2460848, 32'h40a59368} /* (20, 4, 5) {real, imag} */,
  {32'h411aa442, 32'hc1d16654} /* (20, 4, 4) {real, imag} */,
  {32'hc13ef348, 32'h423922df} /* (20, 4, 3) {real, imag} */,
  {32'hc240c5f9, 32'hc1d73330} /* (20, 4, 2) {real, imag} */,
  {32'hc1745042, 32'hc1b34316} /* (20, 4, 1) {real, imag} */,
  {32'h41748423, 32'hc2456c40} /* (20, 4, 0) {real, imag} */,
  {32'h41940647, 32'h428c643a} /* (20, 3, 31) {real, imag} */,
  {32'h41e4cc6e, 32'hc19b2150} /* (20, 3, 30) {real, imag} */,
  {32'hc189feb5, 32'h42e99495} /* (20, 3, 29) {real, imag} */,
  {32'h4218e52e, 32'hc27ca830} /* (20, 3, 28) {real, imag} */,
  {32'hc1d076a6, 32'h40e7a043} /* (20, 3, 27) {real, imag} */,
  {32'h40b30e4b, 32'h41fe2def} /* (20, 3, 26) {real, imag} */,
  {32'h41adaa8f, 32'h428001d8} /* (20, 3, 25) {real, imag} */,
  {32'hc1e663f8, 32'h40dd3ef0} /* (20, 3, 24) {real, imag} */,
  {32'hc0da6118, 32'hbf313f50} /* (20, 3, 23) {real, imag} */,
  {32'hc211d986, 32'hc1883252} /* (20, 3, 22) {real, imag} */,
  {32'h3c9eb000, 32'h410bc22a} /* (20, 3, 21) {real, imag} */,
  {32'h418868ae, 32'h40cb1d0c} /* (20, 3, 20) {real, imag} */,
  {32'hc0e67350, 32'h410d4d98} /* (20, 3, 19) {real, imag} */,
  {32'hc0ea52fd, 32'h416bde98} /* (20, 3, 18) {real, imag} */,
  {32'hbf818870, 32'h40a0165e} /* (20, 3, 17) {real, imag} */,
  {32'h403f083c, 32'hc0ad7157} /* (20, 3, 16) {real, imag} */,
  {32'hc198f64b, 32'hc1abca4c} /* (20, 3, 15) {real, imag} */,
  {32'h4068627a, 32'hc0196b00} /* (20, 3, 14) {real, imag} */,
  {32'hc1d4b3ce, 32'hc12162f8} /* (20, 3, 13) {real, imag} */,
  {32'hc0ce242a, 32'h41d11cbd} /* (20, 3, 12) {real, imag} */,
  {32'hc0a2b904, 32'hc0215dde} /* (20, 3, 11) {real, imag} */,
  {32'hc0a754ec, 32'hc238dd26} /* (20, 3, 10) {real, imag} */,
  {32'h41b4d338, 32'h4191baf8} /* (20, 3, 9) {real, imag} */,
  {32'h420daa80, 32'hc1c95422} /* (20, 3, 8) {real, imag} */,
  {32'hc093e394, 32'h41b416a6} /* (20, 3, 7) {real, imag} */,
  {32'hc052e726, 32'hc0381568} /* (20, 3, 6) {real, imag} */,
  {32'h40bfbafa, 32'hc15f09e4} /* (20, 3, 5) {real, imag} */,
  {32'h42274c3c, 32'h42100140} /* (20, 3, 4) {real, imag} */,
  {32'h4240fe1e, 32'h425505ea} /* (20, 3, 3) {real, imag} */,
  {32'h4251410b, 32'h41a0ac20} /* (20, 3, 2) {real, imag} */,
  {32'h4141b302, 32'hc301c2bd} /* (20, 3, 1) {real, imag} */,
  {32'h413ddd3f, 32'h40cafd35} /* (20, 3, 0) {real, imag} */,
  {32'h4233d0a6, 32'hc3053a3a} /* (20, 2, 31) {real, imag} */,
  {32'hc1c48315, 32'hc01d80e4} /* (20, 2, 30) {real, imag} */,
  {32'h42987cd0, 32'h425017d9} /* (20, 2, 29) {real, imag} */,
  {32'h3fb43b14, 32'h4257f5cc} /* (20, 2, 28) {real, imag} */,
  {32'h42009e99, 32'h41b5b21f} /* (20, 2, 27) {real, imag} */,
  {32'h41f5041a, 32'hc1a28595} /* (20, 2, 26) {real, imag} */,
  {32'h42a11acc, 32'h41869d34} /* (20, 2, 25) {real, imag} */,
  {32'hc0d222ed, 32'h402b23b2} /* (20, 2, 24) {real, imag} */,
  {32'hc12e4afe, 32'hc1a72802} /* (20, 2, 23) {real, imag} */,
  {32'hbf968cb0, 32'hc0ad53ce} /* (20, 2, 22) {real, imag} */,
  {32'hbfb28d90, 32'hc15278e2} /* (20, 2, 21) {real, imag} */,
  {32'h40d86208, 32'h3ffe3f18} /* (20, 2, 20) {real, imag} */,
  {32'hc110c4a5, 32'hc0040707} /* (20, 2, 19) {real, imag} */,
  {32'h415c412b, 32'h41418702} /* (20, 2, 18) {real, imag} */,
  {32'h4116d29c, 32'h4135a2cc} /* (20, 2, 17) {real, imag} */,
  {32'hc1133fa6, 32'h413dd3c9} /* (20, 2, 16) {real, imag} */,
  {32'hc115ba30, 32'hc0487010} /* (20, 2, 15) {real, imag} */,
  {32'hc1878150, 32'hc1125f24} /* (20, 2, 14) {real, imag} */,
  {32'hc0f178e6, 32'h40990aec} /* (20, 2, 13) {real, imag} */,
  {32'h4210c0db, 32'hc1cbe5ca} /* (20, 2, 12) {real, imag} */,
  {32'hc1c96da2, 32'hc0a1ae0c} /* (20, 2, 11) {real, imag} */,
  {32'hc0e6d228, 32'hc0437b90} /* (20, 2, 10) {real, imag} */,
  {32'h41db5c19, 32'hc0df6792} /* (20, 2, 9) {real, imag} */,
  {32'h41b339fe, 32'hc0e9ab35} /* (20, 2, 8) {real, imag} */,
  {32'h420a7a81, 32'hc234483f} /* (20, 2, 7) {real, imag} */,
  {32'h41a6f16e, 32'h40571e78} /* (20, 2, 6) {real, imag} */,
  {32'h420b3e31, 32'h41aadd2d} /* (20, 2, 5) {real, imag} */,
  {32'h41096464, 32'h41920623} /* (20, 2, 4) {real, imag} */,
  {32'h4228863a, 32'hc208be41} /* (20, 2, 3) {real, imag} */,
  {32'hc26c803e, 32'hc1a26fb8} /* (20, 2, 2) {real, imag} */,
  {32'hc1b2582b, 32'h41494ad4} /* (20, 2, 1) {real, imag} */,
  {32'h41611dda, 32'h42271ca0} /* (20, 2, 0) {real, imag} */,
  {32'hc218ae52, 32'h411d7160} /* (20, 1, 31) {real, imag} */,
  {32'hc0711300, 32'hc19f8579} /* (20, 1, 30) {real, imag} */,
  {32'h42020460, 32'hc16679fa} /* (20, 1, 29) {real, imag} */,
  {32'hc1f44a9b, 32'h40cc5364} /* (20, 1, 28) {real, imag} */,
  {32'h424c33b0, 32'h42078deb} /* (20, 1, 27) {real, imag} */,
  {32'h418bbb7a, 32'hc20d0d5b} /* (20, 1, 26) {real, imag} */,
  {32'hc18b7cfb, 32'hc176c98c} /* (20, 1, 25) {real, imag} */,
  {32'h41e8fb15, 32'hc1056a99} /* (20, 1, 24) {real, imag} */,
  {32'h422ff1b2, 32'hc042511c} /* (20, 1, 23) {real, imag} */,
  {32'h421afefa, 32'h40f624fc} /* (20, 1, 22) {real, imag} */,
  {32'hc187ed2f, 32'hc25b4cac} /* (20, 1, 21) {real, imag} */,
  {32'h40f48bc2, 32'h40b8c476} /* (20, 1, 20) {real, imag} */,
  {32'h418eb496, 32'hc202ff30} /* (20, 1, 19) {real, imag} */,
  {32'h3eaada40, 32'hbf23ccf8} /* (20, 1, 18) {real, imag} */,
  {32'hc1ae7d66, 32'hc196c1ff} /* (20, 1, 17) {real, imag} */,
  {32'hbd0ddc00, 32'h4122eb34} /* (20, 1, 16) {real, imag} */,
  {32'hc108f3f0, 32'hc064b118} /* (20, 1, 15) {real, imag} */,
  {32'h41b56a59, 32'hc0f6e921} /* (20, 1, 14) {real, imag} */,
  {32'h4091d598, 32'hc19b58ba} /* (20, 1, 13) {real, imag} */,
  {32'h3fe84380, 32'h40a23d7e} /* (20, 1, 12) {real, imag} */,
  {32'h422dadb2, 32'h413bbbc8} /* (20, 1, 11) {real, imag} */,
  {32'hc1f701cc, 32'h414dd36c} /* (20, 1, 10) {real, imag} */,
  {32'hc0e91ccc, 32'hc128adb5} /* (20, 1, 9) {real, imag} */,
  {32'hc1f837c5, 32'hc1308fb3} /* (20, 1, 8) {real, imag} */,
  {32'h42163420, 32'hc28b13e6} /* (20, 1, 7) {real, imag} */,
  {32'hc286789e, 32'h3fddd920} /* (20, 1, 6) {real, imag} */,
  {32'hc1440f2a, 32'hc168d44b} /* (20, 1, 5) {real, imag} */,
  {32'h402091e8, 32'h427102e6} /* (20, 1, 4) {real, imag} */,
  {32'hc210b7a4, 32'h41d27d33} /* (20, 1, 3) {real, imag} */,
  {32'hc2a2b510, 32'hc0e25b8d} /* (20, 1, 2) {real, imag} */,
  {32'hc2967151, 32'hc1c40f14} /* (20, 1, 1) {real, imag} */,
  {32'h4230e4db, 32'hc2134f86} /* (20, 1, 0) {real, imag} */,
  {32'h4132baaa, 32'h4233e55a} /* (20, 0, 31) {real, imag} */,
  {32'hc1d3c8bc, 32'hc26e0460} /* (20, 0, 30) {real, imag} */,
  {32'hc274e2b8, 32'hc128141c} /* (20, 0, 29) {real, imag} */,
  {32'h4204e0c6, 32'h41abb39f} /* (20, 0, 28) {real, imag} */,
  {32'hc252234c, 32'h4112f848} /* (20, 0, 27) {real, imag} */,
  {32'h42c8835c, 32'hc23dc4e6} /* (20, 0, 26) {real, imag} */,
  {32'hc145886c, 32'h40771538} /* (20, 0, 25) {real, imag} */,
  {32'h41e5130a, 32'h40b9eb54} /* (20, 0, 24) {real, imag} */,
  {32'h4253d6fc, 32'h42457802} /* (20, 0, 23) {real, imag} */,
  {32'h41367f90, 32'h41eec6ed} /* (20, 0, 22) {real, imag} */,
  {32'h40ced4e2, 32'h418def90} /* (20, 0, 21) {real, imag} */,
  {32'hc1a80b64, 32'h41a30765} /* (20, 0, 20) {real, imag} */,
  {32'hc09af6a0, 32'h4124209c} /* (20, 0, 19) {real, imag} */,
  {32'h414e65d9, 32'h40cbff82} /* (20, 0, 18) {real, imag} */,
  {32'h40574e54, 32'hc183d1fc} /* (20, 0, 17) {real, imag} */,
  {32'hbff37480, 32'h4090c840} /* (20, 0, 16) {real, imag} */,
  {32'hc0897280, 32'h40c294e6} /* (20, 0, 15) {real, imag} */,
  {32'h3f84ce18, 32'hc1c17ca0} /* (20, 0, 14) {real, imag} */,
  {32'h40d54f30, 32'h42070339} /* (20, 0, 13) {real, imag} */,
  {32'h40b3f464, 32'h41670b7a} /* (20, 0, 12) {real, imag} */,
  {32'hc20fc0dc, 32'hbff5fd08} /* (20, 0, 11) {real, imag} */,
  {32'h417df618, 32'h405c6c78} /* (20, 0, 10) {real, imag} */,
  {32'hc1905050, 32'hc1a4f143} /* (20, 0, 9) {real, imag} */,
  {32'h427f22e7, 32'hc213374e} /* (20, 0, 8) {real, imag} */,
  {32'hc0b52918, 32'hc210fd68} /* (20, 0, 7) {real, imag} */,
  {32'h42024de7, 32'h421f8c36} /* (20, 0, 6) {real, imag} */,
  {32'h429641c2, 32'h42b6d1fb} /* (20, 0, 5) {real, imag} */,
  {32'h3e877540, 32'hc1e91c41} /* (20, 0, 4) {real, imag} */,
  {32'h41470246, 32'h410980dc} /* (20, 0, 3) {real, imag} */,
  {32'hc24f7bba, 32'h41ab0200} /* (20, 0, 2) {real, imag} */,
  {32'hc0e9a333, 32'hc07bb528} /* (20, 0, 1) {real, imag} */,
  {32'hc2073d8b, 32'h42455be4} /* (20, 0, 0) {real, imag} */,
  {32'hc28d9a11, 32'h40a786bb} /* (19, 31, 31) {real, imag} */,
  {32'hc180ed1c, 32'hc2775b3c} /* (19, 31, 30) {real, imag} */,
  {32'h418b0954, 32'h42000aac} /* (19, 31, 29) {real, imag} */,
  {32'hc1304500, 32'hc2201a04} /* (19, 31, 28) {real, imag} */,
  {32'hc1a02c73, 32'hc0f85674} /* (19, 31, 27) {real, imag} */,
  {32'h42048814, 32'hc0c4c7ac} /* (19, 31, 26) {real, imag} */,
  {32'hc1fb0602, 32'h40c1d230} /* (19, 31, 25) {real, imag} */,
  {32'hc15316dc, 32'hc02d40a8} /* (19, 31, 24) {real, imag} */,
  {32'hc1aab0e3, 32'h4295ce25} /* (19, 31, 23) {real, imag} */,
  {32'h4161840c, 32'hc0fc6b4c} /* (19, 31, 22) {real, imag} */,
  {32'h424b101b, 32'h401813dc} /* (19, 31, 21) {real, imag} */,
  {32'hc110ccb0, 32'h410c7944} /* (19, 31, 20) {real, imag} */,
  {32'h40ae2d58, 32'h4035f39a} /* (19, 31, 19) {real, imag} */,
  {32'h4022b69a, 32'h4153c7d4} /* (19, 31, 18) {real, imag} */,
  {32'hc05a1b00, 32'hc0fc1b90} /* (19, 31, 17) {real, imag} */,
  {32'h41945099, 32'h41f0762a} /* (19, 31, 16) {real, imag} */,
  {32'hc15e9898, 32'h3fce7d58} /* (19, 31, 15) {real, imag} */,
  {32'h4039d6c2, 32'hc0fee6d0} /* (19, 31, 14) {real, imag} */,
  {32'h41169e28, 32'hbf86998c} /* (19, 31, 13) {real, imag} */,
  {32'hc20f09d0, 32'hc09075ab} /* (19, 31, 12) {real, imag} */,
  {32'hc17f26a4, 32'hc0c3247a} /* (19, 31, 11) {real, imag} */,
  {32'h41754de4, 32'hc08e50e8} /* (19, 31, 10) {real, imag} */,
  {32'h4130ee5a, 32'hc1fecf0c} /* (19, 31, 9) {real, imag} */,
  {32'h42101195, 32'hc22c4078} /* (19, 31, 8) {real, imag} */,
  {32'h414112ac, 32'hc1daea74} /* (19, 31, 7) {real, imag} */,
  {32'h4191a471, 32'hc0709518} /* (19, 31, 6) {real, imag} */,
  {32'hc18e4b49, 32'hc259f97c} /* (19, 31, 5) {real, imag} */,
  {32'h4190f338, 32'h404e5080} /* (19, 31, 4) {real, imag} */,
  {32'h42c3cca7, 32'hc1205c62} /* (19, 31, 3) {real, imag} */,
  {32'h421ab010, 32'hc1e082cf} /* (19, 31, 2) {real, imag} */,
  {32'h428355ff, 32'hc19bcb1f} /* (19, 31, 1) {real, imag} */,
  {32'h423cd08e, 32'hc1a86d96} /* (19, 31, 0) {real, imag} */,
  {32'h4211e092, 32'h42c23ad2} /* (19, 30, 31) {real, imag} */,
  {32'hc1e45859, 32'hc26647bd} /* (19, 30, 30) {real, imag} */,
  {32'h41c5c003, 32'h4101fc64} /* (19, 30, 29) {real, imag} */,
  {32'h4109dac6, 32'hc2826a2d} /* (19, 30, 28) {real, imag} */,
  {32'hc1b799a0, 32'h4269a9aa} /* (19, 30, 27) {real, imag} */,
  {32'hc236a86c, 32'h41efa946} /* (19, 30, 26) {real, imag} */,
  {32'hc18ee4c6, 32'h41f3459e} /* (19, 30, 25) {real, imag} */,
  {32'hc255adae, 32'hc205816e} /* (19, 30, 24) {real, imag} */,
  {32'hc1bd2ed2, 32'h4130871c} /* (19, 30, 23) {real, imag} */,
  {32'hc10d1ce4, 32'hc07b1434} /* (19, 30, 22) {real, imag} */,
  {32'h3fc76f78, 32'hc18bb919} /* (19, 30, 21) {real, imag} */,
  {32'hc19b7f35, 32'h41b0e660} /* (19, 30, 20) {real, imag} */,
  {32'hbfb42e10, 32'h41893b3c} /* (19, 30, 19) {real, imag} */,
  {32'h41143d06, 32'hc19fe072} /* (19, 30, 18) {real, imag} */,
  {32'h4164df02, 32'h411ed1fc} /* (19, 30, 17) {real, imag} */,
  {32'h40b148dc, 32'hbfa3e6d8} /* (19, 30, 16) {real, imag} */,
  {32'hc0029888, 32'h40be8b38} /* (19, 30, 15) {real, imag} */,
  {32'h41839c9f, 32'hc155d1ec} /* (19, 30, 14) {real, imag} */,
  {32'hc1095f7e, 32'hc0d303b7} /* (19, 30, 13) {real, imag} */,
  {32'hc078a498, 32'hc1024f20} /* (19, 30, 12) {real, imag} */,
  {32'hc1deef58, 32'hc1295c2a} /* (19, 30, 11) {real, imag} */,
  {32'hc1ee4a72, 32'h4109b2bd} /* (19, 30, 10) {real, imag} */,
  {32'h4175ae69, 32'hc2123e1c} /* (19, 30, 9) {real, imag} */,
  {32'hc2103480, 32'h42150106} /* (19, 30, 8) {real, imag} */,
  {32'h41f4e828, 32'h415a3aa0} /* (19, 30, 7) {real, imag} */,
  {32'hc0ce2a80, 32'h428986ae} /* (19, 30, 6) {real, imag} */,
  {32'hc25fe6d0, 32'hc08720fc} /* (19, 30, 5) {real, imag} */,
  {32'h4267c22e, 32'hc1aeb67c} /* (19, 30, 4) {real, imag} */,
  {32'h42acb6a7, 32'h41db8910} /* (19, 30, 3) {real, imag} */,
  {32'h426d9666, 32'hc29ec4be} /* (19, 30, 2) {real, imag} */,
  {32'hc1d12ce9, 32'hc1f17230} /* (19, 30, 1) {real, imag} */,
  {32'h42836aef, 32'hc16f48bf} /* (19, 30, 0) {real, imag} */,
  {32'hc1e02977, 32'h41d11260} /* (19, 29, 31) {real, imag} */,
  {32'hc20a07c7, 32'hc1626e38} /* (19, 29, 30) {real, imag} */,
  {32'hc1b24e63, 32'h404e1f70} /* (19, 29, 29) {real, imag} */,
  {32'h4218d848, 32'hc1c9e4d7} /* (19, 29, 28) {real, imag} */,
  {32'hc153e4a4, 32'hc1c80f21} /* (19, 29, 27) {real, imag} */,
  {32'hc1233aa7, 32'hc117ff88} /* (19, 29, 26) {real, imag} */,
  {32'h40de330c, 32'hc1ee1d0b} /* (19, 29, 25) {real, imag} */,
  {32'hc124082c, 32'hc2618739} /* (19, 29, 24) {real, imag} */,
  {32'h41d01c0d, 32'h4110b7ba} /* (19, 29, 23) {real, imag} */,
  {32'h40417a7d, 32'hc1a287ca} /* (19, 29, 22) {real, imag} */,
  {32'hc19ff200, 32'hc0710f3d} /* (19, 29, 21) {real, imag} */,
  {32'h40a84f28, 32'hc0c2db3a} /* (19, 29, 20) {real, imag} */,
  {32'h4087af02, 32'hc19164c6} /* (19, 29, 19) {real, imag} */,
  {32'hc1ba4e48, 32'h40b17250} /* (19, 29, 18) {real, imag} */,
  {32'h40871fab, 32'h409708a4} /* (19, 29, 17) {real, imag} */,
  {32'hc0fbfc2c, 32'h403e02ae} /* (19, 29, 16) {real, imag} */,
  {32'hc0ec2b3b, 32'hbf6e25e4} /* (19, 29, 15) {real, imag} */,
  {32'hc01827f0, 32'hc1448004} /* (19, 29, 14) {real, imag} */,
  {32'hbebe7848, 32'hc18367ea} /* (19, 29, 13) {real, imag} */,
  {32'hc1711172, 32'hc0f3e84a} /* (19, 29, 12) {real, imag} */,
  {32'hc0500b9c, 32'h402c0173} /* (19, 29, 11) {real, imag} */,
  {32'h410b60db, 32'h41e3e1ca} /* (19, 29, 10) {real, imag} */,
  {32'h40caac34, 32'h3f804a94} /* (19, 29, 9) {real, imag} */,
  {32'hc132e930, 32'hbe6baf00} /* (19, 29, 8) {real, imag} */,
  {32'h41ee4b2f, 32'hc02a47b8} /* (19, 29, 7) {real, imag} */,
  {32'hc085116e, 32'hc2558f00} /* (19, 29, 6) {real, imag} */,
  {32'hc005db36, 32'h416ffc52} /* (19, 29, 5) {real, imag} */,
  {32'h41992750, 32'h41257892} /* (19, 29, 4) {real, imag} */,
  {32'hc14c00aa, 32'h427ef4cd} /* (19, 29, 3) {real, imag} */,
  {32'hc1f38fd1, 32'h41fc867e} /* (19, 29, 2) {real, imag} */,
  {32'hc16d60ca, 32'hc15345e9} /* (19, 29, 1) {real, imag} */,
  {32'hc2274ae4, 32'h3e7e2ca0} /* (19, 29, 0) {real, imag} */,
  {32'h417dfb86, 32'hc214c260} /* (19, 28, 31) {real, imag} */,
  {32'h41ff86f6, 32'h402ab660} /* (19, 28, 30) {real, imag} */,
  {32'hc05f9aec, 32'hc1fd3a7e} /* (19, 28, 29) {real, imag} */,
  {32'hc22b0d6c, 32'hc2bd0410} /* (19, 28, 28) {real, imag} */,
  {32'h400f8720, 32'h422526ee} /* (19, 28, 27) {real, imag} */,
  {32'hc06df71b, 32'h415a1c62} /* (19, 28, 26) {real, imag} */,
  {32'h4181487e, 32'h415212ea} /* (19, 28, 25) {real, imag} */,
  {32'hbe818f80, 32'h421a2134} /* (19, 28, 24) {real, imag} */,
  {32'h410a3239, 32'h3e7d9040} /* (19, 28, 23) {real, imag} */,
  {32'hc14eede9, 32'hc1a9288d} /* (19, 28, 22) {real, imag} */,
  {32'h4027d608, 32'h414b2d94} /* (19, 28, 21) {real, imag} */,
  {32'hbeef4860, 32'h412e486a} /* (19, 28, 20) {real, imag} */,
  {32'h41813513, 32'hc144d988} /* (19, 28, 19) {real, imag} */,
  {32'h402deb7a, 32'hc0980ec0} /* (19, 28, 18) {real, imag} */,
  {32'hbfc675b4, 32'hc031ded0} /* (19, 28, 17) {real, imag} */,
  {32'h40e0318e, 32'hc014ea70} /* (19, 28, 16) {real, imag} */,
  {32'hc10136d2, 32'hc0ddc850} /* (19, 28, 15) {real, imag} */,
  {32'h3f78c2aa, 32'h41a77ab1} /* (19, 28, 14) {real, imag} */,
  {32'h40e17ae1, 32'h40ab22a4} /* (19, 28, 13) {real, imag} */,
  {32'hc14aa7fb, 32'h40dc2734} /* (19, 28, 12) {real, imag} */,
  {32'h409208a4, 32'hc0be9ca8} /* (19, 28, 11) {real, imag} */,
  {32'h40e8644e, 32'h405d3178} /* (19, 28, 10) {real, imag} */,
  {32'h412d0ba7, 32'h41b6d01e} /* (19, 28, 9) {real, imag} */,
  {32'h4157aa8a, 32'h4141cbee} /* (19, 28, 8) {real, imag} */,
  {32'h413f485b, 32'h41572556} /* (19, 28, 7) {real, imag} */,
  {32'hc026f8bb, 32'hc1c57bcd} /* (19, 28, 6) {real, imag} */,
  {32'hc201d55f, 32'h42163c94} /* (19, 28, 5) {real, imag} */,
  {32'h42083a76, 32'h420e8068} /* (19, 28, 4) {real, imag} */,
  {32'h41c2211a, 32'hc126a045} /* (19, 28, 3) {real, imag} */,
  {32'hc1f49b78, 32'hc255440a} /* (19, 28, 2) {real, imag} */,
  {32'h4174b59a, 32'h42220750} /* (19, 28, 1) {real, imag} */,
  {32'h419f657a, 32'h426701c5} /* (19, 28, 0) {real, imag} */,
  {32'hc1ec5dd7, 32'hc2248796} /* (19, 27, 31) {real, imag} */,
  {32'h4075a1b8, 32'hc2623ce6} /* (19, 27, 30) {real, imag} */,
  {32'h429cd1a7, 32'hc104e18e} /* (19, 27, 29) {real, imag} */,
  {32'h4185a212, 32'hc0290000} /* (19, 27, 28) {real, imag} */,
  {32'h404b8b28, 32'hbcfd1980} /* (19, 27, 27) {real, imag} */,
  {32'h42bbe5cf, 32'hc01ff71e} /* (19, 27, 26) {real, imag} */,
  {32'hc287f624, 32'h421341d4} /* (19, 27, 25) {real, imag} */,
  {32'h4217798f, 32'h4172db4d} /* (19, 27, 24) {real, imag} */,
  {32'hc1a3d982, 32'hc04f2174} /* (19, 27, 23) {real, imag} */,
  {32'hc124df38, 32'h408427ec} /* (19, 27, 22) {real, imag} */,
  {32'hc209b9db, 32'h41614aff} /* (19, 27, 21) {real, imag} */,
  {32'hc13cfe16, 32'h415f8974} /* (19, 27, 20) {real, imag} */,
  {32'h406ae5c0, 32'h409d5957} /* (19, 27, 19) {real, imag} */,
  {32'h4157e6fa, 32'h3ef34fa0} /* (19, 27, 18) {real, imag} */,
  {32'h3fb611f0, 32'hc10215e4} /* (19, 27, 17) {real, imag} */,
  {32'h4148b368, 32'hc083a96c} /* (19, 27, 16) {real, imag} */,
  {32'hc0f99c6e, 32'hc0981550} /* (19, 27, 15) {real, imag} */,
  {32'hc041f356, 32'h40418884} /* (19, 27, 14) {real, imag} */,
  {32'hc1731474, 32'h408eb9ef} /* (19, 27, 13) {real, imag} */,
  {32'hc07efdae, 32'h41243f78} /* (19, 27, 12) {real, imag} */,
  {32'hc20b3fed, 32'hc19e0ca8} /* (19, 27, 11) {real, imag} */,
  {32'hc21cc9b6, 32'h41f8a5ab} /* (19, 27, 10) {real, imag} */,
  {32'h3f11f040, 32'hc115981b} /* (19, 27, 9) {real, imag} */,
  {32'hc1f107ca, 32'hc1cae5c2} /* (19, 27, 8) {real, imag} */,
  {32'hc1d126ce, 32'h41657302} /* (19, 27, 7) {real, imag} */,
  {32'h3fbd0fc0, 32'hc159487c} /* (19, 27, 6) {real, imag} */,
  {32'hc1973909, 32'hbfff2de6} /* (19, 27, 5) {real, imag} */,
  {32'hc1acccf4, 32'hc1e6b030} /* (19, 27, 4) {real, imag} */,
  {32'hc1913925, 32'h42137600} /* (19, 27, 3) {real, imag} */,
  {32'h42047a24, 32'h422dbefa} /* (19, 27, 2) {real, imag} */,
  {32'h40d9e8fc, 32'h4209b17a} /* (19, 27, 1) {real, imag} */,
  {32'h424c4466, 32'h416a7796} /* (19, 27, 0) {real, imag} */,
  {32'h40057f50, 32'h411b0356} /* (19, 26, 31) {real, imag} */,
  {32'h427ac746, 32'h4201504c} /* (19, 26, 30) {real, imag} */,
  {32'hc1f9dc89, 32'h40759120} /* (19, 26, 29) {real, imag} */,
  {32'hc1dc1b5a, 32'h410320b2} /* (19, 26, 28) {real, imag} */,
  {32'h42395c4e, 32'hc0c5e408} /* (19, 26, 27) {real, imag} */,
  {32'h41adaf09, 32'hc23ebde7} /* (19, 26, 26) {real, imag} */,
  {32'hc109175e, 32'hc1d90c89} /* (19, 26, 25) {real, imag} */,
  {32'hc1e5cdc2, 32'h415d07a8} /* (19, 26, 24) {real, imag} */,
  {32'h41a2cadc, 32'h4193c210} /* (19, 26, 23) {real, imag} */,
  {32'hc107a37d, 32'h419f9360} /* (19, 26, 22) {real, imag} */,
  {32'hc16a540d, 32'hc199b06a} /* (19, 26, 21) {real, imag} */,
  {32'h409e8226, 32'h40c8641f} /* (19, 26, 20) {real, imag} */,
  {32'h40f106e8, 32'hc08b59b4} /* (19, 26, 19) {real, imag} */,
  {32'h41424ef4, 32'hbf2d3f00} /* (19, 26, 18) {real, imag} */,
  {32'hc14be329, 32'h418f2043} /* (19, 26, 17) {real, imag} */,
  {32'hc081f41e, 32'hc011bb60} /* (19, 26, 16) {real, imag} */,
  {32'hc13154e7, 32'hbfd98830} /* (19, 26, 15) {real, imag} */,
  {32'h411e65dc, 32'h411adda8} /* (19, 26, 14) {real, imag} */,
  {32'h415a5868, 32'hc1e04feb} /* (19, 26, 13) {real, imag} */,
  {32'hbfc68d7a, 32'h3fb72d3c} /* (19, 26, 12) {real, imag} */,
  {32'h4097c7ee, 32'hc0a9d852} /* (19, 26, 11) {real, imag} */,
  {32'hc0f91946, 32'hbf3d7770} /* (19, 26, 10) {real, imag} */,
  {32'h41d53764, 32'h41d0bce6} /* (19, 26, 9) {real, imag} */,
  {32'hc207ae2b, 32'h428e892f} /* (19, 26, 8) {real, imag} */,
  {32'hc0c1f204, 32'hc19c52d1} /* (19, 26, 7) {real, imag} */,
  {32'hc1adf493, 32'h4221acd7} /* (19, 26, 6) {real, imag} */,
  {32'h4157b6b0, 32'h41fc5896} /* (19, 26, 5) {real, imag} */,
  {32'hc1607631, 32'hc2032814} /* (19, 26, 4) {real, imag} */,
  {32'h414aab26, 32'h41a349e8} /* (19, 26, 3) {real, imag} */,
  {32'hc1e6f911, 32'hc2410e0a} /* (19, 26, 2) {real, imag} */,
  {32'hc234c8af, 32'hc16052b6} /* (19, 26, 1) {real, imag} */,
  {32'h41c27510, 32'hc1c2dff2} /* (19, 26, 0) {real, imag} */,
  {32'h4220e64a, 32'hc17161c7} /* (19, 25, 31) {real, imag} */,
  {32'hc27356bd, 32'hc1a434b4} /* (19, 25, 30) {real, imag} */,
  {32'hc1392151, 32'hc0b7a262} /* (19, 25, 29) {real, imag} */,
  {32'h411e8c4e, 32'h40e0bfd2} /* (19, 25, 28) {real, imag} */,
  {32'hc071c658, 32'hc2296933} /* (19, 25, 27) {real, imag} */,
  {32'h41024e22, 32'hc182c681} /* (19, 25, 26) {real, imag} */,
  {32'h422c323e, 32'h42565212} /* (19, 25, 25) {real, imag} */,
  {32'hc045946c, 32'h41a1628e} /* (19, 25, 24) {real, imag} */,
  {32'hbf35b750, 32'hc22027aa} /* (19, 25, 23) {real, imag} */,
  {32'hc0b57fc3, 32'hc18a4268} /* (19, 25, 22) {real, imag} */,
  {32'hc1176bec, 32'h41a66a8e} /* (19, 25, 21) {real, imag} */,
  {32'h40dea38f, 32'hc0ef0732} /* (19, 25, 20) {real, imag} */,
  {32'h3f91e708, 32'hc026cf4b} /* (19, 25, 19) {real, imag} */,
  {32'h40431834, 32'h414741d1} /* (19, 25, 18) {real, imag} */,
  {32'h3fe30c78, 32'hc01ee70b} /* (19, 25, 17) {real, imag} */,
  {32'h41315920, 32'hc0da8302} /* (19, 25, 16) {real, imag} */,
  {32'hbf37f810, 32'h3dd831a0} /* (19, 25, 15) {real, imag} */,
  {32'h40e8be66, 32'h40aaa63a} /* (19, 25, 14) {real, imag} */,
  {32'hc18ba264, 32'h3f075904} /* (19, 25, 13) {real, imag} */,
  {32'hc14ebeb0, 32'hbfd33848} /* (19, 25, 12) {real, imag} */,
  {32'h41aa851e, 32'hc18323b6} /* (19, 25, 11) {real, imag} */,
  {32'h41134ff4, 32'h412323d9} /* (19, 25, 10) {real, imag} */,
  {32'hc0b48816, 32'h41548b2e} /* (19, 25, 9) {real, imag} */,
  {32'hbf990b00, 32'hc0e09a52} /* (19, 25, 8) {real, imag} */,
  {32'hc1bd481c, 32'hc115d4d2} /* (19, 25, 7) {real, imag} */,
  {32'hbe02c320, 32'h41ca53fb} /* (19, 25, 6) {real, imag} */,
  {32'hc1e33cd1, 32'h4170363d} /* (19, 25, 5) {real, imag} */,
  {32'h4128b17a, 32'h414bff33} /* (19, 25, 4) {real, imag} */,
  {32'hc14f44b7, 32'h3fba6f72} /* (19, 25, 3) {real, imag} */,
  {32'hc0ef9238, 32'h41ae0f1a} /* (19, 25, 2) {real, imag} */,
  {32'h41b32a9f, 32'h4186afa8} /* (19, 25, 1) {real, imag} */,
  {32'hc232e4eb, 32'h41954272} /* (19, 25, 0) {real, imag} */,
  {32'h40b35834, 32'h3f9c2d2c} /* (19, 24, 31) {real, imag} */,
  {32'h40707090, 32'h420818fc} /* (19, 24, 30) {real, imag} */,
  {32'hc24b45ee, 32'hc15c696a} /* (19, 24, 29) {real, imag} */,
  {32'hbdab9300, 32'hc20eeac7} /* (19, 24, 28) {real, imag} */,
  {32'hc1a06ec2, 32'hc1c2fb2d} /* (19, 24, 27) {real, imag} */,
  {32'hc187e65b, 32'h4143768d} /* (19, 24, 26) {real, imag} */,
  {32'hc0894af9, 32'h4015532c} /* (19, 24, 25) {real, imag} */,
  {32'h3f2a0380, 32'h4189098c} /* (19, 24, 24) {real, imag} */,
  {32'hc15600c7, 32'hc17b8f56} /* (19, 24, 23) {real, imag} */,
  {32'h41a2026f, 32'h41ca077f} /* (19, 24, 22) {real, imag} */,
  {32'hbffbc0e0, 32'h418b5c5e} /* (19, 24, 21) {real, imag} */,
  {32'h4009096e, 32'hc151304f} /* (19, 24, 20) {real, imag} */,
  {32'hc0cb6350, 32'hc139f41e} /* (19, 24, 19) {real, imag} */,
  {32'hc10d5a49, 32'h40c0141f} /* (19, 24, 18) {real, imag} */,
  {32'h4047c7aa, 32'hc0466802} /* (19, 24, 17) {real, imag} */,
  {32'h3d97c700, 32'hbde85880} /* (19, 24, 16) {real, imag} */,
  {32'hbfac5f14, 32'h40bebebf} /* (19, 24, 15) {real, imag} */,
  {32'h3fa67238, 32'hbfafffb4} /* (19, 24, 14) {real, imag} */,
  {32'hc0fc1608, 32'h414f0468} /* (19, 24, 13) {real, imag} */,
  {32'h3f1f4ca8, 32'hc14b9657} /* (19, 24, 12) {real, imag} */,
  {32'hc1b2c2f6, 32'hc0a095c1} /* (19, 24, 11) {real, imag} */,
  {32'h40e55844, 32'hc11869e2} /* (19, 24, 10) {real, imag} */,
  {32'h4097b20a, 32'h42002ca4} /* (19, 24, 9) {real, imag} */,
  {32'h40a6bff8, 32'h404df824} /* (19, 24, 8) {real, imag} */,
  {32'hc13c9e58, 32'hc113208d} /* (19, 24, 7) {real, imag} */,
  {32'h420c485e, 32'h4179e0c7} /* (19, 24, 6) {real, imag} */,
  {32'h4142eb2c, 32'hc0c5c2e4} /* (19, 24, 5) {real, imag} */,
  {32'h4202c5ae, 32'h41f0ce1e} /* (19, 24, 4) {real, imag} */,
  {32'h42387eda, 32'h421d1cc2} /* (19, 24, 3) {real, imag} */,
  {32'hc22e2a27, 32'hc1989e8c} /* (19, 24, 2) {real, imag} */,
  {32'h4207bcea, 32'h41119026} /* (19, 24, 1) {real, imag} */,
  {32'h422dc21e, 32'h41a2c810} /* (19, 24, 0) {real, imag} */,
  {32'h421da2d3, 32'h40c267f0} /* (19, 23, 31) {real, imag} */,
  {32'hc2150173, 32'h409ee512} /* (19, 23, 30) {real, imag} */,
  {32'hc1c7b2d0, 32'h419f6624} /* (19, 23, 29) {real, imag} */,
  {32'h40928ba7, 32'h413370b0} /* (19, 23, 28) {real, imag} */,
  {32'hc2143dba, 32'hc1d8aa5f} /* (19, 23, 27) {real, imag} */,
  {32'hc1c1fa8e, 32'hc157a0e9} /* (19, 23, 26) {real, imag} */,
  {32'hc12ab9a5, 32'hc0c8e394} /* (19, 23, 25) {real, imag} */,
  {32'h41c34b98, 32'hc11fcd90} /* (19, 23, 24) {real, imag} */,
  {32'h41ba4580, 32'h3f6fa340} /* (19, 23, 23) {real, imag} */,
  {32'hc18b8da8, 32'hbeed3500} /* (19, 23, 22) {real, imag} */,
  {32'h40663d4c, 32'h4020dc9d} /* (19, 23, 21) {real, imag} */,
  {32'hbe5d09a0, 32'h412a3881} /* (19, 23, 20) {real, imag} */,
  {32'hbf6d8270, 32'h3fc22218} /* (19, 23, 19) {real, imag} */,
  {32'hc0ba8c88, 32'h4085588e} /* (19, 23, 18) {real, imag} */,
  {32'h40a6913a, 32'hc0f6fd4c} /* (19, 23, 17) {real, imag} */,
  {32'h401d3258, 32'h40691d39} /* (19, 23, 16) {real, imag} */,
  {32'hbff75a48, 32'hc0ddca58} /* (19, 23, 15) {real, imag} */,
  {32'hc13189bc, 32'hbfb3a108} /* (19, 23, 14) {real, imag} */,
  {32'hc02540c4, 32'hc01ae544} /* (19, 23, 13) {real, imag} */,
  {32'h4062502e, 32'h41e01b78} /* (19, 23, 12) {real, imag} */,
  {32'h41c05970, 32'h40b90bc2} /* (19, 23, 11) {real, imag} */,
  {32'h412ce87b, 32'hc198151f} /* (19, 23, 10) {real, imag} */,
  {32'h41585ca5, 32'h41c5b182} /* (19, 23, 9) {real, imag} */,
  {32'h408e966a, 32'h420d68ad} /* (19, 23, 8) {real, imag} */,
  {32'hc10b7e93, 32'h41868553} /* (19, 23, 7) {real, imag} */,
  {32'hc2192375, 32'hc1a0aa10} /* (19, 23, 6) {real, imag} */,
  {32'h400d74e8, 32'hc1c97f7f} /* (19, 23, 5) {real, imag} */,
  {32'hc19d4591, 32'hc185f4d7} /* (19, 23, 4) {real, imag} */,
  {32'hc009894c, 32'hc28371b3} /* (19, 23, 3) {real, imag} */,
  {32'h40a895b0, 32'h41c78fca} /* (19, 23, 2) {real, imag} */,
  {32'hc1f750ce, 32'h425da62e} /* (19, 23, 1) {real, imag} */,
  {32'hc19e68d3, 32'hc07e415d} /* (19, 23, 0) {real, imag} */,
  {32'hc123f02d, 32'h412fe73e} /* (19, 22, 31) {real, imag} */,
  {32'hc196cc0a, 32'hc1aa3198} /* (19, 22, 30) {real, imag} */,
  {32'h418ebf4e, 32'h3ea80df0} /* (19, 22, 29) {real, imag} */,
  {32'hc154df42, 32'h4233fbe8} /* (19, 22, 28) {real, imag} */,
  {32'hc0581600, 32'hc2157ac9} /* (19, 22, 27) {real, imag} */,
  {32'hc0fe9a1a, 32'hc1f24f39} /* (19, 22, 26) {real, imag} */,
  {32'h415bc9ab, 32'h41138f1a} /* (19, 22, 25) {real, imag} */,
  {32'h415e0fe1, 32'hc10939fb} /* (19, 22, 24) {real, imag} */,
  {32'hc14d2470, 32'h414f3cdc} /* (19, 22, 23) {real, imag} */,
  {32'h3f7029fe, 32'h409bb313} /* (19, 22, 22) {real, imag} */,
  {32'h40e81ac8, 32'h3f06d1f0} /* (19, 22, 21) {real, imag} */,
  {32'hc176a5ef, 32'h4070e1f8} /* (19, 22, 20) {real, imag} */,
  {32'h413adecd, 32'h40bc8744} /* (19, 22, 19) {real, imag} */,
  {32'hc0ab75e1, 32'h3f29b760} /* (19, 22, 18) {real, imag} */,
  {32'hbfc267ce, 32'hbf9b371a} /* (19, 22, 17) {real, imag} */,
  {32'h40f08b42, 32'h400c4870} /* (19, 22, 16) {real, imag} */,
  {32'hbf856a8e, 32'h410375c7} /* (19, 22, 15) {real, imag} */,
  {32'hc025a91e, 32'hc0ead9f4} /* (19, 22, 14) {real, imag} */,
  {32'h40e456b6, 32'h412cb7de} /* (19, 22, 13) {real, imag} */,
  {32'h402428d4, 32'hc15ccd4e} /* (19, 22, 12) {real, imag} */,
  {32'h40ef7da8, 32'hc1b1da0c} /* (19, 22, 11) {real, imag} */,
  {32'hc093f0b2, 32'h416e126c} /* (19, 22, 10) {real, imag} */,
  {32'h40ac04eb, 32'h4164dda0} /* (19, 22, 9) {real, imag} */,
  {32'h4093eee6, 32'h41aa303a} /* (19, 22, 8) {real, imag} */,
  {32'h418834f8, 32'hc0dc0833} /* (19, 22, 7) {real, imag} */,
  {32'h3fdd6a80, 32'hc1310b16} /* (19, 22, 6) {real, imag} */,
  {32'h423a0954, 32'h40daafb6} /* (19, 22, 5) {real, imag} */,
  {32'hc25a3a1e, 32'h41a6eab5} /* (19, 22, 4) {real, imag} */,
  {32'hc1c39a52, 32'h40924f47} /* (19, 22, 3) {real, imag} */,
  {32'hc1e1bffa, 32'hbfef67d8} /* (19, 22, 2) {real, imag} */,
  {32'h41acbfe4, 32'hc1ae0a01} /* (19, 22, 1) {real, imag} */,
  {32'h419366d6, 32'h4227e895} /* (19, 22, 0) {real, imag} */,
  {32'hc032729a, 32'h41f96659} /* (19, 21, 31) {real, imag} */,
  {32'h411b1c5e, 32'hc1382028} /* (19, 21, 30) {real, imag} */,
  {32'h41dd4e01, 32'h41c4bc11} /* (19, 21, 29) {real, imag} */,
  {32'hc0a37a5d, 32'hc00cf604} /* (19, 21, 28) {real, imag} */,
  {32'hc222bad6, 32'hc104e3de} /* (19, 21, 27) {real, imag} */,
  {32'hc219a564, 32'hc061160e} /* (19, 21, 26) {real, imag} */,
  {32'h3ebdb1a0, 32'hc0ba5764} /* (19, 21, 25) {real, imag} */,
  {32'hc1253a74, 32'h419802e7} /* (19, 21, 24) {real, imag} */,
  {32'hc0de25ec, 32'hc16aca51} /* (19, 21, 23) {real, imag} */,
  {32'hbf8a263c, 32'hc0e5d056} /* (19, 21, 22) {real, imag} */,
  {32'h4126a134, 32'h4175b186} /* (19, 21, 21) {real, imag} */,
  {32'h4093422b, 32'hc1128cca} /* (19, 21, 20) {real, imag} */,
  {32'h40a47574, 32'hbf913852} /* (19, 21, 19) {real, imag} */,
  {32'h3fc80fae, 32'hbfc4b354} /* (19, 21, 18) {real, imag} */,
  {32'hc0270716, 32'h40318e90} /* (19, 21, 17) {real, imag} */,
  {32'hc03e89a2, 32'hbfec8550} /* (19, 21, 16) {real, imag} */,
  {32'h409e5417, 32'h408e6668} /* (19, 21, 15) {real, imag} */,
  {32'h40f0a58c, 32'hc03e44d2} /* (19, 21, 14) {real, imag} */,
  {32'h3eb10920, 32'hc088e4fe} /* (19, 21, 13) {real, imag} */,
  {32'h412dfa5e, 32'hbeb61340} /* (19, 21, 12) {real, imag} */,
  {32'hc128ed18, 32'h3f909514} /* (19, 21, 11) {real, imag} */,
  {32'hc1395956, 32'h40f4f024} /* (19, 21, 10) {real, imag} */,
  {32'hc202f5f8, 32'hc0058dd4} /* (19, 21, 9) {real, imag} */,
  {32'hc0cbd748, 32'hbfdacfb0} /* (19, 21, 8) {real, imag} */,
  {32'hc1700e97, 32'h41738ff2} /* (19, 21, 7) {real, imag} */,
  {32'h40b60d80, 32'hc0f03ef9} /* (19, 21, 6) {real, imag} */,
  {32'h4109224a, 32'hbe3301a0} /* (19, 21, 5) {real, imag} */,
  {32'h40cfd567, 32'h40a79e5e} /* (19, 21, 4) {real, imag} */,
  {32'hc103e2ba, 32'hc0d6ad1c} /* (19, 21, 3) {real, imag} */,
  {32'h40ee9fd4, 32'h411d29f0} /* (19, 21, 2) {real, imag} */,
  {32'h409f0fd5, 32'hc08bfdb4} /* (19, 21, 1) {real, imag} */,
  {32'hc0f3fbcf, 32'hc16363f6} /* (19, 21, 0) {real, imag} */,
  {32'h41c0b7b4, 32'hc157460a} /* (19, 20, 31) {real, imag} */,
  {32'h4172b416, 32'h40d43b08} /* (19, 20, 30) {real, imag} */,
  {32'h40363556, 32'h420de662} /* (19, 20, 29) {real, imag} */,
  {32'hc1f4f345, 32'hc0e8d0ea} /* (19, 20, 28) {real, imag} */,
  {32'hc10494e2, 32'hbfa24008} /* (19, 20, 27) {real, imag} */,
  {32'hc01fc4d8, 32'hc014201a} /* (19, 20, 26) {real, imag} */,
  {32'h410ba8e3, 32'hbfe3ff7e} /* (19, 20, 25) {real, imag} */,
  {32'hc01ee683, 32'h4132cf27} /* (19, 20, 24) {real, imag} */,
  {32'hbf82a688, 32'hbf743f14} /* (19, 20, 23) {real, imag} */,
  {32'hbfe17484, 32'hbfa88d90} /* (19, 20, 22) {real, imag} */,
  {32'h4133708d, 32'h40018e5d} /* (19, 20, 21) {real, imag} */,
  {32'h4120764c, 32'hc016e693} /* (19, 20, 20) {real, imag} */,
  {32'hc05d1c8e, 32'h40083e52} /* (19, 20, 19) {real, imag} */,
  {32'h402a6298, 32'hbea5c928} /* (19, 20, 18) {real, imag} */,
  {32'h40236c94, 32'h410b8017} /* (19, 20, 17) {real, imag} */,
  {32'hbf9c68d8, 32'hc015aaac} /* (19, 20, 16) {real, imag} */,
  {32'h4012c45c, 32'hc08c3272} /* (19, 20, 15) {real, imag} */,
  {32'hc0841f04, 32'hc044f69f} /* (19, 20, 14) {real, imag} */,
  {32'hbf600530, 32'h4093329b} /* (19, 20, 13) {real, imag} */,
  {32'h40850080, 32'hc015d1cf} /* (19, 20, 12) {real, imag} */,
  {32'h41177a23, 32'h40ff1e82} /* (19, 20, 11) {real, imag} */,
  {32'h41014fa8, 32'hbf60871d} /* (19, 20, 10) {real, imag} */,
  {32'h4110972d, 32'hbd247040} /* (19, 20, 9) {real, imag} */,
  {32'hc120ba73, 32'h3f20d3d0} /* (19, 20, 8) {real, imag} */,
  {32'h41e04284, 32'h3fbf22da} /* (19, 20, 7) {real, imag} */,
  {32'hc1b61c25, 32'hbfefc48c} /* (19, 20, 6) {real, imag} */,
  {32'h40f4923f, 32'hc179780b} /* (19, 20, 5) {real, imag} */,
  {32'h4102b212, 32'h40a73bb0} /* (19, 20, 4) {real, imag} */,
  {32'h3fd71368, 32'h40acca00} /* (19, 20, 3) {real, imag} */,
  {32'hc18c66e7, 32'hc112db28} /* (19, 20, 2) {real, imag} */,
  {32'h3f9ace30, 32'h408040a8} /* (19, 20, 1) {real, imag} */,
  {32'hc16ff401, 32'hc13c5549} /* (19, 20, 0) {real, imag} */,
  {32'h41721160, 32'hbf97ee98} /* (19, 19, 31) {real, imag} */,
  {32'h413c2710, 32'h41583910} /* (19, 19, 30) {real, imag} */,
  {32'h41055026, 32'hc0929ad6} /* (19, 19, 29) {real, imag} */,
  {32'h40196aa0, 32'h41329b4a} /* (19, 19, 28) {real, imag} */,
  {32'h41210367, 32'hc12ee57e} /* (19, 19, 27) {real, imag} */,
  {32'h41c4ef91, 32'h4163afba} /* (19, 19, 26) {real, imag} */,
  {32'h409fe9e5, 32'hc13c4f2f} /* (19, 19, 25) {real, imag} */,
  {32'hc16c4838, 32'h40d89a65} /* (19, 19, 24) {real, imag} */,
  {32'hc0f9004e, 32'h3eee5a30} /* (19, 19, 23) {real, imag} */,
  {32'h4086177e, 32'h3ff11634} /* (19, 19, 22) {real, imag} */,
  {32'hc0e80742, 32'h3f470d38} /* (19, 19, 21) {real, imag} */,
  {32'hbf59c450, 32'hc046247a} /* (19, 19, 20) {real, imag} */,
  {32'h4104abe8, 32'h3e622140} /* (19, 19, 19) {real, imag} */,
  {32'hc0397408, 32'h4085bd29} /* (19, 19, 18) {real, imag} */,
  {32'hc03cb85a, 32'hc08edfca} /* (19, 19, 17) {real, imag} */,
  {32'h402a059c, 32'h407b15e4} /* (19, 19, 16) {real, imag} */,
  {32'hbf5bb068, 32'h3ef8a198} /* (19, 19, 15) {real, imag} */,
  {32'hbfb63f90, 32'h3febe034} /* (19, 19, 14) {real, imag} */,
  {32'hc08081f0, 32'h402738f4} /* (19, 19, 13) {real, imag} */,
  {32'h4009b01a, 32'h40ab493b} /* (19, 19, 12) {real, imag} */,
  {32'hc07bc3b3, 32'hc0d4643d} /* (19, 19, 11) {real, imag} */,
  {32'hc094578e, 32'hc101aa38} /* (19, 19, 10) {real, imag} */,
  {32'hc1541fe1, 32'h40d5eddb} /* (19, 19, 9) {real, imag} */,
  {32'h414d2af6, 32'hc10c9770} /* (19, 19, 8) {real, imag} */,
  {32'hc0981b9b, 32'h41059745} /* (19, 19, 7) {real, imag} */,
  {32'h40a3032c, 32'hc18eb3c7} /* (19, 19, 6) {real, imag} */,
  {32'h3f463d50, 32'h41b4c5c5} /* (19, 19, 5) {real, imag} */,
  {32'hc1533598, 32'h41199086} /* (19, 19, 4) {real, imag} */,
  {32'hc1b92535, 32'h41b0d56e} /* (19, 19, 3) {real, imag} */,
  {32'h41ac6668, 32'hc011462a} /* (19, 19, 2) {real, imag} */,
  {32'hc17b4330, 32'hc154eb75} /* (19, 19, 1) {real, imag} */,
  {32'hc197f6b6, 32'h41419067} /* (19, 19, 0) {real, imag} */,
  {32'hbf1d6fe8, 32'hc1418462} /* (19, 18, 31) {real, imag} */,
  {32'hc0fdaf45, 32'hc00a07e8} /* (19, 18, 30) {real, imag} */,
  {32'h40b819af, 32'h40c23b7e} /* (19, 18, 29) {real, imag} */,
  {32'hc0f593bb, 32'h40b159e3} /* (19, 18, 28) {real, imag} */,
  {32'h40e1a588, 32'h400fdeb4} /* (19, 18, 27) {real, imag} */,
  {32'h403c23e4, 32'h40729ce8} /* (19, 18, 26) {real, imag} */,
  {32'h4062985b, 32'h40aa8c34} /* (19, 18, 25) {real, imag} */,
  {32'h410e9e99, 32'h410597c6} /* (19, 18, 24) {real, imag} */,
  {32'hc055b93e, 32'hc0333908} /* (19, 18, 23) {real, imag} */,
  {32'hc0c02ef2, 32'h4023a434} /* (19, 18, 22) {real, imag} */,
  {32'h40a665fc, 32'hc0788c22} /* (19, 18, 21) {real, imag} */,
  {32'h3f795d42, 32'h40447da3} /* (19, 18, 20) {real, imag} */,
  {32'hbec75210, 32'h409b70fa} /* (19, 18, 19) {real, imag} */,
  {32'h3f97ae24, 32'hc04b6db0} /* (19, 18, 18) {real, imag} */,
  {32'hbe626b20, 32'h3fb9c0cc} /* (19, 18, 17) {real, imag} */,
  {32'h3fcd232c, 32'hc0684b7c} /* (19, 18, 16) {real, imag} */,
  {32'h3f1ba428, 32'h3fcae7cc} /* (19, 18, 15) {real, imag} */,
  {32'hbe005720, 32'hbde80800} /* (19, 18, 14) {real, imag} */,
  {32'hc0af33a1, 32'h3fba75c6} /* (19, 18, 13) {real, imag} */,
  {32'h403a5d40, 32'h406e8529} /* (19, 18, 12) {real, imag} */,
  {32'h4073e389, 32'h40d67915} /* (19, 18, 11) {real, imag} */,
  {32'h409de2d2, 32'h3fc50e48} /* (19, 18, 10) {real, imag} */,
  {32'h4106cde4, 32'hc0bd5322} /* (19, 18, 9) {real, imag} */,
  {32'hbf508640, 32'hbfc9b544} /* (19, 18, 8) {real, imag} */,
  {32'hbe912c98, 32'h4106bcdd} /* (19, 18, 7) {real, imag} */,
  {32'hbf4dd812, 32'hc1338d5a} /* (19, 18, 6) {real, imag} */,
  {32'hc1045dbe, 32'h3eb04204} /* (19, 18, 5) {real, imag} */,
  {32'hc1077aa8, 32'h3ec00c30} /* (19, 18, 4) {real, imag} */,
  {32'h41760910, 32'hc12da377} /* (19, 18, 3) {real, imag} */,
  {32'h40e5aa01, 32'h4198cebd} /* (19, 18, 2) {real, imag} */,
  {32'hc17d7328, 32'hc01a4e42} /* (19, 18, 1) {real, imag} */,
  {32'h416df062, 32'h41628ac1} /* (19, 18, 0) {real, imag} */,
  {32'hc10462c1, 32'h40ccba71} /* (19, 17, 31) {real, imag} */,
  {32'hbf3e729a, 32'h4140ab01} /* (19, 17, 30) {real, imag} */,
  {32'hc1483a60, 32'hc15abdb5} /* (19, 17, 29) {real, imag} */,
  {32'h413910da, 32'hc0a54a84} /* (19, 17, 28) {real, imag} */,
  {32'h411ec0c6, 32'h40fff61d} /* (19, 17, 27) {real, imag} */,
  {32'hc0f49748, 32'hc0c7681f} /* (19, 17, 26) {real, imag} */,
  {32'hc1032b64, 32'h40faa994} /* (19, 17, 25) {real, imag} */,
  {32'h3f9ab80c, 32'hbeb4900c} /* (19, 17, 24) {real, imag} */,
  {32'hc1307f40, 32'h404e2e42} /* (19, 17, 23) {real, imag} */,
  {32'h40c3d2ac, 32'hc00013a6} /* (19, 17, 22) {real, imag} */,
  {32'h405ce304, 32'hc0f1ff0e} /* (19, 17, 21) {real, imag} */,
  {32'h401df50c, 32'hc01f3c67} /* (19, 17, 20) {real, imag} */,
  {32'hbf630566, 32'hc03d7e80} /* (19, 17, 19) {real, imag} */,
  {32'h401ec2bc, 32'h3fa0cb0a} /* (19, 17, 18) {real, imag} */,
  {32'hc00346e7, 32'h4093249f} /* (19, 17, 17) {real, imag} */,
  {32'h402d2668, 32'h3fbdcaee} /* (19, 17, 16) {real, imag} */,
  {32'h3f6720ec, 32'hc01d77b6} /* (19, 17, 15) {real, imag} */,
  {32'hbfcac988, 32'hbed295d8} /* (19, 17, 14) {real, imag} */,
  {32'h3f6aaf7a, 32'hc033e07e} /* (19, 17, 13) {real, imag} */,
  {32'hc09fd7be, 32'hc058d5b1} /* (19, 17, 12) {real, imag} */,
  {32'h4021fd26, 32'hc0431ef8} /* (19, 17, 11) {real, imag} */,
  {32'hc09483d8, 32'hbf4c3bba} /* (19, 17, 10) {real, imag} */,
  {32'hbda01b40, 32'hbebfcf70} /* (19, 17, 9) {real, imag} */,
  {32'h406e6f30, 32'hc0371244} /* (19, 17, 8) {real, imag} */,
  {32'hc01bb04e, 32'hc0aed174} /* (19, 17, 7) {real, imag} */,
  {32'hc05fbd9f, 32'h408b1ea9} /* (19, 17, 6) {real, imag} */,
  {32'h40cf9f04, 32'hc03c235a} /* (19, 17, 5) {real, imag} */,
  {32'h417657a2, 32'h3f668aa4} /* (19, 17, 4) {real, imag} */,
  {32'h40ce5c5b, 32'hc06ea5bc} /* (19, 17, 3) {real, imag} */,
  {32'h3f2858da, 32'h3f76c8b0} /* (19, 17, 2) {real, imag} */,
  {32'hc11c8087, 32'h40c90277} /* (19, 17, 1) {real, imag} */,
  {32'h4182e734, 32'h4041e529} /* (19, 17, 0) {real, imag} */,
  {32'hc102e189, 32'hc0812f98} /* (19, 16, 31) {real, imag} */,
  {32'h418bac76, 32'h414e8087} /* (19, 16, 30) {real, imag} */,
  {32'h3fd723b8, 32'h40c4aa54} /* (19, 16, 29) {real, imag} */,
  {32'hbfb2c3ca, 32'h4103745c} /* (19, 16, 28) {real, imag} */,
  {32'h3f099858, 32'h41371fee} /* (19, 16, 27) {real, imag} */,
  {32'h4074337e, 32'h410df8c8} /* (19, 16, 26) {real, imag} */,
  {32'hc05560d9, 32'hc128ee92} /* (19, 16, 25) {real, imag} */,
  {32'hbf9c1604, 32'hbfe2feac} /* (19, 16, 24) {real, imag} */,
  {32'h412128e4, 32'hc0923b5e} /* (19, 16, 23) {real, imag} */,
  {32'hbff05c12, 32'h40518cab} /* (19, 16, 22) {real, imag} */,
  {32'hbfa0858c, 32'h40bb141e} /* (19, 16, 21) {real, imag} */,
  {32'hc0b02c26, 32'hbe8275bf} /* (19, 16, 20) {real, imag} */,
  {32'hc059b4bd, 32'hbdc99020} /* (19, 16, 19) {real, imag} */,
  {32'hc0070190, 32'hbf7279ac} /* (19, 16, 18) {real, imag} */,
  {32'h3f8e36b4, 32'h3f89a508} /* (19, 16, 17) {real, imag} */,
  {32'hbf97bc84, 32'h4011f05d} /* (19, 16, 16) {real, imag} */,
  {32'hbe782aa4, 32'h3f8e5dee} /* (19, 16, 15) {real, imag} */,
  {32'hbc9db040, 32'hc0cdab9e} /* (19, 16, 14) {real, imag} */,
  {32'h408fecba, 32'hc003a035} /* (19, 16, 13) {real, imag} */,
  {32'h3f8a99fe, 32'hbf051b80} /* (19, 16, 12) {real, imag} */,
  {32'h40c32dc7, 32'h3ffe8d12} /* (19, 16, 11) {real, imag} */,
  {32'hc0a606aa, 32'h40f3c604} /* (19, 16, 10) {real, imag} */,
  {32'hc075d805, 32'hc13293c0} /* (19, 16, 9) {real, imag} */,
  {32'hc04f06f4, 32'h4081f48e} /* (19, 16, 8) {real, imag} */,
  {32'hc015e63d, 32'hc17183da} /* (19, 16, 7) {real, imag} */,
  {32'h40d0beb1, 32'hbf9d15f4} /* (19, 16, 6) {real, imag} */,
  {32'h412d7dbc, 32'hc1715b7a} /* (19, 16, 5) {real, imag} */,
  {32'h3e64cc2c, 32'hc1138462} /* (19, 16, 4) {real, imag} */,
  {32'hc117cb07, 32'hc08841b6} /* (19, 16, 3) {real, imag} */,
  {32'h4156a9e0, 32'hc174f1bd} /* (19, 16, 2) {real, imag} */,
  {32'h409d066c, 32'hbea67bdc} /* (19, 16, 1) {real, imag} */,
  {32'h40cb4200, 32'h41089d9b} /* (19, 16, 0) {real, imag} */,
  {32'hbfc30062, 32'hc1343a96} /* (19, 15, 31) {real, imag} */,
  {32'hbe8bc628, 32'hc047e738} /* (19, 15, 30) {real, imag} */,
  {32'hc19e6e1e, 32'hc090fe22} /* (19, 15, 29) {real, imag} */,
  {32'hc0deaea0, 32'h4105827a} /* (19, 15, 28) {real, imag} */,
  {32'hc05d67dc, 32'hbfff069c} /* (19, 15, 27) {real, imag} */,
  {32'hc0c0fa23, 32'h3fa31c72} /* (19, 15, 26) {real, imag} */,
  {32'h410efca0, 32'hc02cae40} /* (19, 15, 25) {real, imag} */,
  {32'h40295959, 32'hc0b8bab0} /* (19, 15, 24) {real, imag} */,
  {32'h401da048, 32'h403fab71} /* (19, 15, 23) {real, imag} */,
  {32'h408f1dcc, 32'h3e4a29a0} /* (19, 15, 22) {real, imag} */,
  {32'h4095c9e5, 32'h3e616180} /* (19, 15, 21) {real, imag} */,
  {32'h3f0a55a0, 32'h40326d9a} /* (19, 15, 20) {real, imag} */,
  {32'hbf47bef8, 32'h3d9e2b80} /* (19, 15, 19) {real, imag} */,
  {32'hbfecfd51, 32'h3cddbb80} /* (19, 15, 18) {real, imag} */,
  {32'hc0a1e142, 32'h3d8c7620} /* (19, 15, 17) {real, imag} */,
  {32'hbff44410, 32'hc0085937} /* (19, 15, 16) {real, imag} */,
  {32'h3f2e7d44, 32'hbed8d428} /* (19, 15, 15) {real, imag} */,
  {32'h4087b6a9, 32'hbe822828} /* (19, 15, 14) {real, imag} */,
  {32'h40424c3e, 32'h4054fd74} /* (19, 15, 13) {real, imag} */,
  {32'hc009595a, 32'h3f4908b6} /* (19, 15, 12) {real, imag} */,
  {32'h3fbdc914, 32'h3e57f040} /* (19, 15, 11) {real, imag} */,
  {32'h40572091, 32'h3e9fc2c0} /* (19, 15, 10) {real, imag} */,
  {32'hc02348e0, 32'hc0479b4f} /* (19, 15, 9) {real, imag} */,
  {32'h3f9908dc, 32'h40bb327c} /* (19, 15, 8) {real, imag} */,
  {32'hc0796500, 32'hc07ffe7e} /* (19, 15, 7) {real, imag} */,
  {32'hc08cded5, 32'h40632305} /* (19, 15, 6) {real, imag} */,
  {32'hbfa08068, 32'hc12135c4} /* (19, 15, 5) {real, imag} */,
  {32'h40fde070, 32'hc055c7de} /* (19, 15, 4) {real, imag} */,
  {32'h40720040, 32'hc1d79666} /* (19, 15, 3) {real, imag} */,
  {32'h40d6ecf6, 32'h415fe71a} /* (19, 15, 2) {real, imag} */,
  {32'hc0a7f25a, 32'hbfdafa50} /* (19, 15, 1) {real, imag} */,
  {32'h40ce3858, 32'h3fc8ec94} /* (19, 15, 0) {real, imag} */,
  {32'h3eb43400, 32'h408505e3} /* (19, 14, 31) {real, imag} */,
  {32'hc1ad5aef, 32'hc09513a9} /* (19, 14, 30) {real, imag} */,
  {32'hc18e2802, 32'hc17cb2a4} /* (19, 14, 29) {real, imag} */,
  {32'h413676cd, 32'hbf142164} /* (19, 14, 28) {real, imag} */,
  {32'h40d992d4, 32'h40ee6555} /* (19, 14, 27) {real, imag} */,
  {32'h3ff20de8, 32'hc145775c} /* (19, 14, 26) {real, imag} */,
  {32'hbf8189cc, 32'hc14e3dc9} /* (19, 14, 25) {real, imag} */,
  {32'hc0499692, 32'h411c92c0} /* (19, 14, 24) {real, imag} */,
  {32'hc0c899e2, 32'h40921df2} /* (19, 14, 23) {real, imag} */,
  {32'h4020feec, 32'hc1048eaf} /* (19, 14, 22) {real, imag} */,
  {32'hc11cf14c, 32'hc0d65785} /* (19, 14, 21) {real, imag} */,
  {32'hc06c08e8, 32'h404e7440} /* (19, 14, 20) {real, imag} */,
  {32'h3fac20fe, 32'h403631e0} /* (19, 14, 19) {real, imag} */,
  {32'hc08d1994, 32'h40620606} /* (19, 14, 18) {real, imag} */,
  {32'h3fb722b2, 32'hc01d8d03} /* (19, 14, 17) {real, imag} */,
  {32'h4051d35a, 32'hc084dfe5} /* (19, 14, 16) {real, imag} */,
  {32'h3f79a74c, 32'hbe31de70} /* (19, 14, 15) {real, imag} */,
  {32'hbec78e88, 32'h40206606} /* (19, 14, 14) {real, imag} */,
  {32'hc02eb493, 32'hc02bb7c6} /* (19, 14, 13) {real, imag} */,
  {32'hc0775afc, 32'h3febebec} /* (19, 14, 12) {real, imag} */,
  {32'h3ef021c0, 32'h3f996474} /* (19, 14, 11) {real, imag} */,
  {32'hc19cdcdc, 32'hc003850d} /* (19, 14, 10) {real, imag} */,
  {32'h4087d78c, 32'hc118d965} /* (19, 14, 9) {real, imag} */,
  {32'h412fd6da, 32'h412afc24} /* (19, 14, 8) {real, imag} */,
  {32'h414f3d98, 32'h41636891} /* (19, 14, 7) {real, imag} */,
  {32'h413b2851, 32'h401565a0} /* (19, 14, 6) {real, imag} */,
  {32'hc0c0b928, 32'h417a872c} /* (19, 14, 5) {real, imag} */,
  {32'h40138330, 32'hc0b0637a} /* (19, 14, 4) {real, imag} */,
  {32'hc15ac989, 32'h407b5c40} /* (19, 14, 3) {real, imag} */,
  {32'h406c1400, 32'h412a2e44} /* (19, 14, 2) {real, imag} */,
  {32'hbffd83d0, 32'h413a0548} /* (19, 14, 1) {real, imag} */,
  {32'hc036fb32, 32'h411be248} /* (19, 14, 0) {real, imag} */,
  {32'h40dbeb07, 32'h4187a0c7} /* (19, 13, 31) {real, imag} */,
  {32'h40ccdcc2, 32'hc0b2dd63} /* (19, 13, 30) {real, imag} */,
  {32'hc1c775e6, 32'h41068c06} /* (19, 13, 29) {real, imag} */,
  {32'hc189d566, 32'h40c584b0} /* (19, 13, 28) {real, imag} */,
  {32'hc07529ea, 32'h40061d12} /* (19, 13, 27) {real, imag} */,
  {32'h40106216, 32'h3f268318} /* (19, 13, 26) {real, imag} */,
  {32'h3fd9c450, 32'hc16d0c2c} /* (19, 13, 25) {real, imag} */,
  {32'hbff5973e, 32'h4140a702} /* (19, 13, 24) {real, imag} */,
  {32'h40b57194, 32'h40ba7b45} /* (19, 13, 23) {real, imag} */,
  {32'hbebcb63c, 32'h4104fc6e} /* (19, 13, 22) {real, imag} */,
  {32'h409932cd, 32'hc117bdc2} /* (19, 13, 21) {real, imag} */,
  {32'hc0246608, 32'hc04ef71a} /* (19, 13, 20) {real, imag} */,
  {32'hbe8245b0, 32'h40852f0c} /* (19, 13, 19) {real, imag} */,
  {32'hc09a9da8, 32'hbf694c76} /* (19, 13, 18) {real, imag} */,
  {32'hbf5a9330, 32'h3f182ddc} /* (19, 13, 17) {real, imag} */,
  {32'hbfe72e20, 32'hc011dac6} /* (19, 13, 16) {real, imag} */,
  {32'h40d4cdb2, 32'h3fd634aa} /* (19, 13, 15) {real, imag} */,
  {32'hc04e2214, 32'h4099c319} /* (19, 13, 14) {real, imag} */,
  {32'h3fc72b8c, 32'h3d12d600} /* (19, 13, 13) {real, imag} */,
  {32'hbf5b461e, 32'hbd42d600} /* (19, 13, 12) {real, imag} */,
  {32'hc0d81709, 32'hbea32930} /* (19, 13, 11) {real, imag} */,
  {32'hc029fcd0, 32'hc004999a} /* (19, 13, 10) {real, imag} */,
  {32'h3fefd0c2, 32'hc0e8e283} /* (19, 13, 9) {real, imag} */,
  {32'h406318b5, 32'h409332fc} /* (19, 13, 8) {real, imag} */,
  {32'hc1730c2e, 32'h40ea58ef} /* (19, 13, 7) {real, imag} */,
  {32'h411faae0, 32'hc0c93c5f} /* (19, 13, 6) {real, imag} */,
  {32'hc1925f72, 32'h41134244} /* (19, 13, 5) {real, imag} */,
  {32'h40c8a516, 32'h40654c37} /* (19, 13, 4) {real, imag} */,
  {32'h405f6c10, 32'hc0a3fe24} /* (19, 13, 3) {real, imag} */,
  {32'hbfc29b88, 32'h4021d7da} /* (19, 13, 2) {real, imag} */,
  {32'hbf8cc994, 32'h41401885} /* (19, 13, 1) {real, imag} */,
  {32'hc1255440, 32'h4144002e} /* (19, 13, 0) {real, imag} */,
  {32'hc1088ada, 32'h411893a9} /* (19, 12, 31) {real, imag} */,
  {32'hc0fe7b64, 32'hc1891c46} /* (19, 12, 30) {real, imag} */,
  {32'h41c51b12, 32'h3f78e550} /* (19, 12, 29) {real, imag} */,
  {32'hc08f0954, 32'hc0f7d29b} /* (19, 12, 28) {real, imag} */,
  {32'hc19e96f6, 32'h41177db2} /* (19, 12, 27) {real, imag} */,
  {32'h41cd5185, 32'hc04d01e3} /* (19, 12, 26) {real, imag} */,
  {32'hbfb78606, 32'hc0d47560} /* (19, 12, 25) {real, imag} */,
  {32'h41124bd7, 32'h40cf18ea} /* (19, 12, 24) {real, imag} */,
  {32'hc01c0221, 32'h40d28ad9} /* (19, 12, 23) {real, imag} */,
  {32'hc0d4c7f5, 32'hc0a0a159} /* (19, 12, 22) {real, imag} */,
  {32'hc0aac336, 32'hc1372391} /* (19, 12, 21) {real, imag} */,
  {32'h40aa235c, 32'hbf3b3442} /* (19, 12, 20) {real, imag} */,
  {32'h3f066580, 32'hc01ebf46} /* (19, 12, 19) {real, imag} */,
  {32'h4035be61, 32'h3fb413f4} /* (19, 12, 18) {real, imag} */,
  {32'h40836802, 32'h403da1f8} /* (19, 12, 17) {real, imag} */,
  {32'h4002f44f, 32'h3fd0f660} /* (19, 12, 16) {real, imag} */,
  {32'h3f9799cf, 32'h403a2dc0} /* (19, 12, 15) {real, imag} */,
  {32'hbed2d128, 32'hc0ab452d} /* (19, 12, 14) {real, imag} */,
  {32'h401d76e8, 32'h406c78b6} /* (19, 12, 13) {real, imag} */,
  {32'hbfd407e6, 32'h3f596cb2} /* (19, 12, 12) {real, imag} */,
  {32'hc04361a4, 32'hc0be89b2} /* (19, 12, 11) {real, imag} */,
  {32'h413ec38a, 32'h40acbb67} /* (19, 12, 10) {real, imag} */,
  {32'h40eac590, 32'hc0a0f92f} /* (19, 12, 9) {real, imag} */,
  {32'hc0a91dde, 32'hc073cf5b} /* (19, 12, 8) {real, imag} */,
  {32'h410a3b2b, 32'h41d3bf42} /* (19, 12, 7) {real, imag} */,
  {32'hc11b11ba, 32'hbe535ed0} /* (19, 12, 6) {real, imag} */,
  {32'h411382d1, 32'h3fd59aec} /* (19, 12, 5) {real, imag} */,
  {32'hc17f237a, 32'h3f9d7604} /* (19, 12, 4) {real, imag} */,
  {32'h418ccb86, 32'hc0e79158} /* (19, 12, 3) {real, imag} */,
  {32'hc162523a, 32'h40829f28} /* (19, 12, 2) {real, imag} */,
  {32'hc1295c3e, 32'h404e27f4} /* (19, 12, 1) {real, imag} */,
  {32'hc0cca9f0, 32'hc12e28d0} /* (19, 12, 0) {real, imag} */,
  {32'h3f2d49a7, 32'h40ac8fe1} /* (19, 11, 31) {real, imag} */,
  {32'h419d6848, 32'h401ee290} /* (19, 11, 30) {real, imag} */,
  {32'h412a9569, 32'hbf445ae0} /* (19, 11, 29) {real, imag} */,
  {32'h3ebfc180, 32'hc14ef28b} /* (19, 11, 28) {real, imag} */,
  {32'hc0c7d4cd, 32'hc115e6bd} /* (19, 11, 27) {real, imag} */,
  {32'h410cf8d2, 32'h4231f584} /* (19, 11, 26) {real, imag} */,
  {32'hc1a6f7ae, 32'hbf4b1fec} /* (19, 11, 25) {real, imag} */,
  {32'h4166db6a, 32'h4125b160} /* (19, 11, 24) {real, imag} */,
  {32'h4102064c, 32'h4141bf68} /* (19, 11, 23) {real, imag} */,
  {32'hc0519572, 32'hc09afa06} /* (19, 11, 22) {real, imag} */,
  {32'h401fac0a, 32'hc1708564} /* (19, 11, 21) {real, imag} */,
  {32'h40d6cf44, 32'hc011c6d3} /* (19, 11, 20) {real, imag} */,
  {32'h413534e0, 32'hbfc4acd8} /* (19, 11, 19) {real, imag} */,
  {32'hbf4ad5f0, 32'h4052e208} /* (19, 11, 18) {real, imag} */,
  {32'hc09a3e3f, 32'h40b15b2e} /* (19, 11, 17) {real, imag} */,
  {32'hbf7e7ed0, 32'hc03e1204} /* (19, 11, 16) {real, imag} */,
  {32'h3e6111a0, 32'h3f92638e} /* (19, 11, 15) {real, imag} */,
  {32'h3fc2a688, 32'hc0574c30} /* (19, 11, 14) {real, imag} */,
  {32'hc0f13644, 32'hbff13048} /* (19, 11, 13) {real, imag} */,
  {32'h3f6462f0, 32'h40ee046a} /* (19, 11, 12) {real, imag} */,
  {32'h41580d64, 32'h40b0520c} /* (19, 11, 11) {real, imag} */,
  {32'hc00e8d72, 32'h3fec0bd8} /* (19, 11, 10) {real, imag} */,
  {32'hbf304de0, 32'h3f1aff28} /* (19, 11, 9) {real, imag} */,
  {32'hc0cf6c55, 32'hc1526128} /* (19, 11, 8) {real, imag} */,
  {32'h41c539ae, 32'hbf3ee764} /* (19, 11, 7) {real, imag} */,
  {32'hc1909627, 32'hc0c24a14} /* (19, 11, 6) {real, imag} */,
  {32'hc08a81ab, 32'h41c7007e} /* (19, 11, 5) {real, imag} */,
  {32'h40867204, 32'h3e7e8b40} /* (19, 11, 4) {real, imag} */,
  {32'h42216c5a, 32'hc2214c5a} /* (19, 11, 3) {real, imag} */,
  {32'hc120af1d, 32'hc21fe89b} /* (19, 11, 2) {real, imag} */,
  {32'hbfa65a5a, 32'hc1188f4c} /* (19, 11, 1) {real, imag} */,
  {32'hc04dded4, 32'h3fc69a60} /* (19, 11, 0) {real, imag} */,
  {32'hc1d04290, 32'h41519d3d} /* (19, 10, 31) {real, imag} */,
  {32'hc18f9a6b, 32'h3f28b630} /* (19, 10, 30) {real, imag} */,
  {32'h419471b0, 32'h3f4fb8f0} /* (19, 10, 29) {real, imag} */,
  {32'h4166d43a, 32'h41907283} /* (19, 10, 28) {real, imag} */,
  {32'h41a79cfe, 32'hc1adcb2c} /* (19, 10, 27) {real, imag} */,
  {32'hc1f18157, 32'hc1b277ea} /* (19, 10, 26) {real, imag} */,
  {32'h40e2a103, 32'hc1829a6a} /* (19, 10, 25) {real, imag} */,
  {32'h4089f0e6, 32'hc0454ea0} /* (19, 10, 24) {real, imag} */,
  {32'h410df51a, 32'hbf6b7480} /* (19, 10, 23) {real, imag} */,
  {32'h410c5dba, 32'hbf9b87e8} /* (19, 10, 22) {real, imag} */,
  {32'hc12a6530, 32'hc11f46f6} /* (19, 10, 21) {real, imag} */,
  {32'h40300dda, 32'hc06a8b2c} /* (19, 10, 20) {real, imag} */,
  {32'hc0e2d437, 32'h3fb6f8b4} /* (19, 10, 19) {real, imag} */,
  {32'h4068b86a, 32'h410e6339} /* (19, 10, 18) {real, imag} */,
  {32'hc0efac7e, 32'h403b0971} /* (19, 10, 17) {real, imag} */,
  {32'hc002d5b8, 32'hbcfd0e00} /* (19, 10, 16) {real, imag} */,
  {32'hc001e863, 32'hbe65eaf0} /* (19, 10, 15) {real, imag} */,
  {32'h3f7eabd8, 32'hc16b22c5} /* (19, 10, 14) {real, imag} */,
  {32'h40d0b8bf, 32'hc0029782} /* (19, 10, 13) {real, imag} */,
  {32'h40098444, 32'hc1519425} /* (19, 10, 12) {real, imag} */,
  {32'hc1c03572, 32'hc01158bb} /* (19, 10, 11) {real, imag} */,
  {32'hc1925cd3, 32'h4121a3db} /* (19, 10, 10) {real, imag} */,
  {32'h4070155b, 32'h41aa69f2} /* (19, 10, 9) {real, imag} */,
  {32'h4192b98e, 32'h4074515c} /* (19, 10, 8) {real, imag} */,
  {32'hc15afe80, 32'h40afaaae} /* (19, 10, 7) {real, imag} */,
  {32'hc09c222c, 32'hc1040946} /* (19, 10, 6) {real, imag} */,
  {32'hc10bcc40, 32'hc11c1f30} /* (19, 10, 5) {real, imag} */,
  {32'h404e9450, 32'h4186ce0d} /* (19, 10, 4) {real, imag} */,
  {32'h41bcacce, 32'h419ca188} /* (19, 10, 3) {real, imag} */,
  {32'hc13d43b2, 32'h40d1feee} /* (19, 10, 2) {real, imag} */,
  {32'hc0fe1020, 32'hc1e02036} /* (19, 10, 1) {real, imag} */,
  {32'h41bf4c73, 32'h41cc3f1a} /* (19, 10, 0) {real, imag} */,
  {32'h41724138, 32'hc220bc8f} /* (19, 9, 31) {real, imag} */,
  {32'h421ff4f4, 32'h41ba4892} /* (19, 9, 30) {real, imag} */,
  {32'hc03c7dea, 32'h412f1272} /* (19, 9, 29) {real, imag} */,
  {32'h4008a14d, 32'hbee0d890} /* (19, 9, 28) {real, imag} */,
  {32'h41d1bad9, 32'hc167fcf0} /* (19, 9, 27) {real, imag} */,
  {32'hc1174f81, 32'h422793ea} /* (19, 9, 26) {real, imag} */,
  {32'h40fe0732, 32'hc177aa06} /* (19, 9, 25) {real, imag} */,
  {32'hc012945c, 32'hc1a11d9e} /* (19, 9, 24) {real, imag} */,
  {32'hc1798ba0, 32'h416f9882} /* (19, 9, 23) {real, imag} */,
  {32'hc06d8918, 32'h416a4dde} /* (19, 9, 22) {real, imag} */,
  {32'h4141b23d, 32'h41b25bf5} /* (19, 9, 21) {real, imag} */,
  {32'h3f6890c1, 32'h4048fd40} /* (19, 9, 20) {real, imag} */,
  {32'h419662e1, 32'hc0cbeebe} /* (19, 9, 19) {real, imag} */,
  {32'hc11df989, 32'hc181dcd4} /* (19, 9, 18) {real, imag} */,
  {32'hc112de78, 32'h3fa3b92c} /* (19, 9, 17) {real, imag} */,
  {32'hc0a6bce0, 32'h40b3473a} /* (19, 9, 16) {real, imag} */,
  {32'hc0c0574c, 32'h3fc10b14} /* (19, 9, 15) {real, imag} */,
  {32'h4096364a, 32'hc0065ebc} /* (19, 9, 14) {real, imag} */,
  {32'h401c7568, 32'hbcc87780} /* (19, 9, 13) {real, imag} */,
  {32'h3df5f4b8, 32'h415ab8f4} /* (19, 9, 12) {real, imag} */,
  {32'h40b10b9a, 32'hc047f3d0} /* (19, 9, 11) {real, imag} */,
  {32'h3ecf7ae0, 32'hbf643420} /* (19, 9, 10) {real, imag} */,
  {32'hc094fe44, 32'hc1a2cdc5} /* (19, 9, 9) {real, imag} */,
  {32'h41218131, 32'h4219ad1d} /* (19, 9, 8) {real, imag} */,
  {32'hc0e86f92, 32'h41039d6a} /* (19, 9, 7) {real, imag} */,
  {32'h40c732cc, 32'h4225db16} /* (19, 9, 6) {real, imag} */,
  {32'hc1b1d137, 32'hbf7fc9e0} /* (19, 9, 5) {real, imag} */,
  {32'h40d7d2de, 32'h4133faba} /* (19, 9, 4) {real, imag} */,
  {32'h4187cdd3, 32'hc01f8fbe} /* (19, 9, 3) {real, imag} */,
  {32'h40bd9524, 32'hc1f4d942} /* (19, 9, 2) {real, imag} */,
  {32'hc1ef9e28, 32'hc229d11f} /* (19, 9, 1) {real, imag} */,
  {32'hc0ed1c54, 32'hc1a16f7e} /* (19, 9, 0) {real, imag} */,
  {32'hc0e7e31a, 32'h42095833} /* (19, 8, 31) {real, imag} */,
  {32'h418831b0, 32'h41b35838} /* (19, 8, 30) {real, imag} */,
  {32'hc0816d28, 32'h408ff155} /* (19, 8, 29) {real, imag} */,
  {32'h41f752e3, 32'hc1fd0ef8} /* (19, 8, 28) {real, imag} */,
  {32'hc15725bf, 32'hc13cb3b4} /* (19, 8, 27) {real, imag} */,
  {32'h40d75c98, 32'hc1546172} /* (19, 8, 26) {real, imag} */,
  {32'hc12e6702, 32'h41c5cb34} /* (19, 8, 25) {real, imag} */,
  {32'h410fc706, 32'h419acb85} /* (19, 8, 24) {real, imag} */,
  {32'h4105d3de, 32'hc0976630} /* (19, 8, 23) {real, imag} */,
  {32'hc10705a8, 32'hc089fe47} /* (19, 8, 22) {real, imag} */,
  {32'h402c7f88, 32'hc0746874} /* (19, 8, 21) {real, imag} */,
  {32'hc08f4483, 32'hc0f065c7} /* (19, 8, 20) {real, imag} */,
  {32'h411c395c, 32'h41b10ee4} /* (19, 8, 19) {real, imag} */,
  {32'h3faebb80, 32'hc0c712d4} /* (19, 8, 18) {real, imag} */,
  {32'h404f9692, 32'hc07330b8} /* (19, 8, 17) {real, imag} */,
  {32'hbf0abff8, 32'hc0725a22} /* (19, 8, 16) {real, imag} */,
  {32'hc122716a, 32'hbf416100} /* (19, 8, 15) {real, imag} */,
  {32'h3fe2e970, 32'hc1542c46} /* (19, 8, 14) {real, imag} */,
  {32'hc0cb5119, 32'h40e660a8} /* (19, 8, 13) {real, imag} */,
  {32'hc10f8ab2, 32'h3f2c6838} /* (19, 8, 12) {real, imag} */,
  {32'h41966c9a, 32'h41680f85} /* (19, 8, 11) {real, imag} */,
  {32'h405255f2, 32'h4119a1cc} /* (19, 8, 10) {real, imag} */,
  {32'hc0e8f5c4, 32'h40b8b4b4} /* (19, 8, 9) {real, imag} */,
  {32'h4238235e, 32'h40900205} /* (19, 8, 8) {real, imag} */,
  {32'h40296a88, 32'h408a1e2c} /* (19, 8, 7) {real, imag} */,
  {32'hc194b5ac, 32'hc1c7d2f9} /* (19, 8, 6) {real, imag} */,
  {32'hbf83fc98, 32'h41d7abe6} /* (19, 8, 5) {real, imag} */,
  {32'hc086398c, 32'hc1670990} /* (19, 8, 4) {real, imag} */,
  {32'hc1a64ba6, 32'hc0c366f7} /* (19, 8, 3) {real, imag} */,
  {32'hc203b23c, 32'h41d73604} /* (19, 8, 2) {real, imag} */,
  {32'hc12d7d9b, 32'hbf5beb40} /* (19, 8, 1) {real, imag} */,
  {32'h410942d4, 32'h4132ce08} /* (19, 8, 0) {real, imag} */,
  {32'hc1b7af84, 32'hc12b557b} /* (19, 7, 31) {real, imag} */,
  {32'h4005a880, 32'hc26301fc} /* (19, 7, 30) {real, imag} */,
  {32'hc0aa03e4, 32'h426204cb} /* (19, 7, 29) {real, imag} */,
  {32'hbfd326e0, 32'h408c2a8c} /* (19, 7, 28) {real, imag} */,
  {32'hc1c2c6ba, 32'hc25de9e8} /* (19, 7, 27) {real, imag} */,
  {32'hc0a5cfe9, 32'h41a3abab} /* (19, 7, 26) {real, imag} */,
  {32'h421b3110, 32'h41d564f6} /* (19, 7, 25) {real, imag} */,
  {32'hc1ac6340, 32'h41948720} /* (19, 7, 24) {real, imag} */,
  {32'h3ee92300, 32'h40642e6e} /* (19, 7, 23) {real, imag} */,
  {32'h41fb719a, 32'hc0bc6344} /* (19, 7, 22) {real, imag} */,
  {32'h4152ca82, 32'hc1494436} /* (19, 7, 21) {real, imag} */,
  {32'h4045ded8, 32'hc15e1455} /* (19, 7, 20) {real, imag} */,
  {32'h40f0e5d4, 32'hc183688e} /* (19, 7, 19) {real, imag} */,
  {32'h40758eb0, 32'h40148cf8} /* (19, 7, 18) {real, imag} */,
  {32'hc0ac83d4, 32'hbfbe512f} /* (19, 7, 17) {real, imag} */,
  {32'h405fa8c6, 32'h405d4cbc} /* (19, 7, 16) {real, imag} */,
  {32'h4065ad90, 32'hbf0740c2} /* (19, 7, 15) {real, imag} */,
  {32'hc06487c0, 32'h40ebdae4} /* (19, 7, 14) {real, imag} */,
  {32'h40bf27a6, 32'hbff10a58} /* (19, 7, 13) {real, imag} */,
  {32'h4167ed78, 32'h417d0a83} /* (19, 7, 12) {real, imag} */,
  {32'h4072c2c8, 32'h41059e88} /* (19, 7, 11) {real, imag} */,
  {32'h4186fa6e, 32'hc0b73d2c} /* (19, 7, 10) {real, imag} */,
  {32'h41503856, 32'hc130307a} /* (19, 7, 9) {real, imag} */,
  {32'h403d913c, 32'hc09951ca} /* (19, 7, 8) {real, imag} */,
  {32'hc1d913db, 32'h40da6c58} /* (19, 7, 7) {real, imag} */,
  {32'hc151e5f6, 32'hc22f8f32} /* (19, 7, 6) {real, imag} */,
  {32'hc21b6246, 32'hc0441a80} /* (19, 7, 5) {real, imag} */,
  {32'h413e8c6c, 32'h41c64c8d} /* (19, 7, 4) {real, imag} */,
  {32'hc1b219a9, 32'hc0f8bb28} /* (19, 7, 3) {real, imag} */,
  {32'hc2a67b00, 32'h41a10a10} /* (19, 7, 2) {real, imag} */,
  {32'hc19e51e8, 32'hc129d61b} /* (19, 7, 1) {real, imag} */,
  {32'h4180cc83, 32'h4136bca5} /* (19, 7, 0) {real, imag} */,
  {32'h42636e3d, 32'hc26521cc} /* (19, 6, 31) {real, imag} */,
  {32'h4157d0be, 32'hc166d754} /* (19, 6, 30) {real, imag} */,
  {32'h421e2fb1, 32'hc1cddde2} /* (19, 6, 29) {real, imag} */,
  {32'hc1495c67, 32'h41a61684} /* (19, 6, 28) {real, imag} */,
  {32'h40c8b1f8, 32'h41136b5a} /* (19, 6, 27) {real, imag} */,
  {32'hc1b4eb07, 32'hc18bc687} /* (19, 6, 26) {real, imag} */,
  {32'h414a942e, 32'h420e62cb} /* (19, 6, 25) {real, imag} */,
  {32'h3f561558, 32'hc1fbc8e8} /* (19, 6, 24) {real, imag} */,
  {32'h4186e14f, 32'h4192b7ba} /* (19, 6, 23) {real, imag} */,
  {32'hc1cdb85d, 32'h40558f0a} /* (19, 6, 22) {real, imag} */,
  {32'h414335ce, 32'h40c7e742} /* (19, 6, 21) {real, imag} */,
  {32'h40b0e3c8, 32'hbf0c41a0} /* (19, 6, 20) {real, imag} */,
  {32'hc0bf06ac, 32'hc09d932e} /* (19, 6, 19) {real, imag} */,
  {32'h40b0d030, 32'h4119f39e} /* (19, 6, 18) {real, imag} */,
  {32'h4078f1e4, 32'h41401b3c} /* (19, 6, 17) {real, imag} */,
  {32'h4050dd28, 32'h414ddcd0} /* (19, 6, 16) {real, imag} */,
  {32'hc0cf3572, 32'hc11d7df8} /* (19, 6, 15) {real, imag} */,
  {32'hc1c73388, 32'h4169ff72} /* (19, 6, 14) {real, imag} */,
  {32'h4058ec67, 32'h40d19c5a} /* (19, 6, 13) {real, imag} */,
  {32'h4143e3c4, 32'h40ecd832} /* (19, 6, 12) {real, imag} */,
  {32'h41523b24, 32'h418ddf3e} /* (19, 6, 11) {real, imag} */,
  {32'hc0b1e8a4, 32'hc0b61073} /* (19, 6, 10) {real, imag} */,
  {32'hc21adefe, 32'hc19bf8d4} /* (19, 6, 9) {real, imag} */,
  {32'hc075b47e, 32'h414ddacd} /* (19, 6, 8) {real, imag} */,
  {32'hc222e1b6, 32'hc11765c1} /* (19, 6, 7) {real, imag} */,
  {32'hc215ea8e, 32'h40267f4a} /* (19, 6, 6) {real, imag} */,
  {32'h418e9e95, 32'hc1f68cff} /* (19, 6, 5) {real, imag} */,
  {32'h41ae122a, 32'hc100c694} /* (19, 6, 4) {real, imag} */,
  {32'hc1d172ca, 32'hc1e144d6} /* (19, 6, 3) {real, imag} */,
  {32'hc203f322, 32'hc1bb2a56} /* (19, 6, 2) {real, imag} */,
  {32'h4233a089, 32'hc27a79c4} /* (19, 6, 1) {real, imag} */,
  {32'h3f885270, 32'h422927f0} /* (19, 6, 0) {real, imag} */,
  {32'h41618fe5, 32'hc218e667} /* (19, 5, 31) {real, imag} */,
  {32'hc2050bee, 32'hc18b97d3} /* (19, 5, 30) {real, imag} */,
  {32'hc0cc5b40, 32'hc1878785} /* (19, 5, 29) {real, imag} */,
  {32'hbf4ffb00, 32'h42902283} /* (19, 5, 28) {real, imag} */,
  {32'hc22b4d18, 32'h41baef4a} /* (19, 5, 27) {real, imag} */,
  {32'h420c3d3d, 32'hc148df9a} /* (19, 5, 26) {real, imag} */,
  {32'hc1d09d97, 32'h40c5056c} /* (19, 5, 25) {real, imag} */,
  {32'hc1e738bf, 32'h41b41b4d} /* (19, 5, 24) {real, imag} */,
  {32'hc2075444, 32'h40f346ca} /* (19, 5, 23) {real, imag} */,
  {32'h3facefa0, 32'hc1e2d8c3} /* (19, 5, 22) {real, imag} */,
  {32'h41e446aa, 32'hbe334380} /* (19, 5, 21) {real, imag} */,
  {32'hc04c811e, 32'hc13b5bf7} /* (19, 5, 20) {real, imag} */,
  {32'hc0870a60, 32'hc05c7bb0} /* (19, 5, 19) {real, imag} */,
  {32'hc17a555e, 32'hc1a8d2e4} /* (19, 5, 18) {real, imag} */,
  {32'h40998be4, 32'hc18c3e8f} /* (19, 5, 17) {real, imag} */,
  {32'h40496dd8, 32'hc1152ad4} /* (19, 5, 16) {real, imag} */,
  {32'hc07ef2b8, 32'h40390fd8} /* (19, 5, 15) {real, imag} */,
  {32'hc164c26a, 32'h40870cb8} /* (19, 5, 14) {real, imag} */,
  {32'h402543b0, 32'h411e1ee6} /* (19, 5, 13) {real, imag} */,
  {32'h40526ede, 32'hc0f4b422} /* (19, 5, 12) {real, imag} */,
  {32'h4094ff70, 32'hc12ee958} /* (19, 5, 11) {real, imag} */,
  {32'h41ffa662, 32'hc14b497a} /* (19, 5, 10) {real, imag} */,
  {32'h41fe3029, 32'h3f6c68c0} /* (19, 5, 9) {real, imag} */,
  {32'hc259efc8, 32'h4145050e} /* (19, 5, 8) {real, imag} */,
  {32'hc23d0bb4, 32'h40235ea4} /* (19, 5, 7) {real, imag} */,
  {32'h40b19d38, 32'hc21fa36a} /* (19, 5, 6) {real, imag} */,
  {32'h42431334, 32'h4211f4c9} /* (19, 5, 5) {real, imag} */,
  {32'hc21ab6d2, 32'h418f4e54} /* (19, 5, 4) {real, imag} */,
  {32'h42557809, 32'hc1a0e9ef} /* (19, 5, 3) {real, imag} */,
  {32'h40c6cecc, 32'hbfc1ac70} /* (19, 5, 2) {real, imag} */,
  {32'h41562475, 32'h42651bad} /* (19, 5, 1) {real, imag} */,
  {32'hc22349c8, 32'h41db2dc6} /* (19, 5, 0) {real, imag} */,
  {32'h418233fa, 32'hc1db9452} /* (19, 4, 31) {real, imag} */,
  {32'hc29fcda6, 32'h4239402f} /* (19, 4, 30) {real, imag} */,
  {32'h3fb93468, 32'h41bcc8ea} /* (19, 4, 29) {real, imag} */,
  {32'h41b01521, 32'h404cfd84} /* (19, 4, 28) {real, imag} */,
  {32'h40324f56, 32'h3ffa7ed8} /* (19, 4, 27) {real, imag} */,
  {32'hc199210a, 32'h42219f7a} /* (19, 4, 26) {real, imag} */,
  {32'h425211bb, 32'hc1b78175} /* (19, 4, 25) {real, imag} */,
  {32'h41bc8c54, 32'hc20e1e16} /* (19, 4, 24) {real, imag} */,
  {32'hc1e0bf5c, 32'hc0e5970a} /* (19, 4, 23) {real, imag} */,
  {32'h41f24db4, 32'hc1d2ee66} /* (19, 4, 22) {real, imag} */,
  {32'h416dd658, 32'hc1860b3c} /* (19, 4, 21) {real, imag} */,
  {32'hc1faffb0, 32'h3f91c868} /* (19, 4, 20) {real, imag} */,
  {32'hc1bdd478, 32'h41904bbf} /* (19, 4, 19) {real, imag} */,
  {32'hc1037d2f, 32'h41997fa4} /* (19, 4, 18) {real, imag} */,
  {32'h40c40faa, 32'hc0d5ede6} /* (19, 4, 17) {real, imag} */,
  {32'h40b6ed1c, 32'h40cfb836} /* (19, 4, 16) {real, imag} */,
  {32'hc13967a5, 32'h4160c815} /* (19, 4, 15) {real, imag} */,
  {32'h411bfdc1, 32'h40e3a310} /* (19, 4, 14) {real, imag} */,
  {32'hbf83a448, 32'h41217ab4} /* (19, 4, 13) {real, imag} */,
  {32'hc1283424, 32'h41a5d4b2} /* (19, 4, 12) {real, imag} */,
  {32'hc1c0ed5e, 32'h41b8a550} /* (19, 4, 11) {real, imag} */,
  {32'h416ad018, 32'hc04a7228} /* (19, 4, 10) {real, imag} */,
  {32'hbf6a8d70, 32'hc1e1b676} /* (19, 4, 9) {real, imag} */,
  {32'h4105875b, 32'h4119e130} /* (19, 4, 8) {real, imag} */,
  {32'h406d2eb0, 32'h414f3666} /* (19, 4, 7) {real, imag} */,
  {32'hc1d0d1be, 32'hc1609ac7} /* (19, 4, 6) {real, imag} */,
  {32'hc181a909, 32'h418f66c0} /* (19, 4, 5) {real, imag} */,
  {32'h4166e09a, 32'hc20343c2} /* (19, 4, 4) {real, imag} */,
  {32'hc200536f, 32'h4202570b} /* (19, 4, 3) {real, imag} */,
  {32'h42118777, 32'hc2a80a86} /* (19, 4, 2) {real, imag} */,
  {32'hbf49d130, 32'h42a90e1a} /* (19, 4, 1) {real, imag} */,
  {32'hc2504e6a, 32'hc038f1bc} /* (19, 4, 0) {real, imag} */,
  {32'hbfcfbe80, 32'hc244a4bc} /* (19, 3, 31) {real, imag} */,
  {32'h4181fbee, 32'h426aa7a0} /* (19, 3, 30) {real, imag} */,
  {32'hc01f3a80, 32'hc26a2548} /* (19, 3, 29) {real, imag} */,
  {32'h40d67384, 32'hc23859fc} /* (19, 3, 28) {real, imag} */,
  {32'hc207326c, 32'h41982eb1} /* (19, 3, 27) {real, imag} */,
  {32'h414511b0, 32'h419b9abf} /* (19, 3, 26) {real, imag} */,
  {32'h41a014d5, 32'h41b29730} /* (19, 3, 25) {real, imag} */,
  {32'hc1b1cd64, 32'h411a33b4} /* (19, 3, 24) {real, imag} */,
  {32'h41051e08, 32'h415dec75} /* (19, 3, 23) {real, imag} */,
  {32'hc1c5bdb7, 32'h41cb977d} /* (19, 3, 22) {real, imag} */,
  {32'hc1e0f7c1, 32'h41a00bc0} /* (19, 3, 21) {real, imag} */,
  {32'h3f952c20, 32'hc12c8b1a} /* (19, 3, 20) {real, imag} */,
  {32'hc09aa6d3, 32'h41834fc5} /* (19, 3, 19) {real, imag} */,
  {32'hc0cda5de, 32'h41240ca6} /* (19, 3, 18) {real, imag} */,
  {32'hc0da2e52, 32'hc141efa8} /* (19, 3, 17) {real, imag} */,
  {32'hc13b332b, 32'hc15e914a} /* (19, 3, 16) {real, imag} */,
  {32'h3f01af90, 32'hc14c8338} /* (19, 3, 15) {real, imag} */,
  {32'hbfbfc618, 32'hc1bd75c1} /* (19, 3, 14) {real, imag} */,
  {32'h411b65aa, 32'h41bc544b} /* (19, 3, 13) {real, imag} */,
  {32'h41bba3a0, 32'hc1c26e7f} /* (19, 3, 12) {real, imag} */,
  {32'hc1bf9a07, 32'h40ab6b55} /* (19, 3, 11) {real, imag} */,
  {32'h41b294c9, 32'hc0a4803c} /* (19, 3, 10) {real, imag} */,
  {32'h4092bf56, 32'hc0a802ae} /* (19, 3, 9) {real, imag} */,
  {32'h420b1ea9, 32'h420aaf8b} /* (19, 3, 8) {real, imag} */,
  {32'hc163588a, 32'hc160436d} /* (19, 3, 7) {real, imag} */,
  {32'h42a57790, 32'hc18dde0d} /* (19, 3, 6) {real, imag} */,
  {32'h3fe1cf50, 32'h40e146e7} /* (19, 3, 5) {real, imag} */,
  {32'hc2307a30, 32'h42204b78} /* (19, 3, 4) {real, imag} */,
  {32'hc1f09cce, 32'h3f6989e0} /* (19, 3, 3) {real, imag} */,
  {32'hc2351a62, 32'h418b51f8} /* (19, 3, 2) {real, imag} */,
  {32'h422a0944, 32'hc1e78e64} /* (19, 3, 1) {real, imag} */,
  {32'h4113e865, 32'hc1d2ce63} /* (19, 3, 0) {real, imag} */,
  {32'h414b0825, 32'h41c0255a} /* (19, 2, 31) {real, imag} */,
  {32'h418b6715, 32'h42a4f534} /* (19, 2, 30) {real, imag} */,
  {32'h419376b6, 32'hc234a153} /* (19, 2, 29) {real, imag} */,
  {32'hc1a8ed1a, 32'hc219dcca} /* (19, 2, 28) {real, imag} */,
  {32'hc21c8a00, 32'hc211e4a9} /* (19, 2, 27) {real, imag} */,
  {32'hc28b9b98, 32'h409ec968} /* (19, 2, 26) {real, imag} */,
  {32'hc1b651fa, 32'h42792f49} /* (19, 2, 25) {real, imag} */,
  {32'h420910a9, 32'hc1f9a41a} /* (19, 2, 24) {real, imag} */,
  {32'hc172fb24, 32'hc2052936} /* (19, 2, 23) {real, imag} */,
  {32'h41f6df79, 32'hc023e720} /* (19, 2, 22) {real, imag} */,
  {32'h41ff2a66, 32'hc18e6562} /* (19, 2, 21) {real, imag} */,
  {32'hc09d6aee, 32'h412f4319} /* (19, 2, 20) {real, imag} */,
  {32'hc156fb6e, 32'h40f775f6} /* (19, 2, 19) {real, imag} */,
  {32'h3fe1f960, 32'hc03e5d18} /* (19, 2, 18) {real, imag} */,
  {32'h408792f6, 32'hbffe2c78} /* (19, 2, 17) {real, imag} */,
  {32'hc12d0de2, 32'hc1870bcc} /* (19, 2, 16) {real, imag} */,
  {32'h4091415e, 32'h4071345c} /* (19, 2, 15) {real, imag} */,
  {32'hc0fab378, 32'hc12b41be} /* (19, 2, 14) {real, imag} */,
  {32'h3ec43170, 32'hc1571e53} /* (19, 2, 13) {real, imag} */,
  {32'h41b9c572, 32'hc0ff76e6} /* (19, 2, 12) {real, imag} */,
  {32'hc0af60a8, 32'hc05bdfd2} /* (19, 2, 11) {real, imag} */,
  {32'h41dc41dd, 32'hc18f5b45} /* (19, 2, 10) {real, imag} */,
  {32'h4149466a, 32'h416e3762} /* (19, 2, 9) {real, imag} */,
  {32'hc06c0ab0, 32'hbfbf1a60} /* (19, 2, 8) {real, imag} */,
  {32'h403df698, 32'h421b541b} /* (19, 2, 7) {real, imag} */,
  {32'hc0fc6720, 32'hc2212537} /* (19, 2, 6) {real, imag} */,
  {32'h41807e2b, 32'hc00ec270} /* (19, 2, 5) {real, imag} */,
  {32'h4116ed59, 32'h41a09145} /* (19, 2, 4) {real, imag} */,
  {32'hc1d9ceca, 32'h3f4f58c0} /* (19, 2, 3) {real, imag} */,
  {32'h41ca372d, 32'hc20ccc22} /* (19, 2, 2) {real, imag} */,
  {32'hc1e32800, 32'h4253c18f} /* (19, 2, 1) {real, imag} */,
  {32'hc21d3e66, 32'h41900828} /* (19, 2, 0) {real, imag} */,
  {32'h418d7f79, 32'h41378f74} /* (19, 1, 31) {real, imag} */,
  {32'h42441bee, 32'h40e06380} /* (19, 1, 30) {real, imag} */,
  {32'hc27412fe, 32'hc202defc} /* (19, 1, 29) {real, imag} */,
  {32'h408541d0, 32'h418cebdf} /* (19, 1, 28) {real, imag} */,
  {32'h41d93ba4, 32'h428a4640} /* (19, 1, 27) {real, imag} */,
  {32'h417ab1de, 32'h428b91f6} /* (19, 1, 26) {real, imag} */,
  {32'hc1ba47fa, 32'hc084b456} /* (19, 1, 25) {real, imag} */,
  {32'hbfc14b38, 32'hc0d9daa6} /* (19, 1, 24) {real, imag} */,
  {32'hc0e56e6a, 32'hc252e547} /* (19, 1, 23) {real, imag} */,
  {32'h3f731a48, 32'hc2004812} /* (19, 1, 22) {real, imag} */,
  {32'hc18041ba, 32'h41912946} /* (19, 1, 21) {real, imag} */,
  {32'h4195d5f2, 32'h4195dc0c} /* (19, 1, 20) {real, imag} */,
  {32'hbea79680, 32'h40201e70} /* (19, 1, 19) {real, imag} */,
  {32'h3fb69ae8, 32'hc0d4d927} /* (19, 1, 18) {real, imag} */,
  {32'h41295e0a, 32'h4095d2b5} /* (19, 1, 17) {real, imag} */,
  {32'hbff6f1b8, 32'h40bf2f66} /* (19, 1, 16) {real, imag} */,
  {32'h40f4dce4, 32'hbfd96644} /* (19, 1, 15) {real, imag} */,
  {32'hbf08c870, 32'h4143df64} /* (19, 1, 14) {real, imag} */,
  {32'hc1a2a7c8, 32'hc11146e8} /* (19, 1, 13) {real, imag} */,
  {32'hc0d897a0, 32'hc16f81b4} /* (19, 1, 12) {real, imag} */,
  {32'h40df4191, 32'hc2303ee6} /* (19, 1, 11) {real, imag} */,
  {32'h4130fa24, 32'h41deaddd} /* (19, 1, 10) {real, imag} */,
  {32'hc1a3d024, 32'h417459ac} /* (19, 1, 9) {real, imag} */,
  {32'h42052297, 32'h41ddae50} /* (19, 1, 8) {real, imag} */,
  {32'hc1d9b5e4, 32'hc0b97626} /* (19, 1, 7) {real, imag} */,
  {32'h3f068258, 32'h41f26d51} /* (19, 1, 6) {real, imag} */,
  {32'hc2690222, 32'hc1b4fedd} /* (19, 1, 5) {real, imag} */,
  {32'h4259ef19, 32'h413432fa} /* (19, 1, 4) {real, imag} */,
  {32'hc14d14c6, 32'hc1cf42ce} /* (19, 1, 3) {real, imag} */,
  {32'hc1a0f614, 32'h403fce4d} /* (19, 1, 2) {real, imag} */,
  {32'hc101ef12, 32'h42090c5b} /* (19, 1, 1) {real, imag} */,
  {32'h419db050, 32'hc1890f24} /* (19, 1, 0) {real, imag} */,
  {32'h41a0cb7a, 32'h4298099b} /* (19, 0, 31) {real, imag} */,
  {32'hc0f27e74, 32'h420e2426} /* (19, 0, 30) {real, imag} */,
  {32'h422ad396, 32'h420c947d} /* (19, 0, 29) {real, imag} */,
  {32'h41daa25c, 32'h4269a50a} /* (19, 0, 28) {real, imag} */,
  {32'h400abfa0, 32'h41c68406} /* (19, 0, 27) {real, imag} */,
  {32'hc240ff91, 32'h41de28e8} /* (19, 0, 26) {real, imag} */,
  {32'hc14c5098, 32'hc1cf34be} /* (19, 0, 25) {real, imag} */,
  {32'hc1ba6ced, 32'hc075d840} /* (19, 0, 24) {real, imag} */,
  {32'h3f8f91a0, 32'h417b145b} /* (19, 0, 23) {real, imag} */,
  {32'hc1dcb7a0, 32'h418affcc} /* (19, 0, 22) {real, imag} */,
  {32'h4120acb0, 32'hc12bf725} /* (19, 0, 21) {real, imag} */,
  {32'h40b7e6b2, 32'h40988ff2} /* (19, 0, 20) {real, imag} */,
  {32'h40a048d4, 32'hc0830e4a} /* (19, 0, 19) {real, imag} */,
  {32'h3eaf2760, 32'hbf9197c4} /* (19, 0, 18) {real, imag} */,
  {32'hbff91998, 32'h4008c230} /* (19, 0, 17) {real, imag} */,
  {32'hc19ebea2, 32'hc19b8b0d} /* (19, 0, 16) {real, imag} */,
  {32'h4172ddad, 32'h40a14d70} /* (19, 0, 15) {real, imag} */,
  {32'h3ffce298, 32'hc0b8a8d9} /* (19, 0, 14) {real, imag} */,
  {32'hc18f230d, 32'hc10e4a17} /* (19, 0, 13) {real, imag} */,
  {32'hc182640a, 32'hc0972cc6} /* (19, 0, 12) {real, imag} */,
  {32'h423e5785, 32'h418d2ca8} /* (19, 0, 11) {real, imag} */,
  {32'hc183d93c, 32'hc216e713} /* (19, 0, 10) {real, imag} */,
  {32'h42510d8e, 32'h408dec56} /* (19, 0, 9) {real, imag} */,
  {32'hc20a6b1c, 32'hc2264f5f} /* (19, 0, 8) {real, imag} */,
  {32'hc1fc47ea, 32'h40b024c2} /* (19, 0, 7) {real, imag} */,
  {32'hc1c40cfa, 32'h41bafeca} /* (19, 0, 6) {real, imag} */,
  {32'hc1fd0802, 32'h40c36c1a} /* (19, 0, 5) {real, imag} */,
  {32'h41133f01, 32'hc25952aa} /* (19, 0, 4) {real, imag} */,
  {32'h411f4130, 32'h429c8ba0} /* (19, 0, 3) {real, imag} */,
  {32'h425006d0, 32'hc22b453e} /* (19, 0, 2) {real, imag} */,
  {32'hc244a753, 32'hc13c05e8} /* (19, 0, 1) {real, imag} */,
  {32'hc0d19e62, 32'h3f990f30} /* (19, 0, 0) {real, imag} */,
  {32'hc32b7951, 32'h429f7b0e} /* (18, 31, 31) {real, imag} */,
  {32'h42da18ac, 32'hc0c5013c} /* (18, 31, 30) {real, imag} */,
  {32'hc1339686, 32'hc154872b} /* (18, 31, 29) {real, imag} */,
  {32'hc1f99f92, 32'hc2502b8e} /* (18, 31, 28) {real, imag} */,
  {32'hc0b50de0, 32'hc0b53fd8} /* (18, 31, 27) {real, imag} */,
  {32'hc13195fc, 32'h41fdc886} /* (18, 31, 26) {real, imag} */,
  {32'h419175fa, 32'hbdc64880} /* (18, 31, 25) {real, imag} */,
  {32'hc102a49a, 32'h413c3d78} /* (18, 31, 24) {real, imag} */,
  {32'h4220e4ac, 32'hc0d088b6} /* (18, 31, 23) {real, imag} */,
  {32'h4154adc1, 32'hc2007656} /* (18, 31, 22) {real, imag} */,
  {32'h413f5fee, 32'h410cc58b} /* (18, 31, 21) {real, imag} */,
  {32'hbeaec420, 32'h40c78ee0} /* (18, 31, 20) {real, imag} */,
  {32'h4177ca02, 32'h40e9dd50} /* (18, 31, 19) {real, imag} */,
  {32'hc13840c8, 32'hc1428f44} /* (18, 31, 18) {real, imag} */,
  {32'hc1511036, 32'h41739426} /* (18, 31, 17) {real, imag} */,
  {32'h3eb90200, 32'h3f402c00} /* (18, 31, 16) {real, imag} */,
  {32'h3fefc2ac, 32'h41923a07} /* (18, 31, 15) {real, imag} */,
  {32'h40540f80, 32'h3f146198} /* (18, 31, 14) {real, imag} */,
  {32'h408d2308, 32'h40246eb8} /* (18, 31, 13) {real, imag} */,
  {32'hc15f4d9b, 32'h410c39c0} /* (18, 31, 12) {real, imag} */,
  {32'h4176d9b6, 32'hc1481a2f} /* (18, 31, 11) {real, imag} */,
  {32'h40f02dc6, 32'hc125e043} /* (18, 31, 10) {real, imag} */,
  {32'h413ccc13, 32'h41c2ca28} /* (18, 31, 9) {real, imag} */,
  {32'hc253fa28, 32'hc1feb2c0} /* (18, 31, 8) {real, imag} */,
  {32'h41b35e80, 32'hc1cffa1e} /* (18, 31, 7) {real, imag} */,
  {32'h4122a668, 32'h3f69aaf0} /* (18, 31, 6) {real, imag} */,
  {32'h42400a93, 32'h428e044c} /* (18, 31, 5) {real, imag} */,
  {32'hc1d93ad8, 32'h4223eac6} /* (18, 31, 4) {real, imag} */,
  {32'h41427370, 32'h420126ed} /* (18, 31, 3) {real, imag} */,
  {32'h42a94d2c, 32'h41f41075} /* (18, 31, 2) {real, imag} */,
  {32'hc2fca6ae, 32'hc2a6307a} /* (18, 31, 1) {real, imag} */,
  {32'hc2e06979, 32'hc156e893} /* (18, 31, 0) {real, imag} */,
  {32'h422c118c, 32'hc0aac367} /* (18, 30, 31) {real, imag} */,
  {32'hc1b249bc, 32'hc24bb07a} /* (18, 30, 30) {real, imag} */,
  {32'hbbbfa000, 32'hc2250fc0} /* (18, 30, 29) {real, imag} */,
  {32'h4184e2e4, 32'hc188640d} /* (18, 30, 28) {real, imag} */,
  {32'h4281f57b, 32'h421bea8d} /* (18, 30, 27) {real, imag} */,
  {32'h411f98c4, 32'h418796ba} /* (18, 30, 26) {real, imag} */,
  {32'h41ba03a7, 32'hbe857218} /* (18, 30, 25) {real, imag} */,
  {32'h418f62fe, 32'h3fe509e0} /* (18, 30, 24) {real, imag} */,
  {32'h41cae17b, 32'hc133e1d5} /* (18, 30, 23) {real, imag} */,
  {32'hc1de18da, 32'hc1426842} /* (18, 30, 22) {real, imag} */,
  {32'h41a4aaf2, 32'h41b9f1ed} /* (18, 30, 21) {real, imag} */,
  {32'hc1ce539f, 32'h4082370a} /* (18, 30, 20) {real, imag} */,
  {32'h402ef99a, 32'hc1cbacfc} /* (18, 30, 19) {real, imag} */,
  {32'hc12698b2, 32'h418c3c0a} /* (18, 30, 18) {real, imag} */,
  {32'h41355f66, 32'hc0e3ed7f} /* (18, 30, 17) {real, imag} */,
  {32'h4100e620, 32'h3f5cf280} /* (18, 30, 16) {real, imag} */,
  {32'h40bf4674, 32'h402b98de} /* (18, 30, 15) {real, imag} */,
  {32'hc0f7707c, 32'h418cc8a6} /* (18, 30, 14) {real, imag} */,
  {32'h4038e156, 32'h407d7ba4} /* (18, 30, 13) {real, imag} */,
  {32'hbfc85290, 32'h3eead898} /* (18, 30, 12) {real, imag} */,
  {32'hc1701998, 32'hc1987487} /* (18, 30, 11) {real, imag} */,
  {32'h41b0b3e0, 32'hbf836a4c} /* (18, 30, 10) {real, imag} */,
  {32'h3f0a7fa0, 32'hc145b349} /* (18, 30, 9) {real, imag} */,
  {32'hc1b18d9a, 32'hc263d807} /* (18, 30, 8) {real, imag} */,
  {32'hc1ce443f, 32'h40f5fd56} /* (18, 30, 7) {real, imag} */,
  {32'h422e3f50, 32'h40aa51e7} /* (18, 30, 6) {real, imag} */,
  {32'h4166e5e6, 32'hc22f26b3} /* (18, 30, 5) {real, imag} */,
  {32'h41a75b84, 32'h41b6230d} /* (18, 30, 4) {real, imag} */,
  {32'h419d49c4, 32'h42481238} /* (18, 30, 3) {real, imag} */,
  {32'hc305758c, 32'hc295ea05} /* (18, 30, 2) {real, imag} */,
  {32'h432ab3b5, 32'hc1a12e7a} /* (18, 30, 1) {real, imag} */,
  {32'h429b45a9, 32'hc196b0bf} /* (18, 30, 0) {real, imag} */,
  {32'hc1a01039, 32'h41d4b34f} /* (18, 29, 31) {real, imag} */,
  {32'hc07538ac, 32'h402c499b} /* (18, 29, 30) {real, imag} */,
  {32'h40115cd0, 32'h4203e9af} /* (18, 29, 29) {real, imag} */,
  {32'h424e69c4, 32'h41ccbb0c} /* (18, 29, 28) {real, imag} */,
  {32'h421c1090, 32'h4161ac36} /* (18, 29, 27) {real, imag} */,
  {32'h40dd5290, 32'hc14d6e0c} /* (18, 29, 26) {real, imag} */,
  {32'h411d4d69, 32'h417009e0} /* (18, 29, 25) {real, imag} */,
  {32'h4135d0af, 32'hbeb9c8c0} /* (18, 29, 24) {real, imag} */,
  {32'hc17e2874, 32'hc0e2e464} /* (18, 29, 23) {real, imag} */,
  {32'hbd2df5c0, 32'h41ae9cbe} /* (18, 29, 22) {real, imag} */,
  {32'hc127b534, 32'hc0751538} /* (18, 29, 21) {real, imag} */,
  {32'hc15d2b40, 32'hc1420f43} /* (18, 29, 20) {real, imag} */,
  {32'hc01e4bc8, 32'hc1556499} /* (18, 29, 19) {real, imag} */,
  {32'hc0fe5cbc, 32'h40319164} /* (18, 29, 18) {real, imag} */,
  {32'h41920f2c, 32'hc0d64475} /* (18, 29, 17) {real, imag} */,
  {32'h414d3a92, 32'hbf284478} /* (18, 29, 16) {real, imag} */,
  {32'hc130b5f7, 32'h40c7f59d} /* (18, 29, 15) {real, imag} */,
  {32'hc130f698, 32'hc14f65b7} /* (18, 29, 14) {real, imag} */,
  {32'h40b208b4, 32'h409d2976} /* (18, 29, 13) {real, imag} */,
  {32'hbf065840, 32'h410d2ee3} /* (18, 29, 12) {real, imag} */,
  {32'h41547a12, 32'h415b8e1a} /* (18, 29, 11) {real, imag} */,
  {32'hc0d8e278, 32'hc1338db8} /* (18, 29, 10) {real, imag} */,
  {32'h41c2ca56, 32'h41742748} /* (18, 29, 9) {real, imag} */,
  {32'h416d7425, 32'h4076959c} /* (18, 29, 8) {real, imag} */,
  {32'h40f38e36, 32'hc240a902} /* (18, 29, 7) {real, imag} */,
  {32'hbfe00630, 32'h41954ee0} /* (18, 29, 6) {real, imag} */,
  {32'hbd527600, 32'h4215d4e0} /* (18, 29, 5) {real, imag} */,
  {32'hc1868897, 32'h4135ea09} /* (18, 29, 4) {real, imag} */,
  {32'hc293c3d2, 32'hc2395aed} /* (18, 29, 3) {real, imag} */,
  {32'h41e4b1d6, 32'hc115307d} /* (18, 29, 2) {real, imag} */,
  {32'h4264313c, 32'h42338894} /* (18, 29, 1) {real, imag} */,
  {32'h41a1dd25, 32'h410fc854} /* (18, 29, 0) {real, imag} */,
  {32'hc2ccb1ee, 32'hc23c2b47} /* (18, 28, 31) {real, imag} */,
  {32'h41749a6e, 32'hc1539620} /* (18, 28, 30) {real, imag} */,
  {32'h4152bb66, 32'hc0ab2f98} /* (18, 28, 29) {real, imag} */,
  {32'h4095065a, 32'h40e0700b} /* (18, 28, 28) {real, imag} */,
  {32'h421045c0, 32'h41e4d5dd} /* (18, 28, 27) {real, imag} */,
  {32'hc1156b5b, 32'h3fc0c114} /* (18, 28, 26) {real, imag} */,
  {32'hc18dc2d4, 32'hc1a48b2e} /* (18, 28, 25) {real, imag} */,
  {32'h404718aa, 32'hc01021f2} /* (18, 28, 24) {real, imag} */,
  {32'hc114c6a7, 32'hc0020a30} /* (18, 28, 23) {real, imag} */,
  {32'h41b51b5e, 32'hc00010fc} /* (18, 28, 22) {real, imag} */,
  {32'hc1d93d9c, 32'h418cb16d} /* (18, 28, 21) {real, imag} */,
  {32'hc099b834, 32'hc13bd900} /* (18, 28, 20) {real, imag} */,
  {32'hc088ab9b, 32'hc11af58a} /* (18, 28, 19) {real, imag} */,
  {32'hc04bc92e, 32'hc0224948} /* (18, 28, 18) {real, imag} */,
  {32'h40e4d764, 32'h3f85d7a0} /* (18, 28, 17) {real, imag} */,
  {32'hbfe14e94, 32'h3f8d3dd0} /* (18, 28, 16) {real, imag} */,
  {32'hbf03b9a0, 32'hbf210c00} /* (18, 28, 15) {real, imag} */,
  {32'h40b8b3cf, 32'hc15237be} /* (18, 28, 14) {real, imag} */,
  {32'hc0dea28d, 32'hc19d7614} /* (18, 28, 13) {real, imag} */,
  {32'h41a9f6f7, 32'hc14e9474} /* (18, 28, 12) {real, imag} */,
  {32'hc0550290, 32'h40e3acb4} /* (18, 28, 11) {real, imag} */,
  {32'h3f521230, 32'hc1812abc} /* (18, 28, 10) {real, imag} */,
  {32'h412b2eb7, 32'h3eeb5a00} /* (18, 28, 9) {real, imag} */,
  {32'h418c37e0, 32'h415dc794} /* (18, 28, 8) {real, imag} */,
  {32'h4135c979, 32'h41886524} /* (18, 28, 7) {real, imag} */,
  {32'h414a3c75, 32'h3e1c2b20} /* (18, 28, 6) {real, imag} */,
  {32'hc17bdaba, 32'h41fdb769} /* (18, 28, 5) {real, imag} */,
  {32'h4035b848, 32'hc1149d9e} /* (18, 28, 4) {real, imag} */,
  {32'h41862c59, 32'h424a711b} /* (18, 28, 3) {real, imag} */,
  {32'h41a667bb, 32'h4212d76a} /* (18, 28, 2) {real, imag} */,
  {32'hc235c1bc, 32'h426b7f31} /* (18, 28, 1) {real, imag} */,
  {32'h4135d7b4, 32'h41c223d9} /* (18, 28, 0) {real, imag} */,
  {32'hc05f5464, 32'hc297fee4} /* (18, 27, 31) {real, imag} */,
  {32'hc12a2348, 32'h41276e1e} /* (18, 27, 30) {real, imag} */,
  {32'hbf39f4a8, 32'h41ae8874} /* (18, 27, 29) {real, imag} */,
  {32'h410a968e, 32'hc2213374} /* (18, 27, 28) {real, imag} */,
  {32'h421f2ad5, 32'hc1c3f95b} /* (18, 27, 27) {real, imag} */,
  {32'hc0b96dcb, 32'hc159a2a0} /* (18, 27, 26) {real, imag} */,
  {32'hc02ff38c, 32'h413e7d42} /* (18, 27, 25) {real, imag} */,
  {32'hc115bfdc, 32'hc197aca6} /* (18, 27, 24) {real, imag} */,
  {32'h41822f90, 32'h4237ca3c} /* (18, 27, 23) {real, imag} */,
  {32'hc0a950f6, 32'hc08f9d50} /* (18, 27, 22) {real, imag} */,
  {32'h413d7d1b, 32'h3fa2b864} /* (18, 27, 21) {real, imag} */,
  {32'h413cdec1, 32'hc0f062c0} /* (18, 27, 20) {real, imag} */,
  {32'h41019b88, 32'h40b2261a} /* (18, 27, 19) {real, imag} */,
  {32'h413975b4, 32'hc0d63b7a} /* (18, 27, 18) {real, imag} */,
  {32'hc0f91d98, 32'hc0bf8f8e} /* (18, 27, 17) {real, imag} */,
  {32'h4140f604, 32'hc111016c} /* (18, 27, 16) {real, imag} */,
  {32'hc1830dea, 32'h3e14eb40} /* (18, 27, 15) {real, imag} */,
  {32'hc13fa938, 32'hc1238731} /* (18, 27, 14) {real, imag} */,
  {32'h410bbe48, 32'hc104d81f} /* (18, 27, 13) {real, imag} */,
  {32'hc1404665, 32'hc0e1dcb8} /* (18, 27, 12) {real, imag} */,
  {32'hc16da5c3, 32'hbf9d030c} /* (18, 27, 11) {real, imag} */,
  {32'hc1b48aca, 32'h415b2828} /* (18, 27, 10) {real, imag} */,
  {32'h417ad287, 32'h4120bc02} /* (18, 27, 9) {real, imag} */,
  {32'hc182091e, 32'hc21194db} /* (18, 27, 8) {real, imag} */,
  {32'h41c129fa, 32'h419b3b07} /* (18, 27, 7) {real, imag} */,
  {32'hbfc2d3e4, 32'hc1b7da92} /* (18, 27, 6) {real, imag} */,
  {32'hc21244a9, 32'hc0ea2874} /* (18, 27, 5) {real, imag} */,
  {32'h422e80c8, 32'h412bfde2} /* (18, 27, 4) {real, imag} */,
  {32'hc16c8bb6, 32'hc1df3fb6} /* (18, 27, 3) {real, imag} */,
  {32'hc00daf26, 32'h4252ce48} /* (18, 27, 2) {real, imag} */,
  {32'hc17c054f, 32'h41923db0} /* (18, 27, 1) {real, imag} */,
  {32'h429d92f8, 32'hc2ab31da} /* (18, 27, 0) {real, imag} */,
  {32'h402fcb28, 32'h42065b4c} /* (18, 26, 31) {real, imag} */,
  {32'hc04f0968, 32'hc15ceeca} /* (18, 26, 30) {real, imag} */,
  {32'h41c74096, 32'hc1edce56} /* (18, 26, 29) {real, imag} */,
  {32'h41a95118, 32'h41c0659a} /* (18, 26, 28) {real, imag} */,
  {32'hc138d5ee, 32'h416969f5} /* (18, 26, 27) {real, imag} */,
  {32'h40e25b8e, 32'hc1f25d56} /* (18, 26, 26) {real, imag} */,
  {32'h4159c418, 32'h418cfb8d} /* (18, 26, 25) {real, imag} */,
  {32'hc14d6dc8, 32'h41af868f} /* (18, 26, 24) {real, imag} */,
  {32'hc22f6774, 32'hc1986b22} /* (18, 26, 23) {real, imag} */,
  {32'h3ff2a738, 32'hc12d5ba6} /* (18, 26, 22) {real, imag} */,
  {32'hc1667e62, 32'hc05efc74} /* (18, 26, 21) {real, imag} */,
  {32'hc0c939ab, 32'hc03ae772} /* (18, 26, 20) {real, imag} */,
  {32'h3faad948, 32'hc126cca0} /* (18, 26, 19) {real, imag} */,
  {32'hc08b1208, 32'h40c153fd} /* (18, 26, 18) {real, imag} */,
  {32'h40e95710, 32'hc1145d4a} /* (18, 26, 17) {real, imag} */,
  {32'hc0fedc6c, 32'h409ebc74} /* (18, 26, 16) {real, imag} */,
  {32'h40aa947c, 32'h3ffe50b2} /* (18, 26, 15) {real, imag} */,
  {32'hc0b6f3e0, 32'hc01dddf2} /* (18, 26, 14) {real, imag} */,
  {32'h40d8266a, 32'h40140ce8} /* (18, 26, 13) {real, imag} */,
  {32'h415b79b2, 32'h40527a62} /* (18, 26, 12) {real, imag} */,
  {32'h40250462, 32'hc1030e21} /* (18, 26, 11) {real, imag} */,
  {32'hc13a19b7, 32'h41b07863} /* (18, 26, 10) {real, imag} */,
  {32'h41875c58, 32'hc1852b96} /* (18, 26, 9) {real, imag} */,
  {32'hc07e78d8, 32'h3f22b120} /* (18, 26, 8) {real, imag} */,
  {32'hc1268a90, 32'h41e076e3} /* (18, 26, 7) {real, imag} */,
  {32'h41b689e6, 32'h40a2af40} /* (18, 26, 6) {real, imag} */,
  {32'h41243aa8, 32'hc2196b1b} /* (18, 26, 5) {real, imag} */,
  {32'h418b26ec, 32'hc12d31c7} /* (18, 26, 4) {real, imag} */,
  {32'hc27690f1, 32'h41dff7ae} /* (18, 26, 3) {real, imag} */,
  {32'h42283904, 32'hc1eabbbb} /* (18, 26, 2) {real, imag} */,
  {32'h4198770c, 32'hc1a8aae8} /* (18, 26, 1) {real, imag} */,
  {32'h42326254, 32'h41affb87} /* (18, 26, 0) {real, imag} */,
  {32'hc245538e, 32'h42007ea7} /* (18, 25, 31) {real, imag} */,
  {32'h41f9b7ef, 32'hc1c33774} /* (18, 25, 30) {real, imag} */,
  {32'h41ba8384, 32'hc1446da5} /* (18, 25, 29) {real, imag} */,
  {32'h4165da20, 32'hc279425e} /* (18, 25, 28) {real, imag} */,
  {32'h41a54073, 32'hc1831469} /* (18, 25, 27) {real, imag} */,
  {32'h4190c4ec, 32'hc1545875} /* (18, 25, 26) {real, imag} */,
  {32'hc0b09b9c, 32'h40d7d499} /* (18, 25, 25) {real, imag} */,
  {32'hc1603b78, 32'h421d8c69} /* (18, 25, 24) {real, imag} */,
  {32'hc1958e64, 32'h4036923a} /* (18, 25, 23) {real, imag} */,
  {32'h4197b982, 32'hc18d8eaa} /* (18, 25, 22) {real, imag} */,
  {32'hc098a76b, 32'h41c078b1} /* (18, 25, 21) {real, imag} */,
  {32'hc149c301, 32'hc10de97b} /* (18, 25, 20) {real, imag} */,
  {32'h41252d20, 32'hbe4186b0} /* (18, 25, 19) {real, imag} */,
  {32'hc1488a55, 32'h4045c41a} /* (18, 25, 18) {real, imag} */,
  {32'h4036de9c, 32'h40d9ccdc} /* (18, 25, 17) {real, imag} */,
  {32'hbf9cf140, 32'h40ddf545} /* (18, 25, 16) {real, imag} */,
  {32'h3fcb2a18, 32'hbf0d4c5c} /* (18, 25, 15) {real, imag} */,
  {32'h3e89ec60, 32'hc08c9dd3} /* (18, 25, 14) {real, imag} */,
  {32'hbfbc3a9c, 32'h3fd236f6} /* (18, 25, 13) {real, imag} */,
  {32'hc09c1102, 32'h404baa35} /* (18, 25, 12) {real, imag} */,
  {32'hbfbac11c, 32'h41848e6f} /* (18, 25, 11) {real, imag} */,
  {32'hc11ebf94, 32'h41a26062} /* (18, 25, 10) {real, imag} */,
  {32'hc0269d90, 32'hc10c85fc} /* (18, 25, 9) {real, imag} */,
  {32'h4126156c, 32'h418c1546} /* (18, 25, 8) {real, imag} */,
  {32'hc1e99501, 32'hc160abd2} /* (18, 25, 7) {real, imag} */,
  {32'h416dee50, 32'hc20cad43} /* (18, 25, 6) {real, imag} */,
  {32'hc1b416a1, 32'hc1c76963} /* (18, 25, 5) {real, imag} */,
  {32'h421e3124, 32'h4266278c} /* (18, 25, 4) {real, imag} */,
  {32'h4177edac, 32'hc176dd4b} /* (18, 25, 3) {real, imag} */,
  {32'hc230008a, 32'h41939bb4} /* (18, 25, 2) {real, imag} */,
  {32'h41abdf84, 32'h415d3e7c} /* (18, 25, 1) {real, imag} */,
  {32'hc1b81300, 32'h4130d0dc} /* (18, 25, 0) {real, imag} */,
  {32'h41da3a56, 32'h3f15be80} /* (18, 24, 31) {real, imag} */,
  {32'h41747096, 32'hc01ce8f9} /* (18, 24, 30) {real, imag} */,
  {32'hc0867848, 32'h416fb314} /* (18, 24, 29) {real, imag} */,
  {32'hc177f7da, 32'h41926c68} /* (18, 24, 28) {real, imag} */,
  {32'hc03f1490, 32'h41908372} /* (18, 24, 27) {real, imag} */,
  {32'hc1cdc9d3, 32'h41ae9da4} /* (18, 24, 26) {real, imag} */,
  {32'hc0ab610e, 32'hc0602480} /* (18, 24, 25) {real, imag} */,
  {32'hc1e12805, 32'hc0b383ff} /* (18, 24, 24) {real, imag} */,
  {32'hc13c84d2, 32'h41c6f341} /* (18, 24, 23) {real, imag} */,
  {32'h409aa03a, 32'h3ff59f68} /* (18, 24, 22) {real, imag} */,
  {32'hc1c2829b, 32'h402797b1} /* (18, 24, 21) {real, imag} */,
  {32'hc0916d8d, 32'h40dea326} /* (18, 24, 20) {real, imag} */,
  {32'hbf785718, 32'hc110a4be} /* (18, 24, 19) {real, imag} */,
  {32'hbfa20c1c, 32'hc0e11300} /* (18, 24, 18) {real, imag} */,
  {32'hc02da076, 32'h40871ae4} /* (18, 24, 17) {real, imag} */,
  {32'hc11c8314, 32'hbf148448} /* (18, 24, 16) {real, imag} */,
  {32'hbf81eab4, 32'h400dafa0} /* (18, 24, 15) {real, imag} */,
  {32'h410f9926, 32'hbe1a74e0} /* (18, 24, 14) {real, imag} */,
  {32'hc0ec0927, 32'hc10b6b6e} /* (18, 24, 13) {real, imag} */,
  {32'h411fb21c, 32'h412421bd} /* (18, 24, 12) {real, imag} */,
  {32'hc023f4a8, 32'h4015ee17} /* (18, 24, 11) {real, imag} */,
  {32'hc1431d4d, 32'h415cd6a5} /* (18, 24, 10) {real, imag} */,
  {32'hc11d0398, 32'h41a90171} /* (18, 24, 9) {real, imag} */,
  {32'h40842854, 32'hc18ef6d4} /* (18, 24, 8) {real, imag} */,
  {32'h4185c5cc, 32'h41a2d598} /* (18, 24, 7) {real, imag} */,
  {32'h41bacaed, 32'hbf026810} /* (18, 24, 6) {real, imag} */,
  {32'h402fd98c, 32'h41a87052} /* (18, 24, 5) {real, imag} */,
  {32'hbfe01cbc, 32'hc1c904c4} /* (18, 24, 4) {real, imag} */,
  {32'hbee233c8, 32'h41d98284} /* (18, 24, 3) {real, imag} */,
  {32'hc108b960, 32'hc10d5ef0} /* (18, 24, 2) {real, imag} */,
  {32'h42273cb1, 32'hc239affc} /* (18, 24, 1) {real, imag} */,
  {32'hc025899c, 32'hc0207912} /* (18, 24, 0) {real, imag} */,
  {32'hc134b197, 32'h41a93116} /* (18, 23, 31) {real, imag} */,
  {32'hc0a37e9a, 32'h3fe0a9b0} /* (18, 23, 30) {real, imag} */,
  {32'hc1a57691, 32'hc0112448} /* (18, 23, 29) {real, imag} */,
  {32'hc19dd99e, 32'hc193e862} /* (18, 23, 28) {real, imag} */,
  {32'h41775cd0, 32'hc0293c8e} /* (18, 23, 27) {real, imag} */,
  {32'hc148e5ac, 32'hbe9f63e0} /* (18, 23, 26) {real, imag} */,
  {32'h40b5be4b, 32'h41196729} /* (18, 23, 25) {real, imag} */,
  {32'h3f9826f4, 32'hc181961c} /* (18, 23, 24) {real, imag} */,
  {32'hc154c1d2, 32'h40cfa950} /* (18, 23, 23) {real, imag} */,
  {32'h41522dfa, 32'h40a49b6a} /* (18, 23, 22) {real, imag} */,
  {32'hbf4c2508, 32'hc1789bfc} /* (18, 23, 21) {real, imag} */,
  {32'hc024e228, 32'hc14ed96e} /* (18, 23, 20) {real, imag} */,
  {32'hc11460c4, 32'h40ec1e93} /* (18, 23, 19) {real, imag} */,
  {32'h40ae4b9f, 32'hc0f49f06} /* (18, 23, 18) {real, imag} */,
  {32'hbf312930, 32'h410a078a} /* (18, 23, 17) {real, imag} */,
  {32'h40e67b37, 32'h40d8aa65} /* (18, 23, 16) {real, imag} */,
  {32'hc0e004d2, 32'hbf72cb78} /* (18, 23, 15) {real, imag} */,
  {32'hbfa069f4, 32'h405a3ae4} /* (18, 23, 14) {real, imag} */,
  {32'h403446fe, 32'h40ce2263} /* (18, 23, 13) {real, imag} */,
  {32'hc07d7e08, 32'hc101989c} /* (18, 23, 12) {real, imag} */,
  {32'hc109e0f0, 32'hc03dd1ce} /* (18, 23, 11) {real, imag} */,
  {32'h4188eb49, 32'h4132685d} /* (18, 23, 10) {real, imag} */,
  {32'h4101eb7a, 32'hbf83ce6e} /* (18, 23, 9) {real, imag} */,
  {32'hbfefd034, 32'h412298ec} /* (18, 23, 8) {real, imag} */,
  {32'h40c6e94f, 32'h3ffa68a8} /* (18, 23, 7) {real, imag} */,
  {32'h41806a20, 32'h41246a27} /* (18, 23, 6) {real, imag} */,
  {32'hc21ebaac, 32'hc188b142} /* (18, 23, 5) {real, imag} */,
  {32'hc2570671, 32'h41bef99e} /* (18, 23, 4) {real, imag} */,
  {32'hc144a272, 32'hc21050b0} /* (18, 23, 3) {real, imag} */,
  {32'h41ae7d6a, 32'h414cc1e2} /* (18, 23, 2) {real, imag} */,
  {32'h41e5095c, 32'h41669d9c} /* (18, 23, 1) {real, imag} */,
  {32'h415f3a98, 32'h41919c7d} /* (18, 23, 0) {real, imag} */,
  {32'hc1cc04cb, 32'hc20d763a} /* (18, 22, 31) {real, imag} */,
  {32'hc1c30b1d, 32'h3e247400} /* (18, 22, 30) {real, imag} */,
  {32'hbc215a00, 32'hc0dbdd30} /* (18, 22, 29) {real, imag} */,
  {32'h40128cca, 32'h41b789e6} /* (18, 22, 28) {real, imag} */,
  {32'h40aad1f7, 32'hc08beb28} /* (18, 22, 27) {real, imag} */,
  {32'h415f4c78, 32'h40f95896} /* (18, 22, 26) {real, imag} */,
  {32'h41860416, 32'hc08b90b8} /* (18, 22, 25) {real, imag} */,
  {32'hc12870bb, 32'h4094654b} /* (18, 22, 24) {real, imag} */,
  {32'h3f9caf3e, 32'h4017db09} /* (18, 22, 23) {real, imag} */,
  {32'h41a44774, 32'hc0454328} /* (18, 22, 22) {real, imag} */,
  {32'h40d0a715, 32'hc05da29e} /* (18, 22, 21) {real, imag} */,
  {32'h3f344fb8, 32'h40b75336} /* (18, 22, 20) {real, imag} */,
  {32'hc0c95651, 32'h418b209e} /* (18, 22, 19) {real, imag} */,
  {32'hc0d37ac8, 32'hc10e90bc} /* (18, 22, 18) {real, imag} */,
  {32'h401aaad2, 32'h4088e9c1} /* (18, 22, 17) {real, imag} */,
  {32'hc11df1ae, 32'h3fd5019f} /* (18, 22, 16) {real, imag} */,
  {32'hc10ff578, 32'hc085459f} /* (18, 22, 15) {real, imag} */,
  {32'hbee706f8, 32'h40c9cdfe} /* (18, 22, 14) {real, imag} */,
  {32'h412d76dc, 32'h409ddd86} /* (18, 22, 13) {real, imag} */,
  {32'h4023a0a5, 32'hc0b28afc} /* (18, 22, 12) {real, imag} */,
  {32'hbf27f5f8, 32'h41186854} /* (18, 22, 11) {real, imag} */,
  {32'hc129f330, 32'h417ff76e} /* (18, 22, 10) {real, imag} */,
  {32'hc044606b, 32'h4042e71f} /* (18, 22, 9) {real, imag} */,
  {32'hbfe9b918, 32'hbe77bda0} /* (18, 22, 8) {real, imag} */,
  {32'h40022c64, 32'hbfd39e92} /* (18, 22, 7) {real, imag} */,
  {32'h4228dd18, 32'hc097c1c2} /* (18, 22, 6) {real, imag} */,
  {32'h3d67e180, 32'hc1011433} /* (18, 22, 5) {real, imag} */,
  {32'hc0ed9091, 32'hc0f022cf} /* (18, 22, 4) {real, imag} */,
  {32'hc133e438, 32'h3e59f490} /* (18, 22, 3) {real, imag} */,
  {32'h41f198c1, 32'hc18db334} /* (18, 22, 2) {real, imag} */,
  {32'hc0ffc66c, 32'h41883e31} /* (18, 22, 1) {real, imag} */,
  {32'h41e4cd87, 32'h3fcd6373} /* (18, 22, 0) {real, imag} */,
  {32'h3f3aac38, 32'h3ea28180} /* (18, 21, 31) {real, imag} */,
  {32'hc14dd2f4, 32'h41f71732} /* (18, 21, 30) {real, imag} */,
  {32'hbfc5d460, 32'h419b1398} /* (18, 21, 29) {real, imag} */,
  {32'hc13d5404, 32'h41b43420} /* (18, 21, 28) {real, imag} */,
  {32'hc1294e60, 32'h3fd1bca8} /* (18, 21, 27) {real, imag} */,
  {32'h4199fce8, 32'hc033246b} /* (18, 21, 26) {real, imag} */,
  {32'h4124338a, 32'hc08fb6a6} /* (18, 21, 25) {real, imag} */,
  {32'h414e68f6, 32'hc16b2bc0} /* (18, 21, 24) {real, imag} */,
  {32'hbfd5f52e, 32'hc083bb6c} /* (18, 21, 23) {real, imag} */,
  {32'hbf282970, 32'h3ff6ee9e} /* (18, 21, 22) {real, imag} */,
  {32'h417dd46a, 32'h406a289c} /* (18, 21, 21) {real, imag} */,
  {32'h400d2524, 32'hc0075b59} /* (18, 21, 20) {real, imag} */,
  {32'h407d82b8, 32'h4102a9b0} /* (18, 21, 19) {real, imag} */,
  {32'h40286519, 32'h40936177} /* (18, 21, 18) {real, imag} */,
  {32'hc080ea2e, 32'h4047ca95} /* (18, 21, 17) {real, imag} */,
  {32'hc0ab0e25, 32'hc100e6d4} /* (18, 21, 16) {real, imag} */,
  {32'hbffd2e81, 32'h411c835d} /* (18, 21, 15) {real, imag} */,
  {32'h401413fb, 32'hc0c1b1eb} /* (18, 21, 14) {real, imag} */,
  {32'hc00018a0, 32'hc13b1fe2} /* (18, 21, 13) {real, imag} */,
  {32'h401c9e74, 32'hc0f99d44} /* (18, 21, 12) {real, imag} */,
  {32'h40a3507c, 32'h40cebb12} /* (18, 21, 11) {real, imag} */,
  {32'h403d9b4c, 32'h3fd74b42} /* (18, 21, 10) {real, imag} */,
  {32'hbf2a2404, 32'h410c9954} /* (18, 21, 9) {real, imag} */,
  {32'h401f8142, 32'hc1439bd2} /* (18, 21, 8) {real, imag} */,
  {32'hc096a2a3, 32'hc136f8ef} /* (18, 21, 7) {real, imag} */,
  {32'hc1083f68, 32'h40a4bd30} /* (18, 21, 6) {real, imag} */,
  {32'h40f54c61, 32'hc1bb6ce6} /* (18, 21, 5) {real, imag} */,
  {32'h40477a2a, 32'h415677cf} /* (18, 21, 4) {real, imag} */,
  {32'h41aacc23, 32'hc113787d} /* (18, 21, 3) {real, imag} */,
  {32'hc015005a, 32'h40f32458} /* (18, 21, 2) {real, imag} */,
  {32'hc0f3c933, 32'hc113c4a6} /* (18, 21, 1) {real, imag} */,
  {32'hbf3a3d48, 32'hc14fb3aa} /* (18, 21, 0) {real, imag} */,
  {32'h410ab55c, 32'h4165a37a} /* (18, 20, 31) {real, imag} */,
  {32'hc004776c, 32'h414b7f29} /* (18, 20, 30) {real, imag} */,
  {32'h407e7344, 32'h404d8388} /* (18, 20, 29) {real, imag} */,
  {32'h4172722c, 32'hbf7230e0} /* (18, 20, 28) {real, imag} */,
  {32'hc18280fd, 32'hbf43a98a} /* (18, 20, 27) {real, imag} */,
  {32'h3f8382c8, 32'h4105af0c} /* (18, 20, 26) {real, imag} */,
  {32'h40fab21c, 32'h411da2a8} /* (18, 20, 25) {real, imag} */,
  {32'hc1a57d30, 32'h40b9ce95} /* (18, 20, 24) {real, imag} */,
  {32'hc094d7f8, 32'hbf41dd50} /* (18, 20, 23) {real, imag} */,
  {32'h41817ebc, 32'h404d691f} /* (18, 20, 22) {real, imag} */,
  {32'hc09b5367, 32'hc0e9a71f} /* (18, 20, 21) {real, imag} */,
  {32'h3fe853f8, 32'hc00635fa} /* (18, 20, 20) {real, imag} */,
  {32'hc03cd214, 32'h3eff9b38} /* (18, 20, 19) {real, imag} */,
  {32'hc02bba72, 32'h41256598} /* (18, 20, 18) {real, imag} */,
  {32'hc0b029cb, 32'hc070e2c8} /* (18, 20, 17) {real, imag} */,
  {32'hbdfe4460, 32'hc07f2a90} /* (18, 20, 16) {real, imag} */,
  {32'hbeee5b30, 32'hbef4f47c} /* (18, 20, 15) {real, imag} */,
  {32'h3fb0b168, 32'h3f1a3c60} /* (18, 20, 14) {real, imag} */,
  {32'hbffa26e8, 32'h3f82e13a} /* (18, 20, 13) {real, imag} */,
  {32'hc0e2416a, 32'hc06dbbd6} /* (18, 20, 12) {real, imag} */,
  {32'h401581b2, 32'h40a85071} /* (18, 20, 11) {real, imag} */,
  {32'h40505ebc, 32'h41100f3c} /* (18, 20, 10) {real, imag} */,
  {32'h40a378bc, 32'hc12ab7ea} /* (18, 20, 9) {real, imag} */,
  {32'h40431194, 32'hc0adc25b} /* (18, 20, 8) {real, imag} */,
  {32'h40e49d74, 32'h3e5d5940} /* (18, 20, 7) {real, imag} */,
  {32'hc0fbd38e, 32'hc1459bc8} /* (18, 20, 6) {real, imag} */,
  {32'h418db6ff, 32'hbfef8f11} /* (18, 20, 5) {real, imag} */,
  {32'h412f7218, 32'hc202c070} /* (18, 20, 4) {real, imag} */,
  {32'hc1fc7274, 32'h4121a4b5} /* (18, 20, 3) {real, imag} */,
  {32'hc14b7425, 32'h3fa6ff48} /* (18, 20, 2) {real, imag} */,
  {32'hc1105b9c, 32'h4131431a} /* (18, 20, 1) {real, imag} */,
  {32'hc003c2f5, 32'h41f8b1ba} /* (18, 20, 0) {real, imag} */,
  {32'h408eb0c5, 32'h3f0b40a0} /* (18, 19, 31) {real, imag} */,
  {32'hc032e400, 32'hc1960721} /* (18, 19, 30) {real, imag} */,
  {32'hc0d9cba6, 32'hc118f551} /* (18, 19, 29) {real, imag} */,
  {32'hbe8477aa, 32'hc0c276df} /* (18, 19, 28) {real, imag} */,
  {32'h4120ef3e, 32'h410721d5} /* (18, 19, 27) {real, imag} */,
  {32'hc124c599, 32'h4070c758} /* (18, 19, 26) {real, imag} */,
  {32'hc16febc5, 32'h3fe319b0} /* (18, 19, 25) {real, imag} */,
  {32'hc1049abd, 32'h408f004a} /* (18, 19, 24) {real, imag} */,
  {32'hbf9ee380, 32'hc14be64c} /* (18, 19, 23) {real, imag} */,
  {32'hc09e60b8, 32'h3f4cd2e8} /* (18, 19, 22) {real, imag} */,
  {32'h3fcd45a0, 32'h4072f9d6} /* (18, 19, 21) {real, imag} */,
  {32'h410bc418, 32'h3f9e4bee} /* (18, 19, 20) {real, imag} */,
  {32'h40984c93, 32'h40d20ab1} /* (18, 19, 19) {real, imag} */,
  {32'hc019e1be, 32'hbfb991f4} /* (18, 19, 18) {real, imag} */,
  {32'h40638951, 32'hbf885ccf} /* (18, 19, 17) {real, imag} */,
  {32'hbf885740, 32'h3f0a5638} /* (18, 19, 16) {real, imag} */,
  {32'hbff19e46, 32'hc0900ede} /* (18, 19, 15) {real, imag} */,
  {32'h3f164890, 32'hbfbd45fc} /* (18, 19, 14) {real, imag} */,
  {32'h3e81d470, 32'h3f94ac60} /* (18, 19, 13) {real, imag} */,
  {32'h40bfa732, 32'h40921384} /* (18, 19, 12) {real, imag} */,
  {32'hc0bfb6f6, 32'hc0530a0e} /* (18, 19, 11) {real, imag} */,
  {32'h414487c8, 32'h40bb2421} /* (18, 19, 10) {real, imag} */,
  {32'hbfd394e8, 32'hc1875cde} /* (18, 19, 9) {real, imag} */,
  {32'hc137d929, 32'hbed3ba20} /* (18, 19, 8) {real, imag} */,
  {32'h41197dd3, 32'h40f556bc} /* (18, 19, 7) {real, imag} */,
  {32'hc0e3966a, 32'h4151f7fe} /* (18, 19, 6) {real, imag} */,
  {32'h40c2fe8c, 32'hc065a048} /* (18, 19, 5) {real, imag} */,
  {32'h3f6464c5, 32'h4117a7c4} /* (18, 19, 4) {real, imag} */,
  {32'hc07459bf, 32'h3f47af50} /* (18, 19, 3) {real, imag} */,
  {32'h4160d038, 32'hc17586ce} /* (18, 19, 2) {real, imag} */,
  {32'h40bf97d7, 32'h3f2a9a00} /* (18, 19, 1) {real, imag} */,
  {32'hc1ed5bc9, 32'h4110658a} /* (18, 19, 0) {real, imag} */,
  {32'h40d15b78, 32'h40952510} /* (18, 18, 31) {real, imag} */,
  {32'h40b36650, 32'hc0038fa6} /* (18, 18, 30) {real, imag} */,
  {32'hc0e6927c, 32'h4118af02} /* (18, 18, 29) {real, imag} */,
  {32'hc0b080b4, 32'hc13c73eb} /* (18, 18, 28) {real, imag} */,
  {32'h4061ff9c, 32'h40cba264} /* (18, 18, 27) {real, imag} */,
  {32'h41795701, 32'hc0b0ef26} /* (18, 18, 26) {real, imag} */,
  {32'hc058c722, 32'h4098595e} /* (18, 18, 25) {real, imag} */,
  {32'hc1285392, 32'hc0412636} /* (18, 18, 24) {real, imag} */,
  {32'h3f592a20, 32'hc1598930} /* (18, 18, 23) {real, imag} */,
  {32'h3f25068c, 32'hbfd57b2c} /* (18, 18, 22) {real, imag} */,
  {32'h40b22edb, 32'h40872b84} /* (18, 18, 21) {real, imag} */,
  {32'h3f9c3acb, 32'h401f7900} /* (18, 18, 20) {real, imag} */,
  {32'h401a4a78, 32'h40b93e09} /* (18, 18, 19) {real, imag} */,
  {32'hbeee2b74, 32'h402bfbf9} /* (18, 18, 18) {real, imag} */,
  {32'h3ee681fc, 32'h3f8299f8} /* (18, 18, 17) {real, imag} */,
  {32'hbf90226a, 32'h4054a43e} /* (18, 18, 16) {real, imag} */,
  {32'h3fa4d937, 32'hbfe526e8} /* (18, 18, 15) {real, imag} */,
  {32'h4044f9d4, 32'hbfc1cac6} /* (18, 18, 14) {real, imag} */,
  {32'h3e8cc4d0, 32'hbfc5a16c} /* (18, 18, 13) {real, imag} */,
  {32'hbfac07cd, 32'h408dc24d} /* (18, 18, 12) {real, imag} */,
  {32'h407b1e2e, 32'h3f384994} /* (18, 18, 11) {real, imag} */,
  {32'hc0257ecb, 32'hbf2d6f70} /* (18, 18, 10) {real, imag} */,
  {32'hc0d17072, 32'h4140c914} /* (18, 18, 9) {real, imag} */,
  {32'h40fbf163, 32'h40b34ead} /* (18, 18, 8) {real, imag} */,
  {32'hc024d132, 32'h3c085d00} /* (18, 18, 7) {real, imag} */,
  {32'h401b47d4, 32'h411b11db} /* (18, 18, 6) {real, imag} */,
  {32'h4187bf7c, 32'hc1453ea6} /* (18, 18, 5) {real, imag} */,
  {32'h40928544, 32'h3fe8b9b8} /* (18, 18, 4) {real, imag} */,
  {32'hbff2f8f0, 32'hc089c4b5} /* (18, 18, 3) {real, imag} */,
  {32'hc0620150, 32'h4142f1de} /* (18, 18, 2) {real, imag} */,
  {32'h3f2e5d90, 32'hc10f50f0} /* (18, 18, 1) {real, imag} */,
  {32'hbf095234, 32'h3f9a8604} /* (18, 18, 0) {real, imag} */,
  {32'h411ddb5d, 32'h4091b79b} /* (18, 17, 31) {real, imag} */,
  {32'h40021c4e, 32'hc18696af} /* (18, 17, 30) {real, imag} */,
  {32'h409295de, 32'hbfcb50ac} /* (18, 17, 29) {real, imag} */,
  {32'h4101efdf, 32'hc130e602} /* (18, 17, 28) {real, imag} */,
  {32'hc00ea75b, 32'h3f96b805} /* (18, 17, 27) {real, imag} */,
  {32'h4147f1d9, 32'h41231c54} /* (18, 17, 26) {real, imag} */,
  {32'h4071c9bc, 32'h3e4eb058} /* (18, 17, 25) {real, imag} */,
  {32'hc0031940, 32'hc15593d1} /* (18, 17, 24) {real, imag} */,
  {32'h403e43bc, 32'h3f5904b8} /* (18, 17, 23) {real, imag} */,
  {32'h408ef217, 32'h3f26c18c} /* (18, 17, 22) {real, imag} */,
  {32'hc0909653, 32'h40d51d4e} /* (18, 17, 21) {real, imag} */,
  {32'hc061ac90, 32'h3eda7fa8} /* (18, 17, 20) {real, imag} */,
  {32'hc0685d00, 32'hc094bac2} /* (18, 17, 19) {real, imag} */,
  {32'h3fc4f7dd, 32'h4071c559} /* (18, 17, 18) {real, imag} */,
  {32'h3fc36cd1, 32'h400d152c} /* (18, 17, 17) {real, imag} */,
  {32'hbf020c90, 32'h406afc5a} /* (18, 17, 16) {real, imag} */,
  {32'h3ead6604, 32'hbf3befb0} /* (18, 17, 15) {real, imag} */,
  {32'h3f267ad6, 32'hbec8d218} /* (18, 17, 14) {real, imag} */,
  {32'hc028ec8c, 32'hbfbc10c2} /* (18, 17, 13) {real, imag} */,
  {32'h3f3673d0, 32'h402191bf} /* (18, 17, 12) {real, imag} */,
  {32'h40940a4b, 32'hc08e044a} /* (18, 17, 11) {real, imag} */,
  {32'h4103ffb4, 32'h40d1094c} /* (18, 17, 10) {real, imag} */,
  {32'hbfbf4b0f, 32'hc0a0aa4b} /* (18, 17, 9) {real, imag} */,
  {32'hc0b3f0bc, 32'h407afc14} /* (18, 17, 8) {real, imag} */,
  {32'h405f6030, 32'hc07ca96a} /* (18, 17, 7) {real, imag} */,
  {32'hc0dcf07e, 32'hc005c958} /* (18, 17, 6) {real, imag} */,
  {32'h40b05918, 32'h3fb17f39} /* (18, 17, 5) {real, imag} */,
  {32'hc13d646d, 32'hbf6ccd18} /* (18, 17, 4) {real, imag} */,
  {32'h411b52ac, 32'h40fe3601} /* (18, 17, 3) {real, imag} */,
  {32'h3e217d48, 32'h40040b68} /* (18, 17, 2) {real, imag} */,
  {32'hc0d41623, 32'h41814241} /* (18, 17, 1) {real, imag} */,
  {32'hc1583cfd, 32'h40c0124f} /* (18, 17, 0) {real, imag} */,
  {32'h3f926ebe, 32'h419ae01e} /* (18, 16, 31) {real, imag} */,
  {32'hc10a7411, 32'hc1643791} /* (18, 16, 30) {real, imag} */,
  {32'h40bbb40d, 32'h408cc296} /* (18, 16, 29) {real, imag} */,
  {32'h40952286, 32'hbeca04a0} /* (18, 16, 28) {real, imag} */,
  {32'h4107e0e9, 32'hc0daf037} /* (18, 16, 27) {real, imag} */,
  {32'hbf869ab4, 32'hc048965a} /* (18, 16, 26) {real, imag} */,
  {32'hc02245f0, 32'h3fb385dc} /* (18, 16, 25) {real, imag} */,
  {32'hbfee4743, 32'hbff7f919} /* (18, 16, 24) {real, imag} */,
  {32'h3fa57430, 32'h405e0442} /* (18, 16, 23) {real, imag} */,
  {32'hbf27d5d0, 32'h4127c720} /* (18, 16, 22) {real, imag} */,
  {32'hbf9d130e, 32'h3e61fa72} /* (18, 16, 21) {real, imag} */,
  {32'h3fe1f3f7, 32'hbf998608} /* (18, 16, 20) {real, imag} */,
  {32'hc02ec959, 32'h3fd5bbeb} /* (18, 16, 19) {real, imag} */,
  {32'h3f733e98, 32'h3f566c2c} /* (18, 16, 18) {real, imag} */,
  {32'h3e03c0a4, 32'hbf3e4d10} /* (18, 16, 17) {real, imag} */,
  {32'h3e1f7620, 32'h3fa84858} /* (18, 16, 16) {real, imag} */,
  {32'hbebde55e, 32'h3f16bcd0} /* (18, 16, 15) {real, imag} */,
  {32'hc036276a, 32'hc00ec761} /* (18, 16, 14) {real, imag} */,
  {32'h40668a1f, 32'hc0784b70} /* (18, 16, 13) {real, imag} */,
  {32'h403b200c, 32'hbe2cbb20} /* (18, 16, 12) {real, imag} */,
  {32'hbe247430, 32'h3f6fc0d4} /* (18, 16, 11) {real, imag} */,
  {32'h403798d8, 32'h40821c39} /* (18, 16, 10) {real, imag} */,
  {32'h4074ce1e, 32'hc06760e2} /* (18, 16, 9) {real, imag} */,
  {32'hc0515860, 32'h402b1222} /* (18, 16, 8) {real, imag} */,
  {32'h40a40e23, 32'h40dcf4a3} /* (18, 16, 7) {real, imag} */,
  {32'hc100986c, 32'hc0e7c143} /* (18, 16, 6) {real, imag} */,
  {32'hc01c081f, 32'hc0d88f0f} /* (18, 16, 5) {real, imag} */,
  {32'h40c0a79a, 32'hc0ec62bf} /* (18, 16, 4) {real, imag} */,
  {32'hc0467e7e, 32'h40ad62f8} /* (18, 16, 3) {real, imag} */,
  {32'hc0839d3c, 32'h40c3112e} /* (18, 16, 2) {real, imag} */,
  {32'hc08410c2, 32'hbf6e71d0} /* (18, 16, 1) {real, imag} */,
  {32'h40575fb0, 32'hc02b3397} /* (18, 16, 0) {real, imag} */,
  {32'h4064ba17, 32'h405ce27e} /* (18, 15, 31) {real, imag} */,
  {32'h4090855c, 32'hc09bed90} /* (18, 15, 30) {real, imag} */,
  {32'h415fe12a, 32'h3ff6e3e3} /* (18, 15, 29) {real, imag} */,
  {32'h40a0691e, 32'h419574c8} /* (18, 15, 28) {real, imag} */,
  {32'hbed58efc, 32'hc0676386} /* (18, 15, 27) {real, imag} */,
  {32'h40b3172d, 32'hc161406a} /* (18, 15, 26) {real, imag} */,
  {32'hc1000e7a, 32'hbf81899a} /* (18, 15, 25) {real, imag} */,
  {32'h407510fc, 32'hc0b9e12e} /* (18, 15, 24) {real, imag} */,
  {32'h4022e062, 32'hc083a412} /* (18, 15, 23) {real, imag} */,
  {32'h409bc94d, 32'h4085958a} /* (18, 15, 22) {real, imag} */,
  {32'hc05c3b7e, 32'h3dbc5f00} /* (18, 15, 21) {real, imag} */,
  {32'hc00fb926, 32'h40160fea} /* (18, 15, 20) {real, imag} */,
  {32'hbfd9edc5, 32'hc0a4a4be} /* (18, 15, 19) {real, imag} */,
  {32'h3fb6ad8a, 32'hbf2a78a0} /* (18, 15, 18) {real, imag} */,
  {32'hbf7216bc, 32'h400adbbc} /* (18, 15, 17) {real, imag} */,
  {32'h3f5f29ae, 32'hbfd7993c} /* (18, 15, 16) {real, imag} */,
  {32'hc05eed6f, 32'hbfcb8449} /* (18, 15, 15) {real, imag} */,
  {32'hc05f9deb, 32'hc09babdc} /* (18, 15, 14) {real, imag} */,
  {32'hc05c9780, 32'h3ec2a780} /* (18, 15, 13) {real, imag} */,
  {32'hc0159e9c, 32'hc12b848a} /* (18, 15, 12) {real, imag} */,
  {32'hc08cfcc0, 32'hc01d9108} /* (18, 15, 11) {real, imag} */,
  {32'h411183ce, 32'h3f8c502e} /* (18, 15, 10) {real, imag} */,
  {32'h4110424c, 32'h40a5d4b6} /* (18, 15, 9) {real, imag} */,
  {32'h404d5a6c, 32'h404b59d7} /* (18, 15, 8) {real, imag} */,
  {32'hc0b1e0b1, 32'hc0b19a2e} /* (18, 15, 7) {real, imag} */,
  {32'hc049f6ee, 32'hbe9dd730} /* (18, 15, 6) {real, imag} */,
  {32'h402fd12a, 32'h40a0eb6b} /* (18, 15, 5) {real, imag} */,
  {32'hc119f91d, 32'h40b6d2e9} /* (18, 15, 4) {real, imag} */,
  {32'h409c709b, 32'h3feec043} /* (18, 15, 3) {real, imag} */,
  {32'hc0c68e40, 32'h4087309c} /* (18, 15, 2) {real, imag} */,
  {32'hc12ccf6a, 32'hbfdff703} /* (18, 15, 1) {real, imag} */,
  {32'h407f7684, 32'h3f96eb84} /* (18, 15, 0) {real, imag} */,
  {32'hbf59323c, 32'h415739b0} /* (18, 14, 31) {real, imag} */,
  {32'h410194a2, 32'h40975b94} /* (18, 14, 30) {real, imag} */,
  {32'hc0adb3c9, 32'h40ed9f4c} /* (18, 14, 29) {real, imag} */,
  {32'h418bba08, 32'h40af7e1a} /* (18, 14, 28) {real, imag} */,
  {32'hc088d089, 32'hbe400760} /* (18, 14, 27) {real, imag} */,
  {32'hc1083e84, 32'h407aee4f} /* (18, 14, 26) {real, imag} */,
  {32'hc0e4cf06, 32'h3ffcc732} /* (18, 14, 25) {real, imag} */,
  {32'hbf4c6ce4, 32'hc01e5cd4} /* (18, 14, 24) {real, imag} */,
  {32'hc0ba8aaa, 32'h3f20c520} /* (18, 14, 23) {real, imag} */,
  {32'hc0feb9b8, 32'hbfd2ca0c} /* (18, 14, 22) {real, imag} */,
  {32'hbfab59a8, 32'hc0d2db3d} /* (18, 14, 21) {real, imag} */,
  {32'hc0bdff5a, 32'hc0b5565f} /* (18, 14, 20) {real, imag} */,
  {32'hc0c74fd0, 32'h408953e8} /* (18, 14, 19) {real, imag} */,
  {32'hc02c1248, 32'hbfcb172c} /* (18, 14, 18) {real, imag} */,
  {32'h3fb781ba, 32'hbf9f82f2} /* (18, 14, 17) {real, imag} */,
  {32'h401d55e6, 32'hbf016bc6} /* (18, 14, 16) {real, imag} */,
  {32'h3f4b326c, 32'h3fd72022} /* (18, 14, 15) {real, imag} */,
  {32'h3f533d80, 32'h3f7e47d1} /* (18, 14, 14) {real, imag} */,
  {32'h4057bbc8, 32'hc0a31c6c} /* (18, 14, 13) {real, imag} */,
  {32'h4065a253, 32'h40bee161} /* (18, 14, 12) {real, imag} */,
  {32'h40b4df8d, 32'h3ecebdf0} /* (18, 14, 11) {real, imag} */,
  {32'h412e3570, 32'hbf84c46c} /* (18, 14, 10) {real, imag} */,
  {32'hc16042e1, 32'hc11d284a} /* (18, 14, 9) {real, imag} */,
  {32'h4011790b, 32'h4032c5d2} /* (18, 14, 8) {real, imag} */,
  {32'h412d1db1, 32'h409e74bc} /* (18, 14, 7) {real, imag} */,
  {32'h408dbdd3, 32'h3fe54e5a} /* (18, 14, 6) {real, imag} */,
  {32'h3f9311d0, 32'hc14931f0} /* (18, 14, 5) {real, imag} */,
  {32'hbfebf4f0, 32'h40a90304} /* (18, 14, 4) {real, imag} */,
  {32'h3fb0148c, 32'hc15c921c} /* (18, 14, 3) {real, imag} */,
  {32'h3f9c8fc0, 32'hc08d4e14} /* (18, 14, 2) {real, imag} */,
  {32'h3f9284c6, 32'h410b68f2} /* (18, 14, 1) {real, imag} */,
  {32'hc07ba1a4, 32'h40852b1a} /* (18, 14, 0) {real, imag} */,
  {32'hc17d65e9, 32'h40b5b886} /* (18, 13, 31) {real, imag} */,
  {32'hc034fde8, 32'hbd6047f0} /* (18, 13, 30) {real, imag} */,
  {32'h40f75a79, 32'h40b2a339} /* (18, 13, 29) {real, imag} */,
  {32'h3fa9698c, 32'hc10b6abb} /* (18, 13, 28) {real, imag} */,
  {32'hc08412e6, 32'hc112ab98} /* (18, 13, 27) {real, imag} */,
  {32'h411b440a, 32'hc122fea4} /* (18, 13, 26) {real, imag} */,
  {32'hc1123de0, 32'h4102d312} /* (18, 13, 25) {real, imag} */,
  {32'hc04d0d2a, 32'hc0dd1a6c} /* (18, 13, 24) {real, imag} */,
  {32'h3e89ea2a, 32'hc03a9006} /* (18, 13, 23) {real, imag} */,
  {32'h40477fc6, 32'h3e2ceae0} /* (18, 13, 22) {real, imag} */,
  {32'hbef83f28, 32'hc0af6764} /* (18, 13, 21) {real, imag} */,
  {32'hbfb50fa8, 32'h3e8fe0b0} /* (18, 13, 20) {real, imag} */,
  {32'hc0be6bb3, 32'hbf849378} /* (18, 13, 19) {real, imag} */,
  {32'hc06eb6a8, 32'h3f366fd9} /* (18, 13, 18) {real, imag} */,
  {32'h3ffdacd6, 32'h3fd90d78} /* (18, 13, 17) {real, imag} */,
  {32'hc0614010, 32'hbffa029c} /* (18, 13, 16) {real, imag} */,
  {32'h3ffe971e, 32'hbeb214a0} /* (18, 13, 15) {real, imag} */,
  {32'h409d9a78, 32'h402655f7} /* (18, 13, 14) {real, imag} */,
  {32'h408af11d, 32'h3fb58a40} /* (18, 13, 13) {real, imag} */,
  {32'hc0e64fb2, 32'h40a812ed} /* (18, 13, 12) {real, imag} */,
  {32'hc0c56c5e, 32'h4025a658} /* (18, 13, 11) {real, imag} */,
  {32'h3fbb5044, 32'h40c394db} /* (18, 13, 10) {real, imag} */,
  {32'h3ffcd9ca, 32'hc0ee8f1f} /* (18, 13, 9) {real, imag} */,
  {32'h41170980, 32'h411c0854} /* (18, 13, 8) {real, imag} */,
  {32'hc0e328f9, 32'h400fa14e} /* (18, 13, 7) {real, imag} */,
  {32'hc1746756, 32'h417d4e2e} /* (18, 13, 6) {real, imag} */,
  {32'h408adb4e, 32'h4139b1b8} /* (18, 13, 5) {real, imag} */,
  {32'h4120fa94, 32'h4029be98} /* (18, 13, 4) {real, imag} */,
  {32'hc163d9a4, 32'h417dd720} /* (18, 13, 3) {real, imag} */,
  {32'hc18244c6, 32'h3e77044c} /* (18, 13, 2) {real, imag} */,
  {32'h40e9c486, 32'hc1223e83} /* (18, 13, 1) {real, imag} */,
  {32'hc180a651, 32'hc1708c86} /* (18, 13, 0) {real, imag} */,
  {32'h40d12cbe, 32'h410fa7b2} /* (18, 12, 31) {real, imag} */,
  {32'hc15d39ad, 32'hc0b90418} /* (18, 12, 30) {real, imag} */,
  {32'h41564e1e, 32'h400be748} /* (18, 12, 29) {real, imag} */,
  {32'hc1af53fd, 32'hc143d64e} /* (18, 12, 28) {real, imag} */,
  {32'hc1286c3a, 32'hc18edf7c} /* (18, 12, 27) {real, imag} */,
  {32'h3f984122, 32'hbf94edee} /* (18, 12, 26) {real, imag} */,
  {32'h4168a3bc, 32'hc1748101} /* (18, 12, 25) {real, imag} */,
  {32'h4150e024, 32'hbdf9eba0} /* (18, 12, 24) {real, imag} */,
  {32'h40ce73d9, 32'h411c8212} /* (18, 12, 23) {real, imag} */,
  {32'hc146f6b2, 32'hc14413a8} /* (18, 12, 22) {real, imag} */,
  {32'h3ff03280, 32'hc10c85c2} /* (18, 12, 21) {real, imag} */,
  {32'h40940c28, 32'h405f9ec6} /* (18, 12, 20) {real, imag} */,
  {32'h3fc1cd0c, 32'hbf0c8d50} /* (18, 12, 19) {real, imag} */,
  {32'h3f070f6a, 32'hc08ef018} /* (18, 12, 18) {real, imag} */,
  {32'hbf5ecc04, 32'h3e805002} /* (18, 12, 17) {real, imag} */,
  {32'hbde7a400, 32'h400d9d59} /* (18, 12, 16) {real, imag} */,
  {32'h40d4ee0c, 32'h3fb772a4} /* (18, 12, 15) {real, imag} */,
  {32'hc06f4c7a, 32'h3ff7d8c4} /* (18, 12, 14) {real, imag} */,
  {32'h3fd8eccc, 32'h3f86fa78} /* (18, 12, 13) {real, imag} */,
  {32'h408d7e94, 32'h406df75e} /* (18, 12, 12) {real, imag} */,
  {32'hc19a1712, 32'h40434f76} /* (18, 12, 11) {real, imag} */,
  {32'h406d5ef2, 32'hc0ca9e88} /* (18, 12, 10) {real, imag} */,
  {32'hc0b0d6c1, 32'h3f656b80} /* (18, 12, 9) {real, imag} */,
  {32'hc0e86827, 32'hc0d1ed48} /* (18, 12, 8) {real, imag} */,
  {32'hc14024dc, 32'hc038b33c} /* (18, 12, 7) {real, imag} */,
  {32'hc0d39302, 32'hc0583885} /* (18, 12, 6) {real, imag} */,
  {32'hc1e09401, 32'hc1818b0a} /* (18, 12, 5) {real, imag} */,
  {32'h40686cd0, 32'h411205b8} /* (18, 12, 4) {real, imag} */,
  {32'hc16a8842, 32'h41236584} /* (18, 12, 3) {real, imag} */,
  {32'h41a3676e, 32'h4117628c} /* (18, 12, 2) {real, imag} */,
  {32'hc10d5e21, 32'h40b34e40} /* (18, 12, 1) {real, imag} */,
  {32'h4159a941, 32'hbf8f82ce} /* (18, 12, 0) {real, imag} */,
  {32'h4193774f, 32'h4104321a} /* (18, 11, 31) {real, imag} */,
  {32'h4059a0ac, 32'h41b744fa} /* (18, 11, 30) {real, imag} */,
  {32'hc147f9b9, 32'hc032514c} /* (18, 11, 29) {real, imag} */,
  {32'h3d367600, 32'hc1832b68} /* (18, 11, 28) {real, imag} */,
  {32'hc1868aa2, 32'h4035935c} /* (18, 11, 27) {real, imag} */,
  {32'h3fba97dc, 32'h41358ad9} /* (18, 11, 26) {real, imag} */,
  {32'hc028078d, 32'hc0b723fa} /* (18, 11, 25) {real, imag} */,
  {32'hbe348780, 32'h414c2284} /* (18, 11, 24) {real, imag} */,
  {32'h3f33aa82, 32'h3f5b9c6c} /* (18, 11, 23) {real, imag} */,
  {32'h41896121, 32'h40a5a77d} /* (18, 11, 22) {real, imag} */,
  {32'hc0c5f8fb, 32'hbf5b54b8} /* (18, 11, 21) {real, imag} */,
  {32'h40d4b522, 32'hc0e65099} /* (18, 11, 20) {real, imag} */,
  {32'hc0b53b82, 32'h414513e5} /* (18, 11, 19) {real, imag} */,
  {32'h40ee94cc, 32'h407f8daa} /* (18, 11, 18) {real, imag} */,
  {32'hc0cb1f52, 32'hbfda5ea4} /* (18, 11, 17) {real, imag} */,
  {32'h3ebda570, 32'h408c3baf} /* (18, 11, 16) {real, imag} */,
  {32'h40a6a79a, 32'h400febae} /* (18, 11, 15) {real, imag} */,
  {32'hc09663b8, 32'hc1070a40} /* (18, 11, 14) {real, imag} */,
  {32'h4016d4ad, 32'h40da063e} /* (18, 11, 13) {real, imag} */,
  {32'hbfcfff1a, 32'hbe0fa9e0} /* (18, 11, 12) {real, imag} */,
  {32'h41139e9e, 32'h40358cda} /* (18, 11, 11) {real, imag} */,
  {32'hc15032ca, 32'hc14f8878} /* (18, 11, 10) {real, imag} */,
  {32'hc04f884a, 32'hc104e2b3} /* (18, 11, 9) {real, imag} */,
  {32'h41aca665, 32'h404a3aca} /* (18, 11, 8) {real, imag} */,
  {32'h40586b47, 32'h413ea96b} /* (18, 11, 7) {real, imag} */,
  {32'h40f70e47, 32'hbfcb4bd0} /* (18, 11, 6) {real, imag} */,
  {32'h41e78e9c, 32'h419f58dc} /* (18, 11, 5) {real, imag} */,
  {32'h41a0ff57, 32'hc1ca945e} /* (18, 11, 4) {real, imag} */,
  {32'h41e531fe, 32'h41ba20b2} /* (18, 11, 3) {real, imag} */,
  {32'hc115f363, 32'h400a9e9c} /* (18, 11, 2) {real, imag} */,
  {32'h41be58c3, 32'hc1bd8457} /* (18, 11, 1) {real, imag} */,
  {32'hc0b2027d, 32'h416d2690} /* (18, 11, 0) {real, imag} */,
  {32'h41fd6594, 32'hc134e454} /* (18, 10, 31) {real, imag} */,
  {32'h41d72d9c, 32'h41967a33} /* (18, 10, 30) {real, imag} */,
  {32'hc0b87d7f, 32'hc017b160} /* (18, 10, 29) {real, imag} */,
  {32'hc21f6271, 32'hc0cf53be} /* (18, 10, 28) {real, imag} */,
  {32'hc1ccd3d6, 32'hc042bfb6} /* (18, 10, 27) {real, imag} */,
  {32'h3fb20294, 32'h411e2885} /* (18, 10, 26) {real, imag} */,
  {32'h413c67cd, 32'h412c2e0c} /* (18, 10, 25) {real, imag} */,
  {32'hc180bf2b, 32'hbf48ec70} /* (18, 10, 24) {real, imag} */,
  {32'h41034b5c, 32'h3fd12ee9} /* (18, 10, 23) {real, imag} */,
  {32'hc153c5c2, 32'hc0dd5bb7} /* (18, 10, 22) {real, imag} */,
  {32'h410a3540, 32'h40b9bdb8} /* (18, 10, 21) {real, imag} */,
  {32'h414e1834, 32'hbfb2ace0} /* (18, 10, 20) {real, imag} */,
  {32'h3f6eb638, 32'h402709a0} /* (18, 10, 19) {real, imag} */,
  {32'h40894ab7, 32'h4017cd13} /* (18, 10, 18) {real, imag} */,
  {32'h40310f1a, 32'h407d0ace} /* (18, 10, 17) {real, imag} */,
  {32'h40b54c6a, 32'hbf0e2ef0} /* (18, 10, 16) {real, imag} */,
  {32'hbe76e960, 32'hc04bcb7e} /* (18, 10, 15) {real, imag} */,
  {32'h3e8c14f0, 32'h4021402d} /* (18, 10, 14) {real, imag} */,
  {32'h4122601c, 32'h3d350b00} /* (18, 10, 13) {real, imag} */,
  {32'h40933250, 32'hc0b09346} /* (18, 10, 12) {real, imag} */,
  {32'h40ad476d, 32'hc1b171ae} /* (18, 10, 11) {real, imag} */,
  {32'h40c758fb, 32'hc09e62dd} /* (18, 10, 10) {real, imag} */,
  {32'h40989b9f, 32'hc07436ea} /* (18, 10, 9) {real, imag} */,
  {32'h40a12b80, 32'hc0493116} /* (18, 10, 8) {real, imag} */,
  {32'hc1785757, 32'hc1263ee2} /* (18, 10, 7) {real, imag} */,
  {32'h4127c34a, 32'hc1a5c21c} /* (18, 10, 6) {real, imag} */,
  {32'h4199d796, 32'hc0860c9f} /* (18, 10, 5) {real, imag} */,
  {32'hc15ca608, 32'hc1661eb1} /* (18, 10, 4) {real, imag} */,
  {32'hbf83cfbc, 32'h41c51cd2} /* (18, 10, 3) {real, imag} */,
  {32'hc06894d0, 32'h406bcfe8} /* (18, 10, 2) {real, imag} */,
  {32'hc072f1c0, 32'h405880b6} /* (18, 10, 1) {real, imag} */,
  {32'h4194af34, 32'hc1882a32} /* (18, 10, 0) {real, imag} */,
  {32'h41612040, 32'hc145c7d1} /* (18, 9, 31) {real, imag} */,
  {32'hc09d2ce0, 32'hc22a9dfd} /* (18, 9, 30) {real, imag} */,
  {32'hc1fac1f0, 32'hc16d3ee8} /* (18, 9, 29) {real, imag} */,
  {32'h41d9bfdd, 32'hc0797614} /* (18, 9, 28) {real, imag} */,
  {32'h41cd4a2c, 32'hc1114c99} /* (18, 9, 27) {real, imag} */,
  {32'h412914dd, 32'hc0a76f16} /* (18, 9, 26) {real, imag} */,
  {32'h41a890e7, 32'h411967e8} /* (18, 9, 25) {real, imag} */,
  {32'h3faf6108, 32'hc1c484c3} /* (18, 9, 24) {real, imag} */,
  {32'hc0704a02, 32'hc1023f92} /* (18, 9, 23) {real, imag} */,
  {32'hc0ab68c0, 32'h40927a1c} /* (18, 9, 22) {real, imag} */,
  {32'hc0e11d6a, 32'hbf58b120} /* (18, 9, 21) {real, imag} */,
  {32'h3f5695e8, 32'h409f7007} /* (18, 9, 20) {real, imag} */,
  {32'h40abf908, 32'h40211bae} /* (18, 9, 19) {real, imag} */,
  {32'h40eb82c9, 32'h400e8456} /* (18, 9, 18) {real, imag} */,
  {32'h40ab7f9b, 32'h409faea6} /* (18, 9, 17) {real, imag} */,
  {32'hbfe08a30, 32'h40f60c40} /* (18, 9, 16) {real, imag} */,
  {32'h402a0fba, 32'hbf806d96} /* (18, 9, 15) {real, imag} */,
  {32'hbfcbc74c, 32'hbf9991b4} /* (18, 9, 14) {real, imag} */,
  {32'h3d39e600, 32'h3fb3efd4} /* (18, 9, 13) {real, imag} */,
  {32'hc07f9116, 32'h4058577e} /* (18, 9, 12) {real, imag} */,
  {32'hc097f2ee, 32'h40fa3fa4} /* (18, 9, 11) {real, imag} */,
  {32'h40e41b90, 32'h41b8ab6c} /* (18, 9, 10) {real, imag} */,
  {32'hc0b1d39f, 32'h4117eaf6} /* (18, 9, 9) {real, imag} */,
  {32'h4116728e, 32'hc0dd870c} /* (18, 9, 8) {real, imag} */,
  {32'h3fe917f0, 32'hc1311f08} /* (18, 9, 7) {real, imag} */,
  {32'h41cbdfc2, 32'hc129ad27} /* (18, 9, 6) {real, imag} */,
  {32'hc1c3c124, 32'h3f3775b0} /* (18, 9, 5) {real, imag} */,
  {32'hc22a1862, 32'h41c95798} /* (18, 9, 4) {real, imag} */,
  {32'h41a2634c, 32'hc0fdecf0} /* (18, 9, 3) {real, imag} */,
  {32'hc1dd7684, 32'h4140a068} /* (18, 9, 2) {real, imag} */,
  {32'hc16c1cf4, 32'h401e6984} /* (18, 9, 1) {real, imag} */,
  {32'hc13f021d, 32'hc1c470fe} /* (18, 9, 0) {real, imag} */,
  {32'h40c34254, 32'h41d999bd} /* (18, 8, 31) {real, imag} */,
  {32'hc1930a9d, 32'h41770254} /* (18, 8, 30) {real, imag} */,
  {32'h411db214, 32'h4021bb2d} /* (18, 8, 29) {real, imag} */,
  {32'h412e3e17, 32'hc20a3d1f} /* (18, 8, 28) {real, imag} */,
  {32'hc1bf4843, 32'hc0eac990} /* (18, 8, 27) {real, imag} */,
  {32'hc113b029, 32'h4121492b} /* (18, 8, 26) {real, imag} */,
  {32'hc11ea04c, 32'hc0d378b8} /* (18, 8, 25) {real, imag} */,
  {32'hc1dc5735, 32'hc12e7d9e} /* (18, 8, 24) {real, imag} */,
  {32'h40a75eed, 32'hc145e574} /* (18, 8, 23) {real, imag} */,
  {32'h40bd2271, 32'hc162a5f8} /* (18, 8, 22) {real, imag} */,
  {32'h4071b7b2, 32'hc0f545fe} /* (18, 8, 21) {real, imag} */,
  {32'hbf090e50, 32'hc1a342e2} /* (18, 8, 20) {real, imag} */,
  {32'h41aad25a, 32'h411a8a7c} /* (18, 8, 19) {real, imag} */,
  {32'hc074de0a, 32'h4100c900} /* (18, 8, 18) {real, imag} */,
  {32'hc0694c26, 32'hc0c9c27d} /* (18, 8, 17) {real, imag} */,
  {32'h40b75aad, 32'hbe9a1900} /* (18, 8, 16) {real, imag} */,
  {32'hc032e4d6, 32'h4080f8fd} /* (18, 8, 15) {real, imag} */,
  {32'h3fa33964, 32'hc0800e7b} /* (18, 8, 14) {real, imag} */,
  {32'hc1431fd4, 32'hc11f004c} /* (18, 8, 13) {real, imag} */,
  {32'hc0e5beba, 32'hc0fbfbf2} /* (18, 8, 12) {real, imag} */,
  {32'h3fc6c6a4, 32'hc0eb5b82} /* (18, 8, 11) {real, imag} */,
  {32'hc16d7fd4, 32'hc0a9b8ec} /* (18, 8, 10) {real, imag} */,
  {32'h40ee5b1d, 32'hc119457a} /* (18, 8, 9) {real, imag} */,
  {32'h404bd748, 32'h4213306c} /* (18, 8, 8) {real, imag} */,
  {32'h417907cc, 32'h417a449a} /* (18, 8, 7) {real, imag} */,
  {32'h40372ab0, 32'h420d1bb5} /* (18, 8, 6) {real, imag} */,
  {32'h41cbefe5, 32'h41c713e4} /* (18, 8, 5) {real, imag} */,
  {32'hc17fa235, 32'h4190a510} /* (18, 8, 4) {real, imag} */,
  {32'hc1f613f6, 32'hc0c80ab2} /* (18, 8, 3) {real, imag} */,
  {32'hc2335068, 32'hc128696e} /* (18, 8, 2) {real, imag} */,
  {32'h41bfd57d, 32'h41df244b} /* (18, 8, 1) {real, imag} */,
  {32'h41209ff8, 32'h3fcb71f8} /* (18, 8, 0) {real, imag} */,
  {32'h41c14228, 32'hc158be4e} /* (18, 7, 31) {real, imag} */,
  {32'h4254611c, 32'hc24367b8} /* (18, 7, 30) {real, imag} */,
  {32'hc20a65a3, 32'hc168a8c4} /* (18, 7, 29) {real, imag} */,
  {32'h4041a97c, 32'h4193bee0} /* (18, 7, 28) {real, imag} */,
  {32'hc13f30c0, 32'hc1df0030} /* (18, 7, 27) {real, imag} */,
  {32'hc0aa2a58, 32'h41af5f15} /* (18, 7, 26) {real, imag} */,
  {32'hc20bd4e4, 32'h412f40b6} /* (18, 7, 25) {real, imag} */,
  {32'hc027dcda, 32'hc091f28e} /* (18, 7, 24) {real, imag} */,
  {32'h3fcdb4e4, 32'hc172dab4} /* (18, 7, 23) {real, imag} */,
  {32'h40942224, 32'hc019e462} /* (18, 7, 22) {real, imag} */,
  {32'h4193cf9c, 32'h3fed3f88} /* (18, 7, 21) {real, imag} */,
  {32'h400cf592, 32'hbdd80180} /* (18, 7, 20) {real, imag} */,
  {32'h416d3fb4, 32'hc0b8c0c9} /* (18, 7, 19) {real, imag} */,
  {32'hbf8e98a0, 32'hc00bc302} /* (18, 7, 18) {real, imag} */,
  {32'hc11b90cc, 32'hc02659aa} /* (18, 7, 17) {real, imag} */,
  {32'h40151c82, 32'hc0520b96} /* (18, 7, 16) {real, imag} */,
  {32'hc0ddb868, 32'h40fe704d} /* (18, 7, 15) {real, imag} */,
  {32'hc0311e40, 32'hc1068d54} /* (18, 7, 14) {real, imag} */,
  {32'h3e408d60, 32'h40b50bed} /* (18, 7, 13) {real, imag} */,
  {32'hc093a225, 32'h3f083b00} /* (18, 7, 12) {real, imag} */,
  {32'h3e69d440, 32'hc06c8cac} /* (18, 7, 11) {real, imag} */,
  {32'h41a375d8, 32'h40524206} /* (18, 7, 10) {real, imag} */,
  {32'hc089d17f, 32'hc1849e6c} /* (18, 7, 9) {real, imag} */,
  {32'hc0f1f903, 32'h407ff880} /* (18, 7, 8) {real, imag} */,
  {32'h40e2dff4, 32'hc12ef672} /* (18, 7, 7) {real, imag} */,
  {32'hc1a3b02d, 32'hc00d24f8} /* (18, 7, 6) {real, imag} */,
  {32'h41f41a74, 32'h41fbe372} /* (18, 7, 5) {real, imag} */,
  {32'h40ac97d0, 32'h40a620f9} /* (18, 7, 4) {real, imag} */,
  {32'h4193202a, 32'hc1ce4c56} /* (18, 7, 3) {real, imag} */,
  {32'h41968db7, 32'hc20826a8} /* (18, 7, 2) {real, imag} */,
  {32'hc2509d2e, 32'hc1e54aa3} /* (18, 7, 1) {real, imag} */,
  {32'hc157d4a8, 32'hc192183b} /* (18, 7, 0) {real, imag} */,
  {32'h40cc86d2, 32'hc1d12699} /* (18, 6, 31) {real, imag} */,
  {32'hc209cb54, 32'hbfd2a058} /* (18, 6, 30) {real, imag} */,
  {32'h410c3fc3, 32'hc222207b} /* (18, 6, 29) {real, imag} */,
  {32'hc1a5b53c, 32'h3ed9c3e0} /* (18, 6, 28) {real, imag} */,
  {32'h41c1e024, 32'hbf8e31ae} /* (18, 6, 27) {real, imag} */,
  {32'hc0ff7cbc, 32'h406df7df} /* (18, 6, 26) {real, imag} */,
  {32'h41104bf6, 32'hc0247fe4} /* (18, 6, 25) {real, imag} */,
  {32'h41597f08, 32'h41068f7f} /* (18, 6, 24) {real, imag} */,
  {32'hc06bd782, 32'h4146ea97} /* (18, 6, 23) {real, imag} */,
  {32'h41786304, 32'hc10534fd} /* (18, 6, 22) {real, imag} */,
  {32'hc0b5452e, 32'h410d647c} /* (18, 6, 21) {real, imag} */,
  {32'h408a11a2, 32'h40d8cc40} /* (18, 6, 20) {real, imag} */,
  {32'hc0eb728a, 32'h3f34594e} /* (18, 6, 19) {real, imag} */,
  {32'hc0b72e80, 32'hc0bf4f92} /* (18, 6, 18) {real, imag} */,
  {32'h40a4fb2e, 32'h40f5448b} /* (18, 6, 17) {real, imag} */,
  {32'h415564f4, 32'hc0d5ff2c} /* (18, 6, 16) {real, imag} */,
  {32'hbf97fafe, 32'h40923c3d} /* (18, 6, 15) {real, imag} */,
  {32'hc11f2b7a, 32'h418b1126} /* (18, 6, 14) {real, imag} */,
  {32'hbf6a3a30, 32'hc04e1b9c} /* (18, 6, 13) {real, imag} */,
  {32'hc0ca721c, 32'hc0ba0e20} /* (18, 6, 12) {real, imag} */,
  {32'h41454b31, 32'h409aadfc} /* (18, 6, 11) {real, imag} */,
  {32'h41bb45f0, 32'h416e66f3} /* (18, 6, 10) {real, imag} */,
  {32'hc09e4e55, 32'hc1469bd9} /* (18, 6, 9) {real, imag} */,
  {32'h4145aed0, 32'hc0b71b16} /* (18, 6, 8) {real, imag} */,
  {32'h4160210e, 32'h41d9f358} /* (18, 6, 7) {real, imag} */,
  {32'hc226ad94, 32'h406c4493} /* (18, 6, 6) {real, imag} */,
  {32'hc037b704, 32'hc0ac2ed8} /* (18, 6, 5) {real, imag} */,
  {32'h414c7701, 32'hc10fcc85} /* (18, 6, 4) {real, imag} */,
  {32'hc19ed956, 32'h42117e6d} /* (18, 6, 3) {real, imag} */,
  {32'h41b7ddb0, 32'hc1d6e740} /* (18, 6, 2) {real, imag} */,
  {32'h418d7114, 32'hbf78cf20} /* (18, 6, 1) {real, imag} */,
  {32'hc21de751, 32'hc1f81637} /* (18, 6, 0) {real, imag} */,
  {32'h42616efb, 32'h4255f649} /* (18, 5, 31) {real, imag} */,
  {32'hc1e7866f, 32'hc0c2ed40} /* (18, 5, 30) {real, imag} */,
  {32'h4152ad22, 32'hc046bc50} /* (18, 5, 29) {real, imag} */,
  {32'h4258e4ff, 32'h417048b0} /* (18, 5, 28) {real, imag} */,
  {32'hc1b74686, 32'hc23407ac} /* (18, 5, 27) {real, imag} */,
  {32'hc0b7f7b8, 32'hc1cef181} /* (18, 5, 26) {real, imag} */,
  {32'h419fde41, 32'h404bd294} /* (18, 5, 25) {real, imag} */,
  {32'h418d9e40, 32'h41daa027} /* (18, 5, 24) {real, imag} */,
  {32'hbfdf8490, 32'hc11c2381} /* (18, 5, 23) {real, imag} */,
  {32'h41b15646, 32'h40c1935a} /* (18, 5, 22) {real, imag} */,
  {32'h404cfe44, 32'h41152b4c} /* (18, 5, 21) {real, imag} */,
  {32'hc19ab3a6, 32'h416ceb48} /* (18, 5, 20) {real, imag} */,
  {32'hc17db195, 32'h4109293f} /* (18, 5, 19) {real, imag} */,
  {32'hc064941a, 32'hc05e8150} /* (18, 5, 18) {real, imag} */,
  {32'h416bdb82, 32'h418fbe64} /* (18, 5, 17) {real, imag} */,
  {32'h40baad40, 32'h3fe1cec0} /* (18, 5, 16) {real, imag} */,
  {32'h4075b388, 32'h403a0784} /* (18, 5, 15) {real, imag} */,
  {32'h3e8a4750, 32'hc0f15750} /* (18, 5, 14) {real, imag} */,
  {32'h408e286a, 32'h407f65bc} /* (18, 5, 13) {real, imag} */,
  {32'hc19881da, 32'h418ae662} /* (18, 5, 12) {real, imag} */,
  {32'hc1ad0f4e, 32'hc1cf4c48} /* (18, 5, 11) {real, imag} */,
  {32'hc0f45f80, 32'h4035227c} /* (18, 5, 10) {real, imag} */,
  {32'hc223866e, 32'h418f772a} /* (18, 5, 9) {real, imag} */,
  {32'hbeaf7f60, 32'hc0a474ac} /* (18, 5, 8) {real, imag} */,
  {32'hc0be6a8b, 32'h41cbba70} /* (18, 5, 7) {real, imag} */,
  {32'h41c5bfb8, 32'h419d0f4b} /* (18, 5, 6) {real, imag} */,
  {32'hc1a866b2, 32'hc1757dfc} /* (18, 5, 5) {real, imag} */,
  {32'h40a59f98, 32'hc09a0208} /* (18, 5, 4) {real, imag} */,
  {32'hc1d82b3b, 32'hc215bc71} /* (18, 5, 3) {real, imag} */,
  {32'hc1057eee, 32'hc2b26d8a} /* (18, 5, 2) {real, imag} */,
  {32'h41160314, 32'hbfd112e0} /* (18, 5, 1) {real, imag} */,
  {32'h42121a10, 32'hc224b1ac} /* (18, 5, 0) {real, imag} */,
  {32'hc23bc6ca, 32'hc255ceac} /* (18, 4, 31) {real, imag} */,
  {32'hbe335800, 32'h4186dffc} /* (18, 4, 30) {real, imag} */,
  {32'h425caa11, 32'h41ee2600} /* (18, 4, 29) {real, imag} */,
  {32'hc28e99af, 32'h42627a87} /* (18, 4, 28) {real, imag} */,
  {32'h4285d6d4, 32'h41ad325a} /* (18, 4, 27) {real, imag} */,
  {32'hc07fc7d4, 32'hc07d8f9c} /* (18, 4, 26) {real, imag} */,
  {32'hc196c4a5, 32'h4177e828} /* (18, 4, 25) {real, imag} */,
  {32'h41fac93d, 32'h401e2ec0} /* (18, 4, 24) {real, imag} */,
  {32'hc20485ae, 32'hbfdd6a1c} /* (18, 4, 23) {real, imag} */,
  {32'hbf1ccd14, 32'hc0ab7a96} /* (18, 4, 22) {real, imag} */,
  {32'hc11c4873, 32'hc1c1b50a} /* (18, 4, 21) {real, imag} */,
  {32'hc11d96e9, 32'h417b86c3} /* (18, 4, 20) {real, imag} */,
  {32'hc0853cb0, 32'hbf5be2a0} /* (18, 4, 19) {real, imag} */,
  {32'hc1921c2a, 32'h411b838a} /* (18, 4, 18) {real, imag} */,
  {32'h3f772188, 32'hc0a408b8} /* (18, 4, 17) {real, imag} */,
  {32'hc093bc7c, 32'hbff1e690} /* (18, 4, 16) {real, imag} */,
  {32'h413d4744, 32'hc06445b0} /* (18, 4, 15) {real, imag} */,
  {32'hc0e650f0, 32'hbfd2b890} /* (18, 4, 14) {real, imag} */,
  {32'hc193a2cc, 32'hc0b05764} /* (18, 4, 13) {real, imag} */,
  {32'h40f815b6, 32'h3f91cc58} /* (18, 4, 12) {real, imag} */,
  {32'hc190679a, 32'hbfe4b910} /* (18, 4, 11) {real, imag} */,
  {32'h3f97cb4e, 32'h41ef710e} /* (18, 4, 10) {real, imag} */,
  {32'hc0a3a688, 32'hc0e34a1f} /* (18, 4, 9) {real, imag} */,
  {32'h41bbcc6b, 32'h428cb7da} /* (18, 4, 8) {real, imag} */,
  {32'hc2586fda, 32'hc1d77372} /* (18, 4, 7) {real, imag} */,
  {32'h4167afeb, 32'h420ad95c} /* (18, 4, 6) {real, imag} */,
  {32'hc03a53d0, 32'h4206d083} /* (18, 4, 5) {real, imag} */,
  {32'h421ac65e, 32'hc03a1190} /* (18, 4, 4) {real, imag} */,
  {32'h424fb1cf, 32'hc1474808} /* (18, 4, 3) {real, imag} */,
  {32'h4281c2ea, 32'hc207011d} /* (18, 4, 2) {real, imag} */,
  {32'hc213a276, 32'hc2b85cb2} /* (18, 4, 1) {real, imag} */,
  {32'hc1d766b5, 32'h417c154a} /* (18, 4, 0) {real, imag} */,
  {32'hc10e8bfc, 32'hc1e2e9c9} /* (18, 3, 31) {real, imag} */,
  {32'h41d63ba2, 32'h4057d95c} /* (18, 3, 30) {real, imag} */,
  {32'hc25e1f45, 32'h42388236} /* (18, 3, 29) {real, imag} */,
  {32'hc206fe83, 32'hbfb7af00} /* (18, 3, 28) {real, imag} */,
  {32'h40ef743c, 32'hc17271f2} /* (18, 3, 27) {real, imag} */,
  {32'h427769a4, 32'hc015170e} /* (18, 3, 26) {real, imag} */,
  {32'hc1769c0a, 32'hc2491928} /* (18, 3, 25) {real, imag} */,
  {32'h40ab3e94, 32'h418e6d93} /* (18, 3, 24) {real, imag} */,
  {32'hc0f1fc3e, 32'hc110b296} /* (18, 3, 23) {real, imag} */,
  {32'hc1ab41fe, 32'hc1b6465b} /* (18, 3, 22) {real, imag} */,
  {32'h4095d7d4, 32'hbf67b8c8} /* (18, 3, 21) {real, imag} */,
  {32'hc057f45c, 32'h40f47869} /* (18, 3, 20) {real, imag} */,
  {32'h40151b4c, 32'h40dca010} /* (18, 3, 19) {real, imag} */,
  {32'h419e7c02, 32'h3e8c6410} /* (18, 3, 18) {real, imag} */,
  {32'hc1042cdb, 32'hc12a5a24} /* (18, 3, 17) {real, imag} */,
  {32'h4080a2b8, 32'hc0e1b858} /* (18, 3, 16) {real, imag} */,
  {32'h4193def8, 32'h41872b74} /* (18, 3, 15) {real, imag} */,
  {32'h404c31ac, 32'h4095b393} /* (18, 3, 14) {real, imag} */,
  {32'h417f9007, 32'hc090a470} /* (18, 3, 13) {real, imag} */,
  {32'hc1a56816, 32'hc128c500} /* (18, 3, 12) {real, imag} */,
  {32'hbfff37d6, 32'hc176fb82} /* (18, 3, 11) {real, imag} */,
  {32'h41646724, 32'hbfd0a8d0} /* (18, 3, 10) {real, imag} */,
  {32'hc16b84bd, 32'h41c52425} /* (18, 3, 9) {real, imag} */,
  {32'hc2265c5a, 32'h411f28f2} /* (18, 3, 8) {real, imag} */,
  {32'h4258da0a, 32'hc1f1ef80} /* (18, 3, 7) {real, imag} */,
  {32'hc05552c0, 32'h407b0ade} /* (18, 3, 6) {real, imag} */,
  {32'hc1c56c85, 32'hc20f4e24} /* (18, 3, 5) {real, imag} */,
  {32'h3eb16180, 32'h419ab2b6} /* (18, 3, 4) {real, imag} */,
  {32'h4141edec, 32'h4269c802} /* (18, 3, 3) {real, imag} */,
  {32'h41c57256, 32'h41c3e5f2} /* (18, 3, 2) {real, imag} */,
  {32'hc271a031, 32'h3ff1cbd0} /* (18, 3, 1) {real, imag} */,
  {32'hc209587a, 32'hc211a707} /* (18, 3, 0) {real, imag} */,
  {32'h4307faef, 32'h4255b956} /* (18, 2, 31) {real, imag} */,
  {32'hc2b43ad5, 32'hc0e68e0e} /* (18, 2, 30) {real, imag} */,
  {32'h4242dbff, 32'h41cbcf74} /* (18, 2, 29) {real, imag} */,
  {32'h4244916a, 32'hc1c13c2a} /* (18, 2, 28) {real, imag} */,
  {32'hc1d06310, 32'hc12be5f9} /* (18, 2, 27) {real, imag} */,
  {32'h415cfd92, 32'hc1004900} /* (18, 2, 26) {real, imag} */,
  {32'hc195720a, 32'hc172cc07} /* (18, 2, 25) {real, imag} */,
  {32'hc1c3dd0f, 32'hc00e3452} /* (18, 2, 24) {real, imag} */,
  {32'h42035dac, 32'h40ea6afe} /* (18, 2, 23) {real, imag} */,
  {32'h41b43420, 32'h41d056da} /* (18, 2, 22) {real, imag} */,
  {32'hc15aa4fc, 32'hc0c5688a} /* (18, 2, 21) {real, imag} */,
  {32'h419a9ef7, 32'h40ed7035} /* (18, 2, 20) {real, imag} */,
  {32'hbf73a5b0, 32'hc1064c2b} /* (18, 2, 19) {real, imag} */,
  {32'hbeb9dfc0, 32'hc17e7f0f} /* (18, 2, 18) {real, imag} */,
  {32'hc158edf8, 32'hc0bbe112} /* (18, 2, 17) {real, imag} */,
  {32'hc12db39c, 32'h4099773b} /* (18, 2, 16) {real, imag} */,
  {32'hc005ab60, 32'h4027fe14} /* (18, 2, 15) {real, imag} */,
  {32'h40c0de2c, 32'h3fd68c48} /* (18, 2, 14) {real, imag} */,
  {32'hc1ca3012, 32'hc08f08d2} /* (18, 2, 13) {real, imag} */,
  {32'hc046e078, 32'hc0338b42} /* (18, 2, 12) {real, imag} */,
  {32'hc0468150, 32'hc1223103} /* (18, 2, 11) {real, imag} */,
  {32'h41f9be04, 32'h4093ba2c} /* (18, 2, 10) {real, imag} */,
  {32'h3f0bbc40, 32'h416eb8b1} /* (18, 2, 9) {real, imag} */,
  {32'hc1ffbb01, 32'h412fbf84} /* (18, 2, 8) {real, imag} */,
  {32'h419d59b0, 32'hc1b2a24c} /* (18, 2, 7) {real, imag} */,
  {32'hc1aba52f, 32'h403b8598} /* (18, 2, 6) {real, imag} */,
  {32'hc212a630, 32'hc20dfb27} /* (18, 2, 5) {real, imag} */,
  {32'hc02502b8, 32'hc227b6df} /* (18, 2, 4) {real, imag} */,
  {32'hc09bc238, 32'hc17f7408} /* (18, 2, 3) {real, imag} */,
  {32'hc2ae5a27, 32'hc1887442} /* (18, 2, 2) {real, imag} */,
  {32'h430be65d, 32'h411f0f42} /* (18, 2, 1) {real, imag} */,
  {32'h427fa7d3, 32'hc12bedb0} /* (18, 2, 0) {real, imag} */,
  {32'hc2cdac70, 32'hc1b1966e} /* (18, 1, 31) {real, imag} */,
  {32'h420e3cee, 32'h41b9bae7} /* (18, 1, 30) {real, imag} */,
  {32'h41987af8, 32'hbd96b200} /* (18, 1, 29) {real, imag} */,
  {32'hbf1613b8, 32'hc1a501e5} /* (18, 1, 28) {real, imag} */,
  {32'h41ea0312, 32'hc1a7ae7d} /* (18, 1, 27) {real, imag} */,
  {32'hc11c2ff0, 32'hc24b98c1} /* (18, 1, 26) {real, imag} */,
  {32'h41f64893, 32'h414f0b26} /* (18, 1, 25) {real, imag} */,
  {32'h4031ee88, 32'h4208800c} /* (18, 1, 24) {real, imag} */,
  {32'h412ca4aa, 32'h41776daa} /* (18, 1, 23) {real, imag} */,
  {32'hc2114bcc, 32'h415465a2} /* (18, 1, 22) {real, imag} */,
  {32'h42077aa7, 32'hbec7bdc0} /* (18, 1, 21) {real, imag} */,
  {32'hc0ba5bcf, 32'h3e106bb0} /* (18, 1, 20) {real, imag} */,
  {32'hc1796ee0, 32'h40011f80} /* (18, 1, 19) {real, imag} */,
  {32'h40497be0, 32'h40c06db8} /* (18, 1, 18) {real, imag} */,
  {32'hc10843e5, 32'hc0b68db1} /* (18, 1, 17) {real, imag} */,
  {32'h40570fa0, 32'h4164d9e0} /* (18, 1, 16) {real, imag} */,
  {32'hc12a8f6b, 32'h40388022} /* (18, 1, 15) {real, imag} */,
  {32'h41325dd2, 32'hbe856500} /* (18, 1, 14) {real, imag} */,
  {32'h407ee090, 32'hc0d23c04} /* (18, 1, 13) {real, imag} */,
  {32'h40cb3911, 32'hc01f7393} /* (18, 1, 12) {real, imag} */,
  {32'h41bd18ea, 32'h41da864b} /* (18, 1, 11) {real, imag} */,
  {32'h41fb2bac, 32'hc1507db4} /* (18, 1, 10) {real, imag} */,
  {32'h414c9cd2, 32'h418d4437} /* (18, 1, 9) {real, imag} */,
  {32'h400ff948, 32'h421c323e} /* (18, 1, 8) {real, imag} */,
  {32'hc266ef98, 32'h418405fc} /* (18, 1, 7) {real, imag} */,
  {32'hc144b968, 32'h421c5833} /* (18, 1, 6) {real, imag} */,
  {32'hc20c9295, 32'h416208da} /* (18, 1, 5) {real, imag} */,
  {32'hc0a749d7, 32'hc1a2f83b} /* (18, 1, 4) {real, imag} */,
  {32'h421fd2bf, 32'hc201ea4f} /* (18, 1, 3) {real, imag} */,
  {32'h41bb4add, 32'h42a96aa2} /* (18, 1, 2) {real, imag} */,
  {32'hc30e95ab, 32'hc20522dd} /* (18, 1, 1) {real, imag} */,
  {32'hc2999639, 32'h406a7200} /* (18, 1, 0) {real, imag} */,
  {32'hc21e3d8e, 32'h42b34091} /* (18, 0, 31) {real, imag} */,
  {32'h4294e903, 32'hc1a95ec6} /* (18, 0, 30) {real, imag} */,
  {32'hc263bdd5, 32'h4143442a} /* (18, 0, 29) {real, imag} */,
  {32'hc1de15b2, 32'hbf8b99a6} /* (18, 0, 28) {real, imag} */,
  {32'h3f98dac0, 32'hc081c35c} /* (18, 0, 27) {real, imag} */,
  {32'hc1a6c093, 32'h4161dc0e} /* (18, 0, 26) {real, imag} */,
  {32'hc206919f, 32'h3fca0660} /* (18, 0, 25) {real, imag} */,
  {32'hc1ccfba0, 32'hc07500c8} /* (18, 0, 24) {real, imag} */,
  {32'h418d1bd1, 32'h426f3701} /* (18, 0, 23) {real, imag} */,
  {32'hc1466030, 32'hc1c09cb0} /* (18, 0, 22) {real, imag} */,
  {32'h404da090, 32'hc196d160} /* (18, 0, 21) {real, imag} */,
  {32'h4104f96d, 32'hbecf3a80} /* (18, 0, 20) {real, imag} */,
  {32'hc11b2b86, 32'hc0d8fc5a} /* (18, 0, 19) {real, imag} */,
  {32'h409590d8, 32'hc0a9458a} /* (18, 0, 18) {real, imag} */,
  {32'h40dff56c, 32'hc1a70e08} /* (18, 0, 17) {real, imag} */,
  {32'hc128eae2, 32'h410d94e6} /* (18, 0, 16) {real, imag} */,
  {32'h405a9538, 32'hbf3d2c00} /* (18, 0, 15) {real, imag} */,
  {32'hc1018854, 32'h4028dd4c} /* (18, 0, 14) {real, imag} */,
  {32'h3f08d618, 32'hc128d9af} /* (18, 0, 13) {real, imag} */,
  {32'hbe447bc0, 32'hbf9342ac} /* (18, 0, 12) {real, imag} */,
  {32'h4126328a, 32'h4098fa11} /* (18, 0, 11) {real, imag} */,
  {32'h40233ace, 32'hc112b67c} /* (18, 0, 10) {real, imag} */,
  {32'h42061494, 32'h41bc802e} /* (18, 0, 9) {real, imag} */,
  {32'hc1f0da00, 32'h417bda82} /* (18, 0, 8) {real, imag} */,
  {32'h4210f4f5, 32'hc2638933} /* (18, 0, 7) {real, imag} */,
  {32'hc236c1fa, 32'hc26b7280} /* (18, 0, 6) {real, imag} */,
  {32'h42269f66, 32'h3f6ee2b0} /* (18, 0, 5) {real, imag} */,
  {32'h426446d7, 32'h410cf8cf} /* (18, 0, 4) {real, imag} */,
  {32'h41a2559a, 32'h423155fa} /* (18, 0, 3) {real, imag} */,
  {32'h416c6190, 32'hc1ce87e6} /* (18, 0, 2) {real, imag} */,
  {32'hc1cb43bc, 32'hc2311036} /* (18, 0, 1) {real, imag} */,
  {32'hc24937ec, 32'hc2330ea4} /* (18, 0, 0) {real, imag} */,
  {32'h42b1dec2, 32'hc1a9d806} /* (17, 31, 31) {real, imag} */,
  {32'hc24eddb5, 32'h424de0f7} /* (17, 31, 30) {real, imag} */,
  {32'hc1c8c8a9, 32'h41629b04} /* (17, 31, 29) {real, imag} */,
  {32'h419febd8, 32'hc1cbe7a6} /* (17, 31, 28) {real, imag} */,
  {32'hc223e6eb, 32'hc16ad068} /* (17, 31, 27) {real, imag} */,
  {32'h40681a8c, 32'hc1458912} /* (17, 31, 26) {real, imag} */,
  {32'h414a795a, 32'hc1cab5f8} /* (17, 31, 25) {real, imag} */,
  {32'hc18cdff5, 32'h4133a344} /* (17, 31, 24) {real, imag} */,
  {32'h41cc4d8a, 32'hc1bbd139} /* (17, 31, 23) {real, imag} */,
  {32'h41350b3b, 32'h4148b548} /* (17, 31, 22) {real, imag} */,
  {32'h41281ce3, 32'hc18a7be1} /* (17, 31, 21) {real, imag} */,
  {32'h411bad05, 32'h4179ac8b} /* (17, 31, 20) {real, imag} */,
  {32'h40fe649c, 32'h4094c054} /* (17, 31, 19) {real, imag} */,
  {32'h3ffbad18, 32'h4148bbf4} /* (17, 31, 18) {real, imag} */,
  {32'h4086f5e6, 32'h402bb5c1} /* (17, 31, 17) {real, imag} */,
  {32'hc1805b87, 32'h417c0f00} /* (17, 31, 16) {real, imag} */,
  {32'h3f8e0e68, 32'h40acbaac} /* (17, 31, 15) {real, imag} */,
  {32'h403fb664, 32'h407d3670} /* (17, 31, 14) {real, imag} */,
  {32'hc0b5a940, 32'h412ef524} /* (17, 31, 13) {real, imag} */,
  {32'h4169d503, 32'hc1866192} /* (17, 31, 12) {real, imag} */,
  {32'h3fb72558, 32'h40dc11b3} /* (17, 31, 11) {real, imag} */,
  {32'h402b904c, 32'hc10f86ec} /* (17, 31, 10) {real, imag} */,
  {32'h42279d03, 32'hc17cfac6} /* (17, 31, 9) {real, imag} */,
  {32'hc0cd060c, 32'hc1d4617a} /* (17, 31, 8) {real, imag} */,
  {32'h415eb236, 32'hbe34de40} /* (17, 31, 7) {real, imag} */,
  {32'hc1c54d22, 32'hc099319c} /* (17, 31, 6) {real, imag} */,
  {32'h413f8119, 32'h4018c212} /* (17, 31, 5) {real, imag} */,
  {32'h41396320, 32'h3f71c690} /* (17, 31, 4) {real, imag} */,
  {32'h41c5c113, 32'hc1687822} /* (17, 31, 3) {real, imag} */,
  {32'hc1c7d8e6, 32'hc1ae1526} /* (17, 31, 2) {real, imag} */,
  {32'h42469869, 32'hc138f75b} /* (17, 31, 1) {real, imag} */,
  {32'h4218a34a, 32'hc1f1fbb6} /* (17, 31, 0) {real, imag} */,
  {32'hc23d9c06, 32'h421d0f36} /* (17, 30, 31) {real, imag} */,
  {32'h41e95acf, 32'h41cac6a3} /* (17, 30, 30) {real, imag} */,
  {32'hc278218a, 32'hc1bc7d52} /* (17, 30, 29) {real, imag} */,
  {32'hc18c4f24, 32'hbe988980} /* (17, 30, 28) {real, imag} */,
  {32'h41b0c5f2, 32'h416daa2c} /* (17, 30, 27) {real, imag} */,
  {32'hc0ea12f7, 32'h4268c436} /* (17, 30, 26) {real, imag} */,
  {32'hc0713374, 32'h3f1e9c60} /* (17, 30, 25) {real, imag} */,
  {32'hc15a19e4, 32'hc10a58d2} /* (17, 30, 24) {real, imag} */,
  {32'h400c63dc, 32'hc13e0e84} /* (17, 30, 23) {real, imag} */,
  {32'hc0296eda, 32'hc1044100} /* (17, 30, 22) {real, imag} */,
  {32'h4002017a, 32'h415684aa} /* (17, 30, 21) {real, imag} */,
  {32'h4120863d, 32'h4117678e} /* (17, 30, 20) {real, imag} */,
  {32'h3f125510, 32'hc1726972} /* (17, 30, 19) {real, imag} */,
  {32'hc13e7a58, 32'h408b4e3d} /* (17, 30, 18) {real, imag} */,
  {32'hc0a2ec58, 32'hc05edf26} /* (17, 30, 17) {real, imag} */,
  {32'h402c825e, 32'h414f1a90} /* (17, 30, 16) {real, imag} */,
  {32'h40c4d590, 32'h4144e766} /* (17, 30, 15) {real, imag} */,
  {32'h3fd0ad84, 32'h4090a903} /* (17, 30, 14) {real, imag} */,
  {32'h4080268a, 32'hc16fbd82} /* (17, 30, 13) {real, imag} */,
  {32'hc1255b09, 32'hbecbe330} /* (17, 30, 12) {real, imag} */,
  {32'hc006528a, 32'h420d816a} /* (17, 30, 11) {real, imag} */,
  {32'h40f59383, 32'h412c1528} /* (17, 30, 10) {real, imag} */,
  {32'hc1bb208e, 32'h41f5412e} /* (17, 30, 9) {real, imag} */,
  {32'hc1248334, 32'h41bf25cd} /* (17, 30, 8) {real, imag} */,
  {32'hc0d1ad06, 32'hc2024dd0} /* (17, 30, 7) {real, imag} */,
  {32'h4108867c, 32'hc26ecc00} /* (17, 30, 6) {real, imag} */,
  {32'h422b0643, 32'hc19b5330} /* (17, 30, 5) {real, imag} */,
  {32'hc0c7238c, 32'h41b7b5b8} /* (17, 30, 4) {real, imag} */,
  {32'h41fbd38c, 32'hc1515bb0} /* (17, 30, 3) {real, imag} */,
  {32'hc1fac8bd, 32'h40cee664} /* (17, 30, 2) {real, imag} */,
  {32'hc1c19774, 32'h4116898e} /* (17, 30, 1) {real, imag} */,
  {32'h40fab447, 32'hc28bf07e} /* (17, 30, 0) {real, imag} */,
  {32'h4226a9ce, 32'hc10c46a2} /* (17, 29, 31) {real, imag} */,
  {32'hc0afcb38, 32'hc07635e0} /* (17, 29, 30) {real, imag} */,
  {32'h40d2e673, 32'hc1c620bd} /* (17, 29, 29) {real, imag} */,
  {32'h411ddbaf, 32'hbfb86634} /* (17, 29, 28) {real, imag} */,
  {32'h42174626, 32'h3fb017a4} /* (17, 29, 27) {real, imag} */,
  {32'h3fff3d80, 32'hc1b06954} /* (17, 29, 26) {real, imag} */,
  {32'h407df3fe, 32'h4178f0ee} /* (17, 29, 25) {real, imag} */,
  {32'h41ac7219, 32'h413b9a24} /* (17, 29, 24) {real, imag} */,
  {32'hc17e682c, 32'hbf581d14} /* (17, 29, 23) {real, imag} */,
  {32'hc1a9a7dc, 32'hc201e607} /* (17, 29, 22) {real, imag} */,
  {32'hc118678a, 32'hc12a47ac} /* (17, 29, 21) {real, imag} */,
  {32'h415354f2, 32'h416a51f9} /* (17, 29, 20) {real, imag} */,
  {32'h40d47a7d, 32'hc17d7d74} /* (17, 29, 19) {real, imag} */,
  {32'hc0fceb15, 32'hc0e76ec4} /* (17, 29, 18) {real, imag} */,
  {32'h3edd5c70, 32'h40c7c20a} /* (17, 29, 17) {real, imag} */,
  {32'hc0525620, 32'hbfab8c48} /* (17, 29, 16) {real, imag} */,
  {32'h417b2da8, 32'hc11da4b5} /* (17, 29, 15) {real, imag} */,
  {32'h409214dd, 32'h40bf6b24} /* (17, 29, 14) {real, imag} */,
  {32'hc19d801a, 32'hbfa78440} /* (17, 29, 13) {real, imag} */,
  {32'hc17a30ca, 32'hc0cbffd2} /* (17, 29, 12) {real, imag} */,
  {32'hc2079ad6, 32'hc159d5d2} /* (17, 29, 11) {real, imag} */,
  {32'h4199af08, 32'h4003e510} /* (17, 29, 10) {real, imag} */,
  {32'h40c6ded9, 32'hbf4ef2d4} /* (17, 29, 9) {real, imag} */,
  {32'hc162d92a, 32'h4184eadf} /* (17, 29, 8) {real, imag} */,
  {32'hc18867c4, 32'hc1dc03eb} /* (17, 29, 7) {real, imag} */,
  {32'h41b66056, 32'hc177e451} /* (17, 29, 6) {real, imag} */,
  {32'h423f587a, 32'hc0e23aed} /* (17, 29, 5) {real, imag} */,
  {32'hc0b092ea, 32'h401b4e1e} /* (17, 29, 4) {real, imag} */,
  {32'h3f0bd938, 32'h42252466} /* (17, 29, 3) {real, imag} */,
  {32'hc23be015, 32'h425b277d} /* (17, 29, 2) {real, imag} */,
  {32'h41b5a643, 32'hc088da44} /* (17, 29, 1) {real, imag} */,
  {32'hc21f7192, 32'hc18cf4ce} /* (17, 29, 0) {real, imag} */,
  {32'h40223302, 32'h42399962} /* (17, 28, 31) {real, imag} */,
  {32'hbe00cbf0, 32'h423d65ae} /* (17, 28, 30) {real, imag} */,
  {32'hc06e7254, 32'h424c808a} /* (17, 28, 29) {real, imag} */,
  {32'h41e4462c, 32'hc2229067} /* (17, 28, 28) {real, imag} */,
  {32'h41e17fc6, 32'hc1046f81} /* (17, 28, 27) {real, imag} */,
  {32'hbf2c6410, 32'h41c492c1} /* (17, 28, 26) {real, imag} */,
  {32'hc18f5db0, 32'hc150d64e} /* (17, 28, 25) {real, imag} */,
  {32'hc1514337, 32'h40b95f14} /* (17, 28, 24) {real, imag} */,
  {32'hc12f33d5, 32'hbe932470} /* (17, 28, 23) {real, imag} */,
  {32'hc224b478, 32'h40b19de4} /* (17, 28, 22) {real, imag} */,
  {32'h41837ad9, 32'h41a3e541} /* (17, 28, 21) {real, imag} */,
  {32'hc0dc12ac, 32'hc1ac61b9} /* (17, 28, 20) {real, imag} */,
  {32'h4148ad83, 32'h3fc9a908} /* (17, 28, 19) {real, imag} */,
  {32'h40908be7, 32'h4061a619} /* (17, 28, 18) {real, imag} */,
  {32'h407a688e, 32'hc0dbfd28} /* (17, 28, 17) {real, imag} */,
  {32'h40446710, 32'hc0bba56c} /* (17, 28, 16) {real, imag} */,
  {32'h403e717a, 32'h418c253e} /* (17, 28, 15) {real, imag} */,
  {32'h40952a35, 32'hc1235ca2} /* (17, 28, 14) {real, imag} */,
  {32'hc0f8dcf2, 32'h4034dd94} /* (17, 28, 13) {real, imag} */,
  {32'h40469520, 32'h4186b83b} /* (17, 28, 12) {real, imag} */,
  {32'h3f0dafa0, 32'hc18de56b} /* (17, 28, 11) {real, imag} */,
  {32'h415e0948, 32'h3f827ece} /* (17, 28, 10) {real, imag} */,
  {32'h409f3cee, 32'h40341d16} /* (17, 28, 9) {real, imag} */,
  {32'hbf3b21b0, 32'h41618528} /* (17, 28, 8) {real, imag} */,
  {32'h4257af30, 32'hc1c34dd5} /* (17, 28, 7) {real, imag} */,
  {32'hc1c4b06c, 32'h41f02fd5} /* (17, 28, 6) {real, imag} */,
  {32'h409033e0, 32'h40e3289a} /* (17, 28, 5) {real, imag} */,
  {32'h41483ad7, 32'h420ae23d} /* (17, 28, 4) {real, imag} */,
  {32'hc08f3a4a, 32'hbfc7cc90} /* (17, 28, 3) {real, imag} */,
  {32'hbf5fc0cc, 32'hc2277768} /* (17, 28, 2) {real, imag} */,
  {32'h4116863e, 32'hc23a956a} /* (17, 28, 1) {real, imag} */,
  {32'hc27d6b29, 32'hc16504b8} /* (17, 28, 0) {real, imag} */,
  {32'h42370517, 32'h41190c7a} /* (17, 27, 31) {real, imag} */,
  {32'hc17190a4, 32'hc210f957} /* (17, 27, 30) {real, imag} */,
  {32'h4196894f, 32'hc21e0bee} /* (17, 27, 29) {real, imag} */,
  {32'h425e2b7a, 32'h41c2d317} /* (17, 27, 28) {real, imag} */,
  {32'hc1d0869e, 32'h416a042a} /* (17, 27, 27) {real, imag} */,
  {32'hc04be458, 32'hc11188ec} /* (17, 27, 26) {real, imag} */,
  {32'h41884e6e, 32'h4181414e} /* (17, 27, 25) {real, imag} */,
  {32'h4125e46e, 32'h41a1599a} /* (17, 27, 24) {real, imag} */,
  {32'hc07bc3e6, 32'h4162a110} /* (17, 27, 23) {real, imag} */,
  {32'hc10a0730, 32'hc04cd342} /* (17, 27, 22) {real, imag} */,
  {32'h416d0a29, 32'hc14c131c} /* (17, 27, 21) {real, imag} */,
  {32'h40347636, 32'h400b45a2} /* (17, 27, 20) {real, imag} */,
  {32'hc163a7c2, 32'hc08956da} /* (17, 27, 19) {real, imag} */,
  {32'hc0ca0885, 32'h41246674} /* (17, 27, 18) {real, imag} */,
  {32'h3f2726c8, 32'hc02955be} /* (17, 27, 17) {real, imag} */,
  {32'hc082a2ed, 32'hbfee8920} /* (17, 27, 16) {real, imag} */,
  {32'h40096e1e, 32'h40e98cb1} /* (17, 27, 15) {real, imag} */,
  {32'h3f9bf6fc, 32'hc07aea72} /* (17, 27, 14) {real, imag} */,
  {32'hc09a532c, 32'hbe006cc0} /* (17, 27, 13) {real, imag} */,
  {32'hc08bbebb, 32'hc14d7722} /* (17, 27, 12) {real, imag} */,
  {32'h40a1f602, 32'hc066fe50} /* (17, 27, 11) {real, imag} */,
  {32'h3f3d00b8, 32'hc1071dde} /* (17, 27, 10) {real, imag} */,
  {32'hc1300710, 32'hc1b1fbca} /* (17, 27, 9) {real, imag} */,
  {32'hc10ecbaa, 32'h40a18c51} /* (17, 27, 8) {real, imag} */,
  {32'h4167aa91, 32'hc1eaa384} /* (17, 27, 7) {real, imag} */,
  {32'h4218fdfe, 32'h42431e41} /* (17, 27, 6) {real, imag} */,
  {32'h41b71596, 32'h40084368} /* (17, 27, 5) {real, imag} */,
  {32'h41b6810c, 32'hc1077fe6} /* (17, 27, 4) {real, imag} */,
  {32'h4015b4a8, 32'hc26a615e} /* (17, 27, 3) {real, imag} */,
  {32'h414d6cfa, 32'hc1b1620d} /* (17, 27, 2) {real, imag} */,
  {32'h41ec2212, 32'h400c5356} /* (17, 27, 1) {real, imag} */,
  {32'h419cf64b, 32'h41e966fc} /* (17, 27, 0) {real, imag} */,
  {32'hc18dff4a, 32'hc1acde4d} /* (17, 26, 31) {real, imag} */,
  {32'h414d02ea, 32'h413938d0} /* (17, 26, 30) {real, imag} */,
  {32'h41953a10, 32'h4197e1b4} /* (17, 26, 29) {real, imag} */,
  {32'h4203c1b3, 32'hc029f8fe} /* (17, 26, 28) {real, imag} */,
  {32'hc13b55fe, 32'hc134ddd8} /* (17, 26, 27) {real, imag} */,
  {32'hc1b106be, 32'hc0040258} /* (17, 26, 26) {real, imag} */,
  {32'h409c0377, 32'h409762ae} /* (17, 26, 25) {real, imag} */,
  {32'hc260e66e, 32'h41b05446} /* (17, 26, 24) {real, imag} */,
  {32'hc06f4126, 32'h41d7c494} /* (17, 26, 23) {real, imag} */,
  {32'h3e9e7fc0, 32'hc1c58a0e} /* (17, 26, 22) {real, imag} */,
  {32'h4180f398, 32'hc07256c2} /* (17, 26, 21) {real, imag} */,
  {32'hc1334a23, 32'hc0084312} /* (17, 26, 20) {real, imag} */,
  {32'h40cc71cc, 32'hc102b224} /* (17, 26, 19) {real, imag} */,
  {32'h416c4c9c, 32'h41344d52} /* (17, 26, 18) {real, imag} */,
  {32'hbf03fbf2, 32'h3fb5e070} /* (17, 26, 17) {real, imag} */,
  {32'hc03a9b50, 32'h4045e57e} /* (17, 26, 16) {real, imag} */,
  {32'h3e39aa48, 32'hc0d787c4} /* (17, 26, 15) {real, imag} */,
  {32'h40e41189, 32'hc0a978c4} /* (17, 26, 14) {real, imag} */,
  {32'hbd1d6600, 32'h411b18d8} /* (17, 26, 13) {real, imag} */,
  {32'hc0119d7c, 32'h406104e2} /* (17, 26, 12) {real, imag} */,
  {32'h41000456, 32'hc112bf88} /* (17, 26, 11) {real, imag} */,
  {32'h41b8127f, 32'hc1a23ca2} /* (17, 26, 10) {real, imag} */,
  {32'hc16005bc, 32'h3f9bd448} /* (17, 26, 9) {real, imag} */,
  {32'hc034b998, 32'h418daa1e} /* (17, 26, 8) {real, imag} */,
  {32'hc08591cb, 32'hc17dad03} /* (17, 26, 7) {real, imag} */,
  {32'h423dadf1, 32'hbf9ddf80} /* (17, 26, 6) {real, imag} */,
  {32'h411f66f2, 32'h4221c100} /* (17, 26, 5) {real, imag} */,
  {32'h41bb9d46, 32'hc0f92619} /* (17, 26, 4) {real, imag} */,
  {32'h413f1131, 32'hc06a91ac} /* (17, 26, 3) {real, imag} */,
  {32'h40029c6a, 32'hc1d7e9ce} /* (17, 26, 2) {real, imag} */,
  {32'hc169af8c, 32'hc0e248cc} /* (17, 26, 1) {real, imag} */,
  {32'hc19b076e, 32'h4095f8ef} /* (17, 26, 0) {real, imag} */,
  {32'h40ebd674, 32'hc2161c40} /* (17, 25, 31) {real, imag} */,
  {32'h4238be99, 32'hc1b5097b} /* (17, 25, 30) {real, imag} */,
  {32'h412acfa6, 32'h40224268} /* (17, 25, 29) {real, imag} */,
  {32'h4164cc2b, 32'h42110a6d} /* (17, 25, 28) {real, imag} */,
  {32'h420fec58, 32'hbf9db0d0} /* (17, 25, 27) {real, imag} */,
  {32'hc202ec25, 32'hbfa30ad4} /* (17, 25, 26) {real, imag} */,
  {32'h3ea20010, 32'hc15de53f} /* (17, 25, 25) {real, imag} */,
  {32'hc12c932c, 32'h3f9efe60} /* (17, 25, 24) {real, imag} */,
  {32'h4198709e, 32'hc1356ede} /* (17, 25, 23) {real, imag} */,
  {32'h4127fbb9, 32'h41ac6c6e} /* (17, 25, 22) {real, imag} */,
  {32'h4085c0c4, 32'hc0fa40e3} /* (17, 25, 21) {real, imag} */,
  {32'hc055dfc9, 32'h4118fc7c} /* (17, 25, 20) {real, imag} */,
  {32'hbfbf8f44, 32'h3f515280} /* (17, 25, 19) {real, imag} */,
  {32'hc06567c8, 32'h407805d6} /* (17, 25, 18) {real, imag} */,
  {32'h409fa4ac, 32'h40028a0c} /* (17, 25, 17) {real, imag} */,
  {32'h3f399078, 32'hc00f79c0} /* (17, 25, 16) {real, imag} */,
  {32'h3f4c9b20, 32'h40e6da1a} /* (17, 25, 15) {real, imag} */,
  {32'h4043e398, 32'hc0873a1f} /* (17, 25, 14) {real, imag} */,
  {32'h41849b38, 32'hc1373ac4} /* (17, 25, 13) {real, imag} */,
  {32'h40ee0c3a, 32'h40523e32} /* (17, 25, 12) {real, imag} */,
  {32'h40893438, 32'hc17cf0aa} /* (17, 25, 11) {real, imag} */,
  {32'hc1a0c636, 32'hbfbc5ee0} /* (17, 25, 10) {real, imag} */,
  {32'hc0a3b319, 32'h41292504} /* (17, 25, 9) {real, imag} */,
  {32'hc0c2a40c, 32'h3f3e2810} /* (17, 25, 8) {real, imag} */,
  {32'hc0d3f0df, 32'h41ab6301} /* (17, 25, 7) {real, imag} */,
  {32'hc2181047, 32'hc0c97461} /* (17, 25, 6) {real, imag} */,
  {32'h409dde4e, 32'h3f5d3010} /* (17, 25, 5) {real, imag} */,
  {32'hc10fe179, 32'hc0c84ec8} /* (17, 25, 4) {real, imag} */,
  {32'hc08d659e, 32'h41934cd7} /* (17, 25, 3) {real, imag} */,
  {32'h41ed63f6, 32'hc1969601} /* (17, 25, 2) {real, imag} */,
  {32'hc1ce8ecd, 32'hc243b38a} /* (17, 25, 1) {real, imag} */,
  {32'hbf0fbb18, 32'hc17f60b0} /* (17, 25, 0) {real, imag} */,
  {32'hc22418d4, 32'h40f628e5} /* (17, 24, 31) {real, imag} */,
  {32'hc1528d7b, 32'h418c81e8} /* (17, 24, 30) {real, imag} */,
  {32'h4138d054, 32'hc10380f5} /* (17, 24, 29) {real, imag} */,
  {32'h421e4462, 32'h419f981d} /* (17, 24, 28) {real, imag} */,
  {32'h40c76d7e, 32'hc1548ac4} /* (17, 24, 27) {real, imag} */,
  {32'hbfaf6798, 32'h41b74079} /* (17, 24, 26) {real, imag} */,
  {32'hc1b9cb62, 32'hc1008718} /* (17, 24, 25) {real, imag} */,
  {32'hc0e2b65c, 32'hc175b060} /* (17, 24, 24) {real, imag} */,
  {32'hc102f645, 32'hc11babdc} /* (17, 24, 23) {real, imag} */,
  {32'h400111fc, 32'hc18e78a1} /* (17, 24, 22) {real, imag} */,
  {32'h408d74da, 32'h40e027d5} /* (17, 24, 21) {real, imag} */,
  {32'hc126b045, 32'hc0f10fac} /* (17, 24, 20) {real, imag} */,
  {32'h4075ceb4, 32'h40d42fde} /* (17, 24, 19) {real, imag} */,
  {32'h4112ee55, 32'h4031e48d} /* (17, 24, 18) {real, imag} */,
  {32'hc0156894, 32'hc0358e12} /* (17, 24, 17) {real, imag} */,
  {32'h40def9f4, 32'hc10c661a} /* (17, 24, 16) {real, imag} */,
  {32'hc02eb4a4, 32'hbf51db1e} /* (17, 24, 15) {real, imag} */,
  {32'h3e864860, 32'h405eec0d} /* (17, 24, 14) {real, imag} */,
  {32'hbfb05b10, 32'hbfcda9b6} /* (17, 24, 13) {real, imag} */,
  {32'h415a0145, 32'hc0a3b5fc} /* (17, 24, 12) {real, imag} */,
  {32'h40c0142e, 32'hc02a77aa} /* (17, 24, 11) {real, imag} */,
  {32'h41922848, 32'hc0dd5364} /* (17, 24, 10) {real, imag} */,
  {32'hc11dfeaf, 32'hc18e9e4c} /* (17, 24, 9) {real, imag} */,
  {32'hc115078a, 32'h41958126} /* (17, 24, 8) {real, imag} */,
  {32'hc1523057, 32'h4179f242} /* (17, 24, 7) {real, imag} */,
  {32'h41bed170, 32'hc19e27c5} /* (17, 24, 6) {real, imag} */,
  {32'h4151fa0f, 32'hc17d1794} /* (17, 24, 5) {real, imag} */,
  {32'h41b743ec, 32'hc2134666} /* (17, 24, 4) {real, imag} */,
  {32'h3f8a5598, 32'h41b8d5e2} /* (17, 24, 3) {real, imag} */,
  {32'hbe338c40, 32'h403fe330} /* (17, 24, 2) {real, imag} */,
  {32'h40c0147c, 32'h410472df} /* (17, 24, 1) {real, imag} */,
  {32'hc210fdca, 32'hbfa8f78c} /* (17, 24, 0) {real, imag} */,
  {32'h419ad64f, 32'hc1735024} /* (17, 23, 31) {real, imag} */,
  {32'h40edd4a8, 32'h41c124d2} /* (17, 23, 30) {real, imag} */,
  {32'h416cb420, 32'h414519fe} /* (17, 23, 29) {real, imag} */,
  {32'hc08f001d, 32'h419047eb} /* (17, 23, 28) {real, imag} */,
  {32'h3f5dc7b0, 32'h41236626} /* (17, 23, 27) {real, imag} */,
  {32'h41095fd3, 32'hc1fe1d78} /* (17, 23, 26) {real, imag} */,
  {32'h413332bf, 32'h401c427e} /* (17, 23, 25) {real, imag} */,
  {32'hc1b396ff, 32'h412e99ce} /* (17, 23, 24) {real, imag} */,
  {32'h412d3d2e, 32'hc1ac5179} /* (17, 23, 23) {real, imag} */,
  {32'h41f253e5, 32'h411402c3} /* (17, 23, 22) {real, imag} */,
  {32'hc0ec90f1, 32'h40b621b2} /* (17, 23, 21) {real, imag} */,
  {32'hc1345b68, 32'h405ac882} /* (17, 23, 20) {real, imag} */,
  {32'h402f6b2e, 32'hc0b634d4} /* (17, 23, 19) {real, imag} */,
  {32'hc0a07c24, 32'hc121f29b} /* (17, 23, 18) {real, imag} */,
  {32'hc0a7e33c, 32'h40aab2a7} /* (17, 23, 17) {real, imag} */,
  {32'hc08a0177, 32'h4029cfc9} /* (17, 23, 16) {real, imag} */,
  {32'hc051061c, 32'h401f463a} /* (17, 23, 15) {real, imag} */,
  {32'h3e5c41c0, 32'hc04b600b} /* (17, 23, 14) {real, imag} */,
  {32'hbf9120bc, 32'hc0420b0c} /* (17, 23, 13) {real, imag} */,
  {32'hbeb423d0, 32'hc0ec1d79} /* (17, 23, 12) {real, imag} */,
  {32'hc1930623, 32'hc10b66ac} /* (17, 23, 11) {real, imag} */,
  {32'h4187ee97, 32'h41a84bb2} /* (17, 23, 10) {real, imag} */,
  {32'h40cbe9f5, 32'hc11aaa5e} /* (17, 23, 9) {real, imag} */,
  {32'hc1b37fe9, 32'hc178333e} /* (17, 23, 8) {real, imag} */,
  {32'hc0a7a8e2, 32'hbef24770} /* (17, 23, 7) {real, imag} */,
  {32'h403dd8dc, 32'h40b94a0e} /* (17, 23, 6) {real, imag} */,
  {32'h41d0ace8, 32'hc0e97765} /* (17, 23, 5) {real, imag} */,
  {32'h3eae0190, 32'h41495b9a} /* (17, 23, 4) {real, imag} */,
  {32'hc0cf658f, 32'hc08f1bf3} /* (17, 23, 3) {real, imag} */,
  {32'h3f825288, 32'h411760a4} /* (17, 23, 2) {real, imag} */,
  {32'h3fbf4f90, 32'hc16696aa} /* (17, 23, 1) {real, imag} */,
  {32'h40aab087, 32'hbf74f050} /* (17, 23, 0) {real, imag} */,
  {32'hc11a2328, 32'hc0dd6659} /* (17, 22, 31) {real, imag} */,
  {32'h40081adc, 32'h411eea7e} /* (17, 22, 30) {real, imag} */,
  {32'h3ec91100, 32'h40c6f83c} /* (17, 22, 29) {real, imag} */,
  {32'hc0b9b534, 32'hc1b01eed} /* (17, 22, 28) {real, imag} */,
  {32'h40580328, 32'h4129e04c} /* (17, 22, 27) {real, imag} */,
  {32'h41441e7e, 32'hc178cd72} /* (17, 22, 26) {real, imag} */,
  {32'hc0e532eb, 32'hc08634cc} /* (17, 22, 25) {real, imag} */,
  {32'hc126218f, 32'hc0890ce9} /* (17, 22, 24) {real, imag} */,
  {32'h40fe433a, 32'h406a4732} /* (17, 22, 23) {real, imag} */,
  {32'hbf9cbe30, 32'hc1515d84} /* (17, 22, 22) {real, imag} */,
  {32'hc04c31a6, 32'hbf905730} /* (17, 22, 21) {real, imag} */,
  {32'hbfcf99ec, 32'hc0e72448} /* (17, 22, 20) {real, imag} */,
  {32'h408b28b2, 32'h410f1552} /* (17, 22, 19) {real, imag} */,
  {32'hc02e230a, 32'h4093db21} /* (17, 22, 18) {real, imag} */,
  {32'hc064fa80, 32'h3aafa000} /* (17, 22, 17) {real, imag} */,
  {32'h406c1904, 32'h4011887c} /* (17, 22, 16) {real, imag} */,
  {32'hc086e2f1, 32'hbfa404f8} /* (17, 22, 15) {real, imag} */,
  {32'hc09297f7, 32'hc0062266} /* (17, 22, 14) {real, imag} */,
  {32'h4052e6f8, 32'h3f631700} /* (17, 22, 13) {real, imag} */,
  {32'h40cc2659, 32'hc0b7c0dc} /* (17, 22, 12) {real, imag} */,
  {32'h3f46a52e, 32'hbf2df840} /* (17, 22, 11) {real, imag} */,
  {32'hc1a88363, 32'h40c42463} /* (17, 22, 10) {real, imag} */,
  {32'h413a5cad, 32'h41927758} /* (17, 22, 9) {real, imag} */,
  {32'hc0b005ce, 32'hc0bb27ff} /* (17, 22, 8) {real, imag} */,
  {32'hc100b448, 32'h41a24bc5} /* (17, 22, 7) {real, imag} */,
  {32'h407d38b8, 32'hc141e89a} /* (17, 22, 6) {real, imag} */,
  {32'h4081bed4, 32'hc18da79b} /* (17, 22, 5) {real, imag} */,
  {32'h4000aaab, 32'hc0d65818} /* (17, 22, 4) {real, imag} */,
  {32'hc0b495a2, 32'h40f0be48} /* (17, 22, 3) {real, imag} */,
  {32'h41c091b4, 32'h4115d072} /* (17, 22, 2) {real, imag} */,
  {32'h4092f1f8, 32'hc15db832} /* (17, 22, 1) {real, imag} */,
  {32'hc1534347, 32'h3f140369} /* (17, 22, 0) {real, imag} */,
  {32'h414a1a09, 32'hc0aa126e} /* (17, 21, 31) {real, imag} */,
  {32'h4047bc5c, 32'hc029d754} /* (17, 21, 30) {real, imag} */,
  {32'hbddd1040, 32'h40f3d840} /* (17, 21, 29) {real, imag} */,
  {32'hc118f0b0, 32'h4196e1a0} /* (17, 21, 28) {real, imag} */,
  {32'h4186364c, 32'h4115dbe2} /* (17, 21, 27) {real, imag} */,
  {32'h41641e3e, 32'hc0571546} /* (17, 21, 26) {real, imag} */,
  {32'h4137bb5c, 32'hc005fd55} /* (17, 21, 25) {real, imag} */,
  {32'hc16cdf14, 32'h414f5e60} /* (17, 21, 24) {real, imag} */,
  {32'h410ff8a1, 32'h3faae68e} /* (17, 21, 23) {real, imag} */,
  {32'hbeaf66a0, 32'hc00d9fe2} /* (17, 21, 22) {real, imag} */,
  {32'hbf91d7c4, 32'hbf0a678c} /* (17, 21, 21) {real, imag} */,
  {32'hc09574b2, 32'hc11538d8} /* (17, 21, 20) {real, imag} */,
  {32'h400dc297, 32'h4000ce51} /* (17, 21, 19) {real, imag} */,
  {32'h4067fe98, 32'h3d523980} /* (17, 21, 18) {real, imag} */,
  {32'h3f827380, 32'h3f2cffbc} /* (17, 21, 17) {real, imag} */,
  {32'h4084ffc4, 32'h40c87aa7} /* (17, 21, 16) {real, imag} */,
  {32'h3efa5540, 32'h40289721} /* (17, 21, 15) {real, imag} */,
  {32'h3fccbce8, 32'h3edcb930} /* (17, 21, 14) {real, imag} */,
  {32'hbfe499ca, 32'hc10d36d5} /* (17, 21, 13) {real, imag} */,
  {32'h40a2d600, 32'h3f817254} /* (17, 21, 12) {real, imag} */,
  {32'hc0bb3a81, 32'h3f80de3e} /* (17, 21, 11) {real, imag} */,
  {32'hc153985e, 32'h3eedda4a} /* (17, 21, 10) {real, imag} */,
  {32'hc11f4d93, 32'hc0d07df8} /* (17, 21, 9) {real, imag} */,
  {32'hc03ada6e, 32'hc11fb3f2} /* (17, 21, 8) {real, imag} */,
  {32'h4174e2f2, 32'h40b762ee} /* (17, 21, 7) {real, imag} */,
  {32'hc046e69a, 32'hbed1aed4} /* (17, 21, 6) {real, imag} */,
  {32'hc0ba78d1, 32'h3e0353e0} /* (17, 21, 5) {real, imag} */,
  {32'hc150a06c, 32'h3ff3dc38} /* (17, 21, 4) {real, imag} */,
  {32'h4140c32c, 32'hc14f7738} /* (17, 21, 3) {real, imag} */,
  {32'h3febae11, 32'h40d5d1da} /* (17, 21, 2) {real, imag} */,
  {32'hbf8ad5f8, 32'hc16b9aa5} /* (17, 21, 1) {real, imag} */,
  {32'h40bc15c4, 32'hc151c4e4} /* (17, 21, 0) {real, imag} */,
  {32'h41269e82, 32'h405f5138} /* (17, 20, 31) {real, imag} */,
  {32'h41686beb, 32'h411d7a3c} /* (17, 20, 30) {real, imag} */,
  {32'h40b2573c, 32'hbee77940} /* (17, 20, 29) {real, imag} */,
  {32'hc12edad2, 32'h40c04a91} /* (17, 20, 28) {real, imag} */,
  {32'hc124743d, 32'h408f3774} /* (17, 20, 27) {real, imag} */,
  {32'h40a22592, 32'hbfeeb7ea} /* (17, 20, 26) {real, imag} */,
  {32'hc0fe0c8b, 32'h409d3a41} /* (17, 20, 25) {real, imag} */,
  {32'h41110df0, 32'h40075130} /* (17, 20, 24) {real, imag} */,
  {32'hc0b036fa, 32'hc09f34cd} /* (17, 20, 23) {real, imag} */,
  {32'hc0f4981e, 32'h4096240d} /* (17, 20, 22) {real, imag} */,
  {32'hbee9a1b8, 32'hc0045543} /* (17, 20, 21) {real, imag} */,
  {32'hbe1c8b88, 32'hc047cdae} /* (17, 20, 20) {real, imag} */,
  {32'h3e2512f0, 32'h3ecb8188} /* (17, 20, 19) {real, imag} */,
  {32'hc04b4441, 32'hbfd1a44c} /* (17, 20, 18) {real, imag} */,
  {32'hbf1a9b90, 32'h3ed0c290} /* (17, 20, 17) {real, imag} */,
  {32'hbfc4a72c, 32'hc043971e} /* (17, 20, 16) {real, imag} */,
  {32'h3dd37580, 32'hc0f6f35f} /* (17, 20, 15) {real, imag} */,
  {32'hc05bc15b, 32'h3cdfe300} /* (17, 20, 14) {real, imag} */,
  {32'hc026f219, 32'hc052352f} /* (17, 20, 13) {real, imag} */,
  {32'h40580a60, 32'h4100f72e} /* (17, 20, 12) {real, imag} */,
  {32'hbfd45fde, 32'hc080330e} /* (17, 20, 11) {real, imag} */,
  {32'h40fa0baa, 32'hc0820c03} /* (17, 20, 10) {real, imag} */,
  {32'h40b0eca2, 32'h40d3228b} /* (17, 20, 9) {real, imag} */,
  {32'hc004bd5a, 32'hc11d393d} /* (17, 20, 8) {real, imag} */,
  {32'hc093f9b9, 32'h40ec2209} /* (17, 20, 7) {real, imag} */,
  {32'h410e056d, 32'hbed0a268} /* (17, 20, 6) {real, imag} */,
  {32'h41940d62, 32'hc0acd334} /* (17, 20, 5) {real, imag} */,
  {32'h40a2b800, 32'hc0d2fead} /* (17, 20, 4) {real, imag} */,
  {32'hc0964508, 32'h4142716e} /* (17, 20, 3) {real, imag} */,
  {32'h410ccbe9, 32'h4001f282} /* (17, 20, 2) {real, imag} */,
  {32'h41f319ab, 32'h3f1c7280} /* (17, 20, 1) {real, imag} */,
  {32'hc1881fa9, 32'hc131c26c} /* (17, 20, 0) {real, imag} */,
  {32'hc159559d, 32'hbf10f290} /* (17, 19, 31) {real, imag} */,
  {32'hc1e3c120, 32'hc02986a4} /* (17, 19, 30) {real, imag} */,
  {32'h40c6242f, 32'h40516406} /* (17, 19, 29) {real, imag} */,
  {32'hbed40ae0, 32'h412da23a} /* (17, 19, 28) {real, imag} */,
  {32'h3ec68ba4, 32'hc0bd3f3e} /* (17, 19, 27) {real, imag} */,
  {32'h40b45a58, 32'h41458e3d} /* (17, 19, 26) {real, imag} */,
  {32'hc03889cf, 32'h404867ec} /* (17, 19, 25) {real, imag} */,
  {32'hc0544af5, 32'hc1034fbe} /* (17, 19, 24) {real, imag} */,
  {32'h41065441, 32'h410318f8} /* (17, 19, 23) {real, imag} */,
  {32'hc067dfb9, 32'hbfaa2f5c} /* (17, 19, 22) {real, imag} */,
  {32'h40a891cc, 32'h40536f91} /* (17, 19, 21) {real, imag} */,
  {32'hc0ca6f68, 32'hc0146cbc} /* (17, 19, 20) {real, imag} */,
  {32'hc0a1bd06, 32'hc01bd7e0} /* (17, 19, 19) {real, imag} */,
  {32'hbfb55f58, 32'hc0c70855} /* (17, 19, 18) {real, imag} */,
  {32'h40b53fdf, 32'h400c9830} /* (17, 19, 17) {real, imag} */,
  {32'h3fb0a4bc, 32'hbe559b20} /* (17, 19, 16) {real, imag} */,
  {32'hbfc80a3c, 32'hc030d76c} /* (17, 19, 15) {real, imag} */,
  {32'hbe2cc080, 32'hc09b7817} /* (17, 19, 14) {real, imag} */,
  {32'hc0a1b610, 32'h401db244} /* (17, 19, 13) {real, imag} */,
  {32'hbff07e88, 32'hc00e34aa} /* (17, 19, 12) {real, imag} */,
  {32'hc07aa538, 32'h3f7fda1c} /* (17, 19, 11) {real, imag} */,
  {32'h3fa61d82, 32'h40cd9171} /* (17, 19, 10) {real, imag} */,
  {32'hc113c685, 32'h3fcec384} /* (17, 19, 9) {real, imag} */,
  {32'hbf5d053c, 32'hc0e68f3b} /* (17, 19, 8) {real, imag} */,
  {32'hc0abd664, 32'hc03b48e4} /* (17, 19, 7) {real, imag} */,
  {32'h4094edac, 32'h4088086e} /* (17, 19, 6) {real, imag} */,
  {32'h403d6996, 32'h40a21b9e} /* (17, 19, 5) {real, imag} */,
  {32'h414aa0d2, 32'hc008dcc0} /* (17, 19, 4) {real, imag} */,
  {32'h3d1db980, 32'h410b66ec} /* (17, 19, 3) {real, imag} */,
  {32'h3fc14980, 32'h41737f57} /* (17, 19, 2) {real, imag} */,
  {32'hc13b4c4f, 32'hc0c355d4} /* (17, 19, 1) {real, imag} */,
  {32'h404785c6, 32'hc10d2e44} /* (17, 19, 0) {real, imag} */,
  {32'h408dea9b, 32'hbf25b1c4} /* (17, 18, 31) {real, imag} */,
  {32'hc140a308, 32'hbf3c58b0} /* (17, 18, 30) {real, imag} */,
  {32'hc1767073, 32'h3fad5106} /* (17, 18, 29) {real, imag} */,
  {32'h40bb77d2, 32'h410d38a7} /* (17, 18, 28) {real, imag} */,
  {32'hc0616ef0, 32'h41539c01} /* (17, 18, 27) {real, imag} */,
  {32'hbf84262a, 32'hc01d5f3a} /* (17, 18, 26) {real, imag} */,
  {32'h402d4b41, 32'h4053a480} /* (17, 18, 25) {real, imag} */,
  {32'h3e4bc220, 32'h404cdb96} /* (17, 18, 24) {real, imag} */,
  {32'h40affc84, 32'hc1142e74} /* (17, 18, 23) {real, imag} */,
  {32'hc046e41e, 32'hc08d64e6} /* (17, 18, 22) {real, imag} */,
  {32'hc035ba7a, 32'h402eaef9} /* (17, 18, 21) {real, imag} */,
  {32'h4078b120, 32'h3fe0e75a} /* (17, 18, 20) {real, imag} */,
  {32'h3f48585c, 32'hc017f613} /* (17, 18, 19) {real, imag} */,
  {32'hbfaa9998, 32'hbfaee6e8} /* (17, 18, 18) {real, imag} */,
  {32'h3fd23beb, 32'h3fac5c42} /* (17, 18, 17) {real, imag} */,
  {32'hbff461cc, 32'h4098a922} /* (17, 18, 16) {real, imag} */,
  {32'hbfee9d3d, 32'h3f8faf8e} /* (17, 18, 15) {real, imag} */,
  {32'hbf0f3498, 32'hc07b46b4} /* (17, 18, 14) {real, imag} */,
  {32'hbf118e54, 32'h403f6031} /* (17, 18, 13) {real, imag} */,
  {32'hc084b930, 32'h3f956492} /* (17, 18, 12) {real, imag} */,
  {32'hbf4b0756, 32'hbe3ae910} /* (17, 18, 11) {real, imag} */,
  {32'hbf6ed842, 32'h3fdf8a81} /* (17, 18, 10) {real, imag} */,
  {32'h40d295d8, 32'h3dff7b00} /* (17, 18, 9) {real, imag} */,
  {32'h3d4c3f00, 32'hc0fa2e7f} /* (17, 18, 8) {real, imag} */,
  {32'hc0e1ca20, 32'h40a54cac} /* (17, 18, 7) {real, imag} */,
  {32'hc0a2c1fe, 32'h40d5b55f} /* (17, 18, 6) {real, imag} */,
  {32'h404537ec, 32'h4152f985} /* (17, 18, 5) {real, imag} */,
  {32'hbfa6e180, 32'hc0bfc562} /* (17, 18, 4) {real, imag} */,
  {32'h40b378f2, 32'h402572db} /* (17, 18, 3) {real, imag} */,
  {32'hc01b3b80, 32'hc185be9a} /* (17, 18, 2) {real, imag} */,
  {32'h3f5bfd58, 32'hc04fa6a7} /* (17, 18, 1) {real, imag} */,
  {32'h413b8b06, 32'h4182a1ba} /* (17, 18, 0) {real, imag} */,
  {32'hbffdf6ba, 32'hc1009bd4} /* (17, 17, 31) {real, imag} */,
  {32'hc0a67f2c, 32'hc09c316f} /* (17, 17, 30) {real, imag} */,
  {32'hbf0fd9e8, 32'h3f92467c} /* (17, 17, 29) {real, imag} */,
  {32'h403591fd, 32'h3c95f000} /* (17, 17, 28) {real, imag} */,
  {32'h40874fd4, 32'h410c567e} /* (17, 17, 27) {real, imag} */,
  {32'h4034da2e, 32'hc1521087} /* (17, 17, 26) {real, imag} */,
  {32'hbff42824, 32'h402aa355} /* (17, 17, 25) {real, imag} */,
  {32'h3f5d6d9a, 32'h4046871e} /* (17, 17, 24) {real, imag} */,
  {32'hbf9d745a, 32'hbff2c91e} /* (17, 17, 23) {real, imag} */,
  {32'h40cf0fd6, 32'hc0a68552} /* (17, 17, 22) {real, imag} */,
  {32'hc07ab32a, 32'hc02f0866} /* (17, 17, 21) {real, imag} */,
  {32'h408aa7ee, 32'hc08626c4} /* (17, 17, 20) {real, imag} */,
  {32'h3fae2386, 32'hbfa83b08} /* (17, 17, 19) {real, imag} */,
  {32'h402037ce, 32'h3fc187f3} /* (17, 17, 18) {real, imag} */,
  {32'h3f5f2fd2, 32'hc05ec708} /* (17, 17, 17) {real, imag} */,
  {32'h3f04aada, 32'h3da70390} /* (17, 17, 16) {real, imag} */,
  {32'h3f8342dd, 32'h3f92db0b} /* (17, 17, 15) {real, imag} */,
  {32'h3f6c9010, 32'hc0536822} /* (17, 17, 14) {real, imag} */,
  {32'h3f783d0c, 32'hbfcbc8d8} /* (17, 17, 13) {real, imag} */,
  {32'h40899fb0, 32'h3fa20859} /* (17, 17, 12) {real, imag} */,
  {32'hc073d6aa, 32'h408f2006} /* (17, 17, 11) {real, imag} */,
  {32'hc0544bf9, 32'h3f8d7738} /* (17, 17, 10) {real, imag} */,
  {32'h3f141f44, 32'hc05b322f} /* (17, 17, 9) {real, imag} */,
  {32'h3fafacb3, 32'h407aa89a} /* (17, 17, 8) {real, imag} */,
  {32'h40c07fa0, 32'hc109f24c} /* (17, 17, 7) {real, imag} */,
  {32'hbfe52c74, 32'hc0630084} /* (17, 17, 6) {real, imag} */,
  {32'h4103ffb5, 32'hc0bfeaf7} /* (17, 17, 5) {real, imag} */,
  {32'h4053b7e3, 32'h40a9ad82} /* (17, 17, 4) {real, imag} */,
  {32'h4081e70f, 32'hc092940d} /* (17, 17, 3) {real, imag} */,
  {32'hbf179358, 32'hbf8f928b} /* (17, 17, 2) {real, imag} */,
  {32'hbfb90338, 32'h409cf01f} /* (17, 17, 1) {real, imag} */,
  {32'hbfc4d5f5, 32'h404e0c4c} /* (17, 17, 0) {real, imag} */,
  {32'h4072de22, 32'hc0862dc2} /* (17, 16, 31) {real, imag} */,
  {32'h40497eb4, 32'hc0ab11a0} /* (17, 16, 30) {real, imag} */,
  {32'h4002fc19, 32'h412b8318} /* (17, 16, 29) {real, imag} */,
  {32'h4000eeca, 32'hc0729a01} /* (17, 16, 28) {real, imag} */,
  {32'h40f09a2a, 32'hc12d740a} /* (17, 16, 27) {real, imag} */,
  {32'h40eeab40, 32'h3fb67866} /* (17, 16, 26) {real, imag} */,
  {32'hc01cc458, 32'h4074730a} /* (17, 16, 25) {real, imag} */,
  {32'h40de7adf, 32'h4011b1f4} /* (17, 16, 24) {real, imag} */,
  {32'hc0985777, 32'hbfb8910c} /* (17, 16, 23) {real, imag} */,
  {32'h40012270, 32'hc115ab0c} /* (17, 16, 22) {real, imag} */,
  {32'h3fa40ee4, 32'h40fd03c1} /* (17, 16, 21) {real, imag} */,
  {32'hc02f8352, 32'h404f514e} /* (17, 16, 20) {real, imag} */,
  {32'hc03f1d66, 32'h3fdc6c28} /* (17, 16, 19) {real, imag} */,
  {32'hc0286602, 32'hc0445d32} /* (17, 16, 18) {real, imag} */,
  {32'hbf369a0c, 32'h3e5e1ef8} /* (17, 16, 17) {real, imag} */,
  {32'h3f5f4498, 32'hbe5aae10} /* (17, 16, 16) {real, imag} */,
  {32'hbf40b66c, 32'hbe3dcae8} /* (17, 16, 15) {real, imag} */,
  {32'hbf1be3ae, 32'hbefe83cc} /* (17, 16, 14) {real, imag} */,
  {32'h4047c620, 32'h402da9c0} /* (17, 16, 13) {real, imag} */,
  {32'h3fe0dda5, 32'hc005a646} /* (17, 16, 12) {real, imag} */,
  {32'hbfa161e4, 32'hbebaa8b0} /* (17, 16, 11) {real, imag} */,
  {32'h412ca1ea, 32'h40c74f42} /* (17, 16, 10) {real, imag} */,
  {32'hbe72d760, 32'h411f6176} /* (17, 16, 9) {real, imag} */,
  {32'hc08bc24d, 32'h408310a4} /* (17, 16, 8) {real, imag} */,
  {32'hc090cc36, 32'hbe8423cc} /* (17, 16, 7) {real, imag} */,
  {32'hc08b3cf4, 32'hc0e75c10} /* (17, 16, 6) {real, imag} */,
  {32'hc0749aaf, 32'h40b5482f} /* (17, 16, 5) {real, imag} */,
  {32'hc107d0a8, 32'h40b45150} /* (17, 16, 4) {real, imag} */,
  {32'hc068b4d1, 32'h41361be0} /* (17, 16, 3) {real, imag} */,
  {32'hbfe82fd7, 32'h3fdd02ef} /* (17, 16, 2) {real, imag} */,
  {32'hc10c98be, 32'h3dbf9680} /* (17, 16, 1) {real, imag} */,
  {32'h4005e3f9, 32'hc092a30a} /* (17, 16, 0) {real, imag} */,
  {32'h40ad6f9b, 32'hc13cda9e} /* (17, 15, 31) {real, imag} */,
  {32'hc07c0806, 32'h3fe24975} /* (17, 15, 30) {real, imag} */,
  {32'h409c2837, 32'h3eaa9610} /* (17, 15, 29) {real, imag} */,
  {32'hbfdb1f72, 32'hbf689278} /* (17, 15, 28) {real, imag} */,
  {32'h3e64c793, 32'h3fa98d5a} /* (17, 15, 27) {real, imag} */,
  {32'h4084164e, 32'h3fd7c90c} /* (17, 15, 26) {real, imag} */,
  {32'hc12c7cb8, 32'h3fe4e752} /* (17, 15, 25) {real, imag} */,
  {32'hbfccfabb, 32'h3fd02244} /* (17, 15, 24) {real, imag} */,
  {32'hbff101bc, 32'h3fd20a3e} /* (17, 15, 23) {real, imag} */,
  {32'hc0dec768, 32'hbfabb7b4} /* (17, 15, 22) {real, imag} */,
  {32'hc0194324, 32'h3f89c484} /* (17, 15, 21) {real, imag} */,
  {32'h4109914b, 32'hc05f3c30} /* (17, 15, 20) {real, imag} */,
  {32'h3ff272de, 32'hc05f5dae} /* (17, 15, 19) {real, imag} */,
  {32'h40051822, 32'h3eb238d4} /* (17, 15, 18) {real, imag} */,
  {32'h4022d08c, 32'h3f82f522} /* (17, 15, 17) {real, imag} */,
  {32'h40134f2c, 32'h3f346b10} /* (17, 15, 16) {real, imag} */,
  {32'h3f84a017, 32'h3f84716e} /* (17, 15, 15) {real, imag} */,
  {32'hc06597ae, 32'h3f2ca10e} /* (17, 15, 14) {real, imag} */,
  {32'hbeb856f6, 32'h3f0b701a} /* (17, 15, 13) {real, imag} */,
  {32'hbfea5e88, 32'hbf6fbbe0} /* (17, 15, 12) {real, imag} */,
  {32'hbfc50878, 32'hbf9f7790} /* (17, 15, 11) {real, imag} */,
  {32'hbef9d098, 32'hc1035078} /* (17, 15, 10) {real, imag} */,
  {32'hc101efac, 32'hbf36f47c} /* (17, 15, 9) {real, imag} */,
  {32'h3e5798e8, 32'h40bc46eb} /* (17, 15, 8) {real, imag} */,
  {32'hbefd6370, 32'hc0a023a4} /* (17, 15, 7) {real, imag} */,
  {32'h40299dc9, 32'hc04ca372} /* (17, 15, 6) {real, imag} */,
  {32'h3eadfe5a, 32'h40faa9d6} /* (17, 15, 5) {real, imag} */,
  {32'hbdda24e0, 32'h405cfac6} /* (17, 15, 4) {real, imag} */,
  {32'h3ef6a490, 32'hc0a3e25d} /* (17, 15, 3) {real, imag} */,
  {32'h40b2369d, 32'hbf713e7a} /* (17, 15, 2) {real, imag} */,
  {32'hc0bae42d, 32'hc1167908} /* (17, 15, 1) {real, imag} */,
  {32'hbf1bb390, 32'hc10fdfbc} /* (17, 15, 0) {real, imag} */,
  {32'h4178aa4f, 32'hc0be1b36} /* (17, 14, 31) {real, imag} */,
  {32'h413debc6, 32'h40a09a96} /* (17, 14, 30) {real, imag} */,
  {32'hc0d3f2ca, 32'h40dc3a55} /* (17, 14, 29) {real, imag} */,
  {32'hbf512cf0, 32'h40dae5f8} /* (17, 14, 28) {real, imag} */,
  {32'h41576054, 32'hc0fdbd9b} /* (17, 14, 27) {real, imag} */,
  {32'h40b05d38, 32'h412b407e} /* (17, 14, 26) {real, imag} */,
  {32'h414b6070, 32'h4119c908} /* (17, 14, 25) {real, imag} */,
  {32'h3eb297b8, 32'h40aed2b8} /* (17, 14, 24) {real, imag} */,
  {32'hc08a2b20, 32'h40a1a2ef} /* (17, 14, 23) {real, imag} */,
  {32'h3ff6acbd, 32'h40dc22be} /* (17, 14, 22) {real, imag} */,
  {32'h3f022cf0, 32'h40dabce3} /* (17, 14, 21) {real, imag} */,
  {32'h3f153d88, 32'h3e7da9c0} /* (17, 14, 20) {real, imag} */,
  {32'hbf890a96, 32'hbeb0d220} /* (17, 14, 19) {real, imag} */,
  {32'hbfec72c1, 32'hc01366ac} /* (17, 14, 18) {real, imag} */,
  {32'h3fba7bb8, 32'hbf59f9ec} /* (17, 14, 17) {real, imag} */,
  {32'hbff4173c, 32'h3f992676} /* (17, 14, 16) {real, imag} */,
  {32'hc0bda902, 32'hc02da07f} /* (17, 14, 15) {real, imag} */,
  {32'h3ff0c539, 32'h3f33b07a} /* (17, 14, 14) {real, imag} */,
  {32'hc0e0e024, 32'hc06d10fc} /* (17, 14, 13) {real, imag} */,
  {32'hbed1eb60, 32'hc0b6077a} /* (17, 14, 12) {real, imag} */,
  {32'h40b368d7, 32'hc0085022} /* (17, 14, 11) {real, imag} */,
  {32'hbf45b102, 32'h408a93c6} /* (17, 14, 10) {real, imag} */,
  {32'hc00050bf, 32'h3f77b240} /* (17, 14, 9) {real, imag} */,
  {32'h409b878a, 32'h40b7b1dc} /* (17, 14, 8) {real, imag} */,
  {32'h4186b59a, 32'hbeb1d800} /* (17, 14, 7) {real, imag} */,
  {32'h412c52b4, 32'hbfd536c0} /* (17, 14, 6) {real, imag} */,
  {32'h40032cc0, 32'hc0420812} /* (17, 14, 5) {real, imag} */,
  {32'h41210ccb, 32'hc11df6ae} /* (17, 14, 4) {real, imag} */,
  {32'hbfa42044, 32'hbfcca574} /* (17, 14, 3) {real, imag} */,
  {32'h4135d21a, 32'hc08e3c6e} /* (17, 14, 2) {real, imag} */,
  {32'h3fe25118, 32'hbf2cfaa4} /* (17, 14, 1) {real, imag} */,
  {32'h3d93d598, 32'h40eff366} /* (17, 14, 0) {real, imag} */,
  {32'h40bbb3d5, 32'h404e4fdd} /* (17, 13, 31) {real, imag} */,
  {32'hc110097e, 32'hc0a05338} /* (17, 13, 30) {real, imag} */,
  {32'hc10d8946, 32'hc0b893b8} /* (17, 13, 29) {real, imag} */,
  {32'hc0915716, 32'hc15c8e66} /* (17, 13, 28) {real, imag} */,
  {32'h4095197a, 32'h41402e22} /* (17, 13, 27) {real, imag} */,
  {32'h40131171, 32'hbfe615d0} /* (17, 13, 26) {real, imag} */,
  {32'h40a9d8a0, 32'h3fc4869f} /* (17, 13, 25) {real, imag} */,
  {32'h410b27b5, 32'hc0d9ec70} /* (17, 13, 24) {real, imag} */,
  {32'h408840e2, 32'hc039576c} /* (17, 13, 23) {real, imag} */,
  {32'h3fffad60, 32'hc111b793} /* (17, 13, 22) {real, imag} */,
  {32'h407a70d8, 32'h3e985694} /* (17, 13, 21) {real, imag} */,
  {32'h3d1eabf0, 32'hc00e9250} /* (17, 13, 20) {real, imag} */,
  {32'hc0a2b6da, 32'h4102a52a} /* (17, 13, 19) {real, imag} */,
  {32'hc0292892, 32'h3ff61718} /* (17, 13, 18) {real, imag} */,
  {32'hc09dc075, 32'h4001d056} /* (17, 13, 17) {real, imag} */,
  {32'h3f39c920, 32'h3f445c58} /* (17, 13, 16) {real, imag} */,
  {32'h4043fe86, 32'hc02f7fe4} /* (17, 13, 15) {real, imag} */,
  {32'hc0a24aea, 32'hc0843535} /* (17, 13, 14) {real, imag} */,
  {32'h3f251f34, 32'h3ff46b84} /* (17, 13, 13) {real, imag} */,
  {32'hbf707c87, 32'hc0d33fb0} /* (17, 13, 12) {real, imag} */,
  {32'hbfd59a10, 32'hc0295666} /* (17, 13, 11) {real, imag} */,
  {32'hbfc44480, 32'hc04b9454} /* (17, 13, 10) {real, imag} */,
  {32'hc0bc329a, 32'h3f427846} /* (17, 13, 9) {real, imag} */,
  {32'h4103d429, 32'h403bfcd0} /* (17, 13, 8) {real, imag} */,
  {32'h4091e9d0, 32'h3fbf4295} /* (17, 13, 7) {real, imag} */,
  {32'h4055e3b3, 32'hc186a049} /* (17, 13, 6) {real, imag} */,
  {32'hbfb7b036, 32'hc0cc6d40} /* (17, 13, 5) {real, imag} */,
  {32'hbd8f4ec0, 32'hc1213d06} /* (17, 13, 4) {real, imag} */,
  {32'hc03040ca, 32'h41098d4f} /* (17, 13, 3) {real, imag} */,
  {32'h40aa2494, 32'h417d310c} /* (17, 13, 2) {real, imag} */,
  {32'h415c23de, 32'h40ebd156} /* (17, 13, 1) {real, imag} */,
  {32'hbfee2104, 32'hc0626a8e} /* (17, 13, 0) {real, imag} */,
  {32'hc12f4f97, 32'h4161ed7d} /* (17, 12, 31) {real, imag} */,
  {32'hc1381674, 32'h40d1d6e8} /* (17, 12, 30) {real, imag} */,
  {32'hc0dcc8d1, 32'hbff4a1ab} /* (17, 12, 29) {real, imag} */,
  {32'hc10f2d26, 32'h4129463e} /* (17, 12, 28) {real, imag} */,
  {32'hc1217ab6, 32'hc139d070} /* (17, 12, 27) {real, imag} */,
  {32'h40e230f9, 32'hc0225045} /* (17, 12, 26) {real, imag} */,
  {32'hc0e8bce0, 32'hbf3c9638} /* (17, 12, 25) {real, imag} */,
  {32'hc0cf3d06, 32'hbee9a6c0} /* (17, 12, 24) {real, imag} */,
  {32'hbbb63a00, 32'hc0f1f2bf} /* (17, 12, 23) {real, imag} */,
  {32'h4072b480, 32'hc0b03212} /* (17, 12, 22) {real, imag} */,
  {32'h4116b410, 32'hc042034a} /* (17, 12, 21) {real, imag} */,
  {32'hc1501716, 32'h4083ce94} /* (17, 12, 20) {real, imag} */,
  {32'h405b24e2, 32'hc02fc9ca} /* (17, 12, 19) {real, imag} */,
  {32'h409c568b, 32'hc09d8b7d} /* (17, 12, 18) {real, imag} */,
  {32'h3fec863e, 32'hbf9518fd} /* (17, 12, 17) {real, imag} */,
  {32'h405eff31, 32'h40182e24} /* (17, 12, 16) {real, imag} */,
  {32'h3ff23eb2, 32'h40a45db5} /* (17, 12, 15) {real, imag} */,
  {32'h40a4d367, 32'h3ff56908} /* (17, 12, 14) {real, imag} */,
  {32'hbf851041, 32'h408b16aa} /* (17, 12, 13) {real, imag} */,
  {32'h3fddf820, 32'hc0e71742} /* (17, 12, 12) {real, imag} */,
  {32'h3fbf423c, 32'h3eb9d054} /* (17, 12, 11) {real, imag} */,
  {32'h40b3d58c, 32'hc04ce943} /* (17, 12, 10) {real, imag} */,
  {32'h4065ecbf, 32'hc130795a} /* (17, 12, 9) {real, imag} */,
  {32'h416ce63d, 32'hc13b6a52} /* (17, 12, 8) {real, imag} */,
  {32'hc096dbbc, 32'h412f2e9c} /* (17, 12, 7) {real, imag} */,
  {32'hbfa0d1d4, 32'h408e2848} /* (17, 12, 6) {real, imag} */,
  {32'hc02a9a58, 32'hc0e974e0} /* (17, 12, 5) {real, imag} */,
  {32'h4107ae24, 32'h415e0e16} /* (17, 12, 4) {real, imag} */,
  {32'h40b03c37, 32'h408455d6} /* (17, 12, 3) {real, imag} */,
  {32'h41803be3, 32'h40ff1044} /* (17, 12, 2) {real, imag} */,
  {32'hc1321773, 32'hc13077ff} /* (17, 12, 1) {real, imag} */,
  {32'h40a96a6c, 32'hc0fa78ba} /* (17, 12, 0) {real, imag} */,
  {32'h4081dd97, 32'h410e7dc0} /* (17, 11, 31) {real, imag} */,
  {32'h413ac3b6, 32'h4215962f} /* (17, 11, 30) {real, imag} */,
  {32'h4077802f, 32'h407ea009} /* (17, 11, 29) {real, imag} */,
  {32'h40a66d8c, 32'hc113dba7} /* (17, 11, 28) {real, imag} */,
  {32'hc088919f, 32'h4183a56e} /* (17, 11, 27) {real, imag} */,
  {32'hc1766694, 32'h40ea9d76} /* (17, 11, 26) {real, imag} */,
  {32'hc0d171b0, 32'hc0e5ab17} /* (17, 11, 25) {real, imag} */,
  {32'hbfaff020, 32'h40d4cf12} /* (17, 11, 24) {real, imag} */,
  {32'hc0d96c32, 32'hc1528fcb} /* (17, 11, 23) {real, imag} */,
  {32'h410157f4, 32'hbfc8dd2e} /* (17, 11, 22) {real, imag} */,
  {32'hc04be066, 32'h40eef24e} /* (17, 11, 21) {real, imag} */,
  {32'h41014a0e, 32'hbff0c678} /* (17, 11, 20) {real, imag} */,
  {32'hc0eb0a50, 32'hc056e1c9} /* (17, 11, 19) {real, imag} */,
  {32'hbf3b5abc, 32'hbf5c2f18} /* (17, 11, 18) {real, imag} */,
  {32'hc073b1c0, 32'h3f971360} /* (17, 11, 17) {real, imag} */,
  {32'hc0597ddc, 32'h403fe38c} /* (17, 11, 16) {real, imag} */,
  {32'h40798ffc, 32'h40842056} /* (17, 11, 15) {real, imag} */,
  {32'h40a0536e, 32'h40a1dbd5} /* (17, 11, 14) {real, imag} */,
  {32'h4064524d, 32'hbe672d30} /* (17, 11, 13) {real, imag} */,
  {32'hbf0d7aec, 32'h411ba321} /* (17, 11, 12) {real, imag} */,
  {32'hc101e31e, 32'hc08969be} /* (17, 11, 11) {real, imag} */,
  {32'hbeaa7ec0, 32'hc085cc78} /* (17, 11, 10) {real, imag} */,
  {32'h3e902f98, 32'h408553fa} /* (17, 11, 9) {real, imag} */,
  {32'hc02888a0, 32'hc07acdb7} /* (17, 11, 8) {real, imag} */,
  {32'hc1222c6a, 32'hc182008d} /* (17, 11, 7) {real, imag} */,
  {32'hc0fb3290, 32'hc103530b} /* (17, 11, 6) {real, imag} */,
  {32'h4185dc3d, 32'h41baa324} /* (17, 11, 5) {real, imag} */,
  {32'h414b1bc6, 32'hc1b5e98c} /* (17, 11, 4) {real, imag} */,
  {32'hc1126ba3, 32'h40c671a2} /* (17, 11, 3) {real, imag} */,
  {32'hbe62b460, 32'hc177df70} /* (17, 11, 2) {real, imag} */,
  {32'hc1a00e52, 32'h3f79a348} /* (17, 11, 1) {real, imag} */,
  {32'h4092ed8c, 32'hc135d1a9} /* (17, 11, 0) {real, imag} */,
  {32'h4022f880, 32'h4175c933} /* (17, 10, 31) {real, imag} */,
  {32'h4096c2c8, 32'hc1a4ce11} /* (17, 10, 30) {real, imag} */,
  {32'h40f81fa2, 32'hc02b91d5} /* (17, 10, 29) {real, imag} */,
  {32'h41923445, 32'hc14e75b8} /* (17, 10, 28) {real, imag} */,
  {32'h41b09f30, 32'h417184d6} /* (17, 10, 27) {real, imag} */,
  {32'h3f0f45e4, 32'hc02f8bf8} /* (17, 10, 26) {real, imag} */,
  {32'h41206578, 32'hc0d7b87c} /* (17, 10, 25) {real, imag} */,
  {32'hc1663139, 32'hc07fbf37} /* (17, 10, 24) {real, imag} */,
  {32'hc103e431, 32'hc16a3a20} /* (17, 10, 23) {real, imag} */,
  {32'h4092cf70, 32'h3fc77370} /* (17, 10, 22) {real, imag} */,
  {32'h40f31388, 32'h3f7c9ff8} /* (17, 10, 21) {real, imag} */,
  {32'hc1000867, 32'h3fcfa52e} /* (17, 10, 20) {real, imag} */,
  {32'hc1036764, 32'hc0025b69} /* (17, 10, 19) {real, imag} */,
  {32'h40fe25e6, 32'hc0782e62} /* (17, 10, 18) {real, imag} */,
  {32'h41013a03, 32'h40ae2570} /* (17, 10, 17) {real, imag} */,
  {32'h408801f4, 32'h3fbdcf38} /* (17, 10, 16) {real, imag} */,
  {32'hc0896c0a, 32'hbe307310} /* (17, 10, 15) {real, imag} */,
  {32'h4036726b, 32'h403d22ba} /* (17, 10, 14) {real, imag} */,
  {32'h4108c2a8, 32'h40182483} /* (17, 10, 13) {real, imag} */,
  {32'hc095839a, 32'hc1180c48} /* (17, 10, 12) {real, imag} */,
  {32'hc0e698b8, 32'h3f31dce8} /* (17, 10, 11) {real, imag} */,
  {32'h4114cc8a, 32'hc1618b02} /* (17, 10, 10) {real, imag} */,
  {32'hc037ea39, 32'hc12b4e60} /* (17, 10, 9) {real, imag} */,
  {32'hc04b815c, 32'h40e41d20} /* (17, 10, 8) {real, imag} */,
  {32'hc0d0354b, 32'h4187479f} /* (17, 10, 7) {real, imag} */,
  {32'h409acc64, 32'hc143f8b4} /* (17, 10, 6) {real, imag} */,
  {32'hc1299ea9, 32'hc1242fb2} /* (17, 10, 5) {real, imag} */,
  {32'h41284ee3, 32'h420221a2} /* (17, 10, 4) {real, imag} */,
  {32'h406115d3, 32'h40ac8b88} /* (17, 10, 3) {real, imag} */,
  {32'hc17260f8, 32'hc105bd2e} /* (17, 10, 2) {real, imag} */,
  {32'hc27968f2, 32'h41527e41} /* (17, 10, 1) {real, imag} */,
  {32'h40987fa0, 32'h4173f3d3} /* (17, 10, 0) {real, imag} */,
  {32'hbfac32c8, 32'hc10871dc} /* (17, 9, 31) {real, imag} */,
  {32'h4073b6c0, 32'hc183ff48} /* (17, 9, 30) {real, imag} */,
  {32'hc1b465e1, 32'h41f28b3f} /* (17, 9, 29) {real, imag} */,
  {32'hc1879364, 32'hc1097645} /* (17, 9, 28) {real, imag} */,
  {32'h404d3028, 32'hc11ea304} /* (17, 9, 27) {real, imag} */,
  {32'hc0f635de, 32'h40abb388} /* (17, 9, 26) {real, imag} */,
  {32'h41755be0, 32'h3fcfbf9c} /* (17, 9, 25) {real, imag} */,
  {32'h411cb89a, 32'h42169eee} /* (17, 9, 24) {real, imag} */,
  {32'h4179d2c2, 32'hc1758197} /* (17, 9, 23) {real, imag} */,
  {32'hc0d9c426, 32'h40eed0a6} /* (17, 9, 22) {real, imag} */,
  {32'h412c4bfc, 32'hbf075de8} /* (17, 9, 21) {real, imag} */,
  {32'hbf7f1d2c, 32'hc0dddfb2} /* (17, 9, 20) {real, imag} */,
  {32'hc0fd02e2, 32'h41440541} /* (17, 9, 19) {real, imag} */,
  {32'hc089d876, 32'hc0e69d87} /* (17, 9, 18) {real, imag} */,
  {32'hc0812345, 32'hbf576138} /* (17, 9, 17) {real, imag} */,
  {32'hc053dc1f, 32'h402d26d8} /* (17, 9, 16) {real, imag} */,
  {32'h3fa9327c, 32'h3ff1fda0} /* (17, 9, 15) {real, imag} */,
  {32'h3f592350, 32'h4056888e} /* (17, 9, 14) {real, imag} */,
  {32'hbeab4d08, 32'hc012598c} /* (17, 9, 13) {real, imag} */,
  {32'h401d29fb, 32'h40cbc08e} /* (17, 9, 12) {real, imag} */,
  {32'hbfccb9a8, 32'hc077618e} /* (17, 9, 11) {real, imag} */,
  {32'hc13f3801, 32'hc11aed43} /* (17, 9, 10) {real, imag} */,
  {32'h3f718da8, 32'h4106abed} /* (17, 9, 9) {real, imag} */,
  {32'h3fae4d7c, 32'h3f3eac00} /* (17, 9, 8) {real, imag} */,
  {32'hc0920ac0, 32'hc0e2fc5b} /* (17, 9, 7) {real, imag} */,
  {32'h40a3105e, 32'h40c422e0} /* (17, 9, 6) {real, imag} */,
  {32'h413b77cd, 32'hc139bd5a} /* (17, 9, 5) {real, imag} */,
  {32'hc1e7f52c, 32'h419429c8} /* (17, 9, 4) {real, imag} */,
  {32'hc17879c6, 32'hc1d3ee57} /* (17, 9, 3) {real, imag} */,
  {32'h41f53148, 32'hc10073dc} /* (17, 9, 2) {real, imag} */,
  {32'hc19a3d40, 32'hc04c7687} /* (17, 9, 1) {real, imag} */,
  {32'hbf8875ce, 32'h420f0304} /* (17, 9, 0) {real, imag} */,
  {32'hc1078620, 32'hc1334ce1} /* (17, 8, 31) {real, imag} */,
  {32'hc10d9384, 32'h41d5f112} /* (17, 8, 30) {real, imag} */,
  {32'h402d1c58, 32'hc09f419d} /* (17, 8, 29) {real, imag} */,
  {32'hc1899a9e, 32'h421e5f7c} /* (17, 8, 28) {real, imag} */,
  {32'hbf248970, 32'hc1d146fa} /* (17, 8, 27) {real, imag} */,
  {32'h40d935a0, 32'h402701ee} /* (17, 8, 26) {real, imag} */,
  {32'hc0a9fca2, 32'h3f1a5a20} /* (17, 8, 25) {real, imag} */,
  {32'h418ecf5c, 32'h3f7d4184} /* (17, 8, 24) {real, imag} */,
  {32'h400eb549, 32'h415a0574} /* (17, 8, 23) {real, imag} */,
  {32'hbf65d548, 32'hc1171dc8} /* (17, 8, 22) {real, imag} */,
  {32'h411b2871, 32'hc1621c5c} /* (17, 8, 21) {real, imag} */,
  {32'h40e1c37c, 32'hc0a85efe} /* (17, 8, 20) {real, imag} */,
  {32'h40e4330b, 32'h41072bd4} /* (17, 8, 19) {real, imag} */,
  {32'hc0d12f27, 32'h40fa1b6a} /* (17, 8, 18) {real, imag} */,
  {32'hbe581680, 32'hc13193a1} /* (17, 8, 17) {real, imag} */,
  {32'h407d44c7, 32'hc11169f8} /* (17, 8, 16) {real, imag} */,
  {32'h3fb2c0e0, 32'hbfebd1b8} /* (17, 8, 15) {real, imag} */,
  {32'h40034292, 32'h40874dba} /* (17, 8, 14) {real, imag} */,
  {32'hbf91dc64, 32'hc0614cb6} /* (17, 8, 13) {real, imag} */,
  {32'h40dfabd0, 32'hc06764cc} /* (17, 8, 12) {real, imag} */,
  {32'hc08f1ff2, 32'hc0946631} /* (17, 8, 11) {real, imag} */,
  {32'h3fd019dc, 32'hc093d4d7} /* (17, 8, 10) {real, imag} */,
  {32'hc0c9f612, 32'h4093c6a8} /* (17, 8, 9) {real, imag} */,
  {32'hc055714c, 32'h402f3feb} /* (17, 8, 8) {real, imag} */,
  {32'h4103c7b4, 32'hc1a32dc9} /* (17, 8, 7) {real, imag} */,
  {32'hbf737330, 32'h416bae22} /* (17, 8, 6) {real, imag} */,
  {32'hc1a1d312, 32'hc1b7bedc} /* (17, 8, 5) {real, imag} */,
  {32'h418bb8da, 32'h41544d22} /* (17, 8, 4) {real, imag} */,
  {32'h4192929f, 32'h414fa0b8} /* (17, 8, 3) {real, imag} */,
  {32'h3fac56ac, 32'hc187ffe2} /* (17, 8, 2) {real, imag} */,
  {32'hc1850367, 32'h41f11e8c} /* (17, 8, 1) {real, imag} */,
  {32'h3bb3e200, 32'h412eaef8} /* (17, 8, 0) {real, imag} */,
  {32'hc1e1c723, 32'h41bee3a0} /* (17, 7, 31) {real, imag} */,
  {32'h40b69bbf, 32'h41753024} /* (17, 7, 30) {real, imag} */,
  {32'h40f53f48, 32'h4190a26c} /* (17, 7, 29) {real, imag} */,
  {32'h41b7cec8, 32'h3de30b00} /* (17, 7, 28) {real, imag} */,
  {32'hc0ea8fb0, 32'hc05f65b6} /* (17, 7, 27) {real, imag} */,
  {32'hc1a57580, 32'h40c1ff2a} /* (17, 7, 26) {real, imag} */,
  {32'hc18214a3, 32'h408dfecc} /* (17, 7, 25) {real, imag} */,
  {32'hc0479a48, 32'hc13892d6} /* (17, 7, 24) {real, imag} */,
  {32'hc18db6e0, 32'h4067fc48} /* (17, 7, 23) {real, imag} */,
  {32'h400b9d94, 32'h40a20bbc} /* (17, 7, 22) {real, imag} */,
  {32'h409b2a42, 32'hc1a457de} /* (17, 7, 21) {real, imag} */,
  {32'hc02e1f80, 32'h411233ab} /* (17, 7, 20) {real, imag} */,
  {32'h400ac9a6, 32'h3e519970} /* (17, 7, 19) {real, imag} */,
  {32'hc14d4dad, 32'hc0ff02a8} /* (17, 7, 18) {real, imag} */,
  {32'hc04a6044, 32'h40489662} /* (17, 7, 17) {real, imag} */,
  {32'hc0e3a21c, 32'hc1465780} /* (17, 7, 16) {real, imag} */,
  {32'hc10d2f2b, 32'hc0e5e04b} /* (17, 7, 15) {real, imag} */,
  {32'hc0a63076, 32'hc0ce7888} /* (17, 7, 14) {real, imag} */,
  {32'h41523c0a, 32'h3d5631c0} /* (17, 7, 13) {real, imag} */,
  {32'hbfd15f70, 32'h4116c6e5} /* (17, 7, 12) {real, imag} */,
  {32'hc1428e99, 32'hc13663ab} /* (17, 7, 11) {real, imag} */,
  {32'hc193326c, 32'h3f448344} /* (17, 7, 10) {real, imag} */,
  {32'hc10b7634, 32'h41c79fec} /* (17, 7, 9) {real, imag} */,
  {32'h4144b1ce, 32'hc106ca84} /* (17, 7, 8) {real, imag} */,
  {32'h41d551a7, 32'h4188df50} /* (17, 7, 7) {real, imag} */,
  {32'hc1651e68, 32'hc0fa36be} /* (17, 7, 6) {real, imag} */,
  {32'h4080a650, 32'h410f0c24} /* (17, 7, 5) {real, imag} */,
  {32'hc0ec344e, 32'hc19de8a1} /* (17, 7, 4) {real, imag} */,
  {32'h41e808b2, 32'hc07a69ac} /* (17, 7, 3) {real, imag} */,
  {32'h40e010db, 32'hc1edf526} /* (17, 7, 2) {real, imag} */,
  {32'h40ee10c4, 32'h40ec5cb6} /* (17, 7, 1) {real, imag} */,
  {32'hc23a0930, 32'hc15abdb2} /* (17, 7, 0) {real, imag} */,
  {32'hc2854e12, 32'hbfa1e680} /* (17, 6, 31) {real, imag} */,
  {32'h40a3ae76, 32'hc1968494} /* (17, 6, 30) {real, imag} */,
  {32'h41d485b6, 32'hc0ce5636} /* (17, 6, 29) {real, imag} */,
  {32'h415f84ea, 32'h40852c1e} /* (17, 6, 28) {real, imag} */,
  {32'h4195a11c, 32'h4113f509} /* (17, 6, 27) {real, imag} */,
  {32'hc18141ac, 32'h400dec0f} /* (17, 6, 26) {real, imag} */,
  {32'h40befbe3, 32'hc0e8cdb2} /* (17, 6, 25) {real, imag} */,
  {32'h4170d766, 32'h41e4b09e} /* (17, 6, 24) {real, imag} */,
  {32'h404f8738, 32'hc130d69d} /* (17, 6, 23) {real, imag} */,
  {32'hc15de21e, 32'h416440a0} /* (17, 6, 22) {real, imag} */,
  {32'hbd94b3a0, 32'h3fdcb504} /* (17, 6, 21) {real, imag} */,
  {32'hc18f2fc4, 32'h418cab0a} /* (17, 6, 20) {real, imag} */,
  {32'hc16a410c, 32'h3f1ee0ba} /* (17, 6, 19) {real, imag} */,
  {32'hc0a1328b, 32'hbfa0f4c0} /* (17, 6, 18) {real, imag} */,
  {32'h40819af8, 32'h3fcc16b4} /* (17, 6, 17) {real, imag} */,
  {32'h40691ac8, 32'hc0978778} /* (17, 6, 16) {real, imag} */,
  {32'hbff0cc40, 32'h40af7fa6} /* (17, 6, 15) {real, imag} */,
  {32'hc13607b4, 32'hc13d863e} /* (17, 6, 14) {real, imag} */,
  {32'h3f95b870, 32'h3f9946d1} /* (17, 6, 13) {real, imag} */,
  {32'hc139e54f, 32'hc106a495} /* (17, 6, 12) {real, imag} */,
  {32'h4100d289, 32'h4185d481} /* (17, 6, 11) {real, imag} */,
  {32'hc079d3ae, 32'hbf5229a0} /* (17, 6, 10) {real, imag} */,
  {32'h41a652e7, 32'h40e33b7e} /* (17, 6, 9) {real, imag} */,
  {32'h3fbf8630, 32'h416ee094} /* (17, 6, 8) {real, imag} */,
  {32'hc16b5ec6, 32'h41c95296} /* (17, 6, 7) {real, imag} */,
  {32'h412497eb, 32'h407fe3d9} /* (17, 6, 6) {real, imag} */,
  {32'hc1007b5b, 32'hc03eba07} /* (17, 6, 5) {real, imag} */,
  {32'hc21857ac, 32'hc1095f3d} /* (17, 6, 4) {real, imag} */,
  {32'h41892842, 32'h406949ac} /* (17, 6, 3) {real, imag} */,
  {32'hc1e19e5c, 32'h4203c978} /* (17, 6, 2) {real, imag} */,
  {32'h3cbd4000, 32'hc138e58a} /* (17, 6, 1) {real, imag} */,
  {32'hc222fd44, 32'h420dc417} /* (17, 6, 0) {real, imag} */,
  {32'hbffb1910, 32'h40ddead0} /* (17, 5, 31) {real, imag} */,
  {32'h41ddf1c4, 32'hc1c47225} /* (17, 5, 30) {real, imag} */,
  {32'h41391925, 32'h41667326} /* (17, 5, 29) {real, imag} */,
  {32'h40d2a460, 32'hc1c9e232} /* (17, 5, 28) {real, imag} */,
  {32'hc1ca57cf, 32'hbfa89d50} /* (17, 5, 27) {real, imag} */,
  {32'h40263700, 32'h41dc0c69} /* (17, 5, 26) {real, imag} */,
  {32'hbff7b2f0, 32'hc1fad2c7} /* (17, 5, 25) {real, imag} */,
  {32'h41b84f0e, 32'hc154d808} /* (17, 5, 24) {real, imag} */,
  {32'h3e537c00, 32'h4020da42} /* (17, 5, 23) {real, imag} */,
  {32'h412ca3af, 32'hc19e6c52} /* (17, 5, 22) {real, imag} */,
  {32'hc0c9a21c, 32'hbffdc470} /* (17, 5, 21) {real, imag} */,
  {32'hc0e78cb2, 32'h4014ace5} /* (17, 5, 20) {real, imag} */,
  {32'h3fd03cfc, 32'h4049d5e6} /* (17, 5, 19) {real, imag} */,
  {32'h3f4d7eb0, 32'hbf82ffb4} /* (17, 5, 18) {real, imag} */,
  {32'h3facba24, 32'hc096c53e} /* (17, 5, 17) {real, imag} */,
  {32'h412c7eb0, 32'hc0b996b4} /* (17, 5, 16) {real, imag} */,
  {32'h412b979c, 32'hc0a2539e} /* (17, 5, 15) {real, imag} */,
  {32'h411cffe9, 32'hc0b521ed} /* (17, 5, 14) {real, imag} */,
  {32'hc0649a02, 32'h3f51b118} /* (17, 5, 13) {real, imag} */,
  {32'hc02033ec, 32'hc0886550} /* (17, 5, 12) {real, imag} */,
  {32'hc1b6f817, 32'h41caa9cd} /* (17, 5, 11) {real, imag} */,
  {32'h40d711f2, 32'h4173ccc3} /* (17, 5, 10) {real, imag} */,
  {32'h41158b94, 32'hbf0b96b8} /* (17, 5, 9) {real, imag} */,
  {32'hc11dcb44, 32'hc174889c} /* (17, 5, 8) {real, imag} */,
  {32'hc15c527a, 32'h418752b3} /* (17, 5, 7) {real, imag} */,
  {32'hc213c94e, 32'hc213cce2} /* (17, 5, 6) {real, imag} */,
  {32'h418c908d, 32'hc1ebe905} /* (17, 5, 5) {real, imag} */,
  {32'hc19270e0, 32'h413ac30b} /* (17, 5, 4) {real, imag} */,
  {32'h414fa263, 32'hc2235ba2} /* (17, 5, 3) {real, imag} */,
  {32'h424ff69e, 32'h424ef002} /* (17, 5, 2) {real, imag} */,
  {32'hc1feb2c3, 32'hc2705746} /* (17, 5, 1) {real, imag} */,
  {32'h4197e192, 32'hc1afe501} /* (17, 5, 0) {real, imag} */,
  {32'h403cb7a4, 32'h40452c0c} /* (17, 4, 31) {real, imag} */,
  {32'hc1e0f423, 32'hc20337fc} /* (17, 4, 30) {real, imag} */,
  {32'h4256ff43, 32'hc188c24a} /* (17, 4, 29) {real, imag} */,
  {32'h40ac2d4a, 32'h4231ae41} /* (17, 4, 28) {real, imag} */,
  {32'h413f8428, 32'h41bc684e} /* (17, 4, 27) {real, imag} */,
  {32'h4164dbcb, 32'hc175be52} /* (17, 4, 26) {real, imag} */,
  {32'h41249d4d, 32'h42044bc6} /* (17, 4, 25) {real, imag} */,
  {32'h40be8b6e, 32'hc19d54d0} /* (17, 4, 24) {real, imag} */,
  {32'h415491c0, 32'h3f614138} /* (17, 4, 23) {real, imag} */,
  {32'hc1832c77, 32'h4101f693} /* (17, 4, 22) {real, imag} */,
  {32'hc0532b2c, 32'h3f22a910} /* (17, 4, 21) {real, imag} */,
  {32'hc0c63cd6, 32'hc17aeb99} /* (17, 4, 20) {real, imag} */,
  {32'hbfc00978, 32'hc029d6dc} /* (17, 4, 19) {real, imag} */,
  {32'h41192f09, 32'hbe3a04e0} /* (17, 4, 18) {real, imag} */,
  {32'h406994c8, 32'hc09b8df2} /* (17, 4, 17) {real, imag} */,
  {32'hbf23ece0, 32'hbffe8ef8} /* (17, 4, 16) {real, imag} */,
  {32'hbf949460, 32'h410c3bcb} /* (17, 4, 15) {real, imag} */,
  {32'hc08d35d6, 32'hc0fa20cb} /* (17, 4, 14) {real, imag} */,
  {32'h413ca839, 32'hc1316825} /* (17, 4, 13) {real, imag} */,
  {32'h4139c187, 32'h3e6077c0} /* (17, 4, 12) {real, imag} */,
  {32'h40fa124a, 32'h4152ab4b} /* (17, 4, 11) {real, imag} */,
  {32'h4102c308, 32'hbfd638d8} /* (17, 4, 10) {real, imag} */,
  {32'h400f52f0, 32'h415e0e10} /* (17, 4, 9) {real, imag} */,
  {32'hc0dca96e, 32'hc1832228} /* (17, 4, 8) {real, imag} */,
  {32'hc0b92fe6, 32'h421f4296} /* (17, 4, 7) {real, imag} */,
  {32'h410deec1, 32'hc16a2ba6} /* (17, 4, 6) {real, imag} */,
  {32'hc280ba21, 32'hc018ce0c} /* (17, 4, 5) {real, imag} */,
  {32'hbf0a2558, 32'hc236a5e9} /* (17, 4, 4) {real, imag} */,
  {32'hc2291603, 32'h41234cfd} /* (17, 4, 3) {real, imag} */,
  {32'h421f4e4a, 32'h41a26ce8} /* (17, 4, 2) {real, imag} */,
  {32'hc1ce6510, 32'hc16cc1e1} /* (17, 4, 1) {real, imag} */,
  {32'h41a92d35, 32'h415778cb} /* (17, 4, 0) {real, imag} */,
  {32'h416ba6ee, 32'hc0c80124} /* (17, 3, 31) {real, imag} */,
  {32'hc1a9840e, 32'hc20466ff} /* (17, 3, 30) {real, imag} */,
  {32'hc1321609, 32'hc2190269} /* (17, 3, 29) {real, imag} */,
  {32'hc186645f, 32'hc1e66ccf} /* (17, 3, 28) {real, imag} */,
  {32'hc1087c4b, 32'h41576652} /* (17, 3, 27) {real, imag} */,
  {32'h41539410, 32'h3fb26e60} /* (17, 3, 26) {real, imag} */,
  {32'hc13c56e0, 32'hc16cb6a7} /* (17, 3, 25) {real, imag} */,
  {32'h411911a0, 32'h40ca91a1} /* (17, 3, 24) {real, imag} */,
  {32'hc1c825e6, 32'hc16fa6bf} /* (17, 3, 23) {real, imag} */,
  {32'hc1b5d915, 32'h40b4b1c0} /* (17, 3, 22) {real, imag} */,
  {32'h4182382c, 32'h41924dbc} /* (17, 3, 21) {real, imag} */,
  {32'hc094d9b5, 32'h416ea776} /* (17, 3, 20) {real, imag} */,
  {32'h40e3e772, 32'hbebb8840} /* (17, 3, 19) {real, imag} */,
  {32'hc13316f4, 32'h411843d6} /* (17, 3, 18) {real, imag} */,
  {32'h40eb3a0d, 32'h4017203c} /* (17, 3, 17) {real, imag} */,
  {32'h41315400, 32'hc03162ba} /* (17, 3, 16) {real, imag} */,
  {32'hbf21a3e8, 32'hc0ce5206} /* (17, 3, 15) {real, imag} */,
  {32'hc14ef9a8, 32'h40cf2973} /* (17, 3, 14) {real, imag} */,
  {32'h4135d999, 32'hc00908b8} /* (17, 3, 13) {real, imag} */,
  {32'hbfdb131d, 32'hc19cb7fb} /* (17, 3, 12) {real, imag} */,
  {32'h41851560, 32'hc0c9d959} /* (17, 3, 11) {real, imag} */,
  {32'hc17018e6, 32'h41ca5351} /* (17, 3, 10) {real, imag} */,
  {32'hc172442c, 32'hc1325543} /* (17, 3, 9) {real, imag} */,
  {32'h4218ca32, 32'hc13cb4be} /* (17, 3, 8) {real, imag} */,
  {32'hc182c380, 32'h41d315e6} /* (17, 3, 7) {real, imag} */,
  {32'hc16ec588, 32'h41ef1c6d} /* (17, 3, 6) {real, imag} */,
  {32'h41f451b2, 32'hc0d32723} /* (17, 3, 5) {real, imag} */,
  {32'hc1c1d459, 32'hbf928150} /* (17, 3, 4) {real, imag} */,
  {32'hc0058df4, 32'h41f8965e} /* (17, 3, 3) {real, imag} */,
  {32'hc06a3500, 32'hc1ddcb62} /* (17, 3, 2) {real, imag} */,
  {32'h414fb73a, 32'h4213574a} /* (17, 3, 1) {real, imag} */,
  {32'h4248183a, 32'h418831d5} /* (17, 3, 0) {real, imag} */,
  {32'h3f559cd0, 32'hc23c3a38} /* (17, 2, 31) {real, imag} */,
  {32'h419d2250, 32'hbf65d740} /* (17, 2, 30) {real, imag} */,
  {32'h4200e592, 32'h41eda484} /* (17, 2, 29) {real, imag} */,
  {32'hc14732ad, 32'h4161772e} /* (17, 2, 28) {real, imag} */,
  {32'hc1ec83e9, 32'hc056b57f} /* (17, 2, 27) {real, imag} */,
  {32'hc07acf4a, 32'h417a7416} /* (17, 2, 26) {real, imag} */,
  {32'hc1633cdc, 32'hbfd9b9e0} /* (17, 2, 25) {real, imag} */,
  {32'h41e327dc, 32'h414f6ba2} /* (17, 2, 24) {real, imag} */,
  {32'h3ee10530, 32'h421fa7d4} /* (17, 2, 23) {real, imag} */,
  {32'hc0301a08, 32'h41af8946} /* (17, 2, 22) {real, imag} */,
  {32'hc1e71907, 32'hc082fab0} /* (17, 2, 21) {real, imag} */,
  {32'h40ce90b4, 32'hbf2997d8} /* (17, 2, 20) {real, imag} */,
  {32'h3f189a80, 32'hc0ba36e4} /* (17, 2, 19) {real, imag} */,
  {32'h3e8bf0a0, 32'h40b230ec} /* (17, 2, 18) {real, imag} */,
  {32'hc0ae4576, 32'hc13b528e} /* (17, 2, 17) {real, imag} */,
  {32'h41169d51, 32'h40ca0776} /* (17, 2, 16) {real, imag} */,
  {32'h40e8905e, 32'h40cfbefc} /* (17, 2, 15) {real, imag} */,
  {32'hc13a3ac5, 32'hc11b7860} /* (17, 2, 14) {real, imag} */,
  {32'hc086e540, 32'h3fe59e40} /* (17, 2, 13) {real, imag} */,
  {32'h40cce708, 32'hc0cc4859} /* (17, 2, 12) {real, imag} */,
  {32'h410b82ae, 32'h411dc089} /* (17, 2, 11) {real, imag} */,
  {32'h41857789, 32'hc0eb7dae} /* (17, 2, 10) {real, imag} */,
  {32'hc11493da, 32'hc19c270c} /* (17, 2, 9) {real, imag} */,
  {32'h41aa52d0, 32'h40750cee} /* (17, 2, 8) {real, imag} */,
  {32'hc1bdb84c, 32'hc1509ca4} /* (17, 2, 7) {real, imag} */,
  {32'h412a1b96, 32'h4174e124} /* (17, 2, 6) {real, imag} */,
  {32'hc1f8f4cf, 32'h41353f1b} /* (17, 2, 5) {real, imag} */,
  {32'h41302ef5, 32'h41e52825} /* (17, 2, 4) {real, imag} */,
  {32'hc1a53470, 32'h418c4450} /* (17, 2, 3) {real, imag} */,
  {32'h428e8fb8, 32'h42230bb9} /* (17, 2, 2) {real, imag} */,
  {32'h3fe88018, 32'hc1ebf940} /* (17, 2, 1) {real, imag} */,
  {32'hc0fcb8d6, 32'hc1e986b6} /* (17, 2, 0) {real, imag} */,
  {32'h42723857, 32'hc235f722} /* (17, 1, 31) {real, imag} */,
  {32'hc134d626, 32'h426c5508} /* (17, 1, 30) {real, imag} */,
  {32'h3ed111c0, 32'hc1ab04a8} /* (17, 1, 29) {real, imag} */,
  {32'h3f8a1bc8, 32'hc1f33fc7} /* (17, 1, 28) {real, imag} */,
  {32'h41caeadc, 32'h421baf10} /* (17, 1, 27) {real, imag} */,
  {32'hc125a578, 32'hc23f0837} /* (17, 1, 26) {real, imag} */,
  {32'h4230dab0, 32'hc2102416} /* (17, 1, 25) {real, imag} */,
  {32'hc0462312, 32'h42107454} /* (17, 1, 24) {real, imag} */,
  {32'h416d570c, 32'h41f85790} /* (17, 1, 23) {real, imag} */,
  {32'h3fc709c4, 32'hc01cabdc} /* (17, 1, 22) {real, imag} */,
  {32'h416d634e, 32'h40837b04} /* (17, 1, 21) {real, imag} */,
  {32'h41f9f917, 32'hbfd3f31c} /* (17, 1, 20) {real, imag} */,
  {32'h4003b896, 32'hbfb63f30} /* (17, 1, 19) {real, imag} */,
  {32'hc0a2c9b2, 32'h3fb6d6f8} /* (17, 1, 18) {real, imag} */,
  {32'h4150377a, 32'hc15a14d5} /* (17, 1, 17) {real, imag} */,
  {32'h3e5a77c0, 32'hbe7cd400} /* (17, 1, 16) {real, imag} */,
  {32'hc0be9474, 32'hc113db3d} /* (17, 1, 15) {real, imag} */,
  {32'hc10803d5, 32'h40b9f01e} /* (17, 1, 14) {real, imag} */,
  {32'hc060ea3a, 32'hc141808e} /* (17, 1, 13) {real, imag} */,
  {32'h41054962, 32'h410c711e} /* (17, 1, 12) {real, imag} */,
  {32'hc00d4a5a, 32'h418002e3} /* (17, 1, 11) {real, imag} */,
  {32'h4153ec4e, 32'hc1b8bcac} /* (17, 1, 10) {real, imag} */,
  {32'hc13c6114, 32'hc1b9bbf8} /* (17, 1, 9) {real, imag} */,
  {32'hc1896dab, 32'h40a59ec6} /* (17, 1, 8) {real, imag} */,
  {32'h418d3c54, 32'h413afc9a} /* (17, 1, 7) {real, imag} */,
  {32'hc06d6eba, 32'hc2028b75} /* (17, 1, 6) {real, imag} */,
  {32'hc2815ef1, 32'hc215a27c} /* (17, 1, 5) {real, imag} */,
  {32'h418f4fb6, 32'hc1b7cdcd} /* (17, 1, 4) {real, imag} */,
  {32'hc1ef08c3, 32'hc2c19a1c} /* (17, 1, 3) {real, imag} */,
  {32'hc25115ea, 32'hc1c182a8} /* (17, 1, 2) {real, imag} */,
  {32'h41f15082, 32'h41d1e678} /* (17, 1, 1) {real, imag} */,
  {32'h3f65c290, 32'h41bf2a16} /* (17, 1, 0) {real, imag} */,
  {32'hc1d23cd4, 32'h412b8af4} /* (17, 0, 31) {real, imag} */,
  {32'h3e9a2c00, 32'h3c936800} /* (17, 0, 30) {real, imag} */,
  {32'hc21e20df, 32'h424bc56e} /* (17, 0, 29) {real, imag} */,
  {32'hc2273da2, 32'h4107c44e} /* (17, 0, 28) {real, imag} */,
  {32'hc090f723, 32'h40a5d2ca} /* (17, 0, 27) {real, imag} */,
  {32'h41852530, 32'hc117dfcb} /* (17, 0, 26) {real, imag} */,
  {32'h41650b4a, 32'h422e64d8} /* (17, 0, 25) {real, imag} */,
  {32'h4254212b, 32'h41973f89} /* (17, 0, 24) {real, imag} */,
  {32'h3f7d4180, 32'hc2008206} /* (17, 0, 23) {real, imag} */,
  {32'hc101c80b, 32'hc12a8751} /* (17, 0, 22) {real, imag} */,
  {32'hc12dae1e, 32'hc198d722} /* (17, 0, 21) {real, imag} */,
  {32'h40edd4c3, 32'hc0067698} /* (17, 0, 20) {real, imag} */,
  {32'h418cf347, 32'hc0ad30b2} /* (17, 0, 19) {real, imag} */,
  {32'hc12f1a24, 32'h40bf3fa6} /* (17, 0, 18) {real, imag} */,
  {32'hbebd18a0, 32'h40f2efce} /* (17, 0, 17) {real, imag} */,
  {32'h4097d490, 32'hc02b0c28} /* (17, 0, 16) {real, imag} */,
  {32'h4085df1e, 32'hc101f5a7} /* (17, 0, 15) {real, imag} */,
  {32'h41c193ea, 32'h407769d4} /* (17, 0, 14) {real, imag} */,
  {32'hc14b7212, 32'hc18bf8c4} /* (17, 0, 13) {real, imag} */,
  {32'h402945ca, 32'h40e5f484} /* (17, 0, 12) {real, imag} */,
  {32'hc0fa804b, 32'hc09a8436} /* (17, 0, 11) {real, imag} */,
  {32'h41699969, 32'h411d0ad1} /* (17, 0, 10) {real, imag} */,
  {32'h413c58a6, 32'hc133ab36} /* (17, 0, 9) {real, imag} */,
  {32'hc1b4afaa, 32'h3e1e6180} /* (17, 0, 8) {real, imag} */,
  {32'h413672b8, 32'hc0363898} /* (17, 0, 7) {real, imag} */,
  {32'hc12dd133, 32'h41ae0c5a} /* (17, 0, 6) {real, imag} */,
  {32'hc181ce13, 32'hc1ac20b8} /* (17, 0, 5) {real, imag} */,
  {32'hc22e96a2, 32'h41c61ce7} /* (17, 0, 4) {real, imag} */,
  {32'hc11b3b94, 32'h4242c5fa} /* (17, 0, 3) {real, imag} */,
  {32'h415278b8, 32'hc2043447} /* (17, 0, 2) {real, imag} */,
  {32'h402ba7ec, 32'h42784f4f} /* (17, 0, 1) {real, imag} */,
  {32'h419a3e68, 32'hc1d0595f} /* (17, 0, 0) {real, imag} */,
  {32'hc0c55bb2, 32'h3d71a200} /* (16, 31, 31) {real, imag} */,
  {32'hc1c34dae, 32'hc219aaa7} /* (16, 31, 30) {real, imag} */,
  {32'hc1434df5, 32'h4201f0d8} /* (16, 31, 29) {real, imag} */,
  {32'hc23ffe78, 32'h41a226b0} /* (16, 31, 28) {real, imag} */,
  {32'h4206b842, 32'h411b7764} /* (16, 31, 27) {real, imag} */,
  {32'h40c3f5c4, 32'hc11e1a46} /* (16, 31, 26) {real, imag} */,
  {32'hc0c9ab50, 32'h40fc6930} /* (16, 31, 25) {real, imag} */,
  {32'h3ff30c20, 32'h3fc4bb40} /* (16, 31, 24) {real, imag} */,
  {32'h418973c6, 32'h41b6c708} /* (16, 31, 23) {real, imag} */,
  {32'hc1c6d3ca, 32'hc0fb726a} /* (16, 31, 22) {real, imag} */,
  {32'hc0aa44d2, 32'h41b6e5ea} /* (16, 31, 21) {real, imag} */,
  {32'h40017dc8, 32'h41132bb4} /* (16, 31, 20) {real, imag} */,
  {32'h40827518, 32'hc16cd054} /* (16, 31, 19) {real, imag} */,
  {32'hbec1c350, 32'hc032d4f0} /* (16, 31, 18) {real, imag} */,
  {32'h3f12c010, 32'hbd5cb500} /* (16, 31, 17) {real, imag} */,
  {32'h3f841960, 32'hc1141b32} /* (16, 31, 16) {real, imag} */,
  {32'hbf350610, 32'h3e6169c0} /* (16, 31, 15) {real, imag} */,
  {32'h40920a31, 32'hc0862f80} /* (16, 31, 14) {real, imag} */,
  {32'h40e75994, 32'h4119f870} /* (16, 31, 13) {real, imag} */,
  {32'hc1b61bb7, 32'h3f8a9624} /* (16, 31, 12) {real, imag} */,
  {32'hc11323f1, 32'hc024b0a0} /* (16, 31, 11) {real, imag} */,
  {32'hc14bdbad, 32'hc1054671} /* (16, 31, 10) {real, imag} */,
  {32'hc12838bc, 32'h4076b798} /* (16, 31, 9) {real, imag} */,
  {32'hc068d040, 32'h41910d2a} /* (16, 31, 8) {real, imag} */,
  {32'hc034217c, 32'h3fe8b6ae} /* (16, 31, 7) {real, imag} */,
  {32'h4153e140, 32'hc1ae2aa6} /* (16, 31, 6) {real, imag} */,
  {32'hc04dc5c4, 32'h42075c54} /* (16, 31, 5) {real, imag} */,
  {32'h3fff6990, 32'h40059620} /* (16, 31, 4) {real, imag} */,
  {32'h41388991, 32'hc2251e74} /* (16, 31, 3) {real, imag} */,
  {32'hc18ff5f2, 32'hc22f777d} /* (16, 31, 2) {real, imag} */,
  {32'h41a20dee, 32'hc216608e} /* (16, 31, 1) {real, imag} */,
  {32'h41f65d90, 32'h4120a604} /* (16, 31, 0) {real, imag} */,
  {32'hc2389c54, 32'hc1882350} /* (16, 30, 31) {real, imag} */,
  {32'hc170449c, 32'hc1a0012e} /* (16, 30, 30) {real, imag} */,
  {32'hc194d7ef, 32'h41b97954} /* (16, 30, 29) {real, imag} */,
  {32'hc1452a54, 32'hc2128f21} /* (16, 30, 28) {real, imag} */,
  {32'h420a7dcd, 32'h40c3b62c} /* (16, 30, 27) {real, imag} */,
  {32'h4112b07d, 32'hc2003ec2} /* (16, 30, 26) {real, imag} */,
  {32'hc0e68ab9, 32'hbf9fe8e0} /* (16, 30, 25) {real, imag} */,
  {32'hc17075f9, 32'hc1916e24} /* (16, 30, 24) {real, imag} */,
  {32'hbf078470, 32'hc06614a4} /* (16, 30, 23) {real, imag} */,
  {32'h41c08963, 32'hc061e906} /* (16, 30, 22) {real, imag} */,
  {32'h41cb1142, 32'hc1280bc1} /* (16, 30, 21) {real, imag} */,
  {32'hbf1548b2, 32'h41224e64} /* (16, 30, 20) {real, imag} */,
  {32'hc108a1cd, 32'h3ffadaf0} /* (16, 30, 19) {real, imag} */,
  {32'hc0735166, 32'h406a4954} /* (16, 30, 18) {real, imag} */,
  {32'hc0f100b4, 32'h40a7b904} /* (16, 30, 17) {real, imag} */,
  {32'h3f049302, 32'h3fdd621c} /* (16, 30, 16) {real, imag} */,
  {32'hc00ceee8, 32'hc154e116} /* (16, 30, 15) {real, imag} */,
  {32'hbe8ea8b0, 32'h408e3536} /* (16, 30, 14) {real, imag} */,
  {32'hc1a66c34, 32'hc17c1ec4} /* (16, 30, 13) {real, imag} */,
  {32'hbfcee6d1, 32'hc04629ea} /* (16, 30, 12) {real, imag} */,
  {32'h40cdfff8, 32'hc02502cd} /* (16, 30, 11) {real, imag} */,
  {32'hc2138934, 32'hc11c454e} /* (16, 30, 10) {real, imag} */,
  {32'h41b1d8cc, 32'h4146d713} /* (16, 30, 9) {real, imag} */,
  {32'h4103f8ff, 32'hc1a45254} /* (16, 30, 8) {real, imag} */,
  {32'hbdae7e40, 32'h4191d5dc} /* (16, 30, 7) {real, imag} */,
  {32'h40d76aae, 32'hc12566fe} /* (16, 30, 6) {real, imag} */,
  {32'hc1b03a63, 32'h3d3a31c0} /* (16, 30, 5) {real, imag} */,
  {32'h41847134, 32'h4110643c} /* (16, 30, 4) {real, imag} */,
  {32'hc190ec47, 32'h419d296c} /* (16, 30, 3) {real, imag} */,
  {32'h41d43918, 32'hc11c49a7} /* (16, 30, 2) {real, imag} */,
  {32'h3f881170, 32'h4138adc7} /* (16, 30, 1) {real, imag} */,
  {32'h40058fda, 32'hc104b9ae} /* (16, 30, 0) {real, imag} */,
  {32'hc24ccecc, 32'hc2044ff5} /* (16, 29, 31) {real, imag} */,
  {32'h40d364d4, 32'h42265f0c} /* (16, 29, 30) {real, imag} */,
  {32'hc1ef874e, 32'hc0dd7030} /* (16, 29, 29) {real, imag} */,
  {32'hc097e75c, 32'h414d3aac} /* (16, 29, 28) {real, imag} */,
  {32'h41b90a87, 32'hc1499512} /* (16, 29, 27) {real, imag} */,
  {32'hc106b22f, 32'h41492f6b} /* (16, 29, 26) {real, imag} */,
  {32'h407f88c0, 32'hc20a868f} /* (16, 29, 25) {real, imag} */,
  {32'h41604a40, 32'h4060924c} /* (16, 29, 24) {real, imag} */,
  {32'hc1603ac0, 32'h4170e0a2} /* (16, 29, 23) {real, imag} */,
  {32'h417e4585, 32'h400a47fc} /* (16, 29, 22) {real, imag} */,
  {32'h41b56ca2, 32'hc1d3e23f} /* (16, 29, 21) {real, imag} */,
  {32'h3f7a2560, 32'h40f08c9f} /* (16, 29, 20) {real, imag} */,
  {32'hc08d6c87, 32'h41aac82e} /* (16, 29, 19) {real, imag} */,
  {32'h40a834d6, 32'h4141f2f8} /* (16, 29, 18) {real, imag} */,
  {32'hc0b69a08, 32'hc0f3b438} /* (16, 29, 17) {real, imag} */,
  {32'hbf4ca5f0, 32'hc061df8c} /* (16, 29, 16) {real, imag} */,
  {32'h41321a50, 32'h40d08b10} /* (16, 29, 15) {real, imag} */,
  {32'hc154be4f, 32'h3fcaae34} /* (16, 29, 14) {real, imag} */,
  {32'h40d30bc7, 32'h4063ea00} /* (16, 29, 13) {real, imag} */,
  {32'hc0da5114, 32'hc0d1bc6d} /* (16, 29, 12) {real, imag} */,
  {32'hc154c910, 32'hc0a1e81c} /* (16, 29, 11) {real, imag} */,
  {32'h412ecc73, 32'hbf118b72} /* (16, 29, 10) {real, imag} */,
  {32'hc0746b82, 32'h4119f790} /* (16, 29, 9) {real, imag} */,
  {32'hc106fcc8, 32'h41b72940} /* (16, 29, 8) {real, imag} */,
  {32'hc1d9fba0, 32'h416df2eb} /* (16, 29, 7) {real, imag} */,
  {32'h419bf740, 32'h41619d55} /* (16, 29, 6) {real, imag} */,
  {32'hc0cff16c, 32'h41b558e7} /* (16, 29, 5) {real, imag} */,
  {32'h42176de8, 32'hc15cc37a} /* (16, 29, 4) {real, imag} */,
  {32'hc21d7df9, 32'hc250da55} /* (16, 29, 3) {real, imag} */,
  {32'hc1589dbc, 32'h41892a23} /* (16, 29, 2) {real, imag} */,
  {32'hc2581394, 32'hc202e067} /* (16, 29, 1) {real, imag} */,
  {32'hc1196ac5, 32'h3fa939d0} /* (16, 29, 0) {real, imag} */,
  {32'h3e4d8540, 32'h4194e2dc} /* (16, 28, 31) {real, imag} */,
  {32'hc0cf7d14, 32'hc25388a0} /* (16, 28, 30) {real, imag} */,
  {32'h41d33394, 32'h40c76559} /* (16, 28, 29) {real, imag} */,
  {32'h418e8ffa, 32'h424ce00a} /* (16, 28, 28) {real, imag} */,
  {32'h413af707, 32'hc1bf0c20} /* (16, 28, 27) {real, imag} */,
  {32'hc1e59722, 32'hc161c07a} /* (16, 28, 26) {real, imag} */,
  {32'hc1aa64c6, 32'hc1408190} /* (16, 28, 25) {real, imag} */,
  {32'h41319e46, 32'h41658468} /* (16, 28, 24) {real, imag} */,
  {32'h41349c22, 32'hc18a3fb6} /* (16, 28, 23) {real, imag} */,
  {32'h41494f1b, 32'hc2079f4a} /* (16, 28, 22) {real, imag} */,
  {32'hc145e5ea, 32'h4189f10a} /* (16, 28, 21) {real, imag} */,
  {32'h4110d217, 32'h40faf578} /* (16, 28, 20) {real, imag} */,
  {32'hc0b6acbd, 32'hc1159970} /* (16, 28, 19) {real, imag} */,
  {32'h41099216, 32'h403a0bba} /* (16, 28, 18) {real, imag} */,
  {32'hc116cc1f, 32'h40c0d12e} /* (16, 28, 17) {real, imag} */,
  {32'hbf46eb00, 32'h40f81ffa} /* (16, 28, 16) {real, imag} */,
  {32'hc180dc7e, 32'hc188629e} /* (16, 28, 15) {real, imag} */,
  {32'hc132477e, 32'h4007a876} /* (16, 28, 14) {real, imag} */,
  {32'hc025f902, 32'h40a44511} /* (16, 28, 13) {real, imag} */,
  {32'h4040833c, 32'h418012ae} /* (16, 28, 12) {real, imag} */,
  {32'h40b7bed4, 32'hc0cee74a} /* (16, 28, 11) {real, imag} */,
  {32'h408eb392, 32'hc11861b6} /* (16, 28, 10) {real, imag} */,
  {32'h41d9fa1b, 32'h4024c830} /* (16, 28, 9) {real, imag} */,
  {32'hc187d90e, 32'hc087bc2f} /* (16, 28, 8) {real, imag} */,
  {32'h41c98960, 32'h41915324} /* (16, 28, 7) {real, imag} */,
  {32'h41c26742, 32'h3fe0bb48} /* (16, 28, 6) {real, imag} */,
  {32'hc116e611, 32'hc20974e4} /* (16, 28, 5) {real, imag} */,
  {32'hc233be43, 32'hc0cf39f0} /* (16, 28, 4) {real, imag} */,
  {32'hbf8143f8, 32'hc0f0a443} /* (16, 28, 3) {real, imag} */,
  {32'hc1968cb9, 32'hc202c5cc} /* (16, 28, 2) {real, imag} */,
  {32'h41be198c, 32'h426c7076} /* (16, 28, 1) {real, imag} */,
  {32'hc1b19894, 32'h418eb0be} /* (16, 28, 0) {real, imag} */,
  {32'hc15f6fec, 32'h4184061a} /* (16, 27, 31) {real, imag} */,
  {32'hc1f11b9c, 32'hc0de47f8} /* (16, 27, 30) {real, imag} */,
  {32'h419d18d9, 32'hc2047708} /* (16, 27, 29) {real, imag} */,
  {32'hc0be0072, 32'h41fb08d0} /* (16, 27, 28) {real, imag} */,
  {32'hc08128ae, 32'hc221a0d1} /* (16, 27, 27) {real, imag} */,
  {32'hc012e0f4, 32'hc1334fe6} /* (16, 27, 26) {real, imag} */,
  {32'hc0e31610, 32'hc112925c} /* (16, 27, 25) {real, imag} */,
  {32'h41aa9c18, 32'h40d6eab8} /* (16, 27, 24) {real, imag} */,
  {32'hc11c47b4, 32'hc13bded9} /* (16, 27, 23) {real, imag} */,
  {32'h409118d2, 32'hbe555ee0} /* (16, 27, 22) {real, imag} */,
  {32'h41797219, 32'hc0ae4458} /* (16, 27, 21) {real, imag} */,
  {32'hc0b779ee, 32'h405e23da} /* (16, 27, 20) {real, imag} */,
  {32'hbf6de518, 32'hc032a2d8} /* (16, 27, 19) {real, imag} */,
  {32'h409605ca, 32'hc07eaf4c} /* (16, 27, 18) {real, imag} */,
  {32'h400d35d6, 32'hc131c8ce} /* (16, 27, 17) {real, imag} */,
  {32'h3ed29620, 32'h40729ac4} /* (16, 27, 16) {real, imag} */,
  {32'hc095f913, 32'hbf0c08c8} /* (16, 27, 15) {real, imag} */,
  {32'hc0feb4ca, 32'h3fb93d18} /* (16, 27, 14) {real, imag} */,
  {32'h3ff4663c, 32'h41578600} /* (16, 27, 13) {real, imag} */,
  {32'hc1684f8d, 32'h3fde4814} /* (16, 27, 12) {real, imag} */,
  {32'h40a6d4a6, 32'h41515756} /* (16, 27, 11) {real, imag} */,
  {32'h40bac756, 32'hbefa1010} /* (16, 27, 10) {real, imag} */,
  {32'h3eed7440, 32'h41031fab} /* (16, 27, 9) {real, imag} */,
  {32'h4150d697, 32'hc07f8b50} /* (16, 27, 8) {real, imag} */,
  {32'hbebcbec8, 32'hbff865d4} /* (16, 27, 7) {real, imag} */,
  {32'hc1462dd1, 32'hc185ac53} /* (16, 27, 6) {real, imag} */,
  {32'hc138e10d, 32'hc19dfee2} /* (16, 27, 5) {real, imag} */,
  {32'h411f1ded, 32'hc19a05dc} /* (16, 27, 4) {real, imag} */,
  {32'h4200105e, 32'h3e7f3a00} /* (16, 27, 3) {real, imag} */,
  {32'hc0d39eb2, 32'hc239d613} /* (16, 27, 2) {real, imag} */,
  {32'hc0eeb7e8, 32'h418ef3be} /* (16, 27, 1) {real, imag} */,
  {32'hc0bbf20e, 32'h4200cc8b} /* (16, 27, 0) {real, imag} */,
  {32'hc1f5e7f4, 32'h42391a02} /* (16, 26, 31) {real, imag} */,
  {32'hc15814ff, 32'h414fdb9c} /* (16, 26, 30) {real, imag} */,
  {32'hc0208aaa, 32'hc1c0cc97} /* (16, 26, 29) {real, imag} */,
  {32'h419989e8, 32'hbf537240} /* (16, 26, 28) {real, imag} */,
  {32'h41ef02f9, 32'hc106009a} /* (16, 26, 27) {real, imag} */,
  {32'h40d94506, 32'h414346f6} /* (16, 26, 26) {real, imag} */,
  {32'hc12bb1f6, 32'hc18df19c} /* (16, 26, 25) {real, imag} */,
  {32'h41cd0336, 32'h3fe20658} /* (16, 26, 24) {real, imag} */,
  {32'h4093323c, 32'h414f79c2} /* (16, 26, 23) {real, imag} */,
  {32'hc156c5bd, 32'hbf51ab10} /* (16, 26, 22) {real, imag} */,
  {32'h41440a4d, 32'h41a306eb} /* (16, 26, 21) {real, imag} */,
  {32'h40b60816, 32'h3f94ced8} /* (16, 26, 20) {real, imag} */,
  {32'hbe763660, 32'h4027c72e} /* (16, 26, 19) {real, imag} */,
  {32'h402276aa, 32'hbffbe23a} /* (16, 26, 18) {real, imag} */,
  {32'h40d85626, 32'hc09285f5} /* (16, 26, 17) {real, imag} */,
  {32'hbefef700, 32'h3d2a9400} /* (16, 26, 16) {real, imag} */,
  {32'hc04571e4, 32'h411146f4} /* (16, 26, 15) {real, imag} */,
  {32'hc061f836, 32'h40dade9e} /* (16, 26, 14) {real, imag} */,
  {32'h410f307c, 32'h410f5b50} /* (16, 26, 13) {real, imag} */,
  {32'h414ffdf5, 32'hc0d731ee} /* (16, 26, 12) {real, imag} */,
  {32'h40dce1d6, 32'h40ae823f} /* (16, 26, 11) {real, imag} */,
  {32'h4081a052, 32'h41719a29} /* (16, 26, 10) {real, imag} */,
  {32'hc1290c3b, 32'h3fd8d0b4} /* (16, 26, 9) {real, imag} */,
  {32'h413d5044, 32'hc028a91c} /* (16, 26, 8) {real, imag} */,
  {32'hc1910515, 32'h41956568} /* (16, 26, 7) {real, imag} */,
  {32'hc1890a94, 32'h3f2064a0} /* (16, 26, 6) {real, imag} */,
  {32'hc1a2792b, 32'hc1bc6196} /* (16, 26, 5) {real, imag} */,
  {32'hc1e9e7ac, 32'hbf48ba7c} /* (16, 26, 4) {real, imag} */,
  {32'hc155fa1c, 32'hc2070b2e} /* (16, 26, 3) {real, imag} */,
  {32'h4149b8a9, 32'hc1b74eaa} /* (16, 26, 2) {real, imag} */,
  {32'hc19a43f8, 32'h4130680a} /* (16, 26, 1) {real, imag} */,
  {32'h402655c0, 32'h41f219f6} /* (16, 26, 0) {real, imag} */,
  {32'h4190e8de, 32'h3ed15e80} /* (16, 25, 31) {real, imag} */,
  {32'hc1874915, 32'hbfc7af28} /* (16, 25, 30) {real, imag} */,
  {32'hc07b29f8, 32'hc1e2bf52} /* (16, 25, 29) {real, imag} */,
  {32'hc1d51300, 32'hc193f527} /* (16, 25, 28) {real, imag} */,
  {32'hc137aaaa, 32'hc20a4b89} /* (16, 25, 27) {real, imag} */,
  {32'h3fafbbd4, 32'hc0d28115} /* (16, 25, 26) {real, imag} */,
  {32'hc1cab4ab, 32'h40007078} /* (16, 25, 25) {real, imag} */,
  {32'h408294bc, 32'h40e39cde} /* (16, 25, 24) {real, imag} */,
  {32'hbfe9a2ec, 32'h41a1a7a8} /* (16, 25, 23) {real, imag} */,
  {32'hc0719784, 32'h409a4ee6} /* (16, 25, 22) {real, imag} */,
  {32'h402f9840, 32'hbd5a5400} /* (16, 25, 21) {real, imag} */,
  {32'hbf37f7b8, 32'hc123d956} /* (16, 25, 20) {real, imag} */,
  {32'hc0c5f088, 32'hc0905af8} /* (16, 25, 19) {real, imag} */,
  {32'h4086a61f, 32'hc0a90c56} /* (16, 25, 18) {real, imag} */,
  {32'h3f6dbc74, 32'h403dc972} /* (16, 25, 17) {real, imag} */,
  {32'hc083d98f, 32'hc0a7be04} /* (16, 25, 16) {real, imag} */,
  {32'hc00b5057, 32'h40930d6d} /* (16, 25, 15) {real, imag} */,
  {32'h3eb4af50, 32'hbf8c9f6e} /* (16, 25, 14) {real, imag} */,
  {32'hc028b348, 32'h405b1798} /* (16, 25, 13) {real, imag} */,
  {32'hc0ca9e7d, 32'h40aa97b4} /* (16, 25, 12) {real, imag} */,
  {32'h4110ea84, 32'h3f6fcc80} /* (16, 25, 11) {real, imag} */,
  {32'hc19516f6, 32'h4147163d} /* (16, 25, 10) {real, imag} */,
  {32'h40b41e13, 32'h3e9e9760} /* (16, 25, 9) {real, imag} */,
  {32'hc0c8415a, 32'hbf082bf0} /* (16, 25, 8) {real, imag} */,
  {32'hc18e67a7, 32'hc133e7ab} /* (16, 25, 7) {real, imag} */,
  {32'h41479c88, 32'h41047630} /* (16, 25, 6) {real, imag} */,
  {32'h40d79c54, 32'hc11132f8} /* (16, 25, 5) {real, imag} */,
  {32'hc12f6230, 32'h4033c5a8} /* (16, 25, 4) {real, imag} */,
  {32'hc12d8080, 32'hc141f233} /* (16, 25, 3) {real, imag} */,
  {32'hbf6a06f8, 32'hc16c927b} /* (16, 25, 2) {real, imag} */,
  {32'hc0de19fe, 32'h418b55d4} /* (16, 25, 1) {real, imag} */,
  {32'h40aeb359, 32'hc1e530a9} /* (16, 25, 0) {real, imag} */,
  {32'hc17db0e0, 32'hc1f4048c} /* (16, 24, 31) {real, imag} */,
  {32'hc11d2129, 32'hc1b55160} /* (16, 24, 30) {real, imag} */,
  {32'hc1d4039d, 32'hc1982f26} /* (16, 24, 29) {real, imag} */,
  {32'hc17591aa, 32'h41ed88b8} /* (16, 24, 28) {real, imag} */,
  {32'h41c5adfe, 32'h41cce61d} /* (16, 24, 27) {real, imag} */,
  {32'h41a3aa82, 32'h41d4960a} /* (16, 24, 26) {real, imag} */,
  {32'h4107a7cf, 32'hc112292a} /* (16, 24, 25) {real, imag} */,
  {32'hc1a11386, 32'h404a7104} /* (16, 24, 24) {real, imag} */,
  {32'hc03b29ef, 32'hc1d385bc} /* (16, 24, 23) {real, imag} */,
  {32'hc1135286, 32'hc1061ae2} /* (16, 24, 22) {real, imag} */,
  {32'hc0483eda, 32'h40aab916} /* (16, 24, 21) {real, imag} */,
  {32'h41070767, 32'hc0434eb7} /* (16, 24, 20) {real, imag} */,
  {32'hc0e55e2c, 32'hbfc4d23a} /* (16, 24, 19) {real, imag} */,
  {32'h3f701230, 32'hbeed1ea0} /* (16, 24, 18) {real, imag} */,
  {32'h4017bb30, 32'hbef2ce00} /* (16, 24, 17) {real, imag} */,
  {32'hc0f2592e, 32'hbefb1540} /* (16, 24, 16) {real, imag} */,
  {32'h40e96b78, 32'hc05b46c0} /* (16, 24, 15) {real, imag} */,
  {32'h3dec9700, 32'h41298573} /* (16, 24, 14) {real, imag} */,
  {32'h4023b938, 32'hc0b48a9c} /* (16, 24, 13) {real, imag} */,
  {32'h40b9cce4, 32'h40532bf7} /* (16, 24, 12) {real, imag} */,
  {32'hc0bbc295, 32'h40d997a2} /* (16, 24, 11) {real, imag} */,
  {32'hc1141a3a, 32'hc11816e0} /* (16, 24, 10) {real, imag} */,
  {32'h400f9cd9, 32'h413fd570} /* (16, 24, 9) {real, imag} */,
  {32'h413b2378, 32'hc03d1fd6} /* (16, 24, 8) {real, imag} */,
  {32'hbf27346c, 32'hc0a027b5} /* (16, 24, 7) {real, imag} */,
  {32'hc16d2ae0, 32'h40254d24} /* (16, 24, 6) {real, imag} */,
  {32'hc156f450, 32'hc1311f8e} /* (16, 24, 5) {real, imag} */,
  {32'h40505a46, 32'h4195b578} /* (16, 24, 4) {real, imag} */,
  {32'hc1e48477, 32'h3e8362e0} /* (16, 24, 3) {real, imag} */,
  {32'hbf10dd40, 32'h41ec85f4} /* (16, 24, 2) {real, imag} */,
  {32'h41f3d08c, 32'hc22d602e} /* (16, 24, 1) {real, imag} */,
  {32'hc118f6bd, 32'hc0a365a4} /* (16, 24, 0) {real, imag} */,
  {32'hc1a2bdd5, 32'hc16d6620} /* (16, 23, 31) {real, imag} */,
  {32'h41111679, 32'hc1ed7817} /* (16, 23, 30) {real, imag} */,
  {32'h41b6c5d8, 32'hc175b06e} /* (16, 23, 29) {real, imag} */,
  {32'hbf7a91f0, 32'h40da6fc8} /* (16, 23, 28) {real, imag} */,
  {32'h3f9e5650, 32'h4158e5ba} /* (16, 23, 27) {real, imag} */,
  {32'h419ac2cc, 32'hc0cf07ae} /* (16, 23, 26) {real, imag} */,
  {32'h4102d1ff, 32'hbfe5ddfc} /* (16, 23, 25) {real, imag} */,
  {32'hc1800206, 32'hc1af3618} /* (16, 23, 24) {real, imag} */,
  {32'h408431fa, 32'h40c6624b} /* (16, 23, 23) {real, imag} */,
  {32'hc133d7ed, 32'h3f48c870} /* (16, 23, 22) {real, imag} */,
  {32'hc0f65989, 32'hc08b0642} /* (16, 23, 21) {real, imag} */,
  {32'h40249e4a, 32'h40b1d67e} /* (16, 23, 20) {real, imag} */,
  {32'hc012cf1c, 32'h40e0a412} /* (16, 23, 19) {real, imag} */,
  {32'hc135fd72, 32'hbee23fa8} /* (16, 23, 18) {real, imag} */,
  {32'h3facdbac, 32'hc10c354e} /* (16, 23, 17) {real, imag} */,
  {32'hc0a263a1, 32'h402f1020} /* (16, 23, 16) {real, imag} */,
  {32'hbf4d52a9, 32'hc0377f82} /* (16, 23, 15) {real, imag} */,
  {32'h40ff578c, 32'h3e4ca450} /* (16, 23, 14) {real, imag} */,
  {32'hc15f5e0f, 32'h40b804c0} /* (16, 23, 13) {real, imag} */,
  {32'h3f5f6cb8, 32'hc153d3dd} /* (16, 23, 12) {real, imag} */,
  {32'hc15a1b14, 32'hc11e71ca} /* (16, 23, 11) {real, imag} */,
  {32'h3e66f580, 32'hc1792c91} /* (16, 23, 10) {real, imag} */,
  {32'hc107b960, 32'hc097af8b} /* (16, 23, 9) {real, imag} */,
  {32'hc189fde6, 32'h414349b0} /* (16, 23, 8) {real, imag} */,
  {32'h40d7a33c, 32'hc0bfdb99} /* (16, 23, 7) {real, imag} */,
  {32'h3f6fab80, 32'h41132435} /* (16, 23, 6) {real, imag} */,
  {32'h41982895, 32'h41308a8e} /* (16, 23, 5) {real, imag} */,
  {32'hc1283420, 32'h3fd4c452} /* (16, 23, 4) {real, imag} */,
  {32'hc18af91e, 32'hc09d60b3} /* (16, 23, 3) {real, imag} */,
  {32'hc1ac29ee, 32'hc190d8e7} /* (16, 23, 2) {real, imag} */,
  {32'h41be2f9f, 32'hc200f10a} /* (16, 23, 1) {real, imag} */,
  {32'h3ecb5410, 32'hc1addd9a} /* (16, 23, 0) {real, imag} */,
  {32'hc1b1e0a6, 32'h412d78a9} /* (16, 22, 31) {real, imag} */,
  {32'hc0a9827e, 32'hc1668ab0} /* (16, 22, 30) {real, imag} */,
  {32'hc1c03608, 32'h3f9a3ed8} /* (16, 22, 29) {real, imag} */,
  {32'hc105318c, 32'h4188b9ca} /* (16, 22, 28) {real, imag} */,
  {32'hbfb10ff6, 32'hc13d3804} /* (16, 22, 27) {real, imag} */,
  {32'h3fe5aa34, 32'hc1f358e4} /* (16, 22, 26) {real, imag} */,
  {32'h3fb68208, 32'hc0c6ad38} /* (16, 22, 25) {real, imag} */,
  {32'h40aee09f, 32'h41094ca8} /* (16, 22, 24) {real, imag} */,
  {32'hc1505442, 32'hc0e18806} /* (16, 22, 23) {real, imag} */,
  {32'hbfc846b5, 32'hc00e8a4e} /* (16, 22, 22) {real, imag} */,
  {32'h41532d6e, 32'h40a6d723} /* (16, 22, 21) {real, imag} */,
  {32'h3ffa3b58, 32'h40ed9f16} /* (16, 22, 20) {real, imag} */,
  {32'h409403d3, 32'hc0ab4e81} /* (16, 22, 19) {real, imag} */,
  {32'hbf3f5d54, 32'hc0ad6239} /* (16, 22, 18) {real, imag} */,
  {32'hbf045c60, 32'hc016ce7e} /* (16, 22, 17) {real, imag} */,
  {32'hbdc41e00, 32'hc0aa9dab} /* (16, 22, 16) {real, imag} */,
  {32'h3f7bcf50, 32'h408a4727} /* (16, 22, 15) {real, imag} */,
  {32'hc00b8cdb, 32'hc05c1092} /* (16, 22, 14) {real, imag} */,
  {32'hbe1ce4e0, 32'hc0e1ccb1} /* (16, 22, 13) {real, imag} */,
  {32'h40fe3416, 32'h40355d6c} /* (16, 22, 12) {real, imag} */,
  {32'hbf98b054, 32'h4182448d} /* (16, 22, 11) {real, imag} */,
  {32'h405c1d48, 32'h40a220bd} /* (16, 22, 10) {real, imag} */,
  {32'h40abd7e3, 32'hc112db07} /* (16, 22, 9) {real, imag} */,
  {32'hc0b8c339, 32'h40ce9db6} /* (16, 22, 8) {real, imag} */,
  {32'hc13de1f6, 32'h40c07120} /* (16, 22, 7) {real, imag} */,
  {32'hc0ff9eaf, 32'h41a42528} /* (16, 22, 6) {real, imag} */,
  {32'h40c4ec00, 32'hc1152c90} /* (16, 22, 5) {real, imag} */,
  {32'hc1c0520e, 32'h40903b94} /* (16, 22, 4) {real, imag} */,
  {32'hc182f780, 32'hc10adb0c} /* (16, 22, 3) {real, imag} */,
  {32'hc0b90a6e, 32'h413482f4} /* (16, 22, 2) {real, imag} */,
  {32'hc0c75ec0, 32'hc1612f43} /* (16, 22, 1) {real, imag} */,
  {32'h41f15d1a, 32'h41a03faf} /* (16, 22, 0) {real, imag} */,
  {32'hc08473bb, 32'hc1478a12} /* (16, 21, 31) {real, imag} */,
  {32'h418e6b05, 32'hc094e6ca} /* (16, 21, 30) {real, imag} */,
  {32'hc11b550a, 32'hc1de55a5} /* (16, 21, 29) {real, imag} */,
  {32'h3f8914b0, 32'hc197abaa} /* (16, 21, 28) {real, imag} */,
  {32'hc0c6827f, 32'h410bab55} /* (16, 21, 27) {real, imag} */,
  {32'hbea62630, 32'h4036ddf8} /* (16, 21, 26) {real, imag} */,
  {32'h414c407f, 32'hbf366b58} /* (16, 21, 25) {real, imag} */,
  {32'hc0f4bbb4, 32'h40f0a5b2} /* (16, 21, 24) {real, imag} */,
  {32'hc10423dd, 32'hc10d2cfc} /* (16, 21, 23) {real, imag} */,
  {32'hc082f83e, 32'hc128df5e} /* (16, 21, 22) {real, imag} */,
  {32'h3e7da890, 32'h40d03046} /* (16, 21, 21) {real, imag} */,
  {32'h3e25b3a0, 32'hc0393fde} /* (16, 21, 20) {real, imag} */,
  {32'hc08a14d6, 32'hc0443946} /* (16, 21, 19) {real, imag} */,
  {32'h410b0b9b, 32'hc0d2f494} /* (16, 21, 18) {real, imag} */,
  {32'h4032d77d, 32'h3e87ea28} /* (16, 21, 17) {real, imag} */,
  {32'hbff09942, 32'hbd83f700} /* (16, 21, 16) {real, imag} */,
  {32'hc007d4c3, 32'hc02b5019} /* (16, 21, 15) {real, imag} */,
  {32'hbf7b85a0, 32'h3f178af0} /* (16, 21, 14) {real, imag} */,
  {32'h3fcbf50a, 32'hbf4f41d8} /* (16, 21, 13) {real, imag} */,
  {32'hc0a14c59, 32'hbd800540} /* (16, 21, 12) {real, imag} */,
  {32'hbf859f0a, 32'h4063cfc4} /* (16, 21, 11) {real, imag} */,
  {32'h3f1e6504, 32'h40611e54} /* (16, 21, 10) {real, imag} */,
  {32'h4094e06a, 32'h3e3a9de0} /* (16, 21, 9) {real, imag} */,
  {32'h40bd9786, 32'hc1127fb7} /* (16, 21, 8) {real, imag} */,
  {32'h4111d979, 32'h4090aa51} /* (16, 21, 7) {real, imag} */,
  {32'h410f64d0, 32'h413ff487} /* (16, 21, 6) {real, imag} */,
  {32'h40ae4a35, 32'h40518f0c} /* (16, 21, 5) {real, imag} */,
  {32'h3e05ef90, 32'hc0399cec} /* (16, 21, 4) {real, imag} */,
  {32'hc199d796, 32'h415ba87a} /* (16, 21, 3) {real, imag} */,
  {32'hc0ad519d, 32'hc101e67c} /* (16, 21, 2) {real, imag} */,
  {32'hc0bde68d, 32'hc053b316} /* (16, 21, 1) {real, imag} */,
  {32'hc011af8d, 32'h41844f28} /* (16, 21, 0) {real, imag} */,
  {32'hc1450fc5, 32'h4121a660} /* (16, 20, 31) {real, imag} */,
  {32'hc10bbcde, 32'hc12440f6} /* (16, 20, 30) {real, imag} */,
  {32'h40fa6850, 32'hbea5fb40} /* (16, 20, 29) {real, imag} */,
  {32'hbf448dc0, 32'hc1a0b5da} /* (16, 20, 28) {real, imag} */,
  {32'hc08acd9b, 32'hc13e8245} /* (16, 20, 27) {real, imag} */,
  {32'hc080b7ab, 32'hbf97b678} /* (16, 20, 26) {real, imag} */,
  {32'h4198bc1c, 32'hc1467e43} /* (16, 20, 25) {real, imag} */,
  {32'h3e6ec3b0, 32'hc1adbeff} /* (16, 20, 24) {real, imag} */,
  {32'hc02cec60, 32'hc100ec4a} /* (16, 20, 23) {real, imag} */,
  {32'h3f6ae72c, 32'h4054caa7} /* (16, 20, 22) {real, imag} */,
  {32'hc1319804, 32'hbfb3c144} /* (16, 20, 21) {real, imag} */,
  {32'h40c4164a, 32'h3fbfb5ce} /* (16, 20, 20) {real, imag} */,
  {32'h40c13a62, 32'hc01a4b9a} /* (16, 20, 19) {real, imag} */,
  {32'hbff5fb40, 32'h4098e09c} /* (16, 20, 18) {real, imag} */,
  {32'hc0990a12, 32'h3fdb62b2} /* (16, 20, 17) {real, imag} */,
  {32'hbfe1b638, 32'hbf0e5180} /* (16, 20, 16) {real, imag} */,
  {32'hbf3db34c, 32'h3f2a913c} /* (16, 20, 15) {real, imag} */,
  {32'hbf811a66, 32'hc0a84392} /* (16, 20, 14) {real, imag} */,
  {32'h404a773d, 32'hc0dd8573} /* (16, 20, 13) {real, imag} */,
  {32'h400c477b, 32'h411137d8} /* (16, 20, 12) {real, imag} */,
  {32'h403b6c3a, 32'h3df86740} /* (16, 20, 11) {real, imag} */,
  {32'h40d5e4a6, 32'hbd15e9c0} /* (16, 20, 10) {real, imag} */,
  {32'hc1360326, 32'hc0873f90} /* (16, 20, 9) {real, imag} */,
  {32'hbf4cdcac, 32'hc0905850} /* (16, 20, 8) {real, imag} */,
  {32'hc122e38e, 32'hc13cc06b} /* (16, 20, 7) {real, imag} */,
  {32'hc0fb9e11, 32'h40441954} /* (16, 20, 6) {real, imag} */,
  {32'hc1540d54, 32'h3f773000} /* (16, 20, 5) {real, imag} */,
  {32'h418f1696, 32'hc0af0cb6} /* (16, 20, 4) {real, imag} */,
  {32'h3eaac088, 32'h417e1236} /* (16, 20, 3) {real, imag} */,
  {32'hbf1e2b88, 32'hc1429eea} /* (16, 20, 2) {real, imag} */,
  {32'hc1198715, 32'h3f0d4338} /* (16, 20, 1) {real, imag} */,
  {32'h41c5055e, 32'h412c5442} /* (16, 20, 0) {real, imag} */,
  {32'h41889d91, 32'hc1b5f55e} /* (16, 19, 31) {real, imag} */,
  {32'h41664cdf, 32'h41611ca0} /* (16, 19, 30) {real, imag} */,
  {32'h40dd276e, 32'h3f877602} /* (16, 19, 29) {real, imag} */,
  {32'hc1871ae8, 32'hc14b8cf6} /* (16, 19, 28) {real, imag} */,
  {32'h40b779ee, 32'h40c3a549} /* (16, 19, 27) {real, imag} */,
  {32'h41226351, 32'h408b97b6} /* (16, 19, 26) {real, imag} */,
  {32'hc0b95a3e, 32'h40080ffc} /* (16, 19, 25) {real, imag} */,
  {32'h40ad5c08, 32'hbfafc04c} /* (16, 19, 24) {real, imag} */,
  {32'h3f956fd4, 32'hc08f0446} /* (16, 19, 23) {real, imag} */,
  {32'h401c69c1, 32'h40c26e22} /* (16, 19, 22) {real, imag} */,
  {32'hc04271f6, 32'h40c45ceb} /* (16, 19, 21) {real, imag} */,
  {32'hc09bf653, 32'hbf8df1dc} /* (16, 19, 20) {real, imag} */,
  {32'hc01319c6, 32'hc103127d} /* (16, 19, 19) {real, imag} */,
  {32'hbd107f80, 32'h3ae5f000} /* (16, 19, 18) {real, imag} */,
  {32'hc0097964, 32'h40c28909} /* (16, 19, 17) {real, imag} */,
  {32'h405ea862, 32'hbf7f8d82} /* (16, 19, 16) {real, imag} */,
  {32'h3ee3b1c0, 32'hbfa9b30c} /* (16, 19, 15) {real, imag} */,
  {32'h400fc6fa, 32'h3e273480} /* (16, 19, 14) {real, imag} */,
  {32'hc02cf160, 32'h40140454} /* (16, 19, 13) {real, imag} */,
  {32'hbfffd4c5, 32'h40385b3c} /* (16, 19, 12) {real, imag} */,
  {32'h40eeafc9, 32'h40b664a5} /* (16, 19, 11) {real, imag} */,
  {32'hbfe50c56, 32'hc00ff0d9} /* (16, 19, 10) {real, imag} */,
  {32'hc0c580ac, 32'h3fd1bc48} /* (16, 19, 9) {real, imag} */,
  {32'h404da530, 32'hc0b8dd2b} /* (16, 19, 8) {real, imag} */,
  {32'h414a46d3, 32'hc1c04894} /* (16, 19, 7) {real, imag} */,
  {32'hc14cdbb3, 32'h3f5d847c} /* (16, 19, 6) {real, imag} */,
  {32'hc15c6973, 32'h405a547e} /* (16, 19, 5) {real, imag} */,
  {32'hc12c994d, 32'h40113980} /* (16, 19, 4) {real, imag} */,
  {32'h414f7b87, 32'h3f87d61e} /* (16, 19, 3) {real, imag} */,
  {32'h418ec774, 32'hbf949220} /* (16, 19, 2) {real, imag} */,
  {32'hc1258152, 32'h419f0416} /* (16, 19, 1) {real, imag} */,
  {32'hbde57cf0, 32'hc097b200} /* (16, 19, 0) {real, imag} */,
  {32'hc09050aa, 32'hc17769de} /* (16, 18, 31) {real, imag} */,
  {32'hc1579108, 32'hc0956685} /* (16, 18, 30) {real, imag} */,
  {32'h4150f089, 32'hc0e31398} /* (16, 18, 29) {real, imag} */,
  {32'hc113b2c6, 32'hc0a000e9} /* (16, 18, 28) {real, imag} */,
  {32'hc03262a6, 32'h4109de10} /* (16, 18, 27) {real, imag} */,
  {32'hc0f84b69, 32'hc093e4c2} /* (16, 18, 26) {real, imag} */,
  {32'hc0098a57, 32'h40fd0bba} /* (16, 18, 25) {real, imag} */,
  {32'hc1715ddd, 32'h408868cc} /* (16, 18, 24) {real, imag} */,
  {32'h4087d10a, 32'h3f627dea} /* (16, 18, 23) {real, imag} */,
  {32'hc089a576, 32'h3f88826e} /* (16, 18, 22) {real, imag} */,
  {32'hbf940035, 32'hc0a2d521} /* (16, 18, 21) {real, imag} */,
  {32'h3f70bfa4, 32'h409bbd63} /* (16, 18, 20) {real, imag} */,
  {32'h4008cc5d, 32'h3fb2ad62} /* (16, 18, 19) {real, imag} */,
  {32'h405ef0dd, 32'h3f5171fe} /* (16, 18, 18) {real, imag} */,
  {32'h3f942e23, 32'hc06a842e} /* (16, 18, 17) {real, imag} */,
  {32'hbf9f9504, 32'h4032bfde} /* (16, 18, 16) {real, imag} */,
  {32'h4005b322, 32'hbe880610} /* (16, 18, 15) {real, imag} */,
  {32'hbfd1584e, 32'hbfe7a6a7} /* (16, 18, 14) {real, imag} */,
  {32'hbfc9ee96, 32'hc0196ac3} /* (16, 18, 13) {real, imag} */,
  {32'h3fe8547e, 32'hbfd16b37} /* (16, 18, 12) {real, imag} */,
  {32'hc0026b2e, 32'h40184e32} /* (16, 18, 11) {real, imag} */,
  {32'hc0a836e8, 32'h3ea473e8} /* (16, 18, 10) {real, imag} */,
  {32'hbed864f8, 32'h3fb330eb} /* (16, 18, 9) {real, imag} */,
  {32'hc03e5694, 32'h4069ac20} /* (16, 18, 8) {real, imag} */,
  {32'h40f67056, 32'h408de9c6} /* (16, 18, 7) {real, imag} */,
  {32'h4003d656, 32'h4045ab59} /* (16, 18, 6) {real, imag} */,
  {32'h4035c242, 32'h40d5556d} /* (16, 18, 5) {real, imag} */,
  {32'h40e3fd94, 32'h414bac1e} /* (16, 18, 4) {real, imag} */,
  {32'hbed53ae0, 32'hc068c26f} /* (16, 18, 3) {real, imag} */,
  {32'h404a6d00, 32'h4013a8ea} /* (16, 18, 2) {real, imag} */,
  {32'h3fd1a1d9, 32'h40fb2254} /* (16, 18, 1) {real, imag} */,
  {32'h41440ce4, 32'hc0a1438a} /* (16, 18, 0) {real, imag} */,
  {32'hbf6a7038, 32'h4135b3f3} /* (16, 17, 31) {real, imag} */,
  {32'hc0f1803a, 32'h40e110e4} /* (16, 17, 30) {real, imag} */,
  {32'h4082966d, 32'hc0075dba} /* (16, 17, 29) {real, imag} */,
  {32'h40b9e3c0, 32'h409a4890} /* (16, 17, 28) {real, imag} */,
  {32'hc0be446d, 32'h4092f428} /* (16, 17, 27) {real, imag} */,
  {32'hc0ac012c, 32'hc08ddacb} /* (16, 17, 26) {real, imag} */,
  {32'h3f2a835c, 32'hc1209632} /* (16, 17, 25) {real, imag} */,
  {32'h3f29afe2, 32'hc01fe6ca} /* (16, 17, 24) {real, imag} */,
  {32'hc03eef9a, 32'hbf1b4968} /* (16, 17, 23) {real, imag} */,
  {32'hbf7b5c4a, 32'hc00be4a4} /* (16, 17, 22) {real, imag} */,
  {32'h4010806e, 32'h40a94bab} /* (16, 17, 21) {real, imag} */,
  {32'h3dcc5a20, 32'h3f168d76} /* (16, 17, 20) {real, imag} */,
  {32'h3ffdcfbe, 32'hbee8a434} /* (16, 17, 19) {real, imag} */,
  {32'hc056a5b8, 32'h3faf62fa} /* (16, 17, 18) {real, imag} */,
  {32'hc006cb56, 32'h3ef15fc4} /* (16, 17, 17) {real, imag} */,
  {32'h3fcdd5a8, 32'h3f248bd0} /* (16, 17, 16) {real, imag} */,
  {32'hbf3f35d0, 32'h3ff52e91} /* (16, 17, 15) {real, imag} */,
  {32'hbf4de750, 32'h3ff5f602} /* (16, 17, 14) {real, imag} */,
  {32'hbf5e7a01, 32'hc07e700c} /* (16, 17, 13) {real, imag} */,
  {32'hbfd42a2e, 32'h3fb1986f} /* (16, 17, 12) {real, imag} */,
  {32'h3fa6a88d, 32'hc0525bfa} /* (16, 17, 11) {real, imag} */,
  {32'h3f8286af, 32'hbd4b6e60} /* (16, 17, 10) {real, imag} */,
  {32'h40bf479d, 32'hbf3ee088} /* (16, 17, 9) {real, imag} */,
  {32'h404325ea, 32'h40b813a3} /* (16, 17, 8) {real, imag} */,
  {32'hc0e3f360, 32'h40027f26} /* (16, 17, 7) {real, imag} */,
  {32'hbf49a7dc, 32'hc084cac9} /* (16, 17, 6) {real, imag} */,
  {32'h41216e28, 32'h40ac4e92} /* (16, 17, 5) {real, imag} */,
  {32'hc1321398, 32'hc1133808} /* (16, 17, 4) {real, imag} */,
  {32'hc0866363, 32'hbea00b54} /* (16, 17, 3) {real, imag} */,
  {32'hc124179f, 32'hc04e300c} /* (16, 17, 2) {real, imag} */,
  {32'h40b3fbfe, 32'hc11faf0b} /* (16, 17, 1) {real, imag} */,
  {32'hc16dfa23, 32'h40ca04d0} /* (16, 17, 0) {real, imag} */,
  {32'hc08972c8, 32'hc09bd368} /* (16, 16, 31) {real, imag} */,
  {32'h408d97fa, 32'hc004c75d} /* (16, 16, 30) {real, imag} */,
  {32'hc1aa2bd0, 32'h403b666e} /* (16, 16, 29) {real, imag} */,
  {32'h4090ea75, 32'h4114b927} /* (16, 16, 28) {real, imag} */,
  {32'h3f59767c, 32'hbfc71e60} /* (16, 16, 27) {real, imag} */,
  {32'h3fefb737, 32'hbfa1e8c0} /* (16, 16, 26) {real, imag} */,
  {32'h40927f98, 32'h405f5c2b} /* (16, 16, 25) {real, imag} */,
  {32'hbf2e5296, 32'h3f4ecc44} /* (16, 16, 24) {real, imag} */,
  {32'hbe599740, 32'h3f6ee044} /* (16, 16, 23) {real, imag} */,
  {32'hbf5fde1e, 32'hbf585610} /* (16, 16, 22) {real, imag} */,
  {32'h3ff08672, 32'hbf09568f} /* (16, 16, 21) {real, imag} */,
  {32'h3db50dc0, 32'hc02b266d} /* (16, 16, 20) {real, imag} */,
  {32'h4034c50c, 32'h4019d3fc} /* (16, 16, 19) {real, imag} */,
  {32'hbf90e0c4, 32'hbfa20feb} /* (16, 16, 18) {real, imag} */,
  {32'h3fb96c0f, 32'hbf94f056} /* (16, 16, 17) {real, imag} */,
  {32'hc0500d44, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h3fb96c0f, 32'h3f94f056} /* (16, 16, 15) {real, imag} */,
  {32'hbf90e0c4, 32'h3fa20feb} /* (16, 16, 14) {real, imag} */,
  {32'h4034c50c, 32'hc019d3fc} /* (16, 16, 13) {real, imag} */,
  {32'h3db50dc0, 32'h402b266d} /* (16, 16, 12) {real, imag} */,
  {32'h3ff08672, 32'h3f09568f} /* (16, 16, 11) {real, imag} */,
  {32'hbf5fde1e, 32'h3f585610} /* (16, 16, 10) {real, imag} */,
  {32'hbe599740, 32'hbf6ee044} /* (16, 16, 9) {real, imag} */,
  {32'hbf2e5296, 32'hbf4ecc44} /* (16, 16, 8) {real, imag} */,
  {32'h40927f98, 32'hc05f5c2b} /* (16, 16, 7) {real, imag} */,
  {32'h3fefb737, 32'h3fa1e8c0} /* (16, 16, 6) {real, imag} */,
  {32'h3f59767c, 32'h3fc71e60} /* (16, 16, 5) {real, imag} */,
  {32'h4090ea75, 32'hc114b927} /* (16, 16, 4) {real, imag} */,
  {32'hc1aa2bd0, 32'hc03b666e} /* (16, 16, 3) {real, imag} */,
  {32'h408d97fa, 32'h4004c75d} /* (16, 16, 2) {real, imag} */,
  {32'hc08972c8, 32'h409bd368} /* (16, 16, 1) {real, imag} */,
  {32'h410522bb, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h40b3fbfe, 32'h411faf0b} /* (16, 15, 31) {real, imag} */,
  {32'hc124179f, 32'h404e300c} /* (16, 15, 30) {real, imag} */,
  {32'hc0866363, 32'h3ea00b54} /* (16, 15, 29) {real, imag} */,
  {32'hc1321398, 32'h41133808} /* (16, 15, 28) {real, imag} */,
  {32'h41216e28, 32'hc0ac4e92} /* (16, 15, 27) {real, imag} */,
  {32'hbf49a7dc, 32'h4084cac9} /* (16, 15, 26) {real, imag} */,
  {32'hc0e3f360, 32'hc0027f26} /* (16, 15, 25) {real, imag} */,
  {32'h404325ea, 32'hc0b813a3} /* (16, 15, 24) {real, imag} */,
  {32'h40bf479d, 32'h3f3ee088} /* (16, 15, 23) {real, imag} */,
  {32'h3f8286af, 32'h3d4b6e60} /* (16, 15, 22) {real, imag} */,
  {32'h3fa6a88d, 32'h40525bfa} /* (16, 15, 21) {real, imag} */,
  {32'hbfd42a2e, 32'hbfb1986f} /* (16, 15, 20) {real, imag} */,
  {32'hbf5e7a01, 32'h407e700c} /* (16, 15, 19) {real, imag} */,
  {32'hbf4de750, 32'hbff5f602} /* (16, 15, 18) {real, imag} */,
  {32'hbf3f35d0, 32'hbff52e91} /* (16, 15, 17) {real, imag} */,
  {32'h3fcdd5a8, 32'hbf248bd0} /* (16, 15, 16) {real, imag} */,
  {32'hc006cb56, 32'hbef15fc4} /* (16, 15, 15) {real, imag} */,
  {32'hc056a5b8, 32'hbfaf62fa} /* (16, 15, 14) {real, imag} */,
  {32'h3ffdcfbe, 32'h3ee8a434} /* (16, 15, 13) {real, imag} */,
  {32'h3dcc5a20, 32'hbf168d76} /* (16, 15, 12) {real, imag} */,
  {32'h4010806e, 32'hc0a94bab} /* (16, 15, 11) {real, imag} */,
  {32'hbf7b5c4a, 32'h400be4a4} /* (16, 15, 10) {real, imag} */,
  {32'hc03eef9a, 32'h3f1b4968} /* (16, 15, 9) {real, imag} */,
  {32'h3f29afe2, 32'h401fe6ca} /* (16, 15, 8) {real, imag} */,
  {32'h3f2a835c, 32'h41209632} /* (16, 15, 7) {real, imag} */,
  {32'hc0ac012c, 32'h408ddacb} /* (16, 15, 6) {real, imag} */,
  {32'hc0be446d, 32'hc092f428} /* (16, 15, 5) {real, imag} */,
  {32'h40b9e3c0, 32'hc09a4890} /* (16, 15, 4) {real, imag} */,
  {32'h4082966d, 32'h40075dba} /* (16, 15, 3) {real, imag} */,
  {32'hc0f1803a, 32'hc0e110e4} /* (16, 15, 2) {real, imag} */,
  {32'hbf6a7038, 32'hc135b3f3} /* (16, 15, 1) {real, imag} */,
  {32'hc16dfa23, 32'hc0ca04d0} /* (16, 15, 0) {real, imag} */,
  {32'h3fd1a1d9, 32'hc0fb2254} /* (16, 14, 31) {real, imag} */,
  {32'h404a6d00, 32'hc013a8ea} /* (16, 14, 30) {real, imag} */,
  {32'hbed53ae0, 32'h4068c26f} /* (16, 14, 29) {real, imag} */,
  {32'h40e3fd94, 32'hc14bac1e} /* (16, 14, 28) {real, imag} */,
  {32'h4035c242, 32'hc0d5556d} /* (16, 14, 27) {real, imag} */,
  {32'h4003d656, 32'hc045ab59} /* (16, 14, 26) {real, imag} */,
  {32'h40f67056, 32'hc08de9c6} /* (16, 14, 25) {real, imag} */,
  {32'hc03e5694, 32'hc069ac20} /* (16, 14, 24) {real, imag} */,
  {32'hbed864f8, 32'hbfb330eb} /* (16, 14, 23) {real, imag} */,
  {32'hc0a836e8, 32'hbea473e8} /* (16, 14, 22) {real, imag} */,
  {32'hc0026b2e, 32'hc0184e32} /* (16, 14, 21) {real, imag} */,
  {32'h3fe8547e, 32'h3fd16b37} /* (16, 14, 20) {real, imag} */,
  {32'hbfc9ee96, 32'h40196ac3} /* (16, 14, 19) {real, imag} */,
  {32'hbfd1584e, 32'h3fe7a6a7} /* (16, 14, 18) {real, imag} */,
  {32'h4005b322, 32'h3e880610} /* (16, 14, 17) {real, imag} */,
  {32'hbf9f9504, 32'hc032bfde} /* (16, 14, 16) {real, imag} */,
  {32'h3f942e23, 32'h406a842e} /* (16, 14, 15) {real, imag} */,
  {32'h405ef0dd, 32'hbf5171fe} /* (16, 14, 14) {real, imag} */,
  {32'h4008cc5d, 32'hbfb2ad62} /* (16, 14, 13) {real, imag} */,
  {32'h3f70bfa4, 32'hc09bbd63} /* (16, 14, 12) {real, imag} */,
  {32'hbf940035, 32'h40a2d521} /* (16, 14, 11) {real, imag} */,
  {32'hc089a576, 32'hbf88826e} /* (16, 14, 10) {real, imag} */,
  {32'h4087d10a, 32'hbf627dea} /* (16, 14, 9) {real, imag} */,
  {32'hc1715ddd, 32'hc08868cc} /* (16, 14, 8) {real, imag} */,
  {32'hc0098a57, 32'hc0fd0bba} /* (16, 14, 7) {real, imag} */,
  {32'hc0f84b69, 32'h4093e4c2} /* (16, 14, 6) {real, imag} */,
  {32'hc03262a6, 32'hc109de10} /* (16, 14, 5) {real, imag} */,
  {32'hc113b2c6, 32'h40a000e9} /* (16, 14, 4) {real, imag} */,
  {32'h4150f089, 32'h40e31398} /* (16, 14, 3) {real, imag} */,
  {32'hc1579108, 32'h40956685} /* (16, 14, 2) {real, imag} */,
  {32'hc09050aa, 32'h417769de} /* (16, 14, 1) {real, imag} */,
  {32'h41440ce4, 32'h40a1438a} /* (16, 14, 0) {real, imag} */,
  {32'hc1258152, 32'hc19f0416} /* (16, 13, 31) {real, imag} */,
  {32'h418ec774, 32'h3f949220} /* (16, 13, 30) {real, imag} */,
  {32'h414f7b87, 32'hbf87d61e} /* (16, 13, 29) {real, imag} */,
  {32'hc12c994d, 32'hc0113980} /* (16, 13, 28) {real, imag} */,
  {32'hc15c6973, 32'hc05a547e} /* (16, 13, 27) {real, imag} */,
  {32'hc14cdbb3, 32'hbf5d847c} /* (16, 13, 26) {real, imag} */,
  {32'h414a46d3, 32'h41c04894} /* (16, 13, 25) {real, imag} */,
  {32'h404da530, 32'h40b8dd2b} /* (16, 13, 24) {real, imag} */,
  {32'hc0c580ac, 32'hbfd1bc48} /* (16, 13, 23) {real, imag} */,
  {32'hbfe50c56, 32'h400ff0d9} /* (16, 13, 22) {real, imag} */,
  {32'h40eeafc9, 32'hc0b664a5} /* (16, 13, 21) {real, imag} */,
  {32'hbfffd4c5, 32'hc0385b3c} /* (16, 13, 20) {real, imag} */,
  {32'hc02cf160, 32'hc0140454} /* (16, 13, 19) {real, imag} */,
  {32'h400fc6fa, 32'hbe273480} /* (16, 13, 18) {real, imag} */,
  {32'h3ee3b1c0, 32'h3fa9b30c} /* (16, 13, 17) {real, imag} */,
  {32'h405ea862, 32'h3f7f8d82} /* (16, 13, 16) {real, imag} */,
  {32'hc0097964, 32'hc0c28909} /* (16, 13, 15) {real, imag} */,
  {32'hbd107f80, 32'hbae5f000} /* (16, 13, 14) {real, imag} */,
  {32'hc01319c6, 32'h4103127d} /* (16, 13, 13) {real, imag} */,
  {32'hc09bf653, 32'h3f8df1dc} /* (16, 13, 12) {real, imag} */,
  {32'hc04271f6, 32'hc0c45ceb} /* (16, 13, 11) {real, imag} */,
  {32'h401c69c1, 32'hc0c26e22} /* (16, 13, 10) {real, imag} */,
  {32'h3f956fd4, 32'h408f0446} /* (16, 13, 9) {real, imag} */,
  {32'h40ad5c08, 32'h3fafc04c} /* (16, 13, 8) {real, imag} */,
  {32'hc0b95a3e, 32'hc0080ffc} /* (16, 13, 7) {real, imag} */,
  {32'h41226351, 32'hc08b97b6} /* (16, 13, 6) {real, imag} */,
  {32'h40b779ee, 32'hc0c3a549} /* (16, 13, 5) {real, imag} */,
  {32'hc1871ae8, 32'h414b8cf6} /* (16, 13, 4) {real, imag} */,
  {32'h40dd276e, 32'hbf877602} /* (16, 13, 3) {real, imag} */,
  {32'h41664cdf, 32'hc1611ca0} /* (16, 13, 2) {real, imag} */,
  {32'h41889d91, 32'h41b5f55e} /* (16, 13, 1) {real, imag} */,
  {32'hbde57cf0, 32'h4097b200} /* (16, 13, 0) {real, imag} */,
  {32'hc1198715, 32'hbf0d4338} /* (16, 12, 31) {real, imag} */,
  {32'hbf1e2b88, 32'h41429eea} /* (16, 12, 30) {real, imag} */,
  {32'h3eaac088, 32'hc17e1236} /* (16, 12, 29) {real, imag} */,
  {32'h418f1696, 32'h40af0cb6} /* (16, 12, 28) {real, imag} */,
  {32'hc1540d54, 32'hbf773000} /* (16, 12, 27) {real, imag} */,
  {32'hc0fb9e11, 32'hc0441954} /* (16, 12, 26) {real, imag} */,
  {32'hc122e38e, 32'h413cc06b} /* (16, 12, 25) {real, imag} */,
  {32'hbf4cdcac, 32'h40905850} /* (16, 12, 24) {real, imag} */,
  {32'hc1360326, 32'h40873f90} /* (16, 12, 23) {real, imag} */,
  {32'h40d5e4a6, 32'h3d15e9c0} /* (16, 12, 22) {real, imag} */,
  {32'h403b6c3a, 32'hbdf86740} /* (16, 12, 21) {real, imag} */,
  {32'h400c477b, 32'hc11137d8} /* (16, 12, 20) {real, imag} */,
  {32'h404a773d, 32'h40dd8573} /* (16, 12, 19) {real, imag} */,
  {32'hbf811a66, 32'h40a84392} /* (16, 12, 18) {real, imag} */,
  {32'hbf3db34c, 32'hbf2a913c} /* (16, 12, 17) {real, imag} */,
  {32'hbfe1b638, 32'h3f0e5180} /* (16, 12, 16) {real, imag} */,
  {32'hc0990a12, 32'hbfdb62b2} /* (16, 12, 15) {real, imag} */,
  {32'hbff5fb40, 32'hc098e09c} /* (16, 12, 14) {real, imag} */,
  {32'h40c13a62, 32'h401a4b9a} /* (16, 12, 13) {real, imag} */,
  {32'h40c4164a, 32'hbfbfb5ce} /* (16, 12, 12) {real, imag} */,
  {32'hc1319804, 32'h3fb3c144} /* (16, 12, 11) {real, imag} */,
  {32'h3f6ae72c, 32'hc054caa7} /* (16, 12, 10) {real, imag} */,
  {32'hc02cec60, 32'h4100ec4a} /* (16, 12, 9) {real, imag} */,
  {32'h3e6ec3b0, 32'h41adbeff} /* (16, 12, 8) {real, imag} */,
  {32'h4198bc1c, 32'h41467e43} /* (16, 12, 7) {real, imag} */,
  {32'hc080b7ab, 32'h3f97b678} /* (16, 12, 6) {real, imag} */,
  {32'hc08acd9b, 32'h413e8245} /* (16, 12, 5) {real, imag} */,
  {32'hbf448dc0, 32'h41a0b5da} /* (16, 12, 4) {real, imag} */,
  {32'h40fa6850, 32'h3ea5fb40} /* (16, 12, 3) {real, imag} */,
  {32'hc10bbcde, 32'h412440f6} /* (16, 12, 2) {real, imag} */,
  {32'hc1450fc5, 32'hc121a660} /* (16, 12, 1) {real, imag} */,
  {32'h41c5055e, 32'hc12c5442} /* (16, 12, 0) {real, imag} */,
  {32'hc0bde68d, 32'h4053b316} /* (16, 11, 31) {real, imag} */,
  {32'hc0ad519d, 32'h4101e67c} /* (16, 11, 30) {real, imag} */,
  {32'hc199d796, 32'hc15ba87a} /* (16, 11, 29) {real, imag} */,
  {32'h3e05ef90, 32'h40399cec} /* (16, 11, 28) {real, imag} */,
  {32'h40ae4a35, 32'hc0518f0c} /* (16, 11, 27) {real, imag} */,
  {32'h410f64d0, 32'hc13ff487} /* (16, 11, 26) {real, imag} */,
  {32'h4111d979, 32'hc090aa51} /* (16, 11, 25) {real, imag} */,
  {32'h40bd9786, 32'h41127fb7} /* (16, 11, 24) {real, imag} */,
  {32'h4094e06a, 32'hbe3a9de0} /* (16, 11, 23) {real, imag} */,
  {32'h3f1e6504, 32'hc0611e54} /* (16, 11, 22) {real, imag} */,
  {32'hbf859f0a, 32'hc063cfc4} /* (16, 11, 21) {real, imag} */,
  {32'hc0a14c59, 32'h3d800540} /* (16, 11, 20) {real, imag} */,
  {32'h3fcbf50a, 32'h3f4f41d8} /* (16, 11, 19) {real, imag} */,
  {32'hbf7b85a0, 32'hbf178af0} /* (16, 11, 18) {real, imag} */,
  {32'hc007d4c3, 32'h402b5019} /* (16, 11, 17) {real, imag} */,
  {32'hbff09942, 32'h3d83f700} /* (16, 11, 16) {real, imag} */,
  {32'h4032d77d, 32'hbe87ea28} /* (16, 11, 15) {real, imag} */,
  {32'h410b0b9b, 32'h40d2f494} /* (16, 11, 14) {real, imag} */,
  {32'hc08a14d6, 32'h40443946} /* (16, 11, 13) {real, imag} */,
  {32'h3e25b3a0, 32'h40393fde} /* (16, 11, 12) {real, imag} */,
  {32'h3e7da890, 32'hc0d03046} /* (16, 11, 11) {real, imag} */,
  {32'hc082f83e, 32'h4128df5e} /* (16, 11, 10) {real, imag} */,
  {32'hc10423dd, 32'h410d2cfc} /* (16, 11, 9) {real, imag} */,
  {32'hc0f4bbb4, 32'hc0f0a5b2} /* (16, 11, 8) {real, imag} */,
  {32'h414c407f, 32'h3f366b58} /* (16, 11, 7) {real, imag} */,
  {32'hbea62630, 32'hc036ddf8} /* (16, 11, 6) {real, imag} */,
  {32'hc0c6827f, 32'hc10bab55} /* (16, 11, 5) {real, imag} */,
  {32'h3f8914b0, 32'h4197abaa} /* (16, 11, 4) {real, imag} */,
  {32'hc11b550a, 32'h41de55a5} /* (16, 11, 3) {real, imag} */,
  {32'h418e6b05, 32'h4094e6ca} /* (16, 11, 2) {real, imag} */,
  {32'hc08473bb, 32'h41478a12} /* (16, 11, 1) {real, imag} */,
  {32'hc011af8d, 32'hc1844f28} /* (16, 11, 0) {real, imag} */,
  {32'hc0c75ec0, 32'h41612f43} /* (16, 10, 31) {real, imag} */,
  {32'hc0b90a6e, 32'hc13482f4} /* (16, 10, 30) {real, imag} */,
  {32'hc182f780, 32'h410adb0c} /* (16, 10, 29) {real, imag} */,
  {32'hc1c0520e, 32'hc0903b94} /* (16, 10, 28) {real, imag} */,
  {32'h40c4ec00, 32'h41152c90} /* (16, 10, 27) {real, imag} */,
  {32'hc0ff9eaf, 32'hc1a42528} /* (16, 10, 26) {real, imag} */,
  {32'hc13de1f6, 32'hc0c07120} /* (16, 10, 25) {real, imag} */,
  {32'hc0b8c339, 32'hc0ce9db6} /* (16, 10, 24) {real, imag} */,
  {32'h40abd7e3, 32'h4112db07} /* (16, 10, 23) {real, imag} */,
  {32'h405c1d48, 32'hc0a220bd} /* (16, 10, 22) {real, imag} */,
  {32'hbf98b054, 32'hc182448d} /* (16, 10, 21) {real, imag} */,
  {32'h40fe3416, 32'hc0355d6c} /* (16, 10, 20) {real, imag} */,
  {32'hbe1ce4e0, 32'h40e1ccb1} /* (16, 10, 19) {real, imag} */,
  {32'hc00b8cdb, 32'h405c1092} /* (16, 10, 18) {real, imag} */,
  {32'h3f7bcf50, 32'hc08a4727} /* (16, 10, 17) {real, imag} */,
  {32'hbdc41e00, 32'h40aa9dab} /* (16, 10, 16) {real, imag} */,
  {32'hbf045c60, 32'h4016ce7e} /* (16, 10, 15) {real, imag} */,
  {32'hbf3f5d54, 32'h40ad6239} /* (16, 10, 14) {real, imag} */,
  {32'h409403d3, 32'h40ab4e81} /* (16, 10, 13) {real, imag} */,
  {32'h3ffa3b58, 32'hc0ed9f16} /* (16, 10, 12) {real, imag} */,
  {32'h41532d6e, 32'hc0a6d723} /* (16, 10, 11) {real, imag} */,
  {32'hbfc846b5, 32'h400e8a4e} /* (16, 10, 10) {real, imag} */,
  {32'hc1505442, 32'h40e18806} /* (16, 10, 9) {real, imag} */,
  {32'h40aee09f, 32'hc1094ca8} /* (16, 10, 8) {real, imag} */,
  {32'h3fb68208, 32'h40c6ad38} /* (16, 10, 7) {real, imag} */,
  {32'h3fe5aa34, 32'h41f358e4} /* (16, 10, 6) {real, imag} */,
  {32'hbfb10ff6, 32'h413d3804} /* (16, 10, 5) {real, imag} */,
  {32'hc105318c, 32'hc188b9ca} /* (16, 10, 4) {real, imag} */,
  {32'hc1c03608, 32'hbf9a3ed8} /* (16, 10, 3) {real, imag} */,
  {32'hc0a9827e, 32'h41668ab0} /* (16, 10, 2) {real, imag} */,
  {32'hc1b1e0a6, 32'hc12d78a9} /* (16, 10, 1) {real, imag} */,
  {32'h41f15d1a, 32'hc1a03faf} /* (16, 10, 0) {real, imag} */,
  {32'h41be2f9f, 32'h4200f10a} /* (16, 9, 31) {real, imag} */,
  {32'hc1ac29ee, 32'h4190d8e7} /* (16, 9, 30) {real, imag} */,
  {32'hc18af91e, 32'h409d60b3} /* (16, 9, 29) {real, imag} */,
  {32'hc1283420, 32'hbfd4c452} /* (16, 9, 28) {real, imag} */,
  {32'h41982895, 32'hc1308a8e} /* (16, 9, 27) {real, imag} */,
  {32'h3f6fab80, 32'hc1132435} /* (16, 9, 26) {real, imag} */,
  {32'h40d7a33c, 32'h40bfdb99} /* (16, 9, 25) {real, imag} */,
  {32'hc189fde6, 32'hc14349b0} /* (16, 9, 24) {real, imag} */,
  {32'hc107b960, 32'h4097af8b} /* (16, 9, 23) {real, imag} */,
  {32'h3e66f580, 32'h41792c91} /* (16, 9, 22) {real, imag} */,
  {32'hc15a1b14, 32'h411e71ca} /* (16, 9, 21) {real, imag} */,
  {32'h3f5f6cb8, 32'h4153d3dd} /* (16, 9, 20) {real, imag} */,
  {32'hc15f5e0f, 32'hc0b804c0} /* (16, 9, 19) {real, imag} */,
  {32'h40ff578c, 32'hbe4ca450} /* (16, 9, 18) {real, imag} */,
  {32'hbf4d52a9, 32'h40377f82} /* (16, 9, 17) {real, imag} */,
  {32'hc0a263a1, 32'hc02f1020} /* (16, 9, 16) {real, imag} */,
  {32'h3facdbac, 32'h410c354e} /* (16, 9, 15) {real, imag} */,
  {32'hc135fd72, 32'h3ee23fa8} /* (16, 9, 14) {real, imag} */,
  {32'hc012cf1c, 32'hc0e0a412} /* (16, 9, 13) {real, imag} */,
  {32'h40249e4a, 32'hc0b1d67e} /* (16, 9, 12) {real, imag} */,
  {32'hc0f65989, 32'h408b0642} /* (16, 9, 11) {real, imag} */,
  {32'hc133d7ed, 32'hbf48c870} /* (16, 9, 10) {real, imag} */,
  {32'h408431fa, 32'hc0c6624b} /* (16, 9, 9) {real, imag} */,
  {32'hc1800206, 32'h41af3618} /* (16, 9, 8) {real, imag} */,
  {32'h4102d1ff, 32'h3fe5ddfc} /* (16, 9, 7) {real, imag} */,
  {32'h419ac2cc, 32'h40cf07ae} /* (16, 9, 6) {real, imag} */,
  {32'h3f9e5650, 32'hc158e5ba} /* (16, 9, 5) {real, imag} */,
  {32'hbf7a91f0, 32'hc0da6fc8} /* (16, 9, 4) {real, imag} */,
  {32'h41b6c5d8, 32'h4175b06e} /* (16, 9, 3) {real, imag} */,
  {32'h41111679, 32'h41ed7817} /* (16, 9, 2) {real, imag} */,
  {32'hc1a2bdd5, 32'h416d6620} /* (16, 9, 1) {real, imag} */,
  {32'h3ecb5410, 32'h41addd9a} /* (16, 9, 0) {real, imag} */,
  {32'h41f3d08c, 32'h422d602e} /* (16, 8, 31) {real, imag} */,
  {32'hbf10dd40, 32'hc1ec85f4} /* (16, 8, 30) {real, imag} */,
  {32'hc1e48477, 32'hbe8362e0} /* (16, 8, 29) {real, imag} */,
  {32'h40505a46, 32'hc195b578} /* (16, 8, 28) {real, imag} */,
  {32'hc156f450, 32'h41311f8e} /* (16, 8, 27) {real, imag} */,
  {32'hc16d2ae0, 32'hc0254d24} /* (16, 8, 26) {real, imag} */,
  {32'hbf27346c, 32'h40a027b5} /* (16, 8, 25) {real, imag} */,
  {32'h413b2378, 32'h403d1fd6} /* (16, 8, 24) {real, imag} */,
  {32'h400f9cd9, 32'hc13fd570} /* (16, 8, 23) {real, imag} */,
  {32'hc1141a3a, 32'h411816e0} /* (16, 8, 22) {real, imag} */,
  {32'hc0bbc295, 32'hc0d997a2} /* (16, 8, 21) {real, imag} */,
  {32'h40b9cce4, 32'hc0532bf7} /* (16, 8, 20) {real, imag} */,
  {32'h4023b938, 32'h40b48a9c} /* (16, 8, 19) {real, imag} */,
  {32'h3dec9700, 32'hc1298573} /* (16, 8, 18) {real, imag} */,
  {32'h40e96b78, 32'h405b46c0} /* (16, 8, 17) {real, imag} */,
  {32'hc0f2592e, 32'h3efb1540} /* (16, 8, 16) {real, imag} */,
  {32'h4017bb30, 32'h3ef2ce00} /* (16, 8, 15) {real, imag} */,
  {32'h3f701230, 32'h3eed1ea0} /* (16, 8, 14) {real, imag} */,
  {32'hc0e55e2c, 32'h3fc4d23a} /* (16, 8, 13) {real, imag} */,
  {32'h41070767, 32'h40434eb7} /* (16, 8, 12) {real, imag} */,
  {32'hc0483eda, 32'hc0aab916} /* (16, 8, 11) {real, imag} */,
  {32'hc1135286, 32'h41061ae2} /* (16, 8, 10) {real, imag} */,
  {32'hc03b29ef, 32'h41d385bc} /* (16, 8, 9) {real, imag} */,
  {32'hc1a11386, 32'hc04a7104} /* (16, 8, 8) {real, imag} */,
  {32'h4107a7cf, 32'h4112292a} /* (16, 8, 7) {real, imag} */,
  {32'h41a3aa82, 32'hc1d4960a} /* (16, 8, 6) {real, imag} */,
  {32'h41c5adfe, 32'hc1cce61d} /* (16, 8, 5) {real, imag} */,
  {32'hc17591aa, 32'hc1ed88b8} /* (16, 8, 4) {real, imag} */,
  {32'hc1d4039d, 32'h41982f26} /* (16, 8, 3) {real, imag} */,
  {32'hc11d2129, 32'h41b55160} /* (16, 8, 2) {real, imag} */,
  {32'hc17db0e0, 32'h41f4048c} /* (16, 8, 1) {real, imag} */,
  {32'hc118f6bd, 32'h40a365a4} /* (16, 8, 0) {real, imag} */,
  {32'hc0de19fe, 32'hc18b55d4} /* (16, 7, 31) {real, imag} */,
  {32'hbf6a06f8, 32'h416c927b} /* (16, 7, 30) {real, imag} */,
  {32'hc12d8080, 32'h4141f233} /* (16, 7, 29) {real, imag} */,
  {32'hc12f6230, 32'hc033c5a8} /* (16, 7, 28) {real, imag} */,
  {32'h40d79c54, 32'h411132f8} /* (16, 7, 27) {real, imag} */,
  {32'h41479c88, 32'hc1047630} /* (16, 7, 26) {real, imag} */,
  {32'hc18e67a7, 32'h4133e7ab} /* (16, 7, 25) {real, imag} */,
  {32'hc0c8415a, 32'h3f082bf0} /* (16, 7, 24) {real, imag} */,
  {32'h40b41e13, 32'hbe9e9760} /* (16, 7, 23) {real, imag} */,
  {32'hc19516f6, 32'hc147163d} /* (16, 7, 22) {real, imag} */,
  {32'h4110ea84, 32'hbf6fcc80} /* (16, 7, 21) {real, imag} */,
  {32'hc0ca9e7d, 32'hc0aa97b4} /* (16, 7, 20) {real, imag} */,
  {32'hc028b348, 32'hc05b1798} /* (16, 7, 19) {real, imag} */,
  {32'h3eb4af50, 32'h3f8c9f6e} /* (16, 7, 18) {real, imag} */,
  {32'hc00b5057, 32'hc0930d6d} /* (16, 7, 17) {real, imag} */,
  {32'hc083d98f, 32'h40a7be04} /* (16, 7, 16) {real, imag} */,
  {32'h3f6dbc74, 32'hc03dc972} /* (16, 7, 15) {real, imag} */,
  {32'h4086a61f, 32'h40a90c56} /* (16, 7, 14) {real, imag} */,
  {32'hc0c5f088, 32'h40905af8} /* (16, 7, 13) {real, imag} */,
  {32'hbf37f7b8, 32'h4123d956} /* (16, 7, 12) {real, imag} */,
  {32'h402f9840, 32'h3d5a5400} /* (16, 7, 11) {real, imag} */,
  {32'hc0719784, 32'hc09a4ee6} /* (16, 7, 10) {real, imag} */,
  {32'hbfe9a2ec, 32'hc1a1a7a8} /* (16, 7, 9) {real, imag} */,
  {32'h408294bc, 32'hc0e39cde} /* (16, 7, 8) {real, imag} */,
  {32'hc1cab4ab, 32'hc0007078} /* (16, 7, 7) {real, imag} */,
  {32'h3fafbbd4, 32'h40d28115} /* (16, 7, 6) {real, imag} */,
  {32'hc137aaaa, 32'h420a4b89} /* (16, 7, 5) {real, imag} */,
  {32'hc1d51300, 32'h4193f527} /* (16, 7, 4) {real, imag} */,
  {32'hc07b29f8, 32'h41e2bf52} /* (16, 7, 3) {real, imag} */,
  {32'hc1874915, 32'h3fc7af28} /* (16, 7, 2) {real, imag} */,
  {32'h4190e8de, 32'hbed15e80} /* (16, 7, 1) {real, imag} */,
  {32'h40aeb359, 32'h41e530a9} /* (16, 7, 0) {real, imag} */,
  {32'hc19a43f8, 32'hc130680a} /* (16, 6, 31) {real, imag} */,
  {32'h4149b8a9, 32'h41b74eaa} /* (16, 6, 30) {real, imag} */,
  {32'hc155fa1c, 32'h42070b2e} /* (16, 6, 29) {real, imag} */,
  {32'hc1e9e7ac, 32'h3f48ba7c} /* (16, 6, 28) {real, imag} */,
  {32'hc1a2792b, 32'h41bc6196} /* (16, 6, 27) {real, imag} */,
  {32'hc1890a94, 32'hbf2064a0} /* (16, 6, 26) {real, imag} */,
  {32'hc1910515, 32'hc1956568} /* (16, 6, 25) {real, imag} */,
  {32'h413d5044, 32'h4028a91c} /* (16, 6, 24) {real, imag} */,
  {32'hc1290c3b, 32'hbfd8d0b4} /* (16, 6, 23) {real, imag} */,
  {32'h4081a052, 32'hc1719a29} /* (16, 6, 22) {real, imag} */,
  {32'h40dce1d6, 32'hc0ae823f} /* (16, 6, 21) {real, imag} */,
  {32'h414ffdf5, 32'h40d731ee} /* (16, 6, 20) {real, imag} */,
  {32'h410f307c, 32'hc10f5b50} /* (16, 6, 19) {real, imag} */,
  {32'hc061f836, 32'hc0dade9e} /* (16, 6, 18) {real, imag} */,
  {32'hc04571e4, 32'hc11146f4} /* (16, 6, 17) {real, imag} */,
  {32'hbefef700, 32'hbd2a9400} /* (16, 6, 16) {real, imag} */,
  {32'h40d85626, 32'h409285f5} /* (16, 6, 15) {real, imag} */,
  {32'h402276aa, 32'h3ffbe23a} /* (16, 6, 14) {real, imag} */,
  {32'hbe763660, 32'hc027c72e} /* (16, 6, 13) {real, imag} */,
  {32'h40b60816, 32'hbf94ced8} /* (16, 6, 12) {real, imag} */,
  {32'h41440a4d, 32'hc1a306eb} /* (16, 6, 11) {real, imag} */,
  {32'hc156c5bd, 32'h3f51ab10} /* (16, 6, 10) {real, imag} */,
  {32'h4093323c, 32'hc14f79c2} /* (16, 6, 9) {real, imag} */,
  {32'h41cd0336, 32'hbfe20658} /* (16, 6, 8) {real, imag} */,
  {32'hc12bb1f6, 32'h418df19c} /* (16, 6, 7) {real, imag} */,
  {32'h40d94506, 32'hc14346f6} /* (16, 6, 6) {real, imag} */,
  {32'h41ef02f9, 32'h4106009a} /* (16, 6, 5) {real, imag} */,
  {32'h419989e8, 32'h3f537240} /* (16, 6, 4) {real, imag} */,
  {32'hc0208aaa, 32'h41c0cc97} /* (16, 6, 3) {real, imag} */,
  {32'hc15814ff, 32'hc14fdb9c} /* (16, 6, 2) {real, imag} */,
  {32'hc1f5e7f4, 32'hc2391a02} /* (16, 6, 1) {real, imag} */,
  {32'h402655c0, 32'hc1f219f6} /* (16, 6, 0) {real, imag} */,
  {32'hc0eeb7e8, 32'hc18ef3be} /* (16, 5, 31) {real, imag} */,
  {32'hc0d39eb2, 32'h4239d613} /* (16, 5, 30) {real, imag} */,
  {32'h4200105e, 32'hbe7f3a00} /* (16, 5, 29) {real, imag} */,
  {32'h411f1ded, 32'h419a05dc} /* (16, 5, 28) {real, imag} */,
  {32'hc138e10d, 32'h419dfee2} /* (16, 5, 27) {real, imag} */,
  {32'hc1462dd1, 32'h4185ac53} /* (16, 5, 26) {real, imag} */,
  {32'hbebcbec8, 32'h3ff865d4} /* (16, 5, 25) {real, imag} */,
  {32'h4150d697, 32'h407f8b50} /* (16, 5, 24) {real, imag} */,
  {32'h3eed7440, 32'hc1031fab} /* (16, 5, 23) {real, imag} */,
  {32'h40bac756, 32'h3efa1010} /* (16, 5, 22) {real, imag} */,
  {32'h40a6d4a6, 32'hc1515756} /* (16, 5, 21) {real, imag} */,
  {32'hc1684f8d, 32'hbfde4814} /* (16, 5, 20) {real, imag} */,
  {32'h3ff4663c, 32'hc1578600} /* (16, 5, 19) {real, imag} */,
  {32'hc0feb4ca, 32'hbfb93d18} /* (16, 5, 18) {real, imag} */,
  {32'hc095f913, 32'h3f0c08c8} /* (16, 5, 17) {real, imag} */,
  {32'h3ed29620, 32'hc0729ac4} /* (16, 5, 16) {real, imag} */,
  {32'h400d35d6, 32'h4131c8ce} /* (16, 5, 15) {real, imag} */,
  {32'h409605ca, 32'h407eaf4c} /* (16, 5, 14) {real, imag} */,
  {32'hbf6de518, 32'h4032a2d8} /* (16, 5, 13) {real, imag} */,
  {32'hc0b779ee, 32'hc05e23da} /* (16, 5, 12) {real, imag} */,
  {32'h41797219, 32'h40ae4458} /* (16, 5, 11) {real, imag} */,
  {32'h409118d2, 32'h3e555ee0} /* (16, 5, 10) {real, imag} */,
  {32'hc11c47b4, 32'h413bded9} /* (16, 5, 9) {real, imag} */,
  {32'h41aa9c18, 32'hc0d6eab8} /* (16, 5, 8) {real, imag} */,
  {32'hc0e31610, 32'h4112925c} /* (16, 5, 7) {real, imag} */,
  {32'hc012e0f4, 32'h41334fe6} /* (16, 5, 6) {real, imag} */,
  {32'hc08128ae, 32'h4221a0d1} /* (16, 5, 5) {real, imag} */,
  {32'hc0be0072, 32'hc1fb08d0} /* (16, 5, 4) {real, imag} */,
  {32'h419d18d9, 32'h42047708} /* (16, 5, 3) {real, imag} */,
  {32'hc1f11b9c, 32'h40de47f8} /* (16, 5, 2) {real, imag} */,
  {32'hc15f6fec, 32'hc184061a} /* (16, 5, 1) {real, imag} */,
  {32'hc0bbf20e, 32'hc200cc8b} /* (16, 5, 0) {real, imag} */,
  {32'h41be198c, 32'hc26c7076} /* (16, 4, 31) {real, imag} */,
  {32'hc1968cb9, 32'h4202c5cc} /* (16, 4, 30) {real, imag} */,
  {32'hbf8143f8, 32'h40f0a443} /* (16, 4, 29) {real, imag} */,
  {32'hc233be43, 32'h40cf39f0} /* (16, 4, 28) {real, imag} */,
  {32'hc116e611, 32'h420974e4} /* (16, 4, 27) {real, imag} */,
  {32'h41c26742, 32'hbfe0bb48} /* (16, 4, 26) {real, imag} */,
  {32'h41c98960, 32'hc1915324} /* (16, 4, 25) {real, imag} */,
  {32'hc187d90e, 32'h4087bc2f} /* (16, 4, 24) {real, imag} */,
  {32'h41d9fa1b, 32'hc024c830} /* (16, 4, 23) {real, imag} */,
  {32'h408eb392, 32'h411861b6} /* (16, 4, 22) {real, imag} */,
  {32'h40b7bed4, 32'h40cee74a} /* (16, 4, 21) {real, imag} */,
  {32'h4040833c, 32'hc18012ae} /* (16, 4, 20) {real, imag} */,
  {32'hc025f902, 32'hc0a44511} /* (16, 4, 19) {real, imag} */,
  {32'hc132477e, 32'hc007a876} /* (16, 4, 18) {real, imag} */,
  {32'hc180dc7e, 32'h4188629e} /* (16, 4, 17) {real, imag} */,
  {32'hbf46eb00, 32'hc0f81ffa} /* (16, 4, 16) {real, imag} */,
  {32'hc116cc1f, 32'hc0c0d12e} /* (16, 4, 15) {real, imag} */,
  {32'h41099216, 32'hc03a0bba} /* (16, 4, 14) {real, imag} */,
  {32'hc0b6acbd, 32'h41159970} /* (16, 4, 13) {real, imag} */,
  {32'h4110d217, 32'hc0faf578} /* (16, 4, 12) {real, imag} */,
  {32'hc145e5ea, 32'hc189f10a} /* (16, 4, 11) {real, imag} */,
  {32'h41494f1b, 32'h42079f4a} /* (16, 4, 10) {real, imag} */,
  {32'h41349c22, 32'h418a3fb6} /* (16, 4, 9) {real, imag} */,
  {32'h41319e46, 32'hc1658468} /* (16, 4, 8) {real, imag} */,
  {32'hc1aa64c6, 32'h41408190} /* (16, 4, 7) {real, imag} */,
  {32'hc1e59722, 32'h4161c07a} /* (16, 4, 6) {real, imag} */,
  {32'h413af707, 32'h41bf0c20} /* (16, 4, 5) {real, imag} */,
  {32'h418e8ffa, 32'hc24ce00a} /* (16, 4, 4) {real, imag} */,
  {32'h41d33394, 32'hc0c76559} /* (16, 4, 3) {real, imag} */,
  {32'hc0cf7d14, 32'h425388a0} /* (16, 4, 2) {real, imag} */,
  {32'h3e4d8540, 32'hc194e2dc} /* (16, 4, 1) {real, imag} */,
  {32'hc1b19894, 32'hc18eb0be} /* (16, 4, 0) {real, imag} */,
  {32'hc2581394, 32'h4202e067} /* (16, 3, 31) {real, imag} */,
  {32'hc1589dbc, 32'hc1892a23} /* (16, 3, 30) {real, imag} */,
  {32'hc21d7df9, 32'h4250da55} /* (16, 3, 29) {real, imag} */,
  {32'h42176de8, 32'h415cc37a} /* (16, 3, 28) {real, imag} */,
  {32'hc0cff16c, 32'hc1b558e7} /* (16, 3, 27) {real, imag} */,
  {32'h419bf740, 32'hc1619d55} /* (16, 3, 26) {real, imag} */,
  {32'hc1d9fba0, 32'hc16df2eb} /* (16, 3, 25) {real, imag} */,
  {32'hc106fcc8, 32'hc1b72940} /* (16, 3, 24) {real, imag} */,
  {32'hc0746b82, 32'hc119f790} /* (16, 3, 23) {real, imag} */,
  {32'h412ecc73, 32'h3f118b72} /* (16, 3, 22) {real, imag} */,
  {32'hc154c910, 32'h40a1e81c} /* (16, 3, 21) {real, imag} */,
  {32'hc0da5114, 32'h40d1bc6d} /* (16, 3, 20) {real, imag} */,
  {32'h40d30bc7, 32'hc063ea00} /* (16, 3, 19) {real, imag} */,
  {32'hc154be4f, 32'hbfcaae34} /* (16, 3, 18) {real, imag} */,
  {32'h41321a50, 32'hc0d08b10} /* (16, 3, 17) {real, imag} */,
  {32'hbf4ca5f0, 32'h4061df8c} /* (16, 3, 16) {real, imag} */,
  {32'hc0b69a08, 32'h40f3b438} /* (16, 3, 15) {real, imag} */,
  {32'h40a834d6, 32'hc141f2f8} /* (16, 3, 14) {real, imag} */,
  {32'hc08d6c87, 32'hc1aac82e} /* (16, 3, 13) {real, imag} */,
  {32'h3f7a2560, 32'hc0f08c9f} /* (16, 3, 12) {real, imag} */,
  {32'h41b56ca2, 32'h41d3e23f} /* (16, 3, 11) {real, imag} */,
  {32'h417e4585, 32'hc00a47fc} /* (16, 3, 10) {real, imag} */,
  {32'hc1603ac0, 32'hc170e0a2} /* (16, 3, 9) {real, imag} */,
  {32'h41604a40, 32'hc060924c} /* (16, 3, 8) {real, imag} */,
  {32'h407f88c0, 32'h420a868f} /* (16, 3, 7) {real, imag} */,
  {32'hc106b22f, 32'hc1492f6b} /* (16, 3, 6) {real, imag} */,
  {32'h41b90a87, 32'h41499512} /* (16, 3, 5) {real, imag} */,
  {32'hc097e75c, 32'hc14d3aac} /* (16, 3, 4) {real, imag} */,
  {32'hc1ef874e, 32'h40dd7030} /* (16, 3, 3) {real, imag} */,
  {32'h40d364d4, 32'hc2265f0c} /* (16, 3, 2) {real, imag} */,
  {32'hc24ccecc, 32'h42044ff5} /* (16, 3, 1) {real, imag} */,
  {32'hc1196ac5, 32'hbfa939d0} /* (16, 3, 0) {real, imag} */,
  {32'h3f881170, 32'hc138adc7} /* (16, 2, 31) {real, imag} */,
  {32'h41d43918, 32'h411c49a7} /* (16, 2, 30) {real, imag} */,
  {32'hc190ec47, 32'hc19d296c} /* (16, 2, 29) {real, imag} */,
  {32'h41847134, 32'hc110643c} /* (16, 2, 28) {real, imag} */,
  {32'hc1b03a63, 32'hbd3a31c0} /* (16, 2, 27) {real, imag} */,
  {32'h40d76aae, 32'h412566fe} /* (16, 2, 26) {real, imag} */,
  {32'hbdae7e40, 32'hc191d5dc} /* (16, 2, 25) {real, imag} */,
  {32'h4103f8ff, 32'h41a45254} /* (16, 2, 24) {real, imag} */,
  {32'h41b1d8cc, 32'hc146d713} /* (16, 2, 23) {real, imag} */,
  {32'hc2138934, 32'h411c454e} /* (16, 2, 22) {real, imag} */,
  {32'h40cdfff8, 32'h402502cd} /* (16, 2, 21) {real, imag} */,
  {32'hbfcee6d1, 32'h404629ea} /* (16, 2, 20) {real, imag} */,
  {32'hc1a66c34, 32'h417c1ec4} /* (16, 2, 19) {real, imag} */,
  {32'hbe8ea8b0, 32'hc08e3536} /* (16, 2, 18) {real, imag} */,
  {32'hc00ceee8, 32'h4154e116} /* (16, 2, 17) {real, imag} */,
  {32'h3f049302, 32'hbfdd621c} /* (16, 2, 16) {real, imag} */,
  {32'hc0f100b4, 32'hc0a7b904} /* (16, 2, 15) {real, imag} */,
  {32'hc0735166, 32'hc06a4954} /* (16, 2, 14) {real, imag} */,
  {32'hc108a1cd, 32'hbffadaf0} /* (16, 2, 13) {real, imag} */,
  {32'hbf1548b2, 32'hc1224e64} /* (16, 2, 12) {real, imag} */,
  {32'h41cb1142, 32'h41280bc1} /* (16, 2, 11) {real, imag} */,
  {32'h41c08963, 32'h4061e906} /* (16, 2, 10) {real, imag} */,
  {32'hbf078470, 32'h406614a4} /* (16, 2, 9) {real, imag} */,
  {32'hc17075f9, 32'h41916e24} /* (16, 2, 8) {real, imag} */,
  {32'hc0e68ab9, 32'h3f9fe8e0} /* (16, 2, 7) {real, imag} */,
  {32'h4112b07d, 32'h42003ec2} /* (16, 2, 6) {real, imag} */,
  {32'h420a7dcd, 32'hc0c3b62c} /* (16, 2, 5) {real, imag} */,
  {32'hc1452a54, 32'h42128f21} /* (16, 2, 4) {real, imag} */,
  {32'hc194d7ef, 32'hc1b97954} /* (16, 2, 3) {real, imag} */,
  {32'hc170449c, 32'h41a0012e} /* (16, 2, 2) {real, imag} */,
  {32'hc2389c54, 32'h41882350} /* (16, 2, 1) {real, imag} */,
  {32'h40058fda, 32'h4104b9ae} /* (16, 2, 0) {real, imag} */,
  {32'h41a20dee, 32'h4216608e} /* (16, 1, 31) {real, imag} */,
  {32'hc18ff5f2, 32'h422f777d} /* (16, 1, 30) {real, imag} */,
  {32'h41388991, 32'h42251e74} /* (16, 1, 29) {real, imag} */,
  {32'h3fff6990, 32'hc0059620} /* (16, 1, 28) {real, imag} */,
  {32'hc04dc5c4, 32'hc2075c54} /* (16, 1, 27) {real, imag} */,
  {32'h4153e140, 32'h41ae2aa6} /* (16, 1, 26) {real, imag} */,
  {32'hc034217c, 32'hbfe8b6ae} /* (16, 1, 25) {real, imag} */,
  {32'hc068d040, 32'hc1910d2a} /* (16, 1, 24) {real, imag} */,
  {32'hc12838bc, 32'hc076b798} /* (16, 1, 23) {real, imag} */,
  {32'hc14bdbad, 32'h41054671} /* (16, 1, 22) {real, imag} */,
  {32'hc11323f1, 32'h4024b0a0} /* (16, 1, 21) {real, imag} */,
  {32'hc1b61bb7, 32'hbf8a9624} /* (16, 1, 20) {real, imag} */,
  {32'h40e75994, 32'hc119f870} /* (16, 1, 19) {real, imag} */,
  {32'h40920a31, 32'h40862f80} /* (16, 1, 18) {real, imag} */,
  {32'hbf350610, 32'hbe6169c0} /* (16, 1, 17) {real, imag} */,
  {32'h3f841960, 32'h41141b32} /* (16, 1, 16) {real, imag} */,
  {32'h3f12c010, 32'h3d5cb500} /* (16, 1, 15) {real, imag} */,
  {32'hbec1c350, 32'h4032d4f0} /* (16, 1, 14) {real, imag} */,
  {32'h40827518, 32'h416cd054} /* (16, 1, 13) {real, imag} */,
  {32'h40017dc8, 32'hc1132bb4} /* (16, 1, 12) {real, imag} */,
  {32'hc0aa44d2, 32'hc1b6e5ea} /* (16, 1, 11) {real, imag} */,
  {32'hc1c6d3ca, 32'h40fb726a} /* (16, 1, 10) {real, imag} */,
  {32'h418973c6, 32'hc1b6c708} /* (16, 1, 9) {real, imag} */,
  {32'h3ff30c20, 32'hbfc4bb40} /* (16, 1, 8) {real, imag} */,
  {32'hc0c9ab50, 32'hc0fc6930} /* (16, 1, 7) {real, imag} */,
  {32'h40c3f5c4, 32'h411e1a46} /* (16, 1, 6) {real, imag} */,
  {32'h4206b842, 32'hc11b7764} /* (16, 1, 5) {real, imag} */,
  {32'hc23ffe78, 32'hc1a226b0} /* (16, 1, 4) {real, imag} */,
  {32'hc1434df5, 32'hc201f0d8} /* (16, 1, 3) {real, imag} */,
  {32'hc1c34dae, 32'h4219aaa7} /* (16, 1, 2) {real, imag} */,
  {32'hc0c55bb2, 32'hbd71a200} /* (16, 1, 1) {real, imag} */,
  {32'h41f65d90, 32'hc120a604} /* (16, 1, 0) {real, imag} */,
  {32'h41978b04, 32'h40ed2340} /* (16, 0, 31) {real, imag} */,
  {32'hbfda01b8, 32'hc19ae176} /* (16, 0, 30) {real, imag} */,
  {32'h41caac5c, 32'h406c1a1e} /* (16, 0, 29) {real, imag} */,
  {32'hc1334d37, 32'h4147d8a8} /* (16, 0, 28) {real, imag} */,
  {32'hc212a8d0, 32'hc0d6b807} /* (16, 0, 27) {real, imag} */,
  {32'h40893f52, 32'hc183ba14} /* (16, 0, 26) {real, imag} */,
  {32'hc1694cf2, 32'hc1e11a1c} /* (16, 0, 25) {real, imag} */,
  {32'h40b81aa1, 32'hc144dde6} /* (16, 0, 24) {real, imag} */,
  {32'hc224ba0e, 32'hc164e334} /* (16, 0, 23) {real, imag} */,
  {32'hc0e5d43c, 32'hc1aa328c} /* (16, 0, 22) {real, imag} */,
  {32'hc021e610, 32'h4117c560} /* (16, 0, 21) {real, imag} */,
  {32'h4091d01e, 32'hc111dd64} /* (16, 0, 20) {real, imag} */,
  {32'h3f793150, 32'h40e4d251} /* (16, 0, 19) {real, imag} */,
  {32'hc134c0bf, 32'hc1502ebb} /* (16, 0, 18) {real, imag} */,
  {32'h40a55ac0, 32'h402fa2e4} /* (16, 0, 17) {real, imag} */,
  {32'hc0f73ad9, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h40a55ac0, 32'hc02fa2e4} /* (16, 0, 15) {real, imag} */,
  {32'hc134c0bf, 32'h41502ebb} /* (16, 0, 14) {real, imag} */,
  {32'h3f793150, 32'hc0e4d251} /* (16, 0, 13) {real, imag} */,
  {32'h4091d01e, 32'h4111dd64} /* (16, 0, 12) {real, imag} */,
  {32'hc021e610, 32'hc117c560} /* (16, 0, 11) {real, imag} */,
  {32'hc0e5d43c, 32'h41aa328c} /* (16, 0, 10) {real, imag} */,
  {32'hc224ba0e, 32'h4164e334} /* (16, 0, 9) {real, imag} */,
  {32'h40b81aa1, 32'h4144dde6} /* (16, 0, 8) {real, imag} */,
  {32'hc1694cf2, 32'h41e11a1c} /* (16, 0, 7) {real, imag} */,
  {32'h40893f52, 32'h4183ba14} /* (16, 0, 6) {real, imag} */,
  {32'hc212a8d0, 32'h40d6b807} /* (16, 0, 5) {real, imag} */,
  {32'hc1334d37, 32'hc147d8a8} /* (16, 0, 4) {real, imag} */,
  {32'h41caac5c, 32'hc06c1a1e} /* (16, 0, 3) {real, imag} */,
  {32'hbfda01b8, 32'h419ae176} /* (16, 0, 2) {real, imag} */,
  {32'h41978b04, 32'hc0ed2340} /* (16, 0, 1) {real, imag} */,
  {32'hbe3e2a20, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h41f15082, 32'hc1d1e678} /* (15, 31, 31) {real, imag} */,
  {32'hc25115ea, 32'h41c182a8} /* (15, 31, 30) {real, imag} */,
  {32'hc1ef08c3, 32'h42c19a1c} /* (15, 31, 29) {real, imag} */,
  {32'h418f4fb6, 32'h41b7cdcd} /* (15, 31, 28) {real, imag} */,
  {32'hc2815ef1, 32'h4215a27c} /* (15, 31, 27) {real, imag} */,
  {32'hc06d6eba, 32'h42028b75} /* (15, 31, 26) {real, imag} */,
  {32'h418d3c54, 32'hc13afc9a} /* (15, 31, 25) {real, imag} */,
  {32'hc1896dab, 32'hc0a59ec6} /* (15, 31, 24) {real, imag} */,
  {32'hc13c6114, 32'h41b9bbf8} /* (15, 31, 23) {real, imag} */,
  {32'h4153ec4e, 32'h41b8bcac} /* (15, 31, 22) {real, imag} */,
  {32'hc00d4a5a, 32'hc18002e3} /* (15, 31, 21) {real, imag} */,
  {32'h41054962, 32'hc10c711e} /* (15, 31, 20) {real, imag} */,
  {32'hc060ea3a, 32'h4141808e} /* (15, 31, 19) {real, imag} */,
  {32'hc10803d5, 32'hc0b9f01e} /* (15, 31, 18) {real, imag} */,
  {32'hc0be9474, 32'h4113db3d} /* (15, 31, 17) {real, imag} */,
  {32'h3e5a77c0, 32'h3e7cd400} /* (15, 31, 16) {real, imag} */,
  {32'h4150377a, 32'h415a14d5} /* (15, 31, 15) {real, imag} */,
  {32'hc0a2c9b2, 32'hbfb6d6f8} /* (15, 31, 14) {real, imag} */,
  {32'h4003b896, 32'h3fb63f30} /* (15, 31, 13) {real, imag} */,
  {32'h41f9f917, 32'h3fd3f31c} /* (15, 31, 12) {real, imag} */,
  {32'h416d634e, 32'hc0837b04} /* (15, 31, 11) {real, imag} */,
  {32'h3fc709c4, 32'h401cabdc} /* (15, 31, 10) {real, imag} */,
  {32'h416d570c, 32'hc1f85790} /* (15, 31, 9) {real, imag} */,
  {32'hc0462312, 32'hc2107454} /* (15, 31, 8) {real, imag} */,
  {32'h4230dab0, 32'h42102416} /* (15, 31, 7) {real, imag} */,
  {32'hc125a578, 32'h423f0837} /* (15, 31, 6) {real, imag} */,
  {32'h41caeadc, 32'hc21baf10} /* (15, 31, 5) {real, imag} */,
  {32'h3f8a1bc8, 32'h41f33fc7} /* (15, 31, 4) {real, imag} */,
  {32'h3ed111c0, 32'h41ab04a8} /* (15, 31, 3) {real, imag} */,
  {32'hc134d626, 32'hc26c5508} /* (15, 31, 2) {real, imag} */,
  {32'h42723857, 32'h4235f722} /* (15, 31, 1) {real, imag} */,
  {32'h3f65c290, 32'hc1bf2a16} /* (15, 31, 0) {real, imag} */,
  {32'h3fe88018, 32'h41ebf940} /* (15, 30, 31) {real, imag} */,
  {32'h428e8fb8, 32'hc2230bb9} /* (15, 30, 30) {real, imag} */,
  {32'hc1a53470, 32'hc18c4450} /* (15, 30, 29) {real, imag} */,
  {32'h41302ef5, 32'hc1e52825} /* (15, 30, 28) {real, imag} */,
  {32'hc1f8f4cf, 32'hc1353f1b} /* (15, 30, 27) {real, imag} */,
  {32'h412a1b96, 32'hc174e124} /* (15, 30, 26) {real, imag} */,
  {32'hc1bdb84c, 32'h41509ca4} /* (15, 30, 25) {real, imag} */,
  {32'h41aa52d0, 32'hc0750cee} /* (15, 30, 24) {real, imag} */,
  {32'hc11493da, 32'h419c270c} /* (15, 30, 23) {real, imag} */,
  {32'h41857789, 32'h40eb7dae} /* (15, 30, 22) {real, imag} */,
  {32'h410b82ae, 32'hc11dc089} /* (15, 30, 21) {real, imag} */,
  {32'h40cce708, 32'h40cc4859} /* (15, 30, 20) {real, imag} */,
  {32'hc086e540, 32'hbfe59e40} /* (15, 30, 19) {real, imag} */,
  {32'hc13a3ac5, 32'h411b7860} /* (15, 30, 18) {real, imag} */,
  {32'h40e8905e, 32'hc0cfbefc} /* (15, 30, 17) {real, imag} */,
  {32'h41169d51, 32'hc0ca0776} /* (15, 30, 16) {real, imag} */,
  {32'hc0ae4576, 32'h413b528e} /* (15, 30, 15) {real, imag} */,
  {32'h3e8bf0a0, 32'hc0b230ec} /* (15, 30, 14) {real, imag} */,
  {32'h3f189a80, 32'h40ba36e4} /* (15, 30, 13) {real, imag} */,
  {32'h40ce90b4, 32'h3f2997d8} /* (15, 30, 12) {real, imag} */,
  {32'hc1e71907, 32'h4082fab0} /* (15, 30, 11) {real, imag} */,
  {32'hc0301a08, 32'hc1af8946} /* (15, 30, 10) {real, imag} */,
  {32'h3ee10530, 32'hc21fa7d4} /* (15, 30, 9) {real, imag} */,
  {32'h41e327dc, 32'hc14f6ba2} /* (15, 30, 8) {real, imag} */,
  {32'hc1633cdc, 32'h3fd9b9e0} /* (15, 30, 7) {real, imag} */,
  {32'hc07acf4a, 32'hc17a7416} /* (15, 30, 6) {real, imag} */,
  {32'hc1ec83e9, 32'h4056b57f} /* (15, 30, 5) {real, imag} */,
  {32'hc14732ad, 32'hc161772e} /* (15, 30, 4) {real, imag} */,
  {32'h4200e592, 32'hc1eda484} /* (15, 30, 3) {real, imag} */,
  {32'h419d2250, 32'h3f65d740} /* (15, 30, 2) {real, imag} */,
  {32'h3f559cd0, 32'h423c3a38} /* (15, 30, 1) {real, imag} */,
  {32'hc0fcb8d6, 32'h41e986b6} /* (15, 30, 0) {real, imag} */,
  {32'h414fb73a, 32'hc213574a} /* (15, 29, 31) {real, imag} */,
  {32'hc06a3500, 32'h41ddcb62} /* (15, 29, 30) {real, imag} */,
  {32'hc0058df4, 32'hc1f8965e} /* (15, 29, 29) {real, imag} */,
  {32'hc1c1d459, 32'h3f928150} /* (15, 29, 28) {real, imag} */,
  {32'h41f451b2, 32'h40d32723} /* (15, 29, 27) {real, imag} */,
  {32'hc16ec588, 32'hc1ef1c6d} /* (15, 29, 26) {real, imag} */,
  {32'hc182c380, 32'hc1d315e6} /* (15, 29, 25) {real, imag} */,
  {32'h4218ca32, 32'h413cb4be} /* (15, 29, 24) {real, imag} */,
  {32'hc172442c, 32'h41325543} /* (15, 29, 23) {real, imag} */,
  {32'hc17018e6, 32'hc1ca5351} /* (15, 29, 22) {real, imag} */,
  {32'h41851560, 32'h40c9d959} /* (15, 29, 21) {real, imag} */,
  {32'hbfdb131d, 32'h419cb7fb} /* (15, 29, 20) {real, imag} */,
  {32'h4135d999, 32'h400908b8} /* (15, 29, 19) {real, imag} */,
  {32'hc14ef9a8, 32'hc0cf2973} /* (15, 29, 18) {real, imag} */,
  {32'hbf21a3e8, 32'h40ce5206} /* (15, 29, 17) {real, imag} */,
  {32'h41315400, 32'h403162ba} /* (15, 29, 16) {real, imag} */,
  {32'h40eb3a0d, 32'hc017203c} /* (15, 29, 15) {real, imag} */,
  {32'hc13316f4, 32'hc11843d6} /* (15, 29, 14) {real, imag} */,
  {32'h40e3e772, 32'h3ebb8840} /* (15, 29, 13) {real, imag} */,
  {32'hc094d9b5, 32'hc16ea776} /* (15, 29, 12) {real, imag} */,
  {32'h4182382c, 32'hc1924dbc} /* (15, 29, 11) {real, imag} */,
  {32'hc1b5d915, 32'hc0b4b1c0} /* (15, 29, 10) {real, imag} */,
  {32'hc1c825e6, 32'h416fa6bf} /* (15, 29, 9) {real, imag} */,
  {32'h411911a0, 32'hc0ca91a1} /* (15, 29, 8) {real, imag} */,
  {32'hc13c56e0, 32'h416cb6a7} /* (15, 29, 7) {real, imag} */,
  {32'h41539410, 32'hbfb26e60} /* (15, 29, 6) {real, imag} */,
  {32'hc1087c4b, 32'hc1576652} /* (15, 29, 5) {real, imag} */,
  {32'hc186645f, 32'h41e66ccf} /* (15, 29, 4) {real, imag} */,
  {32'hc1321609, 32'h42190269} /* (15, 29, 3) {real, imag} */,
  {32'hc1a9840e, 32'h420466ff} /* (15, 29, 2) {real, imag} */,
  {32'h416ba6ee, 32'h40c80124} /* (15, 29, 1) {real, imag} */,
  {32'h4248183a, 32'hc18831d5} /* (15, 29, 0) {real, imag} */,
  {32'hc1ce6510, 32'h416cc1e1} /* (15, 28, 31) {real, imag} */,
  {32'h421f4e4a, 32'hc1a26ce8} /* (15, 28, 30) {real, imag} */,
  {32'hc2291603, 32'hc1234cfd} /* (15, 28, 29) {real, imag} */,
  {32'hbf0a2558, 32'h4236a5e9} /* (15, 28, 28) {real, imag} */,
  {32'hc280ba21, 32'h4018ce0c} /* (15, 28, 27) {real, imag} */,
  {32'h410deec1, 32'h416a2ba6} /* (15, 28, 26) {real, imag} */,
  {32'hc0b92fe6, 32'hc21f4296} /* (15, 28, 25) {real, imag} */,
  {32'hc0dca96e, 32'h41832228} /* (15, 28, 24) {real, imag} */,
  {32'h400f52f0, 32'hc15e0e10} /* (15, 28, 23) {real, imag} */,
  {32'h4102c308, 32'h3fd638d8} /* (15, 28, 22) {real, imag} */,
  {32'h40fa124a, 32'hc152ab4b} /* (15, 28, 21) {real, imag} */,
  {32'h4139c187, 32'hbe6077c0} /* (15, 28, 20) {real, imag} */,
  {32'h413ca839, 32'h41316825} /* (15, 28, 19) {real, imag} */,
  {32'hc08d35d6, 32'h40fa20cb} /* (15, 28, 18) {real, imag} */,
  {32'hbf949460, 32'hc10c3bcb} /* (15, 28, 17) {real, imag} */,
  {32'hbf23ece0, 32'h3ffe8ef8} /* (15, 28, 16) {real, imag} */,
  {32'h406994c8, 32'h409b8df2} /* (15, 28, 15) {real, imag} */,
  {32'h41192f09, 32'h3e3a04e0} /* (15, 28, 14) {real, imag} */,
  {32'hbfc00978, 32'h4029d6dc} /* (15, 28, 13) {real, imag} */,
  {32'hc0c63cd6, 32'h417aeb99} /* (15, 28, 12) {real, imag} */,
  {32'hc0532b2c, 32'hbf22a910} /* (15, 28, 11) {real, imag} */,
  {32'hc1832c77, 32'hc101f693} /* (15, 28, 10) {real, imag} */,
  {32'h415491c0, 32'hbf614138} /* (15, 28, 9) {real, imag} */,
  {32'h40be8b6e, 32'h419d54d0} /* (15, 28, 8) {real, imag} */,
  {32'h41249d4d, 32'hc2044bc6} /* (15, 28, 7) {real, imag} */,
  {32'h4164dbcb, 32'h4175be52} /* (15, 28, 6) {real, imag} */,
  {32'h413f8428, 32'hc1bc684e} /* (15, 28, 5) {real, imag} */,
  {32'h40ac2d4a, 32'hc231ae41} /* (15, 28, 4) {real, imag} */,
  {32'h4256ff43, 32'h4188c24a} /* (15, 28, 3) {real, imag} */,
  {32'hc1e0f423, 32'h420337fc} /* (15, 28, 2) {real, imag} */,
  {32'h403cb7a4, 32'hc0452c0c} /* (15, 28, 1) {real, imag} */,
  {32'h41a92d35, 32'hc15778cb} /* (15, 28, 0) {real, imag} */,
  {32'hc1feb2c3, 32'h42705746} /* (15, 27, 31) {real, imag} */,
  {32'h424ff69e, 32'hc24ef002} /* (15, 27, 30) {real, imag} */,
  {32'h414fa263, 32'h42235ba2} /* (15, 27, 29) {real, imag} */,
  {32'hc19270e0, 32'hc13ac30b} /* (15, 27, 28) {real, imag} */,
  {32'h418c908d, 32'h41ebe905} /* (15, 27, 27) {real, imag} */,
  {32'hc213c94e, 32'h4213cce2} /* (15, 27, 26) {real, imag} */,
  {32'hc15c527a, 32'hc18752b3} /* (15, 27, 25) {real, imag} */,
  {32'hc11dcb44, 32'h4174889c} /* (15, 27, 24) {real, imag} */,
  {32'h41158b94, 32'h3f0b96b8} /* (15, 27, 23) {real, imag} */,
  {32'h40d711f2, 32'hc173ccc3} /* (15, 27, 22) {real, imag} */,
  {32'hc1b6f817, 32'hc1caa9cd} /* (15, 27, 21) {real, imag} */,
  {32'hc02033ec, 32'h40886550} /* (15, 27, 20) {real, imag} */,
  {32'hc0649a02, 32'hbf51b118} /* (15, 27, 19) {real, imag} */,
  {32'h411cffe9, 32'h40b521ed} /* (15, 27, 18) {real, imag} */,
  {32'h412b979c, 32'h40a2539e} /* (15, 27, 17) {real, imag} */,
  {32'h412c7eb0, 32'h40b996b4} /* (15, 27, 16) {real, imag} */,
  {32'h3facba24, 32'h4096c53e} /* (15, 27, 15) {real, imag} */,
  {32'h3f4d7eb0, 32'h3f82ffb4} /* (15, 27, 14) {real, imag} */,
  {32'h3fd03cfc, 32'hc049d5e6} /* (15, 27, 13) {real, imag} */,
  {32'hc0e78cb2, 32'hc014ace5} /* (15, 27, 12) {real, imag} */,
  {32'hc0c9a21c, 32'h3ffdc470} /* (15, 27, 11) {real, imag} */,
  {32'h412ca3af, 32'h419e6c52} /* (15, 27, 10) {real, imag} */,
  {32'h3e537c00, 32'hc020da42} /* (15, 27, 9) {real, imag} */,
  {32'h41b84f0e, 32'h4154d808} /* (15, 27, 8) {real, imag} */,
  {32'hbff7b2f0, 32'h41fad2c7} /* (15, 27, 7) {real, imag} */,
  {32'h40263700, 32'hc1dc0c69} /* (15, 27, 6) {real, imag} */,
  {32'hc1ca57cf, 32'h3fa89d50} /* (15, 27, 5) {real, imag} */,
  {32'h40d2a460, 32'h41c9e232} /* (15, 27, 4) {real, imag} */,
  {32'h41391925, 32'hc1667326} /* (15, 27, 3) {real, imag} */,
  {32'h41ddf1c4, 32'h41c47225} /* (15, 27, 2) {real, imag} */,
  {32'hbffb1910, 32'hc0ddead0} /* (15, 27, 1) {real, imag} */,
  {32'h4197e192, 32'h41afe501} /* (15, 27, 0) {real, imag} */,
  {32'h3cbd4000, 32'h4138e58a} /* (15, 26, 31) {real, imag} */,
  {32'hc1e19e5c, 32'hc203c978} /* (15, 26, 30) {real, imag} */,
  {32'h41892842, 32'hc06949ac} /* (15, 26, 29) {real, imag} */,
  {32'hc21857ac, 32'h41095f3d} /* (15, 26, 28) {real, imag} */,
  {32'hc1007b5b, 32'h403eba07} /* (15, 26, 27) {real, imag} */,
  {32'h412497eb, 32'hc07fe3d9} /* (15, 26, 26) {real, imag} */,
  {32'hc16b5ec6, 32'hc1c95296} /* (15, 26, 25) {real, imag} */,
  {32'h3fbf8630, 32'hc16ee094} /* (15, 26, 24) {real, imag} */,
  {32'h41a652e7, 32'hc0e33b7e} /* (15, 26, 23) {real, imag} */,
  {32'hc079d3ae, 32'h3f5229a0} /* (15, 26, 22) {real, imag} */,
  {32'h4100d289, 32'hc185d481} /* (15, 26, 21) {real, imag} */,
  {32'hc139e54f, 32'h4106a495} /* (15, 26, 20) {real, imag} */,
  {32'h3f95b870, 32'hbf9946d1} /* (15, 26, 19) {real, imag} */,
  {32'hc13607b4, 32'h413d863e} /* (15, 26, 18) {real, imag} */,
  {32'hbff0cc40, 32'hc0af7fa6} /* (15, 26, 17) {real, imag} */,
  {32'h40691ac8, 32'h40978778} /* (15, 26, 16) {real, imag} */,
  {32'h40819af8, 32'hbfcc16b4} /* (15, 26, 15) {real, imag} */,
  {32'hc0a1328b, 32'h3fa0f4c0} /* (15, 26, 14) {real, imag} */,
  {32'hc16a410c, 32'hbf1ee0ba} /* (15, 26, 13) {real, imag} */,
  {32'hc18f2fc4, 32'hc18cab0a} /* (15, 26, 12) {real, imag} */,
  {32'hbd94b3a0, 32'hbfdcb504} /* (15, 26, 11) {real, imag} */,
  {32'hc15de21e, 32'hc16440a0} /* (15, 26, 10) {real, imag} */,
  {32'h404f8738, 32'h4130d69d} /* (15, 26, 9) {real, imag} */,
  {32'h4170d766, 32'hc1e4b09e} /* (15, 26, 8) {real, imag} */,
  {32'h40befbe3, 32'h40e8cdb2} /* (15, 26, 7) {real, imag} */,
  {32'hc18141ac, 32'hc00dec0f} /* (15, 26, 6) {real, imag} */,
  {32'h4195a11c, 32'hc113f509} /* (15, 26, 5) {real, imag} */,
  {32'h415f84ea, 32'hc0852c1e} /* (15, 26, 4) {real, imag} */,
  {32'h41d485b6, 32'h40ce5636} /* (15, 26, 3) {real, imag} */,
  {32'h40a3ae76, 32'h41968494} /* (15, 26, 2) {real, imag} */,
  {32'hc2854e12, 32'h3fa1e680} /* (15, 26, 1) {real, imag} */,
  {32'hc222fd44, 32'hc20dc417} /* (15, 26, 0) {real, imag} */,
  {32'h40ee10c4, 32'hc0ec5cb6} /* (15, 25, 31) {real, imag} */,
  {32'h40e010db, 32'h41edf526} /* (15, 25, 30) {real, imag} */,
  {32'h41e808b2, 32'h407a69ac} /* (15, 25, 29) {real, imag} */,
  {32'hc0ec344e, 32'h419de8a1} /* (15, 25, 28) {real, imag} */,
  {32'h4080a650, 32'hc10f0c24} /* (15, 25, 27) {real, imag} */,
  {32'hc1651e68, 32'h40fa36be} /* (15, 25, 26) {real, imag} */,
  {32'h41d551a7, 32'hc188df50} /* (15, 25, 25) {real, imag} */,
  {32'h4144b1ce, 32'h4106ca84} /* (15, 25, 24) {real, imag} */,
  {32'hc10b7634, 32'hc1c79fec} /* (15, 25, 23) {real, imag} */,
  {32'hc193326c, 32'hbf448344} /* (15, 25, 22) {real, imag} */,
  {32'hc1428e99, 32'h413663ab} /* (15, 25, 21) {real, imag} */,
  {32'hbfd15f70, 32'hc116c6e5} /* (15, 25, 20) {real, imag} */,
  {32'h41523c0a, 32'hbd5631c0} /* (15, 25, 19) {real, imag} */,
  {32'hc0a63076, 32'h40ce7888} /* (15, 25, 18) {real, imag} */,
  {32'hc10d2f2b, 32'h40e5e04b} /* (15, 25, 17) {real, imag} */,
  {32'hc0e3a21c, 32'h41465780} /* (15, 25, 16) {real, imag} */,
  {32'hc04a6044, 32'hc0489662} /* (15, 25, 15) {real, imag} */,
  {32'hc14d4dad, 32'h40ff02a8} /* (15, 25, 14) {real, imag} */,
  {32'h400ac9a6, 32'hbe519970} /* (15, 25, 13) {real, imag} */,
  {32'hc02e1f80, 32'hc11233ab} /* (15, 25, 12) {real, imag} */,
  {32'h409b2a42, 32'h41a457de} /* (15, 25, 11) {real, imag} */,
  {32'h400b9d94, 32'hc0a20bbc} /* (15, 25, 10) {real, imag} */,
  {32'hc18db6e0, 32'hc067fc48} /* (15, 25, 9) {real, imag} */,
  {32'hc0479a48, 32'h413892d6} /* (15, 25, 8) {real, imag} */,
  {32'hc18214a3, 32'hc08dfecc} /* (15, 25, 7) {real, imag} */,
  {32'hc1a57580, 32'hc0c1ff2a} /* (15, 25, 6) {real, imag} */,
  {32'hc0ea8fb0, 32'h405f65b6} /* (15, 25, 5) {real, imag} */,
  {32'h41b7cec8, 32'hbde30b00} /* (15, 25, 4) {real, imag} */,
  {32'h40f53f48, 32'hc190a26c} /* (15, 25, 3) {real, imag} */,
  {32'h40b69bbf, 32'hc1753024} /* (15, 25, 2) {real, imag} */,
  {32'hc1e1c723, 32'hc1bee3a0} /* (15, 25, 1) {real, imag} */,
  {32'hc23a0930, 32'h415abdb2} /* (15, 25, 0) {real, imag} */,
  {32'hc1850367, 32'hc1f11e8c} /* (15, 24, 31) {real, imag} */,
  {32'h3fac56ac, 32'h4187ffe2} /* (15, 24, 30) {real, imag} */,
  {32'h4192929f, 32'hc14fa0b8} /* (15, 24, 29) {real, imag} */,
  {32'h418bb8da, 32'hc1544d22} /* (15, 24, 28) {real, imag} */,
  {32'hc1a1d312, 32'h41b7bedc} /* (15, 24, 27) {real, imag} */,
  {32'hbf737330, 32'hc16bae22} /* (15, 24, 26) {real, imag} */,
  {32'h4103c7b4, 32'h41a32dc9} /* (15, 24, 25) {real, imag} */,
  {32'hc055714c, 32'hc02f3feb} /* (15, 24, 24) {real, imag} */,
  {32'hc0c9f612, 32'hc093c6a8} /* (15, 24, 23) {real, imag} */,
  {32'h3fd019dc, 32'h4093d4d7} /* (15, 24, 22) {real, imag} */,
  {32'hc08f1ff2, 32'h40946631} /* (15, 24, 21) {real, imag} */,
  {32'h40dfabd0, 32'h406764cc} /* (15, 24, 20) {real, imag} */,
  {32'hbf91dc64, 32'h40614cb6} /* (15, 24, 19) {real, imag} */,
  {32'h40034292, 32'hc0874dba} /* (15, 24, 18) {real, imag} */,
  {32'h3fb2c0e0, 32'h3febd1b8} /* (15, 24, 17) {real, imag} */,
  {32'h407d44c7, 32'h411169f8} /* (15, 24, 16) {real, imag} */,
  {32'hbe581680, 32'h413193a1} /* (15, 24, 15) {real, imag} */,
  {32'hc0d12f27, 32'hc0fa1b6a} /* (15, 24, 14) {real, imag} */,
  {32'h40e4330b, 32'hc1072bd4} /* (15, 24, 13) {real, imag} */,
  {32'h40e1c37c, 32'h40a85efe} /* (15, 24, 12) {real, imag} */,
  {32'h411b2871, 32'h41621c5c} /* (15, 24, 11) {real, imag} */,
  {32'hbf65d548, 32'h41171dc8} /* (15, 24, 10) {real, imag} */,
  {32'h400eb549, 32'hc15a0574} /* (15, 24, 9) {real, imag} */,
  {32'h418ecf5c, 32'hbf7d4184} /* (15, 24, 8) {real, imag} */,
  {32'hc0a9fca2, 32'hbf1a5a20} /* (15, 24, 7) {real, imag} */,
  {32'h40d935a0, 32'hc02701ee} /* (15, 24, 6) {real, imag} */,
  {32'hbf248970, 32'h41d146fa} /* (15, 24, 5) {real, imag} */,
  {32'hc1899a9e, 32'hc21e5f7c} /* (15, 24, 4) {real, imag} */,
  {32'h402d1c58, 32'h409f419d} /* (15, 24, 3) {real, imag} */,
  {32'hc10d9384, 32'hc1d5f112} /* (15, 24, 2) {real, imag} */,
  {32'hc1078620, 32'h41334ce1} /* (15, 24, 1) {real, imag} */,
  {32'h3bb3e200, 32'hc12eaef8} /* (15, 24, 0) {real, imag} */,
  {32'hc19a3d40, 32'h404c7687} /* (15, 23, 31) {real, imag} */,
  {32'h41f53148, 32'h410073dc} /* (15, 23, 30) {real, imag} */,
  {32'hc17879c6, 32'h41d3ee57} /* (15, 23, 29) {real, imag} */,
  {32'hc1e7f52c, 32'hc19429c8} /* (15, 23, 28) {real, imag} */,
  {32'h413b77cd, 32'h4139bd5a} /* (15, 23, 27) {real, imag} */,
  {32'h40a3105e, 32'hc0c422e0} /* (15, 23, 26) {real, imag} */,
  {32'hc0920ac0, 32'h40e2fc5b} /* (15, 23, 25) {real, imag} */,
  {32'h3fae4d7c, 32'hbf3eac00} /* (15, 23, 24) {real, imag} */,
  {32'h3f718da8, 32'hc106abed} /* (15, 23, 23) {real, imag} */,
  {32'hc13f3801, 32'h411aed43} /* (15, 23, 22) {real, imag} */,
  {32'hbfccb9a8, 32'h4077618e} /* (15, 23, 21) {real, imag} */,
  {32'h401d29fb, 32'hc0cbc08e} /* (15, 23, 20) {real, imag} */,
  {32'hbeab4d08, 32'h4012598c} /* (15, 23, 19) {real, imag} */,
  {32'h3f592350, 32'hc056888e} /* (15, 23, 18) {real, imag} */,
  {32'h3fa9327c, 32'hbff1fda0} /* (15, 23, 17) {real, imag} */,
  {32'hc053dc1f, 32'hc02d26d8} /* (15, 23, 16) {real, imag} */,
  {32'hc0812345, 32'h3f576138} /* (15, 23, 15) {real, imag} */,
  {32'hc089d876, 32'h40e69d87} /* (15, 23, 14) {real, imag} */,
  {32'hc0fd02e2, 32'hc1440541} /* (15, 23, 13) {real, imag} */,
  {32'hbf7f1d2c, 32'h40dddfb2} /* (15, 23, 12) {real, imag} */,
  {32'h412c4bfc, 32'h3f075de8} /* (15, 23, 11) {real, imag} */,
  {32'hc0d9c426, 32'hc0eed0a6} /* (15, 23, 10) {real, imag} */,
  {32'h4179d2c2, 32'h41758197} /* (15, 23, 9) {real, imag} */,
  {32'h411cb89a, 32'hc2169eee} /* (15, 23, 8) {real, imag} */,
  {32'h41755be0, 32'hbfcfbf9c} /* (15, 23, 7) {real, imag} */,
  {32'hc0f635de, 32'hc0abb388} /* (15, 23, 6) {real, imag} */,
  {32'h404d3028, 32'h411ea304} /* (15, 23, 5) {real, imag} */,
  {32'hc1879364, 32'h41097645} /* (15, 23, 4) {real, imag} */,
  {32'hc1b465e1, 32'hc1f28b3f} /* (15, 23, 3) {real, imag} */,
  {32'h4073b6c0, 32'h4183ff48} /* (15, 23, 2) {real, imag} */,
  {32'hbfac32c8, 32'h410871dc} /* (15, 23, 1) {real, imag} */,
  {32'hbf8875ce, 32'hc20f0304} /* (15, 23, 0) {real, imag} */,
  {32'hc27968f2, 32'hc1527e41} /* (15, 22, 31) {real, imag} */,
  {32'hc17260f8, 32'h4105bd2e} /* (15, 22, 30) {real, imag} */,
  {32'h406115d3, 32'hc0ac8b88} /* (15, 22, 29) {real, imag} */,
  {32'h41284ee3, 32'hc20221a2} /* (15, 22, 28) {real, imag} */,
  {32'hc1299ea9, 32'h41242fb2} /* (15, 22, 27) {real, imag} */,
  {32'h409acc64, 32'h4143f8b4} /* (15, 22, 26) {real, imag} */,
  {32'hc0d0354b, 32'hc187479f} /* (15, 22, 25) {real, imag} */,
  {32'hc04b815c, 32'hc0e41d20} /* (15, 22, 24) {real, imag} */,
  {32'hc037ea39, 32'h412b4e60} /* (15, 22, 23) {real, imag} */,
  {32'h4114cc8a, 32'h41618b02} /* (15, 22, 22) {real, imag} */,
  {32'hc0e698b8, 32'hbf31dce8} /* (15, 22, 21) {real, imag} */,
  {32'hc095839a, 32'h41180c48} /* (15, 22, 20) {real, imag} */,
  {32'h4108c2a8, 32'hc0182483} /* (15, 22, 19) {real, imag} */,
  {32'h4036726b, 32'hc03d22ba} /* (15, 22, 18) {real, imag} */,
  {32'hc0896c0a, 32'h3e307310} /* (15, 22, 17) {real, imag} */,
  {32'h408801f4, 32'hbfbdcf38} /* (15, 22, 16) {real, imag} */,
  {32'h41013a03, 32'hc0ae2570} /* (15, 22, 15) {real, imag} */,
  {32'h40fe25e6, 32'h40782e62} /* (15, 22, 14) {real, imag} */,
  {32'hc1036764, 32'h40025b69} /* (15, 22, 13) {real, imag} */,
  {32'hc1000867, 32'hbfcfa52e} /* (15, 22, 12) {real, imag} */,
  {32'h40f31388, 32'hbf7c9ff8} /* (15, 22, 11) {real, imag} */,
  {32'h4092cf70, 32'hbfc77370} /* (15, 22, 10) {real, imag} */,
  {32'hc103e431, 32'h416a3a20} /* (15, 22, 9) {real, imag} */,
  {32'hc1663139, 32'h407fbf37} /* (15, 22, 8) {real, imag} */,
  {32'h41206578, 32'h40d7b87c} /* (15, 22, 7) {real, imag} */,
  {32'h3f0f45e4, 32'h402f8bf8} /* (15, 22, 6) {real, imag} */,
  {32'h41b09f30, 32'hc17184d6} /* (15, 22, 5) {real, imag} */,
  {32'h41923445, 32'h414e75b8} /* (15, 22, 4) {real, imag} */,
  {32'h40f81fa2, 32'h402b91d5} /* (15, 22, 3) {real, imag} */,
  {32'h4096c2c8, 32'h41a4ce11} /* (15, 22, 2) {real, imag} */,
  {32'h4022f880, 32'hc175c933} /* (15, 22, 1) {real, imag} */,
  {32'h40987fa0, 32'hc173f3d3} /* (15, 22, 0) {real, imag} */,
  {32'hc1a00e52, 32'hbf79a348} /* (15, 21, 31) {real, imag} */,
  {32'hbe62b460, 32'h4177df70} /* (15, 21, 30) {real, imag} */,
  {32'hc1126ba3, 32'hc0c671a2} /* (15, 21, 29) {real, imag} */,
  {32'h414b1bc6, 32'h41b5e98c} /* (15, 21, 28) {real, imag} */,
  {32'h4185dc3d, 32'hc1baa324} /* (15, 21, 27) {real, imag} */,
  {32'hc0fb3290, 32'h4103530b} /* (15, 21, 26) {real, imag} */,
  {32'hc1222c6a, 32'h4182008d} /* (15, 21, 25) {real, imag} */,
  {32'hc02888a0, 32'h407acdb7} /* (15, 21, 24) {real, imag} */,
  {32'h3e902f98, 32'hc08553fa} /* (15, 21, 23) {real, imag} */,
  {32'hbeaa7ec0, 32'h4085cc78} /* (15, 21, 22) {real, imag} */,
  {32'hc101e31e, 32'h408969be} /* (15, 21, 21) {real, imag} */,
  {32'hbf0d7aec, 32'hc11ba321} /* (15, 21, 20) {real, imag} */,
  {32'h4064524d, 32'h3e672d30} /* (15, 21, 19) {real, imag} */,
  {32'h40a0536e, 32'hc0a1dbd5} /* (15, 21, 18) {real, imag} */,
  {32'h40798ffc, 32'hc0842056} /* (15, 21, 17) {real, imag} */,
  {32'hc0597ddc, 32'hc03fe38c} /* (15, 21, 16) {real, imag} */,
  {32'hc073b1c0, 32'hbf971360} /* (15, 21, 15) {real, imag} */,
  {32'hbf3b5abc, 32'h3f5c2f18} /* (15, 21, 14) {real, imag} */,
  {32'hc0eb0a50, 32'h4056e1c9} /* (15, 21, 13) {real, imag} */,
  {32'h41014a0e, 32'h3ff0c678} /* (15, 21, 12) {real, imag} */,
  {32'hc04be066, 32'hc0eef24e} /* (15, 21, 11) {real, imag} */,
  {32'h410157f4, 32'h3fc8dd2e} /* (15, 21, 10) {real, imag} */,
  {32'hc0d96c32, 32'h41528fcb} /* (15, 21, 9) {real, imag} */,
  {32'hbfaff020, 32'hc0d4cf12} /* (15, 21, 8) {real, imag} */,
  {32'hc0d171b0, 32'h40e5ab17} /* (15, 21, 7) {real, imag} */,
  {32'hc1766694, 32'hc0ea9d76} /* (15, 21, 6) {real, imag} */,
  {32'hc088919f, 32'hc183a56e} /* (15, 21, 5) {real, imag} */,
  {32'h40a66d8c, 32'h4113dba7} /* (15, 21, 4) {real, imag} */,
  {32'h4077802f, 32'hc07ea009} /* (15, 21, 3) {real, imag} */,
  {32'h413ac3b6, 32'hc215962f} /* (15, 21, 2) {real, imag} */,
  {32'h4081dd97, 32'hc10e7dc0} /* (15, 21, 1) {real, imag} */,
  {32'h4092ed8c, 32'h4135d1a9} /* (15, 21, 0) {real, imag} */,
  {32'hc1321773, 32'h413077ff} /* (15, 20, 31) {real, imag} */,
  {32'h41803be3, 32'hc0ff1044} /* (15, 20, 30) {real, imag} */,
  {32'h40b03c37, 32'hc08455d6} /* (15, 20, 29) {real, imag} */,
  {32'h4107ae24, 32'hc15e0e16} /* (15, 20, 28) {real, imag} */,
  {32'hc02a9a58, 32'h40e974e0} /* (15, 20, 27) {real, imag} */,
  {32'hbfa0d1d4, 32'hc08e2848} /* (15, 20, 26) {real, imag} */,
  {32'hc096dbbc, 32'hc12f2e9c} /* (15, 20, 25) {real, imag} */,
  {32'h416ce63d, 32'h413b6a52} /* (15, 20, 24) {real, imag} */,
  {32'h4065ecbf, 32'h4130795a} /* (15, 20, 23) {real, imag} */,
  {32'h40b3d58c, 32'h404ce943} /* (15, 20, 22) {real, imag} */,
  {32'h3fbf423c, 32'hbeb9d054} /* (15, 20, 21) {real, imag} */,
  {32'h3fddf820, 32'h40e71742} /* (15, 20, 20) {real, imag} */,
  {32'hbf851041, 32'hc08b16aa} /* (15, 20, 19) {real, imag} */,
  {32'h40a4d367, 32'hbff56908} /* (15, 20, 18) {real, imag} */,
  {32'h3ff23eb2, 32'hc0a45db5} /* (15, 20, 17) {real, imag} */,
  {32'h405eff31, 32'hc0182e24} /* (15, 20, 16) {real, imag} */,
  {32'h3fec863e, 32'h3f9518fd} /* (15, 20, 15) {real, imag} */,
  {32'h409c568b, 32'h409d8b7d} /* (15, 20, 14) {real, imag} */,
  {32'h405b24e2, 32'h402fc9ca} /* (15, 20, 13) {real, imag} */,
  {32'hc1501716, 32'hc083ce94} /* (15, 20, 12) {real, imag} */,
  {32'h4116b410, 32'h4042034a} /* (15, 20, 11) {real, imag} */,
  {32'h4072b480, 32'h40b03212} /* (15, 20, 10) {real, imag} */,
  {32'hbbb63a00, 32'h40f1f2bf} /* (15, 20, 9) {real, imag} */,
  {32'hc0cf3d06, 32'h3ee9a6c0} /* (15, 20, 8) {real, imag} */,
  {32'hc0e8bce0, 32'h3f3c9638} /* (15, 20, 7) {real, imag} */,
  {32'h40e230f9, 32'h40225045} /* (15, 20, 6) {real, imag} */,
  {32'hc1217ab6, 32'h4139d070} /* (15, 20, 5) {real, imag} */,
  {32'hc10f2d26, 32'hc129463e} /* (15, 20, 4) {real, imag} */,
  {32'hc0dcc8d1, 32'h3ff4a1ab} /* (15, 20, 3) {real, imag} */,
  {32'hc1381674, 32'hc0d1d6e8} /* (15, 20, 2) {real, imag} */,
  {32'hc12f4f97, 32'hc161ed7d} /* (15, 20, 1) {real, imag} */,
  {32'h40a96a6c, 32'h40fa78ba} /* (15, 20, 0) {real, imag} */,
  {32'h415c23de, 32'hc0ebd156} /* (15, 19, 31) {real, imag} */,
  {32'h40aa2494, 32'hc17d310c} /* (15, 19, 30) {real, imag} */,
  {32'hc03040ca, 32'hc1098d4f} /* (15, 19, 29) {real, imag} */,
  {32'hbd8f4ec0, 32'h41213d06} /* (15, 19, 28) {real, imag} */,
  {32'hbfb7b036, 32'h40cc6d40} /* (15, 19, 27) {real, imag} */,
  {32'h4055e3b3, 32'h4186a049} /* (15, 19, 26) {real, imag} */,
  {32'h4091e9d0, 32'hbfbf4295} /* (15, 19, 25) {real, imag} */,
  {32'h4103d429, 32'hc03bfcd0} /* (15, 19, 24) {real, imag} */,
  {32'hc0bc329a, 32'hbf427846} /* (15, 19, 23) {real, imag} */,
  {32'hbfc44480, 32'h404b9454} /* (15, 19, 22) {real, imag} */,
  {32'hbfd59a10, 32'h40295666} /* (15, 19, 21) {real, imag} */,
  {32'hbf707c87, 32'h40d33fb0} /* (15, 19, 20) {real, imag} */,
  {32'h3f251f34, 32'hbff46b84} /* (15, 19, 19) {real, imag} */,
  {32'hc0a24aea, 32'h40843535} /* (15, 19, 18) {real, imag} */,
  {32'h4043fe86, 32'h402f7fe4} /* (15, 19, 17) {real, imag} */,
  {32'h3f39c920, 32'hbf445c58} /* (15, 19, 16) {real, imag} */,
  {32'hc09dc075, 32'hc001d056} /* (15, 19, 15) {real, imag} */,
  {32'hc0292892, 32'hbff61718} /* (15, 19, 14) {real, imag} */,
  {32'hc0a2b6da, 32'hc102a52a} /* (15, 19, 13) {real, imag} */,
  {32'h3d1eabf0, 32'h400e9250} /* (15, 19, 12) {real, imag} */,
  {32'h407a70d8, 32'hbe985694} /* (15, 19, 11) {real, imag} */,
  {32'h3fffad60, 32'h4111b793} /* (15, 19, 10) {real, imag} */,
  {32'h408840e2, 32'h4039576c} /* (15, 19, 9) {real, imag} */,
  {32'h410b27b5, 32'h40d9ec70} /* (15, 19, 8) {real, imag} */,
  {32'h40a9d8a0, 32'hbfc4869f} /* (15, 19, 7) {real, imag} */,
  {32'h40131171, 32'h3fe615d0} /* (15, 19, 6) {real, imag} */,
  {32'h4095197a, 32'hc1402e22} /* (15, 19, 5) {real, imag} */,
  {32'hc0915716, 32'h415c8e66} /* (15, 19, 4) {real, imag} */,
  {32'hc10d8946, 32'h40b893b8} /* (15, 19, 3) {real, imag} */,
  {32'hc110097e, 32'h40a05338} /* (15, 19, 2) {real, imag} */,
  {32'h40bbb3d5, 32'hc04e4fdd} /* (15, 19, 1) {real, imag} */,
  {32'hbfee2104, 32'h40626a8e} /* (15, 19, 0) {real, imag} */,
  {32'h3fe25118, 32'h3f2cfaa4} /* (15, 18, 31) {real, imag} */,
  {32'h4135d21a, 32'h408e3c6e} /* (15, 18, 30) {real, imag} */,
  {32'hbfa42044, 32'h3fcca574} /* (15, 18, 29) {real, imag} */,
  {32'h41210ccb, 32'h411df6ae} /* (15, 18, 28) {real, imag} */,
  {32'h40032cc0, 32'h40420812} /* (15, 18, 27) {real, imag} */,
  {32'h412c52b4, 32'h3fd536c0} /* (15, 18, 26) {real, imag} */,
  {32'h4186b59a, 32'h3eb1d800} /* (15, 18, 25) {real, imag} */,
  {32'h409b878a, 32'hc0b7b1dc} /* (15, 18, 24) {real, imag} */,
  {32'hc00050bf, 32'hbf77b240} /* (15, 18, 23) {real, imag} */,
  {32'hbf45b102, 32'hc08a93c6} /* (15, 18, 22) {real, imag} */,
  {32'h40b368d7, 32'h40085022} /* (15, 18, 21) {real, imag} */,
  {32'hbed1eb60, 32'h40b6077a} /* (15, 18, 20) {real, imag} */,
  {32'hc0e0e024, 32'h406d10fc} /* (15, 18, 19) {real, imag} */,
  {32'h3ff0c539, 32'hbf33b07a} /* (15, 18, 18) {real, imag} */,
  {32'hc0bda902, 32'h402da07f} /* (15, 18, 17) {real, imag} */,
  {32'hbff4173c, 32'hbf992676} /* (15, 18, 16) {real, imag} */,
  {32'h3fba7bb8, 32'h3f59f9ec} /* (15, 18, 15) {real, imag} */,
  {32'hbfec72c1, 32'h401366ac} /* (15, 18, 14) {real, imag} */,
  {32'hbf890a96, 32'h3eb0d220} /* (15, 18, 13) {real, imag} */,
  {32'h3f153d88, 32'hbe7da9c0} /* (15, 18, 12) {real, imag} */,
  {32'h3f022cf0, 32'hc0dabce3} /* (15, 18, 11) {real, imag} */,
  {32'h3ff6acbd, 32'hc0dc22be} /* (15, 18, 10) {real, imag} */,
  {32'hc08a2b20, 32'hc0a1a2ef} /* (15, 18, 9) {real, imag} */,
  {32'h3eb297b8, 32'hc0aed2b8} /* (15, 18, 8) {real, imag} */,
  {32'h414b6070, 32'hc119c908} /* (15, 18, 7) {real, imag} */,
  {32'h40b05d38, 32'hc12b407e} /* (15, 18, 6) {real, imag} */,
  {32'h41576054, 32'h40fdbd9b} /* (15, 18, 5) {real, imag} */,
  {32'hbf512cf0, 32'hc0dae5f8} /* (15, 18, 4) {real, imag} */,
  {32'hc0d3f2ca, 32'hc0dc3a55} /* (15, 18, 3) {real, imag} */,
  {32'h413debc6, 32'hc0a09a96} /* (15, 18, 2) {real, imag} */,
  {32'h4178aa4f, 32'h40be1b36} /* (15, 18, 1) {real, imag} */,
  {32'h3d93d598, 32'hc0eff366} /* (15, 18, 0) {real, imag} */,
  {32'hc0bae42d, 32'h41167908} /* (15, 17, 31) {real, imag} */,
  {32'h40b2369d, 32'h3f713e7a} /* (15, 17, 30) {real, imag} */,
  {32'h3ef6a490, 32'h40a3e25d} /* (15, 17, 29) {real, imag} */,
  {32'hbdda24e0, 32'hc05cfac6} /* (15, 17, 28) {real, imag} */,
  {32'h3eadfe5a, 32'hc0faa9d6} /* (15, 17, 27) {real, imag} */,
  {32'h40299dc9, 32'h404ca372} /* (15, 17, 26) {real, imag} */,
  {32'hbefd6370, 32'h40a023a4} /* (15, 17, 25) {real, imag} */,
  {32'h3e5798e8, 32'hc0bc46eb} /* (15, 17, 24) {real, imag} */,
  {32'hc101efac, 32'h3f36f47c} /* (15, 17, 23) {real, imag} */,
  {32'hbef9d098, 32'h41035078} /* (15, 17, 22) {real, imag} */,
  {32'hbfc50878, 32'h3f9f7790} /* (15, 17, 21) {real, imag} */,
  {32'hbfea5e88, 32'h3f6fbbe0} /* (15, 17, 20) {real, imag} */,
  {32'hbeb856f6, 32'hbf0b701a} /* (15, 17, 19) {real, imag} */,
  {32'hc06597ae, 32'hbf2ca10e} /* (15, 17, 18) {real, imag} */,
  {32'h3f84a017, 32'hbf84716e} /* (15, 17, 17) {real, imag} */,
  {32'h40134f2c, 32'hbf346b10} /* (15, 17, 16) {real, imag} */,
  {32'h4022d08c, 32'hbf82f522} /* (15, 17, 15) {real, imag} */,
  {32'h40051822, 32'hbeb238d4} /* (15, 17, 14) {real, imag} */,
  {32'h3ff272de, 32'h405f5dae} /* (15, 17, 13) {real, imag} */,
  {32'h4109914b, 32'h405f3c30} /* (15, 17, 12) {real, imag} */,
  {32'hc0194324, 32'hbf89c484} /* (15, 17, 11) {real, imag} */,
  {32'hc0dec768, 32'h3fabb7b4} /* (15, 17, 10) {real, imag} */,
  {32'hbff101bc, 32'hbfd20a3e} /* (15, 17, 9) {real, imag} */,
  {32'hbfccfabb, 32'hbfd02244} /* (15, 17, 8) {real, imag} */,
  {32'hc12c7cb8, 32'hbfe4e752} /* (15, 17, 7) {real, imag} */,
  {32'h4084164e, 32'hbfd7c90c} /* (15, 17, 6) {real, imag} */,
  {32'h3e64c793, 32'hbfa98d5a} /* (15, 17, 5) {real, imag} */,
  {32'hbfdb1f72, 32'h3f689278} /* (15, 17, 4) {real, imag} */,
  {32'h409c2837, 32'hbeaa9610} /* (15, 17, 3) {real, imag} */,
  {32'hc07c0806, 32'hbfe24975} /* (15, 17, 2) {real, imag} */,
  {32'h40ad6f9b, 32'h413cda9e} /* (15, 17, 1) {real, imag} */,
  {32'hbf1bb390, 32'h410fdfbc} /* (15, 17, 0) {real, imag} */,
  {32'hc10c98be, 32'hbdbf9680} /* (15, 16, 31) {real, imag} */,
  {32'hbfe82fd7, 32'hbfdd02ef} /* (15, 16, 30) {real, imag} */,
  {32'hc068b4d1, 32'hc1361be0} /* (15, 16, 29) {real, imag} */,
  {32'hc107d0a8, 32'hc0b45150} /* (15, 16, 28) {real, imag} */,
  {32'hc0749aaf, 32'hc0b5482f} /* (15, 16, 27) {real, imag} */,
  {32'hc08b3cf4, 32'h40e75c10} /* (15, 16, 26) {real, imag} */,
  {32'hc090cc36, 32'h3e8423cc} /* (15, 16, 25) {real, imag} */,
  {32'hc08bc24d, 32'hc08310a4} /* (15, 16, 24) {real, imag} */,
  {32'hbe72d760, 32'hc11f6176} /* (15, 16, 23) {real, imag} */,
  {32'h412ca1ea, 32'hc0c74f42} /* (15, 16, 22) {real, imag} */,
  {32'hbfa161e4, 32'h3ebaa8b0} /* (15, 16, 21) {real, imag} */,
  {32'h3fe0dda5, 32'h4005a646} /* (15, 16, 20) {real, imag} */,
  {32'h4047c620, 32'hc02da9c0} /* (15, 16, 19) {real, imag} */,
  {32'hbf1be3ae, 32'h3efe83cc} /* (15, 16, 18) {real, imag} */,
  {32'hbf40b66c, 32'h3e3dcae8} /* (15, 16, 17) {real, imag} */,
  {32'h3f5f4498, 32'h3e5aae10} /* (15, 16, 16) {real, imag} */,
  {32'hbf369a0c, 32'hbe5e1ef8} /* (15, 16, 15) {real, imag} */,
  {32'hc0286602, 32'h40445d32} /* (15, 16, 14) {real, imag} */,
  {32'hc03f1d66, 32'hbfdc6c28} /* (15, 16, 13) {real, imag} */,
  {32'hc02f8352, 32'hc04f514e} /* (15, 16, 12) {real, imag} */,
  {32'h3fa40ee4, 32'hc0fd03c1} /* (15, 16, 11) {real, imag} */,
  {32'h40012270, 32'h4115ab0c} /* (15, 16, 10) {real, imag} */,
  {32'hc0985777, 32'h3fb8910c} /* (15, 16, 9) {real, imag} */,
  {32'h40de7adf, 32'hc011b1f4} /* (15, 16, 8) {real, imag} */,
  {32'hc01cc458, 32'hc074730a} /* (15, 16, 7) {real, imag} */,
  {32'h40eeab40, 32'hbfb67866} /* (15, 16, 6) {real, imag} */,
  {32'h40f09a2a, 32'h412d740a} /* (15, 16, 5) {real, imag} */,
  {32'h4000eeca, 32'h40729a01} /* (15, 16, 4) {real, imag} */,
  {32'h4002fc19, 32'hc12b8318} /* (15, 16, 3) {real, imag} */,
  {32'h40497eb4, 32'h40ab11a0} /* (15, 16, 2) {real, imag} */,
  {32'h4072de22, 32'h40862dc2} /* (15, 16, 1) {real, imag} */,
  {32'h4005e3f9, 32'h4092a30a} /* (15, 16, 0) {real, imag} */,
  {32'hbfb90338, 32'hc09cf01f} /* (15, 15, 31) {real, imag} */,
  {32'hbf179358, 32'h3f8f928b} /* (15, 15, 30) {real, imag} */,
  {32'h4081e70f, 32'h4092940d} /* (15, 15, 29) {real, imag} */,
  {32'h4053b7e3, 32'hc0a9ad82} /* (15, 15, 28) {real, imag} */,
  {32'h4103ffb5, 32'h40bfeaf7} /* (15, 15, 27) {real, imag} */,
  {32'hbfe52c74, 32'h40630084} /* (15, 15, 26) {real, imag} */,
  {32'h40c07fa0, 32'h4109f24c} /* (15, 15, 25) {real, imag} */,
  {32'h3fafacb3, 32'hc07aa89a} /* (15, 15, 24) {real, imag} */,
  {32'h3f141f44, 32'h405b322f} /* (15, 15, 23) {real, imag} */,
  {32'hc0544bf9, 32'hbf8d7738} /* (15, 15, 22) {real, imag} */,
  {32'hc073d6aa, 32'hc08f2006} /* (15, 15, 21) {real, imag} */,
  {32'h40899fb0, 32'hbfa20859} /* (15, 15, 20) {real, imag} */,
  {32'h3f783d0c, 32'h3fcbc8d8} /* (15, 15, 19) {real, imag} */,
  {32'h3f6c9010, 32'h40536822} /* (15, 15, 18) {real, imag} */,
  {32'h3f8342dd, 32'hbf92db0b} /* (15, 15, 17) {real, imag} */,
  {32'h3f04aada, 32'hbda70390} /* (15, 15, 16) {real, imag} */,
  {32'h3f5f2fd2, 32'h405ec708} /* (15, 15, 15) {real, imag} */,
  {32'h402037ce, 32'hbfc187f3} /* (15, 15, 14) {real, imag} */,
  {32'h3fae2386, 32'h3fa83b08} /* (15, 15, 13) {real, imag} */,
  {32'h408aa7ee, 32'h408626c4} /* (15, 15, 12) {real, imag} */,
  {32'hc07ab32a, 32'h402f0866} /* (15, 15, 11) {real, imag} */,
  {32'h40cf0fd6, 32'h40a68552} /* (15, 15, 10) {real, imag} */,
  {32'hbf9d745a, 32'h3ff2c91e} /* (15, 15, 9) {real, imag} */,
  {32'h3f5d6d9a, 32'hc046871e} /* (15, 15, 8) {real, imag} */,
  {32'hbff42824, 32'hc02aa355} /* (15, 15, 7) {real, imag} */,
  {32'h4034da2e, 32'h41521087} /* (15, 15, 6) {real, imag} */,
  {32'h40874fd4, 32'hc10c567e} /* (15, 15, 5) {real, imag} */,
  {32'h403591fd, 32'hbc95f000} /* (15, 15, 4) {real, imag} */,
  {32'hbf0fd9e8, 32'hbf92467c} /* (15, 15, 3) {real, imag} */,
  {32'hc0a67f2c, 32'h409c316f} /* (15, 15, 2) {real, imag} */,
  {32'hbffdf6ba, 32'h41009bd4} /* (15, 15, 1) {real, imag} */,
  {32'hbfc4d5f5, 32'hc04e0c4c} /* (15, 15, 0) {real, imag} */,
  {32'h3f5bfd58, 32'h404fa6a7} /* (15, 14, 31) {real, imag} */,
  {32'hc01b3b80, 32'h4185be9a} /* (15, 14, 30) {real, imag} */,
  {32'h40b378f2, 32'hc02572db} /* (15, 14, 29) {real, imag} */,
  {32'hbfa6e180, 32'h40bfc562} /* (15, 14, 28) {real, imag} */,
  {32'h404537ec, 32'hc152f985} /* (15, 14, 27) {real, imag} */,
  {32'hc0a2c1fe, 32'hc0d5b55f} /* (15, 14, 26) {real, imag} */,
  {32'hc0e1ca20, 32'hc0a54cac} /* (15, 14, 25) {real, imag} */,
  {32'h3d4c3f00, 32'h40fa2e7f} /* (15, 14, 24) {real, imag} */,
  {32'h40d295d8, 32'hbdff7b00} /* (15, 14, 23) {real, imag} */,
  {32'hbf6ed842, 32'hbfdf8a81} /* (15, 14, 22) {real, imag} */,
  {32'hbf4b0756, 32'h3e3ae910} /* (15, 14, 21) {real, imag} */,
  {32'hc084b930, 32'hbf956492} /* (15, 14, 20) {real, imag} */,
  {32'hbf118e54, 32'hc03f6031} /* (15, 14, 19) {real, imag} */,
  {32'hbf0f3498, 32'h407b46b4} /* (15, 14, 18) {real, imag} */,
  {32'hbfee9d3d, 32'hbf8faf8e} /* (15, 14, 17) {real, imag} */,
  {32'hbff461cc, 32'hc098a922} /* (15, 14, 16) {real, imag} */,
  {32'h3fd23beb, 32'hbfac5c42} /* (15, 14, 15) {real, imag} */,
  {32'hbfaa9998, 32'h3faee6e8} /* (15, 14, 14) {real, imag} */,
  {32'h3f48585c, 32'h4017f613} /* (15, 14, 13) {real, imag} */,
  {32'h4078b120, 32'hbfe0e75a} /* (15, 14, 12) {real, imag} */,
  {32'hc035ba7a, 32'hc02eaef9} /* (15, 14, 11) {real, imag} */,
  {32'hc046e41e, 32'h408d64e6} /* (15, 14, 10) {real, imag} */,
  {32'h40affc84, 32'h41142e74} /* (15, 14, 9) {real, imag} */,
  {32'h3e4bc220, 32'hc04cdb96} /* (15, 14, 8) {real, imag} */,
  {32'h402d4b41, 32'hc053a480} /* (15, 14, 7) {real, imag} */,
  {32'hbf84262a, 32'h401d5f3a} /* (15, 14, 6) {real, imag} */,
  {32'hc0616ef0, 32'hc1539c01} /* (15, 14, 5) {real, imag} */,
  {32'h40bb77d2, 32'hc10d38a7} /* (15, 14, 4) {real, imag} */,
  {32'hc1767073, 32'hbfad5106} /* (15, 14, 3) {real, imag} */,
  {32'hc140a308, 32'h3f3c58b0} /* (15, 14, 2) {real, imag} */,
  {32'h408dea9b, 32'h3f25b1c4} /* (15, 14, 1) {real, imag} */,
  {32'h413b8b06, 32'hc182a1ba} /* (15, 14, 0) {real, imag} */,
  {32'hc13b4c4f, 32'h40c355d4} /* (15, 13, 31) {real, imag} */,
  {32'h3fc14980, 32'hc1737f57} /* (15, 13, 30) {real, imag} */,
  {32'h3d1db980, 32'hc10b66ec} /* (15, 13, 29) {real, imag} */,
  {32'h414aa0d2, 32'h4008dcc0} /* (15, 13, 28) {real, imag} */,
  {32'h403d6996, 32'hc0a21b9e} /* (15, 13, 27) {real, imag} */,
  {32'h4094edac, 32'hc088086e} /* (15, 13, 26) {real, imag} */,
  {32'hc0abd664, 32'h403b48e4} /* (15, 13, 25) {real, imag} */,
  {32'hbf5d053c, 32'h40e68f3b} /* (15, 13, 24) {real, imag} */,
  {32'hc113c685, 32'hbfcec384} /* (15, 13, 23) {real, imag} */,
  {32'h3fa61d82, 32'hc0cd9171} /* (15, 13, 22) {real, imag} */,
  {32'hc07aa538, 32'hbf7fda1c} /* (15, 13, 21) {real, imag} */,
  {32'hbff07e88, 32'h400e34aa} /* (15, 13, 20) {real, imag} */,
  {32'hc0a1b610, 32'hc01db244} /* (15, 13, 19) {real, imag} */,
  {32'hbe2cc080, 32'h409b7817} /* (15, 13, 18) {real, imag} */,
  {32'hbfc80a3c, 32'h4030d76c} /* (15, 13, 17) {real, imag} */,
  {32'h3fb0a4bc, 32'h3e559b20} /* (15, 13, 16) {real, imag} */,
  {32'h40b53fdf, 32'hc00c9830} /* (15, 13, 15) {real, imag} */,
  {32'hbfb55f58, 32'h40c70855} /* (15, 13, 14) {real, imag} */,
  {32'hc0a1bd06, 32'h401bd7e0} /* (15, 13, 13) {real, imag} */,
  {32'hc0ca6f68, 32'h40146cbc} /* (15, 13, 12) {real, imag} */,
  {32'h40a891cc, 32'hc0536f91} /* (15, 13, 11) {real, imag} */,
  {32'hc067dfb9, 32'h3faa2f5c} /* (15, 13, 10) {real, imag} */,
  {32'h41065441, 32'hc10318f8} /* (15, 13, 9) {real, imag} */,
  {32'hc0544af5, 32'h41034fbe} /* (15, 13, 8) {real, imag} */,
  {32'hc03889cf, 32'hc04867ec} /* (15, 13, 7) {real, imag} */,
  {32'h40b45a58, 32'hc1458e3d} /* (15, 13, 6) {real, imag} */,
  {32'h3ec68ba4, 32'h40bd3f3e} /* (15, 13, 5) {real, imag} */,
  {32'hbed40ae0, 32'hc12da23a} /* (15, 13, 4) {real, imag} */,
  {32'h40c6242f, 32'hc0516406} /* (15, 13, 3) {real, imag} */,
  {32'hc1e3c120, 32'h402986a4} /* (15, 13, 2) {real, imag} */,
  {32'hc159559d, 32'h3f10f290} /* (15, 13, 1) {real, imag} */,
  {32'h404785c6, 32'h410d2e44} /* (15, 13, 0) {real, imag} */,
  {32'h41f319ab, 32'hbf1c7280} /* (15, 12, 31) {real, imag} */,
  {32'h410ccbe9, 32'hc001f282} /* (15, 12, 30) {real, imag} */,
  {32'hc0964508, 32'hc142716e} /* (15, 12, 29) {real, imag} */,
  {32'h40a2b800, 32'h40d2fead} /* (15, 12, 28) {real, imag} */,
  {32'h41940d62, 32'h40acd334} /* (15, 12, 27) {real, imag} */,
  {32'h410e056d, 32'h3ed0a268} /* (15, 12, 26) {real, imag} */,
  {32'hc093f9b9, 32'hc0ec2209} /* (15, 12, 25) {real, imag} */,
  {32'hc004bd5a, 32'h411d393d} /* (15, 12, 24) {real, imag} */,
  {32'h40b0eca2, 32'hc0d3228b} /* (15, 12, 23) {real, imag} */,
  {32'h40fa0baa, 32'h40820c03} /* (15, 12, 22) {real, imag} */,
  {32'hbfd45fde, 32'h4080330e} /* (15, 12, 21) {real, imag} */,
  {32'h40580a60, 32'hc100f72e} /* (15, 12, 20) {real, imag} */,
  {32'hc026f219, 32'h4052352f} /* (15, 12, 19) {real, imag} */,
  {32'hc05bc15b, 32'hbcdfe300} /* (15, 12, 18) {real, imag} */,
  {32'h3dd37580, 32'h40f6f35f} /* (15, 12, 17) {real, imag} */,
  {32'hbfc4a72c, 32'h4043971e} /* (15, 12, 16) {real, imag} */,
  {32'hbf1a9b90, 32'hbed0c290} /* (15, 12, 15) {real, imag} */,
  {32'hc04b4441, 32'h3fd1a44c} /* (15, 12, 14) {real, imag} */,
  {32'h3e2512f0, 32'hbecb8188} /* (15, 12, 13) {real, imag} */,
  {32'hbe1c8b88, 32'h4047cdae} /* (15, 12, 12) {real, imag} */,
  {32'hbee9a1b8, 32'h40045543} /* (15, 12, 11) {real, imag} */,
  {32'hc0f4981e, 32'hc096240d} /* (15, 12, 10) {real, imag} */,
  {32'hc0b036fa, 32'h409f34cd} /* (15, 12, 9) {real, imag} */,
  {32'h41110df0, 32'hc0075130} /* (15, 12, 8) {real, imag} */,
  {32'hc0fe0c8b, 32'hc09d3a41} /* (15, 12, 7) {real, imag} */,
  {32'h40a22592, 32'h3feeb7ea} /* (15, 12, 6) {real, imag} */,
  {32'hc124743d, 32'hc08f3774} /* (15, 12, 5) {real, imag} */,
  {32'hc12edad2, 32'hc0c04a91} /* (15, 12, 4) {real, imag} */,
  {32'h40b2573c, 32'h3ee77940} /* (15, 12, 3) {real, imag} */,
  {32'h41686beb, 32'hc11d7a3c} /* (15, 12, 2) {real, imag} */,
  {32'h41269e82, 32'hc05f5138} /* (15, 12, 1) {real, imag} */,
  {32'hc1881fa9, 32'h4131c26c} /* (15, 12, 0) {real, imag} */,
  {32'hbf8ad5f8, 32'h416b9aa5} /* (15, 11, 31) {real, imag} */,
  {32'h3febae11, 32'hc0d5d1da} /* (15, 11, 30) {real, imag} */,
  {32'h4140c32c, 32'h414f7738} /* (15, 11, 29) {real, imag} */,
  {32'hc150a06c, 32'hbff3dc38} /* (15, 11, 28) {real, imag} */,
  {32'hc0ba78d1, 32'hbe0353e0} /* (15, 11, 27) {real, imag} */,
  {32'hc046e69a, 32'h3ed1aed4} /* (15, 11, 26) {real, imag} */,
  {32'h4174e2f2, 32'hc0b762ee} /* (15, 11, 25) {real, imag} */,
  {32'hc03ada6e, 32'h411fb3f2} /* (15, 11, 24) {real, imag} */,
  {32'hc11f4d93, 32'h40d07df8} /* (15, 11, 23) {real, imag} */,
  {32'hc153985e, 32'hbeedda4a} /* (15, 11, 22) {real, imag} */,
  {32'hc0bb3a81, 32'hbf80de3e} /* (15, 11, 21) {real, imag} */,
  {32'h40a2d600, 32'hbf817254} /* (15, 11, 20) {real, imag} */,
  {32'hbfe499ca, 32'h410d36d5} /* (15, 11, 19) {real, imag} */,
  {32'h3fccbce8, 32'hbedcb930} /* (15, 11, 18) {real, imag} */,
  {32'h3efa5540, 32'hc0289721} /* (15, 11, 17) {real, imag} */,
  {32'h4084ffc4, 32'hc0c87aa7} /* (15, 11, 16) {real, imag} */,
  {32'h3f827380, 32'hbf2cffbc} /* (15, 11, 15) {real, imag} */,
  {32'h4067fe98, 32'hbd523980} /* (15, 11, 14) {real, imag} */,
  {32'h400dc297, 32'hc000ce51} /* (15, 11, 13) {real, imag} */,
  {32'hc09574b2, 32'h411538d8} /* (15, 11, 12) {real, imag} */,
  {32'hbf91d7c4, 32'h3f0a678c} /* (15, 11, 11) {real, imag} */,
  {32'hbeaf66a0, 32'h400d9fe2} /* (15, 11, 10) {real, imag} */,
  {32'h410ff8a1, 32'hbfaae68e} /* (15, 11, 9) {real, imag} */,
  {32'hc16cdf14, 32'hc14f5e60} /* (15, 11, 8) {real, imag} */,
  {32'h4137bb5c, 32'h4005fd55} /* (15, 11, 7) {real, imag} */,
  {32'h41641e3e, 32'h40571546} /* (15, 11, 6) {real, imag} */,
  {32'h4186364c, 32'hc115dbe2} /* (15, 11, 5) {real, imag} */,
  {32'hc118f0b0, 32'hc196e1a0} /* (15, 11, 4) {real, imag} */,
  {32'hbddd1040, 32'hc0f3d840} /* (15, 11, 3) {real, imag} */,
  {32'h4047bc5c, 32'h4029d754} /* (15, 11, 2) {real, imag} */,
  {32'h414a1a09, 32'h40aa126e} /* (15, 11, 1) {real, imag} */,
  {32'h40bc15c4, 32'h4151c4e4} /* (15, 11, 0) {real, imag} */,
  {32'h4092f1f8, 32'h415db832} /* (15, 10, 31) {real, imag} */,
  {32'h41c091b4, 32'hc115d072} /* (15, 10, 30) {real, imag} */,
  {32'hc0b495a2, 32'hc0f0be48} /* (15, 10, 29) {real, imag} */,
  {32'h4000aaab, 32'h40d65818} /* (15, 10, 28) {real, imag} */,
  {32'h4081bed4, 32'h418da79b} /* (15, 10, 27) {real, imag} */,
  {32'h407d38b8, 32'h4141e89a} /* (15, 10, 26) {real, imag} */,
  {32'hc100b448, 32'hc1a24bc5} /* (15, 10, 25) {real, imag} */,
  {32'hc0b005ce, 32'h40bb27ff} /* (15, 10, 24) {real, imag} */,
  {32'h413a5cad, 32'hc1927758} /* (15, 10, 23) {real, imag} */,
  {32'hc1a88363, 32'hc0c42463} /* (15, 10, 22) {real, imag} */,
  {32'h3f46a52e, 32'h3f2df840} /* (15, 10, 21) {real, imag} */,
  {32'h40cc2659, 32'h40b7c0dc} /* (15, 10, 20) {real, imag} */,
  {32'h4052e6f8, 32'hbf631700} /* (15, 10, 19) {real, imag} */,
  {32'hc09297f7, 32'h40062266} /* (15, 10, 18) {real, imag} */,
  {32'hc086e2f1, 32'h3fa404f8} /* (15, 10, 17) {real, imag} */,
  {32'h406c1904, 32'hc011887c} /* (15, 10, 16) {real, imag} */,
  {32'hc064fa80, 32'hbaafa000} /* (15, 10, 15) {real, imag} */,
  {32'hc02e230a, 32'hc093db21} /* (15, 10, 14) {real, imag} */,
  {32'h408b28b2, 32'hc10f1552} /* (15, 10, 13) {real, imag} */,
  {32'hbfcf99ec, 32'h40e72448} /* (15, 10, 12) {real, imag} */,
  {32'hc04c31a6, 32'h3f905730} /* (15, 10, 11) {real, imag} */,
  {32'hbf9cbe30, 32'h41515d84} /* (15, 10, 10) {real, imag} */,
  {32'h40fe433a, 32'hc06a4732} /* (15, 10, 9) {real, imag} */,
  {32'hc126218f, 32'h40890ce9} /* (15, 10, 8) {real, imag} */,
  {32'hc0e532eb, 32'h408634cc} /* (15, 10, 7) {real, imag} */,
  {32'h41441e7e, 32'h4178cd72} /* (15, 10, 6) {real, imag} */,
  {32'h40580328, 32'hc129e04c} /* (15, 10, 5) {real, imag} */,
  {32'hc0b9b534, 32'h41b01eed} /* (15, 10, 4) {real, imag} */,
  {32'h3ec91100, 32'hc0c6f83c} /* (15, 10, 3) {real, imag} */,
  {32'h40081adc, 32'hc11eea7e} /* (15, 10, 2) {real, imag} */,
  {32'hc11a2328, 32'h40dd6659} /* (15, 10, 1) {real, imag} */,
  {32'hc1534347, 32'hbf140369} /* (15, 10, 0) {real, imag} */,
  {32'h3fbf4f90, 32'h416696aa} /* (15, 9, 31) {real, imag} */,
  {32'h3f825288, 32'hc11760a4} /* (15, 9, 30) {real, imag} */,
  {32'hc0cf658f, 32'h408f1bf3} /* (15, 9, 29) {real, imag} */,
  {32'h3eae0190, 32'hc1495b9a} /* (15, 9, 28) {real, imag} */,
  {32'h41d0ace8, 32'h40e97765} /* (15, 9, 27) {real, imag} */,
  {32'h403dd8dc, 32'hc0b94a0e} /* (15, 9, 26) {real, imag} */,
  {32'hc0a7a8e2, 32'h3ef24770} /* (15, 9, 25) {real, imag} */,
  {32'hc1b37fe9, 32'h4178333e} /* (15, 9, 24) {real, imag} */,
  {32'h40cbe9f5, 32'h411aaa5e} /* (15, 9, 23) {real, imag} */,
  {32'h4187ee97, 32'hc1a84bb2} /* (15, 9, 22) {real, imag} */,
  {32'hc1930623, 32'h410b66ac} /* (15, 9, 21) {real, imag} */,
  {32'hbeb423d0, 32'h40ec1d79} /* (15, 9, 20) {real, imag} */,
  {32'hbf9120bc, 32'h40420b0c} /* (15, 9, 19) {real, imag} */,
  {32'h3e5c41c0, 32'h404b600b} /* (15, 9, 18) {real, imag} */,
  {32'hc051061c, 32'hc01f463a} /* (15, 9, 17) {real, imag} */,
  {32'hc08a0177, 32'hc029cfc9} /* (15, 9, 16) {real, imag} */,
  {32'hc0a7e33c, 32'hc0aab2a7} /* (15, 9, 15) {real, imag} */,
  {32'hc0a07c24, 32'h4121f29b} /* (15, 9, 14) {real, imag} */,
  {32'h402f6b2e, 32'h40b634d4} /* (15, 9, 13) {real, imag} */,
  {32'hc1345b68, 32'hc05ac882} /* (15, 9, 12) {real, imag} */,
  {32'hc0ec90f1, 32'hc0b621b2} /* (15, 9, 11) {real, imag} */,
  {32'h41f253e5, 32'hc11402c3} /* (15, 9, 10) {real, imag} */,
  {32'h412d3d2e, 32'h41ac5179} /* (15, 9, 9) {real, imag} */,
  {32'hc1b396ff, 32'hc12e99ce} /* (15, 9, 8) {real, imag} */,
  {32'h413332bf, 32'hc01c427e} /* (15, 9, 7) {real, imag} */,
  {32'h41095fd3, 32'h41fe1d78} /* (15, 9, 6) {real, imag} */,
  {32'h3f5dc7b0, 32'hc1236626} /* (15, 9, 5) {real, imag} */,
  {32'hc08f001d, 32'hc19047eb} /* (15, 9, 4) {real, imag} */,
  {32'h416cb420, 32'hc14519fe} /* (15, 9, 3) {real, imag} */,
  {32'h40edd4a8, 32'hc1c124d2} /* (15, 9, 2) {real, imag} */,
  {32'h419ad64f, 32'h41735024} /* (15, 9, 1) {real, imag} */,
  {32'h40aab087, 32'h3f74f050} /* (15, 9, 0) {real, imag} */,
  {32'h40c0147c, 32'hc10472df} /* (15, 8, 31) {real, imag} */,
  {32'hbe338c40, 32'hc03fe330} /* (15, 8, 30) {real, imag} */,
  {32'h3f8a5598, 32'hc1b8d5e2} /* (15, 8, 29) {real, imag} */,
  {32'h41b743ec, 32'h42134666} /* (15, 8, 28) {real, imag} */,
  {32'h4151fa0f, 32'h417d1794} /* (15, 8, 27) {real, imag} */,
  {32'h41bed170, 32'h419e27c5} /* (15, 8, 26) {real, imag} */,
  {32'hc1523057, 32'hc179f242} /* (15, 8, 25) {real, imag} */,
  {32'hc115078a, 32'hc1958126} /* (15, 8, 24) {real, imag} */,
  {32'hc11dfeaf, 32'h418e9e4c} /* (15, 8, 23) {real, imag} */,
  {32'h41922848, 32'h40dd5364} /* (15, 8, 22) {real, imag} */,
  {32'h40c0142e, 32'h402a77aa} /* (15, 8, 21) {real, imag} */,
  {32'h415a0145, 32'h40a3b5fc} /* (15, 8, 20) {real, imag} */,
  {32'hbfb05b10, 32'h3fcda9b6} /* (15, 8, 19) {real, imag} */,
  {32'h3e864860, 32'hc05eec0d} /* (15, 8, 18) {real, imag} */,
  {32'hc02eb4a4, 32'h3f51db1e} /* (15, 8, 17) {real, imag} */,
  {32'h40def9f4, 32'h410c661a} /* (15, 8, 16) {real, imag} */,
  {32'hc0156894, 32'h40358e12} /* (15, 8, 15) {real, imag} */,
  {32'h4112ee55, 32'hc031e48d} /* (15, 8, 14) {real, imag} */,
  {32'h4075ceb4, 32'hc0d42fde} /* (15, 8, 13) {real, imag} */,
  {32'hc126b045, 32'h40f10fac} /* (15, 8, 12) {real, imag} */,
  {32'h408d74da, 32'hc0e027d5} /* (15, 8, 11) {real, imag} */,
  {32'h400111fc, 32'h418e78a1} /* (15, 8, 10) {real, imag} */,
  {32'hc102f645, 32'h411babdc} /* (15, 8, 9) {real, imag} */,
  {32'hc0e2b65c, 32'h4175b060} /* (15, 8, 8) {real, imag} */,
  {32'hc1b9cb62, 32'h41008718} /* (15, 8, 7) {real, imag} */,
  {32'hbfaf6798, 32'hc1b74079} /* (15, 8, 6) {real, imag} */,
  {32'h40c76d7e, 32'h41548ac4} /* (15, 8, 5) {real, imag} */,
  {32'h421e4462, 32'hc19f981d} /* (15, 8, 4) {real, imag} */,
  {32'h4138d054, 32'h410380f5} /* (15, 8, 3) {real, imag} */,
  {32'hc1528d7b, 32'hc18c81e8} /* (15, 8, 2) {real, imag} */,
  {32'hc22418d4, 32'hc0f628e5} /* (15, 8, 1) {real, imag} */,
  {32'hc210fdca, 32'h3fa8f78c} /* (15, 8, 0) {real, imag} */,
  {32'hc1ce8ecd, 32'h4243b38a} /* (15, 7, 31) {real, imag} */,
  {32'h41ed63f6, 32'h41969601} /* (15, 7, 30) {real, imag} */,
  {32'hc08d659e, 32'hc1934cd7} /* (15, 7, 29) {real, imag} */,
  {32'hc10fe179, 32'h40c84ec8} /* (15, 7, 28) {real, imag} */,
  {32'h409dde4e, 32'hbf5d3010} /* (15, 7, 27) {real, imag} */,
  {32'hc2181047, 32'h40c97461} /* (15, 7, 26) {real, imag} */,
  {32'hc0d3f0df, 32'hc1ab6301} /* (15, 7, 25) {real, imag} */,
  {32'hc0c2a40c, 32'hbf3e2810} /* (15, 7, 24) {real, imag} */,
  {32'hc0a3b319, 32'hc1292504} /* (15, 7, 23) {real, imag} */,
  {32'hc1a0c636, 32'h3fbc5ee0} /* (15, 7, 22) {real, imag} */,
  {32'h40893438, 32'h417cf0aa} /* (15, 7, 21) {real, imag} */,
  {32'h40ee0c3a, 32'hc0523e32} /* (15, 7, 20) {real, imag} */,
  {32'h41849b38, 32'h41373ac4} /* (15, 7, 19) {real, imag} */,
  {32'h4043e398, 32'h40873a1f} /* (15, 7, 18) {real, imag} */,
  {32'h3f4c9b20, 32'hc0e6da1a} /* (15, 7, 17) {real, imag} */,
  {32'h3f399078, 32'h400f79c0} /* (15, 7, 16) {real, imag} */,
  {32'h409fa4ac, 32'hc0028a0c} /* (15, 7, 15) {real, imag} */,
  {32'hc06567c8, 32'hc07805d6} /* (15, 7, 14) {real, imag} */,
  {32'hbfbf8f44, 32'hbf515280} /* (15, 7, 13) {real, imag} */,
  {32'hc055dfc9, 32'hc118fc7c} /* (15, 7, 12) {real, imag} */,
  {32'h4085c0c4, 32'h40fa40e3} /* (15, 7, 11) {real, imag} */,
  {32'h4127fbb9, 32'hc1ac6c6e} /* (15, 7, 10) {real, imag} */,
  {32'h4198709e, 32'h41356ede} /* (15, 7, 9) {real, imag} */,
  {32'hc12c932c, 32'hbf9efe60} /* (15, 7, 8) {real, imag} */,
  {32'h3ea20010, 32'h415de53f} /* (15, 7, 7) {real, imag} */,
  {32'hc202ec25, 32'h3fa30ad4} /* (15, 7, 6) {real, imag} */,
  {32'h420fec58, 32'h3f9db0d0} /* (15, 7, 5) {real, imag} */,
  {32'h4164cc2b, 32'hc2110a6d} /* (15, 7, 4) {real, imag} */,
  {32'h412acfa6, 32'hc0224268} /* (15, 7, 3) {real, imag} */,
  {32'h4238be99, 32'h41b5097b} /* (15, 7, 2) {real, imag} */,
  {32'h40ebd674, 32'h42161c40} /* (15, 7, 1) {real, imag} */,
  {32'hbf0fbb18, 32'h417f60b0} /* (15, 7, 0) {real, imag} */,
  {32'hc169af8c, 32'h40e248cc} /* (15, 6, 31) {real, imag} */,
  {32'h40029c6a, 32'h41d7e9ce} /* (15, 6, 30) {real, imag} */,
  {32'h413f1131, 32'h406a91ac} /* (15, 6, 29) {real, imag} */,
  {32'h41bb9d46, 32'h40f92619} /* (15, 6, 28) {real, imag} */,
  {32'h411f66f2, 32'hc221c100} /* (15, 6, 27) {real, imag} */,
  {32'h423dadf1, 32'h3f9ddf80} /* (15, 6, 26) {real, imag} */,
  {32'hc08591cb, 32'h417dad03} /* (15, 6, 25) {real, imag} */,
  {32'hc034b998, 32'hc18daa1e} /* (15, 6, 24) {real, imag} */,
  {32'hc16005bc, 32'hbf9bd448} /* (15, 6, 23) {real, imag} */,
  {32'h41b8127f, 32'h41a23ca2} /* (15, 6, 22) {real, imag} */,
  {32'h41000456, 32'h4112bf88} /* (15, 6, 21) {real, imag} */,
  {32'hc0119d7c, 32'hc06104e2} /* (15, 6, 20) {real, imag} */,
  {32'hbd1d6600, 32'hc11b18d8} /* (15, 6, 19) {real, imag} */,
  {32'h40e41189, 32'h40a978c4} /* (15, 6, 18) {real, imag} */,
  {32'h3e39aa48, 32'h40d787c4} /* (15, 6, 17) {real, imag} */,
  {32'hc03a9b50, 32'hc045e57e} /* (15, 6, 16) {real, imag} */,
  {32'hbf03fbf2, 32'hbfb5e070} /* (15, 6, 15) {real, imag} */,
  {32'h416c4c9c, 32'hc1344d52} /* (15, 6, 14) {real, imag} */,
  {32'h40cc71cc, 32'h4102b224} /* (15, 6, 13) {real, imag} */,
  {32'hc1334a23, 32'h40084312} /* (15, 6, 12) {real, imag} */,
  {32'h4180f398, 32'h407256c2} /* (15, 6, 11) {real, imag} */,
  {32'h3e9e7fc0, 32'h41c58a0e} /* (15, 6, 10) {real, imag} */,
  {32'hc06f4126, 32'hc1d7c494} /* (15, 6, 9) {real, imag} */,
  {32'hc260e66e, 32'hc1b05446} /* (15, 6, 8) {real, imag} */,
  {32'h409c0377, 32'hc09762ae} /* (15, 6, 7) {real, imag} */,
  {32'hc1b106be, 32'h40040258} /* (15, 6, 6) {real, imag} */,
  {32'hc13b55fe, 32'h4134ddd8} /* (15, 6, 5) {real, imag} */,
  {32'h4203c1b3, 32'h4029f8fe} /* (15, 6, 4) {real, imag} */,
  {32'h41953a10, 32'hc197e1b4} /* (15, 6, 3) {real, imag} */,
  {32'h414d02ea, 32'hc13938d0} /* (15, 6, 2) {real, imag} */,
  {32'hc18dff4a, 32'h41acde4d} /* (15, 6, 1) {real, imag} */,
  {32'hc19b076e, 32'hc095f8ef} /* (15, 6, 0) {real, imag} */,
  {32'h41ec2212, 32'hc00c5356} /* (15, 5, 31) {real, imag} */,
  {32'h414d6cfa, 32'h41b1620d} /* (15, 5, 30) {real, imag} */,
  {32'h4015b4a8, 32'h426a615e} /* (15, 5, 29) {real, imag} */,
  {32'h41b6810c, 32'h41077fe6} /* (15, 5, 28) {real, imag} */,
  {32'h41b71596, 32'hc0084368} /* (15, 5, 27) {real, imag} */,
  {32'h4218fdfe, 32'hc2431e41} /* (15, 5, 26) {real, imag} */,
  {32'h4167aa91, 32'h41eaa384} /* (15, 5, 25) {real, imag} */,
  {32'hc10ecbaa, 32'hc0a18c51} /* (15, 5, 24) {real, imag} */,
  {32'hc1300710, 32'h41b1fbca} /* (15, 5, 23) {real, imag} */,
  {32'h3f3d00b8, 32'h41071dde} /* (15, 5, 22) {real, imag} */,
  {32'h40a1f602, 32'h4066fe50} /* (15, 5, 21) {real, imag} */,
  {32'hc08bbebb, 32'h414d7722} /* (15, 5, 20) {real, imag} */,
  {32'hc09a532c, 32'h3e006cc0} /* (15, 5, 19) {real, imag} */,
  {32'h3f9bf6fc, 32'h407aea72} /* (15, 5, 18) {real, imag} */,
  {32'h40096e1e, 32'hc0e98cb1} /* (15, 5, 17) {real, imag} */,
  {32'hc082a2ed, 32'h3fee8920} /* (15, 5, 16) {real, imag} */,
  {32'h3f2726c8, 32'h402955be} /* (15, 5, 15) {real, imag} */,
  {32'hc0ca0885, 32'hc1246674} /* (15, 5, 14) {real, imag} */,
  {32'hc163a7c2, 32'h408956da} /* (15, 5, 13) {real, imag} */,
  {32'h40347636, 32'hc00b45a2} /* (15, 5, 12) {real, imag} */,
  {32'h416d0a29, 32'h414c131c} /* (15, 5, 11) {real, imag} */,
  {32'hc10a0730, 32'h404cd342} /* (15, 5, 10) {real, imag} */,
  {32'hc07bc3e6, 32'hc162a110} /* (15, 5, 9) {real, imag} */,
  {32'h4125e46e, 32'hc1a1599a} /* (15, 5, 8) {real, imag} */,
  {32'h41884e6e, 32'hc181414e} /* (15, 5, 7) {real, imag} */,
  {32'hc04be458, 32'h411188ec} /* (15, 5, 6) {real, imag} */,
  {32'hc1d0869e, 32'hc16a042a} /* (15, 5, 5) {real, imag} */,
  {32'h425e2b7a, 32'hc1c2d317} /* (15, 5, 4) {real, imag} */,
  {32'h4196894f, 32'h421e0bee} /* (15, 5, 3) {real, imag} */,
  {32'hc17190a4, 32'h4210f957} /* (15, 5, 2) {real, imag} */,
  {32'h42370517, 32'hc1190c7a} /* (15, 5, 1) {real, imag} */,
  {32'h419cf64b, 32'hc1e966fc} /* (15, 5, 0) {real, imag} */,
  {32'h4116863e, 32'h423a956a} /* (15, 4, 31) {real, imag} */,
  {32'hbf5fc0cc, 32'h42277768} /* (15, 4, 30) {real, imag} */,
  {32'hc08f3a4a, 32'h3fc7cc90} /* (15, 4, 29) {real, imag} */,
  {32'h41483ad7, 32'hc20ae23d} /* (15, 4, 28) {real, imag} */,
  {32'h409033e0, 32'hc0e3289a} /* (15, 4, 27) {real, imag} */,
  {32'hc1c4b06c, 32'hc1f02fd5} /* (15, 4, 26) {real, imag} */,
  {32'h4257af30, 32'h41c34dd5} /* (15, 4, 25) {real, imag} */,
  {32'hbf3b21b0, 32'hc1618528} /* (15, 4, 24) {real, imag} */,
  {32'h409f3cee, 32'hc0341d16} /* (15, 4, 23) {real, imag} */,
  {32'h415e0948, 32'hbf827ece} /* (15, 4, 22) {real, imag} */,
  {32'h3f0dafa0, 32'h418de56b} /* (15, 4, 21) {real, imag} */,
  {32'h40469520, 32'hc186b83b} /* (15, 4, 20) {real, imag} */,
  {32'hc0f8dcf2, 32'hc034dd94} /* (15, 4, 19) {real, imag} */,
  {32'h40952a35, 32'h41235ca2} /* (15, 4, 18) {real, imag} */,
  {32'h403e717a, 32'hc18c253e} /* (15, 4, 17) {real, imag} */,
  {32'h40446710, 32'h40bba56c} /* (15, 4, 16) {real, imag} */,
  {32'h407a688e, 32'h40dbfd28} /* (15, 4, 15) {real, imag} */,
  {32'h40908be7, 32'hc061a619} /* (15, 4, 14) {real, imag} */,
  {32'h4148ad83, 32'hbfc9a908} /* (15, 4, 13) {real, imag} */,
  {32'hc0dc12ac, 32'h41ac61b9} /* (15, 4, 12) {real, imag} */,
  {32'h41837ad9, 32'hc1a3e541} /* (15, 4, 11) {real, imag} */,
  {32'hc224b478, 32'hc0b19de4} /* (15, 4, 10) {real, imag} */,
  {32'hc12f33d5, 32'h3e932470} /* (15, 4, 9) {real, imag} */,
  {32'hc1514337, 32'hc0b95f14} /* (15, 4, 8) {real, imag} */,
  {32'hc18f5db0, 32'h4150d64e} /* (15, 4, 7) {real, imag} */,
  {32'hbf2c6410, 32'hc1c492c1} /* (15, 4, 6) {real, imag} */,
  {32'h41e17fc6, 32'h41046f81} /* (15, 4, 5) {real, imag} */,
  {32'h41e4462c, 32'h42229067} /* (15, 4, 4) {real, imag} */,
  {32'hc06e7254, 32'hc24c808a} /* (15, 4, 3) {real, imag} */,
  {32'hbe00cbf0, 32'hc23d65ae} /* (15, 4, 2) {real, imag} */,
  {32'h40223302, 32'hc2399962} /* (15, 4, 1) {real, imag} */,
  {32'hc27d6b29, 32'h416504b8} /* (15, 4, 0) {real, imag} */,
  {32'h41b5a643, 32'h4088da44} /* (15, 3, 31) {real, imag} */,
  {32'hc23be015, 32'hc25b277d} /* (15, 3, 30) {real, imag} */,
  {32'h3f0bd938, 32'hc2252466} /* (15, 3, 29) {real, imag} */,
  {32'hc0b092ea, 32'hc01b4e1e} /* (15, 3, 28) {real, imag} */,
  {32'h423f587a, 32'h40e23aed} /* (15, 3, 27) {real, imag} */,
  {32'h41b66056, 32'h4177e451} /* (15, 3, 26) {real, imag} */,
  {32'hc18867c4, 32'h41dc03eb} /* (15, 3, 25) {real, imag} */,
  {32'hc162d92a, 32'hc184eadf} /* (15, 3, 24) {real, imag} */,
  {32'h40c6ded9, 32'h3f4ef2d4} /* (15, 3, 23) {real, imag} */,
  {32'h4199af08, 32'hc003e510} /* (15, 3, 22) {real, imag} */,
  {32'hc2079ad6, 32'h4159d5d2} /* (15, 3, 21) {real, imag} */,
  {32'hc17a30ca, 32'h40cbffd2} /* (15, 3, 20) {real, imag} */,
  {32'hc19d801a, 32'h3fa78440} /* (15, 3, 19) {real, imag} */,
  {32'h409214dd, 32'hc0bf6b24} /* (15, 3, 18) {real, imag} */,
  {32'h417b2da8, 32'h411da4b5} /* (15, 3, 17) {real, imag} */,
  {32'hc0525620, 32'h3fab8c48} /* (15, 3, 16) {real, imag} */,
  {32'h3edd5c70, 32'hc0c7c20a} /* (15, 3, 15) {real, imag} */,
  {32'hc0fceb15, 32'h40e76ec4} /* (15, 3, 14) {real, imag} */,
  {32'h40d47a7d, 32'h417d7d74} /* (15, 3, 13) {real, imag} */,
  {32'h415354f2, 32'hc16a51f9} /* (15, 3, 12) {real, imag} */,
  {32'hc118678a, 32'h412a47ac} /* (15, 3, 11) {real, imag} */,
  {32'hc1a9a7dc, 32'h4201e607} /* (15, 3, 10) {real, imag} */,
  {32'hc17e682c, 32'h3f581d14} /* (15, 3, 9) {real, imag} */,
  {32'h41ac7219, 32'hc13b9a24} /* (15, 3, 8) {real, imag} */,
  {32'h407df3fe, 32'hc178f0ee} /* (15, 3, 7) {real, imag} */,
  {32'h3fff3d80, 32'h41b06954} /* (15, 3, 6) {real, imag} */,
  {32'h42174626, 32'hbfb017a4} /* (15, 3, 5) {real, imag} */,
  {32'h411ddbaf, 32'h3fb86634} /* (15, 3, 4) {real, imag} */,
  {32'h40d2e673, 32'h41c620bd} /* (15, 3, 3) {real, imag} */,
  {32'hc0afcb38, 32'h407635e0} /* (15, 3, 2) {real, imag} */,
  {32'h4226a9ce, 32'h410c46a2} /* (15, 3, 1) {real, imag} */,
  {32'hc21f7192, 32'h418cf4ce} /* (15, 3, 0) {real, imag} */,
  {32'hc1c19774, 32'hc116898e} /* (15, 2, 31) {real, imag} */,
  {32'hc1fac8bd, 32'hc0cee664} /* (15, 2, 30) {real, imag} */,
  {32'h41fbd38c, 32'h41515bb0} /* (15, 2, 29) {real, imag} */,
  {32'hc0c7238c, 32'hc1b7b5b8} /* (15, 2, 28) {real, imag} */,
  {32'h422b0643, 32'h419b5330} /* (15, 2, 27) {real, imag} */,
  {32'h4108867c, 32'h426ecc00} /* (15, 2, 26) {real, imag} */,
  {32'hc0d1ad06, 32'h42024dd0} /* (15, 2, 25) {real, imag} */,
  {32'hc1248334, 32'hc1bf25cd} /* (15, 2, 24) {real, imag} */,
  {32'hc1bb208e, 32'hc1f5412e} /* (15, 2, 23) {real, imag} */,
  {32'h40f59383, 32'hc12c1528} /* (15, 2, 22) {real, imag} */,
  {32'hc006528a, 32'hc20d816a} /* (15, 2, 21) {real, imag} */,
  {32'hc1255b09, 32'h3ecbe330} /* (15, 2, 20) {real, imag} */,
  {32'h4080268a, 32'h416fbd82} /* (15, 2, 19) {real, imag} */,
  {32'h3fd0ad84, 32'hc090a903} /* (15, 2, 18) {real, imag} */,
  {32'h40c4d590, 32'hc144e766} /* (15, 2, 17) {real, imag} */,
  {32'h402c825e, 32'hc14f1a90} /* (15, 2, 16) {real, imag} */,
  {32'hc0a2ec58, 32'h405edf26} /* (15, 2, 15) {real, imag} */,
  {32'hc13e7a58, 32'hc08b4e3d} /* (15, 2, 14) {real, imag} */,
  {32'h3f125510, 32'h41726972} /* (15, 2, 13) {real, imag} */,
  {32'h4120863d, 32'hc117678e} /* (15, 2, 12) {real, imag} */,
  {32'h4002017a, 32'hc15684aa} /* (15, 2, 11) {real, imag} */,
  {32'hc0296eda, 32'h41044100} /* (15, 2, 10) {real, imag} */,
  {32'h400c63dc, 32'h413e0e84} /* (15, 2, 9) {real, imag} */,
  {32'hc15a19e4, 32'h410a58d2} /* (15, 2, 8) {real, imag} */,
  {32'hc0713374, 32'hbf1e9c60} /* (15, 2, 7) {real, imag} */,
  {32'hc0ea12f7, 32'hc268c436} /* (15, 2, 6) {real, imag} */,
  {32'h41b0c5f2, 32'hc16daa2c} /* (15, 2, 5) {real, imag} */,
  {32'hc18c4f24, 32'h3e988980} /* (15, 2, 4) {real, imag} */,
  {32'hc278218a, 32'h41bc7d52} /* (15, 2, 3) {real, imag} */,
  {32'h41e95acf, 32'hc1cac6a3} /* (15, 2, 2) {real, imag} */,
  {32'hc23d9c06, 32'hc21d0f36} /* (15, 2, 1) {real, imag} */,
  {32'h40fab447, 32'h428bf07e} /* (15, 2, 0) {real, imag} */,
  {32'h42469869, 32'h4138f75b} /* (15, 1, 31) {real, imag} */,
  {32'hc1c7d8e6, 32'h41ae1526} /* (15, 1, 30) {real, imag} */,
  {32'h41c5c113, 32'h41687822} /* (15, 1, 29) {real, imag} */,
  {32'h41396320, 32'hbf71c690} /* (15, 1, 28) {real, imag} */,
  {32'h413f8119, 32'hc018c212} /* (15, 1, 27) {real, imag} */,
  {32'hc1c54d22, 32'h4099319c} /* (15, 1, 26) {real, imag} */,
  {32'h415eb236, 32'h3e34de40} /* (15, 1, 25) {real, imag} */,
  {32'hc0cd060c, 32'h41d4617a} /* (15, 1, 24) {real, imag} */,
  {32'h42279d03, 32'h417cfac6} /* (15, 1, 23) {real, imag} */,
  {32'h402b904c, 32'h410f86ec} /* (15, 1, 22) {real, imag} */,
  {32'h3fb72558, 32'hc0dc11b3} /* (15, 1, 21) {real, imag} */,
  {32'h4169d503, 32'h41866192} /* (15, 1, 20) {real, imag} */,
  {32'hc0b5a940, 32'hc12ef524} /* (15, 1, 19) {real, imag} */,
  {32'h403fb664, 32'hc07d3670} /* (15, 1, 18) {real, imag} */,
  {32'h3f8e0e68, 32'hc0acbaac} /* (15, 1, 17) {real, imag} */,
  {32'hc1805b87, 32'hc17c0f00} /* (15, 1, 16) {real, imag} */,
  {32'h4086f5e6, 32'hc02bb5c1} /* (15, 1, 15) {real, imag} */,
  {32'h3ffbad18, 32'hc148bbf4} /* (15, 1, 14) {real, imag} */,
  {32'h40fe649c, 32'hc094c054} /* (15, 1, 13) {real, imag} */,
  {32'h411bad05, 32'hc179ac8b} /* (15, 1, 12) {real, imag} */,
  {32'h41281ce3, 32'h418a7be1} /* (15, 1, 11) {real, imag} */,
  {32'h41350b3b, 32'hc148b548} /* (15, 1, 10) {real, imag} */,
  {32'h41cc4d8a, 32'h41bbd139} /* (15, 1, 9) {real, imag} */,
  {32'hc18cdff5, 32'hc133a344} /* (15, 1, 8) {real, imag} */,
  {32'h414a795a, 32'h41cab5f8} /* (15, 1, 7) {real, imag} */,
  {32'h40681a8c, 32'h41458912} /* (15, 1, 6) {real, imag} */,
  {32'hc223e6eb, 32'h416ad068} /* (15, 1, 5) {real, imag} */,
  {32'h419febd8, 32'h41cbe7a6} /* (15, 1, 4) {real, imag} */,
  {32'hc1c8c8a9, 32'hc1629b04} /* (15, 1, 3) {real, imag} */,
  {32'hc24eddb5, 32'hc24de0f7} /* (15, 1, 2) {real, imag} */,
  {32'h42b1dec2, 32'h41a9d806} /* (15, 1, 1) {real, imag} */,
  {32'h4218a34a, 32'h41f1fbb6} /* (15, 1, 0) {real, imag} */,
  {32'h402ba7ec, 32'hc2784f4f} /* (15, 0, 31) {real, imag} */,
  {32'h415278b8, 32'h42043447} /* (15, 0, 30) {real, imag} */,
  {32'hc11b3b94, 32'hc242c5fa} /* (15, 0, 29) {real, imag} */,
  {32'hc22e96a2, 32'hc1c61ce7} /* (15, 0, 28) {real, imag} */,
  {32'hc181ce13, 32'h41ac20b8} /* (15, 0, 27) {real, imag} */,
  {32'hc12dd133, 32'hc1ae0c5a} /* (15, 0, 26) {real, imag} */,
  {32'h413672b8, 32'h40363898} /* (15, 0, 25) {real, imag} */,
  {32'hc1b4afaa, 32'hbe1e6180} /* (15, 0, 24) {real, imag} */,
  {32'h413c58a6, 32'h4133ab36} /* (15, 0, 23) {real, imag} */,
  {32'h41699969, 32'hc11d0ad1} /* (15, 0, 22) {real, imag} */,
  {32'hc0fa804b, 32'h409a8436} /* (15, 0, 21) {real, imag} */,
  {32'h402945ca, 32'hc0e5f484} /* (15, 0, 20) {real, imag} */,
  {32'hc14b7212, 32'h418bf8c4} /* (15, 0, 19) {real, imag} */,
  {32'h41c193ea, 32'hc07769d4} /* (15, 0, 18) {real, imag} */,
  {32'h4085df1e, 32'h4101f5a7} /* (15, 0, 17) {real, imag} */,
  {32'h4097d490, 32'h402b0c28} /* (15, 0, 16) {real, imag} */,
  {32'hbebd18a0, 32'hc0f2efce} /* (15, 0, 15) {real, imag} */,
  {32'hc12f1a24, 32'hc0bf3fa6} /* (15, 0, 14) {real, imag} */,
  {32'h418cf347, 32'h40ad30b2} /* (15, 0, 13) {real, imag} */,
  {32'h40edd4c3, 32'h40067698} /* (15, 0, 12) {real, imag} */,
  {32'hc12dae1e, 32'h4198d722} /* (15, 0, 11) {real, imag} */,
  {32'hc101c80b, 32'h412a8751} /* (15, 0, 10) {real, imag} */,
  {32'h3f7d4180, 32'h42008206} /* (15, 0, 9) {real, imag} */,
  {32'h4254212b, 32'hc1973f89} /* (15, 0, 8) {real, imag} */,
  {32'h41650b4a, 32'hc22e64d8} /* (15, 0, 7) {real, imag} */,
  {32'h41852530, 32'h4117dfcb} /* (15, 0, 6) {real, imag} */,
  {32'hc090f723, 32'hc0a5d2ca} /* (15, 0, 5) {real, imag} */,
  {32'hc2273da2, 32'hc107c44e} /* (15, 0, 4) {real, imag} */,
  {32'hc21e20df, 32'hc24bc56e} /* (15, 0, 3) {real, imag} */,
  {32'h3e9a2c00, 32'hbc936800} /* (15, 0, 2) {real, imag} */,
  {32'hc1d23cd4, 32'hc12b8af4} /* (15, 0, 1) {real, imag} */,
  {32'h419a3e68, 32'h41d0595f} /* (15, 0, 0) {real, imag} */,
  {32'hc30e95ab, 32'h420522dd} /* (14, 31, 31) {real, imag} */,
  {32'h41bb4add, 32'hc2a96aa2} /* (14, 31, 30) {real, imag} */,
  {32'h421fd2bf, 32'h4201ea4f} /* (14, 31, 29) {real, imag} */,
  {32'hc0a749d7, 32'h41a2f83b} /* (14, 31, 28) {real, imag} */,
  {32'hc20c9295, 32'hc16208da} /* (14, 31, 27) {real, imag} */,
  {32'hc144b968, 32'hc21c5833} /* (14, 31, 26) {real, imag} */,
  {32'hc266ef98, 32'hc18405fc} /* (14, 31, 25) {real, imag} */,
  {32'h400ff948, 32'hc21c323e} /* (14, 31, 24) {real, imag} */,
  {32'h414c9cd2, 32'hc18d4437} /* (14, 31, 23) {real, imag} */,
  {32'h41fb2bac, 32'h41507db4} /* (14, 31, 22) {real, imag} */,
  {32'h41bd18ea, 32'hc1da864b} /* (14, 31, 21) {real, imag} */,
  {32'h40cb3911, 32'h401f7393} /* (14, 31, 20) {real, imag} */,
  {32'h407ee090, 32'h40d23c04} /* (14, 31, 19) {real, imag} */,
  {32'h41325dd2, 32'h3e856500} /* (14, 31, 18) {real, imag} */,
  {32'hc12a8f6b, 32'hc0388022} /* (14, 31, 17) {real, imag} */,
  {32'h40570fa0, 32'hc164d9e0} /* (14, 31, 16) {real, imag} */,
  {32'hc10843e5, 32'h40b68db1} /* (14, 31, 15) {real, imag} */,
  {32'h40497be0, 32'hc0c06db8} /* (14, 31, 14) {real, imag} */,
  {32'hc1796ee0, 32'hc0011f80} /* (14, 31, 13) {real, imag} */,
  {32'hc0ba5bcf, 32'hbe106bb0} /* (14, 31, 12) {real, imag} */,
  {32'h42077aa7, 32'h3ec7bdc0} /* (14, 31, 11) {real, imag} */,
  {32'hc2114bcc, 32'hc15465a2} /* (14, 31, 10) {real, imag} */,
  {32'h412ca4aa, 32'hc1776daa} /* (14, 31, 9) {real, imag} */,
  {32'h4031ee88, 32'hc208800c} /* (14, 31, 8) {real, imag} */,
  {32'h41f64893, 32'hc14f0b26} /* (14, 31, 7) {real, imag} */,
  {32'hc11c2ff0, 32'h424b98c1} /* (14, 31, 6) {real, imag} */,
  {32'h41ea0312, 32'h41a7ae7d} /* (14, 31, 5) {real, imag} */,
  {32'hbf1613b8, 32'h41a501e5} /* (14, 31, 4) {real, imag} */,
  {32'h41987af8, 32'h3d96b200} /* (14, 31, 3) {real, imag} */,
  {32'h420e3cee, 32'hc1b9bae7} /* (14, 31, 2) {real, imag} */,
  {32'hc2cdac70, 32'h41b1966e} /* (14, 31, 1) {real, imag} */,
  {32'hc2999639, 32'hc06a7200} /* (14, 31, 0) {real, imag} */,
  {32'h430be65d, 32'hc11f0f42} /* (14, 30, 31) {real, imag} */,
  {32'hc2ae5a27, 32'h41887442} /* (14, 30, 30) {real, imag} */,
  {32'hc09bc238, 32'h417f7408} /* (14, 30, 29) {real, imag} */,
  {32'hc02502b8, 32'h4227b6df} /* (14, 30, 28) {real, imag} */,
  {32'hc212a630, 32'h420dfb27} /* (14, 30, 27) {real, imag} */,
  {32'hc1aba52f, 32'hc03b8598} /* (14, 30, 26) {real, imag} */,
  {32'h419d59b0, 32'h41b2a24c} /* (14, 30, 25) {real, imag} */,
  {32'hc1ffbb01, 32'hc12fbf84} /* (14, 30, 24) {real, imag} */,
  {32'h3f0bbc40, 32'hc16eb8b1} /* (14, 30, 23) {real, imag} */,
  {32'h41f9be04, 32'hc093ba2c} /* (14, 30, 22) {real, imag} */,
  {32'hc0468150, 32'h41223103} /* (14, 30, 21) {real, imag} */,
  {32'hc046e078, 32'h40338b42} /* (14, 30, 20) {real, imag} */,
  {32'hc1ca3012, 32'h408f08d2} /* (14, 30, 19) {real, imag} */,
  {32'h40c0de2c, 32'hbfd68c48} /* (14, 30, 18) {real, imag} */,
  {32'hc005ab60, 32'hc027fe14} /* (14, 30, 17) {real, imag} */,
  {32'hc12db39c, 32'hc099773b} /* (14, 30, 16) {real, imag} */,
  {32'hc158edf8, 32'h40bbe112} /* (14, 30, 15) {real, imag} */,
  {32'hbeb9dfc0, 32'h417e7f0f} /* (14, 30, 14) {real, imag} */,
  {32'hbf73a5b0, 32'h41064c2b} /* (14, 30, 13) {real, imag} */,
  {32'h419a9ef7, 32'hc0ed7035} /* (14, 30, 12) {real, imag} */,
  {32'hc15aa4fc, 32'h40c5688a} /* (14, 30, 11) {real, imag} */,
  {32'h41b43420, 32'hc1d056da} /* (14, 30, 10) {real, imag} */,
  {32'h42035dac, 32'hc0ea6afe} /* (14, 30, 9) {real, imag} */,
  {32'hc1c3dd0f, 32'h400e3452} /* (14, 30, 8) {real, imag} */,
  {32'hc195720a, 32'h4172cc07} /* (14, 30, 7) {real, imag} */,
  {32'h415cfd92, 32'h41004900} /* (14, 30, 6) {real, imag} */,
  {32'hc1d06310, 32'h412be5f9} /* (14, 30, 5) {real, imag} */,
  {32'h4244916a, 32'h41c13c2a} /* (14, 30, 4) {real, imag} */,
  {32'h4242dbff, 32'hc1cbcf74} /* (14, 30, 3) {real, imag} */,
  {32'hc2b43ad5, 32'h40e68e0e} /* (14, 30, 2) {real, imag} */,
  {32'h4307faef, 32'hc255b956} /* (14, 30, 1) {real, imag} */,
  {32'h427fa7d3, 32'h412bedb0} /* (14, 30, 0) {real, imag} */,
  {32'hc271a031, 32'hbff1cbd0} /* (14, 29, 31) {real, imag} */,
  {32'h41c57256, 32'hc1c3e5f2} /* (14, 29, 30) {real, imag} */,
  {32'h4141edec, 32'hc269c802} /* (14, 29, 29) {real, imag} */,
  {32'h3eb16180, 32'hc19ab2b6} /* (14, 29, 28) {real, imag} */,
  {32'hc1c56c85, 32'h420f4e24} /* (14, 29, 27) {real, imag} */,
  {32'hc05552c0, 32'hc07b0ade} /* (14, 29, 26) {real, imag} */,
  {32'h4258da0a, 32'h41f1ef80} /* (14, 29, 25) {real, imag} */,
  {32'hc2265c5a, 32'hc11f28f2} /* (14, 29, 24) {real, imag} */,
  {32'hc16b84bd, 32'hc1c52425} /* (14, 29, 23) {real, imag} */,
  {32'h41646724, 32'h3fd0a8d0} /* (14, 29, 22) {real, imag} */,
  {32'hbfff37d6, 32'h4176fb82} /* (14, 29, 21) {real, imag} */,
  {32'hc1a56816, 32'h4128c500} /* (14, 29, 20) {real, imag} */,
  {32'h417f9007, 32'h4090a470} /* (14, 29, 19) {real, imag} */,
  {32'h404c31ac, 32'hc095b393} /* (14, 29, 18) {real, imag} */,
  {32'h4193def8, 32'hc1872b74} /* (14, 29, 17) {real, imag} */,
  {32'h4080a2b8, 32'h40e1b858} /* (14, 29, 16) {real, imag} */,
  {32'hc1042cdb, 32'h412a5a24} /* (14, 29, 15) {real, imag} */,
  {32'h419e7c02, 32'hbe8c6410} /* (14, 29, 14) {real, imag} */,
  {32'h40151b4c, 32'hc0dca010} /* (14, 29, 13) {real, imag} */,
  {32'hc057f45c, 32'hc0f47869} /* (14, 29, 12) {real, imag} */,
  {32'h4095d7d4, 32'h3f67b8c8} /* (14, 29, 11) {real, imag} */,
  {32'hc1ab41fe, 32'h41b6465b} /* (14, 29, 10) {real, imag} */,
  {32'hc0f1fc3e, 32'h4110b296} /* (14, 29, 9) {real, imag} */,
  {32'h40ab3e94, 32'hc18e6d93} /* (14, 29, 8) {real, imag} */,
  {32'hc1769c0a, 32'h42491928} /* (14, 29, 7) {real, imag} */,
  {32'h427769a4, 32'h4015170e} /* (14, 29, 6) {real, imag} */,
  {32'h40ef743c, 32'h417271f2} /* (14, 29, 5) {real, imag} */,
  {32'hc206fe83, 32'h3fb7af00} /* (14, 29, 4) {real, imag} */,
  {32'hc25e1f45, 32'hc2388236} /* (14, 29, 3) {real, imag} */,
  {32'h41d63ba2, 32'hc057d95c} /* (14, 29, 2) {real, imag} */,
  {32'hc10e8bfc, 32'h41e2e9c9} /* (14, 29, 1) {real, imag} */,
  {32'hc209587a, 32'h4211a707} /* (14, 29, 0) {real, imag} */,
  {32'hc213a276, 32'h42b85cb2} /* (14, 28, 31) {real, imag} */,
  {32'h4281c2ea, 32'h4207011d} /* (14, 28, 30) {real, imag} */,
  {32'h424fb1cf, 32'h41474808} /* (14, 28, 29) {real, imag} */,
  {32'h421ac65e, 32'h403a1190} /* (14, 28, 28) {real, imag} */,
  {32'hc03a53d0, 32'hc206d083} /* (14, 28, 27) {real, imag} */,
  {32'h4167afeb, 32'hc20ad95c} /* (14, 28, 26) {real, imag} */,
  {32'hc2586fda, 32'h41d77372} /* (14, 28, 25) {real, imag} */,
  {32'h41bbcc6b, 32'hc28cb7da} /* (14, 28, 24) {real, imag} */,
  {32'hc0a3a688, 32'h40e34a1f} /* (14, 28, 23) {real, imag} */,
  {32'h3f97cb4e, 32'hc1ef710e} /* (14, 28, 22) {real, imag} */,
  {32'hc190679a, 32'h3fe4b910} /* (14, 28, 21) {real, imag} */,
  {32'h40f815b6, 32'hbf91cc58} /* (14, 28, 20) {real, imag} */,
  {32'hc193a2cc, 32'h40b05764} /* (14, 28, 19) {real, imag} */,
  {32'hc0e650f0, 32'h3fd2b890} /* (14, 28, 18) {real, imag} */,
  {32'h413d4744, 32'h406445b0} /* (14, 28, 17) {real, imag} */,
  {32'hc093bc7c, 32'h3ff1e690} /* (14, 28, 16) {real, imag} */,
  {32'h3f772188, 32'h40a408b8} /* (14, 28, 15) {real, imag} */,
  {32'hc1921c2a, 32'hc11b838a} /* (14, 28, 14) {real, imag} */,
  {32'hc0853cb0, 32'h3f5be2a0} /* (14, 28, 13) {real, imag} */,
  {32'hc11d96e9, 32'hc17b86c3} /* (14, 28, 12) {real, imag} */,
  {32'hc11c4873, 32'h41c1b50a} /* (14, 28, 11) {real, imag} */,
  {32'hbf1ccd14, 32'h40ab7a96} /* (14, 28, 10) {real, imag} */,
  {32'hc20485ae, 32'h3fdd6a1c} /* (14, 28, 9) {real, imag} */,
  {32'h41fac93d, 32'hc01e2ec0} /* (14, 28, 8) {real, imag} */,
  {32'hc196c4a5, 32'hc177e828} /* (14, 28, 7) {real, imag} */,
  {32'hc07fc7d4, 32'h407d8f9c} /* (14, 28, 6) {real, imag} */,
  {32'h4285d6d4, 32'hc1ad325a} /* (14, 28, 5) {real, imag} */,
  {32'hc28e99af, 32'hc2627a87} /* (14, 28, 4) {real, imag} */,
  {32'h425caa11, 32'hc1ee2600} /* (14, 28, 3) {real, imag} */,
  {32'hbe335800, 32'hc186dffc} /* (14, 28, 2) {real, imag} */,
  {32'hc23bc6ca, 32'h4255ceac} /* (14, 28, 1) {real, imag} */,
  {32'hc1d766b5, 32'hc17c154a} /* (14, 28, 0) {real, imag} */,
  {32'h41160314, 32'h3fd112e0} /* (14, 27, 31) {real, imag} */,
  {32'hc1057eee, 32'h42b26d8a} /* (14, 27, 30) {real, imag} */,
  {32'hc1d82b3b, 32'h4215bc71} /* (14, 27, 29) {real, imag} */,
  {32'h40a59f98, 32'h409a0208} /* (14, 27, 28) {real, imag} */,
  {32'hc1a866b2, 32'h41757dfc} /* (14, 27, 27) {real, imag} */,
  {32'h41c5bfb8, 32'hc19d0f4b} /* (14, 27, 26) {real, imag} */,
  {32'hc0be6a8b, 32'hc1cbba70} /* (14, 27, 25) {real, imag} */,
  {32'hbeaf7f60, 32'h40a474ac} /* (14, 27, 24) {real, imag} */,
  {32'hc223866e, 32'hc18f772a} /* (14, 27, 23) {real, imag} */,
  {32'hc0f45f80, 32'hc035227c} /* (14, 27, 22) {real, imag} */,
  {32'hc1ad0f4e, 32'h41cf4c48} /* (14, 27, 21) {real, imag} */,
  {32'hc19881da, 32'hc18ae662} /* (14, 27, 20) {real, imag} */,
  {32'h408e286a, 32'hc07f65bc} /* (14, 27, 19) {real, imag} */,
  {32'h3e8a4750, 32'h40f15750} /* (14, 27, 18) {real, imag} */,
  {32'h4075b388, 32'hc03a0784} /* (14, 27, 17) {real, imag} */,
  {32'h40baad40, 32'hbfe1cec0} /* (14, 27, 16) {real, imag} */,
  {32'h416bdb82, 32'hc18fbe64} /* (14, 27, 15) {real, imag} */,
  {32'hc064941a, 32'h405e8150} /* (14, 27, 14) {real, imag} */,
  {32'hc17db195, 32'hc109293f} /* (14, 27, 13) {real, imag} */,
  {32'hc19ab3a6, 32'hc16ceb48} /* (14, 27, 12) {real, imag} */,
  {32'h404cfe44, 32'hc1152b4c} /* (14, 27, 11) {real, imag} */,
  {32'h41b15646, 32'hc0c1935a} /* (14, 27, 10) {real, imag} */,
  {32'hbfdf8490, 32'h411c2381} /* (14, 27, 9) {real, imag} */,
  {32'h418d9e40, 32'hc1daa027} /* (14, 27, 8) {real, imag} */,
  {32'h419fde41, 32'hc04bd294} /* (14, 27, 7) {real, imag} */,
  {32'hc0b7f7b8, 32'h41cef181} /* (14, 27, 6) {real, imag} */,
  {32'hc1b74686, 32'h423407ac} /* (14, 27, 5) {real, imag} */,
  {32'h4258e4ff, 32'hc17048b0} /* (14, 27, 4) {real, imag} */,
  {32'h4152ad22, 32'h4046bc50} /* (14, 27, 3) {real, imag} */,
  {32'hc1e7866f, 32'h40c2ed40} /* (14, 27, 2) {real, imag} */,
  {32'h42616efb, 32'hc255f649} /* (14, 27, 1) {real, imag} */,
  {32'h42121a10, 32'h4224b1ac} /* (14, 27, 0) {real, imag} */,
  {32'h418d7114, 32'h3f78cf20} /* (14, 26, 31) {real, imag} */,
  {32'h41b7ddb0, 32'h41d6e740} /* (14, 26, 30) {real, imag} */,
  {32'hc19ed956, 32'hc2117e6d} /* (14, 26, 29) {real, imag} */,
  {32'h414c7701, 32'h410fcc85} /* (14, 26, 28) {real, imag} */,
  {32'hc037b704, 32'h40ac2ed8} /* (14, 26, 27) {real, imag} */,
  {32'hc226ad94, 32'hc06c4493} /* (14, 26, 26) {real, imag} */,
  {32'h4160210e, 32'hc1d9f358} /* (14, 26, 25) {real, imag} */,
  {32'h4145aed0, 32'h40b71b16} /* (14, 26, 24) {real, imag} */,
  {32'hc09e4e55, 32'h41469bd9} /* (14, 26, 23) {real, imag} */,
  {32'h41bb45f0, 32'hc16e66f3} /* (14, 26, 22) {real, imag} */,
  {32'h41454b31, 32'hc09aadfc} /* (14, 26, 21) {real, imag} */,
  {32'hc0ca721c, 32'h40ba0e20} /* (14, 26, 20) {real, imag} */,
  {32'hbf6a3a30, 32'h404e1b9c} /* (14, 26, 19) {real, imag} */,
  {32'hc11f2b7a, 32'hc18b1126} /* (14, 26, 18) {real, imag} */,
  {32'hbf97fafe, 32'hc0923c3d} /* (14, 26, 17) {real, imag} */,
  {32'h415564f4, 32'h40d5ff2c} /* (14, 26, 16) {real, imag} */,
  {32'h40a4fb2e, 32'hc0f5448b} /* (14, 26, 15) {real, imag} */,
  {32'hc0b72e80, 32'h40bf4f92} /* (14, 26, 14) {real, imag} */,
  {32'hc0eb728a, 32'hbf34594e} /* (14, 26, 13) {real, imag} */,
  {32'h408a11a2, 32'hc0d8cc40} /* (14, 26, 12) {real, imag} */,
  {32'hc0b5452e, 32'hc10d647c} /* (14, 26, 11) {real, imag} */,
  {32'h41786304, 32'h410534fd} /* (14, 26, 10) {real, imag} */,
  {32'hc06bd782, 32'hc146ea97} /* (14, 26, 9) {real, imag} */,
  {32'h41597f08, 32'hc1068f7f} /* (14, 26, 8) {real, imag} */,
  {32'h41104bf6, 32'h40247fe4} /* (14, 26, 7) {real, imag} */,
  {32'hc0ff7cbc, 32'hc06df7df} /* (14, 26, 6) {real, imag} */,
  {32'h41c1e024, 32'h3f8e31ae} /* (14, 26, 5) {real, imag} */,
  {32'hc1a5b53c, 32'hbed9c3e0} /* (14, 26, 4) {real, imag} */,
  {32'h410c3fc3, 32'h4222207b} /* (14, 26, 3) {real, imag} */,
  {32'hc209cb54, 32'h3fd2a058} /* (14, 26, 2) {real, imag} */,
  {32'h40cc86d2, 32'h41d12699} /* (14, 26, 1) {real, imag} */,
  {32'hc21de751, 32'h41f81637} /* (14, 26, 0) {real, imag} */,
  {32'hc2509d2e, 32'h41e54aa3} /* (14, 25, 31) {real, imag} */,
  {32'h41968db7, 32'h420826a8} /* (14, 25, 30) {real, imag} */,
  {32'h4193202a, 32'h41ce4c56} /* (14, 25, 29) {real, imag} */,
  {32'h40ac97d0, 32'hc0a620f9} /* (14, 25, 28) {real, imag} */,
  {32'h41f41a74, 32'hc1fbe372} /* (14, 25, 27) {real, imag} */,
  {32'hc1a3b02d, 32'h400d24f8} /* (14, 25, 26) {real, imag} */,
  {32'h40e2dff4, 32'h412ef672} /* (14, 25, 25) {real, imag} */,
  {32'hc0f1f903, 32'hc07ff880} /* (14, 25, 24) {real, imag} */,
  {32'hc089d17f, 32'h41849e6c} /* (14, 25, 23) {real, imag} */,
  {32'h41a375d8, 32'hc0524206} /* (14, 25, 22) {real, imag} */,
  {32'h3e69d440, 32'h406c8cac} /* (14, 25, 21) {real, imag} */,
  {32'hc093a225, 32'hbf083b00} /* (14, 25, 20) {real, imag} */,
  {32'h3e408d60, 32'hc0b50bed} /* (14, 25, 19) {real, imag} */,
  {32'hc0311e40, 32'h41068d54} /* (14, 25, 18) {real, imag} */,
  {32'hc0ddb868, 32'hc0fe704d} /* (14, 25, 17) {real, imag} */,
  {32'h40151c82, 32'h40520b96} /* (14, 25, 16) {real, imag} */,
  {32'hc11b90cc, 32'h402659aa} /* (14, 25, 15) {real, imag} */,
  {32'hbf8e98a0, 32'h400bc302} /* (14, 25, 14) {real, imag} */,
  {32'h416d3fb4, 32'h40b8c0c9} /* (14, 25, 13) {real, imag} */,
  {32'h400cf592, 32'h3dd80180} /* (14, 25, 12) {real, imag} */,
  {32'h4193cf9c, 32'hbfed3f88} /* (14, 25, 11) {real, imag} */,
  {32'h40942224, 32'h4019e462} /* (14, 25, 10) {real, imag} */,
  {32'h3fcdb4e4, 32'h4172dab4} /* (14, 25, 9) {real, imag} */,
  {32'hc027dcda, 32'h4091f28e} /* (14, 25, 8) {real, imag} */,
  {32'hc20bd4e4, 32'hc12f40b6} /* (14, 25, 7) {real, imag} */,
  {32'hc0aa2a58, 32'hc1af5f15} /* (14, 25, 6) {real, imag} */,
  {32'hc13f30c0, 32'h41df0030} /* (14, 25, 5) {real, imag} */,
  {32'h4041a97c, 32'hc193bee0} /* (14, 25, 4) {real, imag} */,
  {32'hc20a65a3, 32'h4168a8c4} /* (14, 25, 3) {real, imag} */,
  {32'h4254611c, 32'h424367b8} /* (14, 25, 2) {real, imag} */,
  {32'h41c14228, 32'h4158be4e} /* (14, 25, 1) {real, imag} */,
  {32'hc157d4a8, 32'h4192183b} /* (14, 25, 0) {real, imag} */,
  {32'h41bfd57d, 32'hc1df244b} /* (14, 24, 31) {real, imag} */,
  {32'hc2335068, 32'h4128696e} /* (14, 24, 30) {real, imag} */,
  {32'hc1f613f6, 32'h40c80ab2} /* (14, 24, 29) {real, imag} */,
  {32'hc17fa235, 32'hc190a510} /* (14, 24, 28) {real, imag} */,
  {32'h41cbefe5, 32'hc1c713e4} /* (14, 24, 27) {real, imag} */,
  {32'h40372ab0, 32'hc20d1bb5} /* (14, 24, 26) {real, imag} */,
  {32'h417907cc, 32'hc17a449a} /* (14, 24, 25) {real, imag} */,
  {32'h404bd748, 32'hc213306c} /* (14, 24, 24) {real, imag} */,
  {32'h40ee5b1d, 32'h4119457a} /* (14, 24, 23) {real, imag} */,
  {32'hc16d7fd4, 32'h40a9b8ec} /* (14, 24, 22) {real, imag} */,
  {32'h3fc6c6a4, 32'h40eb5b82} /* (14, 24, 21) {real, imag} */,
  {32'hc0e5beba, 32'h40fbfbf2} /* (14, 24, 20) {real, imag} */,
  {32'hc1431fd4, 32'h411f004c} /* (14, 24, 19) {real, imag} */,
  {32'h3fa33964, 32'h40800e7b} /* (14, 24, 18) {real, imag} */,
  {32'hc032e4d6, 32'hc080f8fd} /* (14, 24, 17) {real, imag} */,
  {32'h40b75aad, 32'h3e9a1900} /* (14, 24, 16) {real, imag} */,
  {32'hc0694c26, 32'h40c9c27d} /* (14, 24, 15) {real, imag} */,
  {32'hc074de0a, 32'hc100c900} /* (14, 24, 14) {real, imag} */,
  {32'h41aad25a, 32'hc11a8a7c} /* (14, 24, 13) {real, imag} */,
  {32'hbf090e50, 32'h41a342e2} /* (14, 24, 12) {real, imag} */,
  {32'h4071b7b2, 32'h40f545fe} /* (14, 24, 11) {real, imag} */,
  {32'h40bd2271, 32'h4162a5f8} /* (14, 24, 10) {real, imag} */,
  {32'h40a75eed, 32'h4145e574} /* (14, 24, 9) {real, imag} */,
  {32'hc1dc5735, 32'h412e7d9e} /* (14, 24, 8) {real, imag} */,
  {32'hc11ea04c, 32'h40d378b8} /* (14, 24, 7) {real, imag} */,
  {32'hc113b029, 32'hc121492b} /* (14, 24, 6) {real, imag} */,
  {32'hc1bf4843, 32'h40eac990} /* (14, 24, 5) {real, imag} */,
  {32'h412e3e17, 32'h420a3d1f} /* (14, 24, 4) {real, imag} */,
  {32'h411db214, 32'hc021bb2d} /* (14, 24, 3) {real, imag} */,
  {32'hc1930a9d, 32'hc1770254} /* (14, 24, 2) {real, imag} */,
  {32'h40c34254, 32'hc1d999bd} /* (14, 24, 1) {real, imag} */,
  {32'h41209ff8, 32'hbfcb71f8} /* (14, 24, 0) {real, imag} */,
  {32'hc16c1cf4, 32'hc01e6984} /* (14, 23, 31) {real, imag} */,
  {32'hc1dd7684, 32'hc140a068} /* (14, 23, 30) {real, imag} */,
  {32'h41a2634c, 32'h40fdecf0} /* (14, 23, 29) {real, imag} */,
  {32'hc22a1862, 32'hc1c95798} /* (14, 23, 28) {real, imag} */,
  {32'hc1c3c124, 32'hbf3775b0} /* (14, 23, 27) {real, imag} */,
  {32'h41cbdfc2, 32'h4129ad27} /* (14, 23, 26) {real, imag} */,
  {32'h3fe917f0, 32'h41311f08} /* (14, 23, 25) {real, imag} */,
  {32'h4116728e, 32'h40dd870c} /* (14, 23, 24) {real, imag} */,
  {32'hc0b1d39f, 32'hc117eaf6} /* (14, 23, 23) {real, imag} */,
  {32'h40e41b90, 32'hc1b8ab6c} /* (14, 23, 22) {real, imag} */,
  {32'hc097f2ee, 32'hc0fa3fa4} /* (14, 23, 21) {real, imag} */,
  {32'hc07f9116, 32'hc058577e} /* (14, 23, 20) {real, imag} */,
  {32'h3d39e600, 32'hbfb3efd4} /* (14, 23, 19) {real, imag} */,
  {32'hbfcbc74c, 32'h3f9991b4} /* (14, 23, 18) {real, imag} */,
  {32'h402a0fba, 32'h3f806d96} /* (14, 23, 17) {real, imag} */,
  {32'hbfe08a30, 32'hc0f60c40} /* (14, 23, 16) {real, imag} */,
  {32'h40ab7f9b, 32'hc09faea6} /* (14, 23, 15) {real, imag} */,
  {32'h40eb82c9, 32'hc00e8456} /* (14, 23, 14) {real, imag} */,
  {32'h40abf908, 32'hc0211bae} /* (14, 23, 13) {real, imag} */,
  {32'h3f5695e8, 32'hc09f7007} /* (14, 23, 12) {real, imag} */,
  {32'hc0e11d6a, 32'h3f58b120} /* (14, 23, 11) {real, imag} */,
  {32'hc0ab68c0, 32'hc0927a1c} /* (14, 23, 10) {real, imag} */,
  {32'hc0704a02, 32'h41023f92} /* (14, 23, 9) {real, imag} */,
  {32'h3faf6108, 32'h41c484c3} /* (14, 23, 8) {real, imag} */,
  {32'h41a890e7, 32'hc11967e8} /* (14, 23, 7) {real, imag} */,
  {32'h412914dd, 32'h40a76f16} /* (14, 23, 6) {real, imag} */,
  {32'h41cd4a2c, 32'h41114c99} /* (14, 23, 5) {real, imag} */,
  {32'h41d9bfdd, 32'h40797614} /* (14, 23, 4) {real, imag} */,
  {32'hc1fac1f0, 32'h416d3ee8} /* (14, 23, 3) {real, imag} */,
  {32'hc09d2ce0, 32'h422a9dfd} /* (14, 23, 2) {real, imag} */,
  {32'h41612040, 32'h4145c7d1} /* (14, 23, 1) {real, imag} */,
  {32'hc13f021d, 32'h41c470fe} /* (14, 23, 0) {real, imag} */,
  {32'hc072f1c0, 32'hc05880b6} /* (14, 22, 31) {real, imag} */,
  {32'hc06894d0, 32'hc06bcfe8} /* (14, 22, 30) {real, imag} */,
  {32'hbf83cfbc, 32'hc1c51cd2} /* (14, 22, 29) {real, imag} */,
  {32'hc15ca608, 32'h41661eb1} /* (14, 22, 28) {real, imag} */,
  {32'h4199d796, 32'h40860c9f} /* (14, 22, 27) {real, imag} */,
  {32'h4127c34a, 32'h41a5c21c} /* (14, 22, 26) {real, imag} */,
  {32'hc1785757, 32'h41263ee2} /* (14, 22, 25) {real, imag} */,
  {32'h40a12b80, 32'h40493116} /* (14, 22, 24) {real, imag} */,
  {32'h40989b9f, 32'h407436ea} /* (14, 22, 23) {real, imag} */,
  {32'h40c758fb, 32'h409e62dd} /* (14, 22, 22) {real, imag} */,
  {32'h40ad476d, 32'h41b171ae} /* (14, 22, 21) {real, imag} */,
  {32'h40933250, 32'h40b09346} /* (14, 22, 20) {real, imag} */,
  {32'h4122601c, 32'hbd350b00} /* (14, 22, 19) {real, imag} */,
  {32'h3e8c14f0, 32'hc021402d} /* (14, 22, 18) {real, imag} */,
  {32'hbe76e960, 32'h404bcb7e} /* (14, 22, 17) {real, imag} */,
  {32'h40b54c6a, 32'h3f0e2ef0} /* (14, 22, 16) {real, imag} */,
  {32'h40310f1a, 32'hc07d0ace} /* (14, 22, 15) {real, imag} */,
  {32'h40894ab7, 32'hc017cd13} /* (14, 22, 14) {real, imag} */,
  {32'h3f6eb638, 32'hc02709a0} /* (14, 22, 13) {real, imag} */,
  {32'h414e1834, 32'h3fb2ace0} /* (14, 22, 12) {real, imag} */,
  {32'h410a3540, 32'hc0b9bdb8} /* (14, 22, 11) {real, imag} */,
  {32'hc153c5c2, 32'h40dd5bb7} /* (14, 22, 10) {real, imag} */,
  {32'h41034b5c, 32'hbfd12ee9} /* (14, 22, 9) {real, imag} */,
  {32'hc180bf2b, 32'h3f48ec70} /* (14, 22, 8) {real, imag} */,
  {32'h413c67cd, 32'hc12c2e0c} /* (14, 22, 7) {real, imag} */,
  {32'h3fb20294, 32'hc11e2885} /* (14, 22, 6) {real, imag} */,
  {32'hc1ccd3d6, 32'h4042bfb6} /* (14, 22, 5) {real, imag} */,
  {32'hc21f6271, 32'h40cf53be} /* (14, 22, 4) {real, imag} */,
  {32'hc0b87d7f, 32'h4017b160} /* (14, 22, 3) {real, imag} */,
  {32'h41d72d9c, 32'hc1967a33} /* (14, 22, 2) {real, imag} */,
  {32'h41fd6594, 32'h4134e454} /* (14, 22, 1) {real, imag} */,
  {32'h4194af34, 32'h41882a32} /* (14, 22, 0) {real, imag} */,
  {32'h41be58c3, 32'h41bd8457} /* (14, 21, 31) {real, imag} */,
  {32'hc115f363, 32'hc00a9e9c} /* (14, 21, 30) {real, imag} */,
  {32'h41e531fe, 32'hc1ba20b2} /* (14, 21, 29) {real, imag} */,
  {32'h41a0ff57, 32'h41ca945e} /* (14, 21, 28) {real, imag} */,
  {32'h41e78e9c, 32'hc19f58dc} /* (14, 21, 27) {real, imag} */,
  {32'h40f70e47, 32'h3fcb4bd0} /* (14, 21, 26) {real, imag} */,
  {32'h40586b47, 32'hc13ea96b} /* (14, 21, 25) {real, imag} */,
  {32'h41aca665, 32'hc04a3aca} /* (14, 21, 24) {real, imag} */,
  {32'hc04f884a, 32'h4104e2b3} /* (14, 21, 23) {real, imag} */,
  {32'hc15032ca, 32'h414f8878} /* (14, 21, 22) {real, imag} */,
  {32'h41139e9e, 32'hc0358cda} /* (14, 21, 21) {real, imag} */,
  {32'hbfcfff1a, 32'h3e0fa9e0} /* (14, 21, 20) {real, imag} */,
  {32'h4016d4ad, 32'hc0da063e} /* (14, 21, 19) {real, imag} */,
  {32'hc09663b8, 32'h41070a40} /* (14, 21, 18) {real, imag} */,
  {32'h40a6a79a, 32'hc00febae} /* (14, 21, 17) {real, imag} */,
  {32'h3ebda570, 32'hc08c3baf} /* (14, 21, 16) {real, imag} */,
  {32'hc0cb1f52, 32'h3fda5ea4} /* (14, 21, 15) {real, imag} */,
  {32'h40ee94cc, 32'hc07f8daa} /* (14, 21, 14) {real, imag} */,
  {32'hc0b53b82, 32'hc14513e5} /* (14, 21, 13) {real, imag} */,
  {32'h40d4b522, 32'h40e65099} /* (14, 21, 12) {real, imag} */,
  {32'hc0c5f8fb, 32'h3f5b54b8} /* (14, 21, 11) {real, imag} */,
  {32'h41896121, 32'hc0a5a77d} /* (14, 21, 10) {real, imag} */,
  {32'h3f33aa82, 32'hbf5b9c6c} /* (14, 21, 9) {real, imag} */,
  {32'hbe348780, 32'hc14c2284} /* (14, 21, 8) {real, imag} */,
  {32'hc028078d, 32'h40b723fa} /* (14, 21, 7) {real, imag} */,
  {32'h3fba97dc, 32'hc1358ad9} /* (14, 21, 6) {real, imag} */,
  {32'hc1868aa2, 32'hc035935c} /* (14, 21, 5) {real, imag} */,
  {32'h3d367600, 32'h41832b68} /* (14, 21, 4) {real, imag} */,
  {32'hc147f9b9, 32'h4032514c} /* (14, 21, 3) {real, imag} */,
  {32'h4059a0ac, 32'hc1b744fa} /* (14, 21, 2) {real, imag} */,
  {32'h4193774f, 32'hc104321a} /* (14, 21, 1) {real, imag} */,
  {32'hc0b2027d, 32'hc16d2690} /* (14, 21, 0) {real, imag} */,
  {32'hc10d5e21, 32'hc0b34e40} /* (14, 20, 31) {real, imag} */,
  {32'h41a3676e, 32'hc117628c} /* (14, 20, 30) {real, imag} */,
  {32'hc16a8842, 32'hc1236584} /* (14, 20, 29) {real, imag} */,
  {32'h40686cd0, 32'hc11205b8} /* (14, 20, 28) {real, imag} */,
  {32'hc1e09401, 32'h41818b0a} /* (14, 20, 27) {real, imag} */,
  {32'hc0d39302, 32'h40583885} /* (14, 20, 26) {real, imag} */,
  {32'hc14024dc, 32'h4038b33c} /* (14, 20, 25) {real, imag} */,
  {32'hc0e86827, 32'h40d1ed48} /* (14, 20, 24) {real, imag} */,
  {32'hc0b0d6c1, 32'hbf656b80} /* (14, 20, 23) {real, imag} */,
  {32'h406d5ef2, 32'h40ca9e88} /* (14, 20, 22) {real, imag} */,
  {32'hc19a1712, 32'hc0434f76} /* (14, 20, 21) {real, imag} */,
  {32'h408d7e94, 32'hc06df75e} /* (14, 20, 20) {real, imag} */,
  {32'h3fd8eccc, 32'hbf86fa78} /* (14, 20, 19) {real, imag} */,
  {32'hc06f4c7a, 32'hbff7d8c4} /* (14, 20, 18) {real, imag} */,
  {32'h40d4ee0c, 32'hbfb772a4} /* (14, 20, 17) {real, imag} */,
  {32'hbde7a400, 32'hc00d9d59} /* (14, 20, 16) {real, imag} */,
  {32'hbf5ecc04, 32'hbe805002} /* (14, 20, 15) {real, imag} */,
  {32'h3f070f6a, 32'h408ef018} /* (14, 20, 14) {real, imag} */,
  {32'h3fc1cd0c, 32'h3f0c8d50} /* (14, 20, 13) {real, imag} */,
  {32'h40940c28, 32'hc05f9ec6} /* (14, 20, 12) {real, imag} */,
  {32'h3ff03280, 32'h410c85c2} /* (14, 20, 11) {real, imag} */,
  {32'hc146f6b2, 32'h414413a8} /* (14, 20, 10) {real, imag} */,
  {32'h40ce73d9, 32'hc11c8212} /* (14, 20, 9) {real, imag} */,
  {32'h4150e024, 32'h3df9eba0} /* (14, 20, 8) {real, imag} */,
  {32'h4168a3bc, 32'h41748101} /* (14, 20, 7) {real, imag} */,
  {32'h3f984122, 32'h3f94edee} /* (14, 20, 6) {real, imag} */,
  {32'hc1286c3a, 32'h418edf7c} /* (14, 20, 5) {real, imag} */,
  {32'hc1af53fd, 32'h4143d64e} /* (14, 20, 4) {real, imag} */,
  {32'h41564e1e, 32'hc00be748} /* (14, 20, 3) {real, imag} */,
  {32'hc15d39ad, 32'h40b90418} /* (14, 20, 2) {real, imag} */,
  {32'h40d12cbe, 32'hc10fa7b2} /* (14, 20, 1) {real, imag} */,
  {32'h4159a941, 32'h3f8f82ce} /* (14, 20, 0) {real, imag} */,
  {32'h40e9c486, 32'h41223e83} /* (14, 19, 31) {real, imag} */,
  {32'hc18244c6, 32'hbe77044c} /* (14, 19, 30) {real, imag} */,
  {32'hc163d9a4, 32'hc17dd720} /* (14, 19, 29) {real, imag} */,
  {32'h4120fa94, 32'hc029be98} /* (14, 19, 28) {real, imag} */,
  {32'h408adb4e, 32'hc139b1b8} /* (14, 19, 27) {real, imag} */,
  {32'hc1746756, 32'hc17d4e2e} /* (14, 19, 26) {real, imag} */,
  {32'hc0e328f9, 32'hc00fa14e} /* (14, 19, 25) {real, imag} */,
  {32'h41170980, 32'hc11c0854} /* (14, 19, 24) {real, imag} */,
  {32'h3ffcd9ca, 32'h40ee8f1f} /* (14, 19, 23) {real, imag} */,
  {32'h3fbb5044, 32'hc0c394db} /* (14, 19, 22) {real, imag} */,
  {32'hc0c56c5e, 32'hc025a658} /* (14, 19, 21) {real, imag} */,
  {32'hc0e64fb2, 32'hc0a812ed} /* (14, 19, 20) {real, imag} */,
  {32'h408af11d, 32'hbfb58a40} /* (14, 19, 19) {real, imag} */,
  {32'h409d9a78, 32'hc02655f7} /* (14, 19, 18) {real, imag} */,
  {32'h3ffe971e, 32'h3eb214a0} /* (14, 19, 17) {real, imag} */,
  {32'hc0614010, 32'h3ffa029c} /* (14, 19, 16) {real, imag} */,
  {32'h3ffdacd6, 32'hbfd90d78} /* (14, 19, 15) {real, imag} */,
  {32'hc06eb6a8, 32'hbf366fd9} /* (14, 19, 14) {real, imag} */,
  {32'hc0be6bb3, 32'h3f849378} /* (14, 19, 13) {real, imag} */,
  {32'hbfb50fa8, 32'hbe8fe0b0} /* (14, 19, 12) {real, imag} */,
  {32'hbef83f28, 32'h40af6764} /* (14, 19, 11) {real, imag} */,
  {32'h40477fc6, 32'hbe2ceae0} /* (14, 19, 10) {real, imag} */,
  {32'h3e89ea2a, 32'h403a9006} /* (14, 19, 9) {real, imag} */,
  {32'hc04d0d2a, 32'h40dd1a6c} /* (14, 19, 8) {real, imag} */,
  {32'hc1123de0, 32'hc102d312} /* (14, 19, 7) {real, imag} */,
  {32'h411b440a, 32'h4122fea4} /* (14, 19, 6) {real, imag} */,
  {32'hc08412e6, 32'h4112ab98} /* (14, 19, 5) {real, imag} */,
  {32'h3fa9698c, 32'h410b6abb} /* (14, 19, 4) {real, imag} */,
  {32'h40f75a79, 32'hc0b2a339} /* (14, 19, 3) {real, imag} */,
  {32'hc034fde8, 32'h3d6047f0} /* (14, 19, 2) {real, imag} */,
  {32'hc17d65e9, 32'hc0b5b886} /* (14, 19, 1) {real, imag} */,
  {32'hc180a651, 32'h41708c86} /* (14, 19, 0) {real, imag} */,
  {32'h3f9284c6, 32'hc10b68f2} /* (14, 18, 31) {real, imag} */,
  {32'h3f9c8fc0, 32'h408d4e14} /* (14, 18, 30) {real, imag} */,
  {32'h3fb0148c, 32'h415c921c} /* (14, 18, 29) {real, imag} */,
  {32'hbfebf4f0, 32'hc0a90304} /* (14, 18, 28) {real, imag} */,
  {32'h3f9311d0, 32'h414931f0} /* (14, 18, 27) {real, imag} */,
  {32'h408dbdd3, 32'hbfe54e5a} /* (14, 18, 26) {real, imag} */,
  {32'h412d1db1, 32'hc09e74bc} /* (14, 18, 25) {real, imag} */,
  {32'h4011790b, 32'hc032c5d2} /* (14, 18, 24) {real, imag} */,
  {32'hc16042e1, 32'h411d284a} /* (14, 18, 23) {real, imag} */,
  {32'h412e3570, 32'h3f84c46c} /* (14, 18, 22) {real, imag} */,
  {32'h40b4df8d, 32'hbecebdf0} /* (14, 18, 21) {real, imag} */,
  {32'h4065a253, 32'hc0bee161} /* (14, 18, 20) {real, imag} */,
  {32'h4057bbc8, 32'h40a31c6c} /* (14, 18, 19) {real, imag} */,
  {32'h3f533d80, 32'hbf7e47d1} /* (14, 18, 18) {real, imag} */,
  {32'h3f4b326c, 32'hbfd72022} /* (14, 18, 17) {real, imag} */,
  {32'h401d55e6, 32'h3f016bc6} /* (14, 18, 16) {real, imag} */,
  {32'h3fb781ba, 32'h3f9f82f2} /* (14, 18, 15) {real, imag} */,
  {32'hc02c1248, 32'h3fcb172c} /* (14, 18, 14) {real, imag} */,
  {32'hc0c74fd0, 32'hc08953e8} /* (14, 18, 13) {real, imag} */,
  {32'hc0bdff5a, 32'h40b5565f} /* (14, 18, 12) {real, imag} */,
  {32'hbfab59a8, 32'h40d2db3d} /* (14, 18, 11) {real, imag} */,
  {32'hc0feb9b8, 32'h3fd2ca0c} /* (14, 18, 10) {real, imag} */,
  {32'hc0ba8aaa, 32'hbf20c520} /* (14, 18, 9) {real, imag} */,
  {32'hbf4c6ce4, 32'h401e5cd4} /* (14, 18, 8) {real, imag} */,
  {32'hc0e4cf06, 32'hbffcc732} /* (14, 18, 7) {real, imag} */,
  {32'hc1083e84, 32'hc07aee4f} /* (14, 18, 6) {real, imag} */,
  {32'hc088d089, 32'h3e400760} /* (14, 18, 5) {real, imag} */,
  {32'h418bba08, 32'hc0af7e1a} /* (14, 18, 4) {real, imag} */,
  {32'hc0adb3c9, 32'hc0ed9f4c} /* (14, 18, 3) {real, imag} */,
  {32'h410194a2, 32'hc0975b94} /* (14, 18, 2) {real, imag} */,
  {32'hbf59323c, 32'hc15739b0} /* (14, 18, 1) {real, imag} */,
  {32'hc07ba1a4, 32'hc0852b1a} /* (14, 18, 0) {real, imag} */,
  {32'hc12ccf6a, 32'h3fdff703} /* (14, 17, 31) {real, imag} */,
  {32'hc0c68e40, 32'hc087309c} /* (14, 17, 30) {real, imag} */,
  {32'h409c709b, 32'hbfeec043} /* (14, 17, 29) {real, imag} */,
  {32'hc119f91d, 32'hc0b6d2e9} /* (14, 17, 28) {real, imag} */,
  {32'h402fd12a, 32'hc0a0eb6b} /* (14, 17, 27) {real, imag} */,
  {32'hc049f6ee, 32'h3e9dd730} /* (14, 17, 26) {real, imag} */,
  {32'hc0b1e0b1, 32'h40b19a2e} /* (14, 17, 25) {real, imag} */,
  {32'h404d5a6c, 32'hc04b59d7} /* (14, 17, 24) {real, imag} */,
  {32'h4110424c, 32'hc0a5d4b6} /* (14, 17, 23) {real, imag} */,
  {32'h411183ce, 32'hbf8c502e} /* (14, 17, 22) {real, imag} */,
  {32'hc08cfcc0, 32'h401d9108} /* (14, 17, 21) {real, imag} */,
  {32'hc0159e9c, 32'h412b848a} /* (14, 17, 20) {real, imag} */,
  {32'hc05c9780, 32'hbec2a780} /* (14, 17, 19) {real, imag} */,
  {32'hc05f9deb, 32'h409babdc} /* (14, 17, 18) {real, imag} */,
  {32'hc05eed6f, 32'h3fcb8449} /* (14, 17, 17) {real, imag} */,
  {32'h3f5f29ae, 32'h3fd7993c} /* (14, 17, 16) {real, imag} */,
  {32'hbf7216bc, 32'hc00adbbc} /* (14, 17, 15) {real, imag} */,
  {32'h3fb6ad8a, 32'h3f2a78a0} /* (14, 17, 14) {real, imag} */,
  {32'hbfd9edc5, 32'h40a4a4be} /* (14, 17, 13) {real, imag} */,
  {32'hc00fb926, 32'hc0160fea} /* (14, 17, 12) {real, imag} */,
  {32'hc05c3b7e, 32'hbdbc5f00} /* (14, 17, 11) {real, imag} */,
  {32'h409bc94d, 32'hc085958a} /* (14, 17, 10) {real, imag} */,
  {32'h4022e062, 32'h4083a412} /* (14, 17, 9) {real, imag} */,
  {32'h407510fc, 32'h40b9e12e} /* (14, 17, 8) {real, imag} */,
  {32'hc1000e7a, 32'h3f81899a} /* (14, 17, 7) {real, imag} */,
  {32'h40b3172d, 32'h4161406a} /* (14, 17, 6) {real, imag} */,
  {32'hbed58efc, 32'h40676386} /* (14, 17, 5) {real, imag} */,
  {32'h40a0691e, 32'hc19574c8} /* (14, 17, 4) {real, imag} */,
  {32'h415fe12a, 32'hbff6e3e3} /* (14, 17, 3) {real, imag} */,
  {32'h4090855c, 32'h409bed90} /* (14, 17, 2) {real, imag} */,
  {32'h4064ba17, 32'hc05ce27e} /* (14, 17, 1) {real, imag} */,
  {32'h407f7684, 32'hbf96eb84} /* (14, 17, 0) {real, imag} */,
  {32'hc08410c2, 32'h3f6e71d0} /* (14, 16, 31) {real, imag} */,
  {32'hc0839d3c, 32'hc0c3112e} /* (14, 16, 30) {real, imag} */,
  {32'hc0467e7e, 32'hc0ad62f8} /* (14, 16, 29) {real, imag} */,
  {32'h40c0a79a, 32'h40ec62bf} /* (14, 16, 28) {real, imag} */,
  {32'hc01c081f, 32'h40d88f0f} /* (14, 16, 27) {real, imag} */,
  {32'hc100986c, 32'h40e7c143} /* (14, 16, 26) {real, imag} */,
  {32'h40a40e23, 32'hc0dcf4a3} /* (14, 16, 25) {real, imag} */,
  {32'hc0515860, 32'hc02b1222} /* (14, 16, 24) {real, imag} */,
  {32'h4074ce1e, 32'h406760e2} /* (14, 16, 23) {real, imag} */,
  {32'h403798d8, 32'hc0821c39} /* (14, 16, 22) {real, imag} */,
  {32'hbe247430, 32'hbf6fc0d4} /* (14, 16, 21) {real, imag} */,
  {32'h403b200c, 32'h3e2cbb20} /* (14, 16, 20) {real, imag} */,
  {32'h40668a1f, 32'h40784b70} /* (14, 16, 19) {real, imag} */,
  {32'hc036276a, 32'h400ec761} /* (14, 16, 18) {real, imag} */,
  {32'hbebde55e, 32'hbf16bcd0} /* (14, 16, 17) {real, imag} */,
  {32'h3e1f7620, 32'hbfa84858} /* (14, 16, 16) {real, imag} */,
  {32'h3e03c0a4, 32'h3f3e4d10} /* (14, 16, 15) {real, imag} */,
  {32'h3f733e98, 32'hbf566c2c} /* (14, 16, 14) {real, imag} */,
  {32'hc02ec959, 32'hbfd5bbeb} /* (14, 16, 13) {real, imag} */,
  {32'h3fe1f3f7, 32'h3f998608} /* (14, 16, 12) {real, imag} */,
  {32'hbf9d130e, 32'hbe61fa72} /* (14, 16, 11) {real, imag} */,
  {32'hbf27d5d0, 32'hc127c720} /* (14, 16, 10) {real, imag} */,
  {32'h3fa57430, 32'hc05e0442} /* (14, 16, 9) {real, imag} */,
  {32'hbfee4743, 32'h3ff7f919} /* (14, 16, 8) {real, imag} */,
  {32'hc02245f0, 32'hbfb385dc} /* (14, 16, 7) {real, imag} */,
  {32'hbf869ab4, 32'h4048965a} /* (14, 16, 6) {real, imag} */,
  {32'h4107e0e9, 32'h40daf037} /* (14, 16, 5) {real, imag} */,
  {32'h40952286, 32'h3eca04a0} /* (14, 16, 4) {real, imag} */,
  {32'h40bbb40d, 32'hc08cc296} /* (14, 16, 3) {real, imag} */,
  {32'hc10a7411, 32'h41643791} /* (14, 16, 2) {real, imag} */,
  {32'h3f926ebe, 32'hc19ae01e} /* (14, 16, 1) {real, imag} */,
  {32'h40575fb0, 32'h402b3397} /* (14, 16, 0) {real, imag} */,
  {32'hc0d41623, 32'hc1814241} /* (14, 15, 31) {real, imag} */,
  {32'h3e217d48, 32'hc0040b68} /* (14, 15, 30) {real, imag} */,
  {32'h411b52ac, 32'hc0fe3601} /* (14, 15, 29) {real, imag} */,
  {32'hc13d646d, 32'h3f6ccd18} /* (14, 15, 28) {real, imag} */,
  {32'h40b05918, 32'hbfb17f39} /* (14, 15, 27) {real, imag} */,
  {32'hc0dcf07e, 32'h4005c958} /* (14, 15, 26) {real, imag} */,
  {32'h405f6030, 32'h407ca96a} /* (14, 15, 25) {real, imag} */,
  {32'hc0b3f0bc, 32'hc07afc14} /* (14, 15, 24) {real, imag} */,
  {32'hbfbf4b0f, 32'h40a0aa4b} /* (14, 15, 23) {real, imag} */,
  {32'h4103ffb4, 32'hc0d1094c} /* (14, 15, 22) {real, imag} */,
  {32'h40940a4b, 32'h408e044a} /* (14, 15, 21) {real, imag} */,
  {32'h3f3673d0, 32'hc02191bf} /* (14, 15, 20) {real, imag} */,
  {32'hc028ec8c, 32'h3fbc10c2} /* (14, 15, 19) {real, imag} */,
  {32'h3f267ad6, 32'h3ec8d218} /* (14, 15, 18) {real, imag} */,
  {32'h3ead6604, 32'h3f3befb0} /* (14, 15, 17) {real, imag} */,
  {32'hbf020c90, 32'hc06afc5a} /* (14, 15, 16) {real, imag} */,
  {32'h3fc36cd1, 32'hc00d152c} /* (14, 15, 15) {real, imag} */,
  {32'h3fc4f7dd, 32'hc071c559} /* (14, 15, 14) {real, imag} */,
  {32'hc0685d00, 32'h4094bac2} /* (14, 15, 13) {real, imag} */,
  {32'hc061ac90, 32'hbeda7fa8} /* (14, 15, 12) {real, imag} */,
  {32'hc0909653, 32'hc0d51d4e} /* (14, 15, 11) {real, imag} */,
  {32'h408ef217, 32'hbf26c18c} /* (14, 15, 10) {real, imag} */,
  {32'h403e43bc, 32'hbf5904b8} /* (14, 15, 9) {real, imag} */,
  {32'hc0031940, 32'h415593d1} /* (14, 15, 8) {real, imag} */,
  {32'h4071c9bc, 32'hbe4eb058} /* (14, 15, 7) {real, imag} */,
  {32'h4147f1d9, 32'hc1231c54} /* (14, 15, 6) {real, imag} */,
  {32'hc00ea75b, 32'hbf96b805} /* (14, 15, 5) {real, imag} */,
  {32'h4101efdf, 32'h4130e602} /* (14, 15, 4) {real, imag} */,
  {32'h409295de, 32'h3fcb50ac} /* (14, 15, 3) {real, imag} */,
  {32'h40021c4e, 32'h418696af} /* (14, 15, 2) {real, imag} */,
  {32'h411ddb5d, 32'hc091b79b} /* (14, 15, 1) {real, imag} */,
  {32'hc1583cfd, 32'hc0c0124f} /* (14, 15, 0) {real, imag} */,
  {32'h3f2e5d90, 32'h410f50f0} /* (14, 14, 31) {real, imag} */,
  {32'hc0620150, 32'hc142f1de} /* (14, 14, 30) {real, imag} */,
  {32'hbff2f8f0, 32'h4089c4b5} /* (14, 14, 29) {real, imag} */,
  {32'h40928544, 32'hbfe8b9b8} /* (14, 14, 28) {real, imag} */,
  {32'h4187bf7c, 32'h41453ea6} /* (14, 14, 27) {real, imag} */,
  {32'h401b47d4, 32'hc11b11db} /* (14, 14, 26) {real, imag} */,
  {32'hc024d132, 32'hbc085d00} /* (14, 14, 25) {real, imag} */,
  {32'h40fbf163, 32'hc0b34ead} /* (14, 14, 24) {real, imag} */,
  {32'hc0d17072, 32'hc140c914} /* (14, 14, 23) {real, imag} */,
  {32'hc0257ecb, 32'h3f2d6f70} /* (14, 14, 22) {real, imag} */,
  {32'h407b1e2e, 32'hbf384994} /* (14, 14, 21) {real, imag} */,
  {32'hbfac07cd, 32'hc08dc24d} /* (14, 14, 20) {real, imag} */,
  {32'h3e8cc4d0, 32'h3fc5a16c} /* (14, 14, 19) {real, imag} */,
  {32'h4044f9d4, 32'h3fc1cac6} /* (14, 14, 18) {real, imag} */,
  {32'h3fa4d937, 32'h3fe526e8} /* (14, 14, 17) {real, imag} */,
  {32'hbf90226a, 32'hc054a43e} /* (14, 14, 16) {real, imag} */,
  {32'h3ee681fc, 32'hbf8299f8} /* (14, 14, 15) {real, imag} */,
  {32'hbeee2b74, 32'hc02bfbf9} /* (14, 14, 14) {real, imag} */,
  {32'h401a4a78, 32'hc0b93e09} /* (14, 14, 13) {real, imag} */,
  {32'h3f9c3acb, 32'hc01f7900} /* (14, 14, 12) {real, imag} */,
  {32'h40b22edb, 32'hc0872b84} /* (14, 14, 11) {real, imag} */,
  {32'h3f25068c, 32'h3fd57b2c} /* (14, 14, 10) {real, imag} */,
  {32'h3f592a20, 32'h41598930} /* (14, 14, 9) {real, imag} */,
  {32'hc1285392, 32'h40412636} /* (14, 14, 8) {real, imag} */,
  {32'hc058c722, 32'hc098595e} /* (14, 14, 7) {real, imag} */,
  {32'h41795701, 32'h40b0ef26} /* (14, 14, 6) {real, imag} */,
  {32'h4061ff9c, 32'hc0cba264} /* (14, 14, 5) {real, imag} */,
  {32'hc0b080b4, 32'h413c73eb} /* (14, 14, 4) {real, imag} */,
  {32'hc0e6927c, 32'hc118af02} /* (14, 14, 3) {real, imag} */,
  {32'h40b36650, 32'h40038fa6} /* (14, 14, 2) {real, imag} */,
  {32'h40d15b78, 32'hc0952510} /* (14, 14, 1) {real, imag} */,
  {32'hbf095234, 32'hbf9a8604} /* (14, 14, 0) {real, imag} */,
  {32'h40bf97d7, 32'hbf2a9a00} /* (14, 13, 31) {real, imag} */,
  {32'h4160d038, 32'h417586ce} /* (14, 13, 30) {real, imag} */,
  {32'hc07459bf, 32'hbf47af50} /* (14, 13, 29) {real, imag} */,
  {32'h3f6464c5, 32'hc117a7c4} /* (14, 13, 28) {real, imag} */,
  {32'h40c2fe8c, 32'h4065a048} /* (14, 13, 27) {real, imag} */,
  {32'hc0e3966a, 32'hc151f7fe} /* (14, 13, 26) {real, imag} */,
  {32'h41197dd3, 32'hc0f556bc} /* (14, 13, 25) {real, imag} */,
  {32'hc137d929, 32'h3ed3ba20} /* (14, 13, 24) {real, imag} */,
  {32'hbfd394e8, 32'h41875cde} /* (14, 13, 23) {real, imag} */,
  {32'h414487c8, 32'hc0bb2421} /* (14, 13, 22) {real, imag} */,
  {32'hc0bfb6f6, 32'h40530a0e} /* (14, 13, 21) {real, imag} */,
  {32'h40bfa732, 32'hc0921384} /* (14, 13, 20) {real, imag} */,
  {32'h3e81d470, 32'hbf94ac60} /* (14, 13, 19) {real, imag} */,
  {32'h3f164890, 32'h3fbd45fc} /* (14, 13, 18) {real, imag} */,
  {32'hbff19e46, 32'h40900ede} /* (14, 13, 17) {real, imag} */,
  {32'hbf885740, 32'hbf0a5638} /* (14, 13, 16) {real, imag} */,
  {32'h40638951, 32'h3f885ccf} /* (14, 13, 15) {real, imag} */,
  {32'hc019e1be, 32'h3fb991f4} /* (14, 13, 14) {real, imag} */,
  {32'h40984c93, 32'hc0d20ab1} /* (14, 13, 13) {real, imag} */,
  {32'h410bc418, 32'hbf9e4bee} /* (14, 13, 12) {real, imag} */,
  {32'h3fcd45a0, 32'hc072f9d6} /* (14, 13, 11) {real, imag} */,
  {32'hc09e60b8, 32'hbf4cd2e8} /* (14, 13, 10) {real, imag} */,
  {32'hbf9ee380, 32'h414be64c} /* (14, 13, 9) {real, imag} */,
  {32'hc1049abd, 32'hc08f004a} /* (14, 13, 8) {real, imag} */,
  {32'hc16febc5, 32'hbfe319b0} /* (14, 13, 7) {real, imag} */,
  {32'hc124c599, 32'hc070c758} /* (14, 13, 6) {real, imag} */,
  {32'h4120ef3e, 32'hc10721d5} /* (14, 13, 5) {real, imag} */,
  {32'hbe8477aa, 32'h40c276df} /* (14, 13, 4) {real, imag} */,
  {32'hc0d9cba6, 32'h4118f551} /* (14, 13, 3) {real, imag} */,
  {32'hc032e400, 32'h41960721} /* (14, 13, 2) {real, imag} */,
  {32'h408eb0c5, 32'hbf0b40a0} /* (14, 13, 1) {real, imag} */,
  {32'hc1ed5bc9, 32'hc110658a} /* (14, 13, 0) {real, imag} */,
  {32'hc1105b9c, 32'hc131431a} /* (14, 12, 31) {real, imag} */,
  {32'hc14b7425, 32'hbfa6ff48} /* (14, 12, 30) {real, imag} */,
  {32'hc1fc7274, 32'hc121a4b5} /* (14, 12, 29) {real, imag} */,
  {32'h412f7218, 32'h4202c070} /* (14, 12, 28) {real, imag} */,
  {32'h418db6ff, 32'h3fef8f11} /* (14, 12, 27) {real, imag} */,
  {32'hc0fbd38e, 32'h41459bc8} /* (14, 12, 26) {real, imag} */,
  {32'h40e49d74, 32'hbe5d5940} /* (14, 12, 25) {real, imag} */,
  {32'h40431194, 32'h40adc25b} /* (14, 12, 24) {real, imag} */,
  {32'h40a378bc, 32'h412ab7ea} /* (14, 12, 23) {real, imag} */,
  {32'h40505ebc, 32'hc1100f3c} /* (14, 12, 22) {real, imag} */,
  {32'h401581b2, 32'hc0a85071} /* (14, 12, 21) {real, imag} */,
  {32'hc0e2416a, 32'h406dbbd6} /* (14, 12, 20) {real, imag} */,
  {32'hbffa26e8, 32'hbf82e13a} /* (14, 12, 19) {real, imag} */,
  {32'h3fb0b168, 32'hbf1a3c60} /* (14, 12, 18) {real, imag} */,
  {32'hbeee5b30, 32'h3ef4f47c} /* (14, 12, 17) {real, imag} */,
  {32'hbdfe4460, 32'h407f2a90} /* (14, 12, 16) {real, imag} */,
  {32'hc0b029cb, 32'h4070e2c8} /* (14, 12, 15) {real, imag} */,
  {32'hc02bba72, 32'hc1256598} /* (14, 12, 14) {real, imag} */,
  {32'hc03cd214, 32'hbeff9b38} /* (14, 12, 13) {real, imag} */,
  {32'h3fe853f8, 32'h400635fa} /* (14, 12, 12) {real, imag} */,
  {32'hc09b5367, 32'h40e9a71f} /* (14, 12, 11) {real, imag} */,
  {32'h41817ebc, 32'hc04d691f} /* (14, 12, 10) {real, imag} */,
  {32'hc094d7f8, 32'h3f41dd50} /* (14, 12, 9) {real, imag} */,
  {32'hc1a57d30, 32'hc0b9ce95} /* (14, 12, 8) {real, imag} */,
  {32'h40fab21c, 32'hc11da2a8} /* (14, 12, 7) {real, imag} */,
  {32'h3f8382c8, 32'hc105af0c} /* (14, 12, 6) {real, imag} */,
  {32'hc18280fd, 32'h3f43a98a} /* (14, 12, 5) {real, imag} */,
  {32'h4172722c, 32'h3f7230e0} /* (14, 12, 4) {real, imag} */,
  {32'h407e7344, 32'hc04d8388} /* (14, 12, 3) {real, imag} */,
  {32'hc004776c, 32'hc14b7f29} /* (14, 12, 2) {real, imag} */,
  {32'h410ab55c, 32'hc165a37a} /* (14, 12, 1) {real, imag} */,
  {32'hc003c2f5, 32'hc1f8b1ba} /* (14, 12, 0) {real, imag} */,
  {32'hc0f3c933, 32'h4113c4a6} /* (14, 11, 31) {real, imag} */,
  {32'hc015005a, 32'hc0f32458} /* (14, 11, 30) {real, imag} */,
  {32'h41aacc23, 32'h4113787d} /* (14, 11, 29) {real, imag} */,
  {32'h40477a2a, 32'hc15677cf} /* (14, 11, 28) {real, imag} */,
  {32'h40f54c61, 32'h41bb6ce6} /* (14, 11, 27) {real, imag} */,
  {32'hc1083f68, 32'hc0a4bd30} /* (14, 11, 26) {real, imag} */,
  {32'hc096a2a3, 32'h4136f8ef} /* (14, 11, 25) {real, imag} */,
  {32'h401f8142, 32'h41439bd2} /* (14, 11, 24) {real, imag} */,
  {32'hbf2a2404, 32'hc10c9954} /* (14, 11, 23) {real, imag} */,
  {32'h403d9b4c, 32'hbfd74b42} /* (14, 11, 22) {real, imag} */,
  {32'h40a3507c, 32'hc0cebb12} /* (14, 11, 21) {real, imag} */,
  {32'h401c9e74, 32'h40f99d44} /* (14, 11, 20) {real, imag} */,
  {32'hc00018a0, 32'h413b1fe2} /* (14, 11, 19) {real, imag} */,
  {32'h401413fb, 32'h40c1b1eb} /* (14, 11, 18) {real, imag} */,
  {32'hbffd2e81, 32'hc11c835d} /* (14, 11, 17) {real, imag} */,
  {32'hc0ab0e25, 32'h4100e6d4} /* (14, 11, 16) {real, imag} */,
  {32'hc080ea2e, 32'hc047ca95} /* (14, 11, 15) {real, imag} */,
  {32'h40286519, 32'hc0936177} /* (14, 11, 14) {real, imag} */,
  {32'h407d82b8, 32'hc102a9b0} /* (14, 11, 13) {real, imag} */,
  {32'h400d2524, 32'h40075b59} /* (14, 11, 12) {real, imag} */,
  {32'h417dd46a, 32'hc06a289c} /* (14, 11, 11) {real, imag} */,
  {32'hbf282970, 32'hbff6ee9e} /* (14, 11, 10) {real, imag} */,
  {32'hbfd5f52e, 32'h4083bb6c} /* (14, 11, 9) {real, imag} */,
  {32'h414e68f6, 32'h416b2bc0} /* (14, 11, 8) {real, imag} */,
  {32'h4124338a, 32'h408fb6a6} /* (14, 11, 7) {real, imag} */,
  {32'h4199fce8, 32'h4033246b} /* (14, 11, 6) {real, imag} */,
  {32'hc1294e60, 32'hbfd1bca8} /* (14, 11, 5) {real, imag} */,
  {32'hc13d5404, 32'hc1b43420} /* (14, 11, 4) {real, imag} */,
  {32'hbfc5d460, 32'hc19b1398} /* (14, 11, 3) {real, imag} */,
  {32'hc14dd2f4, 32'hc1f71732} /* (14, 11, 2) {real, imag} */,
  {32'h3f3aac38, 32'hbea28180} /* (14, 11, 1) {real, imag} */,
  {32'hbf3a3d48, 32'h414fb3aa} /* (14, 11, 0) {real, imag} */,
  {32'hc0ffc66c, 32'hc1883e31} /* (14, 10, 31) {real, imag} */,
  {32'h41f198c1, 32'h418db334} /* (14, 10, 30) {real, imag} */,
  {32'hc133e438, 32'hbe59f490} /* (14, 10, 29) {real, imag} */,
  {32'hc0ed9091, 32'h40f022cf} /* (14, 10, 28) {real, imag} */,
  {32'h3d67e180, 32'h41011433} /* (14, 10, 27) {real, imag} */,
  {32'h4228dd18, 32'h4097c1c2} /* (14, 10, 26) {real, imag} */,
  {32'h40022c64, 32'h3fd39e92} /* (14, 10, 25) {real, imag} */,
  {32'hbfe9b918, 32'h3e77bda0} /* (14, 10, 24) {real, imag} */,
  {32'hc044606b, 32'hc042e71f} /* (14, 10, 23) {real, imag} */,
  {32'hc129f330, 32'hc17ff76e} /* (14, 10, 22) {real, imag} */,
  {32'hbf27f5f8, 32'hc1186854} /* (14, 10, 21) {real, imag} */,
  {32'h4023a0a5, 32'h40b28afc} /* (14, 10, 20) {real, imag} */,
  {32'h412d76dc, 32'hc09ddd86} /* (14, 10, 19) {real, imag} */,
  {32'hbee706f8, 32'hc0c9cdfe} /* (14, 10, 18) {real, imag} */,
  {32'hc10ff578, 32'h4085459f} /* (14, 10, 17) {real, imag} */,
  {32'hc11df1ae, 32'hbfd5019f} /* (14, 10, 16) {real, imag} */,
  {32'h401aaad2, 32'hc088e9c1} /* (14, 10, 15) {real, imag} */,
  {32'hc0d37ac8, 32'h410e90bc} /* (14, 10, 14) {real, imag} */,
  {32'hc0c95651, 32'hc18b209e} /* (14, 10, 13) {real, imag} */,
  {32'h3f344fb8, 32'hc0b75336} /* (14, 10, 12) {real, imag} */,
  {32'h40d0a715, 32'h405da29e} /* (14, 10, 11) {real, imag} */,
  {32'h41a44774, 32'h40454328} /* (14, 10, 10) {real, imag} */,
  {32'h3f9caf3e, 32'hc017db09} /* (14, 10, 9) {real, imag} */,
  {32'hc12870bb, 32'hc094654b} /* (14, 10, 8) {real, imag} */,
  {32'h41860416, 32'h408b90b8} /* (14, 10, 7) {real, imag} */,
  {32'h415f4c78, 32'hc0f95896} /* (14, 10, 6) {real, imag} */,
  {32'h40aad1f7, 32'h408beb28} /* (14, 10, 5) {real, imag} */,
  {32'h40128cca, 32'hc1b789e6} /* (14, 10, 4) {real, imag} */,
  {32'hbc215a00, 32'h40dbdd30} /* (14, 10, 3) {real, imag} */,
  {32'hc1c30b1d, 32'hbe247400} /* (14, 10, 2) {real, imag} */,
  {32'hc1cc04cb, 32'h420d763a} /* (14, 10, 1) {real, imag} */,
  {32'h41e4cd87, 32'hbfcd6373} /* (14, 10, 0) {real, imag} */,
  {32'h41e5095c, 32'hc1669d9c} /* (14, 9, 31) {real, imag} */,
  {32'h41ae7d6a, 32'hc14cc1e2} /* (14, 9, 30) {real, imag} */,
  {32'hc144a272, 32'h421050b0} /* (14, 9, 29) {real, imag} */,
  {32'hc2570671, 32'hc1bef99e} /* (14, 9, 28) {real, imag} */,
  {32'hc21ebaac, 32'h4188b142} /* (14, 9, 27) {real, imag} */,
  {32'h41806a20, 32'hc1246a27} /* (14, 9, 26) {real, imag} */,
  {32'h40c6e94f, 32'hbffa68a8} /* (14, 9, 25) {real, imag} */,
  {32'hbfefd034, 32'hc12298ec} /* (14, 9, 24) {real, imag} */,
  {32'h4101eb7a, 32'h3f83ce6e} /* (14, 9, 23) {real, imag} */,
  {32'h4188eb49, 32'hc132685d} /* (14, 9, 22) {real, imag} */,
  {32'hc109e0f0, 32'h403dd1ce} /* (14, 9, 21) {real, imag} */,
  {32'hc07d7e08, 32'h4101989c} /* (14, 9, 20) {real, imag} */,
  {32'h403446fe, 32'hc0ce2263} /* (14, 9, 19) {real, imag} */,
  {32'hbfa069f4, 32'hc05a3ae4} /* (14, 9, 18) {real, imag} */,
  {32'hc0e004d2, 32'h3f72cb78} /* (14, 9, 17) {real, imag} */,
  {32'h40e67b37, 32'hc0d8aa65} /* (14, 9, 16) {real, imag} */,
  {32'hbf312930, 32'hc10a078a} /* (14, 9, 15) {real, imag} */,
  {32'h40ae4b9f, 32'h40f49f06} /* (14, 9, 14) {real, imag} */,
  {32'hc11460c4, 32'hc0ec1e93} /* (14, 9, 13) {real, imag} */,
  {32'hc024e228, 32'h414ed96e} /* (14, 9, 12) {real, imag} */,
  {32'hbf4c2508, 32'h41789bfc} /* (14, 9, 11) {real, imag} */,
  {32'h41522dfa, 32'hc0a49b6a} /* (14, 9, 10) {real, imag} */,
  {32'hc154c1d2, 32'hc0cfa950} /* (14, 9, 9) {real, imag} */,
  {32'h3f9826f4, 32'h4181961c} /* (14, 9, 8) {real, imag} */,
  {32'h40b5be4b, 32'hc1196729} /* (14, 9, 7) {real, imag} */,
  {32'hc148e5ac, 32'h3e9f63e0} /* (14, 9, 6) {real, imag} */,
  {32'h41775cd0, 32'h40293c8e} /* (14, 9, 5) {real, imag} */,
  {32'hc19dd99e, 32'h4193e862} /* (14, 9, 4) {real, imag} */,
  {32'hc1a57691, 32'h40112448} /* (14, 9, 3) {real, imag} */,
  {32'hc0a37e9a, 32'hbfe0a9b0} /* (14, 9, 2) {real, imag} */,
  {32'hc134b197, 32'hc1a93116} /* (14, 9, 1) {real, imag} */,
  {32'h415f3a98, 32'hc1919c7d} /* (14, 9, 0) {real, imag} */,
  {32'h42273cb1, 32'h4239affc} /* (14, 8, 31) {real, imag} */,
  {32'hc108b960, 32'h410d5ef0} /* (14, 8, 30) {real, imag} */,
  {32'hbee233c8, 32'hc1d98284} /* (14, 8, 29) {real, imag} */,
  {32'hbfe01cbc, 32'h41c904c4} /* (14, 8, 28) {real, imag} */,
  {32'h402fd98c, 32'hc1a87052} /* (14, 8, 27) {real, imag} */,
  {32'h41bacaed, 32'h3f026810} /* (14, 8, 26) {real, imag} */,
  {32'h4185c5cc, 32'hc1a2d598} /* (14, 8, 25) {real, imag} */,
  {32'h40842854, 32'h418ef6d4} /* (14, 8, 24) {real, imag} */,
  {32'hc11d0398, 32'hc1a90171} /* (14, 8, 23) {real, imag} */,
  {32'hc1431d4d, 32'hc15cd6a5} /* (14, 8, 22) {real, imag} */,
  {32'hc023f4a8, 32'hc015ee17} /* (14, 8, 21) {real, imag} */,
  {32'h411fb21c, 32'hc12421bd} /* (14, 8, 20) {real, imag} */,
  {32'hc0ec0927, 32'h410b6b6e} /* (14, 8, 19) {real, imag} */,
  {32'h410f9926, 32'h3e1a74e0} /* (14, 8, 18) {real, imag} */,
  {32'hbf81eab4, 32'hc00dafa0} /* (14, 8, 17) {real, imag} */,
  {32'hc11c8314, 32'h3f148448} /* (14, 8, 16) {real, imag} */,
  {32'hc02da076, 32'hc0871ae4} /* (14, 8, 15) {real, imag} */,
  {32'hbfa20c1c, 32'h40e11300} /* (14, 8, 14) {real, imag} */,
  {32'hbf785718, 32'h4110a4be} /* (14, 8, 13) {real, imag} */,
  {32'hc0916d8d, 32'hc0dea326} /* (14, 8, 12) {real, imag} */,
  {32'hc1c2829b, 32'hc02797b1} /* (14, 8, 11) {real, imag} */,
  {32'h409aa03a, 32'hbff59f68} /* (14, 8, 10) {real, imag} */,
  {32'hc13c84d2, 32'hc1c6f341} /* (14, 8, 9) {real, imag} */,
  {32'hc1e12805, 32'h40b383ff} /* (14, 8, 8) {real, imag} */,
  {32'hc0ab610e, 32'h40602480} /* (14, 8, 7) {real, imag} */,
  {32'hc1cdc9d3, 32'hc1ae9da4} /* (14, 8, 6) {real, imag} */,
  {32'hc03f1490, 32'hc1908372} /* (14, 8, 5) {real, imag} */,
  {32'hc177f7da, 32'hc1926c68} /* (14, 8, 4) {real, imag} */,
  {32'hc0867848, 32'hc16fb314} /* (14, 8, 3) {real, imag} */,
  {32'h41747096, 32'h401ce8f9} /* (14, 8, 2) {real, imag} */,
  {32'h41da3a56, 32'hbf15be80} /* (14, 8, 1) {real, imag} */,
  {32'hc025899c, 32'h40207912} /* (14, 8, 0) {real, imag} */,
  {32'h41abdf84, 32'hc15d3e7c} /* (14, 7, 31) {real, imag} */,
  {32'hc230008a, 32'hc1939bb4} /* (14, 7, 30) {real, imag} */,
  {32'h4177edac, 32'h4176dd4b} /* (14, 7, 29) {real, imag} */,
  {32'h421e3124, 32'hc266278c} /* (14, 7, 28) {real, imag} */,
  {32'hc1b416a1, 32'h41c76963} /* (14, 7, 27) {real, imag} */,
  {32'h416dee50, 32'h420cad43} /* (14, 7, 26) {real, imag} */,
  {32'hc1e99501, 32'h4160abd2} /* (14, 7, 25) {real, imag} */,
  {32'h4126156c, 32'hc18c1546} /* (14, 7, 24) {real, imag} */,
  {32'hc0269d90, 32'h410c85fc} /* (14, 7, 23) {real, imag} */,
  {32'hc11ebf94, 32'hc1a26062} /* (14, 7, 22) {real, imag} */,
  {32'hbfbac11c, 32'hc1848e6f} /* (14, 7, 21) {real, imag} */,
  {32'hc09c1102, 32'hc04baa35} /* (14, 7, 20) {real, imag} */,
  {32'hbfbc3a9c, 32'hbfd236f6} /* (14, 7, 19) {real, imag} */,
  {32'h3e89ec60, 32'h408c9dd3} /* (14, 7, 18) {real, imag} */,
  {32'h3fcb2a18, 32'h3f0d4c5c} /* (14, 7, 17) {real, imag} */,
  {32'hbf9cf140, 32'hc0ddf545} /* (14, 7, 16) {real, imag} */,
  {32'h4036de9c, 32'hc0d9ccdc} /* (14, 7, 15) {real, imag} */,
  {32'hc1488a55, 32'hc045c41a} /* (14, 7, 14) {real, imag} */,
  {32'h41252d20, 32'h3e4186b0} /* (14, 7, 13) {real, imag} */,
  {32'hc149c301, 32'h410de97b} /* (14, 7, 12) {real, imag} */,
  {32'hc098a76b, 32'hc1c078b1} /* (14, 7, 11) {real, imag} */,
  {32'h4197b982, 32'h418d8eaa} /* (14, 7, 10) {real, imag} */,
  {32'hc1958e64, 32'hc036923a} /* (14, 7, 9) {real, imag} */,
  {32'hc1603b78, 32'hc21d8c69} /* (14, 7, 8) {real, imag} */,
  {32'hc0b09b9c, 32'hc0d7d499} /* (14, 7, 7) {real, imag} */,
  {32'h4190c4ec, 32'h41545875} /* (14, 7, 6) {real, imag} */,
  {32'h41a54073, 32'h41831469} /* (14, 7, 5) {real, imag} */,
  {32'h4165da20, 32'h4279425e} /* (14, 7, 4) {real, imag} */,
  {32'h41ba8384, 32'h41446da5} /* (14, 7, 3) {real, imag} */,
  {32'h41f9b7ef, 32'h41c33774} /* (14, 7, 2) {real, imag} */,
  {32'hc245538e, 32'hc2007ea7} /* (14, 7, 1) {real, imag} */,
  {32'hc1b81300, 32'hc130d0dc} /* (14, 7, 0) {real, imag} */,
  {32'h4198770c, 32'h41a8aae8} /* (14, 6, 31) {real, imag} */,
  {32'h42283904, 32'h41eabbbb} /* (14, 6, 30) {real, imag} */,
  {32'hc27690f1, 32'hc1dff7ae} /* (14, 6, 29) {real, imag} */,
  {32'h418b26ec, 32'h412d31c7} /* (14, 6, 28) {real, imag} */,
  {32'h41243aa8, 32'h42196b1b} /* (14, 6, 27) {real, imag} */,
  {32'h41b689e6, 32'hc0a2af40} /* (14, 6, 26) {real, imag} */,
  {32'hc1268a90, 32'hc1e076e3} /* (14, 6, 25) {real, imag} */,
  {32'hc07e78d8, 32'hbf22b120} /* (14, 6, 24) {real, imag} */,
  {32'h41875c58, 32'h41852b96} /* (14, 6, 23) {real, imag} */,
  {32'hc13a19b7, 32'hc1b07863} /* (14, 6, 22) {real, imag} */,
  {32'h40250462, 32'h41030e21} /* (14, 6, 21) {real, imag} */,
  {32'h415b79b2, 32'hc0527a62} /* (14, 6, 20) {real, imag} */,
  {32'h40d8266a, 32'hc0140ce8} /* (14, 6, 19) {real, imag} */,
  {32'hc0b6f3e0, 32'h401dddf2} /* (14, 6, 18) {real, imag} */,
  {32'h40aa947c, 32'hbffe50b2} /* (14, 6, 17) {real, imag} */,
  {32'hc0fedc6c, 32'hc09ebc74} /* (14, 6, 16) {real, imag} */,
  {32'h40e95710, 32'h41145d4a} /* (14, 6, 15) {real, imag} */,
  {32'hc08b1208, 32'hc0c153fd} /* (14, 6, 14) {real, imag} */,
  {32'h3faad948, 32'h4126cca0} /* (14, 6, 13) {real, imag} */,
  {32'hc0c939ab, 32'h403ae772} /* (14, 6, 12) {real, imag} */,
  {32'hc1667e62, 32'h405efc74} /* (14, 6, 11) {real, imag} */,
  {32'h3ff2a738, 32'h412d5ba6} /* (14, 6, 10) {real, imag} */,
  {32'hc22f6774, 32'h41986b22} /* (14, 6, 9) {real, imag} */,
  {32'hc14d6dc8, 32'hc1af868f} /* (14, 6, 8) {real, imag} */,
  {32'h4159c418, 32'hc18cfb8d} /* (14, 6, 7) {real, imag} */,
  {32'h40e25b8e, 32'h41f25d56} /* (14, 6, 6) {real, imag} */,
  {32'hc138d5ee, 32'hc16969f5} /* (14, 6, 5) {real, imag} */,
  {32'h41a95118, 32'hc1c0659a} /* (14, 6, 4) {real, imag} */,
  {32'h41c74096, 32'h41edce56} /* (14, 6, 3) {real, imag} */,
  {32'hc04f0968, 32'h415ceeca} /* (14, 6, 2) {real, imag} */,
  {32'h402fcb28, 32'hc2065b4c} /* (14, 6, 1) {real, imag} */,
  {32'h42326254, 32'hc1affb87} /* (14, 6, 0) {real, imag} */,
  {32'hc17c054f, 32'hc1923db0} /* (14, 5, 31) {real, imag} */,
  {32'hc00daf26, 32'hc252ce48} /* (14, 5, 30) {real, imag} */,
  {32'hc16c8bb6, 32'h41df3fb6} /* (14, 5, 29) {real, imag} */,
  {32'h422e80c8, 32'hc12bfde2} /* (14, 5, 28) {real, imag} */,
  {32'hc21244a9, 32'h40ea2874} /* (14, 5, 27) {real, imag} */,
  {32'hbfc2d3e4, 32'h41b7da92} /* (14, 5, 26) {real, imag} */,
  {32'h41c129fa, 32'hc19b3b07} /* (14, 5, 25) {real, imag} */,
  {32'hc182091e, 32'h421194db} /* (14, 5, 24) {real, imag} */,
  {32'h417ad287, 32'hc120bc02} /* (14, 5, 23) {real, imag} */,
  {32'hc1b48aca, 32'hc15b2828} /* (14, 5, 22) {real, imag} */,
  {32'hc16da5c3, 32'h3f9d030c} /* (14, 5, 21) {real, imag} */,
  {32'hc1404665, 32'h40e1dcb8} /* (14, 5, 20) {real, imag} */,
  {32'h410bbe48, 32'h4104d81f} /* (14, 5, 19) {real, imag} */,
  {32'hc13fa938, 32'h41238731} /* (14, 5, 18) {real, imag} */,
  {32'hc1830dea, 32'hbe14eb40} /* (14, 5, 17) {real, imag} */,
  {32'h4140f604, 32'h4111016c} /* (14, 5, 16) {real, imag} */,
  {32'hc0f91d98, 32'h40bf8f8e} /* (14, 5, 15) {real, imag} */,
  {32'h413975b4, 32'h40d63b7a} /* (14, 5, 14) {real, imag} */,
  {32'h41019b88, 32'hc0b2261a} /* (14, 5, 13) {real, imag} */,
  {32'h413cdec1, 32'h40f062c0} /* (14, 5, 12) {real, imag} */,
  {32'h413d7d1b, 32'hbfa2b864} /* (14, 5, 11) {real, imag} */,
  {32'hc0a950f6, 32'h408f9d50} /* (14, 5, 10) {real, imag} */,
  {32'h41822f90, 32'hc237ca3c} /* (14, 5, 9) {real, imag} */,
  {32'hc115bfdc, 32'h4197aca6} /* (14, 5, 8) {real, imag} */,
  {32'hc02ff38c, 32'hc13e7d42} /* (14, 5, 7) {real, imag} */,
  {32'hc0b96dcb, 32'h4159a2a0} /* (14, 5, 6) {real, imag} */,
  {32'h421f2ad5, 32'h41c3f95b} /* (14, 5, 5) {real, imag} */,
  {32'h410a968e, 32'h42213374} /* (14, 5, 4) {real, imag} */,
  {32'hbf39f4a8, 32'hc1ae8874} /* (14, 5, 3) {real, imag} */,
  {32'hc12a2348, 32'hc1276e1e} /* (14, 5, 2) {real, imag} */,
  {32'hc05f5464, 32'h4297fee4} /* (14, 5, 1) {real, imag} */,
  {32'h429d92f8, 32'h42ab31da} /* (14, 5, 0) {real, imag} */,
  {32'hc235c1bc, 32'hc26b7f31} /* (14, 4, 31) {real, imag} */,
  {32'h41a667bb, 32'hc212d76a} /* (14, 4, 30) {real, imag} */,
  {32'h41862c59, 32'hc24a711b} /* (14, 4, 29) {real, imag} */,
  {32'h4035b848, 32'h41149d9e} /* (14, 4, 28) {real, imag} */,
  {32'hc17bdaba, 32'hc1fdb769} /* (14, 4, 27) {real, imag} */,
  {32'h414a3c75, 32'hbe1c2b20} /* (14, 4, 26) {real, imag} */,
  {32'h4135c979, 32'hc1886524} /* (14, 4, 25) {real, imag} */,
  {32'h418c37e0, 32'hc15dc794} /* (14, 4, 24) {real, imag} */,
  {32'h412b2eb7, 32'hbeeb5a00} /* (14, 4, 23) {real, imag} */,
  {32'h3f521230, 32'h41812abc} /* (14, 4, 22) {real, imag} */,
  {32'hc0550290, 32'hc0e3acb4} /* (14, 4, 21) {real, imag} */,
  {32'h41a9f6f7, 32'h414e9474} /* (14, 4, 20) {real, imag} */,
  {32'hc0dea28d, 32'h419d7614} /* (14, 4, 19) {real, imag} */,
  {32'h40b8b3cf, 32'h415237be} /* (14, 4, 18) {real, imag} */,
  {32'hbf03b9a0, 32'h3f210c00} /* (14, 4, 17) {real, imag} */,
  {32'hbfe14e94, 32'hbf8d3dd0} /* (14, 4, 16) {real, imag} */,
  {32'h40e4d764, 32'hbf85d7a0} /* (14, 4, 15) {real, imag} */,
  {32'hc04bc92e, 32'h40224948} /* (14, 4, 14) {real, imag} */,
  {32'hc088ab9b, 32'h411af58a} /* (14, 4, 13) {real, imag} */,
  {32'hc099b834, 32'h413bd900} /* (14, 4, 12) {real, imag} */,
  {32'hc1d93d9c, 32'hc18cb16d} /* (14, 4, 11) {real, imag} */,
  {32'h41b51b5e, 32'h400010fc} /* (14, 4, 10) {real, imag} */,
  {32'hc114c6a7, 32'h40020a30} /* (14, 4, 9) {real, imag} */,
  {32'h404718aa, 32'h401021f2} /* (14, 4, 8) {real, imag} */,
  {32'hc18dc2d4, 32'h41a48b2e} /* (14, 4, 7) {real, imag} */,
  {32'hc1156b5b, 32'hbfc0c114} /* (14, 4, 6) {real, imag} */,
  {32'h421045c0, 32'hc1e4d5dd} /* (14, 4, 5) {real, imag} */,
  {32'h4095065a, 32'hc0e0700b} /* (14, 4, 4) {real, imag} */,
  {32'h4152bb66, 32'h40ab2f98} /* (14, 4, 3) {real, imag} */,
  {32'h41749a6e, 32'h41539620} /* (14, 4, 2) {real, imag} */,
  {32'hc2ccb1ee, 32'h423c2b47} /* (14, 4, 1) {real, imag} */,
  {32'h4135d7b4, 32'hc1c223d9} /* (14, 4, 0) {real, imag} */,
  {32'h4264313c, 32'hc2338894} /* (14, 3, 31) {real, imag} */,
  {32'h41e4b1d6, 32'h4115307d} /* (14, 3, 30) {real, imag} */,
  {32'hc293c3d2, 32'h42395aed} /* (14, 3, 29) {real, imag} */,
  {32'hc1868897, 32'hc135ea09} /* (14, 3, 28) {real, imag} */,
  {32'hbd527600, 32'hc215d4e0} /* (14, 3, 27) {real, imag} */,
  {32'hbfe00630, 32'hc1954ee0} /* (14, 3, 26) {real, imag} */,
  {32'h40f38e36, 32'h4240a902} /* (14, 3, 25) {real, imag} */,
  {32'h416d7425, 32'hc076959c} /* (14, 3, 24) {real, imag} */,
  {32'h41c2ca56, 32'hc1742748} /* (14, 3, 23) {real, imag} */,
  {32'hc0d8e278, 32'h41338db8} /* (14, 3, 22) {real, imag} */,
  {32'h41547a12, 32'hc15b8e1a} /* (14, 3, 21) {real, imag} */,
  {32'hbf065840, 32'hc10d2ee3} /* (14, 3, 20) {real, imag} */,
  {32'h40b208b4, 32'hc09d2976} /* (14, 3, 19) {real, imag} */,
  {32'hc130f698, 32'h414f65b7} /* (14, 3, 18) {real, imag} */,
  {32'hc130b5f7, 32'hc0c7f59d} /* (14, 3, 17) {real, imag} */,
  {32'h414d3a92, 32'h3f284478} /* (14, 3, 16) {real, imag} */,
  {32'h41920f2c, 32'h40d64475} /* (14, 3, 15) {real, imag} */,
  {32'hc0fe5cbc, 32'hc0319164} /* (14, 3, 14) {real, imag} */,
  {32'hc01e4bc8, 32'h41556499} /* (14, 3, 13) {real, imag} */,
  {32'hc15d2b40, 32'h41420f43} /* (14, 3, 12) {real, imag} */,
  {32'hc127b534, 32'h40751538} /* (14, 3, 11) {real, imag} */,
  {32'hbd2df5c0, 32'hc1ae9cbe} /* (14, 3, 10) {real, imag} */,
  {32'hc17e2874, 32'h40e2e464} /* (14, 3, 9) {real, imag} */,
  {32'h4135d0af, 32'h3eb9c8c0} /* (14, 3, 8) {real, imag} */,
  {32'h411d4d69, 32'hc17009e0} /* (14, 3, 7) {real, imag} */,
  {32'h40dd5290, 32'h414d6e0c} /* (14, 3, 6) {real, imag} */,
  {32'h421c1090, 32'hc161ac36} /* (14, 3, 5) {real, imag} */,
  {32'h424e69c4, 32'hc1ccbb0c} /* (14, 3, 4) {real, imag} */,
  {32'h40115cd0, 32'hc203e9af} /* (14, 3, 3) {real, imag} */,
  {32'hc07538ac, 32'hc02c499b} /* (14, 3, 2) {real, imag} */,
  {32'hc1a01039, 32'hc1d4b34f} /* (14, 3, 1) {real, imag} */,
  {32'h41a1dd25, 32'hc10fc854} /* (14, 3, 0) {real, imag} */,
  {32'h432ab3b5, 32'h41a12e7a} /* (14, 2, 31) {real, imag} */,
  {32'hc305758c, 32'h4295ea05} /* (14, 2, 30) {real, imag} */,
  {32'h419d49c4, 32'hc2481238} /* (14, 2, 29) {real, imag} */,
  {32'h41a75b84, 32'hc1b6230d} /* (14, 2, 28) {real, imag} */,
  {32'h4166e5e6, 32'h422f26b3} /* (14, 2, 27) {real, imag} */,
  {32'h422e3f50, 32'hc0aa51e7} /* (14, 2, 26) {real, imag} */,
  {32'hc1ce443f, 32'hc0f5fd56} /* (14, 2, 25) {real, imag} */,
  {32'hc1b18d9a, 32'h4263d807} /* (14, 2, 24) {real, imag} */,
  {32'h3f0a7fa0, 32'h4145b349} /* (14, 2, 23) {real, imag} */,
  {32'h41b0b3e0, 32'h3f836a4c} /* (14, 2, 22) {real, imag} */,
  {32'hc1701998, 32'h41987487} /* (14, 2, 21) {real, imag} */,
  {32'hbfc85290, 32'hbeead898} /* (14, 2, 20) {real, imag} */,
  {32'h4038e156, 32'hc07d7ba4} /* (14, 2, 19) {real, imag} */,
  {32'hc0f7707c, 32'hc18cc8a6} /* (14, 2, 18) {real, imag} */,
  {32'h40bf4674, 32'hc02b98de} /* (14, 2, 17) {real, imag} */,
  {32'h4100e620, 32'hbf5cf280} /* (14, 2, 16) {real, imag} */,
  {32'h41355f66, 32'h40e3ed7f} /* (14, 2, 15) {real, imag} */,
  {32'hc12698b2, 32'hc18c3c0a} /* (14, 2, 14) {real, imag} */,
  {32'h402ef99a, 32'h41cbacfc} /* (14, 2, 13) {real, imag} */,
  {32'hc1ce539f, 32'hc082370a} /* (14, 2, 12) {real, imag} */,
  {32'h41a4aaf2, 32'hc1b9f1ed} /* (14, 2, 11) {real, imag} */,
  {32'hc1de18da, 32'h41426842} /* (14, 2, 10) {real, imag} */,
  {32'h41cae17b, 32'h4133e1d5} /* (14, 2, 9) {real, imag} */,
  {32'h418f62fe, 32'hbfe509e0} /* (14, 2, 8) {real, imag} */,
  {32'h41ba03a7, 32'h3e857218} /* (14, 2, 7) {real, imag} */,
  {32'h411f98c4, 32'hc18796ba} /* (14, 2, 6) {real, imag} */,
  {32'h4281f57b, 32'hc21bea8d} /* (14, 2, 5) {real, imag} */,
  {32'h4184e2e4, 32'h4188640d} /* (14, 2, 4) {real, imag} */,
  {32'hbbbfa000, 32'h42250fc0} /* (14, 2, 3) {real, imag} */,
  {32'hc1b249bc, 32'h424bb07a} /* (14, 2, 2) {real, imag} */,
  {32'h422c118c, 32'h40aac367} /* (14, 2, 1) {real, imag} */,
  {32'h429b45a9, 32'h4196b0bf} /* (14, 2, 0) {real, imag} */,
  {32'hc2fca6ae, 32'h42a6307a} /* (14, 1, 31) {real, imag} */,
  {32'h42a94d2c, 32'hc1f41075} /* (14, 1, 30) {real, imag} */,
  {32'h41427370, 32'hc20126ed} /* (14, 1, 29) {real, imag} */,
  {32'hc1d93ad8, 32'hc223eac6} /* (14, 1, 28) {real, imag} */,
  {32'h42400a93, 32'hc28e044c} /* (14, 1, 27) {real, imag} */,
  {32'h4122a668, 32'hbf69aaf0} /* (14, 1, 26) {real, imag} */,
  {32'h41b35e80, 32'h41cffa1e} /* (14, 1, 25) {real, imag} */,
  {32'hc253fa28, 32'h41feb2c0} /* (14, 1, 24) {real, imag} */,
  {32'h413ccc13, 32'hc1c2ca28} /* (14, 1, 23) {real, imag} */,
  {32'h40f02dc6, 32'h4125e043} /* (14, 1, 22) {real, imag} */,
  {32'h4176d9b6, 32'h41481a2f} /* (14, 1, 21) {real, imag} */,
  {32'hc15f4d9b, 32'hc10c39c0} /* (14, 1, 20) {real, imag} */,
  {32'h408d2308, 32'hc0246eb8} /* (14, 1, 19) {real, imag} */,
  {32'h40540f80, 32'hbf146198} /* (14, 1, 18) {real, imag} */,
  {32'h3fefc2ac, 32'hc1923a07} /* (14, 1, 17) {real, imag} */,
  {32'h3eb90200, 32'hbf402c00} /* (14, 1, 16) {real, imag} */,
  {32'hc1511036, 32'hc1739426} /* (14, 1, 15) {real, imag} */,
  {32'hc13840c8, 32'h41428f44} /* (14, 1, 14) {real, imag} */,
  {32'h4177ca02, 32'hc0e9dd50} /* (14, 1, 13) {real, imag} */,
  {32'hbeaec420, 32'hc0c78ee0} /* (14, 1, 12) {real, imag} */,
  {32'h413f5fee, 32'hc10cc58b} /* (14, 1, 11) {real, imag} */,
  {32'h4154adc1, 32'h42007656} /* (14, 1, 10) {real, imag} */,
  {32'h4220e4ac, 32'h40d088b6} /* (14, 1, 9) {real, imag} */,
  {32'hc102a49a, 32'hc13c3d78} /* (14, 1, 8) {real, imag} */,
  {32'h419175fa, 32'h3dc64880} /* (14, 1, 7) {real, imag} */,
  {32'hc13195fc, 32'hc1fdc886} /* (14, 1, 6) {real, imag} */,
  {32'hc0b50de0, 32'h40b53fd8} /* (14, 1, 5) {real, imag} */,
  {32'hc1f99f92, 32'h42502b8e} /* (14, 1, 4) {real, imag} */,
  {32'hc1339686, 32'h4154872b} /* (14, 1, 3) {real, imag} */,
  {32'h42da18ac, 32'h40c5013c} /* (14, 1, 2) {real, imag} */,
  {32'hc32b7951, 32'hc29f7b0e} /* (14, 1, 1) {real, imag} */,
  {32'hc2e06979, 32'h4156e893} /* (14, 1, 0) {real, imag} */,
  {32'hc1cb43bc, 32'h42311036} /* (14, 0, 31) {real, imag} */,
  {32'h416c6190, 32'h41ce87e6} /* (14, 0, 30) {real, imag} */,
  {32'h41a2559a, 32'hc23155fa} /* (14, 0, 29) {real, imag} */,
  {32'h426446d7, 32'hc10cf8cf} /* (14, 0, 28) {real, imag} */,
  {32'h42269f66, 32'hbf6ee2b0} /* (14, 0, 27) {real, imag} */,
  {32'hc236c1fa, 32'h426b7280} /* (14, 0, 26) {real, imag} */,
  {32'h4210f4f5, 32'h42638933} /* (14, 0, 25) {real, imag} */,
  {32'hc1f0da00, 32'hc17bda82} /* (14, 0, 24) {real, imag} */,
  {32'h42061494, 32'hc1bc802e} /* (14, 0, 23) {real, imag} */,
  {32'h40233ace, 32'h4112b67c} /* (14, 0, 22) {real, imag} */,
  {32'h4126328a, 32'hc098fa11} /* (14, 0, 21) {real, imag} */,
  {32'hbe447bc0, 32'h3f9342ac} /* (14, 0, 20) {real, imag} */,
  {32'h3f08d618, 32'h4128d9af} /* (14, 0, 19) {real, imag} */,
  {32'hc1018854, 32'hc028dd4c} /* (14, 0, 18) {real, imag} */,
  {32'h405a9538, 32'h3f3d2c00} /* (14, 0, 17) {real, imag} */,
  {32'hc128eae2, 32'hc10d94e6} /* (14, 0, 16) {real, imag} */,
  {32'h40dff56c, 32'h41a70e08} /* (14, 0, 15) {real, imag} */,
  {32'h409590d8, 32'h40a9458a} /* (14, 0, 14) {real, imag} */,
  {32'hc11b2b86, 32'h40d8fc5a} /* (14, 0, 13) {real, imag} */,
  {32'h4104f96d, 32'h3ecf3a80} /* (14, 0, 12) {real, imag} */,
  {32'h404da090, 32'h4196d160} /* (14, 0, 11) {real, imag} */,
  {32'hc1466030, 32'h41c09cb0} /* (14, 0, 10) {real, imag} */,
  {32'h418d1bd1, 32'hc26f3701} /* (14, 0, 9) {real, imag} */,
  {32'hc1ccfba0, 32'h407500c8} /* (14, 0, 8) {real, imag} */,
  {32'hc206919f, 32'hbfca0660} /* (14, 0, 7) {real, imag} */,
  {32'hc1a6c093, 32'hc161dc0e} /* (14, 0, 6) {real, imag} */,
  {32'h3f98dac0, 32'h4081c35c} /* (14, 0, 5) {real, imag} */,
  {32'hc1de15b2, 32'h3f8b99a6} /* (14, 0, 4) {real, imag} */,
  {32'hc263bdd5, 32'hc143442a} /* (14, 0, 3) {real, imag} */,
  {32'h4294e903, 32'h41a95ec6} /* (14, 0, 2) {real, imag} */,
  {32'hc21e3d8e, 32'hc2b34091} /* (14, 0, 1) {real, imag} */,
  {32'hc24937ec, 32'h42330ea4} /* (14, 0, 0) {real, imag} */,
  {32'hc101ef12, 32'hc2090c5b} /* (13, 31, 31) {real, imag} */,
  {32'hc1a0f614, 32'hc03fce4d} /* (13, 31, 30) {real, imag} */,
  {32'hc14d14c6, 32'h41cf42ce} /* (13, 31, 29) {real, imag} */,
  {32'h4259ef19, 32'hc13432fa} /* (13, 31, 28) {real, imag} */,
  {32'hc2690222, 32'h41b4fedd} /* (13, 31, 27) {real, imag} */,
  {32'h3f068258, 32'hc1f26d51} /* (13, 31, 26) {real, imag} */,
  {32'hc1d9b5e4, 32'h40b97626} /* (13, 31, 25) {real, imag} */,
  {32'h42052297, 32'hc1ddae50} /* (13, 31, 24) {real, imag} */,
  {32'hc1a3d024, 32'hc17459ac} /* (13, 31, 23) {real, imag} */,
  {32'h4130fa24, 32'hc1deaddd} /* (13, 31, 22) {real, imag} */,
  {32'h40df4191, 32'h42303ee6} /* (13, 31, 21) {real, imag} */,
  {32'hc0d897a0, 32'h416f81b4} /* (13, 31, 20) {real, imag} */,
  {32'hc1a2a7c8, 32'h411146e8} /* (13, 31, 19) {real, imag} */,
  {32'hbf08c870, 32'hc143df64} /* (13, 31, 18) {real, imag} */,
  {32'h40f4dce4, 32'h3fd96644} /* (13, 31, 17) {real, imag} */,
  {32'hbff6f1b8, 32'hc0bf2f66} /* (13, 31, 16) {real, imag} */,
  {32'h41295e0a, 32'hc095d2b5} /* (13, 31, 15) {real, imag} */,
  {32'h3fb69ae8, 32'h40d4d927} /* (13, 31, 14) {real, imag} */,
  {32'hbea79680, 32'hc0201e70} /* (13, 31, 13) {real, imag} */,
  {32'h4195d5f2, 32'hc195dc0c} /* (13, 31, 12) {real, imag} */,
  {32'hc18041ba, 32'hc1912946} /* (13, 31, 11) {real, imag} */,
  {32'h3f731a48, 32'h42004812} /* (13, 31, 10) {real, imag} */,
  {32'hc0e56e6a, 32'h4252e547} /* (13, 31, 9) {real, imag} */,
  {32'hbfc14b38, 32'h40d9daa6} /* (13, 31, 8) {real, imag} */,
  {32'hc1ba47fa, 32'h4084b456} /* (13, 31, 7) {real, imag} */,
  {32'h417ab1de, 32'hc28b91f6} /* (13, 31, 6) {real, imag} */,
  {32'h41d93ba4, 32'hc28a4640} /* (13, 31, 5) {real, imag} */,
  {32'h408541d0, 32'hc18cebdf} /* (13, 31, 4) {real, imag} */,
  {32'hc27412fe, 32'h4202defc} /* (13, 31, 3) {real, imag} */,
  {32'h42441bee, 32'hc0e06380} /* (13, 31, 2) {real, imag} */,
  {32'h418d7f79, 32'hc1378f74} /* (13, 31, 1) {real, imag} */,
  {32'h419db050, 32'h41890f24} /* (13, 31, 0) {real, imag} */,
  {32'hc1e32800, 32'hc253c18f} /* (13, 30, 31) {real, imag} */,
  {32'h41ca372d, 32'h420ccc22} /* (13, 30, 30) {real, imag} */,
  {32'hc1d9ceca, 32'hbf4f58c0} /* (13, 30, 29) {real, imag} */,
  {32'h4116ed59, 32'hc1a09145} /* (13, 30, 28) {real, imag} */,
  {32'h41807e2b, 32'h400ec270} /* (13, 30, 27) {real, imag} */,
  {32'hc0fc6720, 32'h42212537} /* (13, 30, 26) {real, imag} */,
  {32'h403df698, 32'hc21b541b} /* (13, 30, 25) {real, imag} */,
  {32'hc06c0ab0, 32'h3fbf1a60} /* (13, 30, 24) {real, imag} */,
  {32'h4149466a, 32'hc16e3762} /* (13, 30, 23) {real, imag} */,
  {32'h41dc41dd, 32'h418f5b45} /* (13, 30, 22) {real, imag} */,
  {32'hc0af60a8, 32'h405bdfd2} /* (13, 30, 21) {real, imag} */,
  {32'h41b9c572, 32'h40ff76e6} /* (13, 30, 20) {real, imag} */,
  {32'h3ec43170, 32'h41571e53} /* (13, 30, 19) {real, imag} */,
  {32'hc0fab378, 32'h412b41be} /* (13, 30, 18) {real, imag} */,
  {32'h4091415e, 32'hc071345c} /* (13, 30, 17) {real, imag} */,
  {32'hc12d0de2, 32'h41870bcc} /* (13, 30, 16) {real, imag} */,
  {32'h408792f6, 32'h3ffe2c78} /* (13, 30, 15) {real, imag} */,
  {32'h3fe1f960, 32'h403e5d18} /* (13, 30, 14) {real, imag} */,
  {32'hc156fb6e, 32'hc0f775f6} /* (13, 30, 13) {real, imag} */,
  {32'hc09d6aee, 32'hc12f4319} /* (13, 30, 12) {real, imag} */,
  {32'h41ff2a66, 32'h418e6562} /* (13, 30, 11) {real, imag} */,
  {32'h41f6df79, 32'h4023e720} /* (13, 30, 10) {real, imag} */,
  {32'hc172fb24, 32'h42052936} /* (13, 30, 9) {real, imag} */,
  {32'h420910a9, 32'h41f9a41a} /* (13, 30, 8) {real, imag} */,
  {32'hc1b651fa, 32'hc2792f49} /* (13, 30, 7) {real, imag} */,
  {32'hc28b9b98, 32'hc09ec968} /* (13, 30, 6) {real, imag} */,
  {32'hc21c8a00, 32'h4211e4a9} /* (13, 30, 5) {real, imag} */,
  {32'hc1a8ed1a, 32'h4219dcca} /* (13, 30, 4) {real, imag} */,
  {32'h419376b6, 32'h4234a153} /* (13, 30, 3) {real, imag} */,
  {32'h418b6715, 32'hc2a4f534} /* (13, 30, 2) {real, imag} */,
  {32'h414b0825, 32'hc1c0255a} /* (13, 30, 1) {real, imag} */,
  {32'hc21d3e66, 32'hc1900828} /* (13, 30, 0) {real, imag} */,
  {32'h422a0944, 32'h41e78e64} /* (13, 29, 31) {real, imag} */,
  {32'hc2351a62, 32'hc18b51f8} /* (13, 29, 30) {real, imag} */,
  {32'hc1f09cce, 32'hbf6989e0} /* (13, 29, 29) {real, imag} */,
  {32'hc2307a30, 32'hc2204b78} /* (13, 29, 28) {real, imag} */,
  {32'h3fe1cf50, 32'hc0e146e7} /* (13, 29, 27) {real, imag} */,
  {32'h42a57790, 32'h418dde0d} /* (13, 29, 26) {real, imag} */,
  {32'hc163588a, 32'h4160436d} /* (13, 29, 25) {real, imag} */,
  {32'h420b1ea9, 32'hc20aaf8b} /* (13, 29, 24) {real, imag} */,
  {32'h4092bf56, 32'h40a802ae} /* (13, 29, 23) {real, imag} */,
  {32'h41b294c9, 32'h40a4803c} /* (13, 29, 22) {real, imag} */,
  {32'hc1bf9a07, 32'hc0ab6b55} /* (13, 29, 21) {real, imag} */,
  {32'h41bba3a0, 32'h41c26e7f} /* (13, 29, 20) {real, imag} */,
  {32'h411b65aa, 32'hc1bc544b} /* (13, 29, 19) {real, imag} */,
  {32'hbfbfc618, 32'h41bd75c1} /* (13, 29, 18) {real, imag} */,
  {32'h3f01af90, 32'h414c8338} /* (13, 29, 17) {real, imag} */,
  {32'hc13b332b, 32'h415e914a} /* (13, 29, 16) {real, imag} */,
  {32'hc0da2e52, 32'h4141efa8} /* (13, 29, 15) {real, imag} */,
  {32'hc0cda5de, 32'hc1240ca6} /* (13, 29, 14) {real, imag} */,
  {32'hc09aa6d3, 32'hc1834fc5} /* (13, 29, 13) {real, imag} */,
  {32'h3f952c20, 32'h412c8b1a} /* (13, 29, 12) {real, imag} */,
  {32'hc1e0f7c1, 32'hc1a00bc0} /* (13, 29, 11) {real, imag} */,
  {32'hc1c5bdb7, 32'hc1cb977d} /* (13, 29, 10) {real, imag} */,
  {32'h41051e08, 32'hc15dec75} /* (13, 29, 9) {real, imag} */,
  {32'hc1b1cd64, 32'hc11a33b4} /* (13, 29, 8) {real, imag} */,
  {32'h41a014d5, 32'hc1b29730} /* (13, 29, 7) {real, imag} */,
  {32'h414511b0, 32'hc19b9abf} /* (13, 29, 6) {real, imag} */,
  {32'hc207326c, 32'hc1982eb1} /* (13, 29, 5) {real, imag} */,
  {32'h40d67384, 32'h423859fc} /* (13, 29, 4) {real, imag} */,
  {32'hc01f3a80, 32'h426a2548} /* (13, 29, 3) {real, imag} */,
  {32'h4181fbee, 32'hc26aa7a0} /* (13, 29, 2) {real, imag} */,
  {32'hbfcfbe80, 32'h4244a4bc} /* (13, 29, 1) {real, imag} */,
  {32'h4113e865, 32'h41d2ce63} /* (13, 29, 0) {real, imag} */,
  {32'hbf49d130, 32'hc2a90e1a} /* (13, 28, 31) {real, imag} */,
  {32'h42118777, 32'h42a80a86} /* (13, 28, 30) {real, imag} */,
  {32'hc200536f, 32'hc202570b} /* (13, 28, 29) {real, imag} */,
  {32'h4166e09a, 32'h420343c2} /* (13, 28, 28) {real, imag} */,
  {32'hc181a909, 32'hc18f66c0} /* (13, 28, 27) {real, imag} */,
  {32'hc1d0d1be, 32'h41609ac7} /* (13, 28, 26) {real, imag} */,
  {32'h406d2eb0, 32'hc14f3666} /* (13, 28, 25) {real, imag} */,
  {32'h4105875b, 32'hc119e130} /* (13, 28, 24) {real, imag} */,
  {32'hbf6a8d70, 32'h41e1b676} /* (13, 28, 23) {real, imag} */,
  {32'h416ad018, 32'h404a7228} /* (13, 28, 22) {real, imag} */,
  {32'hc1c0ed5e, 32'hc1b8a550} /* (13, 28, 21) {real, imag} */,
  {32'hc1283424, 32'hc1a5d4b2} /* (13, 28, 20) {real, imag} */,
  {32'hbf83a448, 32'hc1217ab4} /* (13, 28, 19) {real, imag} */,
  {32'h411bfdc1, 32'hc0e3a310} /* (13, 28, 18) {real, imag} */,
  {32'hc13967a5, 32'hc160c815} /* (13, 28, 17) {real, imag} */,
  {32'h40b6ed1c, 32'hc0cfb836} /* (13, 28, 16) {real, imag} */,
  {32'h40c40faa, 32'h40d5ede6} /* (13, 28, 15) {real, imag} */,
  {32'hc1037d2f, 32'hc1997fa4} /* (13, 28, 14) {real, imag} */,
  {32'hc1bdd478, 32'hc1904bbf} /* (13, 28, 13) {real, imag} */,
  {32'hc1faffb0, 32'hbf91c868} /* (13, 28, 12) {real, imag} */,
  {32'h416dd658, 32'h41860b3c} /* (13, 28, 11) {real, imag} */,
  {32'h41f24db4, 32'h41d2ee66} /* (13, 28, 10) {real, imag} */,
  {32'hc1e0bf5c, 32'h40e5970a} /* (13, 28, 9) {real, imag} */,
  {32'h41bc8c54, 32'h420e1e16} /* (13, 28, 8) {real, imag} */,
  {32'h425211bb, 32'h41b78175} /* (13, 28, 7) {real, imag} */,
  {32'hc199210a, 32'hc2219f7a} /* (13, 28, 6) {real, imag} */,
  {32'h40324f56, 32'hbffa7ed8} /* (13, 28, 5) {real, imag} */,
  {32'h41b01521, 32'hc04cfd84} /* (13, 28, 4) {real, imag} */,
  {32'h3fb93468, 32'hc1bcc8ea} /* (13, 28, 3) {real, imag} */,
  {32'hc29fcda6, 32'hc239402f} /* (13, 28, 2) {real, imag} */,
  {32'h418233fa, 32'h41db9452} /* (13, 28, 1) {real, imag} */,
  {32'hc2504e6a, 32'h4038f1bc} /* (13, 28, 0) {real, imag} */,
  {32'h41562475, 32'hc2651bad} /* (13, 27, 31) {real, imag} */,
  {32'h40c6cecc, 32'h3fc1ac70} /* (13, 27, 30) {real, imag} */,
  {32'h42557809, 32'h41a0e9ef} /* (13, 27, 29) {real, imag} */,
  {32'hc21ab6d2, 32'hc18f4e54} /* (13, 27, 28) {real, imag} */,
  {32'h42431334, 32'hc211f4c9} /* (13, 27, 27) {real, imag} */,
  {32'h40b19d38, 32'h421fa36a} /* (13, 27, 26) {real, imag} */,
  {32'hc23d0bb4, 32'hc0235ea4} /* (13, 27, 25) {real, imag} */,
  {32'hc259efc8, 32'hc145050e} /* (13, 27, 24) {real, imag} */,
  {32'h41fe3029, 32'hbf6c68c0} /* (13, 27, 23) {real, imag} */,
  {32'h41ffa662, 32'h414b497a} /* (13, 27, 22) {real, imag} */,
  {32'h4094ff70, 32'h412ee958} /* (13, 27, 21) {real, imag} */,
  {32'h40526ede, 32'h40f4b422} /* (13, 27, 20) {real, imag} */,
  {32'h402543b0, 32'hc11e1ee6} /* (13, 27, 19) {real, imag} */,
  {32'hc164c26a, 32'hc0870cb8} /* (13, 27, 18) {real, imag} */,
  {32'hc07ef2b8, 32'hc0390fd8} /* (13, 27, 17) {real, imag} */,
  {32'h40496dd8, 32'h41152ad4} /* (13, 27, 16) {real, imag} */,
  {32'h40998be4, 32'h418c3e8f} /* (13, 27, 15) {real, imag} */,
  {32'hc17a555e, 32'h41a8d2e4} /* (13, 27, 14) {real, imag} */,
  {32'hc0870a60, 32'h405c7bb0} /* (13, 27, 13) {real, imag} */,
  {32'hc04c811e, 32'h413b5bf7} /* (13, 27, 12) {real, imag} */,
  {32'h41e446aa, 32'h3e334380} /* (13, 27, 11) {real, imag} */,
  {32'h3facefa0, 32'h41e2d8c3} /* (13, 27, 10) {real, imag} */,
  {32'hc2075444, 32'hc0f346ca} /* (13, 27, 9) {real, imag} */,
  {32'hc1e738bf, 32'hc1b41b4d} /* (13, 27, 8) {real, imag} */,
  {32'hc1d09d97, 32'hc0c5056c} /* (13, 27, 7) {real, imag} */,
  {32'h420c3d3d, 32'h4148df9a} /* (13, 27, 6) {real, imag} */,
  {32'hc22b4d18, 32'hc1baef4a} /* (13, 27, 5) {real, imag} */,
  {32'hbf4ffb00, 32'hc2902283} /* (13, 27, 4) {real, imag} */,
  {32'hc0cc5b40, 32'h41878785} /* (13, 27, 3) {real, imag} */,
  {32'hc2050bee, 32'h418b97d3} /* (13, 27, 2) {real, imag} */,
  {32'h41618fe5, 32'h4218e667} /* (13, 27, 1) {real, imag} */,
  {32'hc22349c8, 32'hc1db2dc6} /* (13, 27, 0) {real, imag} */,
  {32'h4233a089, 32'h427a79c4} /* (13, 26, 31) {real, imag} */,
  {32'hc203f322, 32'h41bb2a56} /* (13, 26, 30) {real, imag} */,
  {32'hc1d172ca, 32'h41e144d6} /* (13, 26, 29) {real, imag} */,
  {32'h41ae122a, 32'h4100c694} /* (13, 26, 28) {real, imag} */,
  {32'h418e9e95, 32'h41f68cff} /* (13, 26, 27) {real, imag} */,
  {32'hc215ea8e, 32'hc0267f4a} /* (13, 26, 26) {real, imag} */,
  {32'hc222e1b6, 32'h411765c1} /* (13, 26, 25) {real, imag} */,
  {32'hc075b47e, 32'hc14ddacd} /* (13, 26, 24) {real, imag} */,
  {32'hc21adefe, 32'h419bf8d4} /* (13, 26, 23) {real, imag} */,
  {32'hc0b1e8a4, 32'h40b61073} /* (13, 26, 22) {real, imag} */,
  {32'h41523b24, 32'hc18ddf3e} /* (13, 26, 21) {real, imag} */,
  {32'h4143e3c4, 32'hc0ecd832} /* (13, 26, 20) {real, imag} */,
  {32'h4058ec67, 32'hc0d19c5a} /* (13, 26, 19) {real, imag} */,
  {32'hc1c73388, 32'hc169ff72} /* (13, 26, 18) {real, imag} */,
  {32'hc0cf3572, 32'h411d7df8} /* (13, 26, 17) {real, imag} */,
  {32'h4050dd28, 32'hc14ddcd0} /* (13, 26, 16) {real, imag} */,
  {32'h4078f1e4, 32'hc1401b3c} /* (13, 26, 15) {real, imag} */,
  {32'h40b0d030, 32'hc119f39e} /* (13, 26, 14) {real, imag} */,
  {32'hc0bf06ac, 32'h409d932e} /* (13, 26, 13) {real, imag} */,
  {32'h40b0e3c8, 32'h3f0c41a0} /* (13, 26, 12) {real, imag} */,
  {32'h414335ce, 32'hc0c7e742} /* (13, 26, 11) {real, imag} */,
  {32'hc1cdb85d, 32'hc0558f0a} /* (13, 26, 10) {real, imag} */,
  {32'h4186e14f, 32'hc192b7ba} /* (13, 26, 9) {real, imag} */,
  {32'h3f561558, 32'h41fbc8e8} /* (13, 26, 8) {real, imag} */,
  {32'h414a942e, 32'hc20e62cb} /* (13, 26, 7) {real, imag} */,
  {32'hc1b4eb07, 32'h418bc687} /* (13, 26, 6) {real, imag} */,
  {32'h40c8b1f8, 32'hc1136b5a} /* (13, 26, 5) {real, imag} */,
  {32'hc1495c67, 32'hc1a61684} /* (13, 26, 4) {real, imag} */,
  {32'h421e2fb1, 32'h41cddde2} /* (13, 26, 3) {real, imag} */,
  {32'h4157d0be, 32'h4166d754} /* (13, 26, 2) {real, imag} */,
  {32'h42636e3d, 32'h426521cc} /* (13, 26, 1) {real, imag} */,
  {32'h3f885270, 32'hc22927f0} /* (13, 26, 0) {real, imag} */,
  {32'hc19e51e8, 32'h4129d61b} /* (13, 25, 31) {real, imag} */,
  {32'hc2a67b00, 32'hc1a10a10} /* (13, 25, 30) {real, imag} */,
  {32'hc1b219a9, 32'h40f8bb28} /* (13, 25, 29) {real, imag} */,
  {32'h413e8c6c, 32'hc1c64c8d} /* (13, 25, 28) {real, imag} */,
  {32'hc21b6246, 32'h40441a80} /* (13, 25, 27) {real, imag} */,
  {32'hc151e5f6, 32'h422f8f32} /* (13, 25, 26) {real, imag} */,
  {32'hc1d913db, 32'hc0da6c58} /* (13, 25, 25) {real, imag} */,
  {32'h403d913c, 32'h409951ca} /* (13, 25, 24) {real, imag} */,
  {32'h41503856, 32'h4130307a} /* (13, 25, 23) {real, imag} */,
  {32'h4186fa6e, 32'h40b73d2c} /* (13, 25, 22) {real, imag} */,
  {32'h4072c2c8, 32'hc1059e88} /* (13, 25, 21) {real, imag} */,
  {32'h4167ed78, 32'hc17d0a83} /* (13, 25, 20) {real, imag} */,
  {32'h40bf27a6, 32'h3ff10a58} /* (13, 25, 19) {real, imag} */,
  {32'hc06487c0, 32'hc0ebdae4} /* (13, 25, 18) {real, imag} */,
  {32'h4065ad90, 32'h3f0740c2} /* (13, 25, 17) {real, imag} */,
  {32'h405fa8c6, 32'hc05d4cbc} /* (13, 25, 16) {real, imag} */,
  {32'hc0ac83d4, 32'h3fbe512f} /* (13, 25, 15) {real, imag} */,
  {32'h40758eb0, 32'hc0148cf8} /* (13, 25, 14) {real, imag} */,
  {32'h40f0e5d4, 32'h4183688e} /* (13, 25, 13) {real, imag} */,
  {32'h4045ded8, 32'h415e1455} /* (13, 25, 12) {real, imag} */,
  {32'h4152ca82, 32'h41494436} /* (13, 25, 11) {real, imag} */,
  {32'h41fb719a, 32'h40bc6344} /* (13, 25, 10) {real, imag} */,
  {32'h3ee92300, 32'hc0642e6e} /* (13, 25, 9) {real, imag} */,
  {32'hc1ac6340, 32'hc1948720} /* (13, 25, 8) {real, imag} */,
  {32'h421b3110, 32'hc1d564f6} /* (13, 25, 7) {real, imag} */,
  {32'hc0a5cfe9, 32'hc1a3abab} /* (13, 25, 6) {real, imag} */,
  {32'hc1c2c6ba, 32'h425de9e8} /* (13, 25, 5) {real, imag} */,
  {32'hbfd326e0, 32'hc08c2a8c} /* (13, 25, 4) {real, imag} */,
  {32'hc0aa03e4, 32'hc26204cb} /* (13, 25, 3) {real, imag} */,
  {32'h4005a880, 32'h426301fc} /* (13, 25, 2) {real, imag} */,
  {32'hc1b7af84, 32'h412b557b} /* (13, 25, 1) {real, imag} */,
  {32'h4180cc83, 32'hc136bca5} /* (13, 25, 0) {real, imag} */,
  {32'hc12d7d9b, 32'h3f5beb40} /* (13, 24, 31) {real, imag} */,
  {32'hc203b23c, 32'hc1d73604} /* (13, 24, 30) {real, imag} */,
  {32'hc1a64ba6, 32'h40c366f7} /* (13, 24, 29) {real, imag} */,
  {32'hc086398c, 32'h41670990} /* (13, 24, 28) {real, imag} */,
  {32'hbf83fc98, 32'hc1d7abe6} /* (13, 24, 27) {real, imag} */,
  {32'hc194b5ac, 32'h41c7d2f9} /* (13, 24, 26) {real, imag} */,
  {32'h40296a88, 32'hc08a1e2c} /* (13, 24, 25) {real, imag} */,
  {32'h4238235e, 32'hc0900205} /* (13, 24, 24) {real, imag} */,
  {32'hc0e8f5c4, 32'hc0b8b4b4} /* (13, 24, 23) {real, imag} */,
  {32'h405255f2, 32'hc119a1cc} /* (13, 24, 22) {real, imag} */,
  {32'h41966c9a, 32'hc1680f85} /* (13, 24, 21) {real, imag} */,
  {32'hc10f8ab2, 32'hbf2c6838} /* (13, 24, 20) {real, imag} */,
  {32'hc0cb5119, 32'hc0e660a8} /* (13, 24, 19) {real, imag} */,
  {32'h3fe2e970, 32'h41542c46} /* (13, 24, 18) {real, imag} */,
  {32'hc122716a, 32'h3f416100} /* (13, 24, 17) {real, imag} */,
  {32'hbf0abff8, 32'h40725a22} /* (13, 24, 16) {real, imag} */,
  {32'h404f9692, 32'h407330b8} /* (13, 24, 15) {real, imag} */,
  {32'h3faebb80, 32'h40c712d4} /* (13, 24, 14) {real, imag} */,
  {32'h411c395c, 32'hc1b10ee4} /* (13, 24, 13) {real, imag} */,
  {32'hc08f4483, 32'h40f065c7} /* (13, 24, 12) {real, imag} */,
  {32'h402c7f88, 32'h40746874} /* (13, 24, 11) {real, imag} */,
  {32'hc10705a8, 32'h4089fe47} /* (13, 24, 10) {real, imag} */,
  {32'h4105d3de, 32'h40976630} /* (13, 24, 9) {real, imag} */,
  {32'h410fc706, 32'hc19acb85} /* (13, 24, 8) {real, imag} */,
  {32'hc12e6702, 32'hc1c5cb34} /* (13, 24, 7) {real, imag} */,
  {32'h40d75c98, 32'h41546172} /* (13, 24, 6) {real, imag} */,
  {32'hc15725bf, 32'h413cb3b4} /* (13, 24, 5) {real, imag} */,
  {32'h41f752e3, 32'h41fd0ef8} /* (13, 24, 4) {real, imag} */,
  {32'hc0816d28, 32'hc08ff155} /* (13, 24, 3) {real, imag} */,
  {32'h418831b0, 32'hc1b35838} /* (13, 24, 2) {real, imag} */,
  {32'hc0e7e31a, 32'hc2095833} /* (13, 24, 1) {real, imag} */,
  {32'h410942d4, 32'hc132ce08} /* (13, 24, 0) {real, imag} */,
  {32'hc1ef9e28, 32'h4229d11f} /* (13, 23, 31) {real, imag} */,
  {32'h40bd9524, 32'h41f4d942} /* (13, 23, 30) {real, imag} */,
  {32'h4187cdd3, 32'h401f8fbe} /* (13, 23, 29) {real, imag} */,
  {32'h40d7d2de, 32'hc133faba} /* (13, 23, 28) {real, imag} */,
  {32'hc1b1d137, 32'h3f7fc9e0} /* (13, 23, 27) {real, imag} */,
  {32'h40c732cc, 32'hc225db16} /* (13, 23, 26) {real, imag} */,
  {32'hc0e86f92, 32'hc1039d6a} /* (13, 23, 25) {real, imag} */,
  {32'h41218131, 32'hc219ad1d} /* (13, 23, 24) {real, imag} */,
  {32'hc094fe44, 32'h41a2cdc5} /* (13, 23, 23) {real, imag} */,
  {32'h3ecf7ae0, 32'h3f643420} /* (13, 23, 22) {real, imag} */,
  {32'h40b10b9a, 32'h4047f3d0} /* (13, 23, 21) {real, imag} */,
  {32'h3df5f4b8, 32'hc15ab8f4} /* (13, 23, 20) {real, imag} */,
  {32'h401c7568, 32'h3cc87780} /* (13, 23, 19) {real, imag} */,
  {32'h4096364a, 32'h40065ebc} /* (13, 23, 18) {real, imag} */,
  {32'hc0c0574c, 32'hbfc10b14} /* (13, 23, 17) {real, imag} */,
  {32'hc0a6bce0, 32'hc0b3473a} /* (13, 23, 16) {real, imag} */,
  {32'hc112de78, 32'hbfa3b92c} /* (13, 23, 15) {real, imag} */,
  {32'hc11df989, 32'h4181dcd4} /* (13, 23, 14) {real, imag} */,
  {32'h419662e1, 32'h40cbeebe} /* (13, 23, 13) {real, imag} */,
  {32'h3f6890c1, 32'hc048fd40} /* (13, 23, 12) {real, imag} */,
  {32'h4141b23d, 32'hc1b25bf5} /* (13, 23, 11) {real, imag} */,
  {32'hc06d8918, 32'hc16a4dde} /* (13, 23, 10) {real, imag} */,
  {32'hc1798ba0, 32'hc16f9882} /* (13, 23, 9) {real, imag} */,
  {32'hc012945c, 32'h41a11d9e} /* (13, 23, 8) {real, imag} */,
  {32'h40fe0732, 32'h4177aa06} /* (13, 23, 7) {real, imag} */,
  {32'hc1174f81, 32'hc22793ea} /* (13, 23, 6) {real, imag} */,
  {32'h41d1bad9, 32'h4167fcf0} /* (13, 23, 5) {real, imag} */,
  {32'h4008a14d, 32'h3ee0d890} /* (13, 23, 4) {real, imag} */,
  {32'hc03c7dea, 32'hc12f1272} /* (13, 23, 3) {real, imag} */,
  {32'h421ff4f4, 32'hc1ba4892} /* (13, 23, 2) {real, imag} */,
  {32'h41724138, 32'h4220bc8f} /* (13, 23, 1) {real, imag} */,
  {32'hc0ed1c54, 32'h41a16f7e} /* (13, 23, 0) {real, imag} */,
  {32'hc0fe1020, 32'h41e02036} /* (13, 22, 31) {real, imag} */,
  {32'hc13d43b2, 32'hc0d1feee} /* (13, 22, 30) {real, imag} */,
  {32'h41bcacce, 32'hc19ca188} /* (13, 22, 29) {real, imag} */,
  {32'h404e9450, 32'hc186ce0d} /* (13, 22, 28) {real, imag} */,
  {32'hc10bcc40, 32'h411c1f30} /* (13, 22, 27) {real, imag} */,
  {32'hc09c222c, 32'h41040946} /* (13, 22, 26) {real, imag} */,
  {32'hc15afe80, 32'hc0afaaae} /* (13, 22, 25) {real, imag} */,
  {32'h4192b98e, 32'hc074515c} /* (13, 22, 24) {real, imag} */,
  {32'h4070155b, 32'hc1aa69f2} /* (13, 22, 23) {real, imag} */,
  {32'hc1925cd3, 32'hc121a3db} /* (13, 22, 22) {real, imag} */,
  {32'hc1c03572, 32'h401158bb} /* (13, 22, 21) {real, imag} */,
  {32'h40098444, 32'h41519425} /* (13, 22, 20) {real, imag} */,
  {32'h40d0b8bf, 32'h40029782} /* (13, 22, 19) {real, imag} */,
  {32'h3f7eabd8, 32'h416b22c5} /* (13, 22, 18) {real, imag} */,
  {32'hc001e863, 32'h3e65eaf0} /* (13, 22, 17) {real, imag} */,
  {32'hc002d5b8, 32'h3cfd0e00} /* (13, 22, 16) {real, imag} */,
  {32'hc0efac7e, 32'hc03b0971} /* (13, 22, 15) {real, imag} */,
  {32'h4068b86a, 32'hc10e6339} /* (13, 22, 14) {real, imag} */,
  {32'hc0e2d437, 32'hbfb6f8b4} /* (13, 22, 13) {real, imag} */,
  {32'h40300dda, 32'h406a8b2c} /* (13, 22, 12) {real, imag} */,
  {32'hc12a6530, 32'h411f46f6} /* (13, 22, 11) {real, imag} */,
  {32'h410c5dba, 32'h3f9b87e8} /* (13, 22, 10) {real, imag} */,
  {32'h410df51a, 32'h3f6b7480} /* (13, 22, 9) {real, imag} */,
  {32'h4089f0e6, 32'h40454ea0} /* (13, 22, 8) {real, imag} */,
  {32'h40e2a103, 32'h41829a6a} /* (13, 22, 7) {real, imag} */,
  {32'hc1f18157, 32'h41b277ea} /* (13, 22, 6) {real, imag} */,
  {32'h41a79cfe, 32'h41adcb2c} /* (13, 22, 5) {real, imag} */,
  {32'h4166d43a, 32'hc1907283} /* (13, 22, 4) {real, imag} */,
  {32'h419471b0, 32'hbf4fb8f0} /* (13, 22, 3) {real, imag} */,
  {32'hc18f9a6b, 32'hbf28b630} /* (13, 22, 2) {real, imag} */,
  {32'hc1d04290, 32'hc1519d3d} /* (13, 22, 1) {real, imag} */,
  {32'h41bf4c73, 32'hc1cc3f1a} /* (13, 22, 0) {real, imag} */,
  {32'hbfa65a5a, 32'h41188f4c} /* (13, 21, 31) {real, imag} */,
  {32'hc120af1d, 32'h421fe89b} /* (13, 21, 30) {real, imag} */,
  {32'h42216c5a, 32'h42214c5a} /* (13, 21, 29) {real, imag} */,
  {32'h40867204, 32'hbe7e8b40} /* (13, 21, 28) {real, imag} */,
  {32'hc08a81ab, 32'hc1c7007e} /* (13, 21, 27) {real, imag} */,
  {32'hc1909627, 32'h40c24a14} /* (13, 21, 26) {real, imag} */,
  {32'h41c539ae, 32'h3f3ee764} /* (13, 21, 25) {real, imag} */,
  {32'hc0cf6c55, 32'h41526128} /* (13, 21, 24) {real, imag} */,
  {32'hbf304de0, 32'hbf1aff28} /* (13, 21, 23) {real, imag} */,
  {32'hc00e8d72, 32'hbfec0bd8} /* (13, 21, 22) {real, imag} */,
  {32'h41580d64, 32'hc0b0520c} /* (13, 21, 21) {real, imag} */,
  {32'h3f6462f0, 32'hc0ee046a} /* (13, 21, 20) {real, imag} */,
  {32'hc0f13644, 32'h3ff13048} /* (13, 21, 19) {real, imag} */,
  {32'h3fc2a688, 32'h40574c30} /* (13, 21, 18) {real, imag} */,
  {32'h3e6111a0, 32'hbf92638e} /* (13, 21, 17) {real, imag} */,
  {32'hbf7e7ed0, 32'h403e1204} /* (13, 21, 16) {real, imag} */,
  {32'hc09a3e3f, 32'hc0b15b2e} /* (13, 21, 15) {real, imag} */,
  {32'hbf4ad5f0, 32'hc052e208} /* (13, 21, 14) {real, imag} */,
  {32'h413534e0, 32'h3fc4acd8} /* (13, 21, 13) {real, imag} */,
  {32'h40d6cf44, 32'h4011c6d3} /* (13, 21, 12) {real, imag} */,
  {32'h401fac0a, 32'h41708564} /* (13, 21, 11) {real, imag} */,
  {32'hc0519572, 32'h409afa06} /* (13, 21, 10) {real, imag} */,
  {32'h4102064c, 32'hc141bf68} /* (13, 21, 9) {real, imag} */,
  {32'h4166db6a, 32'hc125b160} /* (13, 21, 8) {real, imag} */,
  {32'hc1a6f7ae, 32'h3f4b1fec} /* (13, 21, 7) {real, imag} */,
  {32'h410cf8d2, 32'hc231f584} /* (13, 21, 6) {real, imag} */,
  {32'hc0c7d4cd, 32'h4115e6bd} /* (13, 21, 5) {real, imag} */,
  {32'h3ebfc180, 32'h414ef28b} /* (13, 21, 4) {real, imag} */,
  {32'h412a9569, 32'h3f445ae0} /* (13, 21, 3) {real, imag} */,
  {32'h419d6848, 32'hc01ee290} /* (13, 21, 2) {real, imag} */,
  {32'h3f2d49a7, 32'hc0ac8fe1} /* (13, 21, 1) {real, imag} */,
  {32'hc04dded4, 32'hbfc69a60} /* (13, 21, 0) {real, imag} */,
  {32'hc1295c3e, 32'hc04e27f4} /* (13, 20, 31) {real, imag} */,
  {32'hc162523a, 32'hc0829f28} /* (13, 20, 30) {real, imag} */,
  {32'h418ccb86, 32'h40e79158} /* (13, 20, 29) {real, imag} */,
  {32'hc17f237a, 32'hbf9d7604} /* (13, 20, 28) {real, imag} */,
  {32'h411382d1, 32'hbfd59aec} /* (13, 20, 27) {real, imag} */,
  {32'hc11b11ba, 32'h3e535ed0} /* (13, 20, 26) {real, imag} */,
  {32'h410a3b2b, 32'hc1d3bf42} /* (13, 20, 25) {real, imag} */,
  {32'hc0a91dde, 32'h4073cf5b} /* (13, 20, 24) {real, imag} */,
  {32'h40eac590, 32'h40a0f92f} /* (13, 20, 23) {real, imag} */,
  {32'h413ec38a, 32'hc0acbb67} /* (13, 20, 22) {real, imag} */,
  {32'hc04361a4, 32'h40be89b2} /* (13, 20, 21) {real, imag} */,
  {32'hbfd407e6, 32'hbf596cb2} /* (13, 20, 20) {real, imag} */,
  {32'h401d76e8, 32'hc06c78b6} /* (13, 20, 19) {real, imag} */,
  {32'hbed2d128, 32'h40ab452d} /* (13, 20, 18) {real, imag} */,
  {32'h3f9799cf, 32'hc03a2dc0} /* (13, 20, 17) {real, imag} */,
  {32'h4002f44f, 32'hbfd0f660} /* (13, 20, 16) {real, imag} */,
  {32'h40836802, 32'hc03da1f8} /* (13, 20, 15) {real, imag} */,
  {32'h4035be61, 32'hbfb413f4} /* (13, 20, 14) {real, imag} */,
  {32'h3f066580, 32'h401ebf46} /* (13, 20, 13) {real, imag} */,
  {32'h40aa235c, 32'h3f3b3442} /* (13, 20, 12) {real, imag} */,
  {32'hc0aac336, 32'h41372391} /* (13, 20, 11) {real, imag} */,
  {32'hc0d4c7f5, 32'h40a0a159} /* (13, 20, 10) {real, imag} */,
  {32'hc01c0221, 32'hc0d28ad9} /* (13, 20, 9) {real, imag} */,
  {32'h41124bd7, 32'hc0cf18ea} /* (13, 20, 8) {real, imag} */,
  {32'hbfb78606, 32'h40d47560} /* (13, 20, 7) {real, imag} */,
  {32'h41cd5185, 32'h404d01e3} /* (13, 20, 6) {real, imag} */,
  {32'hc19e96f6, 32'hc1177db2} /* (13, 20, 5) {real, imag} */,
  {32'hc08f0954, 32'h40f7d29b} /* (13, 20, 4) {real, imag} */,
  {32'h41c51b12, 32'hbf78e550} /* (13, 20, 3) {real, imag} */,
  {32'hc0fe7b64, 32'h41891c46} /* (13, 20, 2) {real, imag} */,
  {32'hc1088ada, 32'hc11893a9} /* (13, 20, 1) {real, imag} */,
  {32'hc0cca9f0, 32'h412e28d0} /* (13, 20, 0) {real, imag} */,
  {32'hbf8cc994, 32'hc1401885} /* (13, 19, 31) {real, imag} */,
  {32'hbfc29b88, 32'hc021d7da} /* (13, 19, 30) {real, imag} */,
  {32'h405f6c10, 32'h40a3fe24} /* (13, 19, 29) {real, imag} */,
  {32'h40c8a516, 32'hc0654c37} /* (13, 19, 28) {real, imag} */,
  {32'hc1925f72, 32'hc1134244} /* (13, 19, 27) {real, imag} */,
  {32'h411faae0, 32'h40c93c5f} /* (13, 19, 26) {real, imag} */,
  {32'hc1730c2e, 32'hc0ea58ef} /* (13, 19, 25) {real, imag} */,
  {32'h406318b5, 32'hc09332fc} /* (13, 19, 24) {real, imag} */,
  {32'h3fefd0c2, 32'h40e8e283} /* (13, 19, 23) {real, imag} */,
  {32'hc029fcd0, 32'h4004999a} /* (13, 19, 22) {real, imag} */,
  {32'hc0d81709, 32'h3ea32930} /* (13, 19, 21) {real, imag} */,
  {32'hbf5b461e, 32'h3d42d600} /* (13, 19, 20) {real, imag} */,
  {32'h3fc72b8c, 32'hbd12d600} /* (13, 19, 19) {real, imag} */,
  {32'hc04e2214, 32'hc099c319} /* (13, 19, 18) {real, imag} */,
  {32'h40d4cdb2, 32'hbfd634aa} /* (13, 19, 17) {real, imag} */,
  {32'hbfe72e20, 32'h4011dac6} /* (13, 19, 16) {real, imag} */,
  {32'hbf5a9330, 32'hbf182ddc} /* (13, 19, 15) {real, imag} */,
  {32'hc09a9da8, 32'h3f694c76} /* (13, 19, 14) {real, imag} */,
  {32'hbe8245b0, 32'hc0852f0c} /* (13, 19, 13) {real, imag} */,
  {32'hc0246608, 32'h404ef71a} /* (13, 19, 12) {real, imag} */,
  {32'h409932cd, 32'h4117bdc2} /* (13, 19, 11) {real, imag} */,
  {32'hbebcb63c, 32'hc104fc6e} /* (13, 19, 10) {real, imag} */,
  {32'h40b57194, 32'hc0ba7b45} /* (13, 19, 9) {real, imag} */,
  {32'hbff5973e, 32'hc140a702} /* (13, 19, 8) {real, imag} */,
  {32'h3fd9c450, 32'h416d0c2c} /* (13, 19, 7) {real, imag} */,
  {32'h40106216, 32'hbf268318} /* (13, 19, 6) {real, imag} */,
  {32'hc07529ea, 32'hc0061d12} /* (13, 19, 5) {real, imag} */,
  {32'hc189d566, 32'hc0c584b0} /* (13, 19, 4) {real, imag} */,
  {32'hc1c775e6, 32'hc1068c06} /* (13, 19, 3) {real, imag} */,
  {32'h40ccdcc2, 32'h40b2dd63} /* (13, 19, 2) {real, imag} */,
  {32'h40dbeb07, 32'hc187a0c7} /* (13, 19, 1) {real, imag} */,
  {32'hc1255440, 32'hc144002e} /* (13, 19, 0) {real, imag} */,
  {32'hbffd83d0, 32'hc13a0548} /* (13, 18, 31) {real, imag} */,
  {32'h406c1400, 32'hc12a2e44} /* (13, 18, 30) {real, imag} */,
  {32'hc15ac989, 32'hc07b5c40} /* (13, 18, 29) {real, imag} */,
  {32'h40138330, 32'h40b0637a} /* (13, 18, 28) {real, imag} */,
  {32'hc0c0b928, 32'hc17a872c} /* (13, 18, 27) {real, imag} */,
  {32'h413b2851, 32'hc01565a0} /* (13, 18, 26) {real, imag} */,
  {32'h414f3d98, 32'hc1636891} /* (13, 18, 25) {real, imag} */,
  {32'h412fd6da, 32'hc12afc24} /* (13, 18, 24) {real, imag} */,
  {32'h4087d78c, 32'h4118d965} /* (13, 18, 23) {real, imag} */,
  {32'hc19cdcdc, 32'h4003850d} /* (13, 18, 22) {real, imag} */,
  {32'h3ef021c0, 32'hbf996474} /* (13, 18, 21) {real, imag} */,
  {32'hc0775afc, 32'hbfebebec} /* (13, 18, 20) {real, imag} */,
  {32'hc02eb493, 32'h402bb7c6} /* (13, 18, 19) {real, imag} */,
  {32'hbec78e88, 32'hc0206606} /* (13, 18, 18) {real, imag} */,
  {32'h3f79a74c, 32'h3e31de70} /* (13, 18, 17) {real, imag} */,
  {32'h4051d35a, 32'h4084dfe5} /* (13, 18, 16) {real, imag} */,
  {32'h3fb722b2, 32'h401d8d03} /* (13, 18, 15) {real, imag} */,
  {32'hc08d1994, 32'hc0620606} /* (13, 18, 14) {real, imag} */,
  {32'h3fac20fe, 32'hc03631e0} /* (13, 18, 13) {real, imag} */,
  {32'hc06c08e8, 32'hc04e7440} /* (13, 18, 12) {real, imag} */,
  {32'hc11cf14c, 32'h40d65785} /* (13, 18, 11) {real, imag} */,
  {32'h4020feec, 32'h41048eaf} /* (13, 18, 10) {real, imag} */,
  {32'hc0c899e2, 32'hc0921df2} /* (13, 18, 9) {real, imag} */,
  {32'hc0499692, 32'hc11c92c0} /* (13, 18, 8) {real, imag} */,
  {32'hbf8189cc, 32'h414e3dc9} /* (13, 18, 7) {real, imag} */,
  {32'h3ff20de8, 32'h4145775c} /* (13, 18, 6) {real, imag} */,
  {32'h40d992d4, 32'hc0ee6555} /* (13, 18, 5) {real, imag} */,
  {32'h413676cd, 32'h3f142164} /* (13, 18, 4) {real, imag} */,
  {32'hc18e2802, 32'h417cb2a4} /* (13, 18, 3) {real, imag} */,
  {32'hc1ad5aef, 32'h409513a9} /* (13, 18, 2) {real, imag} */,
  {32'h3eb43400, 32'hc08505e3} /* (13, 18, 1) {real, imag} */,
  {32'hc036fb32, 32'hc11be248} /* (13, 18, 0) {real, imag} */,
  {32'hc0a7f25a, 32'h3fdafa50} /* (13, 17, 31) {real, imag} */,
  {32'h40d6ecf6, 32'hc15fe71a} /* (13, 17, 30) {real, imag} */,
  {32'h40720040, 32'h41d79666} /* (13, 17, 29) {real, imag} */,
  {32'h40fde070, 32'h4055c7de} /* (13, 17, 28) {real, imag} */,
  {32'hbfa08068, 32'h412135c4} /* (13, 17, 27) {real, imag} */,
  {32'hc08cded5, 32'hc0632305} /* (13, 17, 26) {real, imag} */,
  {32'hc0796500, 32'h407ffe7e} /* (13, 17, 25) {real, imag} */,
  {32'h3f9908dc, 32'hc0bb327c} /* (13, 17, 24) {real, imag} */,
  {32'hc02348e0, 32'h40479b4f} /* (13, 17, 23) {real, imag} */,
  {32'h40572091, 32'hbe9fc2c0} /* (13, 17, 22) {real, imag} */,
  {32'h3fbdc914, 32'hbe57f040} /* (13, 17, 21) {real, imag} */,
  {32'hc009595a, 32'hbf4908b6} /* (13, 17, 20) {real, imag} */,
  {32'h40424c3e, 32'hc054fd74} /* (13, 17, 19) {real, imag} */,
  {32'h4087b6a9, 32'h3e822828} /* (13, 17, 18) {real, imag} */,
  {32'h3f2e7d44, 32'h3ed8d428} /* (13, 17, 17) {real, imag} */,
  {32'hbff44410, 32'h40085937} /* (13, 17, 16) {real, imag} */,
  {32'hc0a1e142, 32'hbd8c7620} /* (13, 17, 15) {real, imag} */,
  {32'hbfecfd51, 32'hbcddbb80} /* (13, 17, 14) {real, imag} */,
  {32'hbf47bef8, 32'hbd9e2b80} /* (13, 17, 13) {real, imag} */,
  {32'h3f0a55a0, 32'hc0326d9a} /* (13, 17, 12) {real, imag} */,
  {32'h4095c9e5, 32'hbe616180} /* (13, 17, 11) {real, imag} */,
  {32'h408f1dcc, 32'hbe4a29a0} /* (13, 17, 10) {real, imag} */,
  {32'h401da048, 32'hc03fab71} /* (13, 17, 9) {real, imag} */,
  {32'h40295959, 32'h40b8bab0} /* (13, 17, 8) {real, imag} */,
  {32'h410efca0, 32'h402cae40} /* (13, 17, 7) {real, imag} */,
  {32'hc0c0fa23, 32'hbfa31c72} /* (13, 17, 6) {real, imag} */,
  {32'hc05d67dc, 32'h3fff069c} /* (13, 17, 5) {real, imag} */,
  {32'hc0deaea0, 32'hc105827a} /* (13, 17, 4) {real, imag} */,
  {32'hc19e6e1e, 32'h4090fe22} /* (13, 17, 3) {real, imag} */,
  {32'hbe8bc628, 32'h4047e738} /* (13, 17, 2) {real, imag} */,
  {32'hbfc30062, 32'h41343a96} /* (13, 17, 1) {real, imag} */,
  {32'h40ce3858, 32'hbfc8ec94} /* (13, 17, 0) {real, imag} */,
  {32'h409d066c, 32'h3ea67bdc} /* (13, 16, 31) {real, imag} */,
  {32'h4156a9e0, 32'h4174f1bd} /* (13, 16, 30) {real, imag} */,
  {32'hc117cb07, 32'h408841b6} /* (13, 16, 29) {real, imag} */,
  {32'h3e64cc2c, 32'h41138462} /* (13, 16, 28) {real, imag} */,
  {32'h412d7dbc, 32'h41715b7a} /* (13, 16, 27) {real, imag} */,
  {32'h40d0beb1, 32'h3f9d15f4} /* (13, 16, 26) {real, imag} */,
  {32'hc015e63d, 32'h417183da} /* (13, 16, 25) {real, imag} */,
  {32'hc04f06f4, 32'hc081f48e} /* (13, 16, 24) {real, imag} */,
  {32'hc075d805, 32'h413293c0} /* (13, 16, 23) {real, imag} */,
  {32'hc0a606aa, 32'hc0f3c604} /* (13, 16, 22) {real, imag} */,
  {32'h40c32dc7, 32'hbffe8d12} /* (13, 16, 21) {real, imag} */,
  {32'h3f8a99fe, 32'h3f051b80} /* (13, 16, 20) {real, imag} */,
  {32'h408fecba, 32'h4003a035} /* (13, 16, 19) {real, imag} */,
  {32'hbc9db040, 32'h40cdab9e} /* (13, 16, 18) {real, imag} */,
  {32'hbe782aa4, 32'hbf8e5dee} /* (13, 16, 17) {real, imag} */,
  {32'hbf97bc84, 32'hc011f05d} /* (13, 16, 16) {real, imag} */,
  {32'h3f8e36b4, 32'hbf89a508} /* (13, 16, 15) {real, imag} */,
  {32'hc0070190, 32'h3f7279ac} /* (13, 16, 14) {real, imag} */,
  {32'hc059b4bd, 32'h3dc99020} /* (13, 16, 13) {real, imag} */,
  {32'hc0b02c26, 32'h3e8275bf} /* (13, 16, 12) {real, imag} */,
  {32'hbfa0858c, 32'hc0bb141e} /* (13, 16, 11) {real, imag} */,
  {32'hbff05c12, 32'hc0518cab} /* (13, 16, 10) {real, imag} */,
  {32'h412128e4, 32'h40923b5e} /* (13, 16, 9) {real, imag} */,
  {32'hbf9c1604, 32'h3fe2feac} /* (13, 16, 8) {real, imag} */,
  {32'hc05560d9, 32'h4128ee92} /* (13, 16, 7) {real, imag} */,
  {32'h4074337e, 32'hc10df8c8} /* (13, 16, 6) {real, imag} */,
  {32'h3f099858, 32'hc1371fee} /* (13, 16, 5) {real, imag} */,
  {32'hbfb2c3ca, 32'hc103745c} /* (13, 16, 4) {real, imag} */,
  {32'h3fd723b8, 32'hc0c4aa54} /* (13, 16, 3) {real, imag} */,
  {32'h418bac76, 32'hc14e8087} /* (13, 16, 2) {real, imag} */,
  {32'hc102e189, 32'h40812f98} /* (13, 16, 1) {real, imag} */,
  {32'h40cb4200, 32'hc1089d9b} /* (13, 16, 0) {real, imag} */,
  {32'hc11c8087, 32'hc0c90277} /* (13, 15, 31) {real, imag} */,
  {32'h3f2858da, 32'hbf76c8b0} /* (13, 15, 30) {real, imag} */,
  {32'h40ce5c5b, 32'h406ea5bc} /* (13, 15, 29) {real, imag} */,
  {32'h417657a2, 32'hbf668aa4} /* (13, 15, 28) {real, imag} */,
  {32'h40cf9f04, 32'h403c235a} /* (13, 15, 27) {real, imag} */,
  {32'hc05fbd9f, 32'hc08b1ea9} /* (13, 15, 26) {real, imag} */,
  {32'hc01bb04e, 32'h40aed174} /* (13, 15, 25) {real, imag} */,
  {32'h406e6f30, 32'h40371244} /* (13, 15, 24) {real, imag} */,
  {32'hbda01b40, 32'h3ebfcf70} /* (13, 15, 23) {real, imag} */,
  {32'hc09483d8, 32'h3f4c3bba} /* (13, 15, 22) {real, imag} */,
  {32'h4021fd26, 32'h40431ef8} /* (13, 15, 21) {real, imag} */,
  {32'hc09fd7be, 32'h4058d5b1} /* (13, 15, 20) {real, imag} */,
  {32'h3f6aaf7a, 32'h4033e07e} /* (13, 15, 19) {real, imag} */,
  {32'hbfcac988, 32'h3ed295d8} /* (13, 15, 18) {real, imag} */,
  {32'h3f6720ec, 32'h401d77b6} /* (13, 15, 17) {real, imag} */,
  {32'h402d2668, 32'hbfbdcaee} /* (13, 15, 16) {real, imag} */,
  {32'hc00346e7, 32'hc093249f} /* (13, 15, 15) {real, imag} */,
  {32'h401ec2bc, 32'hbfa0cb0a} /* (13, 15, 14) {real, imag} */,
  {32'hbf630566, 32'h403d7e80} /* (13, 15, 13) {real, imag} */,
  {32'h401df50c, 32'h401f3c67} /* (13, 15, 12) {real, imag} */,
  {32'h405ce304, 32'h40f1ff0e} /* (13, 15, 11) {real, imag} */,
  {32'h40c3d2ac, 32'h400013a6} /* (13, 15, 10) {real, imag} */,
  {32'hc1307f40, 32'hc04e2e42} /* (13, 15, 9) {real, imag} */,
  {32'h3f9ab80c, 32'h3eb4900c} /* (13, 15, 8) {real, imag} */,
  {32'hc1032b64, 32'hc0faa994} /* (13, 15, 7) {real, imag} */,
  {32'hc0f49748, 32'h40c7681f} /* (13, 15, 6) {real, imag} */,
  {32'h411ec0c6, 32'hc0fff61d} /* (13, 15, 5) {real, imag} */,
  {32'h413910da, 32'h40a54a84} /* (13, 15, 4) {real, imag} */,
  {32'hc1483a60, 32'h415abdb5} /* (13, 15, 3) {real, imag} */,
  {32'hbf3e729a, 32'hc140ab01} /* (13, 15, 2) {real, imag} */,
  {32'hc10462c1, 32'hc0ccba71} /* (13, 15, 1) {real, imag} */,
  {32'h4182e734, 32'hc041e529} /* (13, 15, 0) {real, imag} */,
  {32'hc17d7328, 32'h401a4e42} /* (13, 14, 31) {real, imag} */,
  {32'h40e5aa01, 32'hc198cebd} /* (13, 14, 30) {real, imag} */,
  {32'h41760910, 32'h412da377} /* (13, 14, 29) {real, imag} */,
  {32'hc1077aa8, 32'hbec00c30} /* (13, 14, 28) {real, imag} */,
  {32'hc1045dbe, 32'hbeb04204} /* (13, 14, 27) {real, imag} */,
  {32'hbf4dd812, 32'h41338d5a} /* (13, 14, 26) {real, imag} */,
  {32'hbe912c98, 32'hc106bcdd} /* (13, 14, 25) {real, imag} */,
  {32'hbf508640, 32'h3fc9b544} /* (13, 14, 24) {real, imag} */,
  {32'h4106cde4, 32'h40bd5322} /* (13, 14, 23) {real, imag} */,
  {32'h409de2d2, 32'hbfc50e48} /* (13, 14, 22) {real, imag} */,
  {32'h4073e389, 32'hc0d67915} /* (13, 14, 21) {real, imag} */,
  {32'h403a5d40, 32'hc06e8529} /* (13, 14, 20) {real, imag} */,
  {32'hc0af33a1, 32'hbfba75c6} /* (13, 14, 19) {real, imag} */,
  {32'hbe005720, 32'h3de80800} /* (13, 14, 18) {real, imag} */,
  {32'h3f1ba428, 32'hbfcae7cc} /* (13, 14, 17) {real, imag} */,
  {32'h3fcd232c, 32'h40684b7c} /* (13, 14, 16) {real, imag} */,
  {32'hbe626b20, 32'hbfb9c0cc} /* (13, 14, 15) {real, imag} */,
  {32'h3f97ae24, 32'h404b6db0} /* (13, 14, 14) {real, imag} */,
  {32'hbec75210, 32'hc09b70fa} /* (13, 14, 13) {real, imag} */,
  {32'h3f795d42, 32'hc0447da3} /* (13, 14, 12) {real, imag} */,
  {32'h40a665fc, 32'h40788c22} /* (13, 14, 11) {real, imag} */,
  {32'hc0c02ef2, 32'hc023a434} /* (13, 14, 10) {real, imag} */,
  {32'hc055b93e, 32'h40333908} /* (13, 14, 9) {real, imag} */,
  {32'h410e9e99, 32'hc10597c6} /* (13, 14, 8) {real, imag} */,
  {32'h4062985b, 32'hc0aa8c34} /* (13, 14, 7) {real, imag} */,
  {32'h403c23e4, 32'hc0729ce8} /* (13, 14, 6) {real, imag} */,
  {32'h40e1a588, 32'hc00fdeb4} /* (13, 14, 5) {real, imag} */,
  {32'hc0f593bb, 32'hc0b159e3} /* (13, 14, 4) {real, imag} */,
  {32'h40b819af, 32'hc0c23b7e} /* (13, 14, 3) {real, imag} */,
  {32'hc0fdaf45, 32'h400a07e8} /* (13, 14, 2) {real, imag} */,
  {32'hbf1d6fe8, 32'h41418462} /* (13, 14, 1) {real, imag} */,
  {32'h416df062, 32'hc1628ac1} /* (13, 14, 0) {real, imag} */,
  {32'hc17b4330, 32'h4154eb75} /* (13, 13, 31) {real, imag} */,
  {32'h41ac6668, 32'h4011462a} /* (13, 13, 30) {real, imag} */,
  {32'hc1b92535, 32'hc1b0d56e} /* (13, 13, 29) {real, imag} */,
  {32'hc1533598, 32'hc1199086} /* (13, 13, 28) {real, imag} */,
  {32'h3f463d50, 32'hc1b4c5c5} /* (13, 13, 27) {real, imag} */,
  {32'h40a3032c, 32'h418eb3c7} /* (13, 13, 26) {real, imag} */,
  {32'hc0981b9b, 32'hc1059745} /* (13, 13, 25) {real, imag} */,
  {32'h414d2af6, 32'h410c9770} /* (13, 13, 24) {real, imag} */,
  {32'hc1541fe1, 32'hc0d5eddb} /* (13, 13, 23) {real, imag} */,
  {32'hc094578e, 32'h4101aa38} /* (13, 13, 22) {real, imag} */,
  {32'hc07bc3b3, 32'h40d4643d} /* (13, 13, 21) {real, imag} */,
  {32'h4009b01a, 32'hc0ab493b} /* (13, 13, 20) {real, imag} */,
  {32'hc08081f0, 32'hc02738f4} /* (13, 13, 19) {real, imag} */,
  {32'hbfb63f90, 32'hbfebe034} /* (13, 13, 18) {real, imag} */,
  {32'hbf5bb068, 32'hbef8a198} /* (13, 13, 17) {real, imag} */,
  {32'h402a059c, 32'hc07b15e4} /* (13, 13, 16) {real, imag} */,
  {32'hc03cb85a, 32'h408edfca} /* (13, 13, 15) {real, imag} */,
  {32'hc0397408, 32'hc085bd29} /* (13, 13, 14) {real, imag} */,
  {32'h4104abe8, 32'hbe622140} /* (13, 13, 13) {real, imag} */,
  {32'hbf59c450, 32'h4046247a} /* (13, 13, 12) {real, imag} */,
  {32'hc0e80742, 32'hbf470d38} /* (13, 13, 11) {real, imag} */,
  {32'h4086177e, 32'hbff11634} /* (13, 13, 10) {real, imag} */,
  {32'hc0f9004e, 32'hbeee5a30} /* (13, 13, 9) {real, imag} */,
  {32'hc16c4838, 32'hc0d89a65} /* (13, 13, 8) {real, imag} */,
  {32'h409fe9e5, 32'h413c4f2f} /* (13, 13, 7) {real, imag} */,
  {32'h41c4ef91, 32'hc163afba} /* (13, 13, 6) {real, imag} */,
  {32'h41210367, 32'h412ee57e} /* (13, 13, 5) {real, imag} */,
  {32'h40196aa0, 32'hc1329b4a} /* (13, 13, 4) {real, imag} */,
  {32'h41055026, 32'h40929ad6} /* (13, 13, 3) {real, imag} */,
  {32'h413c2710, 32'hc1583910} /* (13, 13, 2) {real, imag} */,
  {32'h41721160, 32'h3f97ee98} /* (13, 13, 1) {real, imag} */,
  {32'hc197f6b6, 32'hc1419067} /* (13, 13, 0) {real, imag} */,
  {32'h3f9ace30, 32'hc08040a8} /* (13, 12, 31) {real, imag} */,
  {32'hc18c66e7, 32'h4112db28} /* (13, 12, 30) {real, imag} */,
  {32'h3fd71368, 32'hc0acca00} /* (13, 12, 29) {real, imag} */,
  {32'h4102b212, 32'hc0a73bb0} /* (13, 12, 28) {real, imag} */,
  {32'h40f4923f, 32'h4179780b} /* (13, 12, 27) {real, imag} */,
  {32'hc1b61c25, 32'h3fefc48c} /* (13, 12, 26) {real, imag} */,
  {32'h41e04284, 32'hbfbf22da} /* (13, 12, 25) {real, imag} */,
  {32'hc120ba73, 32'hbf20d3d0} /* (13, 12, 24) {real, imag} */,
  {32'h4110972d, 32'h3d247040} /* (13, 12, 23) {real, imag} */,
  {32'h41014fa8, 32'h3f60871d} /* (13, 12, 22) {real, imag} */,
  {32'h41177a23, 32'hc0ff1e82} /* (13, 12, 21) {real, imag} */,
  {32'h40850080, 32'h4015d1cf} /* (13, 12, 20) {real, imag} */,
  {32'hbf600530, 32'hc093329b} /* (13, 12, 19) {real, imag} */,
  {32'hc0841f04, 32'h4044f69f} /* (13, 12, 18) {real, imag} */,
  {32'h4012c45c, 32'h408c3272} /* (13, 12, 17) {real, imag} */,
  {32'hbf9c68d8, 32'h4015aaac} /* (13, 12, 16) {real, imag} */,
  {32'h40236c94, 32'hc10b8017} /* (13, 12, 15) {real, imag} */,
  {32'h402a6298, 32'h3ea5c928} /* (13, 12, 14) {real, imag} */,
  {32'hc05d1c8e, 32'hc0083e52} /* (13, 12, 13) {real, imag} */,
  {32'h4120764c, 32'h4016e693} /* (13, 12, 12) {real, imag} */,
  {32'h4133708d, 32'hc0018e5d} /* (13, 12, 11) {real, imag} */,
  {32'hbfe17484, 32'h3fa88d90} /* (13, 12, 10) {real, imag} */,
  {32'hbf82a688, 32'h3f743f14} /* (13, 12, 9) {real, imag} */,
  {32'hc01ee683, 32'hc132cf27} /* (13, 12, 8) {real, imag} */,
  {32'h410ba8e3, 32'h3fe3ff7e} /* (13, 12, 7) {real, imag} */,
  {32'hc01fc4d8, 32'h4014201a} /* (13, 12, 6) {real, imag} */,
  {32'hc10494e2, 32'h3fa24008} /* (13, 12, 5) {real, imag} */,
  {32'hc1f4f345, 32'h40e8d0ea} /* (13, 12, 4) {real, imag} */,
  {32'h40363556, 32'hc20de662} /* (13, 12, 3) {real, imag} */,
  {32'h4172b416, 32'hc0d43b08} /* (13, 12, 2) {real, imag} */,
  {32'h41c0b7b4, 32'h4157460a} /* (13, 12, 1) {real, imag} */,
  {32'hc16ff401, 32'h413c5549} /* (13, 12, 0) {real, imag} */,
  {32'h409f0fd5, 32'h408bfdb4} /* (13, 11, 31) {real, imag} */,
  {32'h40ee9fd4, 32'hc11d29f0} /* (13, 11, 30) {real, imag} */,
  {32'hc103e2ba, 32'h40d6ad1c} /* (13, 11, 29) {real, imag} */,
  {32'h40cfd567, 32'hc0a79e5e} /* (13, 11, 28) {real, imag} */,
  {32'h4109224a, 32'h3e3301a0} /* (13, 11, 27) {real, imag} */,
  {32'h40b60d80, 32'h40f03ef9} /* (13, 11, 26) {real, imag} */,
  {32'hc1700e97, 32'hc1738ff2} /* (13, 11, 25) {real, imag} */,
  {32'hc0cbd748, 32'h3fdacfb0} /* (13, 11, 24) {real, imag} */,
  {32'hc202f5f8, 32'h40058dd4} /* (13, 11, 23) {real, imag} */,
  {32'hc1395956, 32'hc0f4f024} /* (13, 11, 22) {real, imag} */,
  {32'hc128ed18, 32'hbf909514} /* (13, 11, 21) {real, imag} */,
  {32'h412dfa5e, 32'h3eb61340} /* (13, 11, 20) {real, imag} */,
  {32'h3eb10920, 32'h4088e4fe} /* (13, 11, 19) {real, imag} */,
  {32'h40f0a58c, 32'h403e44d2} /* (13, 11, 18) {real, imag} */,
  {32'h409e5417, 32'hc08e6668} /* (13, 11, 17) {real, imag} */,
  {32'hc03e89a2, 32'h3fec8550} /* (13, 11, 16) {real, imag} */,
  {32'hc0270716, 32'hc0318e90} /* (13, 11, 15) {real, imag} */,
  {32'h3fc80fae, 32'h3fc4b354} /* (13, 11, 14) {real, imag} */,
  {32'h40a47574, 32'h3f913852} /* (13, 11, 13) {real, imag} */,
  {32'h4093422b, 32'h41128cca} /* (13, 11, 12) {real, imag} */,
  {32'h4126a134, 32'hc175b186} /* (13, 11, 11) {real, imag} */,
  {32'hbf8a263c, 32'h40e5d056} /* (13, 11, 10) {real, imag} */,
  {32'hc0de25ec, 32'h416aca51} /* (13, 11, 9) {real, imag} */,
  {32'hc1253a74, 32'hc19802e7} /* (13, 11, 8) {real, imag} */,
  {32'h3ebdb1a0, 32'h40ba5764} /* (13, 11, 7) {real, imag} */,
  {32'hc219a564, 32'h4061160e} /* (13, 11, 6) {real, imag} */,
  {32'hc222bad6, 32'h4104e3de} /* (13, 11, 5) {real, imag} */,
  {32'hc0a37a5d, 32'h400cf604} /* (13, 11, 4) {real, imag} */,
  {32'h41dd4e01, 32'hc1c4bc11} /* (13, 11, 3) {real, imag} */,
  {32'h411b1c5e, 32'h41382028} /* (13, 11, 2) {real, imag} */,
  {32'hc032729a, 32'hc1f96659} /* (13, 11, 1) {real, imag} */,
  {32'hc0f3fbcf, 32'h416363f6} /* (13, 11, 0) {real, imag} */,
  {32'h41acbfe4, 32'h41ae0a01} /* (13, 10, 31) {real, imag} */,
  {32'hc1e1bffa, 32'h3fef67d8} /* (13, 10, 30) {real, imag} */,
  {32'hc1c39a52, 32'hc0924f47} /* (13, 10, 29) {real, imag} */,
  {32'hc25a3a1e, 32'hc1a6eab5} /* (13, 10, 28) {real, imag} */,
  {32'h423a0954, 32'hc0daafb6} /* (13, 10, 27) {real, imag} */,
  {32'h3fdd6a80, 32'h41310b16} /* (13, 10, 26) {real, imag} */,
  {32'h418834f8, 32'h40dc0833} /* (13, 10, 25) {real, imag} */,
  {32'h4093eee6, 32'hc1aa303a} /* (13, 10, 24) {real, imag} */,
  {32'h40ac04eb, 32'hc164dda0} /* (13, 10, 23) {real, imag} */,
  {32'hc093f0b2, 32'hc16e126c} /* (13, 10, 22) {real, imag} */,
  {32'h40ef7da8, 32'h41b1da0c} /* (13, 10, 21) {real, imag} */,
  {32'h402428d4, 32'h415ccd4e} /* (13, 10, 20) {real, imag} */,
  {32'h40e456b6, 32'hc12cb7de} /* (13, 10, 19) {real, imag} */,
  {32'hc025a91e, 32'h40ead9f4} /* (13, 10, 18) {real, imag} */,
  {32'hbf856a8e, 32'hc10375c7} /* (13, 10, 17) {real, imag} */,
  {32'h40f08b42, 32'hc00c4870} /* (13, 10, 16) {real, imag} */,
  {32'hbfc267ce, 32'h3f9b371a} /* (13, 10, 15) {real, imag} */,
  {32'hc0ab75e1, 32'hbf29b760} /* (13, 10, 14) {real, imag} */,
  {32'h413adecd, 32'hc0bc8744} /* (13, 10, 13) {real, imag} */,
  {32'hc176a5ef, 32'hc070e1f8} /* (13, 10, 12) {real, imag} */,
  {32'h40e81ac8, 32'hbf06d1f0} /* (13, 10, 11) {real, imag} */,
  {32'h3f7029fe, 32'hc09bb313} /* (13, 10, 10) {real, imag} */,
  {32'hc14d2470, 32'hc14f3cdc} /* (13, 10, 9) {real, imag} */,
  {32'h415e0fe1, 32'h410939fb} /* (13, 10, 8) {real, imag} */,
  {32'h415bc9ab, 32'hc1138f1a} /* (13, 10, 7) {real, imag} */,
  {32'hc0fe9a1a, 32'h41f24f39} /* (13, 10, 6) {real, imag} */,
  {32'hc0581600, 32'h42157ac9} /* (13, 10, 5) {real, imag} */,
  {32'hc154df42, 32'hc233fbe8} /* (13, 10, 4) {real, imag} */,
  {32'h418ebf4e, 32'hbea80df0} /* (13, 10, 3) {real, imag} */,
  {32'hc196cc0a, 32'h41aa3198} /* (13, 10, 2) {real, imag} */,
  {32'hc123f02d, 32'hc12fe73e} /* (13, 10, 1) {real, imag} */,
  {32'h419366d6, 32'hc227e895} /* (13, 10, 0) {real, imag} */,
  {32'hc1f750ce, 32'hc25da62e} /* (13, 9, 31) {real, imag} */,
  {32'h40a895b0, 32'hc1c78fca} /* (13, 9, 30) {real, imag} */,
  {32'hc009894c, 32'h428371b3} /* (13, 9, 29) {real, imag} */,
  {32'hc19d4591, 32'h4185f4d7} /* (13, 9, 28) {real, imag} */,
  {32'h400d74e8, 32'h41c97f7f} /* (13, 9, 27) {real, imag} */,
  {32'hc2192375, 32'h41a0aa10} /* (13, 9, 26) {real, imag} */,
  {32'hc10b7e93, 32'hc1868553} /* (13, 9, 25) {real, imag} */,
  {32'h408e966a, 32'hc20d68ad} /* (13, 9, 24) {real, imag} */,
  {32'h41585ca5, 32'hc1c5b182} /* (13, 9, 23) {real, imag} */,
  {32'h412ce87b, 32'h4198151f} /* (13, 9, 22) {real, imag} */,
  {32'h41c05970, 32'hc0b90bc2} /* (13, 9, 21) {real, imag} */,
  {32'h4062502e, 32'hc1e01b78} /* (13, 9, 20) {real, imag} */,
  {32'hc02540c4, 32'h401ae544} /* (13, 9, 19) {real, imag} */,
  {32'hc13189bc, 32'h3fb3a108} /* (13, 9, 18) {real, imag} */,
  {32'hbff75a48, 32'h40ddca58} /* (13, 9, 17) {real, imag} */,
  {32'h401d3258, 32'hc0691d39} /* (13, 9, 16) {real, imag} */,
  {32'h40a6913a, 32'h40f6fd4c} /* (13, 9, 15) {real, imag} */,
  {32'hc0ba8c88, 32'hc085588e} /* (13, 9, 14) {real, imag} */,
  {32'hbf6d8270, 32'hbfc22218} /* (13, 9, 13) {real, imag} */,
  {32'hbe5d09a0, 32'hc12a3881} /* (13, 9, 12) {real, imag} */,
  {32'h40663d4c, 32'hc020dc9d} /* (13, 9, 11) {real, imag} */,
  {32'hc18b8da8, 32'h3eed3500} /* (13, 9, 10) {real, imag} */,
  {32'h41ba4580, 32'hbf6fa340} /* (13, 9, 9) {real, imag} */,
  {32'h41c34b98, 32'h411fcd90} /* (13, 9, 8) {real, imag} */,
  {32'hc12ab9a5, 32'h40c8e394} /* (13, 9, 7) {real, imag} */,
  {32'hc1c1fa8e, 32'h4157a0e9} /* (13, 9, 6) {real, imag} */,
  {32'hc2143dba, 32'h41d8aa5f} /* (13, 9, 5) {real, imag} */,
  {32'h40928ba7, 32'hc13370b0} /* (13, 9, 4) {real, imag} */,
  {32'hc1c7b2d0, 32'hc19f6624} /* (13, 9, 3) {real, imag} */,
  {32'hc2150173, 32'hc09ee512} /* (13, 9, 2) {real, imag} */,
  {32'h421da2d3, 32'hc0c267f0} /* (13, 9, 1) {real, imag} */,
  {32'hc19e68d3, 32'h407e415d} /* (13, 9, 0) {real, imag} */,
  {32'h4207bcea, 32'hc1119026} /* (13, 8, 31) {real, imag} */,
  {32'hc22e2a27, 32'h41989e8c} /* (13, 8, 30) {real, imag} */,
  {32'h42387eda, 32'hc21d1cc2} /* (13, 8, 29) {real, imag} */,
  {32'h4202c5ae, 32'hc1f0ce1e} /* (13, 8, 28) {real, imag} */,
  {32'h4142eb2c, 32'h40c5c2e4} /* (13, 8, 27) {real, imag} */,
  {32'h420c485e, 32'hc179e0c7} /* (13, 8, 26) {real, imag} */,
  {32'hc13c9e58, 32'h4113208d} /* (13, 8, 25) {real, imag} */,
  {32'h40a6bff8, 32'hc04df824} /* (13, 8, 24) {real, imag} */,
  {32'h4097b20a, 32'hc2002ca4} /* (13, 8, 23) {real, imag} */,
  {32'h40e55844, 32'h411869e2} /* (13, 8, 22) {real, imag} */,
  {32'hc1b2c2f6, 32'h40a095c1} /* (13, 8, 21) {real, imag} */,
  {32'h3f1f4ca8, 32'h414b9657} /* (13, 8, 20) {real, imag} */,
  {32'hc0fc1608, 32'hc14f0468} /* (13, 8, 19) {real, imag} */,
  {32'h3fa67238, 32'h3fafffb4} /* (13, 8, 18) {real, imag} */,
  {32'hbfac5f14, 32'hc0bebebf} /* (13, 8, 17) {real, imag} */,
  {32'h3d97c700, 32'h3de85880} /* (13, 8, 16) {real, imag} */,
  {32'h4047c7aa, 32'h40466802} /* (13, 8, 15) {real, imag} */,
  {32'hc10d5a49, 32'hc0c0141f} /* (13, 8, 14) {real, imag} */,
  {32'hc0cb6350, 32'h4139f41e} /* (13, 8, 13) {real, imag} */,
  {32'h4009096e, 32'h4151304f} /* (13, 8, 12) {real, imag} */,
  {32'hbffbc0e0, 32'hc18b5c5e} /* (13, 8, 11) {real, imag} */,
  {32'h41a2026f, 32'hc1ca077f} /* (13, 8, 10) {real, imag} */,
  {32'hc15600c7, 32'h417b8f56} /* (13, 8, 9) {real, imag} */,
  {32'h3f2a0380, 32'hc189098c} /* (13, 8, 8) {real, imag} */,
  {32'hc0894af9, 32'hc015532c} /* (13, 8, 7) {real, imag} */,
  {32'hc187e65b, 32'hc143768d} /* (13, 8, 6) {real, imag} */,
  {32'hc1a06ec2, 32'h41c2fb2d} /* (13, 8, 5) {real, imag} */,
  {32'hbdab9300, 32'h420eeac7} /* (13, 8, 4) {real, imag} */,
  {32'hc24b45ee, 32'h415c696a} /* (13, 8, 3) {real, imag} */,
  {32'h40707090, 32'hc20818fc} /* (13, 8, 2) {real, imag} */,
  {32'h40b35834, 32'hbf9c2d2c} /* (13, 8, 1) {real, imag} */,
  {32'h422dc21e, 32'hc1a2c810} /* (13, 8, 0) {real, imag} */,
  {32'h41b32a9f, 32'hc186afa8} /* (13, 7, 31) {real, imag} */,
  {32'hc0ef9238, 32'hc1ae0f1a} /* (13, 7, 30) {real, imag} */,
  {32'hc14f44b7, 32'hbfba6f72} /* (13, 7, 29) {real, imag} */,
  {32'h4128b17a, 32'hc14bff33} /* (13, 7, 28) {real, imag} */,
  {32'hc1e33cd1, 32'hc170363d} /* (13, 7, 27) {real, imag} */,
  {32'hbe02c320, 32'hc1ca53fb} /* (13, 7, 26) {real, imag} */,
  {32'hc1bd481c, 32'h4115d4d2} /* (13, 7, 25) {real, imag} */,
  {32'hbf990b00, 32'h40e09a52} /* (13, 7, 24) {real, imag} */,
  {32'hc0b48816, 32'hc1548b2e} /* (13, 7, 23) {real, imag} */,
  {32'h41134ff4, 32'hc12323d9} /* (13, 7, 22) {real, imag} */,
  {32'h41aa851e, 32'h418323b6} /* (13, 7, 21) {real, imag} */,
  {32'hc14ebeb0, 32'h3fd33848} /* (13, 7, 20) {real, imag} */,
  {32'hc18ba264, 32'hbf075904} /* (13, 7, 19) {real, imag} */,
  {32'h40e8be66, 32'hc0aaa63a} /* (13, 7, 18) {real, imag} */,
  {32'hbf37f810, 32'hbdd831a0} /* (13, 7, 17) {real, imag} */,
  {32'h41315920, 32'h40da8302} /* (13, 7, 16) {real, imag} */,
  {32'h3fe30c78, 32'h401ee70b} /* (13, 7, 15) {real, imag} */,
  {32'h40431834, 32'hc14741d1} /* (13, 7, 14) {real, imag} */,
  {32'h3f91e708, 32'h4026cf4b} /* (13, 7, 13) {real, imag} */,
  {32'h40dea38f, 32'h40ef0732} /* (13, 7, 12) {real, imag} */,
  {32'hc1176bec, 32'hc1a66a8e} /* (13, 7, 11) {real, imag} */,
  {32'hc0b57fc3, 32'h418a4268} /* (13, 7, 10) {real, imag} */,
  {32'hbf35b750, 32'h422027aa} /* (13, 7, 9) {real, imag} */,
  {32'hc045946c, 32'hc1a1628e} /* (13, 7, 8) {real, imag} */,
  {32'h422c323e, 32'hc2565212} /* (13, 7, 7) {real, imag} */,
  {32'h41024e22, 32'h4182c681} /* (13, 7, 6) {real, imag} */,
  {32'hc071c658, 32'h42296933} /* (13, 7, 5) {real, imag} */,
  {32'h411e8c4e, 32'hc0e0bfd2} /* (13, 7, 4) {real, imag} */,
  {32'hc1392151, 32'h40b7a262} /* (13, 7, 3) {real, imag} */,
  {32'hc27356bd, 32'h41a434b4} /* (13, 7, 2) {real, imag} */,
  {32'h4220e64a, 32'h417161c7} /* (13, 7, 1) {real, imag} */,
  {32'hc232e4eb, 32'hc1954272} /* (13, 7, 0) {real, imag} */,
  {32'hc234c8af, 32'h416052b6} /* (13, 6, 31) {real, imag} */,
  {32'hc1e6f911, 32'h42410e0a} /* (13, 6, 30) {real, imag} */,
  {32'h414aab26, 32'hc1a349e8} /* (13, 6, 29) {real, imag} */,
  {32'hc1607631, 32'h42032814} /* (13, 6, 28) {real, imag} */,
  {32'h4157b6b0, 32'hc1fc5896} /* (13, 6, 27) {real, imag} */,
  {32'hc1adf493, 32'hc221acd7} /* (13, 6, 26) {real, imag} */,
  {32'hc0c1f204, 32'h419c52d1} /* (13, 6, 25) {real, imag} */,
  {32'hc207ae2b, 32'hc28e892f} /* (13, 6, 24) {real, imag} */,
  {32'h41d53764, 32'hc1d0bce6} /* (13, 6, 23) {real, imag} */,
  {32'hc0f91946, 32'h3f3d7770} /* (13, 6, 22) {real, imag} */,
  {32'h4097c7ee, 32'h40a9d852} /* (13, 6, 21) {real, imag} */,
  {32'hbfc68d7a, 32'hbfb72d3c} /* (13, 6, 20) {real, imag} */,
  {32'h415a5868, 32'h41e04feb} /* (13, 6, 19) {real, imag} */,
  {32'h411e65dc, 32'hc11adda8} /* (13, 6, 18) {real, imag} */,
  {32'hc13154e7, 32'h3fd98830} /* (13, 6, 17) {real, imag} */,
  {32'hc081f41e, 32'h4011bb60} /* (13, 6, 16) {real, imag} */,
  {32'hc14be329, 32'hc18f2043} /* (13, 6, 15) {real, imag} */,
  {32'h41424ef4, 32'h3f2d3f00} /* (13, 6, 14) {real, imag} */,
  {32'h40f106e8, 32'h408b59b4} /* (13, 6, 13) {real, imag} */,
  {32'h409e8226, 32'hc0c8641f} /* (13, 6, 12) {real, imag} */,
  {32'hc16a540d, 32'h4199b06a} /* (13, 6, 11) {real, imag} */,
  {32'hc107a37d, 32'hc19f9360} /* (13, 6, 10) {real, imag} */,
  {32'h41a2cadc, 32'hc193c210} /* (13, 6, 9) {real, imag} */,
  {32'hc1e5cdc2, 32'hc15d07a8} /* (13, 6, 8) {real, imag} */,
  {32'hc109175e, 32'h41d90c89} /* (13, 6, 7) {real, imag} */,
  {32'h41adaf09, 32'h423ebde7} /* (13, 6, 6) {real, imag} */,
  {32'h42395c4e, 32'h40c5e408} /* (13, 6, 5) {real, imag} */,
  {32'hc1dc1b5a, 32'hc10320b2} /* (13, 6, 4) {real, imag} */,
  {32'hc1f9dc89, 32'hc0759120} /* (13, 6, 3) {real, imag} */,
  {32'h427ac746, 32'hc201504c} /* (13, 6, 2) {real, imag} */,
  {32'h40057f50, 32'hc11b0356} /* (13, 6, 1) {real, imag} */,
  {32'h41c27510, 32'h41c2dff2} /* (13, 6, 0) {real, imag} */,
  {32'h40d9e8fc, 32'hc209b17a} /* (13, 5, 31) {real, imag} */,
  {32'h42047a24, 32'hc22dbefa} /* (13, 5, 30) {real, imag} */,
  {32'hc1913925, 32'hc2137600} /* (13, 5, 29) {real, imag} */,
  {32'hc1acccf4, 32'h41e6b030} /* (13, 5, 28) {real, imag} */,
  {32'hc1973909, 32'h3fff2de6} /* (13, 5, 27) {real, imag} */,
  {32'h3fbd0fc0, 32'h4159487c} /* (13, 5, 26) {real, imag} */,
  {32'hc1d126ce, 32'hc1657302} /* (13, 5, 25) {real, imag} */,
  {32'hc1f107ca, 32'h41cae5c2} /* (13, 5, 24) {real, imag} */,
  {32'h3f11f040, 32'h4115981b} /* (13, 5, 23) {real, imag} */,
  {32'hc21cc9b6, 32'hc1f8a5ab} /* (13, 5, 22) {real, imag} */,
  {32'hc20b3fed, 32'h419e0ca8} /* (13, 5, 21) {real, imag} */,
  {32'hc07efdae, 32'hc1243f78} /* (13, 5, 20) {real, imag} */,
  {32'hc1731474, 32'hc08eb9ef} /* (13, 5, 19) {real, imag} */,
  {32'hc041f356, 32'hc0418884} /* (13, 5, 18) {real, imag} */,
  {32'hc0f99c6e, 32'h40981550} /* (13, 5, 17) {real, imag} */,
  {32'h4148b368, 32'h4083a96c} /* (13, 5, 16) {real, imag} */,
  {32'h3fb611f0, 32'h410215e4} /* (13, 5, 15) {real, imag} */,
  {32'h4157e6fa, 32'hbef34fa0} /* (13, 5, 14) {real, imag} */,
  {32'h406ae5c0, 32'hc09d5957} /* (13, 5, 13) {real, imag} */,
  {32'hc13cfe16, 32'hc15f8974} /* (13, 5, 12) {real, imag} */,
  {32'hc209b9db, 32'hc1614aff} /* (13, 5, 11) {real, imag} */,
  {32'hc124df38, 32'hc08427ec} /* (13, 5, 10) {real, imag} */,
  {32'hc1a3d982, 32'h404f2174} /* (13, 5, 9) {real, imag} */,
  {32'h4217798f, 32'hc172db4d} /* (13, 5, 8) {real, imag} */,
  {32'hc287f624, 32'hc21341d4} /* (13, 5, 7) {real, imag} */,
  {32'h42bbe5cf, 32'h401ff71e} /* (13, 5, 6) {real, imag} */,
  {32'h404b8b28, 32'h3cfd1980} /* (13, 5, 5) {real, imag} */,
  {32'h4185a212, 32'h40290000} /* (13, 5, 4) {real, imag} */,
  {32'h429cd1a7, 32'h4104e18e} /* (13, 5, 3) {real, imag} */,
  {32'h4075a1b8, 32'h42623ce6} /* (13, 5, 2) {real, imag} */,
  {32'hc1ec5dd7, 32'h42248796} /* (13, 5, 1) {real, imag} */,
  {32'h424c4466, 32'hc16a7796} /* (13, 5, 0) {real, imag} */,
  {32'h4174b59a, 32'hc2220750} /* (13, 4, 31) {real, imag} */,
  {32'hc1f49b78, 32'h4255440a} /* (13, 4, 30) {real, imag} */,
  {32'h41c2211a, 32'h4126a045} /* (13, 4, 29) {real, imag} */,
  {32'h42083a76, 32'hc20e8068} /* (13, 4, 28) {real, imag} */,
  {32'hc201d55f, 32'hc2163c94} /* (13, 4, 27) {real, imag} */,
  {32'hc026f8bb, 32'h41c57bcd} /* (13, 4, 26) {real, imag} */,
  {32'h413f485b, 32'hc1572556} /* (13, 4, 25) {real, imag} */,
  {32'h4157aa8a, 32'hc141cbee} /* (13, 4, 24) {real, imag} */,
  {32'h412d0ba7, 32'hc1b6d01e} /* (13, 4, 23) {real, imag} */,
  {32'h40e8644e, 32'hc05d3178} /* (13, 4, 22) {real, imag} */,
  {32'h409208a4, 32'h40be9ca8} /* (13, 4, 21) {real, imag} */,
  {32'hc14aa7fb, 32'hc0dc2734} /* (13, 4, 20) {real, imag} */,
  {32'h40e17ae1, 32'hc0ab22a4} /* (13, 4, 19) {real, imag} */,
  {32'h3f78c2aa, 32'hc1a77ab1} /* (13, 4, 18) {real, imag} */,
  {32'hc10136d2, 32'h40ddc850} /* (13, 4, 17) {real, imag} */,
  {32'h40e0318e, 32'h4014ea70} /* (13, 4, 16) {real, imag} */,
  {32'hbfc675b4, 32'h4031ded0} /* (13, 4, 15) {real, imag} */,
  {32'h402deb7a, 32'h40980ec0} /* (13, 4, 14) {real, imag} */,
  {32'h41813513, 32'h4144d988} /* (13, 4, 13) {real, imag} */,
  {32'hbeef4860, 32'hc12e486a} /* (13, 4, 12) {real, imag} */,
  {32'h4027d608, 32'hc14b2d94} /* (13, 4, 11) {real, imag} */,
  {32'hc14eede9, 32'h41a9288d} /* (13, 4, 10) {real, imag} */,
  {32'h410a3239, 32'hbe7d9040} /* (13, 4, 9) {real, imag} */,
  {32'hbe818f80, 32'hc21a2134} /* (13, 4, 8) {real, imag} */,
  {32'h4181487e, 32'hc15212ea} /* (13, 4, 7) {real, imag} */,
  {32'hc06df71b, 32'hc15a1c62} /* (13, 4, 6) {real, imag} */,
  {32'h400f8720, 32'hc22526ee} /* (13, 4, 5) {real, imag} */,
  {32'hc22b0d6c, 32'h42bd0410} /* (13, 4, 4) {real, imag} */,
  {32'hc05f9aec, 32'h41fd3a7e} /* (13, 4, 3) {real, imag} */,
  {32'h41ff86f6, 32'hc02ab660} /* (13, 4, 2) {real, imag} */,
  {32'h417dfb86, 32'h4214c260} /* (13, 4, 1) {real, imag} */,
  {32'h419f657a, 32'hc26701c5} /* (13, 4, 0) {real, imag} */,
  {32'hc16d60ca, 32'h415345e9} /* (13, 3, 31) {real, imag} */,
  {32'hc1f38fd1, 32'hc1fc867e} /* (13, 3, 30) {real, imag} */,
  {32'hc14c00aa, 32'hc27ef4cd} /* (13, 3, 29) {real, imag} */,
  {32'h41992750, 32'hc1257892} /* (13, 3, 28) {real, imag} */,
  {32'hc005db36, 32'hc16ffc52} /* (13, 3, 27) {real, imag} */,
  {32'hc085116e, 32'h42558f00} /* (13, 3, 26) {real, imag} */,
  {32'h41ee4b2f, 32'h402a47b8} /* (13, 3, 25) {real, imag} */,
  {32'hc132e930, 32'h3e6baf00} /* (13, 3, 24) {real, imag} */,
  {32'h40caac34, 32'hbf804a94} /* (13, 3, 23) {real, imag} */,
  {32'h410b60db, 32'hc1e3e1ca} /* (13, 3, 22) {real, imag} */,
  {32'hc0500b9c, 32'hc02c0173} /* (13, 3, 21) {real, imag} */,
  {32'hc1711172, 32'h40f3e84a} /* (13, 3, 20) {real, imag} */,
  {32'hbebe7848, 32'h418367ea} /* (13, 3, 19) {real, imag} */,
  {32'hc01827f0, 32'h41448004} /* (13, 3, 18) {real, imag} */,
  {32'hc0ec2b3b, 32'h3f6e25e4} /* (13, 3, 17) {real, imag} */,
  {32'hc0fbfc2c, 32'hc03e02ae} /* (13, 3, 16) {real, imag} */,
  {32'h40871fab, 32'hc09708a4} /* (13, 3, 15) {real, imag} */,
  {32'hc1ba4e48, 32'hc0b17250} /* (13, 3, 14) {real, imag} */,
  {32'h4087af02, 32'h419164c6} /* (13, 3, 13) {real, imag} */,
  {32'h40a84f28, 32'h40c2db3a} /* (13, 3, 12) {real, imag} */,
  {32'hc19ff200, 32'h40710f3d} /* (13, 3, 11) {real, imag} */,
  {32'h40417a7d, 32'h41a287ca} /* (13, 3, 10) {real, imag} */,
  {32'h41d01c0d, 32'hc110b7ba} /* (13, 3, 9) {real, imag} */,
  {32'hc124082c, 32'h42618739} /* (13, 3, 8) {real, imag} */,
  {32'h40de330c, 32'h41ee1d0b} /* (13, 3, 7) {real, imag} */,
  {32'hc1233aa7, 32'h4117ff88} /* (13, 3, 6) {real, imag} */,
  {32'hc153e4a4, 32'h41c80f21} /* (13, 3, 5) {real, imag} */,
  {32'h4218d848, 32'h41c9e4d7} /* (13, 3, 4) {real, imag} */,
  {32'hc1b24e63, 32'hc04e1f70} /* (13, 3, 3) {real, imag} */,
  {32'hc20a07c7, 32'h41626e38} /* (13, 3, 2) {real, imag} */,
  {32'hc1e02977, 32'hc1d11260} /* (13, 3, 1) {real, imag} */,
  {32'hc2274ae4, 32'hbe7e2ca0} /* (13, 3, 0) {real, imag} */,
  {32'hc1d12ce9, 32'h41f17230} /* (13, 2, 31) {real, imag} */,
  {32'h426d9666, 32'h429ec4be} /* (13, 2, 30) {real, imag} */,
  {32'h42acb6a7, 32'hc1db8910} /* (13, 2, 29) {real, imag} */,
  {32'h4267c22e, 32'h41aeb67c} /* (13, 2, 28) {real, imag} */,
  {32'hc25fe6d0, 32'h408720fc} /* (13, 2, 27) {real, imag} */,
  {32'hc0ce2a80, 32'hc28986ae} /* (13, 2, 26) {real, imag} */,
  {32'h41f4e828, 32'hc15a3aa0} /* (13, 2, 25) {real, imag} */,
  {32'hc2103480, 32'hc2150106} /* (13, 2, 24) {real, imag} */,
  {32'h4175ae69, 32'h42123e1c} /* (13, 2, 23) {real, imag} */,
  {32'hc1ee4a72, 32'hc109b2bd} /* (13, 2, 22) {real, imag} */,
  {32'hc1deef58, 32'h41295c2a} /* (13, 2, 21) {real, imag} */,
  {32'hc078a498, 32'h41024f20} /* (13, 2, 20) {real, imag} */,
  {32'hc1095f7e, 32'h40d303b7} /* (13, 2, 19) {real, imag} */,
  {32'h41839c9f, 32'h4155d1ec} /* (13, 2, 18) {real, imag} */,
  {32'hc0029888, 32'hc0be8b38} /* (13, 2, 17) {real, imag} */,
  {32'h40b148dc, 32'h3fa3e6d8} /* (13, 2, 16) {real, imag} */,
  {32'h4164df02, 32'hc11ed1fc} /* (13, 2, 15) {real, imag} */,
  {32'h41143d06, 32'h419fe072} /* (13, 2, 14) {real, imag} */,
  {32'hbfb42e10, 32'hc1893b3c} /* (13, 2, 13) {real, imag} */,
  {32'hc19b7f35, 32'hc1b0e660} /* (13, 2, 12) {real, imag} */,
  {32'h3fc76f78, 32'h418bb919} /* (13, 2, 11) {real, imag} */,
  {32'hc10d1ce4, 32'h407b1434} /* (13, 2, 10) {real, imag} */,
  {32'hc1bd2ed2, 32'hc130871c} /* (13, 2, 9) {real, imag} */,
  {32'hc255adae, 32'h4205816e} /* (13, 2, 8) {real, imag} */,
  {32'hc18ee4c6, 32'hc1f3459e} /* (13, 2, 7) {real, imag} */,
  {32'hc236a86c, 32'hc1efa946} /* (13, 2, 6) {real, imag} */,
  {32'hc1b799a0, 32'hc269a9aa} /* (13, 2, 5) {real, imag} */,
  {32'h4109dac6, 32'h42826a2d} /* (13, 2, 4) {real, imag} */,
  {32'h41c5c003, 32'hc101fc64} /* (13, 2, 3) {real, imag} */,
  {32'hc1e45859, 32'h426647bd} /* (13, 2, 2) {real, imag} */,
  {32'h4211e092, 32'hc2c23ad2} /* (13, 2, 1) {real, imag} */,
  {32'h42836aef, 32'h416f48bf} /* (13, 2, 0) {real, imag} */,
  {32'h428355ff, 32'h419bcb1f} /* (13, 1, 31) {real, imag} */,
  {32'h421ab010, 32'h41e082cf} /* (13, 1, 30) {real, imag} */,
  {32'h42c3cca7, 32'h41205c62} /* (13, 1, 29) {real, imag} */,
  {32'h4190f338, 32'hc04e5080} /* (13, 1, 28) {real, imag} */,
  {32'hc18e4b49, 32'h4259f97c} /* (13, 1, 27) {real, imag} */,
  {32'h4191a471, 32'h40709518} /* (13, 1, 26) {real, imag} */,
  {32'h414112ac, 32'h41daea74} /* (13, 1, 25) {real, imag} */,
  {32'h42101195, 32'h422c4078} /* (13, 1, 24) {real, imag} */,
  {32'h4130ee5a, 32'h41fecf0c} /* (13, 1, 23) {real, imag} */,
  {32'h41754de4, 32'h408e50e8} /* (13, 1, 22) {real, imag} */,
  {32'hc17f26a4, 32'h40c3247a} /* (13, 1, 21) {real, imag} */,
  {32'hc20f09d0, 32'h409075ab} /* (13, 1, 20) {real, imag} */,
  {32'h41169e28, 32'h3f86998c} /* (13, 1, 19) {real, imag} */,
  {32'h4039d6c2, 32'h40fee6d0} /* (13, 1, 18) {real, imag} */,
  {32'hc15e9898, 32'hbfce7d58} /* (13, 1, 17) {real, imag} */,
  {32'h41945099, 32'hc1f0762a} /* (13, 1, 16) {real, imag} */,
  {32'hc05a1b00, 32'h40fc1b90} /* (13, 1, 15) {real, imag} */,
  {32'h4022b69a, 32'hc153c7d4} /* (13, 1, 14) {real, imag} */,
  {32'h40ae2d58, 32'hc035f39a} /* (13, 1, 13) {real, imag} */,
  {32'hc110ccb0, 32'hc10c7944} /* (13, 1, 12) {real, imag} */,
  {32'h424b101b, 32'hc01813dc} /* (13, 1, 11) {real, imag} */,
  {32'h4161840c, 32'h40fc6b4c} /* (13, 1, 10) {real, imag} */,
  {32'hc1aab0e3, 32'hc295ce25} /* (13, 1, 9) {real, imag} */,
  {32'hc15316dc, 32'h402d40a8} /* (13, 1, 8) {real, imag} */,
  {32'hc1fb0602, 32'hc0c1d230} /* (13, 1, 7) {real, imag} */,
  {32'h42048814, 32'h40c4c7ac} /* (13, 1, 6) {real, imag} */,
  {32'hc1a02c73, 32'h40f85674} /* (13, 1, 5) {real, imag} */,
  {32'hc1304500, 32'h42201a04} /* (13, 1, 4) {real, imag} */,
  {32'h418b0954, 32'hc2000aac} /* (13, 1, 3) {real, imag} */,
  {32'hc180ed1c, 32'h42775b3c} /* (13, 1, 2) {real, imag} */,
  {32'hc28d9a11, 32'hc0a786bb} /* (13, 1, 1) {real, imag} */,
  {32'h423cd08e, 32'h41a86d96} /* (13, 1, 0) {real, imag} */,
  {32'hc244a753, 32'h413c05e8} /* (13, 0, 31) {real, imag} */,
  {32'h425006d0, 32'h422b453e} /* (13, 0, 30) {real, imag} */,
  {32'h411f4130, 32'hc29c8ba0} /* (13, 0, 29) {real, imag} */,
  {32'h41133f01, 32'h425952aa} /* (13, 0, 28) {real, imag} */,
  {32'hc1fd0802, 32'hc0c36c1a} /* (13, 0, 27) {real, imag} */,
  {32'hc1c40cfa, 32'hc1bafeca} /* (13, 0, 26) {real, imag} */,
  {32'hc1fc47ea, 32'hc0b024c2} /* (13, 0, 25) {real, imag} */,
  {32'hc20a6b1c, 32'h42264f5f} /* (13, 0, 24) {real, imag} */,
  {32'h42510d8e, 32'hc08dec56} /* (13, 0, 23) {real, imag} */,
  {32'hc183d93c, 32'h4216e713} /* (13, 0, 22) {real, imag} */,
  {32'h423e5785, 32'hc18d2ca8} /* (13, 0, 21) {real, imag} */,
  {32'hc182640a, 32'h40972cc6} /* (13, 0, 20) {real, imag} */,
  {32'hc18f230d, 32'h410e4a17} /* (13, 0, 19) {real, imag} */,
  {32'h3ffce298, 32'h40b8a8d9} /* (13, 0, 18) {real, imag} */,
  {32'h4172ddad, 32'hc0a14d70} /* (13, 0, 17) {real, imag} */,
  {32'hc19ebea2, 32'h419b8b0d} /* (13, 0, 16) {real, imag} */,
  {32'hbff91998, 32'hc008c230} /* (13, 0, 15) {real, imag} */,
  {32'h3eaf2760, 32'h3f9197c4} /* (13, 0, 14) {real, imag} */,
  {32'h40a048d4, 32'h40830e4a} /* (13, 0, 13) {real, imag} */,
  {32'h40b7e6b2, 32'hc0988ff2} /* (13, 0, 12) {real, imag} */,
  {32'h4120acb0, 32'h412bf725} /* (13, 0, 11) {real, imag} */,
  {32'hc1dcb7a0, 32'hc18affcc} /* (13, 0, 10) {real, imag} */,
  {32'h3f8f91a0, 32'hc17b145b} /* (13, 0, 9) {real, imag} */,
  {32'hc1ba6ced, 32'h4075d840} /* (13, 0, 8) {real, imag} */,
  {32'hc14c5098, 32'h41cf34be} /* (13, 0, 7) {real, imag} */,
  {32'hc240ff91, 32'hc1de28e8} /* (13, 0, 6) {real, imag} */,
  {32'h400abfa0, 32'hc1c68406} /* (13, 0, 5) {real, imag} */,
  {32'h41daa25c, 32'hc269a50a} /* (13, 0, 4) {real, imag} */,
  {32'h422ad396, 32'hc20c947d} /* (13, 0, 3) {real, imag} */,
  {32'hc0f27e74, 32'hc20e2426} /* (13, 0, 2) {real, imag} */,
  {32'h41a0cb7a, 32'hc298099b} /* (13, 0, 1) {real, imag} */,
  {32'hc0d19e62, 32'hbf990f30} /* (13, 0, 0) {real, imag} */,
  {32'hc2967151, 32'h41c40f14} /* (12, 31, 31) {real, imag} */,
  {32'hc2a2b510, 32'h40e25b8d} /* (12, 31, 30) {real, imag} */,
  {32'hc210b7a4, 32'hc1d27d33} /* (12, 31, 29) {real, imag} */,
  {32'h402091e8, 32'hc27102e6} /* (12, 31, 28) {real, imag} */,
  {32'hc1440f2a, 32'h4168d44b} /* (12, 31, 27) {real, imag} */,
  {32'hc286789e, 32'hbfddd920} /* (12, 31, 26) {real, imag} */,
  {32'h42163420, 32'h428b13e6} /* (12, 31, 25) {real, imag} */,
  {32'hc1f837c5, 32'h41308fb3} /* (12, 31, 24) {real, imag} */,
  {32'hc0e91ccc, 32'h4128adb5} /* (12, 31, 23) {real, imag} */,
  {32'hc1f701cc, 32'hc14dd36c} /* (12, 31, 22) {real, imag} */,
  {32'h422dadb2, 32'hc13bbbc8} /* (12, 31, 21) {real, imag} */,
  {32'h3fe84380, 32'hc0a23d7e} /* (12, 31, 20) {real, imag} */,
  {32'h4091d598, 32'h419b58ba} /* (12, 31, 19) {real, imag} */,
  {32'h41b56a59, 32'h40f6e921} /* (12, 31, 18) {real, imag} */,
  {32'hc108f3f0, 32'h4064b118} /* (12, 31, 17) {real, imag} */,
  {32'hbd0ddc00, 32'hc122eb34} /* (12, 31, 16) {real, imag} */,
  {32'hc1ae7d66, 32'h4196c1ff} /* (12, 31, 15) {real, imag} */,
  {32'h3eaada40, 32'h3f23ccf8} /* (12, 31, 14) {real, imag} */,
  {32'h418eb496, 32'h4202ff30} /* (12, 31, 13) {real, imag} */,
  {32'h40f48bc2, 32'hc0b8c476} /* (12, 31, 12) {real, imag} */,
  {32'hc187ed2f, 32'h425b4cac} /* (12, 31, 11) {real, imag} */,
  {32'h421afefa, 32'hc0f624fc} /* (12, 31, 10) {real, imag} */,
  {32'h422ff1b2, 32'h4042511c} /* (12, 31, 9) {real, imag} */,
  {32'h41e8fb15, 32'h41056a99} /* (12, 31, 8) {real, imag} */,
  {32'hc18b7cfb, 32'h4176c98c} /* (12, 31, 7) {real, imag} */,
  {32'h418bbb7a, 32'h420d0d5b} /* (12, 31, 6) {real, imag} */,
  {32'h424c33b0, 32'hc2078deb} /* (12, 31, 5) {real, imag} */,
  {32'hc1f44a9b, 32'hc0cc5364} /* (12, 31, 4) {real, imag} */,
  {32'h42020460, 32'h416679fa} /* (12, 31, 3) {real, imag} */,
  {32'hc0711300, 32'h419f8579} /* (12, 31, 2) {real, imag} */,
  {32'hc218ae52, 32'hc11d7160} /* (12, 31, 1) {real, imag} */,
  {32'h4230e4db, 32'h42134f86} /* (12, 31, 0) {real, imag} */,
  {32'hc1b2582b, 32'hc1494ad4} /* (12, 30, 31) {real, imag} */,
  {32'hc26c803e, 32'h41a26fb8} /* (12, 30, 30) {real, imag} */,
  {32'h4228863a, 32'h4208be41} /* (12, 30, 29) {real, imag} */,
  {32'h41096464, 32'hc1920623} /* (12, 30, 28) {real, imag} */,
  {32'h420b3e31, 32'hc1aadd2d} /* (12, 30, 27) {real, imag} */,
  {32'h41a6f16e, 32'hc0571e78} /* (12, 30, 26) {real, imag} */,
  {32'h420a7a81, 32'h4234483f} /* (12, 30, 25) {real, imag} */,
  {32'h41b339fe, 32'h40e9ab35} /* (12, 30, 24) {real, imag} */,
  {32'h41db5c19, 32'h40df6792} /* (12, 30, 23) {real, imag} */,
  {32'hc0e6d228, 32'h40437b90} /* (12, 30, 22) {real, imag} */,
  {32'hc1c96da2, 32'h40a1ae0c} /* (12, 30, 21) {real, imag} */,
  {32'h4210c0db, 32'h41cbe5ca} /* (12, 30, 20) {real, imag} */,
  {32'hc0f178e6, 32'hc0990aec} /* (12, 30, 19) {real, imag} */,
  {32'hc1878150, 32'h41125f24} /* (12, 30, 18) {real, imag} */,
  {32'hc115ba30, 32'h40487010} /* (12, 30, 17) {real, imag} */,
  {32'hc1133fa6, 32'hc13dd3c9} /* (12, 30, 16) {real, imag} */,
  {32'h4116d29c, 32'hc135a2cc} /* (12, 30, 15) {real, imag} */,
  {32'h415c412b, 32'hc1418702} /* (12, 30, 14) {real, imag} */,
  {32'hc110c4a5, 32'h40040707} /* (12, 30, 13) {real, imag} */,
  {32'h40d86208, 32'hbffe3f18} /* (12, 30, 12) {real, imag} */,
  {32'hbfb28d90, 32'h415278e2} /* (12, 30, 11) {real, imag} */,
  {32'hbf968cb0, 32'h40ad53ce} /* (12, 30, 10) {real, imag} */,
  {32'hc12e4afe, 32'h41a72802} /* (12, 30, 9) {real, imag} */,
  {32'hc0d222ed, 32'hc02b23b2} /* (12, 30, 8) {real, imag} */,
  {32'h42a11acc, 32'hc1869d34} /* (12, 30, 7) {real, imag} */,
  {32'h41f5041a, 32'h41a28595} /* (12, 30, 6) {real, imag} */,
  {32'h42009e99, 32'hc1b5b21f} /* (12, 30, 5) {real, imag} */,
  {32'h3fb43b14, 32'hc257f5cc} /* (12, 30, 4) {real, imag} */,
  {32'h42987cd0, 32'hc25017d9} /* (12, 30, 3) {real, imag} */,
  {32'hc1c48315, 32'h401d80e4} /* (12, 30, 2) {real, imag} */,
  {32'h4233d0a6, 32'h43053a3a} /* (12, 30, 1) {real, imag} */,
  {32'h41611dda, 32'hc2271ca0} /* (12, 30, 0) {real, imag} */,
  {32'h4141b302, 32'h4301c2bd} /* (12, 29, 31) {real, imag} */,
  {32'h4251410b, 32'hc1a0ac20} /* (12, 29, 30) {real, imag} */,
  {32'h4240fe1e, 32'hc25505ea} /* (12, 29, 29) {real, imag} */,
  {32'h42274c3c, 32'hc2100140} /* (12, 29, 28) {real, imag} */,
  {32'h40bfbafa, 32'h415f09e4} /* (12, 29, 27) {real, imag} */,
  {32'hc052e726, 32'h40381568} /* (12, 29, 26) {real, imag} */,
  {32'hc093e394, 32'hc1b416a6} /* (12, 29, 25) {real, imag} */,
  {32'h420daa80, 32'h41c95422} /* (12, 29, 24) {real, imag} */,
  {32'h41b4d338, 32'hc191baf8} /* (12, 29, 23) {real, imag} */,
  {32'hc0a754ec, 32'h4238dd26} /* (12, 29, 22) {real, imag} */,
  {32'hc0a2b904, 32'h40215dde} /* (12, 29, 21) {real, imag} */,
  {32'hc0ce242a, 32'hc1d11cbd} /* (12, 29, 20) {real, imag} */,
  {32'hc1d4b3ce, 32'h412162f8} /* (12, 29, 19) {real, imag} */,
  {32'h4068627a, 32'h40196b00} /* (12, 29, 18) {real, imag} */,
  {32'hc198f64b, 32'h41abca4c} /* (12, 29, 17) {real, imag} */,
  {32'h403f083c, 32'h40ad7157} /* (12, 29, 16) {real, imag} */,
  {32'hbf818870, 32'hc0a0165e} /* (12, 29, 15) {real, imag} */,
  {32'hc0ea52fd, 32'hc16bde98} /* (12, 29, 14) {real, imag} */,
  {32'hc0e67350, 32'hc10d4d98} /* (12, 29, 13) {real, imag} */,
  {32'h418868ae, 32'hc0cb1d0c} /* (12, 29, 12) {real, imag} */,
  {32'h3c9eb000, 32'hc10bc22a} /* (12, 29, 11) {real, imag} */,
  {32'hc211d986, 32'h41883252} /* (12, 29, 10) {real, imag} */,
  {32'hc0da6118, 32'h3f313f50} /* (12, 29, 9) {real, imag} */,
  {32'hc1e663f8, 32'hc0dd3ef0} /* (12, 29, 8) {real, imag} */,
  {32'h41adaa8f, 32'hc28001d8} /* (12, 29, 7) {real, imag} */,
  {32'h40b30e4b, 32'hc1fe2def} /* (12, 29, 6) {real, imag} */,
  {32'hc1d076a6, 32'hc0e7a043} /* (12, 29, 5) {real, imag} */,
  {32'h4218e52e, 32'h427ca830} /* (12, 29, 4) {real, imag} */,
  {32'hc189feb5, 32'hc2e99495} /* (12, 29, 3) {real, imag} */,
  {32'h41e4cc6e, 32'h419b2150} /* (12, 29, 2) {real, imag} */,
  {32'h41940647, 32'hc28c643a} /* (12, 29, 1) {real, imag} */,
  {32'h413ddd3f, 32'hc0cafd35} /* (12, 29, 0) {real, imag} */,
  {32'hc1745042, 32'h41b34316} /* (12, 28, 31) {real, imag} */,
  {32'hc240c5f9, 32'h41d73330} /* (12, 28, 30) {real, imag} */,
  {32'hc13ef348, 32'hc23922df} /* (12, 28, 29) {real, imag} */,
  {32'h411aa442, 32'h41d16654} /* (12, 28, 28) {real, imag} */,
  {32'hc2460848, 32'hc0a59368} /* (12, 28, 27) {real, imag} */,
  {32'hc018ab98, 32'h4191cc2a} /* (12, 28, 26) {real, imag} */,
  {32'h40fb45ee, 32'hc20e7933} /* (12, 28, 25) {real, imag} */,
  {32'hc1bfb2f0, 32'hc16cff80} /* (12, 28, 24) {real, imag} */,
  {32'h40d52c82, 32'hc24140e8} /* (12, 28, 23) {real, imag} */,
  {32'hc238aa86, 32'h41c104f8} /* (12, 28, 22) {real, imag} */,
  {32'hc049d940, 32'h410aad3c} /* (12, 28, 21) {real, imag} */,
  {32'h414602f3, 32'hbffcc3d4} /* (12, 28, 20) {real, imag} */,
  {32'hc1685fb9, 32'h41596314} /* (12, 28, 19) {real, imag} */,
  {32'h41262f0b, 32'h401ce264} /* (12, 28, 18) {real, imag} */,
  {32'h40e88ac7, 32'h40abfec0} /* (12, 28, 17) {real, imag} */,
  {32'hc04ed36c, 32'hc082df00} /* (12, 28, 16) {real, imag} */,
  {32'h40d81a03, 32'h412b5204} /* (12, 28, 15) {real, imag} */,
  {32'h40a127ce, 32'hc1b2c29c} /* (12, 28, 14) {real, imag} */,
  {32'h40ba77c2, 32'h3fbd4920} /* (12, 28, 13) {real, imag} */,
  {32'hc1667447, 32'hc0b00097} /* (12, 28, 12) {real, imag} */,
  {32'hc21d9fe8, 32'h412497a4} /* (12, 28, 11) {real, imag} */,
  {32'h41957581, 32'h41b92c28} /* (12, 28, 10) {real, imag} */,
  {32'h42001a50, 32'h41722d48} /* (12, 28, 9) {real, imag} */,
  {32'hc2241a4c, 32'h4224f2cc} /* (12, 28, 8) {real, imag} */,
  {32'h413096c1, 32'hc0a9b1e8} /* (12, 28, 7) {real, imag} */,
  {32'h42369c14, 32'hc1b652ae} /* (12, 28, 6) {real, imag} */,
  {32'h3f0a0600, 32'hc290595e} /* (12, 28, 5) {real, imag} */,
  {32'hc195de12, 32'h41232a70} /* (12, 28, 4) {real, imag} */,
  {32'hc26297c0, 32'hc0995458} /* (12, 28, 3) {real, imag} */,
  {32'h4210b3cb, 32'h41f97558} /* (12, 28, 2) {real, imag} */,
  {32'h41b283a3, 32'h4102ed61} /* (12, 28, 1) {real, imag} */,
  {32'h41748423, 32'h42456c40} /* (12, 28, 0) {real, imag} */,
  {32'h41d5978b, 32'hc24f8085} /* (12, 27, 31) {real, imag} */,
  {32'hc20745ad, 32'h3decc440} /* (12, 27, 30) {real, imag} */,
  {32'hc1b227ce, 32'h41241475} /* (12, 27, 29) {real, imag} */,
  {32'hc12a8280, 32'hc23e9fb0} /* (12, 27, 28) {real, imag} */,
  {32'hc20bf0d0, 32'hc2438245} /* (12, 27, 27) {real, imag} */,
  {32'hc2058488, 32'hc1c6b86f} /* (12, 27, 26) {real, imag} */,
  {32'h421579d2, 32'h42051716} /* (12, 27, 25) {real, imag} */,
  {32'hc01e3080, 32'h424965a0} /* (12, 27, 24) {real, imag} */,
  {32'hc1dee443, 32'hc1a5a288} /* (12, 27, 23) {real, imag} */,
  {32'hc185d7e2, 32'h40b9220d} /* (12, 27, 22) {real, imag} */,
  {32'h41bca24e, 32'hc0a599f0} /* (12, 27, 21) {real, imag} */,
  {32'hbfaa7fcc, 32'h411117ba} /* (12, 27, 20) {real, imag} */,
  {32'h3fdd78f0, 32'hc130b69a} /* (12, 27, 19) {real, imag} */,
  {32'h3f7b8710, 32'hc0c48a45} /* (12, 27, 18) {real, imag} */,
  {32'hbfd3df18, 32'hc132d18d} /* (12, 27, 17) {real, imag} */,
  {32'hc15898c2, 32'hc0293b64} /* (12, 27, 16) {real, imag} */,
  {32'h40a6a39a, 32'hbf5216b0} /* (12, 27, 15) {real, imag} */,
  {32'hc1270463, 32'hc090c23f} /* (12, 27, 14) {real, imag} */,
  {32'h40bb018c, 32'h40bc9f60} /* (12, 27, 13) {real, imag} */,
  {32'hc04c7ce2, 32'hc1940849} /* (12, 27, 12) {real, imag} */,
  {32'hc1a7cffa, 32'h421a1cb0} /* (12, 27, 11) {real, imag} */,
  {32'hc12af941, 32'h40874a7b} /* (12, 27, 10) {real, imag} */,
  {32'h41dfd95f, 32'hc22e80a0} /* (12, 27, 9) {real, imag} */,
  {32'hc248a42e, 32'h41688a0e} /* (12, 27, 8) {real, imag} */,
  {32'hc16c9ba5, 32'hc0f0c6f4} /* (12, 27, 7) {real, imag} */,
  {32'hc129a11d, 32'hc24e09b0} /* (12, 27, 6) {real, imag} */,
  {32'h4189fd8f, 32'hc200789d} /* (12, 27, 5) {real, imag} */,
  {32'hc1a9373b, 32'hc07382e8} /* (12, 27, 4) {real, imag} */,
  {32'hc2771111, 32'h42197907} /* (12, 27, 3) {real, imag} */,
  {32'h403e7b3c, 32'h414c9a02} /* (12, 27, 2) {real, imag} */,
  {32'h41d2775d, 32'h3fa0cfe0} /* (12, 27, 1) {real, imag} */,
  {32'h41e65c8d, 32'hc177df6f} /* (12, 27, 0) {real, imag} */,
  {32'hc1e8409a, 32'h426c382e} /* (12, 26, 31) {real, imag} */,
  {32'h41cfb551, 32'h3f5f2170} /* (12, 26, 30) {real, imag} */,
  {32'h42645546, 32'h41b97037} /* (12, 26, 29) {real, imag} */,
  {32'hc1524626, 32'hc294095b} /* (12, 26, 28) {real, imag} */,
  {32'h408d6e9c, 32'h419ae324} /* (12, 26, 27) {real, imag} */,
  {32'h40457a20, 32'hc1a0f5df} /* (12, 26, 26) {real, imag} */,
  {32'h425192de, 32'hbfb41970} /* (12, 26, 25) {real, imag} */,
  {32'hc1c2fe88, 32'h417b798c} /* (12, 26, 24) {real, imag} */,
  {32'hc1aa1f53, 32'h4165c14c} /* (12, 26, 23) {real, imag} */,
  {32'h40cbe890, 32'hc08bd5ec} /* (12, 26, 22) {real, imag} */,
  {32'hc101ab82, 32'hc0159e62} /* (12, 26, 21) {real, imag} */,
  {32'h4165d1ca, 32'h411cca43} /* (12, 26, 20) {real, imag} */,
  {32'h40be275a, 32'hc0cf61df} /* (12, 26, 19) {real, imag} */,
  {32'h4149c174, 32'h3eec4290} /* (12, 26, 18) {real, imag} */,
  {32'hc11dcef3, 32'h412df1fc} /* (12, 26, 17) {real, imag} */,
  {32'hbef56060, 32'hc0bf9368} /* (12, 26, 16) {real, imag} */,
  {32'h412203e5, 32'hc0cea330} /* (12, 26, 15) {real, imag} */,
  {32'h40409d40, 32'h417729ae} /* (12, 26, 14) {real, imag} */,
  {32'h41a176b8, 32'hbf86c224} /* (12, 26, 13) {real, imag} */,
  {32'hc0f2271d, 32'h41a60ec4} /* (12, 26, 12) {real, imag} */,
  {32'hc0d8ac84, 32'hc14100ea} /* (12, 26, 11) {real, imag} */,
  {32'h4098d558, 32'hc1a8abaf} /* (12, 26, 10) {real, imag} */,
  {32'hc17aca42, 32'h414e4614} /* (12, 26, 9) {real, imag} */,
  {32'h42186740, 32'h416ef5fc} /* (12, 26, 8) {real, imag} */,
  {32'h41474256, 32'hc14e1a5d} /* (12, 26, 7) {real, imag} */,
  {32'hc28b7e81, 32'hc1628d0e} /* (12, 26, 6) {real, imag} */,
  {32'h4233d40c, 32'hc14ad727} /* (12, 26, 5) {real, imag} */,
  {32'h41f494a5, 32'hc1184e48} /* (12, 26, 4) {real, imag} */,
  {32'h41b635bc, 32'h424d3070} /* (12, 26, 3) {real, imag} */,
  {32'hc2a2441a, 32'h41c45bfc} /* (12, 26, 2) {real, imag} */,
  {32'hc1e564ba, 32'hc1388bc6} /* (12, 26, 1) {real, imag} */,
  {32'hc106854b, 32'h40cb1c98} /* (12, 26, 0) {real, imag} */,
  {32'h41ca2416, 32'h42082c49} /* (12, 25, 31) {real, imag} */,
  {32'h42477d48, 32'h41266738} /* (12, 25, 30) {real, imag} */,
  {32'hc0ed0a68, 32'h41704a0e} /* (12, 25, 29) {real, imag} */,
  {32'hc1a8c626, 32'h41998fc7} /* (12, 25, 28) {real, imag} */,
  {32'hc22a5d1e, 32'h41e7fb16} /* (12, 25, 27) {real, imag} */,
  {32'h42208469, 32'h41c85f5f} /* (12, 25, 26) {real, imag} */,
  {32'h4107836b, 32'h411087a3} /* (12, 25, 25) {real, imag} */,
  {32'hc1aed59c, 32'hc23b12b8} /* (12, 25, 24) {real, imag} */,
  {32'h41d6d79e, 32'hc172a30c} /* (12, 25, 23) {real, imag} */,
  {32'hc18bf606, 32'hc19f608e} /* (12, 25, 22) {real, imag} */,
  {32'h40497fbc, 32'hc09b75b6} /* (12, 25, 21) {real, imag} */,
  {32'hc11af35e, 32'h40a526b7} /* (12, 25, 20) {real, imag} */,
  {32'hbfe9ed18, 32'hc1846bdc} /* (12, 25, 19) {real, imag} */,
  {32'h416aa681, 32'hc0beb8e3} /* (12, 25, 18) {real, imag} */,
  {32'hc0d06829, 32'hc0fbf758} /* (12, 25, 17) {real, imag} */,
  {32'hc16b9cd4, 32'hbf3ef690} /* (12, 25, 16) {real, imag} */,
  {32'hc1022b5c, 32'h401d1730} /* (12, 25, 15) {real, imag} */,
  {32'h415491ed, 32'hbfb5aeb4} /* (12, 25, 14) {real, imag} */,
  {32'hc00df9a4, 32'h3fa59460} /* (12, 25, 13) {real, imag} */,
  {32'h40579294, 32'h408c468d} /* (12, 25, 12) {real, imag} */,
  {32'h400385ec, 32'hc14d2a21} /* (12, 25, 11) {real, imag} */,
  {32'h417c08cc, 32'hc192367a} /* (12, 25, 10) {real, imag} */,
  {32'hc196adbe, 32'hc1250b5a} /* (12, 25, 9) {real, imag} */,
  {32'h40d72718, 32'hc11563c2} /* (12, 25, 8) {real, imag} */,
  {32'h4171add5, 32'hc1c20f62} /* (12, 25, 7) {real, imag} */,
  {32'h41e08ce6, 32'h42647b68} /* (12, 25, 6) {real, imag} */,
  {32'h3f9075b0, 32'hc188f546} /* (12, 25, 5) {real, imag} */,
  {32'hc08888c8, 32'h41ae0ffd} /* (12, 25, 4) {real, imag} */,
  {32'hc2165862, 32'hc28c71ce} /* (12, 25, 3) {real, imag} */,
  {32'hc1471d4c, 32'h40a237b9} /* (12, 25, 2) {real, imag} */,
  {32'h412bab34, 32'hc26ae9f5} /* (12, 25, 1) {real, imag} */,
  {32'hc205301e, 32'h41e2fc64} /* (12, 25, 0) {real, imag} */,
  {32'h412df679, 32'hc18fb370} /* (12, 24, 31) {real, imag} */,
  {32'hc19b58fe, 32'h4155917d} /* (12, 24, 30) {real, imag} */,
  {32'h41963555, 32'h428e8f79} /* (12, 24, 29) {real, imag} */,
  {32'hc2030678, 32'h41cdd7c0} /* (12, 24, 28) {real, imag} */,
  {32'hc12f9b23, 32'hc25fb01f} /* (12, 24, 27) {real, imag} */,
  {32'h4153dcc0, 32'h4250d282} /* (12, 24, 26) {real, imag} */,
  {32'hc2237882, 32'hbfe803a0} /* (12, 24, 25) {real, imag} */,
  {32'hbd217d80, 32'h41e02992} /* (12, 24, 24) {real, imag} */,
  {32'hbe5c9860, 32'h414e5394} /* (12, 24, 23) {real, imag} */,
  {32'hc216c919, 32'h41ef0839} /* (12, 24, 22) {real, imag} */,
  {32'hc09b6590, 32'hc15eb99a} /* (12, 24, 21) {real, imag} */,
  {32'h41a7fcef, 32'h41cb9bd0} /* (12, 24, 20) {real, imag} */,
  {32'h41d2889f, 32'h404001e0} /* (12, 24, 19) {real, imag} */,
  {32'hc145a982, 32'hc14673f6} /* (12, 24, 18) {real, imag} */,
  {32'h404707ed, 32'h40786f9f} /* (12, 24, 17) {real, imag} */,
  {32'h407d2040, 32'hc07063f2} /* (12, 24, 16) {real, imag} */,
  {32'hc023b3df, 32'hc00505e9} /* (12, 24, 15) {real, imag} */,
  {32'h3f850500, 32'h41031b30} /* (12, 24, 14) {real, imag} */,
  {32'h4021ad68, 32'h3fd2f860} /* (12, 24, 13) {real, imag} */,
  {32'h3fb58fb0, 32'h40eb77a2} /* (12, 24, 12) {real, imag} */,
  {32'h40b98470, 32'hc1a0ba5f} /* (12, 24, 11) {real, imag} */,
  {32'h40787c00, 32'h41bd8e1f} /* (12, 24, 10) {real, imag} */,
  {32'h414f847a, 32'hc162c1da} /* (12, 24, 9) {real, imag} */,
  {32'hc0beeda5, 32'h42174867} /* (12, 24, 8) {real, imag} */,
  {32'hc13de882, 32'hc15235f2} /* (12, 24, 7) {real, imag} */,
  {32'h3fa84684, 32'hc0a3ca4c} /* (12, 24, 6) {real, imag} */,
  {32'h41100e63, 32'h413a8824} /* (12, 24, 5) {real, imag} */,
  {32'h41bf5e48, 32'h4143bc3f} /* (12, 24, 4) {real, imag} */,
  {32'hc228f174, 32'hc0a07a30} /* (12, 24, 3) {real, imag} */,
  {32'hc1c6da12, 32'h41e5819a} /* (12, 24, 2) {real, imag} */,
  {32'hc19f9f86, 32'h402e17d4} /* (12, 24, 1) {real, imag} */,
  {32'h4286ab94, 32'h403ae1a2} /* (12, 24, 0) {real, imag} */,
  {32'hc112abd2, 32'hc28072bb} /* (12, 23, 31) {real, imag} */,
  {32'hc1759f0f, 32'hbf965e54} /* (12, 23, 30) {real, imag} */,
  {32'h419d46c6, 32'h41d3f7b6} /* (12, 23, 29) {real, imag} */,
  {32'hc1ff466a, 32'hc192e2c5} /* (12, 23, 28) {real, imag} */,
  {32'h424afb41, 32'hc1a0d256} /* (12, 23, 27) {real, imag} */,
  {32'h4046e90a, 32'h42129732} /* (12, 23, 26) {real, imag} */,
  {32'h40d3b699, 32'h40f64a0c} /* (12, 23, 25) {real, imag} */,
  {32'hc192249e, 32'hc16ca85e} /* (12, 23, 24) {real, imag} */,
  {32'hc16b1e28, 32'hc123a358} /* (12, 23, 23) {real, imag} */,
  {32'hc0ea70dd, 32'hc135d9a6} /* (12, 23, 22) {real, imag} */,
  {32'h415a4c7f, 32'hc0de600a} /* (12, 23, 21) {real, imag} */,
  {32'h419dc3e0, 32'hc10c7a29} /* (12, 23, 20) {real, imag} */,
  {32'hc00d84bc, 32'h419d6f50} /* (12, 23, 19) {real, imag} */,
  {32'h409d1012, 32'hc156fb52} /* (12, 23, 18) {real, imag} */,
  {32'hc00f4cb6, 32'hc0c61e9c} /* (12, 23, 17) {real, imag} */,
  {32'h3f87cc40, 32'h40dbae64} /* (12, 23, 16) {real, imag} */,
  {32'hc03119fa, 32'hbfbc53b0} /* (12, 23, 15) {real, imag} */,
  {32'h40333d8d, 32'hc103549e} /* (12, 23, 14) {real, imag} */,
  {32'h415e2e03, 32'h413000d6} /* (12, 23, 13) {real, imag} */,
  {32'hc088bf00, 32'hc1adc85e} /* (12, 23, 12) {real, imag} */,
  {32'hc0832316, 32'hc0cf9aba} /* (12, 23, 11) {real, imag} */,
  {32'h403ded6a, 32'h3dabebc0} /* (12, 23, 10) {real, imag} */,
  {32'h40b08460, 32'hc101f6f4} /* (12, 23, 9) {real, imag} */,
  {32'hbfc07dc0, 32'h40a32db9} /* (12, 23, 8) {real, imag} */,
  {32'h416d0f0c, 32'hc0e18b46} /* (12, 23, 7) {real, imag} */,
  {32'hc0e1f5c9, 32'h41d33324} /* (12, 23, 6) {real, imag} */,
  {32'hbf6df7c0, 32'h42036df9} /* (12, 23, 5) {real, imag} */,
  {32'hc15350e8, 32'h4203f8e5} /* (12, 23, 4) {real, imag} */,
  {32'hc0664f34, 32'h409cc624} /* (12, 23, 3) {real, imag} */,
  {32'h41caec94, 32'hc16aa152} /* (12, 23, 2) {real, imag} */,
  {32'hc1fc0fa5, 32'h4129791e} /* (12, 23, 1) {real, imag} */,
  {32'hc20314a6, 32'h42026f76} /* (12, 23, 0) {real, imag} */,
  {32'hc218aa08, 32'h3fc5b5e0} /* (12, 22, 31) {real, imag} */,
  {32'h4207b5e7, 32'hbe9185ec} /* (12, 22, 30) {real, imag} */,
  {32'hc28b8791, 32'hc10a4d59} /* (12, 22, 29) {real, imag} */,
  {32'h41a1d108, 32'hc1763a06} /* (12, 22, 28) {real, imag} */,
  {32'h4122295c, 32'hc21fe7e5} /* (12, 22, 27) {real, imag} */,
  {32'hbff4a1d8, 32'h41356360} /* (12, 22, 26) {real, imag} */,
  {32'h41a373bf, 32'h41adc391} /* (12, 22, 25) {real, imag} */,
  {32'h415d7b9f, 32'hc12c87f4} /* (12, 22, 24) {real, imag} */,
  {32'hbd8c4640, 32'hc0838368} /* (12, 22, 23) {real, imag} */,
  {32'h4180a38b, 32'h41b62534} /* (12, 22, 22) {real, imag} */,
  {32'h412818f9, 32'hbe9021c0} /* (12, 22, 21) {real, imag} */,
  {32'h4019ef40, 32'h40257d74} /* (12, 22, 20) {real, imag} */,
  {32'hbfcbb170, 32'hc027c3d0} /* (12, 22, 19) {real, imag} */,
  {32'hc0fb242e, 32'h40550cbd} /* (12, 22, 18) {real, imag} */,
  {32'hc00eae98, 32'hbf0e5690} /* (12, 22, 17) {real, imag} */,
  {32'h40ef283c, 32'h415b0e8d} /* (12, 22, 16) {real, imag} */,
  {32'h4097a9c8, 32'hc0e86be2} /* (12, 22, 15) {real, imag} */,
  {32'h3f3941b0, 32'h4085b82a} /* (12, 22, 14) {real, imag} */,
  {32'hc0491438, 32'h3fe03688} /* (12, 22, 13) {real, imag} */,
  {32'hc13f07ba, 32'hc0866c2e} /* (12, 22, 12) {real, imag} */,
  {32'hc0fcaede, 32'h413e21e2} /* (12, 22, 11) {real, imag} */,
  {32'hc11a7bf8, 32'h408c8902} /* (12, 22, 10) {real, imag} */,
  {32'h40b34be7, 32'h3f583920} /* (12, 22, 9) {real, imag} */,
  {32'hc18d17e8, 32'hc0479a2e} /* (12, 22, 8) {real, imag} */,
  {32'hc1229a96, 32'hc1441cc6} /* (12, 22, 7) {real, imag} */,
  {32'h418b7986, 32'hc210d66c} /* (12, 22, 6) {real, imag} */,
  {32'h41a6f207, 32'h40d1f550} /* (12, 22, 5) {real, imag} */,
  {32'hbfe1f5d0, 32'hc1aab24d} /* (12, 22, 4) {real, imag} */,
  {32'h42249596, 32'hc188a290} /* (12, 22, 3) {real, imag} */,
  {32'h4218aa19, 32'h4021c590} /* (12, 22, 2) {real, imag} */,
  {32'hc09affa0, 32'h4238a1bf} /* (12, 22, 1) {real, imag} */,
  {32'hc02ab4e3, 32'h4213de51} /* (12, 22, 0) {real, imag} */,
  {32'h40eeddfe, 32'h41800077} /* (12, 21, 31) {real, imag} */,
  {32'h4175d8f6, 32'hc0bbbdcc} /* (12, 21, 30) {real, imag} */,
  {32'hc166e368, 32'hc18b82d8} /* (12, 21, 29) {real, imag} */,
  {32'h419f4193, 32'hc0c1bdd6} /* (12, 21, 28) {real, imag} */,
  {32'hc1c188d3, 32'h414bbb88} /* (12, 21, 27) {real, imag} */,
  {32'hbf9c4878, 32'hc0a3031a} /* (12, 21, 26) {real, imag} */,
  {32'hc1c1452a, 32'hc0d662f4} /* (12, 21, 25) {real, imag} */,
  {32'h4181ff48, 32'h412c6ca9} /* (12, 21, 24) {real, imag} */,
  {32'h4186d9ca, 32'h416a7714} /* (12, 21, 23) {real, imag} */,
  {32'hbf1076f0, 32'h41195dcc} /* (12, 21, 22) {real, imag} */,
  {32'h4121dde0, 32'h418ac722} /* (12, 21, 21) {real, imag} */,
  {32'hc12d0314, 32'hc11c2962} /* (12, 21, 20) {real, imag} */,
  {32'hc1237dfa, 32'hc12fc60f} /* (12, 21, 19) {real, imag} */,
  {32'h3f27b822, 32'hc0d130df} /* (12, 21, 18) {real, imag} */,
  {32'hc098c970, 32'hbe35a510} /* (12, 21, 17) {real, imag} */,
  {32'h3e2dd810, 32'hbff6a310} /* (12, 21, 16) {real, imag} */,
  {32'h3fdf7880, 32'h402fc419} /* (12, 21, 15) {real, imag} */,
  {32'hbea7a4c4, 32'h40613ec2} /* (12, 21, 14) {real, imag} */,
  {32'h40b5ae55, 32'h403b1368} /* (12, 21, 13) {real, imag} */,
  {32'h40c49534, 32'hc0c61bc7} /* (12, 21, 12) {real, imag} */,
  {32'hc0f7a767, 32'hc04b1168} /* (12, 21, 11) {real, imag} */,
  {32'hc18193a6, 32'h41a7e9c3} /* (12, 21, 10) {real, imag} */,
  {32'h40e28fba, 32'hc129fad4} /* (12, 21, 9) {real, imag} */,
  {32'hc150f038, 32'h4057663b} /* (12, 21, 8) {real, imag} */,
  {32'h41cb0b52, 32'hc16c28ae} /* (12, 21, 7) {real, imag} */,
  {32'hc1aea442, 32'h415d025f} /* (12, 21, 6) {real, imag} */,
  {32'h41e363a3, 32'hc1548f22} /* (12, 21, 5) {real, imag} */,
  {32'h412fb044, 32'hc213ccb1} /* (12, 21, 4) {real, imag} */,
  {32'hbe829310, 32'h41b1e1bc} /* (12, 21, 3) {real, imag} */,
  {32'h419fcb69, 32'hc1de5477} /* (12, 21, 2) {real, imag} */,
  {32'h4182702e, 32'h419aab81} /* (12, 21, 1) {real, imag} */,
  {32'h40b43ba4, 32'hc0e0c874} /* (12, 21, 0) {real, imag} */,
  {32'h4181a10e, 32'hc1632c59} /* (12, 20, 31) {real, imag} */,
  {32'hc0c898e4, 32'hc2411f46} /* (12, 20, 30) {real, imag} */,
  {32'h4181fe97, 32'hc1a9807c} /* (12, 20, 29) {real, imag} */,
  {32'hc181ec95, 32'h3f9f3438} /* (12, 20, 28) {real, imag} */,
  {32'h4164b39e, 32'h40ac9d94} /* (12, 20, 27) {real, imag} */,
  {32'h414a230a, 32'hc0430740} /* (12, 20, 26) {real, imag} */,
  {32'hc036d9cc, 32'hc136cc04} /* (12, 20, 25) {real, imag} */,
  {32'hc1cb1bd0, 32'h3f73c288} /* (12, 20, 24) {real, imag} */,
  {32'h410b20be, 32'h40afd5bf} /* (12, 20, 23) {real, imag} */,
  {32'h3f839d9e, 32'hbfea79e0} /* (12, 20, 22) {real, imag} */,
  {32'hc141b562, 32'h40b33d39} /* (12, 20, 21) {real, imag} */,
  {32'h41308152, 32'h408c9e36} /* (12, 20, 20) {real, imag} */,
  {32'h40a8f5ca, 32'h403c982e} /* (12, 20, 19) {real, imag} */,
  {32'hc09fa490, 32'h409ec4d8} /* (12, 20, 18) {real, imag} */,
  {32'h406f5956, 32'h40b1adaf} /* (12, 20, 17) {real, imag} */,
  {32'hc00a4e8a, 32'h3f873248} /* (12, 20, 16) {real, imag} */,
  {32'hc0607b8e, 32'hbfef1afc} /* (12, 20, 15) {real, imag} */,
  {32'h3e812e28, 32'h409334a8} /* (12, 20, 14) {real, imag} */,
  {32'h40c0c23e, 32'h3fc9b8ac} /* (12, 20, 13) {real, imag} */,
  {32'h4017a438, 32'h418747ac} /* (12, 20, 12) {real, imag} */,
  {32'h4123613a, 32'h3ec55ae0} /* (12, 20, 11) {real, imag} */,
  {32'hc0dee22c, 32'hc1fce9de} /* (12, 20, 10) {real, imag} */,
  {32'hc16bc602, 32'hbff5bd94} /* (12, 20, 9) {real, imag} */,
  {32'hc0e44b30, 32'hc185ee32} /* (12, 20, 8) {real, imag} */,
  {32'h4112cf0e, 32'h41bbdcd6} /* (12, 20, 7) {real, imag} */,
  {32'hc0cab6e4, 32'h3fe90800} /* (12, 20, 6) {real, imag} */,
  {32'hc2345176, 32'h3fbc6354} /* (12, 20, 5) {real, imag} */,
  {32'h41400862, 32'h41e2dd6e} /* (12, 20, 4) {real, imag} */,
  {32'h41884cb3, 32'h41144614} /* (12, 20, 3) {real, imag} */,
  {32'h40881d74, 32'h4053d560} /* (12, 20, 2) {real, imag} */,
  {32'h41a2e12e, 32'hc12f0b79} /* (12, 20, 1) {real, imag} */,
  {32'hbfcaaf8c, 32'h4116774c} /* (12, 20, 0) {real, imag} */,
  {32'h40b4d36c, 32'hc09ad268} /* (12, 19, 31) {real, imag} */,
  {32'hc039f7a0, 32'h41b2e285} /* (12, 19, 30) {real, imag} */,
  {32'h41654690, 32'hc18d261e} /* (12, 19, 29) {real, imag} */,
  {32'h417b3f82, 32'h41c6258e} /* (12, 19, 28) {real, imag} */,
  {32'h3ebb2f30, 32'h41ecd3f4} /* (12, 19, 27) {real, imag} */,
  {32'h4103fe2c, 32'hc1fd1f16} /* (12, 19, 26) {real, imag} */,
  {32'hc08e2fb1, 32'hc12a766c} /* (12, 19, 25) {real, imag} */,
  {32'hc0607e0e, 32'hbdde2780} /* (12, 19, 24) {real, imag} */,
  {32'hc16fa3ca, 32'h3e3efaa0} /* (12, 19, 23) {real, imag} */,
  {32'h41a9986a, 32'hc1737b6d} /* (12, 19, 22) {real, imag} */,
  {32'h3f3b9a34, 32'h40e0bbf2} /* (12, 19, 21) {real, imag} */,
  {32'h3ff7d380, 32'hc07d05ac} /* (12, 19, 20) {real, imag} */,
  {32'h3df06500, 32'h40d62e97} /* (12, 19, 19) {real, imag} */,
  {32'h401eb748, 32'h3ff4e0a2} /* (12, 19, 18) {real, imag} */,
  {32'h408b8e5d, 32'hbf21270c} /* (12, 19, 17) {real, imag} */,
  {32'hc013582e, 32'hbf9e57c8} /* (12, 19, 16) {real, imag} */,
  {32'hc06d628e, 32'hbf98831e} /* (12, 19, 15) {real, imag} */,
  {32'h4000146c, 32'h4055d09f} /* (12, 19, 14) {real, imag} */,
  {32'h40873378, 32'hbea42f30} /* (12, 19, 13) {real, imag} */,
  {32'h411f5390, 32'h405e9ad4} /* (12, 19, 12) {real, imag} */,
  {32'hc0ba4cd2, 32'hc00fe32c} /* (12, 19, 11) {real, imag} */,
  {32'hbe8b1080, 32'h3fdc9128} /* (12, 19, 10) {real, imag} */,
  {32'hc0af24d4, 32'h3f617b40} /* (12, 19, 9) {real, imag} */,
  {32'hc1601d0a, 32'h419599ca} /* (12, 19, 8) {real, imag} */,
  {32'hc0161cd2, 32'hc0114780} /* (12, 19, 7) {real, imag} */,
  {32'hc178f4b4, 32'hc1a8fd5e} /* (12, 19, 6) {real, imag} */,
  {32'hc107de0c, 32'hc1431999} /* (12, 19, 5) {real, imag} */,
  {32'h4087f13c, 32'hc0494bfc} /* (12, 19, 4) {real, imag} */,
  {32'hbea13640, 32'hc18f51d2} /* (12, 19, 3) {real, imag} */,
  {32'h41c3da38, 32'h417687bb} /* (12, 19, 2) {real, imag} */,
  {32'h41591e36, 32'h419f5314} /* (12, 19, 1) {real, imag} */,
  {32'hbfa227f4, 32'hc1deb92a} /* (12, 19, 0) {real, imag} */,
  {32'h40bdb12e, 32'h41096808} /* (12, 18, 31) {real, imag} */,
  {32'hc1486bd4, 32'hbdb75180} /* (12, 18, 30) {real, imag} */,
  {32'h41cf95c4, 32'hc119a6de} /* (12, 18, 29) {real, imag} */,
  {32'h4101f86a, 32'hc10dc740} /* (12, 18, 28) {real, imag} */,
  {32'hc0beabd0, 32'h414859d4} /* (12, 18, 27) {real, imag} */,
  {32'h3ebd1638, 32'h4000e68c} /* (12, 18, 26) {real, imag} */,
  {32'h40afdcca, 32'hc00874b0} /* (12, 18, 25) {real, imag} */,
  {32'hbf8638ba, 32'hc02814aa} /* (12, 18, 24) {real, imag} */,
  {32'h40312828, 32'h412b0986} /* (12, 18, 23) {real, imag} */,
  {32'hc155f348, 32'hc1209e1c} /* (12, 18, 22) {real, imag} */,
  {32'h40ca028e, 32'h40ca765a} /* (12, 18, 21) {real, imag} */,
  {32'hc0a3e476, 32'hbf4d465e} /* (12, 18, 20) {real, imag} */,
  {32'h3fbcd8ba, 32'h409f0874} /* (12, 18, 19) {real, imag} */,
  {32'hc0693ed0, 32'hc1155c32} /* (12, 18, 18) {real, imag} */,
  {32'hbe948658, 32'hc0369d58} /* (12, 18, 17) {real, imag} */,
  {32'hc0b92418, 32'hbf8da028} /* (12, 18, 16) {real, imag} */,
  {32'hc0d4d876, 32'hc00278ec} /* (12, 18, 15) {real, imag} */,
  {32'hbfe9e250, 32'hc118555c} /* (12, 18, 14) {real, imag} */,
  {32'h40cb8df6, 32'h40e9d0f0} /* (12, 18, 13) {real, imag} */,
  {32'hc105c04b, 32'h3faebf67} /* (12, 18, 12) {real, imag} */,
  {32'hc0f0fc12, 32'hc0a81298} /* (12, 18, 11) {real, imag} */,
  {32'h4135e014, 32'h415174e6} /* (12, 18, 10) {real, imag} */,
  {32'h41780dc0, 32'hc05f7101} /* (12, 18, 9) {real, imag} */,
  {32'hc03ef36d, 32'hc0d0be37} /* (12, 18, 8) {real, imag} */,
  {32'h40e76672, 32'h406dea72} /* (12, 18, 7) {real, imag} */,
  {32'hc0379509, 32'hc1c7083a} /* (12, 18, 6) {real, imag} */,
  {32'h40f81fac, 32'h41069888} /* (12, 18, 5) {real, imag} */,
  {32'h3f666bc4, 32'hc1668f84} /* (12, 18, 4) {real, imag} */,
  {32'hc0f58e42, 32'h40b21a10} /* (12, 18, 3) {real, imag} */,
  {32'hc103b7fe, 32'h41cfad36} /* (12, 18, 2) {real, imag} */,
  {32'h41974a42, 32'hbfb2c6f4} /* (12, 18, 1) {real, imag} */,
  {32'h4125a86c, 32'h418b173e} /* (12, 18, 0) {real, imag} */,
  {32'hbf7a1cf0, 32'hc043f46c} /* (12, 17, 31) {real, imag} */,
  {32'h41a2273c, 32'hc09c090b} /* (12, 17, 30) {real, imag} */,
  {32'hc11cc9e7, 32'hbfada294} /* (12, 17, 29) {real, imag} */,
  {32'h413b0ba4, 32'h41b7cdbb} /* (12, 17, 28) {real, imag} */,
  {32'h40851e0f, 32'h408eab44} /* (12, 17, 27) {real, imag} */,
  {32'h3f909230, 32'h41ad1704} /* (12, 17, 26) {real, imag} */,
  {32'hc11a6580, 32'hc1509138} /* (12, 17, 25) {real, imag} */,
  {32'hc0353934, 32'h40560e1a} /* (12, 17, 24) {real, imag} */,
  {32'hc15dacec, 32'hc1192bcd} /* (12, 17, 23) {real, imag} */,
  {32'h410cbb1a, 32'h41209896} /* (12, 17, 22) {real, imag} */,
  {32'h401f7d72, 32'hc067c192} /* (12, 17, 21) {real, imag} */,
  {32'h405bc753, 32'h4033c78e} /* (12, 17, 20) {real, imag} */,
  {32'h401ae5fe, 32'h3f7fb7f2} /* (12, 17, 19) {real, imag} */,
  {32'hbf8cc5a6, 32'h3fb5508c} /* (12, 17, 18) {real, imag} */,
  {32'hbea94280, 32'hbf3cbe30} /* (12, 17, 17) {real, imag} */,
  {32'hbebe0630, 32'h3e2924c0} /* (12, 17, 16) {real, imag} */,
  {32'h4047b71d, 32'hbfed0f38} /* (12, 17, 15) {real, imag} */,
  {32'h40c941ba, 32'h402f32c2} /* (12, 17, 14) {real, imag} */,
  {32'hc00c12c6, 32'h40430bb8} /* (12, 17, 13) {real, imag} */,
  {32'hbf03e524, 32'h400a23e2} /* (12, 17, 12) {real, imag} */,
  {32'hc0045712, 32'h4003d67e} /* (12, 17, 11) {real, imag} */,
  {32'hc06bfdb2, 32'h403a4d26} /* (12, 17, 10) {real, imag} */,
  {32'hc0a83079, 32'h4122e65b} /* (12, 17, 9) {real, imag} */,
  {32'h3dc50a80, 32'hc18a3661} /* (12, 17, 8) {real, imag} */,
  {32'h415a8524, 32'hc04fbefe} /* (12, 17, 7) {real, imag} */,
  {32'h41fe9ef9, 32'hc0d92ba7} /* (12, 17, 6) {real, imag} */,
  {32'hc1223afa, 32'h417d8036} /* (12, 17, 5) {real, imag} */,
  {32'hc0524536, 32'h3dd1df00} /* (12, 17, 4) {real, imag} */,
  {32'h4116ebfd, 32'hc1015206} /* (12, 17, 3) {real, imag} */,
  {32'h409cdcfe, 32'h409b00c5} /* (12, 17, 2) {real, imag} */,
  {32'hc0c078f0, 32'hc1dab440} /* (12, 17, 1) {real, imag} */,
  {32'hc0328d56, 32'hc182c33c} /* (12, 17, 0) {real, imag} */,
  {32'h40d41f96, 32'hc173378c} /* (12, 16, 31) {real, imag} */,
  {32'h41918076, 32'h41b1e0c8} /* (12, 16, 30) {real, imag} */,
  {32'hc12049ff, 32'h413ab6b4} /* (12, 16, 29) {real, imag} */,
  {32'hc18d5939, 32'hc0e0fcbe} /* (12, 16, 28) {real, imag} */,
  {32'h3fbfabae, 32'h418315a3} /* (12, 16, 27) {real, imag} */,
  {32'hc0840686, 32'hc0de0f44} /* (12, 16, 26) {real, imag} */,
  {32'h4054a818, 32'h40b24df2} /* (12, 16, 25) {real, imag} */,
  {32'hc11c97b7, 32'hc0ace780} /* (12, 16, 24) {real, imag} */,
  {32'h4096c746, 32'h3fdf010a} /* (12, 16, 23) {real, imag} */,
  {32'hbf4a9f18, 32'hc0ab3862} /* (12, 16, 22) {real, imag} */,
  {32'h410d164e, 32'hc03717f0} /* (12, 16, 21) {real, imag} */,
  {32'h40f91ba7, 32'hbe5c7178} /* (12, 16, 20) {real, imag} */,
  {32'hc0e90788, 32'h40c34cab} /* (12, 16, 19) {real, imag} */,
  {32'h3fe743c6, 32'hbfe0cdf0} /* (12, 16, 18) {real, imag} */,
  {32'h40089025, 32'h407d4e58} /* (12, 16, 17) {real, imag} */,
  {32'hc053f5fb, 32'h3edfb3dc} /* (12, 16, 16) {real, imag} */,
  {32'hc070e13f, 32'h40914b38} /* (12, 16, 15) {real, imag} */,
  {32'hc059288d, 32'h3fcd9280} /* (12, 16, 14) {real, imag} */,
  {32'hc0d0f7d6, 32'h40a0b47f} /* (12, 16, 13) {real, imag} */,
  {32'hc0a72e31, 32'hbfdb3ccf} /* (12, 16, 12) {real, imag} */,
  {32'h3f1ce440, 32'h3d6e5120} /* (12, 16, 11) {real, imag} */,
  {32'hc07d8e1e, 32'h3fd07cda} /* (12, 16, 10) {real, imag} */,
  {32'h40df778a, 32'h410c40dd} /* (12, 16, 9) {real, imag} */,
  {32'hbf8cd5b8, 32'hc11e23a0} /* (12, 16, 8) {real, imag} */,
  {32'h400328c6, 32'hc12e6f63} /* (12, 16, 7) {real, imag} */,
  {32'hc17b1cc5, 32'hc121137c} /* (12, 16, 6) {real, imag} */,
  {32'h3dacb6e0, 32'h40e321ed} /* (12, 16, 5) {real, imag} */,
  {32'hbe74f780, 32'h411ef7f5} /* (12, 16, 4) {real, imag} */,
  {32'hc17cfb4d, 32'hc03af46a} /* (12, 16, 3) {real, imag} */,
  {32'hc02720cc, 32'h40e3aafc} /* (12, 16, 2) {real, imag} */,
  {32'h40cbe33a, 32'hbe9f1770} /* (12, 16, 1) {real, imag} */,
  {32'h40aceeae, 32'hbfee944b} /* (12, 16, 0) {real, imag} */,
  {32'h41174200, 32'hc0c9a78d} /* (12, 15, 31) {real, imag} */,
  {32'h40e800a4, 32'h41107f54} /* (12, 15, 30) {real, imag} */,
  {32'h41467e48, 32'hc034a0c0} /* (12, 15, 29) {real, imag} */,
  {32'h40e882ea, 32'h403218b6} /* (12, 15, 28) {real, imag} */,
  {32'hc0c3f34e, 32'h404747a0} /* (12, 15, 27) {real, imag} */,
  {32'hc08b48fa, 32'h41388211} /* (12, 15, 26) {real, imag} */,
  {32'hc09f7b93, 32'h40e3e544} /* (12, 15, 25) {real, imag} */,
  {32'h41439faa, 32'h409c41e8} /* (12, 15, 24) {real, imag} */,
  {32'h418ab7ae, 32'hbf5d3be8} /* (12, 15, 23) {real, imag} */,
  {32'h3ec66570, 32'hc0365d30} /* (12, 15, 22) {real, imag} */,
  {32'hc0adcbee, 32'h405c70d2} /* (12, 15, 21) {real, imag} */,
  {32'hc16c3e57, 32'h3f97752c} /* (12, 15, 20) {real, imag} */,
  {32'h3f73bbc0, 32'h3f3c8618} /* (12, 15, 19) {real, imag} */,
  {32'h40182d1b, 32'hbfec4f82} /* (12, 15, 18) {real, imag} */,
  {32'h40655b7a, 32'h40bb8752} /* (12, 15, 17) {real, imag} */,
  {32'hbee378f0, 32'h3fde9b48} /* (12, 15, 16) {real, imag} */,
  {32'hbf87583c, 32'hc023ec44} /* (12, 15, 15) {real, imag} */,
  {32'hbfa09466, 32'h3f42ccb4} /* (12, 15, 14) {real, imag} */,
  {32'h40bde2b6, 32'hc08798bd} /* (12, 15, 13) {real, imag} */,
  {32'h4015a60c, 32'hc123f276} /* (12, 15, 12) {real, imag} */,
  {32'h3fe6c938, 32'h40de610d} /* (12, 15, 11) {real, imag} */,
  {32'hc1129ab0, 32'hbf60f0c2} /* (12, 15, 10) {real, imag} */,
  {32'hbf3143b0, 32'h4023f2bc} /* (12, 15, 9) {real, imag} */,
  {32'h404705aa, 32'hc1485852} /* (12, 15, 8) {real, imag} */,
  {32'h3fdd8a9c, 32'h4105024e} /* (12, 15, 7) {real, imag} */,
  {32'h3ffcc148, 32'hc1a95370} /* (12, 15, 6) {real, imag} */,
  {32'hc0e9bf5a, 32'h41324799} /* (12, 15, 5) {real, imag} */,
  {32'hc17722c9, 32'hc18c301a} /* (12, 15, 4) {real, imag} */,
  {32'hc0d0c5f8, 32'h3f0aa09e} /* (12, 15, 3) {real, imag} */,
  {32'h3f8032be, 32'h4026d445} /* (12, 15, 2) {real, imag} */,
  {32'h4026438c, 32'h40f5a4bb} /* (12, 15, 1) {real, imag} */,
  {32'h4183044d, 32'h3eb41620} /* (12, 15, 0) {real, imag} */,
  {32'hc16be35a, 32'hc11c3f66} /* (12, 14, 31) {real, imag} */,
  {32'hc15892da, 32'h4159f916} /* (12, 14, 30) {real, imag} */,
  {32'h4029d2ae, 32'h40164385} /* (12, 14, 29) {real, imag} */,
  {32'h41caed7a, 32'hbede9060} /* (12, 14, 28) {real, imag} */,
  {32'h3f2dec10, 32'hc16b322a} /* (12, 14, 27) {real, imag} */,
  {32'hc1a17106, 32'h4100ceaa} /* (12, 14, 26) {real, imag} */,
  {32'hc0f0bd42, 32'h400b244b} /* (12, 14, 25) {real, imag} */,
  {32'hbf76663e, 32'h40813107} /* (12, 14, 24) {real, imag} */,
  {32'hc12cded6, 32'h408d6b78} /* (12, 14, 23) {real, imag} */,
  {32'hc1773355, 32'h3f0e94a8} /* (12, 14, 22) {real, imag} */,
  {32'h412f589e, 32'hc0c0d286} /* (12, 14, 21) {real, imag} */,
  {32'h40e57e86, 32'hc035d5b8} /* (12, 14, 20) {real, imag} */,
  {32'h40b37bd5, 32'hc09af46a} /* (12, 14, 19) {real, imag} */,
  {32'h3f1095e8, 32'h3eca6ce0} /* (12, 14, 18) {real, imag} */,
  {32'hbfbb31cc, 32'h3fe79b9e} /* (12, 14, 17) {real, imag} */,
  {32'hbfa05722, 32'hc0a02f22} /* (12, 14, 16) {real, imag} */,
  {32'h411aa41a, 32'hc0cd39f2} /* (12, 14, 15) {real, imag} */,
  {32'h406e5c62, 32'hc10318f3} /* (12, 14, 14) {real, imag} */,
  {32'h408cf067, 32'h408e428e} /* (12, 14, 13) {real, imag} */,
  {32'h3f272dac, 32'h404ed4d8} /* (12, 14, 12) {real, imag} */,
  {32'h40950514, 32'h4074ef44} /* (12, 14, 11) {real, imag} */,
  {32'hc0760eec, 32'h4088740b} /* (12, 14, 10) {real, imag} */,
  {32'hc13df208, 32'h40cea4a6} /* (12, 14, 9) {real, imag} */,
  {32'h40910df6, 32'h3f2485f6} /* (12, 14, 8) {real, imag} */,
  {32'hc1c277dc, 32'hbf2b3f3c} /* (12, 14, 7) {real, imag} */,
  {32'hc0e489ce, 32'hc15bc78a} /* (12, 14, 6) {real, imag} */,
  {32'hc10ce8dd, 32'hc2094244} /* (12, 14, 5) {real, imag} */,
  {32'hc19f6fd0, 32'h416a7e5f} /* (12, 14, 4) {real, imag} */,
  {32'hc14a23aa, 32'hbf3bbedc} /* (12, 14, 3) {real, imag} */,
  {32'h4140ed78, 32'hc10ed85c} /* (12, 14, 2) {real, imag} */,
  {32'h406bc838, 32'hc021daf8} /* (12, 14, 1) {real, imag} */,
  {32'hc01e86bc, 32'h412751c8} /* (12, 14, 0) {real, imag} */,
  {32'hc1d5343d, 32'hc0cd8f66} /* (12, 13, 31) {real, imag} */,
  {32'h4181ce87, 32'h40fc9437} /* (12, 13, 30) {real, imag} */,
  {32'hc1db71f4, 32'h41e05ec7} /* (12, 13, 29) {real, imag} */,
  {32'hc0d1dc3e, 32'hbfb36e00} /* (12, 13, 28) {real, imag} */,
  {32'hc195b5d3, 32'h41b2fd36} /* (12, 13, 27) {real, imag} */,
  {32'hc10864e4, 32'h41b135ff} /* (12, 13, 26) {real, imag} */,
  {32'h3fcb2828, 32'h403f5e78} /* (12, 13, 25) {real, imag} */,
  {32'h410b329c, 32'h3ed43548} /* (12, 13, 24) {real, imag} */,
  {32'h40d3e8d5, 32'hc088deec} /* (12, 13, 23) {real, imag} */,
  {32'h3f6b3010, 32'h3fc294ec} /* (12, 13, 22) {real, imag} */,
  {32'h41502447, 32'h3f627518} /* (12, 13, 21) {real, imag} */,
  {32'hbf901140, 32'h41158dba} /* (12, 13, 20) {real, imag} */,
  {32'hc0936b26, 32'h40246dba} /* (12, 13, 19) {real, imag} */,
  {32'hc0c02a7a, 32'h40b78334} /* (12, 13, 18) {real, imag} */,
  {32'hc020f1a2, 32'hc04b6efc} /* (12, 13, 17) {real, imag} */,
  {32'hc0cec988, 32'h3fa7f470} /* (12, 13, 16) {real, imag} */,
  {32'hc02cfc66, 32'h4030a53c} /* (12, 13, 15) {real, imag} */,
  {32'hc015064c, 32'hbf5e8004} /* (12, 13, 14) {real, imag} */,
  {32'hbf22e850, 32'h3f7e1a08} /* (12, 13, 13) {real, imag} */,
  {32'hbf4786a8, 32'hc0a8ab70} /* (12, 13, 12) {real, imag} */,
  {32'h4110f1cd, 32'h40eb4d13} /* (12, 13, 11) {real, imag} */,
  {32'h40290712, 32'hc0dab8f5} /* (12, 13, 10) {real, imag} */,
  {32'h413f1640, 32'h3f4e4d66} /* (12, 13, 9) {real, imag} */,
  {32'h413f720c, 32'hbec05e78} /* (12, 13, 8) {real, imag} */,
  {32'h4110e149, 32'hc0cfda0c} /* (12, 13, 7) {real, imag} */,
  {32'h3ff6b72e, 32'h4016cf08} /* (12, 13, 6) {real, imag} */,
  {32'h4216a146, 32'hc09693a0} /* (12, 13, 5) {real, imag} */,
  {32'hc12d49a9, 32'hc1d45765} /* (12, 13, 4) {real, imag} */,
  {32'h402b13e4, 32'hc190bc7d} /* (12, 13, 3) {real, imag} */,
  {32'hc089be04, 32'hc0b0506d} /* (12, 13, 2) {real, imag} */,
  {32'hc139e6ee, 32'h41b1a902} /* (12, 13, 1) {real, imag} */,
  {32'h41b03ace, 32'h40022cee} /* (12, 13, 0) {real, imag} */,
  {32'hc1574306, 32'h41b80d84} /* (12, 12, 31) {real, imag} */,
  {32'h402bf773, 32'hc120fe22} /* (12, 12, 30) {real, imag} */,
  {32'h41aa0659, 32'h41aa9620} /* (12, 12, 29) {real, imag} */,
  {32'hc1a94045, 32'h40f8df4d} /* (12, 12, 28) {real, imag} */,
  {32'hc0ac0c2e, 32'hc1217b64} /* (12, 12, 27) {real, imag} */,
  {32'h408293a1, 32'hc155ae55} /* (12, 12, 26) {real, imag} */,
  {32'hc019458c, 32'hc1572e54} /* (12, 12, 25) {real, imag} */,
  {32'h40a0e3e0, 32'hc11b3b90} /* (12, 12, 24) {real, imag} */,
  {32'hc105f4aa, 32'hc117ca08} /* (12, 12, 23) {real, imag} */,
  {32'h40ce2f8b, 32'hc114e336} /* (12, 12, 22) {real, imag} */,
  {32'h3db311a0, 32'h3df0b8e0} /* (12, 12, 21) {real, imag} */,
  {32'h3f978280, 32'h40c43777} /* (12, 12, 20) {real, imag} */,
  {32'hc08cb60e, 32'hc0cbf284} /* (12, 12, 19) {real, imag} */,
  {32'hc0f403d4, 32'h3fd070f4} /* (12, 12, 18) {real, imag} */,
  {32'hc07f106c, 32'hbf0708f0} /* (12, 12, 17) {real, imag} */,
  {32'h40db0d64, 32'h404c3330} /* (12, 12, 16) {real, imag} */,
  {32'h405d53d8, 32'hc064679c} /* (12, 12, 15) {real, imag} */,
  {32'hc0b2b718, 32'hc0c10b81} /* (12, 12, 14) {real, imag} */,
  {32'hc0ec3612, 32'hbee831f8} /* (12, 12, 13) {real, imag} */,
  {32'hc14c25e3, 32'hc0a95589} /* (12, 12, 12) {real, imag} */,
  {32'hbec26fd8, 32'hc0f02378} /* (12, 12, 11) {real, imag} */,
  {32'hc126921a, 32'h417ff454} /* (12, 12, 10) {real, imag} */,
  {32'h41d65059, 32'hc17d7f44} /* (12, 12, 9) {real, imag} */,
  {32'hc0c0d11c, 32'h3fa798d4} /* (12, 12, 8) {real, imag} */,
  {32'hc0494dbc, 32'h406f3602} /* (12, 12, 7) {real, imag} */,
  {32'hc041c6ae, 32'hc1f87afe} /* (12, 12, 6) {real, imag} */,
  {32'h4194e234, 32'hc1355264} /* (12, 12, 5) {real, imag} */,
  {32'hc0dae6a5, 32'hc0378756} /* (12, 12, 4) {real, imag} */,
  {32'h41f80373, 32'h41c3d520} /* (12, 12, 3) {real, imag} */,
  {32'hc086239a, 32'hc196737e} /* (12, 12, 2) {real, imag} */,
  {32'hc0fb4bbb, 32'hc1216ef7} /* (12, 12, 1) {real, imag} */,
  {32'h41ea46bf, 32'h423afaa9} /* (12, 12, 0) {real, imag} */,
  {32'h40d49e78, 32'hc1d62fea} /* (12, 11, 31) {real, imag} */,
  {32'hc200b2a6, 32'hc168972d} /* (12, 11, 30) {real, imag} */,
  {32'h419b6768, 32'hc1334f3c} /* (12, 11, 29) {real, imag} */,
  {32'hc1a363e2, 32'h40b1bfe7} /* (12, 11, 28) {real, imag} */,
  {32'h40ad7d5c, 32'h4180b84e} /* (12, 11, 27) {real, imag} */,
  {32'h410ea860, 32'hbfcbccd0} /* (12, 11, 26) {real, imag} */,
  {32'h4204848b, 32'hc027242c} /* (12, 11, 25) {real, imag} */,
  {32'h40843304, 32'hc18b62ef} /* (12, 11, 24) {real, imag} */,
  {32'hc0cb4fec, 32'h40402e0c} /* (12, 11, 23) {real, imag} */,
  {32'h418574e5, 32'h40c4aa36} /* (12, 11, 22) {real, imag} */,
  {32'h4125a146, 32'hc12168a6} /* (12, 11, 21) {real, imag} */,
  {32'h416f2ac7, 32'h413837b0} /* (12, 11, 20) {real, imag} */,
  {32'hbf641d60, 32'h4143aaee} /* (12, 11, 19) {real, imag} */,
  {32'h40b2af60, 32'hbfbf6286} /* (12, 11, 18) {real, imag} */,
  {32'hbf211cc0, 32'hc04e9432} /* (12, 11, 17) {real, imag} */,
  {32'h3f735d58, 32'h409de0ea} /* (12, 11, 16) {real, imag} */,
  {32'hc03ce3c8, 32'hc0de5ed9} /* (12, 11, 15) {real, imag} */,
  {32'h40927680, 32'h40a3a236} /* (12, 11, 14) {real, imag} */,
  {32'hc0aca3a0, 32'hbf70f618} /* (12, 11, 13) {real, imag} */,
  {32'h412c88d3, 32'hc02626a2} /* (12, 11, 12) {real, imag} */,
  {32'h403b2d98, 32'h40aaffa7} /* (12, 11, 11) {real, imag} */,
  {32'hc17b726e, 32'hc07bc8f3} /* (12, 11, 10) {real, imag} */,
  {32'h41eaa445, 32'h41d280e2} /* (12, 11, 9) {real, imag} */,
  {32'h41913d31, 32'h41282234} /* (12, 11, 8) {real, imag} */,
  {32'hc1879d9a, 32'h415bfce9} /* (12, 11, 7) {real, imag} */,
  {32'hc204c18e, 32'h3f8f3c74} /* (12, 11, 6) {real, imag} */,
  {32'h409c1d24, 32'h413843f3} /* (12, 11, 5) {real, imag} */,
  {32'h3fc7bf28, 32'hc11f73ca} /* (12, 11, 4) {real, imag} */,
  {32'h420704c0, 32'h4193240c} /* (12, 11, 3) {real, imag} */,
  {32'h41e94bfb, 32'h4194b878} /* (12, 11, 2) {real, imag} */,
  {32'hc02a29b8, 32'hc10edc41} /* (12, 11, 1) {real, imag} */,
  {32'hc0d907a1, 32'hc20ba483} /* (12, 11, 0) {real, imag} */,
  {32'hc1e53ee2, 32'h40b135e4} /* (12, 10, 31) {real, imag} */,
  {32'hc0bfa26c, 32'h4137ba58} /* (12, 10, 30) {real, imag} */,
  {32'hc09c46b8, 32'hc17d4672} /* (12, 10, 29) {real, imag} */,
  {32'h40eb5c14, 32'hc0bd88bd} /* (12, 10, 28) {real, imag} */,
  {32'hc1018bcc, 32'h423517fb} /* (12, 10, 27) {real, imag} */,
  {32'hc1c497aa, 32'hc01b359a} /* (12, 10, 26) {real, imag} */,
  {32'h3fffde80, 32'hc10e9424} /* (12, 10, 25) {real, imag} */,
  {32'hc132e70e, 32'hc18e60f1} /* (12, 10, 24) {real, imag} */,
  {32'h3fe7ded0, 32'hc13b98ec} /* (12, 10, 23) {real, imag} */,
  {32'h40c3aa6c, 32'hbfbb240c} /* (12, 10, 22) {real, imag} */,
  {32'h410bf6e2, 32'h3f0a06a8} /* (12, 10, 21) {real, imag} */,
  {32'h404d9916, 32'hc08314ee} /* (12, 10, 20) {real, imag} */,
  {32'h41135e4d, 32'h40cb605e} /* (12, 10, 19) {real, imag} */,
  {32'hc11c0962, 32'hc0ca9830} /* (12, 10, 18) {real, imag} */,
  {32'hbfcd0480, 32'hbca2aa00} /* (12, 10, 17) {real, imag} */,
  {32'hc0ac262b, 32'h3f32db28} /* (12, 10, 16) {real, imag} */,
  {32'h413b1d7e, 32'h4140d8b9} /* (12, 10, 15) {real, imag} */,
  {32'h419ef5c4, 32'hc0aceb1a} /* (12, 10, 14) {real, imag} */,
  {32'hc0b55fba, 32'h3e4bbd00} /* (12, 10, 13) {real, imag} */,
  {32'hc13965c2, 32'h41765e49} /* (12, 10, 12) {real, imag} */,
  {32'hc060d666, 32'hbe759ea0} /* (12, 10, 11) {real, imag} */,
  {32'hc02ed7c0, 32'h407e39b6} /* (12, 10, 10) {real, imag} */,
  {32'hc18783db, 32'hbf98dd24} /* (12, 10, 9) {real, imag} */,
  {32'hc008d782, 32'hc1146cc4} /* (12, 10, 8) {real, imag} */,
  {32'hc1145f90, 32'hc145e860} /* (12, 10, 7) {real, imag} */,
  {32'hc22a6301, 32'hc10bf51a} /* (12, 10, 6) {real, imag} */,
  {32'hc18e7218, 32'h418b040e} /* (12, 10, 5) {real, imag} */,
  {32'h41f14393, 32'hc1166c9a} /* (12, 10, 4) {real, imag} */,
  {32'hc21a9c43, 32'hc16fa0f6} /* (12, 10, 3) {real, imag} */,
  {32'h41a5a12e, 32'h41528338} /* (12, 10, 2) {real, imag} */,
  {32'hc191a8ba, 32'hc20b2100} /* (12, 10, 1) {real, imag} */,
  {32'hc11d75f2, 32'hc10646a4} /* (12, 10, 0) {real, imag} */,
  {32'hc1b634fb, 32'h419457e4} /* (12, 9, 31) {real, imag} */,
  {32'h3ffb895e, 32'h428aa931} /* (12, 9, 30) {real, imag} */,
  {32'h41472062, 32'h41abda62} /* (12, 9, 29) {real, imag} */,
  {32'h3fcf32e0, 32'h414322f0} /* (12, 9, 28) {real, imag} */,
  {32'hc002d600, 32'h4167b4b3} /* (12, 9, 27) {real, imag} */,
  {32'hc0155034, 32'h3fbb2778} /* (12, 9, 26) {real, imag} */,
  {32'hc0d73cfd, 32'hc201e97d} /* (12, 9, 25) {real, imag} */,
  {32'h41501556, 32'h40fcfd58} /* (12, 9, 24) {real, imag} */,
  {32'hc20bc180, 32'h41886a4c} /* (12, 9, 23) {real, imag} */,
  {32'hc05c84ce, 32'hc04934f4} /* (12, 9, 22) {real, imag} */,
  {32'hbf8fe8c0, 32'hbfffc408} /* (12, 9, 21) {real, imag} */,
  {32'hc071bcb0, 32'hc101b488} /* (12, 9, 20) {real, imag} */,
  {32'h415c8446, 32'hc0abf698} /* (12, 9, 19) {real, imag} */,
  {32'h3fac4bda, 32'hc010cbd4} /* (12, 9, 18) {real, imag} */,
  {32'h3f454218, 32'hc108203e} /* (12, 9, 17) {real, imag} */,
  {32'h3fe45a90, 32'h40786a4c} /* (12, 9, 16) {real, imag} */,
  {32'hc09dea4b, 32'h402da198} /* (12, 9, 15) {real, imag} */,
  {32'hc0acbbc4, 32'h415ff24d} /* (12, 9, 14) {real, imag} */,
  {32'hc1378402, 32'h40e2161c} /* (12, 9, 13) {real, imag} */,
  {32'hc0fed9c4, 32'hc0591abf} /* (12, 9, 12) {real, imag} */,
  {32'h40ad698c, 32'h41af96fc} /* (12, 9, 11) {real, imag} */,
  {32'hc18b6ec5, 32'h41404f03} /* (12, 9, 10) {real, imag} */,
  {32'hc139cff2, 32'hc10397c1} /* (12, 9, 9) {real, imag} */,
  {32'hc15fd592, 32'hc031beb8} /* (12, 9, 8) {real, imag} */,
  {32'hc18740c1, 32'hc0872f38} /* (12, 9, 7) {real, imag} */,
  {32'h41a5a5fe, 32'hc0e2b95a} /* (12, 9, 6) {real, imag} */,
  {32'h42329ffe, 32'hc1b15226} /* (12, 9, 5) {real, imag} */,
  {32'hc1b91335, 32'h4164f0b0} /* (12, 9, 4) {real, imag} */,
  {32'hc1a07ca7, 32'hc241984b} /* (12, 9, 3) {real, imag} */,
  {32'hc106f09b, 32'hc0debbb0} /* (12, 9, 2) {real, imag} */,
  {32'hc27032d6, 32'hc1d14cea} /* (12, 9, 1) {real, imag} */,
  {32'h40f5385c, 32'hc1dd4998} /* (12, 9, 0) {real, imag} */,
  {32'hc1744732, 32'h42038520} /* (12, 8, 31) {real, imag} */,
  {32'hc203b15f, 32'hc2116f36} /* (12, 8, 30) {real, imag} */,
  {32'hc1960543, 32'h4185df73} /* (12, 8, 29) {real, imag} */,
  {32'h41aaa77e, 32'h4158b364} /* (12, 8, 28) {real, imag} */,
  {32'hc2014631, 32'h407ac144} /* (12, 8, 27) {real, imag} */,
  {32'h40c81c8c, 32'h41c6ea6d} /* (12, 8, 26) {real, imag} */,
  {32'h418411a2, 32'hc09a69b4} /* (12, 8, 25) {real, imag} */,
  {32'hc0a5acc4, 32'h41e19d64} /* (12, 8, 24) {real, imag} */,
  {32'h3f6bbb70, 32'h413173c0} /* (12, 8, 23) {real, imag} */,
  {32'hc1824fc0, 32'hc07f482e} /* (12, 8, 22) {real, imag} */,
  {32'h3f82461a, 32'h3f626e38} /* (12, 8, 21) {real, imag} */,
  {32'h3fbe9a08, 32'h3f411b68} /* (12, 8, 20) {real, imag} */,
  {32'hc0b0233c, 32'hc00f67ff} /* (12, 8, 19) {real, imag} */,
  {32'h404e792c, 32'hc033dc94} /* (12, 8, 18) {real, imag} */,
  {32'h40985358, 32'h40a81376} /* (12, 8, 17) {real, imag} */,
  {32'hc0889239, 32'h41444d9f} /* (12, 8, 16) {real, imag} */,
  {32'hbfeacf7e, 32'h40d6ab82} /* (12, 8, 15) {real, imag} */,
  {32'hc0cc9782, 32'h413cce85} /* (12, 8, 14) {real, imag} */,
  {32'h40f3c764, 32'hc07c1149} /* (12, 8, 13) {real, imag} */,
  {32'h4182febc, 32'hc0c702b5} /* (12, 8, 12) {real, imag} */,
  {32'h40936dd2, 32'h3f447118} /* (12, 8, 11) {real, imag} */,
  {32'hc12eb3c9, 32'hc0983ae1} /* (12, 8, 10) {real, imag} */,
  {32'hc1cf64e2, 32'hc13adff0} /* (12, 8, 9) {real, imag} */,
  {32'hc08d27be, 32'h4178dd95} /* (12, 8, 8) {real, imag} */,
  {32'h41dbd110, 32'h4141dd06} /* (12, 8, 7) {real, imag} */,
  {32'h41e69a67, 32'h40540888} /* (12, 8, 6) {real, imag} */,
  {32'h412b632c, 32'h41a8c4c2} /* (12, 8, 5) {real, imag} */,
  {32'h422a7147, 32'hc18b2fce} /* (12, 8, 4) {real, imag} */,
  {32'h423fd6ea, 32'h41aca789} /* (12, 8, 3) {real, imag} */,
  {32'h4272d849, 32'hc21bf6fe} /* (12, 8, 2) {real, imag} */,
  {32'h402466a0, 32'hc12f1978} /* (12, 8, 1) {real, imag} */,
  {32'h411412fa, 32'hbfa10db8} /* (12, 8, 0) {real, imag} */,
  {32'h41e1f404, 32'h41985fcc} /* (12, 7, 31) {real, imag} */,
  {32'hc040b2d0, 32'hc1640886} /* (12, 7, 30) {real, imag} */,
  {32'h41428a6b, 32'hc1db7a2c} /* (12, 7, 29) {real, imag} */,
  {32'h41a4ac36, 32'h41b6cb17} /* (12, 7, 28) {real, imag} */,
  {32'h41b8149a, 32'h4241e9ea} /* (12, 7, 27) {real, imag} */,
  {32'hc20d357d, 32'hc135cf71} /* (12, 7, 26) {real, imag} */,
  {32'hc1a9d244, 32'hc1d6ac42} /* (12, 7, 25) {real, imag} */,
  {32'hc1c1807e, 32'h4218e714} /* (12, 7, 24) {real, imag} */,
  {32'h4233a1f4, 32'h3fe66be9} /* (12, 7, 23) {real, imag} */,
  {32'h40cb09a6, 32'hc13a61fa} /* (12, 7, 22) {real, imag} */,
  {32'h40a64bae, 32'hc18a7334} /* (12, 7, 21) {real, imag} */,
  {32'hc0c3d19a, 32'h41263408} /* (12, 7, 20) {real, imag} */,
  {32'h40b56904, 32'h3e5d1500} /* (12, 7, 19) {real, imag} */,
  {32'hc1ae0dc4, 32'hc013d638} /* (12, 7, 18) {real, imag} */,
  {32'hc03e276e, 32'hc10ca5dc} /* (12, 7, 17) {real, imag} */,
  {32'h414fdfad, 32'hc1942e00} /* (12, 7, 16) {real, imag} */,
  {32'h40e3ef11, 32'h410f2618} /* (12, 7, 15) {real, imag} */,
  {32'h411e0a6f, 32'hc115470e} /* (12, 7, 14) {real, imag} */,
  {32'hbf917740, 32'hc13c3252} /* (12, 7, 13) {real, imag} */,
  {32'h41bd04ac, 32'h40c6f1e8} /* (12, 7, 12) {real, imag} */,
  {32'hc1a560ce, 32'h401e3f40} /* (12, 7, 11) {real, imag} */,
  {32'hc16436e7, 32'h413a7a9e} /* (12, 7, 10) {real, imag} */,
  {32'hc1820ddb, 32'hbff7f739} /* (12, 7, 9) {real, imag} */,
  {32'h41f708e6, 32'hc0ed0f32} /* (12, 7, 8) {real, imag} */,
  {32'hc17fbbbb, 32'hc1875cd6} /* (12, 7, 7) {real, imag} */,
  {32'hc1da78b3, 32'h4164cfaf} /* (12, 7, 6) {real, imag} */,
  {32'h4165b99c, 32'hc05414c0} /* (12, 7, 5) {real, imag} */,
  {32'h40efc54e, 32'hc204ac6e} /* (12, 7, 4) {real, imag} */,
  {32'h41f9d726, 32'hc20ec3ea} /* (12, 7, 3) {real, imag} */,
  {32'hc224bed3, 32'h42308b74} /* (12, 7, 2) {real, imag} */,
  {32'hc22ebef6, 32'h421c4eca} /* (12, 7, 1) {real, imag} */,
  {32'h42075487, 32'hc281af11} /* (12, 7, 0) {real, imag} */,
  {32'h41da360c, 32'hc25445b6} /* (12, 6, 31) {real, imag} */,
  {32'h41996a8a, 32'h42242be8} /* (12, 6, 30) {real, imag} */,
  {32'hc22f59e5, 32'hc1178ad6} /* (12, 6, 29) {real, imag} */,
  {32'hc18dd3dc, 32'hc1a463f8} /* (12, 6, 28) {real, imag} */,
  {32'h4195fbe0, 32'hc1f02df8} /* (12, 6, 27) {real, imag} */,
  {32'h41ca7da4, 32'hc23f8fca} /* (12, 6, 26) {real, imag} */,
  {32'h3f0cad60, 32'h41dd9b29} /* (12, 6, 25) {real, imag} */,
  {32'hc221bbf0, 32'hc2025e08} /* (12, 6, 24) {real, imag} */,
  {32'h40fab388, 32'h419b2e65} /* (12, 6, 23) {real, imag} */,
  {32'h4188b800, 32'h3fd28620} /* (12, 6, 22) {real, imag} */,
  {32'h4110bdb8, 32'h417759a6} /* (12, 6, 21) {real, imag} */,
  {32'hc0ed0121, 32'hc15b0fb8} /* (12, 6, 20) {real, imag} */,
  {32'h41050d29, 32'h41677f9e} /* (12, 6, 19) {real, imag} */,
  {32'h40b75c67, 32'hc0f8f8a8} /* (12, 6, 18) {real, imag} */,
  {32'hc13b0966, 32'h3f98bdd0} /* (12, 6, 17) {real, imag} */,
  {32'hc089dc34, 32'h4062eb08} /* (12, 6, 16) {real, imag} */,
  {32'h4042b678, 32'hbf68ade0} /* (12, 6, 15) {real, imag} */,
  {32'h4088a311, 32'h4198e49a} /* (12, 6, 14) {real, imag} */,
  {32'h410a029f, 32'h3fb6b5e4} /* (12, 6, 13) {real, imag} */,
  {32'hc0b01d7d, 32'hc0f0dc19} /* (12, 6, 12) {real, imag} */,
  {32'hc1d6225c, 32'hbea74fa0} /* (12, 6, 11) {real, imag} */,
  {32'h41681896, 32'h400a1f58} /* (12, 6, 10) {real, imag} */,
  {32'h40fbbe28, 32'h41412706} /* (12, 6, 9) {real, imag} */,
  {32'h40f789cc, 32'h4185a4ed} /* (12, 6, 8) {real, imag} */,
  {32'hc21607ae, 32'h41182cc6} /* (12, 6, 7) {real, imag} */,
  {32'h4220c28a, 32'hc11ee3f0} /* (12, 6, 6) {real, imag} */,
  {32'hc280f6f0, 32'hc117dc60} /* (12, 6, 5) {real, imag} */,
  {32'h413568cc, 32'hbfee76c0} /* (12, 6, 4) {real, imag} */,
  {32'h410e339c, 32'h40bd9359} /* (12, 6, 3) {real, imag} */,
  {32'h421c511a, 32'h4226eb6c} /* (12, 6, 2) {real, imag} */,
  {32'hc22e0eca, 32'hc22a172e} /* (12, 6, 1) {real, imag} */,
  {32'hc216b1d2, 32'h42282da2} /* (12, 6, 0) {real, imag} */,
  {32'h4239df72, 32'hc25e4e63} /* (12, 5, 31) {real, imag} */,
  {32'h42110c77, 32'h41043060} /* (12, 5, 30) {real, imag} */,
  {32'h41121b15, 32'h42a357ed} /* (12, 5, 29) {real, imag} */,
  {32'h41bd929d, 32'h42351a83} /* (12, 5, 28) {real, imag} */,
  {32'hc1c8daa0, 32'hc18245e1} /* (12, 5, 27) {real, imag} */,
  {32'h42255d77, 32'h41b86100} /* (12, 5, 26) {real, imag} */,
  {32'h40f7039c, 32'hc21b9558} /* (12, 5, 25) {real, imag} */,
  {32'hc089e0de, 32'hc22e4d36} /* (12, 5, 24) {real, imag} */,
  {32'hc2720b44, 32'h41c33cce} /* (12, 5, 23) {real, imag} */,
  {32'h41b22fb8, 32'h427d8888} /* (12, 5, 22) {real, imag} */,
  {32'hc165daa8, 32'hc16023ea} /* (12, 5, 21) {real, imag} */,
  {32'hc2077136, 32'hc0bba444} /* (12, 5, 20) {real, imag} */,
  {32'h3fbc0b78, 32'hc0ebd217} /* (12, 5, 19) {real, imag} */,
  {32'hbfcd1410, 32'hc18855ee} /* (12, 5, 18) {real, imag} */,
  {32'h4191a691, 32'h4104b59d} /* (12, 5, 17) {real, imag} */,
  {32'h3fdaf0b8, 32'h40721100} /* (12, 5, 16) {real, imag} */,
  {32'hc15f7a22, 32'hc1672171} /* (12, 5, 15) {real, imag} */,
  {32'h412ace6a, 32'hc148905c} /* (12, 5, 14) {real, imag} */,
  {32'hc050f6bc, 32'hc18e712a} /* (12, 5, 13) {real, imag} */,
  {32'h41c9f122, 32'h4185ec98} /* (12, 5, 12) {real, imag} */,
  {32'h41c5200a, 32'hc0e0f3c5} /* (12, 5, 11) {real, imag} */,
  {32'h40dd90da, 32'hc0260348} /* (12, 5, 10) {real, imag} */,
  {32'hc1422232, 32'h41710537} /* (12, 5, 9) {real, imag} */,
  {32'hc17fe42f, 32'h421187ae} /* (12, 5, 8) {real, imag} */,
  {32'h42419fd8, 32'h410e9b36} /* (12, 5, 7) {real, imag} */,
  {32'hc2b2b2dc, 32'hc0e76c58} /* (12, 5, 6) {real, imag} */,
  {32'hc20b0521, 32'h4191010b} /* (12, 5, 5) {real, imag} */,
  {32'hc15a62b2, 32'hc153a6c4} /* (12, 5, 4) {real, imag} */,
  {32'hc14f0e77, 32'h42a6abdb} /* (12, 5, 3) {real, imag} */,
  {32'hc2a26202, 32'hc29ae8d3} /* (12, 5, 2) {real, imag} */,
  {32'h420e17f6, 32'hc2815510} /* (12, 5, 1) {real, imag} */,
  {32'hc1ac6c2c, 32'hc1bdbc9a} /* (12, 5, 0) {real, imag} */,
  {32'h40e90000, 32'hc15b220a} /* (12, 4, 31) {real, imag} */,
  {32'h419042de, 32'hc280179a} /* (12, 4, 30) {real, imag} */,
  {32'hc2873935, 32'h422b9600} /* (12, 4, 29) {real, imag} */,
  {32'hc253e5dc, 32'h42a14448} /* (12, 4, 28) {real, imag} */,
  {32'h41efdf3c, 32'hc18e8a0c} /* (12, 4, 27) {real, imag} */,
  {32'h41715a7e, 32'hc129aa11} /* (12, 4, 26) {real, imag} */,
  {32'hc151e9d4, 32'h40587f34} /* (12, 4, 25) {real, imag} */,
  {32'h414db74c, 32'h4167650e} /* (12, 4, 24) {real, imag} */,
  {32'h4206c0aa, 32'hc11e2e43} /* (12, 4, 23) {real, imag} */,
  {32'hc15692bc, 32'h415e2ca0} /* (12, 4, 22) {real, imag} */,
  {32'h4219e7ae, 32'hc0730d04} /* (12, 4, 21) {real, imag} */,
  {32'hc1ca9093, 32'h4142deea} /* (12, 4, 20) {real, imag} */,
  {32'hc19db474, 32'h410a5643} /* (12, 4, 19) {real, imag} */,
  {32'hc072f778, 32'hc1f502a0} /* (12, 4, 18) {real, imag} */,
  {32'hbd556880, 32'h3f7887a8} /* (12, 4, 17) {real, imag} */,
  {32'h3fb5c180, 32'hc0d51cf8} /* (12, 4, 16) {real, imag} */,
  {32'h4019012a, 32'hc181d299} /* (12, 4, 15) {real, imag} */,
  {32'h3f6c46c0, 32'h400cdca0} /* (12, 4, 14) {real, imag} */,
  {32'h3e18b540, 32'hc0584ab4} /* (12, 4, 13) {real, imag} */,
  {32'h3f5f2c60, 32'h40964cb4} /* (12, 4, 12) {real, imag} */,
  {32'h40c4daa4, 32'h420aa82b} /* (12, 4, 11) {real, imag} */,
  {32'h419709ec, 32'h4160395e} /* (12, 4, 10) {real, imag} */,
  {32'h41909512, 32'hc189028a} /* (12, 4, 9) {real, imag} */,
  {32'h424c3427, 32'h41431b94} /* (12, 4, 8) {real, imag} */,
  {32'hbff15a40, 32'hc1b20e56} /* (12, 4, 7) {real, imag} */,
  {32'h418ca34f, 32'hc1b11b90} /* (12, 4, 6) {real, imag} */,
  {32'hc176bf74, 32'h428acbb7} /* (12, 4, 5) {real, imag} */,
  {32'hc1c941e8, 32'hc1368c40} /* (12, 4, 4) {real, imag} */,
  {32'h4229634e, 32'h41c0f310} /* (12, 4, 3) {real, imag} */,
  {32'h40bd6522, 32'h426bc412} /* (12, 4, 2) {real, imag} */,
  {32'h42214158, 32'h3f2e5918} /* (12, 4, 1) {real, imag} */,
  {32'hc279c51a, 32'hc1fba41a} /* (12, 4, 0) {real, imag} */,
  {32'h42a0e563, 32'hc1cef548} /* (12, 3, 31) {real, imag} */,
  {32'hc230436e, 32'h4134fe0d} /* (12, 3, 30) {real, imag} */,
  {32'h420c9093, 32'hc1dba062} /* (12, 3, 29) {real, imag} */,
  {32'hc2012ba2, 32'h428c25a4} /* (12, 3, 28) {real, imag} */,
  {32'hc1eee0e6, 32'hc16ad374} /* (12, 3, 27) {real, imag} */,
  {32'h41a60446, 32'hc10d2608} /* (12, 3, 26) {real, imag} */,
  {32'hc108c1a1, 32'hc1b164a6} /* (12, 3, 25) {real, imag} */,
  {32'h414b7880, 32'hc10a9a58} /* (12, 3, 24) {real, imag} */,
  {32'h40362a04, 32'h40d731fc} /* (12, 3, 23) {real, imag} */,
  {32'h4174ac5a, 32'hc0503024} /* (12, 3, 22) {real, imag} */,
  {32'h42185788, 32'h41dbd1e6} /* (12, 3, 21) {real, imag} */,
  {32'h410bc5f8, 32'hc11799ec} /* (12, 3, 20) {real, imag} */,
  {32'h4156f3c1, 32'h40b2843b} /* (12, 3, 19) {real, imag} */,
  {32'h4163de78, 32'h402d9658} /* (12, 3, 18) {real, imag} */,
  {32'hc1081c51, 32'h41473904} /* (12, 3, 17) {real, imag} */,
  {32'h3f26e920, 32'h4166657c} /* (12, 3, 16) {real, imag} */,
  {32'h41874b94, 32'h41b61132} /* (12, 3, 15) {real, imag} */,
  {32'hc16cf65c, 32'hbf66f360} /* (12, 3, 14) {real, imag} */,
  {32'h3feea7c8, 32'h3fac148c} /* (12, 3, 13) {real, imag} */,
  {32'hbfa7684c, 32'hc09139b8} /* (12, 3, 12) {real, imag} */,
  {32'h42041b44, 32'hbe7c0900} /* (12, 3, 11) {real, imag} */,
  {32'h3f9e94e0, 32'h418d088e} /* (12, 3, 10) {real, imag} */,
  {32'hbf3eb990, 32'hc22cef0a} /* (12, 3, 9) {real, imag} */,
  {32'h41a66de0, 32'h4082f797} /* (12, 3, 8) {real, imag} */,
  {32'hc1ce4934, 32'hc1b20da8} /* (12, 3, 7) {real, imag} */,
  {32'hc14b6d7d, 32'hc280eeb7} /* (12, 3, 6) {real, imag} */,
  {32'h40b2572a, 32'h4235840f} /* (12, 3, 5) {real, imag} */,
  {32'h417bde26, 32'hc09ce198} /* (12, 3, 4) {real, imag} */,
  {32'hc2ab519a, 32'h42333e0f} /* (12, 3, 3) {real, imag} */,
  {32'h4285df3d, 32'hc15bb1c7} /* (12, 3, 2) {real, imag} */,
  {32'hc1c08d70, 32'hc2071902} /* (12, 3, 1) {real, imag} */,
  {32'h42209e94, 32'h3f307e78} /* (12, 3, 0) {real, imag} */,
  {32'h400cbff8, 32'hc28cfc5c} /* (12, 2, 31) {real, imag} */,
  {32'hc1b59e44, 32'h41ca6282} /* (12, 2, 30) {real, imag} */,
  {32'hc221c840, 32'h4232f214} /* (12, 2, 29) {real, imag} */,
  {32'h420fba02, 32'hc1db6e9a} /* (12, 2, 28) {real, imag} */,
  {32'h423a4e15, 32'h4103b742} /* (12, 2, 27) {real, imag} */,
  {32'hc2b2e8c9, 32'hc1ac2086} /* (12, 2, 26) {real, imag} */,
  {32'h40a84640, 32'hc1259fee} /* (12, 2, 25) {real, imag} */,
  {32'h41873e3a, 32'h421b7c50} /* (12, 2, 24) {real, imag} */,
  {32'hc1f92078, 32'hc06b22b8} /* (12, 2, 23) {real, imag} */,
  {32'hc1e94135, 32'hc1eea461} /* (12, 2, 22) {real, imag} */,
  {32'h40990390, 32'h4235c908} /* (12, 2, 21) {real, imag} */,
  {32'h3f3a0a00, 32'hc1907c3f} /* (12, 2, 20) {real, imag} */,
  {32'hc11a1a77, 32'hc1357e52} /* (12, 2, 19) {real, imag} */,
  {32'hc19de40b, 32'h41a37c7d} /* (12, 2, 18) {real, imag} */,
  {32'h41b36c11, 32'h4127a75b} /* (12, 2, 17) {real, imag} */,
  {32'h404b05d0, 32'hc00f7028} /* (12, 2, 16) {real, imag} */,
  {32'hc0b6c37c, 32'hc0bbe1ea} /* (12, 2, 15) {real, imag} */,
  {32'h4108958a, 32'hc1d9faff} /* (12, 2, 14) {real, imag} */,
  {32'h4159ea97, 32'hc03f81fa} /* (12, 2, 13) {real, imag} */,
  {32'hc1f12470, 32'h415e3cc2} /* (12, 2, 12) {real, imag} */,
  {32'h41032a10, 32'hc11a0bea} /* (12, 2, 11) {real, imag} */,
  {32'hc1acded5, 32'hc18ed25b} /* (12, 2, 10) {real, imag} */,
  {32'h3fdd9f78, 32'hc2077f3a} /* (12, 2, 9) {real, imag} */,
  {32'hc210030d, 32'hc25411ea} /* (12, 2, 8) {real, imag} */,
  {32'h41173ada, 32'hc2942507} /* (12, 2, 7) {real, imag} */,
  {32'h427a63da, 32'h4244f425} /* (12, 2, 6) {real, imag} */,
  {32'hc1b12a42, 32'h41cf2c1b} /* (12, 2, 5) {real, imag} */,
  {32'hc09b192c, 32'hc25f0f8b} /* (12, 2, 4) {real, imag} */,
  {32'h41c3fc98, 32'hc232af90} /* (12, 2, 3) {real, imag} */,
  {32'hc1c7d76a, 32'h427ed7d3} /* (12, 2, 2) {real, imag} */,
  {32'h422892a8, 32'h42975bb0} /* (12, 2, 1) {real, imag} */,
  {32'hc19f942a, 32'h4174a20e} /* (12, 2, 0) {real, imag} */,
  {32'hc20e69fb, 32'hbe98e8a8} /* (12, 1, 31) {real, imag} */,
  {32'h428b096e, 32'hc1774362} /* (12, 1, 30) {real, imag} */,
  {32'h40f8a730, 32'h3f99aee0} /* (12, 1, 29) {real, imag} */,
  {32'hc2a43802, 32'h42238ab3} /* (12, 1, 28) {real, imag} */,
  {32'hc28d3774, 32'hc1853187} /* (12, 1, 27) {real, imag} */,
  {32'hc2270170, 32'hc1e1e575} /* (12, 1, 26) {real, imag} */,
  {32'h417f75ca, 32'h41126538} /* (12, 1, 25) {real, imag} */,
  {32'hc180c506, 32'h41d502be} /* (12, 1, 24) {real, imag} */,
  {32'h41494cee, 32'hc11c767b} /* (12, 1, 23) {real, imag} */,
  {32'hc137ed79, 32'h41e0469c} /* (12, 1, 22) {real, imag} */,
  {32'h4111e588, 32'h413a6dce} /* (12, 1, 21) {real, imag} */,
  {32'hc1b2888b, 32'hc1b86831} /* (12, 1, 20) {real, imag} */,
  {32'h3f2bb800, 32'hc1786197} /* (12, 1, 19) {real, imag} */,
  {32'hc0eec0fc, 32'hc0313dd2} /* (12, 1, 18) {real, imag} */,
  {32'h4146a46c, 32'hc0974420} /* (12, 1, 17) {real, imag} */,
  {32'h4151707c, 32'h407cb834} /* (12, 1, 16) {real, imag} */,
  {32'h406580f0, 32'h4100be9a} /* (12, 1, 15) {real, imag} */,
  {32'h3fa86e90, 32'hc011223e} /* (12, 1, 14) {real, imag} */,
  {32'h418604e7, 32'hc0db34d2} /* (12, 1, 13) {real, imag} */,
  {32'hc199d2c1, 32'h418771ef} /* (12, 1, 12) {real, imag} */,
  {32'h4198a855, 32'hc1d99ad9} /* (12, 1, 11) {real, imag} */,
  {32'hc11d4877, 32'hc1ab14b2} /* (12, 1, 10) {real, imag} */,
  {32'hc19e981d, 32'h41819cb2} /* (12, 1, 9) {real, imag} */,
  {32'h424551e5, 32'h41df6e2a} /* (12, 1, 8) {real, imag} */,
  {32'hc13f3a64, 32'h41f523f8} /* (12, 1, 7) {real, imag} */,
  {32'hc0d1a6f0, 32'h4250536e} /* (12, 1, 6) {real, imag} */,
  {32'hc0fedd18, 32'h42731924} /* (12, 1, 5) {real, imag} */,
  {32'hc2b2205a, 32'h41830164} /* (12, 1, 4) {real, imag} */,
  {32'h421f8336, 32'h420d662b} /* (12, 1, 3) {real, imag} */,
  {32'h4266efe8, 32'hc226b880} /* (12, 1, 2) {real, imag} */,
  {32'h41e34ff2, 32'h3ed40fe8} /* (12, 1, 1) {real, imag} */,
  {32'h426444cd, 32'h406c96b4} /* (12, 1, 0) {real, imag} */,
  {32'hc0e9a333, 32'h407bb528} /* (12, 0, 31) {real, imag} */,
  {32'hc24f7bba, 32'hc1ab0200} /* (12, 0, 30) {real, imag} */,
  {32'h41470246, 32'hc10980dc} /* (12, 0, 29) {real, imag} */,
  {32'h3e877540, 32'h41e91c41} /* (12, 0, 28) {real, imag} */,
  {32'h429641c2, 32'hc2b6d1fb} /* (12, 0, 27) {real, imag} */,
  {32'h42024de7, 32'hc21f8c36} /* (12, 0, 26) {real, imag} */,
  {32'hc0b52918, 32'h4210fd68} /* (12, 0, 25) {real, imag} */,
  {32'h427f22e7, 32'h4213374e} /* (12, 0, 24) {real, imag} */,
  {32'hc1905050, 32'h41a4f143} /* (12, 0, 23) {real, imag} */,
  {32'h417df618, 32'hc05c6c78} /* (12, 0, 22) {real, imag} */,
  {32'hc20fc0dc, 32'h3ff5fd08} /* (12, 0, 21) {real, imag} */,
  {32'h40b3f464, 32'hc1670b7a} /* (12, 0, 20) {real, imag} */,
  {32'h40d54f30, 32'hc2070339} /* (12, 0, 19) {real, imag} */,
  {32'h3f84ce18, 32'h41c17ca0} /* (12, 0, 18) {real, imag} */,
  {32'hc0897280, 32'hc0c294e6} /* (12, 0, 17) {real, imag} */,
  {32'hbff37480, 32'hc090c840} /* (12, 0, 16) {real, imag} */,
  {32'h40574e54, 32'h4183d1fc} /* (12, 0, 15) {real, imag} */,
  {32'h414e65d9, 32'hc0cbff82} /* (12, 0, 14) {real, imag} */,
  {32'hc09af6a0, 32'hc124209c} /* (12, 0, 13) {real, imag} */,
  {32'hc1a80b64, 32'hc1a30765} /* (12, 0, 12) {real, imag} */,
  {32'h40ced4e2, 32'hc18def90} /* (12, 0, 11) {real, imag} */,
  {32'h41367f90, 32'hc1eec6ed} /* (12, 0, 10) {real, imag} */,
  {32'h4253d6fc, 32'hc2457802} /* (12, 0, 9) {real, imag} */,
  {32'h41e5130a, 32'hc0b9eb54} /* (12, 0, 8) {real, imag} */,
  {32'hc145886c, 32'hc0771538} /* (12, 0, 7) {real, imag} */,
  {32'h42c8835c, 32'h423dc4e6} /* (12, 0, 6) {real, imag} */,
  {32'hc252234c, 32'hc112f848} /* (12, 0, 5) {real, imag} */,
  {32'h4204e0c6, 32'hc1abb39f} /* (12, 0, 4) {real, imag} */,
  {32'hc274e2b8, 32'h4128141c} /* (12, 0, 3) {real, imag} */,
  {32'hc1d3c8bc, 32'h426e0460} /* (12, 0, 2) {real, imag} */,
  {32'h4132baaa, 32'hc233e55a} /* (12, 0, 1) {real, imag} */,
  {32'hc2073d8b, 32'hc2455be4} /* (12, 0, 0) {real, imag} */,
  {32'h430d4776, 32'hc320538a} /* (11, 31, 31) {real, imag} */,
  {32'hc289a43c, 32'h43764092} /* (11, 31, 30) {real, imag} */,
  {32'hc0991804, 32'h420d4bd0} /* (11, 31, 29) {real, imag} */,
  {32'hc2bebe7a, 32'hc2d7c4ad} /* (11, 31, 28) {real, imag} */,
  {32'hc1ef38fe, 32'hc1a165d4} /* (11, 31, 27) {real, imag} */,
  {32'h42389141, 32'h41a22481} /* (11, 31, 26) {real, imag} */,
  {32'h4285bdf5, 32'hc22f07c0} /* (11, 31, 25) {real, imag} */,
  {32'h41daf502, 32'h4142eb14} /* (11, 31, 24) {real, imag} */,
  {32'hc2243c4c, 32'hc1cae4a5} /* (11, 31, 23) {real, imag} */,
  {32'hc22c252e, 32'h41ef137a} /* (11, 31, 22) {real, imag} */,
  {32'h41067405, 32'h423658d0} /* (11, 31, 21) {real, imag} */,
  {32'hbf5dc880, 32'h40cf60df} /* (11, 31, 20) {real, imag} */,
  {32'h41d8a5d1, 32'h415ccc25} /* (11, 31, 19) {real, imag} */,
  {32'hc0a76b00, 32'h420280e0} /* (11, 31, 18) {real, imag} */,
  {32'h4112317a, 32'h4196721e} /* (11, 31, 17) {real, imag} */,
  {32'h40e2bd40, 32'h40fc2c00} /* (11, 31, 16) {real, imag} */,
  {32'h4189a693, 32'hc163f0a4} /* (11, 31, 15) {real, imag} */,
  {32'hc1e3a3e4, 32'h3ef21840} /* (11, 31, 14) {real, imag} */,
  {32'h4143dfd2, 32'hc1df5954} /* (11, 31, 13) {real, imag} */,
  {32'hc1fb9914, 32'h40cd5031} /* (11, 31, 12) {real, imag} */,
  {32'hc20b16b5, 32'hc1b81a17} /* (11, 31, 11) {real, imag} */,
  {32'h4191dfb8, 32'hc2297f7f} /* (11, 31, 10) {real, imag} */,
  {32'h4246a48c, 32'h425289b2} /* (11, 31, 9) {real, imag} */,
  {32'hc2096141, 32'hbf546ac0} /* (11, 31, 8) {real, imag} */,
  {32'h416418b8, 32'hc1fef04f} /* (11, 31, 7) {real, imag} */,
  {32'h426435b3, 32'h42124966} /* (11, 31, 6) {real, imag} */,
  {32'hc17f8794, 32'h42caf0b9} /* (11, 31, 5) {real, imag} */,
  {32'h3c5b7000, 32'hc2a6146b} /* (11, 31, 4) {real, imag} */,
  {32'h425760d4, 32'hc2775eac} /* (11, 31, 3) {real, imag} */,
  {32'h4215ff2b, 32'h430131f6} /* (11, 31, 2) {real, imag} */,
  {32'h429548dc, 32'hc2072222} /* (11, 31, 1) {real, imag} */,
  {32'h4306ff40, 32'hc358d560} /* (11, 31, 0) {real, imag} */,
  {32'hc280c310, 32'h4294891f} /* (11, 30, 31) {real, imag} */,
  {32'h42eba64d, 32'hc0ce61f0} /* (11, 30, 30) {real, imag} */,
  {32'hc20e2f6b, 32'hc2732c48} /* (11, 30, 29) {real, imag} */,
  {32'h42ae31b9, 32'h4238a279} /* (11, 30, 28) {real, imag} */,
  {32'hc1d462d0, 32'hc1c3a18e} /* (11, 30, 27) {real, imag} */,
  {32'h41c051ba, 32'hc2dbbbd6} /* (11, 30, 26) {real, imag} */,
  {32'h417297c2, 32'hc2205430} /* (11, 30, 25) {real, imag} */,
  {32'h41db79fb, 32'hc1ff6c82} /* (11, 30, 24) {real, imag} */,
  {32'h4209f95e, 32'hc163660c} /* (11, 30, 23) {real, imag} */,
  {32'h425decc9, 32'h41ce6620} /* (11, 30, 22) {real, imag} */,
  {32'hc0db6ad2, 32'hc1fb6fc6} /* (11, 30, 21) {real, imag} */,
  {32'h410dfc94, 32'hc13959ea} /* (11, 30, 20) {real, imag} */,
  {32'h415358b2, 32'h41c1dbec} /* (11, 30, 19) {real, imag} */,
  {32'h4133eb32, 32'hc1b6815b} /* (11, 30, 18) {real, imag} */,
  {32'h41a4b153, 32'h4182b872} /* (11, 30, 17) {real, imag} */,
  {32'h4000b478, 32'h411af9d4} /* (11, 30, 16) {real, imag} */,
  {32'h3fa37f50, 32'hc17cf38c} /* (11, 30, 15) {real, imag} */,
  {32'h4000a638, 32'h40c77314} /* (11, 30, 14) {real, imag} */,
  {32'h41a049a5, 32'h40cf7880} /* (11, 30, 13) {real, imag} */,
  {32'hc23d0e29, 32'h41118dde} /* (11, 30, 12) {real, imag} */,
  {32'hc10f7f75, 32'hc1ad5d8e} /* (11, 30, 11) {real, imag} */,
  {32'h400d8d50, 32'hc1574148} /* (11, 30, 10) {real, imag} */,
  {32'hc2134392, 32'h40781610} /* (11, 30, 9) {real, imag} */,
  {32'h42106616, 32'hc15a49dc} /* (11, 30, 8) {real, imag} */,
  {32'h42509d80, 32'h40c90990} /* (11, 30, 7) {real, imag} */,
  {32'hc222ce93, 32'h40fdd178} /* (11, 30, 6) {real, imag} */,
  {32'h3ef690a0, 32'hc16465dc} /* (11, 30, 5) {real, imag} */,
  {32'hc22aa37e, 32'hc23a763f} /* (11, 30, 4) {real, imag} */,
  {32'hc2acd15c, 32'h41e1c09c} /* (11, 30, 3) {real, imag} */,
  {32'h432cbf0b, 32'hc2b403f1} /* (11, 30, 2) {real, imag} */,
  {32'hc342f9f4, 32'h429c5ac1} /* (11, 30, 1) {real, imag} */,
  {32'hc203b0f6, 32'h42dd8ec8} /* (11, 30, 0) {real, imag} */,
  {32'h4187a394, 32'hc2bf0c42} /* (11, 29, 31) {real, imag} */,
  {32'h425c8434, 32'h42d60e7f} /* (11, 29, 30) {real, imag} */,
  {32'hc1c972a4, 32'hc131a814} /* (11, 29, 29) {real, imag} */,
  {32'h40fe284c, 32'hc23b74ae} /* (11, 29, 28) {real, imag} */,
  {32'h4299076e, 32'hc23ead4f} /* (11, 29, 27) {real, imag} */,
  {32'h41e08b3c, 32'hc10cbc80} /* (11, 29, 26) {real, imag} */,
  {32'hc06f3524, 32'h41d1bff7} /* (11, 29, 25) {real, imag} */,
  {32'hc19ccc8b, 32'h4259d41a} /* (11, 29, 24) {real, imag} */,
  {32'hc0331c68, 32'hc1d48e92} /* (11, 29, 23) {real, imag} */,
  {32'h41a72fb4, 32'h3f01a550} /* (11, 29, 22) {real, imag} */,
  {32'hc1867d40, 32'hc06e61e4} /* (11, 29, 21) {real, imag} */,
  {32'hc1ad45d0, 32'hc1e9c514} /* (11, 29, 20) {real, imag} */,
  {32'h41144b29, 32'h412725a2} /* (11, 29, 19) {real, imag} */,
  {32'h40a1317a, 32'hbf8f0860} /* (11, 29, 18) {real, imag} */,
  {32'hc1877264, 32'hc1878241} /* (11, 29, 17) {real, imag} */,
  {32'h41b62bef, 32'hc219b96c} /* (11, 29, 16) {real, imag} */,
  {32'h410b1071, 32'hc09ca81c} /* (11, 29, 15) {real, imag} */,
  {32'hc1c31ebc, 32'h40985e28} /* (11, 29, 14) {real, imag} */,
  {32'h4204566e, 32'hc10b65f0} /* (11, 29, 13) {real, imag} */,
  {32'h406a91e0, 32'hc0812f46} /* (11, 29, 12) {real, imag} */,
  {32'hc0e02ae2, 32'hc0fe7556} /* (11, 29, 11) {real, imag} */,
  {32'h424354a6, 32'h402cc80c} /* (11, 29, 10) {real, imag} */,
  {32'hc242363e, 32'h41221d58} /* (11, 29, 9) {real, imag} */,
  {32'hc1b61d0f, 32'h419e34b1} /* (11, 29, 8) {real, imag} */,
  {32'h4120ee15, 32'h42a325d8} /* (11, 29, 7) {real, imag} */,
  {32'hc1efaed4, 32'hc2273786} /* (11, 29, 6) {real, imag} */,
  {32'h41f74d38, 32'hc20ba125} /* (11, 29, 5) {real, imag} */,
  {32'h41469f1e, 32'hc1d09cec} /* (11, 29, 4) {real, imag} */,
  {32'h41d250d0, 32'h418821d1} /* (11, 29, 3) {real, imag} */,
  {32'hc1778c28, 32'h430501ca} /* (11, 29, 2) {real, imag} */,
  {32'hc209c4f8, 32'hc20e8660} /* (11, 29, 1) {real, imag} */,
  {32'h41a25bbb, 32'h42329aaa} /* (11, 29, 0) {real, imag} */,
  {32'h428494e3, 32'h40dd209e} /* (11, 28, 31) {real, imag} */,
  {32'h42cbb9c2, 32'hc200d026} /* (11, 28, 30) {real, imag} */,
  {32'hc168265e, 32'hc25b00d2} /* (11, 28, 29) {real, imag} */,
  {32'hc1b12839, 32'hc161a820} /* (11, 28, 28) {real, imag} */,
  {32'h4155d43a, 32'hc22199c0} /* (11, 28, 27) {real, imag} */,
  {32'h4269aa88, 32'hc220d592} /* (11, 28, 26) {real, imag} */,
  {32'hc0ce6f33, 32'hc0e67b98} /* (11, 28, 25) {real, imag} */,
  {32'hc23b89de, 32'h421fd586} /* (11, 28, 24) {real, imag} */,
  {32'h417140f8, 32'hc1c6dffc} /* (11, 28, 23) {real, imag} */,
  {32'h41c08c6e, 32'hc201a738} /* (11, 28, 22) {real, imag} */,
  {32'hbff88d10, 32'hc09eb260} /* (11, 28, 21) {real, imag} */,
  {32'hc12bfeca, 32'h3f003d7a} /* (11, 28, 20) {real, imag} */,
  {32'h4173d2f2, 32'hc02819c8} /* (11, 28, 19) {real, imag} */,
  {32'h4009709e, 32'h41acfb1c} /* (11, 28, 18) {real, imag} */,
  {32'hc14fa39a, 32'hc106753c} /* (11, 28, 17) {real, imag} */,
  {32'h417597ca, 32'h41c293e5} /* (11, 28, 16) {real, imag} */,
  {32'hbf532120, 32'hc0b45ad4} /* (11, 28, 15) {real, imag} */,
  {32'hc18e983c, 32'hc08dbdae} /* (11, 28, 14) {real, imag} */,
  {32'hc199fa6b, 32'h41af7451} /* (11, 28, 13) {real, imag} */,
  {32'h41550b62, 32'hbe9485b4} /* (11, 28, 12) {real, imag} */,
  {32'h41656e4c, 32'hc0f8da08} /* (11, 28, 11) {real, imag} */,
  {32'hc107a22d, 32'hc098c42a} /* (11, 28, 10) {real, imag} */,
  {32'hc235742b, 32'hbf984040} /* (11, 28, 9) {real, imag} */,
  {32'hc217217a, 32'h4153dfa0} /* (11, 28, 8) {real, imag} */,
  {32'h41b365e9, 32'hc2481fc9} /* (11, 28, 7) {real, imag} */,
  {32'hc12075e8, 32'hc1e891a4} /* (11, 28, 6) {real, imag} */,
  {32'h418cccf6, 32'h41b9b2ea} /* (11, 28, 5) {real, imag} */,
  {32'hc0d9dfdb, 32'hc1041722} /* (11, 28, 4) {real, imag} */,
  {32'h4278e642, 32'hc31af20a} /* (11, 28, 3) {real, imag} */,
  {32'hc292191a, 32'h4213bc2e} /* (11, 28, 2) {real, imag} */,
  {32'hc1091692, 32'h41e1613c} /* (11, 28, 1) {real, imag} */,
  {32'h4029384a, 32'hbf3632a0} /* (11, 28, 0) {real, imag} */,
  {32'hc1befc9c, 32'h42aa75e4} /* (11, 27, 31) {real, imag} */,
  {32'hc2722a9f, 32'hc1d8b8a2} /* (11, 27, 30) {real, imag} */,
  {32'hc1c0c492, 32'hc22b1cfe} /* (11, 27, 29) {real, imag} */,
  {32'h418c2d41, 32'hbd747600} /* (11, 27, 28) {real, imag} */,
  {32'h42d37433, 32'h3f05fc80} /* (11, 27, 27) {real, imag} */,
  {32'hc22bb07a, 32'h41796038} /* (11, 27, 26) {real, imag} */,
  {32'hc18a63b3, 32'hc28b4743} /* (11, 27, 25) {real, imag} */,
  {32'h4242c687, 32'h42104904} /* (11, 27, 24) {real, imag} */,
  {32'h41b24884, 32'h411023e9} /* (11, 27, 23) {real, imag} */,
  {32'h40eeb320, 32'hc20a779c} /* (11, 27, 22) {real, imag} */,
  {32'h3fe8b840, 32'h4193f00e} /* (11, 27, 21) {real, imag} */,
  {32'hc117868e, 32'h41341fde} /* (11, 27, 20) {real, imag} */,
  {32'h409cf91e, 32'hc10ba4db} /* (11, 27, 19) {real, imag} */,
  {32'h40919668, 32'h41342a24} /* (11, 27, 18) {real, imag} */,
  {32'h41ad5810, 32'h41be5300} /* (11, 27, 17) {real, imag} */,
  {32'h41213b06, 32'h3fc92160} /* (11, 27, 16) {real, imag} */,
  {32'hc10a08dd, 32'h3f538650} /* (11, 27, 15) {real, imag} */,
  {32'hc0414ab0, 32'hbebb7680} /* (11, 27, 14) {real, imag} */,
  {32'h413f8c51, 32'hc0bdd6de} /* (11, 27, 13) {real, imag} */,
  {32'h412d9572, 32'hbffe4e90} /* (11, 27, 12) {real, imag} */,
  {32'hc1149908, 32'h414ae0dd} /* (11, 27, 11) {real, imag} */,
  {32'hc1a339e6, 32'hc19b1f30} /* (11, 27, 10) {real, imag} */,
  {32'h41a31bd0, 32'h40e8a2a2} /* (11, 27, 9) {real, imag} */,
  {32'h42157e7d, 32'hc17a71d6} /* (11, 27, 8) {real, imag} */,
  {32'hc1937e91, 32'h42185611} /* (11, 27, 7) {real, imag} */,
  {32'hc0f2b058, 32'h4265d54c} /* (11, 27, 6) {real, imag} */,
  {32'hc1678428, 32'hc25e6348} /* (11, 27, 5) {real, imag} */,
  {32'hc1da71c3, 32'hc1c0ead3} /* (11, 27, 4) {real, imag} */,
  {32'h4114d3bc, 32'h417563fd} /* (11, 27, 3) {real, imag} */,
  {32'h41a61e76, 32'hc31715bf} /* (11, 27, 2) {real, imag} */,
  {32'hc1f9600c, 32'h40b73e48} /* (11, 27, 1) {real, imag} */,
  {32'hc257f2c6, 32'h42c22abe} /* (11, 27, 0) {real, imag} */,
  {32'h4155eff0, 32'hc25212c8} /* (11, 26, 31) {real, imag} */,
  {32'hc289fc6e, 32'hc2b7a09a} /* (11, 26, 30) {real, imag} */,
  {32'hc2073a15, 32'h425e2b1c} /* (11, 26, 29) {real, imag} */,
  {32'h42515cbe, 32'h4248e2d8} /* (11, 26, 28) {real, imag} */,
  {32'h419e81d4, 32'hc0235c08} /* (11, 26, 27) {real, imag} */,
  {32'h41a1969a, 32'hc1582df1} /* (11, 26, 26) {real, imag} */,
  {32'h42277ea5, 32'hc1ff8399} /* (11, 26, 25) {real, imag} */,
  {32'hc1296658, 32'h40fe0046} /* (11, 26, 24) {real, imag} */,
  {32'hc0b39920, 32'hc1ab9bfe} /* (11, 26, 23) {real, imag} */,
  {32'h408a370d, 32'hc04c2974} /* (11, 26, 22) {real, imag} */,
  {32'h41d045e0, 32'h41db22aa} /* (11, 26, 21) {real, imag} */,
  {32'hc18660d4, 32'h41138002} /* (11, 26, 20) {real, imag} */,
  {32'hc13cb9ca, 32'h4128edc8} /* (11, 26, 19) {real, imag} */,
  {32'hc151119c, 32'hc1be564e} /* (11, 26, 18) {real, imag} */,
  {32'h41463c53, 32'h41306b92} /* (11, 26, 17) {real, imag} */,
  {32'hc106efa0, 32'h409e4400} /* (11, 26, 16) {real, imag} */,
  {32'hc18ab08c, 32'hbf64c758} /* (11, 26, 15) {real, imag} */,
  {32'h40eafa18, 32'hc1ae30f6} /* (11, 26, 14) {real, imag} */,
  {32'h411ca126, 32'h414ddaa4} /* (11, 26, 13) {real, imag} */,
  {32'h414395f7, 32'hc0a2916b} /* (11, 26, 12) {real, imag} */,
  {32'hc150d5a8, 32'h4138563c} /* (11, 26, 11) {real, imag} */,
  {32'hc043c252, 32'h41bd28da} /* (11, 26, 10) {real, imag} */,
  {32'h4270e7d0, 32'h41ff895c} /* (11, 26, 9) {real, imag} */,
  {32'h41c67344, 32'hc21db5ab} /* (11, 26, 8) {real, imag} */,
  {32'hc0916fa8, 32'h405432e8} /* (11, 26, 7) {real, imag} */,
  {32'h420d0bd7, 32'hc18a9c4a} /* (11, 26, 6) {real, imag} */,
  {32'hc247138e, 32'hc20bbf44} /* (11, 26, 5) {real, imag} */,
  {32'hc18458dc, 32'hc1b82548} /* (11, 26, 4) {real, imag} */,
  {32'hc205ae7b, 32'h41a82389} /* (11, 26, 3) {real, imag} */,
  {32'hc183f9be, 32'hc208374d} /* (11, 26, 2) {real, imag} */,
  {32'hc1958bb8, 32'h41be6579} /* (11, 26, 1) {real, imag} */,
  {32'h42291b32, 32'h4238cd32} /* (11, 26, 0) {real, imag} */,
  {32'h41ea7214, 32'h40e5e9e9} /* (11, 25, 31) {real, imag} */,
  {32'hbf8de828, 32'hc179348d} /* (11, 25, 30) {real, imag} */,
  {32'hc1a14948, 32'h420bb1f7} /* (11, 25, 29) {real, imag} */,
  {32'hc03a133c, 32'hc140280e} /* (11, 25, 28) {real, imag} */,
  {32'hc1854235, 32'hc1ab69e4} /* (11, 25, 27) {real, imag} */,
  {32'hc222b267, 32'h418a9b8f} /* (11, 25, 26) {real, imag} */,
  {32'hc176e71a, 32'h41870b93} /* (11, 25, 25) {real, imag} */,
  {32'h41438c02, 32'h41b81b47} /* (11, 25, 24) {real, imag} */,
  {32'hc1511aca, 32'hc1a5c251} /* (11, 25, 23) {real, imag} */,
  {32'hc13db709, 32'h4187b74e} /* (11, 25, 22) {real, imag} */,
  {32'hc0307bb6, 32'hc1068599} /* (11, 25, 21) {real, imag} */,
  {32'h41805aba, 32'hc1b9158d} /* (11, 25, 20) {real, imag} */,
  {32'h41359a02, 32'h400b3b80} /* (11, 25, 19) {real, imag} */,
  {32'hc1909170, 32'hc147f7c5} /* (11, 25, 18) {real, imag} */,
  {32'h41275060, 32'h4131d287} /* (11, 25, 17) {real, imag} */,
  {32'h3d8c6d00, 32'h3f9d8c30} /* (11, 25, 16) {real, imag} */,
  {32'hc10f7018, 32'h41ba790c} /* (11, 25, 15) {real, imag} */,
  {32'hc0b6b6c8, 32'h3fe35dc8} /* (11, 25, 14) {real, imag} */,
  {32'hbfa2a45c, 32'hc09b4430} /* (11, 25, 13) {real, imag} */,
  {32'hbdc55280, 32'h41988af7} /* (11, 25, 12) {real, imag} */,
  {32'h402cd07a, 32'h412b2521} /* (11, 25, 11) {real, imag} */,
  {32'h41ba7b48, 32'hc1c1ac10} /* (11, 25, 10) {real, imag} */,
  {32'hc19ab7a5, 32'hc13765de} /* (11, 25, 9) {real, imag} */,
  {32'h41ed3a45, 32'hc18d0b4d} /* (11, 25, 8) {real, imag} */,
  {32'h3e6eed80, 32'h41b3edf9} /* (11, 25, 7) {real, imag} */,
  {32'hc201cd27, 32'hc26d8d9c} /* (11, 25, 6) {real, imag} */,
  {32'h41c26285, 32'hc26e96ba} /* (11, 25, 5) {real, imag} */,
  {32'h41e4aae4, 32'h4198b6c5} /* (11, 25, 4) {real, imag} */,
  {32'hc0e170b6, 32'h412a76db} /* (11, 25, 3) {real, imag} */,
  {32'h40f9421a, 32'hc239d33e} /* (11, 25, 2) {real, imag} */,
  {32'hc20ad1ca, 32'h407d37ae} /* (11, 25, 1) {real, imag} */,
  {32'h426a3984, 32'h41d3deef} /* (11, 25, 0) {real, imag} */,
  {32'hc1a93e84, 32'hc0aa7c48} /* (11, 24, 31) {real, imag} */,
  {32'hc25935be, 32'h41a99542} /* (11, 24, 30) {real, imag} */,
  {32'h420949d2, 32'hc20615c6} /* (11, 24, 29) {real, imag} */,
  {32'h40d5acb6, 32'h4237095b} /* (11, 24, 28) {real, imag} */,
  {32'h42261b36, 32'hc20a68c3} /* (11, 24, 27) {real, imag} */,
  {32'hc217da00, 32'hc027f260} /* (11, 24, 26) {real, imag} */,
  {32'hc1cded48, 32'hc22e9366} /* (11, 24, 25) {real, imag} */,
  {32'hc20654dc, 32'hc15a359e} /* (11, 24, 24) {real, imag} */,
  {32'hc0e5ed30, 32'h40fe76f4} /* (11, 24, 23) {real, imag} */,
  {32'h41864f6b, 32'h41140210} /* (11, 24, 22) {real, imag} */,
  {32'hc0aca659, 32'h404739ac} /* (11, 24, 21) {real, imag} */,
  {32'hc1411c0f, 32'hc0436292} /* (11, 24, 20) {real, imag} */,
  {32'h40fe12d6, 32'hc1921d7c} /* (11, 24, 19) {real, imag} */,
  {32'hc1163667, 32'hc0ffa5ce} /* (11, 24, 18) {real, imag} */,
  {32'hc036f746, 32'hbff916d8} /* (11, 24, 17) {real, imag} */,
  {32'h4145b57c, 32'h414e7ab6} /* (11, 24, 16) {real, imag} */,
  {32'h40bd637b, 32'hc02f4e0c} /* (11, 24, 15) {real, imag} */,
  {32'hbdb6cb80, 32'hbec083a0} /* (11, 24, 14) {real, imag} */,
  {32'h41653eb9, 32'hc0866811} /* (11, 24, 13) {real, imag} */,
  {32'hc08824c2, 32'hc1108fb8} /* (11, 24, 12) {real, imag} */,
  {32'hc18a7adb, 32'hc06d1144} /* (11, 24, 11) {real, imag} */,
  {32'hc12632d2, 32'h41bb1ca2} /* (11, 24, 10) {real, imag} */,
  {32'hc2244e90, 32'h418a12c1} /* (11, 24, 9) {real, imag} */,
  {32'h4129f5f6, 32'hc1b181ff} /* (11, 24, 8) {real, imag} */,
  {32'h41ca8d28, 32'h4221d34c} /* (11, 24, 7) {real, imag} */,
  {32'h428bbc57, 32'hc1218d29} /* (11, 24, 6) {real, imag} */,
  {32'hbfa40a40, 32'h41138048} /* (11, 24, 5) {real, imag} */,
  {32'h4201e131, 32'hc19028e8} /* (11, 24, 4) {real, imag} */,
  {32'h4143f98c, 32'hc00e95b8} /* (11, 24, 3) {real, imag} */,
  {32'h425ef466, 32'h4233c9a3} /* (11, 24, 2) {real, imag} */,
  {32'hc20d9900, 32'h4258d795} /* (11, 24, 1) {real, imag} */,
  {32'hc24ffd39, 32'h4298cf35} /* (11, 24, 0) {real, imag} */,
  {32'hc0b1d9d0, 32'h414d79f0} /* (11, 23, 31) {real, imag} */,
  {32'hc29449a8, 32'h42472b46} /* (11, 23, 30) {real, imag} */,
  {32'h4201c438, 32'hc158ca97} /* (11, 23, 29) {real, imag} */,
  {32'hc1ab045d, 32'hc1497743} /* (11, 23, 28) {real, imag} */,
  {32'hc1eb4770, 32'hc13f9a3c} /* (11, 23, 27) {real, imag} */,
  {32'h41f87a04, 32'hc1ec6153} /* (11, 23, 26) {real, imag} */,
  {32'hc2137219, 32'h417f32c6} /* (11, 23, 25) {real, imag} */,
  {32'h4170bf8a, 32'h415285f4} /* (11, 23, 24) {real, imag} */,
  {32'h4190c7ee, 32'hc132a712} /* (11, 23, 23) {real, imag} */,
  {32'h41eff376, 32'hc14157a8} /* (11, 23, 22) {real, imag} */,
  {32'hc1802b26, 32'h414b884b} /* (11, 23, 21) {real, imag} */,
  {32'h4089abdd, 32'h4038edbe} /* (11, 23, 20) {real, imag} */,
  {32'hc12d6180, 32'hc0a4461a} /* (11, 23, 19) {real, imag} */,
  {32'hc1449150, 32'h3fa06b40} /* (11, 23, 18) {real, imag} */,
  {32'h4075afb4, 32'hc055dd0a} /* (11, 23, 17) {real, imag} */,
  {32'h40d6b485, 32'h40bac172} /* (11, 23, 16) {real, imag} */,
  {32'hc0ccb020, 32'h40b1947d} /* (11, 23, 15) {real, imag} */,
  {32'h400b05b2, 32'h3fb17530} /* (11, 23, 14) {real, imag} */,
  {32'h3fc145a4, 32'h401be8fc} /* (11, 23, 13) {real, imag} */,
  {32'hbf9cfa74, 32'hc0d772a1} /* (11, 23, 12) {real, imag} */,
  {32'h40ae5b1e, 32'hc1855748} /* (11, 23, 11) {real, imag} */,
  {32'h4024f070, 32'h414c64c4} /* (11, 23, 10) {real, imag} */,
  {32'h41d4a82e, 32'h3f26ef88} /* (11, 23, 9) {real, imag} */,
  {32'h41e809a7, 32'h41bf3866} /* (11, 23, 8) {real, imag} */,
  {32'h4127f644, 32'h417007d4} /* (11, 23, 7) {real, imag} */,
  {32'h419c29a4, 32'h4150e76e} /* (11, 23, 6) {real, imag} */,
  {32'hc1fa393c, 32'hc2179d93} /* (11, 23, 5) {real, imag} */,
  {32'hc11a9b86, 32'hc18ab6f8} /* (11, 23, 4) {real, imag} */,
  {32'hc1060800, 32'h423167b7} /* (11, 23, 3) {real, imag} */,
  {32'hc1e6b4f1, 32'h40e85f70} /* (11, 23, 2) {real, imag} */,
  {32'hc1d527e4, 32'h41aa1af6} /* (11, 23, 1) {real, imag} */,
  {32'h4166de3e, 32'hc17134df} /* (11, 23, 0) {real, imag} */,
  {32'h4000e0c2, 32'hc24c660a} /* (11, 22, 31) {real, imag} */,
  {32'h405d647a, 32'hc19ae988} /* (11, 22, 30) {real, imag} */,
  {32'hc12d0ac2, 32'h4170e4ac} /* (11, 22, 29) {real, imag} */,
  {32'hc241173b, 32'h416ead7a} /* (11, 22, 28) {real, imag} */,
  {32'h41f4027c, 32'h41e3d9d9} /* (11, 22, 27) {real, imag} */,
  {32'h41c0743e, 32'h41a58562} /* (11, 22, 26) {real, imag} */,
  {32'h41c3c21a, 32'h403a21e8} /* (11, 22, 25) {real, imag} */,
  {32'h420c3be8, 32'h4090fa8c} /* (11, 22, 24) {real, imag} */,
  {32'hc116cfd8, 32'h422c84c5} /* (11, 22, 23) {real, imag} */,
  {32'hc182a792, 32'hc0158642} /* (11, 22, 22) {real, imag} */,
  {32'hbffecff0, 32'hc1b391b6} /* (11, 22, 21) {real, imag} */,
  {32'hc10d758c, 32'hc08cc6b0} /* (11, 22, 20) {real, imag} */,
  {32'hc0ecfb42, 32'h405d419c} /* (11, 22, 19) {real, imag} */,
  {32'h41ee7dd1, 32'hc11b8c20} /* (11, 22, 18) {real, imag} */,
  {32'hc09afef4, 32'h3d3b9780} /* (11, 22, 17) {real, imag} */,
  {32'hc0f4a720, 32'hbfa52f34} /* (11, 22, 16) {real, imag} */,
  {32'hbefe4f58, 32'h4147a950} /* (11, 22, 15) {real, imag} */,
  {32'hc0e7eecc, 32'h4189c7a1} /* (11, 22, 14) {real, imag} */,
  {32'h3d0d1400, 32'h416de2b5} /* (11, 22, 13) {real, imag} */,
  {32'hc14de526, 32'hbec59a88} /* (11, 22, 12) {real, imag} */,
  {32'h41a22179, 32'hbf2ee670} /* (11, 22, 11) {real, imag} */,
  {32'h4180d530, 32'h3cb6e100} /* (11, 22, 10) {real, imag} */,
  {32'hc1443090, 32'hc20a025d} /* (11, 22, 9) {real, imag} */,
  {32'h41c4d3a0, 32'h41b51c80} /* (11, 22, 8) {real, imag} */,
  {32'h418524bc, 32'hbfd93bf0} /* (11, 22, 7) {real, imag} */,
  {32'h41e4c802, 32'h418c10d6} /* (11, 22, 6) {real, imag} */,
  {32'hc1f32f7c, 32'hc140f8ae} /* (11, 22, 5) {real, imag} */,
  {32'hc18a684e, 32'hbfcb47f0} /* (11, 22, 4) {real, imag} */,
  {32'h414434a6, 32'hbf3e1c08} /* (11, 22, 3) {real, imag} */,
  {32'hc03a644e, 32'hc0d5a9ae} /* (11, 22, 2) {real, imag} */,
  {32'hbfc12aa9, 32'hc11ab53a} /* (11, 22, 1) {real, imag} */,
  {32'h406ae998, 32'h41487578} /* (11, 22, 0) {real, imag} */,
  {32'hc1ceacf7, 32'h42531e3e} /* (11, 21, 31) {real, imag} */,
  {32'h406aae7c, 32'hc1182140} /* (11, 21, 30) {real, imag} */,
  {32'h416bfbee, 32'hc254d5e8} /* (11, 21, 29) {real, imag} */,
  {32'hc1dd5bf5, 32'h3fc66b60} /* (11, 21, 28) {real, imag} */,
  {32'hc0e91212, 32'h411d86eb} /* (11, 21, 27) {real, imag} */,
  {32'h41c84b37, 32'h411a76a3} /* (11, 21, 26) {real, imag} */,
  {32'h417eb9da, 32'hc2239c34} /* (11, 21, 25) {real, imag} */,
  {32'hc2062f36, 32'hc16302e8} /* (11, 21, 24) {real, imag} */,
  {32'h40bce661, 32'h41adf12a} /* (11, 21, 23) {real, imag} */,
  {32'h3d978360, 32'h40a531c7} /* (11, 21, 22) {real, imag} */,
  {32'h40788245, 32'h3e0d7d80} /* (11, 21, 21) {real, imag} */,
  {32'h3fb898ce, 32'h40930e81} /* (11, 21, 20) {real, imag} */,
  {32'h40982b64, 32'hc082a33c} /* (11, 21, 19) {real, imag} */,
  {32'h4019c172, 32'h41358f81} /* (11, 21, 18) {real, imag} */,
  {32'hc09e2f3a, 32'hbf7bfa80} /* (11, 21, 17) {real, imag} */,
  {32'hc132d93a, 32'h40257db6} /* (11, 21, 16) {real, imag} */,
  {32'h4085bb76, 32'hc09c38b0} /* (11, 21, 15) {real, imag} */,
  {32'hc03f1ca6, 32'hbf776760} /* (11, 21, 14) {real, imag} */,
  {32'h409be090, 32'hc0903dc4} /* (11, 21, 13) {real, imag} */,
  {32'hc07e8479, 32'h4175e860} /* (11, 21, 12) {real, imag} */,
  {32'hc1090e1f, 32'hc062ba88} /* (11, 21, 11) {real, imag} */,
  {32'hc0f53d72, 32'hc0d56dff} /* (11, 21, 10) {real, imag} */,
  {32'h4168bc44, 32'hbd168c00} /* (11, 21, 9) {real, imag} */,
  {32'hc0e06018, 32'hbf170580} /* (11, 21, 8) {real, imag} */,
  {32'h41a10039, 32'hbf062260} /* (11, 21, 7) {real, imag} */,
  {32'hc194e0fd, 32'hc186c57c} /* (11, 21, 6) {real, imag} */,
  {32'h40cd5472, 32'h4199b16e} /* (11, 21, 5) {real, imag} */,
  {32'h417e0296, 32'h41b26d3e} /* (11, 21, 4) {real, imag} */,
  {32'hc2110034, 32'hc18cd817} /* (11, 21, 3) {real, imag} */,
  {32'h41ba0e2e, 32'hc12d9754} /* (11, 21, 2) {real, imag} */,
  {32'h41c00fbd, 32'h420bf7ea} /* (11, 21, 1) {real, imag} */,
  {32'hc239f3d6, 32'h3fbcd2e4} /* (11, 21, 0) {real, imag} */,
  {32'h3fb47ff2, 32'h40a7e1b4} /* (11, 20, 31) {real, imag} */,
  {32'h4184859d, 32'h407c7b22} /* (11, 20, 30) {real, imag} */,
  {32'hbf9fadd0, 32'h416a91f0} /* (11, 20, 29) {real, imag} */,
  {32'hc15f6597, 32'hc1005cc2} /* (11, 20, 28) {real, imag} */,
  {32'h41bf2650, 32'hc1018c28} /* (11, 20, 27) {real, imag} */,
  {32'hc1e9a75e, 32'hc14e3ee1} /* (11, 20, 26) {real, imag} */,
  {32'h407249f4, 32'h40684dd0} /* (11, 20, 25) {real, imag} */,
  {32'h40732566, 32'h4158c08d} /* (11, 20, 24) {real, imag} */,
  {32'hc1c34c36, 32'hc0dfc2a0} /* (11, 20, 23) {real, imag} */,
  {32'hc1c458c7, 32'h41544aac} /* (11, 20, 22) {real, imag} */,
  {32'h40d3998e, 32'h3f906f78} /* (11, 20, 21) {real, imag} */,
  {32'hc09ab1da, 32'hc13cee3e} /* (11, 20, 20) {real, imag} */,
  {32'h4107a436, 32'h40a34755} /* (11, 20, 19) {real, imag} */,
  {32'hc0c3d695, 32'h3f15e018} /* (11, 20, 18) {real, imag} */,
  {32'h4065686e, 32'h409c107c} /* (11, 20, 17) {real, imag} */,
  {32'hc09a0e62, 32'hc040c5c4} /* (11, 20, 16) {real, imag} */,
  {32'hc0a5c895, 32'hc0dd82d0} /* (11, 20, 15) {real, imag} */,
  {32'h410c0cee, 32'hc10384f6} /* (11, 20, 14) {real, imag} */,
  {32'h40a8efdd, 32'hc124cd00} /* (11, 20, 13) {real, imag} */,
  {32'h411679ce, 32'hc102d17e} /* (11, 20, 12) {real, imag} */,
  {32'hc0c99786, 32'hc01931b4} /* (11, 20, 11) {real, imag} */,
  {32'hc09e478c, 32'h41def39a} /* (11, 20, 10) {real, imag} */,
  {32'hbe5cecc0, 32'h409ec43c} /* (11, 20, 9) {real, imag} */,
  {32'hc1804592, 32'h412bcc23} /* (11, 20, 8) {real, imag} */,
  {32'h4139c645, 32'hc17fe1be} /* (11, 20, 7) {real, imag} */,
  {32'h40ad8990, 32'h4122fad7} /* (11, 20, 6) {real, imag} */,
  {32'hc1465fc9, 32'h42004b7b} /* (11, 20, 5) {real, imag} */,
  {32'hbf8bdfb0, 32'h410c15ec} /* (11, 20, 4) {real, imag} */,
  {32'h41e28f0b, 32'hbfdc470c} /* (11, 20, 3) {real, imag} */,
  {32'hc1768ade, 32'h416f62b8} /* (11, 20, 2) {real, imag} */,
  {32'hc0bf7c30, 32'hc171cc78} /* (11, 20, 1) {real, imag} */,
  {32'hc1d45020, 32'hc194377c} /* (11, 20, 0) {real, imag} */,
  {32'h420061b8, 32'hc19b7b61} /* (11, 19, 31) {real, imag} */,
  {32'h41a02180, 32'h401ced28} /* (11, 19, 30) {real, imag} */,
  {32'h41b3df28, 32'h41e1d8ea} /* (11, 19, 29) {real, imag} */,
  {32'h42006e3d, 32'hc18c646e} /* (11, 19, 28) {real, imag} */,
  {32'h410550aa, 32'hc184f58a} /* (11, 19, 27) {real, imag} */,
  {32'hc0e7b45d, 32'h41dd7822} /* (11, 19, 26) {real, imag} */,
  {32'hbb599400, 32'hc1202f0a} /* (11, 19, 25) {real, imag} */,
  {32'h4114b044, 32'hc082d394} /* (11, 19, 24) {real, imag} */,
  {32'hc1c9ed0c, 32'h41164f74} /* (11, 19, 23) {real, imag} */,
  {32'h407d8548, 32'h415fe86a} /* (11, 19, 22) {real, imag} */,
  {32'hc17d69f4, 32'hc0b0b02e} /* (11, 19, 21) {real, imag} */,
  {32'hbe4648a0, 32'h4120fa0c} /* (11, 19, 20) {real, imag} */,
  {32'h3f82a570, 32'hbf8f917c} /* (11, 19, 19) {real, imag} */,
  {32'h4089797c, 32'h3fc8d9bc} /* (11, 19, 18) {real, imag} */,
  {32'hbfdbb158, 32'hc0ea7988} /* (11, 19, 17) {real, imag} */,
  {32'h3f6c8304, 32'hc09f61e2} /* (11, 19, 16) {real, imag} */,
  {32'h40b769aa, 32'hc0680468} /* (11, 19, 15) {real, imag} */,
  {32'hc0bc5070, 32'hbfa056c4} /* (11, 19, 14) {real, imag} */,
  {32'h3fbf2d80, 32'hc095f447} /* (11, 19, 13) {real, imag} */,
  {32'hbda015c0, 32'h3ff53af0} /* (11, 19, 12) {real, imag} */,
  {32'hc080f8c0, 32'h3f93bf28} /* (11, 19, 11) {real, imag} */,
  {32'hc08936f8, 32'hc0b9f9dc} /* (11, 19, 10) {real, imag} */,
  {32'h419116a0, 32'hc137c34c} /* (11, 19, 9) {real, imag} */,
  {32'hc056e3d8, 32'hc119afae} /* (11, 19, 8) {real, imag} */,
  {32'hc0dfc442, 32'h41960771} /* (11, 19, 7) {real, imag} */,
  {32'h412f52eb, 32'h4156625c} /* (11, 19, 6) {real, imag} */,
  {32'h4023ad27, 32'h4154e6a8} /* (11, 19, 5) {real, imag} */,
  {32'h4115afc4, 32'h4117ab7f} /* (11, 19, 4) {real, imag} */,
  {32'hc0925fee, 32'hc197f368} /* (11, 19, 3) {real, imag} */,
  {32'hbea0dee0, 32'hc10f43ad} /* (11, 19, 2) {real, imag} */,
  {32'hc11d1837, 32'hc0bc1e38} /* (11, 19, 1) {real, imag} */,
  {32'hbf6157a4, 32'hc1290c3f} /* (11, 19, 0) {real, imag} */,
  {32'h4156df6e, 32'h419ea27f} /* (11, 18, 31) {real, imag} */,
  {32'h419f5c11, 32'h41e38ce6} /* (11, 18, 30) {real, imag} */,
  {32'hc0949984, 32'hc0ac60fc} /* (11, 18, 29) {real, imag} */,
  {32'h4008aefe, 32'hc0d9b87a} /* (11, 18, 28) {real, imag} */,
  {32'hc1164c67, 32'h41797052} /* (11, 18, 27) {real, imag} */,
  {32'h3f4e51f4, 32'hc0e5c16e} /* (11, 18, 26) {real, imag} */,
  {32'h417128df, 32'hbfe98b6c} /* (11, 18, 25) {real, imag} */,
  {32'hc13f1745, 32'h40ceb832} /* (11, 18, 24) {real, imag} */,
  {32'h3f1e89a0, 32'h4197bc89} /* (11, 18, 23) {real, imag} */,
  {32'h4077e4cb, 32'h416ec771} /* (11, 18, 22) {real, imag} */,
  {32'hc096172e, 32'hbf7a0ce8} /* (11, 18, 21) {real, imag} */,
  {32'hc0aa9ec9, 32'hc0127052} /* (11, 18, 20) {real, imag} */,
  {32'h40511fb8, 32'h4101c46a} /* (11, 18, 19) {real, imag} */,
  {32'h4016c336, 32'h40d2912a} /* (11, 18, 18) {real, imag} */,
  {32'hbee32b10, 32'h3f403184} /* (11, 18, 17) {real, imag} */,
  {32'h40c91bbf, 32'hc0008d99} /* (11, 18, 16) {real, imag} */,
  {32'h40a72a7d, 32'h40ae96d4} /* (11, 18, 15) {real, imag} */,
  {32'h41161200, 32'h3f9329a8} /* (11, 18, 14) {real, imag} */,
  {32'hc085d857, 32'hc0225190} /* (11, 18, 13) {real, imag} */,
  {32'h40bc3dff, 32'hc102c698} /* (11, 18, 12) {real, imag} */,
  {32'hbfcfaf4e, 32'h415321ea} /* (11, 18, 11) {real, imag} */,
  {32'h3fe53542, 32'h4103e01d} /* (11, 18, 10) {real, imag} */,
  {32'h41675310, 32'hc109e770} /* (11, 18, 9) {real, imag} */,
  {32'h40a2ec5e, 32'hc0cba430} /* (11, 18, 8) {real, imag} */,
  {32'hc0d3383e, 32'hc11a77b4} /* (11, 18, 7) {real, imag} */,
  {32'hc0d1bbac, 32'h3ebb5a68} /* (11, 18, 6) {real, imag} */,
  {32'hc1662c31, 32'h3f919354} /* (11, 18, 5) {real, imag} */,
  {32'h3f840a18, 32'h408642f6} /* (11, 18, 4) {real, imag} */,
  {32'h40528106, 32'hc194c968} /* (11, 18, 3) {real, imag} */,
  {32'hc031da28, 32'h4110c175} /* (11, 18, 2) {real, imag} */,
  {32'h40e848c3, 32'hc0167220} /* (11, 18, 1) {real, imag} */,
  {32'h41514afe, 32'hc05587a1} /* (11, 18, 0) {real, imag} */,
  {32'h41343e73, 32'hc0a059f3} /* (11, 17, 31) {real, imag} */,
  {32'h413a262a, 32'h40f7b9dc} /* (11, 17, 30) {real, imag} */,
  {32'hc00114ec, 32'h41d7ee0b} /* (11, 17, 29) {real, imag} */,
  {32'hbfb5b466, 32'hc13bb9c6} /* (11, 17, 28) {real, imag} */,
  {32'hc1242da1, 32'hc0dbd6f7} /* (11, 17, 27) {real, imag} */,
  {32'h4023a5be, 32'hc101381d} /* (11, 17, 26) {real, imag} */,
  {32'h40bae8c9, 32'h41108f66} /* (11, 17, 25) {real, imag} */,
  {32'hc135e466, 32'h40002502} /* (11, 17, 24) {real, imag} */,
  {32'hc0bde303, 32'hc11b633c} /* (11, 17, 23) {real, imag} */,
  {32'h4039cb8c, 32'hbd4f5780} /* (11, 17, 22) {real, imag} */,
  {32'hc11d10da, 32'hc15a7120} /* (11, 17, 21) {real, imag} */,
  {32'hbfc2c04e, 32'hc044d05a} /* (11, 17, 20) {real, imag} */,
  {32'h3e1a82e0, 32'hbf16d48c} /* (11, 17, 19) {real, imag} */,
  {32'h4063bbf4, 32'h3e6f4148} /* (11, 17, 18) {real, imag} */,
  {32'hc092fedf, 32'hbe789620} /* (11, 17, 17) {real, imag} */,
  {32'hc0636ad5, 32'h407ada39} /* (11, 17, 16) {real, imag} */,
  {32'hc0921379, 32'h3fefada4} /* (11, 17, 15) {real, imag} */,
  {32'h3ef056e0, 32'h40508806} /* (11, 17, 14) {real, imag} */,
  {32'hc0e7738f, 32'hc0445273} /* (11, 17, 13) {real, imag} */,
  {32'h3f276afc, 32'h408c62cf} /* (11, 17, 12) {real, imag} */,
  {32'hc1031d84, 32'h41149b54} /* (11, 17, 11) {real, imag} */,
  {32'h400f1848, 32'hc07b34f6} /* (11, 17, 10) {real, imag} */,
  {32'hc11d0638, 32'hc0f5c0b8} /* (11, 17, 9) {real, imag} */,
  {32'hbed26b50, 32'h3fc7c3f0} /* (11, 17, 8) {real, imag} */,
  {32'hc18d3db1, 32'hc02cd390} /* (11, 17, 7) {real, imag} */,
  {32'hc1665f34, 32'h41516369} /* (11, 17, 6) {real, imag} */,
  {32'h411d743b, 32'hc1136edc} /* (11, 17, 5) {real, imag} */,
  {32'h4009089b, 32'hc1220a7e} /* (11, 17, 4) {real, imag} */,
  {32'h4101a71c, 32'hc149ecd6} /* (11, 17, 3) {real, imag} */,
  {32'h42330ab0, 32'h401f8278} /* (11, 17, 2) {real, imag} */,
  {32'hc12b4951, 32'h3f740dd8} /* (11, 17, 1) {real, imag} */,
  {32'hc0ec6194, 32'hc13abec6} /* (11, 17, 0) {real, imag} */,
  {32'hbf682f74, 32'h410c0ce1} /* (11, 16, 31) {real, imag} */,
  {32'hbee1d2b0, 32'h3f812298} /* (11, 16, 30) {real, imag} */,
  {32'hc108c33f, 32'hc09f1879} /* (11, 16, 29) {real, imag} */,
  {32'hc106645e, 32'h3f90a2b4} /* (11, 16, 28) {real, imag} */,
  {32'h3ecb6ee0, 32'h41986702} /* (11, 16, 27) {real, imag} */,
  {32'hc1156a8a, 32'hc0cc855a} /* (11, 16, 26) {real, imag} */,
  {32'hc0565d8e, 32'h3fde5e90} /* (11, 16, 25) {real, imag} */,
  {32'h40ec2580, 32'hc066c148} /* (11, 16, 24) {real, imag} */,
  {32'h41ba4087, 32'h40262b28} /* (11, 16, 23) {real, imag} */,
  {32'hbfedd836, 32'h3ffd8946} /* (11, 16, 22) {real, imag} */,
  {32'hc0860c07, 32'h40e50f32} /* (11, 16, 21) {real, imag} */,
  {32'hc08170e5, 32'hc06cbd0d} /* (11, 16, 20) {real, imag} */,
  {32'hc04706f7, 32'h405b7d1c} /* (11, 16, 19) {real, imag} */,
  {32'h3fab025d, 32'h3fa03ffc} /* (11, 16, 18) {real, imag} */,
  {32'h404390af, 32'hbec55a04} /* (11, 16, 17) {real, imag} */,
  {32'h3f87f9d0, 32'h3e550860} /* (11, 16, 16) {real, imag} */,
  {32'hc016980b, 32'hc04702e4} /* (11, 16, 15) {real, imag} */,
  {32'h3d994850, 32'hbf81fe10} /* (11, 16, 14) {real, imag} */,
  {32'h4104780a, 32'hc0414e58} /* (11, 16, 13) {real, imag} */,
  {32'h4008f120, 32'h40877be8} /* (11, 16, 12) {real, imag} */,
  {32'h4048eeb8, 32'hc0c5107e} /* (11, 16, 11) {real, imag} */,
  {32'hc0596a01, 32'hc0918e00} /* (11, 16, 10) {real, imag} */,
  {32'hbe82c040, 32'hc17d325e} /* (11, 16, 9) {real, imag} */,
  {32'h40da1e12, 32'hc13d4982} /* (11, 16, 8) {real, imag} */,
  {32'h41113664, 32'hc1831e6b} /* (11, 16, 7) {real, imag} */,
  {32'h3fa9a860, 32'h414d660f} /* (11, 16, 6) {real, imag} */,
  {32'hc15f1a57, 32'h40b3b07e} /* (11, 16, 5) {real, imag} */,
  {32'h410c168c, 32'hbf82c916} /* (11, 16, 4) {real, imag} */,
  {32'h41501995, 32'hbf811aac} /* (11, 16, 3) {real, imag} */,
  {32'h40a5a11d, 32'h4116f355} /* (11, 16, 2) {real, imag} */,
  {32'hc0f6c0c8, 32'hc0e47a25} /* (11, 16, 1) {real, imag} */,
  {32'h41afffc1, 32'h4093100d} /* (11, 16, 0) {real, imag} */,
  {32'h4194e408, 32'hc11ec813} /* (11, 15, 31) {real, imag} */,
  {32'hc15f2752, 32'h40172b16} /* (11, 15, 30) {real, imag} */,
  {32'hc14f3f4e, 32'h413ffa2c} /* (11, 15, 29) {real, imag} */,
  {32'hc05b131a, 32'hbf8c5964} /* (11, 15, 28) {real, imag} */,
  {32'hc021c112, 32'h418e0fa4} /* (11, 15, 27) {real, imag} */,
  {32'h3f85a1b2, 32'hc088e732} /* (11, 15, 26) {real, imag} */,
  {32'h4036fa50, 32'hc098e85d} /* (11, 15, 25) {real, imag} */,
  {32'hc19004b6, 32'h415775bd} /* (11, 15, 24) {real, imag} */,
  {32'hc0e59cf9, 32'hc01f7d77} /* (11, 15, 23) {real, imag} */,
  {32'h3f911922, 32'h4034a438} /* (11, 15, 22) {real, imag} */,
  {32'h40c72339, 32'h40f9ddd2} /* (11, 15, 21) {real, imag} */,
  {32'hc09578a2, 32'hc0418f44} /* (11, 15, 20) {real, imag} */,
  {32'h3fd436a0, 32'hc0d44423} /* (11, 15, 19) {real, imag} */,
  {32'h3fa8fd50, 32'hc098afbb} /* (11, 15, 18) {real, imag} */,
  {32'h3e81f770, 32'hbf951334} /* (11, 15, 17) {real, imag} */,
  {32'hc06867ae, 32'h3faa93a4} /* (11, 15, 16) {real, imag} */,
  {32'hc00d114a, 32'hbf757828} /* (11, 15, 15) {real, imag} */,
  {32'h3f7d8b60, 32'h40182108} /* (11, 15, 14) {real, imag} */,
  {32'hc0e830ba, 32'hbfd22b74} /* (11, 15, 13) {real, imag} */,
  {32'h4006b81b, 32'hbf9c7be0} /* (11, 15, 12) {real, imag} */,
  {32'h412971cc, 32'hc128a20f} /* (11, 15, 11) {real, imag} */,
  {32'h408bfcee, 32'hc091c0d0} /* (11, 15, 10) {real, imag} */,
  {32'hc0aca517, 32'h3f28b254} /* (11, 15, 9) {real, imag} */,
  {32'hbf4f1e80, 32'h412f0555} /* (11, 15, 8) {real, imag} */,
  {32'h40e03618, 32'hc0b9e03f} /* (11, 15, 7) {real, imag} */,
  {32'hc0ca5a66, 32'h411e1301} /* (11, 15, 6) {real, imag} */,
  {32'h414dd694, 32'h4128419e} /* (11, 15, 5) {real, imag} */,
  {32'h401b3046, 32'hc17ac85c} /* (11, 15, 4) {real, imag} */,
  {32'hbea8d7a0, 32'h4190092a} /* (11, 15, 3) {real, imag} */,
  {32'h3fe00b10, 32'hbe83f764} /* (11, 15, 2) {real, imag} */,
  {32'h411bf155, 32'h40f32162} /* (11, 15, 1) {real, imag} */,
  {32'h41021168, 32'hbfbae174} /* (11, 15, 0) {real, imag} */,
  {32'hc012086c, 32'hc19e9a11} /* (11, 14, 31) {real, imag} */,
  {32'hc1558cac, 32'h4161794d} /* (11, 14, 30) {real, imag} */,
  {32'h411205a3, 32'hc18ea8be} /* (11, 14, 29) {real, imag} */,
  {32'hc0fe1ef7, 32'h410e5f8e} /* (11, 14, 28) {real, imag} */,
  {32'h407e1336, 32'hbea481a0} /* (11, 14, 27) {real, imag} */,
  {32'hc0d3aca6, 32'h3f9bc8aa} /* (11, 14, 26) {real, imag} */,
  {32'hbecced50, 32'h3f4859cc} /* (11, 14, 25) {real, imag} */,
  {32'hc1206836, 32'hc1734532} /* (11, 14, 24) {real, imag} */,
  {32'h41219a8e, 32'h40c7afca} /* (11, 14, 23) {real, imag} */,
  {32'hc1a09585, 32'h3efe9348} /* (11, 14, 22) {real, imag} */,
  {32'hbf1ee46c, 32'h3f40bf80} /* (11, 14, 21) {real, imag} */,
  {32'hbf4bae6c, 32'hbe9d2928} /* (11, 14, 20) {real, imag} */,
  {32'h405f3f39, 32'hc09c6474} /* (11, 14, 19) {real, imag} */,
  {32'h410695bc, 32'h408d2934} /* (11, 14, 18) {real, imag} */,
  {32'h3f9e7908, 32'h400565ec} /* (11, 14, 17) {real, imag} */,
  {32'h40ae5c06, 32'hc0ec268f} /* (11, 14, 16) {real, imag} */,
  {32'hc01d8454, 32'h403f09f4} /* (11, 14, 15) {real, imag} */,
  {32'h400128be, 32'hc009a94f} /* (11, 14, 14) {real, imag} */,
  {32'h40cc4440, 32'h4046ae80} /* (11, 14, 13) {real, imag} */,
  {32'h3f1a0600, 32'hc062efff} /* (11, 14, 12) {real, imag} */,
  {32'hbf3f6238, 32'h40ff275c} /* (11, 14, 11) {real, imag} */,
  {32'hc0c7885d, 32'h3fba4152} /* (11, 14, 10) {real, imag} */,
  {32'hc098407b, 32'hc018e8ac} /* (11, 14, 9) {real, imag} */,
  {32'h3f5f6558, 32'hc0a199ac} /* (11, 14, 8) {real, imag} */,
  {32'hc1302766, 32'hbfd68fb6} /* (11, 14, 7) {real, imag} */,
  {32'hbe82fdc0, 32'hc0d2c890} /* (11, 14, 6) {real, imag} */,
  {32'h3fcb1a33, 32'h41999508} /* (11, 14, 5) {real, imag} */,
  {32'h3f897b2c, 32'hc03c6dd6} /* (11, 14, 4) {real, imag} */,
  {32'h3fb1e486, 32'hc17c81dd} /* (11, 14, 3) {real, imag} */,
  {32'h413416b8, 32'h4087aeda} /* (11, 14, 2) {real, imag} */,
  {32'hc1925b52, 32'h41cd5faf} /* (11, 14, 1) {real, imag} */,
  {32'hc09ef432, 32'hc1969bf8} /* (11, 14, 0) {real, imag} */,
  {32'h411793d8, 32'hc18afc30} /* (11, 13, 31) {real, imag} */,
  {32'h4100580e, 32'h41c3c4f2} /* (11, 13, 30) {real, imag} */,
  {32'h40dd832f, 32'h418d89dc} /* (11, 13, 29) {real, imag} */,
  {32'hc0ae8966, 32'hbee9c6c0} /* (11, 13, 28) {real, imag} */,
  {32'hc12a86c6, 32'h4163f670} /* (11, 13, 27) {real, imag} */,
  {32'h4125c261, 32'h4085b40e} /* (11, 13, 26) {real, imag} */,
  {32'h4198d9d1, 32'hc0f4b6f8} /* (11, 13, 25) {real, imag} */,
  {32'h4087ed93, 32'h3f9a9472} /* (11, 13, 24) {real, imag} */,
  {32'h4173abee, 32'h4135fa88} /* (11, 13, 23) {real, imag} */,
  {32'h4119a15b, 32'hc16f5bf6} /* (11, 13, 22) {real, imag} */,
  {32'hbf07e278, 32'hbfd79df4} /* (11, 13, 21) {real, imag} */,
  {32'h405abd53, 32'h40f383b8} /* (11, 13, 20) {real, imag} */,
  {32'hbfe37404, 32'hc09490f4} /* (11, 13, 19) {real, imag} */,
  {32'h3dd33eb0, 32'h411883fa} /* (11, 13, 18) {real, imag} */,
  {32'hc09d3cd6, 32'h3fa671c4} /* (11, 13, 17) {real, imag} */,
  {32'hc01080bc, 32'hbffd381c} /* (11, 13, 16) {real, imag} */,
  {32'hc012bbf0, 32'hc04e8cea} /* (11, 13, 15) {real, imag} */,
  {32'h3ff44023, 32'hbffa771c} /* (11, 13, 14) {real, imag} */,
  {32'hbf931034, 32'hc0976798} /* (11, 13, 13) {real, imag} */,
  {32'h40a46724, 32'hc09b0c20} /* (11, 13, 12) {real, imag} */,
  {32'h40a84d23, 32'hc123d8f8} /* (11, 13, 11) {real, imag} */,
  {32'h4024010b, 32'h407d64ba} /* (11, 13, 10) {real, imag} */,
  {32'hc08cd97b, 32'hc11da0a0} /* (11, 13, 9) {real, imag} */,
  {32'h41167e56, 32'hc0a04b60} /* (11, 13, 8) {real, imag} */,
  {32'hbfb49970, 32'h408de706} /* (11, 13, 7) {real, imag} */,
  {32'h417dd471, 32'h3e9d5600} /* (11, 13, 6) {real, imag} */,
  {32'h405a364a, 32'hc1ada590} /* (11, 13, 5) {real, imag} */,
  {32'h41299059, 32'h41233ece} /* (11, 13, 4) {real, imag} */,
  {32'hc1a8a4c5, 32'hbfe9e488} /* (11, 13, 3) {real, imag} */,
  {32'hc112da72, 32'h4181f162} /* (11, 13, 2) {real, imag} */,
  {32'hc137c814, 32'h4081df8a} /* (11, 13, 1) {real, imag} */,
  {32'h41a97eaa, 32'h414cad16} /* (11, 13, 0) {real, imag} */,
  {32'h4199a112, 32'h41d3436e} /* (11, 12, 31) {real, imag} */,
  {32'hc2060716, 32'hc02dbaa0} /* (11, 12, 30) {real, imag} */,
  {32'hbeccf630, 32'h3ff00f98} /* (11, 12, 29) {real, imag} */,
  {32'h4196240a, 32'h40827be2} /* (11, 12, 28) {real, imag} */,
  {32'h415deb08, 32'hc16587f5} /* (11, 12, 27) {real, imag} */,
  {32'hc193b0b7, 32'h41f01924} /* (11, 12, 26) {real, imag} */,
  {32'hc1734bcc, 32'h415b8c38} /* (11, 12, 25) {real, imag} */,
  {32'h405dbc4e, 32'h41afd2a6} /* (11, 12, 24) {real, imag} */,
  {32'hc0c9fe91, 32'hc0ca5012} /* (11, 12, 23) {real, imag} */,
  {32'hc13652ac, 32'hc1703060} /* (11, 12, 22) {real, imag} */,
  {32'h3fe52628, 32'hc1738bee} /* (11, 12, 21) {real, imag} */,
  {32'hbfec99d4, 32'hc16e7af4} /* (11, 12, 20) {real, imag} */,
  {32'hc1012023, 32'h411d92aa} /* (11, 12, 19) {real, imag} */,
  {32'h41143300, 32'hc14c125e} /* (11, 12, 18) {real, imag} */,
  {32'hc07b767a, 32'hc1081dfe} /* (11, 12, 17) {real, imag} */,
  {32'hbfc90b2c, 32'hbeb47e80} /* (11, 12, 16) {real, imag} */,
  {32'hc031940a, 32'hc0f36d5c} /* (11, 12, 15) {real, imag} */,
  {32'h3ef6b490, 32'h4095b15b} /* (11, 12, 14) {real, imag} */,
  {32'h406f9a17, 32'hc14d5d62} /* (11, 12, 13) {real, imag} */,
  {32'hbe16cea0, 32'hc0655152} /* (11, 12, 12) {real, imag} */,
  {32'hc09b8ade, 32'hc07a1b20} /* (11, 12, 11) {real, imag} */,
  {32'h4094553f, 32'h3eaf81d0} /* (11, 12, 10) {real, imag} */,
  {32'h40547982, 32'h408506f4} /* (11, 12, 9) {real, imag} */,
  {32'hc1465158, 32'hc12f6e2c} /* (11, 12, 8) {real, imag} */,
  {32'h41b82fea, 32'hc0705898} /* (11, 12, 7) {real, imag} */,
  {32'h40bdd0b3, 32'hc0070c40} /* (11, 12, 6) {real, imag} */,
  {32'hc12c3b6c, 32'hc1a9df1e} /* (11, 12, 5) {real, imag} */,
  {32'h40b6227a, 32'h401de9f0} /* (11, 12, 4) {real, imag} */,
  {32'hc1711350, 32'h40ed6226} /* (11, 12, 3) {real, imag} */,
  {32'hc1cf5b7e, 32'h41eb9ed2} /* (11, 12, 2) {real, imag} */,
  {32'hc1e352b8, 32'hc1c79682} /* (11, 12, 1) {real, imag} */,
  {32'h403ad12a, 32'hc19dfbea} /* (11, 12, 0) {real, imag} */,
  {32'hc26e1b02, 32'h415d07af} /* (11, 11, 31) {real, imag} */,
  {32'hc1cb08c5, 32'h4258e962} /* (11, 11, 30) {real, imag} */,
  {32'hc1e384b6, 32'h4112c29c} /* (11, 11, 29) {real, imag} */,
  {32'hc0afa5e0, 32'hc0bcfe08} /* (11, 11, 28) {real, imag} */,
  {32'hc10512db, 32'hc199862b} /* (11, 11, 27) {real, imag} */,
  {32'h416f1dc9, 32'hc1cc3af3} /* (11, 11, 26) {real, imag} */,
  {32'hc1b173f7, 32'hc13b9ad5} /* (11, 11, 25) {real, imag} */,
  {32'h418bc169, 32'hc17a9df0} /* (11, 11, 24) {real, imag} */,
  {32'hc09fb686, 32'hbfa88f48} /* (11, 11, 23) {real, imag} */,
  {32'h414e2a5f, 32'hc101b3f7} /* (11, 11, 22) {real, imag} */,
  {32'h409389d6, 32'hc0efe075} /* (11, 11, 21) {real, imag} */,
  {32'hc0ca156c, 32'hc1a1f990} /* (11, 11, 20) {real, imag} */,
  {32'hc0c2e03c, 32'hc0964b63} /* (11, 11, 19) {real, imag} */,
  {32'hc15851dd, 32'hc11fd398} /* (11, 11, 18) {real, imag} */,
  {32'hbffcb548, 32'h411e088a} /* (11, 11, 17) {real, imag} */,
  {32'hc0482860, 32'hc071dd88} /* (11, 11, 16) {real, imag} */,
  {32'h3faaaee8, 32'h40848314} /* (11, 11, 15) {real, imag} */,
  {32'hc0635714, 32'hc10fc016} /* (11, 11, 14) {real, imag} */,
  {32'hc074d7b8, 32'hc04cbfb6} /* (11, 11, 13) {real, imag} */,
  {32'h411387b0, 32'h40844574} /* (11, 11, 12) {real, imag} */,
  {32'hbf1f04bc, 32'h419e40c1} /* (11, 11, 11) {real, imag} */,
  {32'h40658cac, 32'hc11e19ed} /* (11, 11, 10) {real, imag} */,
  {32'hc144e6c5, 32'hc0f28020} /* (11, 11, 9) {real, imag} */,
  {32'h40760da8, 32'h41039cc8} /* (11, 11, 8) {real, imag} */,
  {32'hbf686fa0, 32'hc0545900} /* (11, 11, 7) {real, imag} */,
  {32'hc0d73f7a, 32'hc19bb105} /* (11, 11, 6) {real, imag} */,
  {32'hc0929900, 32'hc0adf753} /* (11, 11, 5) {real, imag} */,
  {32'hc236f08a, 32'h423baf8d} /* (11, 11, 4) {real, imag} */,
  {32'hc2200a65, 32'h40d41a0b} /* (11, 11, 3) {real, imag} */,
  {32'hc15926f6, 32'h3fc2df80} /* (11, 11, 2) {real, imag} */,
  {32'hbf9183b0, 32'hc1379aa9} /* (11, 11, 1) {real, imag} */,
  {32'hc1801f6c, 32'hc2030c34} /* (11, 11, 0) {real, imag} */,
  {32'hc0e140c0, 32'h400fb470} /* (11, 10, 31) {real, imag} */,
  {32'hc14c4e18, 32'hc10effc3} /* (11, 10, 30) {real, imag} */,
  {32'h4206a8ec, 32'hc1adadb9} /* (11, 10, 29) {real, imag} */,
  {32'h40d2f94e, 32'h41f01014} /* (11, 10, 28) {real, imag} */,
  {32'h41e3a6be, 32'hc14a8cd0} /* (11, 10, 27) {real, imag} */,
  {32'hc1162522, 32'hc1e8c106} /* (11, 10, 26) {real, imag} */,
  {32'hbfdec9b4, 32'h42537fda} /* (11, 10, 25) {real, imag} */,
  {32'h4261726b, 32'hc239743b} /* (11, 10, 24) {real, imag} */,
  {32'hc21c60c6, 32'h41a540f6} /* (11, 10, 23) {real, imag} */,
  {32'hc13b4282, 32'hbeb72c80} /* (11, 10, 22) {real, imag} */,
  {32'h40eb417a, 32'h40575a67} /* (11, 10, 21) {real, imag} */,
  {32'hc1611595, 32'h40b28a90} /* (11, 10, 20) {real, imag} */,
  {32'h405d9266, 32'hc09311da} /* (11, 10, 19) {real, imag} */,
  {32'hc117e1c5, 32'h411b8bae} /* (11, 10, 18) {real, imag} */,
  {32'h40c51850, 32'hbf6358b8} /* (11, 10, 17) {real, imag} */,
  {32'hbf3c4c78, 32'hc0bdb918} /* (11, 10, 16) {real, imag} */,
  {32'hbf193ec0, 32'h4002aefe} /* (11, 10, 15) {real, imag} */,
  {32'h417482a3, 32'h40bf1ca4} /* (11, 10, 14) {real, imag} */,
  {32'hc17ef62e, 32'hc0e0cfb6} /* (11, 10, 13) {real, imag} */,
  {32'h418f3e36, 32'h40665739} /* (11, 10, 12) {real, imag} */,
  {32'h4088c586, 32'hc000a277} /* (11, 10, 11) {real, imag} */,
  {32'h4139e55a, 32'h41af9005} /* (11, 10, 10) {real, imag} */,
  {32'hc1b49ab5, 32'hc220f379} /* (11, 10, 9) {real, imag} */,
  {32'h416151bc, 32'hc1d7f7be} /* (11, 10, 8) {real, imag} */,
  {32'h40f94dbd, 32'hbf87a480} /* (11, 10, 7) {real, imag} */,
  {32'h4121e4ee, 32'hc120e135} /* (11, 10, 6) {real, imag} */,
  {32'hc1674d95, 32'hc19242f2} /* (11, 10, 5) {real, imag} */,
  {32'hc1878d5c, 32'h41961620} /* (11, 10, 4) {real, imag} */,
  {32'hc145f5e8, 32'h41fd2417} /* (11, 10, 3) {real, imag} */,
  {32'hc1dc5184, 32'hc136f4b1} /* (11, 10, 2) {real, imag} */,
  {32'hc26343a7, 32'h4211863f} /* (11, 10, 1) {real, imag} */,
  {32'hc15440fe, 32'h42886924} /* (11, 10, 0) {real, imag} */,
  {32'hc2186deb, 32'hc1032d98} /* (11, 9, 31) {real, imag} */,
  {32'h42140f38, 32'h420ce794} /* (11, 9, 30) {real, imag} */,
  {32'hc2079940, 32'h4068c1e0} /* (11, 9, 29) {real, imag} */,
  {32'hc24c0964, 32'h40fd98a6} /* (11, 9, 28) {real, imag} */,
  {32'hc1cdff6b, 32'h41ed9620} /* (11, 9, 27) {real, imag} */,
  {32'hbfa9d7f8, 32'hc0e895da} /* (11, 9, 26) {real, imag} */,
  {32'h41c246c5, 32'h42037e88} /* (11, 9, 25) {real, imag} */,
  {32'hc1fa1077, 32'h41d373da} /* (11, 9, 24) {real, imag} */,
  {32'hc1befc44, 32'h41864761} /* (11, 9, 23) {real, imag} */,
  {32'hc1ff6f39, 32'hc1c72342} /* (11, 9, 22) {real, imag} */,
  {32'h411172ff, 32'hc105e283} /* (11, 9, 21) {real, imag} */,
  {32'hc09bb684, 32'hc0dfd809} /* (11, 9, 20) {real, imag} */,
  {32'h40be6e30, 32'h40d35b42} /* (11, 9, 19) {real, imag} */,
  {32'hc08a5c45, 32'h3fabfd52} /* (11, 9, 18) {real, imag} */,
  {32'hc0b03b6a, 32'hc1accc32} /* (11, 9, 17) {real, imag} */,
  {32'h409b815c, 32'hc1122f52} /* (11, 9, 16) {real, imag} */,
  {32'hc0f37ff2, 32'hc003b3b4} /* (11, 9, 15) {real, imag} */,
  {32'hc118af88, 32'h405e0d89} /* (11, 9, 14) {real, imag} */,
  {32'h40874724, 32'h413df535} /* (11, 9, 13) {real, imag} */,
  {32'h4114a55e, 32'h417df5fe} /* (11, 9, 12) {real, imag} */,
  {32'hc18ec6f6, 32'h4096d102} /* (11, 9, 11) {real, imag} */,
  {32'hc181cb4b, 32'hbf8b9448} /* (11, 9, 10) {real, imag} */,
  {32'hc1a132d8, 32'hc01b0978} /* (11, 9, 9) {real, imag} */,
  {32'h41d2f45f, 32'h40b19656} /* (11, 9, 8) {real, imag} */,
  {32'hc01dc0f0, 32'h4103c63c} /* (11, 9, 7) {real, imag} */,
  {32'h41052bb9, 32'h41ea3038} /* (11, 9, 6) {real, imag} */,
  {32'h41d87a97, 32'hc15d5d49} /* (11, 9, 5) {real, imag} */,
  {32'hbf8a6940, 32'h41aed19c} /* (11, 9, 4) {real, imag} */,
  {32'h409c14ae, 32'hc22e87a6} /* (11, 9, 3) {real, imag} */,
  {32'hbfc74650, 32'hc221ac62} /* (11, 9, 2) {real, imag} */,
  {32'h42af45ac, 32'h40d7b8b5} /* (11, 9, 1) {real, imag} */,
  {32'h4245c822, 32'hc258ca22} /* (11, 9, 0) {real, imag} */,
  {32'hc1006968, 32'hc1f117ee} /* (11, 8, 31) {real, imag} */,
  {32'hc1ea198a, 32'h4185e530} /* (11, 8, 30) {real, imag} */,
  {32'hc1a4fa56, 32'h417e8fb5} /* (11, 8, 29) {real, imag} */,
  {32'h42046e3e, 32'hc211a32f} /* (11, 8, 28) {real, imag} */,
  {32'h402d7894, 32'hc202be21} /* (11, 8, 27) {real, imag} */,
  {32'h41071a98, 32'hc0f6709e} /* (11, 8, 26) {real, imag} */,
  {32'hc27fa21e, 32'hc1a8d3bc} /* (11, 8, 25) {real, imag} */,
  {32'hc1a1e6b2, 32'hc1b81ecf} /* (11, 8, 24) {real, imag} */,
  {32'hc0a41e9e, 32'h41bbdbc0} /* (11, 8, 23) {real, imag} */,
  {32'h421e2de9, 32'h419fb6ca} /* (11, 8, 22) {real, imag} */,
  {32'h42174cb0, 32'h3f8b287c} /* (11, 8, 21) {real, imag} */,
  {32'hbff5bad6, 32'hc1368e69} /* (11, 8, 20) {real, imag} */,
  {32'hbf529f18, 32'h405a31c8} /* (11, 8, 19) {real, imag} */,
  {32'h4155d046, 32'hc134d61c} /* (11, 8, 18) {real, imag} */,
  {32'hc0f896a8, 32'hc0e7941c} /* (11, 8, 17) {real, imag} */,
  {32'h40b2782d, 32'hbe6f9600} /* (11, 8, 16) {real, imag} */,
  {32'hc0f8c7f2, 32'h407fd7a0} /* (11, 8, 15) {real, imag} */,
  {32'hc0dd4c60, 32'h40662dc5} /* (11, 8, 14) {real, imag} */,
  {32'h4122bb5a, 32'h4201e31a} /* (11, 8, 13) {real, imag} */,
  {32'hc047c34b, 32'h412f483f} /* (11, 8, 12) {real, imag} */,
  {32'hc05e6608, 32'hc1831428} /* (11, 8, 11) {real, imag} */,
  {32'hc19739e6, 32'hc162f253} /* (11, 8, 10) {real, imag} */,
  {32'hc187f1f8, 32'hc0ef1886} /* (11, 8, 9) {real, imag} */,
  {32'h4221fe79, 32'hc043c548} /* (11, 8, 8) {real, imag} */,
  {32'h4228c906, 32'h401ca0f4} /* (11, 8, 7) {real, imag} */,
  {32'hc256e56c, 32'h41d481d4} /* (11, 8, 6) {real, imag} */,
  {32'hc1af5c64, 32'h4217a92d} /* (11, 8, 5) {real, imag} */,
  {32'hc2188158, 32'h42018e71} /* (11, 8, 4) {real, imag} */,
  {32'h41abb176, 32'h3f417310} /* (11, 8, 3) {real, imag} */,
  {32'hc1ddfc02, 32'h3e8323e0} /* (11, 8, 2) {real, imag} */,
  {32'h3fb5bdb4, 32'hc1a8b976} /* (11, 8, 1) {real, imag} */,
  {32'h418217e1, 32'h41979cdc} /* (11, 8, 0) {real, imag} */,
  {32'h42a40da7, 32'hc1aa4c24} /* (11, 7, 31) {real, imag} */,
  {32'hc23086ba, 32'hc085a918} /* (11, 7, 30) {real, imag} */,
  {32'h425acc6d, 32'h429b9474} /* (11, 7, 29) {real, imag} */,
  {32'h3f858b90, 32'hc1be81e5} /* (11, 7, 28) {real, imag} */,
  {32'hc2693ebd, 32'h415a3f74} /* (11, 7, 27) {real, imag} */,
  {32'hc1bd4545, 32'hc1a1f724} /* (11, 7, 26) {real, imag} */,
  {32'hc0d793f2, 32'hc1686abe} /* (11, 7, 25) {real, imag} */,
  {32'h41f58f4d, 32'hc0b3c5de} /* (11, 7, 24) {real, imag} */,
  {32'hc20d35f2, 32'hc16b32ec} /* (11, 7, 23) {real, imag} */,
  {32'h4026f268, 32'h4229cd6b} /* (11, 7, 22) {real, imag} */,
  {32'hc1cbe38b, 32'hc00590d8} /* (11, 7, 21) {real, imag} */,
  {32'h421af264, 32'h415a7460} /* (11, 7, 20) {real, imag} */,
  {32'hc0fcce48, 32'h41cee1a9} /* (11, 7, 19) {real, imag} */,
  {32'hc026d988, 32'hc0df8708} /* (11, 7, 18) {real, imag} */,
  {32'h4089d22e, 32'h405c8c70} /* (11, 7, 17) {real, imag} */,
  {32'hc16ab8ea, 32'hbfb349a8} /* (11, 7, 16) {real, imag} */,
  {32'hc11aae47, 32'h4162aec2} /* (11, 7, 15) {real, imag} */,
  {32'h40aac27c, 32'hc120d204} /* (11, 7, 14) {real, imag} */,
  {32'hc16f1ffc, 32'hc19f928f} /* (11, 7, 13) {real, imag} */,
  {32'hbffd58b0, 32'hbf1109d0} /* (11, 7, 12) {real, imag} */,
  {32'h41d96dad, 32'h419ff09b} /* (11, 7, 11) {real, imag} */,
  {32'hc0db4f9c, 32'hc1422949} /* (11, 7, 10) {real, imag} */,
  {32'h413702c0, 32'hbb428000} /* (11, 7, 9) {real, imag} */,
  {32'h4219ccc0, 32'h4128c78d} /* (11, 7, 8) {real, imag} */,
  {32'h41aa09e0, 32'h42366414} /* (11, 7, 7) {real, imag} */,
  {32'h428d23f2, 32'hbffcae28} /* (11, 7, 6) {real, imag} */,
  {32'hc2152033, 32'hc2a3ee94} /* (11, 7, 5) {real, imag} */,
  {32'h420cbf1c, 32'h4196921d} /* (11, 7, 4) {real, imag} */,
  {32'hc1cef6be, 32'hc297b1fe} /* (11, 7, 3) {real, imag} */,
  {32'hbf11ad60, 32'h40bfe878} /* (11, 7, 2) {real, imag} */,
  {32'h42b82c73, 32'hc1bc394c} /* (11, 7, 1) {real, imag} */,
  {32'hc28dc3a4, 32'h41e56038} /* (11, 7, 0) {real, imag} */,
  {32'h4304ab5e, 32'h4232539e} /* (11, 6, 31) {real, imag} */,
  {32'hc0b11703, 32'h41ff6ce5} /* (11, 6, 30) {real, imag} */,
  {32'hc26b2781, 32'hc2476f6c} /* (11, 6, 29) {real, imag} */,
  {32'h420f113a, 32'hc18bdce9} /* (11, 6, 28) {real, imag} */,
  {32'hc240c1b7, 32'h41a57ab8} /* (11, 6, 27) {real, imag} */,
  {32'hc213d7e7, 32'hc19b360c} /* (11, 6, 26) {real, imag} */,
  {32'hc0f35ee8, 32'hc1a33882} /* (11, 6, 25) {real, imag} */,
  {32'hc25ac73c, 32'h4218c834} /* (11, 6, 24) {real, imag} */,
  {32'h4136a360, 32'hc0beb5c4} /* (11, 6, 23) {real, imag} */,
  {32'h402537a8, 32'hc1fe6acb} /* (11, 6, 22) {real, imag} */,
  {32'hc1068937, 32'h41715a56} /* (11, 6, 21) {real, imag} */,
  {32'h418b7374, 32'h41e94fad} /* (11, 6, 20) {real, imag} */,
  {32'hc17016ce, 32'hc180c6c6} /* (11, 6, 19) {real, imag} */,
  {32'h41743b85, 32'h414c541a} /* (11, 6, 18) {real, imag} */,
  {32'h41111bc2, 32'hc16b9b59} /* (11, 6, 17) {real, imag} */,
  {32'h414cc1c0, 32'h41631c5b} /* (11, 6, 16) {real, imag} */,
  {32'h40875fdc, 32'hc0de9bde} /* (11, 6, 15) {real, imag} */,
  {32'hc0afad8e, 32'h40ee33ac} /* (11, 6, 14) {real, imag} */,
  {32'hc0ef6664, 32'h40832d4a} /* (11, 6, 13) {real, imag} */,
  {32'hbf586ac0, 32'h41aa7f3f} /* (11, 6, 12) {real, imag} */,
  {32'h40f93b92, 32'h41cf3e61} /* (11, 6, 11) {real, imag} */,
  {32'hbfe84b10, 32'h426821f2} /* (11, 6, 10) {real, imag} */,
  {32'h421d3227, 32'h41e1b873} /* (11, 6, 9) {real, imag} */,
  {32'hc217cde2, 32'hc09b5ab0} /* (11, 6, 8) {real, imag} */,
  {32'hc201cb5a, 32'hc188cfb0} /* (11, 6, 7) {real, imag} */,
  {32'hc20b940b, 32'h423586f2} /* (11, 6, 6) {real, imag} */,
  {32'h420ce183, 32'hc1860b6e} /* (11, 6, 5) {real, imag} */,
  {32'h42515386, 32'hc2236d02} /* (11, 6, 4) {real, imag} */,
  {32'h42159dfb, 32'h4108d300} /* (11, 6, 3) {real, imag} */,
  {32'hc0de3ab1, 32'h421ede22} /* (11, 6, 2) {real, imag} */,
  {32'h423bdffe, 32'h4198627c} /* (11, 6, 1) {real, imag} */,
  {32'hc2af1353, 32'hc179ab3d} /* (11, 6, 0) {real, imag} */,
  {32'hc275a018, 32'h42aaa6d1} /* (11, 5, 31) {real, imag} */,
  {32'h42247aaa, 32'h425b099c} /* (11, 5, 30) {real, imag} */,
  {32'h40e54b19, 32'h3f818d40} /* (11, 5, 29) {real, imag} */,
  {32'h41baaa71, 32'hc28305c6} /* (11, 5, 28) {real, imag} */,
  {32'h421dc434, 32'hc1c85b74} /* (11, 5, 27) {real, imag} */,
  {32'hc1430dab, 32'h41333dd4} /* (11, 5, 26) {real, imag} */,
  {32'hc1bae1f4, 32'h421f0f18} /* (11, 5, 25) {real, imag} */,
  {32'h40f68bec, 32'h40de6c38} /* (11, 5, 24) {real, imag} */,
  {32'h3f8bb1a8, 32'hc1d2a379} /* (11, 5, 23) {real, imag} */,
  {32'hc2043bfe, 32'h40b00560} /* (11, 5, 22) {real, imag} */,
  {32'h4168662a, 32'hc1adbae8} /* (11, 5, 21) {real, imag} */,
  {32'h41254564, 32'h41376e85} /* (11, 5, 20) {real, imag} */,
  {32'hc0cc3ff5, 32'h41e87142} /* (11, 5, 19) {real, imag} */,
  {32'hc10d12e2, 32'hc0dc80b6} /* (11, 5, 18) {real, imag} */,
  {32'hbfc9df90, 32'h40334648} /* (11, 5, 17) {real, imag} */,
  {32'h41852eaf, 32'hbf44f470} /* (11, 5, 16) {real, imag} */,
  {32'h41a08d79, 32'hc0e05b2c} /* (11, 5, 15) {real, imag} */,
  {32'hc1639f9e, 32'h404e1174} /* (11, 5, 14) {real, imag} */,
  {32'hc1ad1de9, 32'h413533c4} /* (11, 5, 13) {real, imag} */,
  {32'hc2096f3c, 32'hc0408c14} /* (11, 5, 12) {real, imag} */,
  {32'h41ae3677, 32'h42034152} /* (11, 5, 11) {real, imag} */,
  {32'hc0901cb4, 32'h41c3e162} /* (11, 5, 10) {real, imag} */,
  {32'h41a090fe, 32'hc22c9ffc} /* (11, 5, 9) {real, imag} */,
  {32'h4236d746, 32'h41818c00} /* (11, 5, 8) {real, imag} */,
  {32'hc22786e4, 32'hc20ff730} /* (11, 5, 7) {real, imag} */,
  {32'hc190b870, 32'hc1807ca4} /* (11, 5, 6) {real, imag} */,
  {32'h418b2413, 32'h427cee78} /* (11, 5, 5) {real, imag} */,
  {32'hc147e23a, 32'hc27ac2eb} /* (11, 5, 4) {real, imag} */,
  {32'hc03f0482, 32'hc25565ba} /* (11, 5, 3) {real, imag} */,
  {32'h425776ec, 32'hc1c023bc} /* (11, 5, 2) {real, imag} */,
  {32'hc31f86ac, 32'hc25b224e} /* (11, 5, 1) {real, imag} */,
  {32'hc264a594, 32'h41b3e218} /* (11, 5, 0) {real, imag} */,
  {32'h41432874, 32'h41b5a6c0} /* (11, 4, 31) {real, imag} */,
  {32'h40040bc0, 32'hc2988b0b} /* (11, 4, 30) {real, imag} */,
  {32'hc0c8a510, 32'h4231dba8} /* (11, 4, 29) {real, imag} */,
  {32'h414260b3, 32'hc232b71a} /* (11, 4, 28) {real, imag} */,
  {32'hc2cae5d3, 32'h424729ce} /* (11, 4, 27) {real, imag} */,
  {32'h422f2550, 32'hc1f67002} /* (11, 4, 26) {real, imag} */,
  {32'hc134f928, 32'h42ae5f8e} /* (11, 4, 25) {real, imag} */,
  {32'h40ef22ec, 32'h4121b6a3} /* (11, 4, 24) {real, imag} */,
  {32'hc1d03338, 32'hc173fe6c} /* (11, 4, 23) {real, imag} */,
  {32'hc23900a9, 32'h402fd0d8} /* (11, 4, 22) {real, imag} */,
  {32'hbf69e2b0, 32'h416d7c78} /* (11, 4, 21) {real, imag} */,
  {32'h418fe336, 32'h41a89796} /* (11, 4, 20) {real, imag} */,
  {32'h41865d81, 32'hc124f8d9} /* (11, 4, 19) {real, imag} */,
  {32'h3fc71a30, 32'hc188727b} /* (11, 4, 18) {real, imag} */,
  {32'hbddfe200, 32'hc1b27574} /* (11, 4, 17) {real, imag} */,
  {32'hc036c8e0, 32'h41934738} /* (11, 4, 16) {real, imag} */,
  {32'h418ae73a, 32'h400262b4} /* (11, 4, 15) {real, imag} */,
  {32'hbfef0e50, 32'h4156cf6e} /* (11, 4, 14) {real, imag} */,
  {32'hc1ea1551, 32'hc092dab2} /* (11, 4, 13) {real, imag} */,
  {32'hc1ee18f2, 32'h41c2f77a} /* (11, 4, 12) {real, imag} */,
  {32'hc1f6ada2, 32'h40bfea69} /* (11, 4, 11) {real, imag} */,
  {32'h4012beb0, 32'hc1f599f7} /* (11, 4, 10) {real, imag} */,
  {32'hc012e9bc, 32'hc2621e07} /* (11, 4, 9) {real, imag} */,
  {32'hc0b12c7c, 32'hc195c978} /* (11, 4, 8) {real, imag} */,
  {32'h42a31da5, 32'hc23af418} /* (11, 4, 7) {real, imag} */,
  {32'hc2986c66, 32'h42484eef} /* (11, 4, 6) {real, imag} */,
  {32'hc25f96ba, 32'h41ec30ec} /* (11, 4, 5) {real, imag} */,
  {32'h4191779c, 32'h4235043c} /* (11, 4, 4) {real, imag} */,
  {32'h42a8b297, 32'hc1f479b8} /* (11, 4, 3) {real, imag} */,
  {32'hc2b50fb4, 32'hc2ef4639} /* (11, 4, 2) {real, imag} */,
  {32'h42f582cc, 32'h3fe1f2c8} /* (11, 4, 1) {real, imag} */,
  {32'h4218446d, 32'hc17c5c5b} /* (11, 4, 0) {real, imag} */,
  {32'h421670dc, 32'h42d18c2c} /* (11, 3, 31) {real, imag} */,
  {32'hc1aecd40, 32'hc2ec4e8c} /* (11, 3, 30) {real, imag} */,
  {32'h425d3192, 32'h421e8724} /* (11, 3, 29) {real, imag} */,
  {32'h423e2f16, 32'hc1fef287} /* (11, 3, 28) {real, imag} */,
  {32'h41e9d9be, 32'hc2d46574} /* (11, 3, 27) {real, imag} */,
  {32'hc2362572, 32'h424bb2fc} /* (11, 3, 26) {real, imag} */,
  {32'hc2177fbe, 32'hc28bf6af} /* (11, 3, 25) {real, imag} */,
  {32'hc0a539ca, 32'hc213462c} /* (11, 3, 24) {real, imag} */,
  {32'h423731ec, 32'hc1d3a409} /* (11, 3, 23) {real, imag} */,
  {32'hc1f15ffb, 32'hc151bf00} /* (11, 3, 22) {real, imag} */,
  {32'hc2193792, 32'hc11ec22a} /* (11, 3, 21) {real, imag} */,
  {32'hc1684522, 32'h424161fe} /* (11, 3, 20) {real, imag} */,
  {32'hc156fe3e, 32'hc07c5114} /* (11, 3, 19) {real, imag} */,
  {32'hc1575624, 32'h4136da06} /* (11, 3, 18) {real, imag} */,
  {32'h40a99eea, 32'h4153fce4} /* (11, 3, 17) {real, imag} */,
  {32'hc1c0b7ca, 32'hc0bc4d74} /* (11, 3, 16) {real, imag} */,
  {32'hc116b1eb, 32'hc126c17c} /* (11, 3, 15) {real, imag} */,
  {32'h41991320, 32'h415a5932} /* (11, 3, 14) {real, imag} */,
  {32'h4153d8ca, 32'hc1037f39} /* (11, 3, 13) {real, imag} */,
  {32'hc17ac052, 32'h41d76bfc} /* (11, 3, 12) {real, imag} */,
  {32'h41c54f95, 32'h41ef5d21} /* (11, 3, 11) {real, imag} */,
  {32'hc1e11319, 32'hc08242f8} /* (11, 3, 10) {real, imag} */,
  {32'h426977fc, 32'hc1455ba2} /* (11, 3, 9) {real, imag} */,
  {32'hc1a04f96, 32'h42465aa8} /* (11, 3, 8) {real, imag} */,
  {32'h41b7b6b3, 32'h403d0ca0} /* (11, 3, 7) {real, imag} */,
  {32'h41a3589c, 32'hc1c78f07} /* (11, 3, 6) {real, imag} */,
  {32'hc1855296, 32'hc1a6675e} /* (11, 3, 5) {real, imag} */,
  {32'hc1def8d5, 32'h41ca4bc5} /* (11, 3, 4) {real, imag} */,
  {32'hc2a4247b, 32'hc22d38b8} /* (11, 3, 3) {real, imag} */,
  {32'hc2cf1c44, 32'hc05ad770} /* (11, 3, 2) {real, imag} */,
  {32'hc1d1ad44, 32'h423b4e40} /* (11, 3, 1) {real, imag} */,
  {32'h42ba135a, 32'h42278902} /* (11, 3, 0) {real, imag} */,
  {32'hc33c3263, 32'h42d1bb7f} /* (11, 2, 31) {real, imag} */,
  {32'h432e0860, 32'hc11b6c78} /* (11, 2, 30) {real, imag} */,
  {32'h40e7fe3c, 32'hbf710e08} /* (11, 2, 29) {real, imag} */,
  {32'h4167d2fe, 32'hc0a60dde} /* (11, 2, 28) {real, imag} */,
  {32'hc08da410, 32'h418e3108} /* (11, 2, 27) {real, imag} */,
  {32'h41809e13, 32'h423d9c0a} /* (11, 2, 26) {real, imag} */,
  {32'hc268fc3e, 32'h42c469b6} /* (11, 2, 25) {real, imag} */,
  {32'h41230510, 32'hc28b3c92} /* (11, 2, 24) {real, imag} */,
  {32'h424b74f4, 32'h4064d758} /* (11, 2, 23) {real, imag} */,
  {32'h40cd9ce0, 32'h4195fafc} /* (11, 2, 22) {real, imag} */,
  {32'h405df680, 32'hc164617d} /* (11, 2, 21) {real, imag} */,
  {32'hc16f5f7e, 32'h41ccaec0} /* (11, 2, 20) {real, imag} */,
  {32'h419c9836, 32'h40a8b91f} /* (11, 2, 19) {real, imag} */,
  {32'hc1164ff8, 32'h40205408} /* (11, 2, 18) {real, imag} */,
  {32'hc07a2250, 32'h41bfc457} /* (11, 2, 17) {real, imag} */,
  {32'h3cfc7000, 32'h4110b940} /* (11, 2, 16) {real, imag} */,
  {32'h410c3aec, 32'hc1f07907} /* (11, 2, 15) {real, imag} */,
  {32'hc1a0dfcc, 32'hc06b7b08} /* (11, 2, 14) {real, imag} */,
  {32'hc198eb9e, 32'hc0d3e1b7} /* (11, 2, 13) {real, imag} */,
  {32'h425e4fb8, 32'h401d8eb8} /* (11, 2, 12) {real, imag} */,
  {32'h41da163a, 32'h42274829} /* (11, 2, 11) {real, imag} */,
  {32'hc298d298, 32'hc0fb2f20} /* (11, 2, 10) {real, imag} */,
  {32'hc210f68e, 32'hc23614c6} /* (11, 2, 9) {real, imag} */,
  {32'hc1b62dc8, 32'h428a358c} /* (11, 2, 8) {real, imag} */,
  {32'h41dc593f, 32'h41dd1c48} /* (11, 2, 7) {real, imag} */,
  {32'h41a9a00f, 32'hc235bbba} /* (11, 2, 6) {real, imag} */,
  {32'h425cdd95, 32'h414addb5} /* (11, 2, 5) {real, imag} */,
  {32'hc24dcc10, 32'hc213aef0} /* (11, 2, 4) {real, imag} */,
  {32'hc1d02ca9, 32'hbf9f7e3c} /* (11, 2, 3) {real, imag} */,
  {32'h41935ba4, 32'hc30d5ed0} /* (11, 2, 2) {real, imag} */,
  {32'hc231cdd4, 32'h41fb0054} /* (11, 2, 1) {real, imag} */,
  {32'hc2c2e52d, 32'h40bf8a2d} /* (11, 2, 0) {real, imag} */,
  {32'h4212ec4a, 32'hc2b65580} /* (11, 1, 31) {real, imag} */,
  {32'hc2e804b2, 32'hc13335a4} /* (11, 1, 30) {real, imag} */,
  {32'hc121a5a4, 32'h423bdbe9} /* (11, 1, 29) {real, imag} */,
  {32'h424e8862, 32'h42fab04b} /* (11, 1, 28) {real, imag} */,
  {32'hc2f962e4, 32'h426499ec} /* (11, 1, 27) {real, imag} */,
  {32'hc25c4764, 32'h415d06a0} /* (11, 1, 26) {real, imag} */,
  {32'hc18e04c8, 32'hc24927b0} /* (11, 1, 25) {real, imag} */,
  {32'h41d3ef76, 32'hc2b8ce42} /* (11, 1, 24) {real, imag} */,
  {32'hc09839b0, 32'hc1711b6a} /* (11, 1, 23) {real, imag} */,
  {32'hc1016f1a, 32'hc1f89d11} /* (11, 1, 22) {real, imag} */,
  {32'hc0d453d8, 32'hc0fa42dd} /* (11, 1, 21) {real, imag} */,
  {32'h41249b5c, 32'h4223fddc} /* (11, 1, 20) {real, imag} */,
  {32'h40eed132, 32'hc1ee6321} /* (11, 1, 19) {real, imag} */,
  {32'hbff87520, 32'hc01077d0} /* (11, 1, 18) {real, imag} */,
  {32'h41f35378, 32'hc1b4b4e9} /* (11, 1, 17) {real, imag} */,
  {32'hc0a58fc0, 32'hc13d3a0c} /* (11, 1, 16) {real, imag} */,
  {32'hc0109d80, 32'h41a39d51} /* (11, 1, 15) {real, imag} */,
  {32'h42368971, 32'hc19a161d} /* (11, 1, 14) {real, imag} */,
  {32'h41859e02, 32'hc1030fb2} /* (11, 1, 13) {real, imag} */,
  {32'hc062a4f2, 32'h41961b9e} /* (11, 1, 12) {real, imag} */,
  {32'hc1ac187a, 32'hc0301426} /* (11, 1, 11) {real, imag} */,
  {32'hbf7d0720, 32'h41325f2e} /* (11, 1, 10) {real, imag} */,
  {32'h42399589, 32'hc1afd4ff} /* (11, 1, 9) {real, imag} */,
  {32'hc29fe38e, 32'h421ae5f3} /* (11, 1, 8) {real, imag} */,
  {32'hc2082297, 32'hc1d363dd} /* (11, 1, 7) {real, imag} */,
  {32'h42871bb1, 32'hc1802080} /* (11, 1, 6) {real, imag} */,
  {32'hc28da48c, 32'h41fb3658} /* (11, 1, 5) {real, imag} */,
  {32'h420b311e, 32'h422c1d86} /* (11, 1, 4) {real, imag} */,
  {32'h427c7ae7, 32'h41afc416} /* (11, 1, 3) {real, imag} */,
  {32'hc34201bd, 32'hc26675ab} /* (11, 1, 2) {real, imag} */,
  {32'h4389bb5d, 32'h41e41548} /* (11, 1, 1) {real, imag} */,
  {32'h432ee17c, 32'hc20d67ab} /* (11, 1, 0) {real, imag} */,
  {32'h42a158cc, 32'hc30f8097} /* (11, 0, 31) {real, imag} */,
  {32'h42f23554, 32'h41367684} /* (11, 0, 30) {real, imag} */,
  {32'h4213ceb4, 32'h42e2f660} /* (11, 0, 29) {real, imag} */,
  {32'h41884cec, 32'hc1822081} /* (11, 0, 28) {real, imag} */,
  {32'hc28d778b, 32'hc259270c} /* (11, 0, 27) {real, imag} */,
  {32'h41ccfd96, 32'hc113d1da} /* (11, 0, 26) {real, imag} */,
  {32'hc1456aa0, 32'h410d1200} /* (11, 0, 25) {real, imag} */,
  {32'h42add182, 32'h4304da6b} /* (11, 0, 24) {real, imag} */,
  {32'hc24b90e2, 32'h42883254} /* (11, 0, 23) {real, imag} */,
  {32'hc151326d, 32'h41dbb43f} /* (11, 0, 22) {real, imag} */,
  {32'h413cc302, 32'h41d0577e} /* (11, 0, 21) {real, imag} */,
  {32'h4137fa45, 32'hc0dd1d5e} /* (11, 0, 20) {real, imag} */,
  {32'hc12e1a53, 32'hc08b0c24} /* (11, 0, 19) {real, imag} */,
  {32'h4112c02a, 32'hc0805108} /* (11, 0, 18) {real, imag} */,
  {32'hc11270e4, 32'hc1936a36} /* (11, 0, 17) {real, imag} */,
  {32'h411fbf1c, 32'hc15a0d68} /* (11, 0, 16) {real, imag} */,
  {32'hc1184d5c, 32'h40d4afda} /* (11, 0, 15) {real, imag} */,
  {32'h3f3eb4a0, 32'hc21e6d29} /* (11, 0, 14) {real, imag} */,
  {32'hc1d44cb6, 32'hc1b1118d} /* (11, 0, 13) {real, imag} */,
  {32'h40e07e9e, 32'hc196b4f6} /* (11, 0, 12) {real, imag} */,
  {32'hc0c4be84, 32'hc16c669b} /* (11, 0, 11) {real, imag} */,
  {32'hc16a44b1, 32'hc108f04e} /* (11, 0, 10) {real, imag} */,
  {32'hc1de587b, 32'hc1f82914} /* (11, 0, 9) {real, imag} */,
  {32'hc1dbc6f8, 32'h418c5472} /* (11, 0, 8) {real, imag} */,
  {32'h420798e9, 32'hc260cba6} /* (11, 0, 7) {real, imag} */,
  {32'hc1da6568, 32'hc0fd54cc} /* (11, 0, 6) {real, imag} */,
  {32'h4202091e, 32'h4228a50e} /* (11, 0, 5) {real, imag} */,
  {32'h42955309, 32'hc15215ed} /* (11, 0, 4) {real, imag} */,
  {32'h420d6d40, 32'hc00c4090} /* (11, 0, 3) {real, imag} */,
  {32'hc1f89900, 32'hc3049586} /* (11, 0, 2) {real, imag} */,
  {32'h430c8344, 32'hc296a9aa} /* (11, 0, 1) {real, imag} */,
  {32'h430043e7, 32'hc29469d9} /* (11, 0, 0) {real, imag} */,
  {32'hc28184be, 32'h430a33cf} /* (10, 31, 31) {real, imag} */,
  {32'h41fbf3a8, 32'hc2bb3bc0} /* (10, 31, 30) {real, imag} */,
  {32'h430b1f1f, 32'hbed19380} /* (10, 31, 29) {real, imag} */,
  {32'hc22c0f48, 32'h4183e2a7} /* (10, 31, 28) {real, imag} */,
  {32'h430e4902, 32'hc233531a} /* (10, 31, 27) {real, imag} */,
  {32'h42209580, 32'hc201f27f} /* (10, 31, 26) {real, imag} */,
  {32'h40f7a0c8, 32'h42cc1d16} /* (10, 31, 25) {real, imag} */,
  {32'hc19d3590, 32'h41f143c3} /* (10, 31, 24) {real, imag} */,
  {32'hc288d1cb, 32'h41c0117e} /* (10, 31, 23) {real, imag} */,
  {32'h4107f248, 32'hc1ee0a9a} /* (10, 31, 22) {real, imag} */,
  {32'h4102383a, 32'h41e15c8e} /* (10, 31, 21) {real, imag} */,
  {32'hc195b554, 32'h3fc3f204} /* (10, 31, 20) {real, imag} */,
  {32'hc10df20c, 32'h40b2cb4c} /* (10, 31, 19) {real, imag} */,
  {32'hc16f7e37, 32'h4129fa84} /* (10, 31, 18) {real, imag} */,
  {32'h41563381, 32'hc12da518} /* (10, 31, 17) {real, imag} */,
  {32'h40f7de74, 32'hc000c740} /* (10, 31, 16) {real, imag} */,
  {32'hc1334ea9, 32'h41ac96c4} /* (10, 31, 15) {real, imag} */,
  {32'hc0e4c852, 32'h410586bc} /* (10, 31, 14) {real, imag} */,
  {32'h41ed6f72, 32'hc21eb2ec} /* (10, 31, 13) {real, imag} */,
  {32'h3feb7df8, 32'hc0f53a61} /* (10, 31, 12) {real, imag} */,
  {32'h4115c1c2, 32'h410a3ecc} /* (10, 31, 11) {real, imag} */,
  {32'h41e28d7c, 32'hc1b8c6da} /* (10, 31, 10) {real, imag} */,
  {32'h417bf7f6, 32'h40eca9d6} /* (10, 31, 9) {real, imag} */,
  {32'hc104b678, 32'hc26b227a} /* (10, 31, 8) {real, imag} */,
  {32'hc1ce67d0, 32'h421863fd} /* (10, 31, 7) {real, imag} */,
  {32'hc1afd438, 32'hc24011cf} /* (10, 31, 6) {real, imag} */,
  {32'hc1c2b6cc, 32'hc322a7d2} /* (10, 31, 5) {real, imag} */,
  {32'hc222c9c2, 32'h3f37d198} /* (10, 31, 4) {real, imag} */,
  {32'h41e55c78, 32'h42c69876} /* (10, 31, 3) {real, imag} */,
  {32'h42926038, 32'hc2d43dec} /* (10, 31, 2) {real, imag} */,
  {32'hc2be1d16, 32'h422c2e28} /* (10, 31, 1) {real, imag} */,
  {32'h428004c0, 32'h431b0ef1} /* (10, 31, 0) {real, imag} */,
  {32'h42072cea, 32'h429b8ce5} /* (10, 30, 31) {real, imag} */,
  {32'hc3260cb8, 32'hc0e2e706} /* (10, 30, 30) {real, imag} */,
  {32'hc157b53c, 32'hc2b74786} /* (10, 30, 29) {real, imag} */,
  {32'h41189127, 32'hc271f38c} /* (10, 30, 28) {real, imag} */,
  {32'hc2a2d138, 32'h422ffe4e} /* (10, 30, 27) {real, imag} */,
  {32'h40f5ad84, 32'h41c53d9c} /* (10, 30, 26) {real, imag} */,
  {32'h40ea310c, 32'hc2847d0a} /* (10, 30, 25) {real, imag} */,
  {32'hc232472e, 32'h42b6dbda} /* (10, 30, 24) {real, imag} */,
  {32'hc1d77a06, 32'h419f8722} /* (10, 30, 23) {real, imag} */,
  {32'hc182ab2e, 32'hc22285d2} /* (10, 30, 22) {real, imag} */,
  {32'hc001d6a8, 32'hc182f820} /* (10, 30, 21) {real, imag} */,
  {32'hc1a983d5, 32'h41d241f5} /* (10, 30, 20) {real, imag} */,
  {32'h40f556f4, 32'h41ed3bb7} /* (10, 30, 19) {real, imag} */,
  {32'h42084250, 32'h41d1461e} /* (10, 30, 18) {real, imag} */,
  {32'h40699422, 32'hc1017a3f} /* (10, 30, 17) {real, imag} */,
  {32'h40b1be10, 32'h3e816c40} /* (10, 30, 16) {real, imag} */,
  {32'hc1369048, 32'hc0b380ae} /* (10, 30, 15) {real, imag} */,
  {32'h416aa472, 32'hc1f2a8be} /* (10, 30, 14) {real, imag} */,
  {32'h410b5a02, 32'hc16836b6} /* (10, 30, 13) {real, imag} */,
  {32'hc1b5faf1, 32'hc2157f50} /* (10, 30, 12) {real, imag} */,
  {32'hc0dc41ec, 32'hc068b10e} /* (10, 30, 11) {real, imag} */,
  {32'h40966752, 32'h40f9ca18} /* (10, 30, 10) {real, imag} */,
  {32'hc207b34b, 32'hc0298230} /* (10, 30, 9) {real, imag} */,
  {32'hc27acf2e, 32'h41e52baa} /* (10, 30, 8) {real, imag} */,
  {32'hc11aaffe, 32'h42286028} /* (10, 30, 7) {real, imag} */,
  {32'h4205d68e, 32'hc2286cb6} /* (10, 30, 6) {real, imag} */,
  {32'hc0a96db8, 32'h427bef32} /* (10, 30, 5) {real, imag} */,
  {32'h418a9b63, 32'h433cd1b3} /* (10, 30, 4) {real, imag} */,
  {32'h42da1d30, 32'hc0c68f20} /* (10, 30, 3) {real, imag} */,
  {32'hc11a1328, 32'hc1616339} /* (10, 30, 2) {real, imag} */,
  {32'h4285900f, 32'hc2b98747} /* (10, 30, 1) {real, imag} */,
  {32'h431715d0, 32'hc1fb8353} /* (10, 30, 0) {real, imag} */,
  {32'hc28f24e1, 32'hc277d3e3} /* (10, 29, 31) {real, imag} */,
  {32'hc1a002b6, 32'hc256a662} /* (10, 29, 30) {real, imag} */,
  {32'hc257537a, 32'hc094999e} /* (10, 29, 29) {real, imag} */,
  {32'hc1ad4735, 32'h4119f237} /* (10, 29, 28) {real, imag} */,
  {32'hc20c7488, 32'h42b0def3} /* (10, 29, 27) {real, imag} */,
  {32'h418b71c2, 32'h42bbf80a} /* (10, 29, 26) {real, imag} */,
  {32'hc2053ce7, 32'hc18b72f0} /* (10, 29, 25) {real, imag} */,
  {32'hc1a6dbd1, 32'hc12751c4} /* (10, 29, 24) {real, imag} */,
  {32'h41d6f078, 32'h41c0e668} /* (10, 29, 23) {real, imag} */,
  {32'hc0398b10, 32'hc17bff1a} /* (10, 29, 22) {real, imag} */,
  {32'hc1a9b5ee, 32'hc10841ae} /* (10, 29, 21) {real, imag} */,
  {32'h4226126a, 32'hc0a6b94a} /* (10, 29, 20) {real, imag} */,
  {32'hc181bb5a, 32'hc0ee7bda} /* (10, 29, 19) {real, imag} */,
  {32'hc13b48bf, 32'hc1ecd170} /* (10, 29, 18) {real, imag} */,
  {32'h4110bb2b, 32'h40c980e0} /* (10, 29, 17) {real, imag} */,
  {32'h419f3a50, 32'hc18687ae} /* (10, 29, 16) {real, imag} */,
  {32'h3e8f32a0, 32'hc1405c78} /* (10, 29, 15) {real, imag} */,
  {32'hc126e4c9, 32'h420b50fe} /* (10, 29, 14) {real, imag} */,
  {32'hc0f04eee, 32'h4165f3eb} /* (10, 29, 13) {real, imag} */,
  {32'h410aa546, 32'h421268a5} /* (10, 29, 12) {real, imag} */,
  {32'hc1a1ec9e, 32'h41164dd2} /* (10, 29, 11) {real, imag} */,
  {32'hc27f76ff, 32'h41cdf09f} /* (10, 29, 10) {real, imag} */,
  {32'h41d70ba4, 32'h406f6330} /* (10, 29, 9) {real, imag} */,
  {32'h40e69854, 32'h42bcca7c} /* (10, 29, 8) {real, imag} */,
  {32'hc10c9c33, 32'h419c701a} /* (10, 29, 7) {real, imag} */,
  {32'h40da5dfa, 32'h41c9d220} /* (10, 29, 6) {real, imag} */,
  {32'h420b3df4, 32'hc2465ae2} /* (10, 29, 5) {real, imag} */,
  {32'h42216f78, 32'hc1d107bc} /* (10, 29, 4) {real, imag} */,
  {32'hc0dee60c, 32'h41b27a50} /* (10, 29, 3) {real, imag} */,
  {32'hc205a4fb, 32'hc2c87cef} /* (10, 29, 2) {real, imag} */,
  {32'hc2d17e2b, 32'hc26a49c3} /* (10, 29, 1) {real, imag} */,
  {32'hc28a40c4, 32'hc2c3f51c} /* (10, 29, 0) {real, imag} */,
  {32'h41bed296, 32'h425a4c6d} /* (10, 28, 31) {real, imag} */,
  {32'hc247f9a3, 32'hc29742a8} /* (10, 28, 30) {real, imag} */,
  {32'h3f95b9c0, 32'h41c25e72} /* (10, 28, 29) {real, imag} */,
  {32'hc3229947, 32'h401dc0e0} /* (10, 28, 28) {real, imag} */,
  {32'h40aa4924, 32'hc2487ac2} /* (10, 28, 27) {real, imag} */,
  {32'hbf782b00, 32'hc021a7f0} /* (10, 28, 26) {real, imag} */,
  {32'h422181dd, 32'h422dfb74} /* (10, 28, 25) {real, imag} */,
  {32'h42267643, 32'h41c1a2aa} /* (10, 28, 24) {real, imag} */,
  {32'h3fa8ab90, 32'hc200aa9f} /* (10, 28, 23) {real, imag} */,
  {32'h3eadaf80, 32'hc1fdbf71} /* (10, 28, 22) {real, imag} */,
  {32'h40b9f5f4, 32'h416d19c7} /* (10, 28, 21) {real, imag} */,
  {32'hc1892b08, 32'hc136c00e} /* (10, 28, 20) {real, imag} */,
  {32'h4130b353, 32'h410d9925} /* (10, 28, 19) {real, imag} */,
  {32'hc19af0fe, 32'h4147c150} /* (10, 28, 18) {real, imag} */,
  {32'h4111c835, 32'hc073593e} /* (10, 28, 17) {real, imag} */,
  {32'hc12d8ecd, 32'hc0ccdb78} /* (10, 28, 16) {real, imag} */,
  {32'h4132ef93, 32'h4183f170} /* (10, 28, 15) {real, imag} */,
  {32'hc180da32, 32'h41383dd8} /* (10, 28, 14) {real, imag} */,
  {32'h418153a6, 32'h40286184} /* (10, 28, 13) {real, imag} */,
  {32'hc28f32ac, 32'h4217e472} /* (10, 28, 12) {real, imag} */,
  {32'h42690be6, 32'hc08dc4b2} /* (10, 28, 11) {real, imag} */,
  {32'hc04a7460, 32'hc22a15e2} /* (10, 28, 10) {real, imag} */,
  {32'hc2260ca4, 32'hc14620e5} /* (10, 28, 9) {real, imag} */,
  {32'h41ced19a, 32'hc0598094} /* (10, 28, 8) {real, imag} */,
  {32'h4201a66b, 32'h41fb6d24} /* (10, 28, 7) {real, imag} */,
  {32'hc2a03e08, 32'h42b008b6} /* (10, 28, 6) {real, imag} */,
  {32'hc1f209fd, 32'hc191dc07} /* (10, 28, 5) {real, imag} */,
  {32'h40786880, 32'h42a18ca5} /* (10, 28, 4) {real, imag} */,
  {32'hc26abdc2, 32'hc287f844} /* (10, 28, 3) {real, imag} */,
  {32'h40cfffe8, 32'hc2815614} /* (10, 28, 2) {real, imag} */,
  {32'h421bb8d1, 32'hc1bb132e} /* (10, 28, 1) {real, imag} */,
  {32'hc15a6e33, 32'h422fd733} /* (10, 28, 0) {real, imag} */,
  {32'hc24cc130, 32'hc10ce612} /* (10, 27, 31) {real, imag} */,
  {32'hc21a64be, 32'h41123346} /* (10, 27, 30) {real, imag} */,
  {32'hc28818f6, 32'hc2370d73} /* (10, 27, 29) {real, imag} */,
  {32'h42563ccc, 32'hc27c0e48} /* (10, 27, 28) {real, imag} */,
  {32'h4121c9e4, 32'h424e569f} /* (10, 27, 27) {real, imag} */,
  {32'hc1fbc0e4, 32'hc2311268} /* (10, 27, 26) {real, imag} */,
  {32'hc10121ec, 32'h420419a2} /* (10, 27, 25) {real, imag} */,
  {32'hbfd0f010, 32'hc0e883e6} /* (10, 27, 24) {real, imag} */,
  {32'h41ae0453, 32'hc1dc963b} /* (10, 27, 23) {real, imag} */,
  {32'hc221da78, 32'h409fb594} /* (10, 27, 22) {real, imag} */,
  {32'h41e13377, 32'hc12f26bb} /* (10, 27, 21) {real, imag} */,
  {32'h40aaeef0, 32'h4134a39c} /* (10, 27, 20) {real, imag} */,
  {32'hc0153414, 32'h40e5d4f6} /* (10, 27, 19) {real, imag} */,
  {32'h410992b8, 32'h4130bff0} /* (10, 27, 18) {real, imag} */,
  {32'hbffb8d8c, 32'h40ac3908} /* (10, 27, 17) {real, imag} */,
  {32'hc1c94a8b, 32'h40eabda8} /* (10, 27, 16) {real, imag} */,
  {32'h40948c55, 32'hbe12c800} /* (10, 27, 15) {real, imag} */,
  {32'h41d98920, 32'hbffd8f84} /* (10, 27, 14) {real, imag} */,
  {32'h40a3c98e, 32'h405bd284} /* (10, 27, 13) {real, imag} */,
  {32'hc0bf2380, 32'hc1ad2a5c} /* (10, 27, 12) {real, imag} */,
  {32'h412179de, 32'hc1919650} /* (10, 27, 11) {real, imag} */,
  {32'h414d6c8c, 32'hc24df6dc} /* (10, 27, 10) {real, imag} */,
  {32'hc062b688, 32'h41a34629} /* (10, 27, 9) {real, imag} */,
  {32'hc200d7e2, 32'h413ba771} /* (10, 27, 8) {real, imag} */,
  {32'h4172ac28, 32'h41c6759b} /* (10, 27, 7) {real, imag} */,
  {32'h42016403, 32'h42820b25} /* (10, 27, 6) {real, imag} */,
  {32'h429e3c7a, 32'hc1babc1a} /* (10, 27, 5) {real, imag} */,
  {32'hc2cf66b6, 32'hc165a3f2} /* (10, 27, 4) {real, imag} */,
  {32'h41975872, 32'hc26c5661} /* (10, 27, 3) {real, imag} */,
  {32'h3fc69f80, 32'hc1cd49c1} /* (10, 27, 2) {real, imag} */,
  {32'h41bf4150, 32'h427353e0} /* (10, 27, 1) {real, imag} */,
  {32'h4240eb7e, 32'h422b54a1} /* (10, 27, 0) {real, imag} */,
  {32'h4024a368, 32'h41adbfa8} /* (10, 26, 31) {real, imag} */,
  {32'hc29951e6, 32'hc22b3936} /* (10, 26, 30) {real, imag} */,
  {32'hc0d54788, 32'h426c1de2} /* (10, 26, 29) {real, imag} */,
  {32'hc1036a54, 32'h41a0c17a} /* (10, 26, 28) {real, imag} */,
  {32'hc29bb504, 32'hc0b5aec8} /* (10, 26, 27) {real, imag} */,
  {32'h422436d6, 32'h4203405a} /* (10, 26, 26) {real, imag} */,
  {32'h415b27b0, 32'hc0efcf9c} /* (10, 26, 25) {real, imag} */,
  {32'h4228b453, 32'h40774134} /* (10, 26, 24) {real, imag} */,
  {32'hc097512a, 32'hc0ee94af} /* (10, 26, 23) {real, imag} */,
  {32'h4195909e, 32'h41b640c7} /* (10, 26, 22) {real, imag} */,
  {32'h40e58646, 32'hc2031486} /* (10, 26, 21) {real, imag} */,
  {32'h411c6ce2, 32'hc22e1455} /* (10, 26, 20) {real, imag} */,
  {32'h4222c31a, 32'hc1819602} /* (10, 26, 19) {real, imag} */,
  {32'hc12be22f, 32'h40a89990} /* (10, 26, 18) {real, imag} */,
  {32'h4180adb7, 32'h407cc022} /* (10, 26, 17) {real, imag} */,
  {32'hc055a100, 32'hc02635c0} /* (10, 26, 16) {real, imag} */,
  {32'hc12b4642, 32'hbf3edc58} /* (10, 26, 15) {real, imag} */,
  {32'hc0819dce, 32'hc1588b88} /* (10, 26, 14) {real, imag} */,
  {32'h41319e68, 32'h406b8800} /* (10, 26, 13) {real, imag} */,
  {32'h41a40041, 32'h405a6e90} /* (10, 26, 12) {real, imag} */,
  {32'hbfb8a3b8, 32'h42069e3e} /* (10, 26, 11) {real, imag} */,
  {32'h413c70d9, 32'h41b8d3f1} /* (10, 26, 10) {real, imag} */,
  {32'hc047b83c, 32'h4095e557} /* (10, 26, 9) {real, imag} */,
  {32'hc127e4bb, 32'h417d9855} /* (10, 26, 8) {real, imag} */,
  {32'h428cb446, 32'hc219968e} /* (10, 26, 7) {real, imag} */,
  {32'h40320b88, 32'h3fae6fc0} /* (10, 26, 6) {real, imag} */,
  {32'hc25e5a24, 32'hc2993b8c} /* (10, 26, 5) {real, imag} */,
  {32'hc2ab636c, 32'h418140a2} /* (10, 26, 4) {real, imag} */,
  {32'h42ad9b34, 32'h4150e2ba} /* (10, 26, 3) {real, imag} */,
  {32'h414e1008, 32'hc07c9ed8} /* (10, 26, 2) {real, imag} */,
  {32'h418f8319, 32'hc10b5302} /* (10, 26, 1) {real, imag} */,
  {32'h426622be, 32'hc2549026} /* (10, 26, 0) {real, imag} */,
  {32'h42818608, 32'hc27eb097} /* (10, 25, 31) {real, imag} */,
  {32'h41c91b39, 32'h418ff699} /* (10, 25, 30) {real, imag} */,
  {32'h427011d1, 32'hc1917bb6} /* (10, 25, 29) {real, imag} */,
  {32'h40cdf324, 32'h41dd2a7f} /* (10, 25, 28) {real, imag} */,
  {32'h4280e2c2, 32'h41c1fb37} /* (10, 25, 27) {real, imag} */,
  {32'h4274b02a, 32'hc2688172} /* (10, 25, 26) {real, imag} */,
  {32'h401274dc, 32'h425a80bc} /* (10, 25, 25) {real, imag} */,
  {32'hc1bab13e, 32'hc0f8c448} /* (10, 25, 24) {real, imag} */,
  {32'hbf19e270, 32'hc23410f4} /* (10, 25, 23) {real, imag} */,
  {32'hc205753b, 32'h42009b0c} /* (10, 25, 22) {real, imag} */,
  {32'hc17b46f9, 32'h417119fc} /* (10, 25, 21) {real, imag} */,
  {32'h411a7ab6, 32'h4137e46c} /* (10, 25, 20) {real, imag} */,
  {32'hc13aade8, 32'h413123f9} /* (10, 25, 19) {real, imag} */,
  {32'h3feb06d0, 32'h41943d1b} /* (10, 25, 18) {real, imag} */,
  {32'h4088ca16, 32'hc19607ab} /* (10, 25, 17) {real, imag} */,
  {32'hc11f2129, 32'hc0d1f640} /* (10, 25, 16) {real, imag} */,
  {32'hc0220b74, 32'h3ecfe2c0} /* (10, 25, 15) {real, imag} */,
  {32'h40b925ac, 32'h403d1798} /* (10, 25, 14) {real, imag} */,
  {32'hc1e8ef78, 32'hc0a66aa2} /* (10, 25, 13) {real, imag} */,
  {32'hc159ab76, 32'hc06916a2} /* (10, 25, 12) {real, imag} */,
  {32'hc1332e9f, 32'h41b2af5c} /* (10, 25, 11) {real, imag} */,
  {32'h41484413, 32'hc20c0556} /* (10, 25, 10) {real, imag} */,
  {32'hc0955cd2, 32'h41271a96} /* (10, 25, 9) {real, imag} */,
  {32'h41663495, 32'hc10b15b4} /* (10, 25, 8) {real, imag} */,
  {32'hc1a9c7a2, 32'h423759ce} /* (10, 25, 7) {real, imag} */,
  {32'hc280e30f, 32'hc16ccac8} /* (10, 25, 6) {real, imag} */,
  {32'h4250c816, 32'hc28113f2} /* (10, 25, 5) {real, imag} */,
  {32'h41cf448f, 32'hc00d63a8} /* (10, 25, 4) {real, imag} */,
  {32'hc27be6ed, 32'hc26c2633} /* (10, 25, 3) {real, imag} */,
  {32'hc1fd016d, 32'hc28808d9} /* (10, 25, 2) {real, imag} */,
  {32'hc1c8a368, 32'h41bbfad2} /* (10, 25, 1) {real, imag} */,
  {32'hc1cdfe28, 32'h420326d4} /* (10, 25, 0) {real, imag} */,
  {32'h4234157d, 32'h416fd780} /* (10, 24, 31) {real, imag} */,
  {32'hc1f399ba, 32'h4220904d} /* (10, 24, 30) {real, imag} */,
  {32'h419c2d02, 32'hc28a0e88} /* (10, 24, 29) {real, imag} */,
  {32'hc129b966, 32'h4221b7f8} /* (10, 24, 28) {real, imag} */,
  {32'h4293e828, 32'h42705e24} /* (10, 24, 27) {real, imag} */,
  {32'hc2a7bb70, 32'hc058eec8} /* (10, 24, 26) {real, imag} */,
  {32'hc2069d96, 32'hc237e284} /* (10, 24, 25) {real, imag} */,
  {32'hc135d876, 32'h3f24e194} /* (10, 24, 24) {real, imag} */,
  {32'h410e9d32, 32'h41827a0d} /* (10, 24, 23) {real, imag} */,
  {32'hc166f717, 32'h41d52a12} /* (10, 24, 22) {real, imag} */,
  {32'hc09d6abe, 32'hc171ab8b} /* (10, 24, 21) {real, imag} */,
  {32'h4184fdba, 32'hc1cd0b68} /* (10, 24, 20) {real, imag} */,
  {32'hc078ccaf, 32'hc135d143} /* (10, 24, 19) {real, imag} */,
  {32'h410913e0, 32'hc0a108b4} /* (10, 24, 18) {real, imag} */,
  {32'h4207ddd4, 32'h40c8622d} /* (10, 24, 17) {real, imag} */,
  {32'h401ed296, 32'h3f862108} /* (10, 24, 16) {real, imag} */,
  {32'hc1eb0244, 32'hbe3ab2e0} /* (10, 24, 15) {real, imag} */,
  {32'h41017004, 32'h3ff0cb60} /* (10, 24, 14) {real, imag} */,
  {32'hc12d6e2a, 32'h40807172} /* (10, 24, 13) {real, imag} */,
  {32'hc2165568, 32'h41105d17} /* (10, 24, 12) {real, imag} */,
  {32'h403c88c4, 32'h400c8cb4} /* (10, 24, 11) {real, imag} */,
  {32'hc0ea010a, 32'hc1101bff} /* (10, 24, 10) {real, imag} */,
  {32'h40bc943a, 32'h414ceed8} /* (10, 24, 9) {real, imag} */,
  {32'h4117813c, 32'hc03ccafb} /* (10, 24, 8) {real, imag} */,
  {32'h3e5e3400, 32'h4121a660} /* (10, 24, 7) {real, imag} */,
  {32'hc2536134, 32'h4216b73a} /* (10, 24, 6) {real, imag} */,
  {32'hc18f2a20, 32'hc22bc408} /* (10, 24, 5) {real, imag} */,
  {32'h40f3133c, 32'hc22d2c96} /* (10, 24, 4) {real, imag} */,
  {32'h418a8b56, 32'h4280052c} /* (10, 24, 3) {real, imag} */,
  {32'h41266b40, 32'h41d27dae} /* (10, 24, 2) {real, imag} */,
  {32'hbfebf4a0, 32'hc21143e8} /* (10, 24, 1) {real, imag} */,
  {32'hc08aa7dd, 32'h41495477} /* (10, 24, 0) {real, imag} */,
  {32'h40ac9fb4, 32'h4253d168} /* (10, 23, 31) {real, imag} */,
  {32'hc227b23f, 32'h417f4592} /* (10, 23, 30) {real, imag} */,
  {32'h41a52384, 32'h41b8906a} /* (10, 23, 29) {real, imag} */,
  {32'hc1edda62, 32'hc1d8ab08} /* (10, 23, 28) {real, imag} */,
  {32'hc1bd633c, 32'hc209aa56} /* (10, 23, 27) {real, imag} */,
  {32'h4235a9b0, 32'hc098b3a0} /* (10, 23, 26) {real, imag} */,
  {32'h414ecb8c, 32'hc1d8d31a} /* (10, 23, 25) {real, imag} */,
  {32'hc0a4e08f, 32'h41163a39} /* (10, 23, 24) {real, imag} */,
  {32'hc25090f2, 32'h3e4fa5a0} /* (10, 23, 23) {real, imag} */,
  {32'h414c4127, 32'h41d640dd} /* (10, 23, 22) {real, imag} */,
  {32'h41eb6f85, 32'hbfbfac68} /* (10, 23, 21) {real, imag} */,
  {32'h411212c2, 32'hc20b7dc5} /* (10, 23, 20) {real, imag} */,
  {32'hc06eda32, 32'h3f81d470} /* (10, 23, 19) {real, imag} */,
  {32'h419f8373, 32'hbf0ca400} /* (10, 23, 18) {real, imag} */,
  {32'h41266638, 32'h40e745e4} /* (10, 23, 17) {real, imag} */,
  {32'h40e52336, 32'h410cafe9} /* (10, 23, 16) {real, imag} */,
  {32'h40b4c529, 32'hc0e8bb28} /* (10, 23, 15) {real, imag} */,
  {32'hc0cc26b8, 32'hc090dd18} /* (10, 23, 14) {real, imag} */,
  {32'h413e552e, 32'hc1be84cb} /* (10, 23, 13) {real, imag} */,
  {32'h41cdac43, 32'hc0759b54} /* (10, 23, 12) {real, imag} */,
  {32'hc19390bf, 32'h4197d3d6} /* (10, 23, 11) {real, imag} */,
  {32'hc1cc9cf4, 32'hc0e101b4} /* (10, 23, 10) {real, imag} */,
  {32'h41d706c9, 32'hc10ab334} /* (10, 23, 9) {real, imag} */,
  {32'h4099ca31, 32'hc1b2b346} /* (10, 23, 8) {real, imag} */,
  {32'hc21fd758, 32'h41a76bf2} /* (10, 23, 7) {real, imag} */,
  {32'hc1cf7588, 32'hc219b4cf} /* (10, 23, 6) {real, imag} */,
  {32'hc154e379, 32'h41e5e518} /* (10, 23, 5) {real, imag} */,
  {32'h4244af63, 32'hc04d91dc} /* (10, 23, 4) {real, imag} */,
  {32'h408a22da, 32'h421a295d} /* (10, 23, 3) {real, imag} */,
  {32'h421e6e61, 32'hc248d728} /* (10, 23, 2) {real, imag} */,
  {32'h41e58b09, 32'hc169b678} /* (10, 23, 1) {real, imag} */,
  {32'hbff2be90, 32'hc1468033} /* (10, 23, 0) {real, imag} */,
  {32'hc1aa401c, 32'h41923bb8} /* (10, 22, 31) {real, imag} */,
  {32'h4188fc70, 32'hc1baf11e} /* (10, 22, 30) {real, imag} */,
  {32'hc1d58716, 32'h403a2c98} /* (10, 22, 29) {real, imag} */,
  {32'h4124be8e, 32'h41f03832} /* (10, 22, 28) {real, imag} */,
  {32'h40ba0b82, 32'hc26301aa} /* (10, 22, 27) {real, imag} */,
  {32'hc1d79f00, 32'hc24b9820} /* (10, 22, 26) {real, imag} */,
  {32'h412f00f0, 32'h41e0ba68} /* (10, 22, 25) {real, imag} */,
  {32'hc17861a6, 32'hc1da4eef} /* (10, 22, 24) {real, imag} */,
  {32'hc17efbb8, 32'h3f9f8580} /* (10, 22, 23) {real, imag} */,
  {32'h40f51834, 32'hc1c9d1b4} /* (10, 22, 22) {real, imag} */,
  {32'h3fd1cc18, 32'hc086c524} /* (10, 22, 21) {real, imag} */,
  {32'hc1837b70, 32'hbfdd15d4} /* (10, 22, 20) {real, imag} */,
  {32'hc196542d, 32'h404dce80} /* (10, 22, 19) {real, imag} */,
  {32'h412230b9, 32'hc08f74ea} /* (10, 22, 18) {real, imag} */,
  {32'h3f9c8f74, 32'h412ea8a6} /* (10, 22, 17) {real, imag} */,
  {32'hc010e1b2, 32'hc0a0f098} /* (10, 22, 16) {real, imag} */,
  {32'hc089b2ad, 32'hc0bc4cc4} /* (10, 22, 15) {real, imag} */,
  {32'hc0e0668e, 32'hc077f234} /* (10, 22, 14) {real, imag} */,
  {32'hc1549d3e, 32'hc1b858fa} /* (10, 22, 13) {real, imag} */,
  {32'h4037d92c, 32'hbfb82084} /* (10, 22, 12) {real, imag} */,
  {32'hc1a0aec6, 32'hbfed6c10} /* (10, 22, 11) {real, imag} */,
  {32'h4135e294, 32'hc0bd1c6e} /* (10, 22, 10) {real, imag} */,
  {32'h4100e9fa, 32'hbf84b2c8} /* (10, 22, 9) {real, imag} */,
  {32'h404050fa, 32'hc179c9be} /* (10, 22, 8) {real, imag} */,
  {32'h407251a8, 32'h40821f60} /* (10, 22, 7) {real, imag} */,
  {32'hc0fbd1f2, 32'hc0960560} /* (10, 22, 6) {real, imag} */,
  {32'h41a88a70, 32'hbf3c0e40} /* (10, 22, 5) {real, imag} */,
  {32'h419b38c0, 32'h404a2610} /* (10, 22, 4) {real, imag} */,
  {32'hc1d6a3d2, 32'h41ad0527} /* (10, 22, 3) {real, imag} */,
  {32'hc1ca27ca, 32'h420a6b11} /* (10, 22, 2) {real, imag} */,
  {32'h41227ac4, 32'h4083080f} /* (10, 22, 1) {real, imag} */,
  {32'h417b6afc, 32'hc22e48de} /* (10, 22, 0) {real, imag} */,
  {32'h40253cc0, 32'hc178a03e} /* (10, 21, 31) {real, imag} */,
  {32'hc1efbda2, 32'hc012548c} /* (10, 21, 30) {real, imag} */,
  {32'h41116f16, 32'h423c75d2} /* (10, 21, 29) {real, imag} */,
  {32'h40ea5390, 32'hc154d069} /* (10, 21, 28) {real, imag} */,
  {32'h414aaec6, 32'h424c3815} /* (10, 21, 27) {real, imag} */,
  {32'hc216e617, 32'hc1830648} /* (10, 21, 26) {real, imag} */,
  {32'hc1e932df, 32'hc1b870d1} /* (10, 21, 25) {real, imag} */,
  {32'hc0c6b70d, 32'hc0fe6d1e} /* (10, 21, 24) {real, imag} */,
  {32'hc0e4bf68, 32'hc093fa9c} /* (10, 21, 23) {real, imag} */,
  {32'hc0e03904, 32'h4188d374} /* (10, 21, 22) {real, imag} */,
  {32'h410bfd20, 32'h3fe39580} /* (10, 21, 21) {real, imag} */,
  {32'h410a420d, 32'hc0b02b94} /* (10, 21, 20) {real, imag} */,
  {32'h4103a818, 32'hc10ca713} /* (10, 21, 19) {real, imag} */,
  {32'hc0f6d778, 32'h40c31b80} /* (10, 21, 18) {real, imag} */,
  {32'hbf4558c0, 32'hc0e3815d} /* (10, 21, 17) {real, imag} */,
  {32'h41179b6c, 32'h4100a64b} /* (10, 21, 16) {real, imag} */,
  {32'h40759a30, 32'h3f172b08} /* (10, 21, 15) {real, imag} */,
  {32'hc1659e50, 32'hc019fef8} /* (10, 21, 14) {real, imag} */,
  {32'hbea5d608, 32'h4185c4cc} /* (10, 21, 13) {real, imag} */,
  {32'hc137a913, 32'h4085ec66} /* (10, 21, 12) {real, imag} */,
  {32'h419b02a0, 32'h41753160} /* (10, 21, 11) {real, imag} */,
  {32'hc0b1ec64, 32'h3ebae660} /* (10, 21, 10) {real, imag} */,
  {32'h4200932a, 32'hc1ca829d} /* (10, 21, 9) {real, imag} */,
  {32'hc0eaf78b, 32'h420fd5e3} /* (10, 21, 8) {real, imag} */,
  {32'h3fcc0af0, 32'hc110589e} /* (10, 21, 7) {real, imag} */,
  {32'h420286c5, 32'h42308b47} /* (10, 21, 6) {real, imag} */,
  {32'hc1a61fa1, 32'h41c05656} /* (10, 21, 5) {real, imag} */,
  {32'hc0b7cd2a, 32'h4123cd8b} /* (10, 21, 4) {real, imag} */,
  {32'h413bf346, 32'hbfa36810} /* (10, 21, 3) {real, imag} */,
  {32'h417f68c4, 32'hc164c3b5} /* (10, 21, 2) {real, imag} */,
  {32'hc228fb60, 32'h41a8bff3} /* (10, 21, 1) {real, imag} */,
  {32'h4226379a, 32'hc198abee} /* (10, 21, 0) {real, imag} */,
  {32'h41a40079, 32'h40b358f0} /* (10, 20, 31) {real, imag} */,
  {32'h3febff34, 32'hc1958b6b} /* (10, 20, 30) {real, imag} */,
  {32'hc20fbef4, 32'hc18f35f8} /* (10, 20, 29) {real, imag} */,
  {32'h41e2f5f4, 32'hc08c6bc2} /* (10, 20, 28) {real, imag} */,
  {32'hbfd6db66, 32'hc000ba04} /* (10, 20, 27) {real, imag} */,
  {32'hc1a5b2a6, 32'hc18536c7} /* (10, 20, 26) {real, imag} */,
  {32'h418a1e34, 32'hc1dbaf9b} /* (10, 20, 25) {real, imag} */,
  {32'h41081732, 32'hc0e96110} /* (10, 20, 24) {real, imag} */,
  {32'h4094bcf0, 32'h411d2172} /* (10, 20, 23) {real, imag} */,
  {32'h4090eb62, 32'hc0ee7821} /* (10, 20, 22) {real, imag} */,
  {32'h40bba370, 32'hc0e759f5} /* (10, 20, 21) {real, imag} */,
  {32'hc11357b2, 32'h40f855cc} /* (10, 20, 20) {real, imag} */,
  {32'h3f3f559c, 32'h40db704f} /* (10, 20, 19) {real, imag} */,
  {32'hc0ad1a2c, 32'hc0004bda} /* (10, 20, 18) {real, imag} */,
  {32'hbfc0bd0e, 32'h3edaec00} /* (10, 20, 17) {real, imag} */,
  {32'h4181d1da, 32'h3f8ffef8} /* (10, 20, 16) {real, imag} */,
  {32'hc058a193, 32'h40ee06e8} /* (10, 20, 15) {real, imag} */,
  {32'h414e5b8e, 32'hc147c4b8} /* (10, 20, 14) {real, imag} */,
  {32'h40cc3fb8, 32'hbf756bf0} /* (10, 20, 13) {real, imag} */,
  {32'hc153377e, 32'h413bd60e} /* (10, 20, 12) {real, imag} */,
  {32'hc1225188, 32'hbf542a58} /* (10, 20, 11) {real, imag} */,
  {32'hc1923d74, 32'h3d8ec740} /* (10, 20, 10) {real, imag} */,
  {32'hc167709c, 32'h4139d1d6} /* (10, 20, 9) {real, imag} */,
  {32'hc088ef0d, 32'h417f0422} /* (10, 20, 8) {real, imag} */,
  {32'hc1896182, 32'h41bce8af} /* (10, 20, 7) {real, imag} */,
  {32'h41fee736, 32'hc2050f00} /* (10, 20, 6) {real, imag} */,
  {32'h3ff8c5c2, 32'hbe9356bc} /* (10, 20, 5) {real, imag} */,
  {32'hc1bcd3f0, 32'hc1eeddc0} /* (10, 20, 4) {real, imag} */,
  {32'hc20298e4, 32'hc042bcd8} /* (10, 20, 3) {real, imag} */,
  {32'h41417b96, 32'h40408922} /* (10, 20, 2) {real, imag} */,
  {32'hc09cadbc, 32'h42046c55} /* (10, 20, 1) {real, imag} */,
  {32'h411ba083, 32'h41e59cc4} /* (10, 20, 0) {real, imag} */,
  {32'hc0b63828, 32'h410de5de} /* (10, 19, 31) {real, imag} */,
  {32'hc1ba7294, 32'h419921cc} /* (10, 19, 30) {real, imag} */,
  {32'h417e5123, 32'hc13158da} /* (10, 19, 29) {real, imag} */,
  {32'h421dc56e, 32'hbfec2024} /* (10, 19, 28) {real, imag} */,
  {32'hc1dc66fb, 32'h41bcb944} /* (10, 19, 27) {real, imag} */,
  {32'h4166bcea, 32'h40987b26} /* (10, 19, 26) {real, imag} */,
  {32'hc18ed20f, 32'h415b4586} /* (10, 19, 25) {real, imag} */,
  {32'h40467a62, 32'h41310aba} /* (10, 19, 24) {real, imag} */,
  {32'hc169bbf2, 32'hc1a52612} /* (10, 19, 23) {real, imag} */,
  {32'h4139a1e6, 32'hc17dc02a} /* (10, 19, 22) {real, imag} */,
  {32'h3ec9a9e0, 32'hc18821e2} /* (10, 19, 21) {real, imag} */,
  {32'h400c8ddc, 32'h4053abee} /* (10, 19, 20) {real, imag} */,
  {32'hc0f64e1a, 32'h40a89cbe} /* (10, 19, 19) {real, imag} */,
  {32'h403fe470, 32'h4100ea52} /* (10, 19, 18) {real, imag} */,
  {32'h41114d60, 32'hc11b1d2c} /* (10, 19, 17) {real, imag} */,
  {32'h410e8131, 32'hc0b321e0} /* (10, 19, 16) {real, imag} */,
  {32'h404dbcf0, 32'h40925c23} /* (10, 19, 15) {real, imag} */,
  {32'h3f8566a0, 32'h41798f22} /* (10, 19, 14) {real, imag} */,
  {32'h40edfbe0, 32'h411d2883} /* (10, 19, 13) {real, imag} */,
  {32'hc0cd0002, 32'hc0eff78f} /* (10, 19, 12) {real, imag} */,
  {32'hc0ec1614, 32'hc0b84dce} /* (10, 19, 11) {real, imag} */,
  {32'h40d324b4, 32'h418748e5} /* (10, 19, 10) {real, imag} */,
  {32'hc19632c9, 32'hc0b4675e} /* (10, 19, 9) {real, imag} */,
  {32'hc0eff44f, 32'h40331848} /* (10, 19, 8) {real, imag} */,
  {32'h413543ae, 32'hc14f8bfc} /* (10, 19, 7) {real, imag} */,
  {32'h426f25ca, 32'hc1b59b84} /* (10, 19, 6) {real, imag} */,
  {32'h406fb538, 32'h3dd8c780} /* (10, 19, 5) {real, imag} */,
  {32'hc18128f0, 32'hc1334de6} /* (10, 19, 4) {real, imag} */,
  {32'hc1e3263e, 32'h3f4a6560} /* (10, 19, 3) {real, imag} */,
  {32'h41d104d4, 32'h415d76c5} /* (10, 19, 2) {real, imag} */,
  {32'h41a961be, 32'hbd8bf640} /* (10, 19, 1) {real, imag} */,
  {32'hc11dec5f, 32'hc091670c} /* (10, 19, 0) {real, imag} */,
  {32'hbeb84500, 32'hc0e5ed09} /* (10, 18, 31) {real, imag} */,
  {32'h4056982e, 32'h41efe047} /* (10, 18, 30) {real, imag} */,
  {32'h3e9a26b0, 32'hc0f36b50} /* (10, 18, 29) {real, imag} */,
  {32'h41aaa660, 32'hc12cc4f1} /* (10, 18, 28) {real, imag} */,
  {32'h413bb12a, 32'h4147d1b2} /* (10, 18, 27) {real, imag} */,
  {32'hc1145ed7, 32'hc082ae28} /* (10, 18, 26) {real, imag} */,
  {32'h411fadb0, 32'h40d4a2e6} /* (10, 18, 25) {real, imag} */,
  {32'hbf08d8dc, 32'h40d2aca1} /* (10, 18, 24) {real, imag} */,
  {32'h41861549, 32'h40f1ac85} /* (10, 18, 23) {real, imag} */,
  {32'h4117150f, 32'h41843ed9} /* (10, 18, 22) {real, imag} */,
  {32'hc0e07a54, 32'hc05d8870} /* (10, 18, 21) {real, imag} */,
  {32'hc11df454, 32'h40eab77e} /* (10, 18, 20) {real, imag} */,
  {32'h3f9258e4, 32'h40607f4f} /* (10, 18, 19) {real, imag} */,
  {32'hc11ec414, 32'h3ff55e76} /* (10, 18, 18) {real, imag} */,
  {32'h40242090, 32'h4052b737} /* (10, 18, 17) {real, imag} */,
  {32'hbfa18bd8, 32'h4001b17c} /* (10, 18, 16) {real, imag} */,
  {32'hc05b1958, 32'hc01c9d93} /* (10, 18, 15) {real, imag} */,
  {32'h4052a716, 32'h408e57c6} /* (10, 18, 14) {real, imag} */,
  {32'hc0c8b249, 32'h408d834c} /* (10, 18, 13) {real, imag} */,
  {32'h41493826, 32'hc1d48af2} /* (10, 18, 12) {real, imag} */,
  {32'hbf4aa6a0, 32'hc0bebfa6} /* (10, 18, 11) {real, imag} */,
  {32'h40f04623, 32'h4178027a} /* (10, 18, 10) {real, imag} */,
  {32'hc11f0cd1, 32'hc0e449fb} /* (10, 18, 9) {real, imag} */,
  {32'h4103e098, 32'hc0af2957} /* (10, 18, 8) {real, imag} */,
  {32'h3fd97cb4, 32'hc0f81dc6} /* (10, 18, 7) {real, imag} */,
  {32'hc1018001, 32'h411f34a8} /* (10, 18, 6) {real, imag} */,
  {32'h41eaa661, 32'hc142d186} /* (10, 18, 5) {real, imag} */,
  {32'h40c7e722, 32'h412408ab} /* (10, 18, 4) {real, imag} */,
  {32'h40f264c9, 32'hc18395c5} /* (10, 18, 3) {real, imag} */,
  {32'h3ee48c4c, 32'h41a77b49} /* (10, 18, 2) {real, imag} */,
  {32'h421b2446, 32'h403904d6} /* (10, 18, 1) {real, imag} */,
  {32'hc12785c3, 32'hc1c5edd4} /* (10, 18, 0) {real, imag} */,
  {32'hc110bc4d, 32'h410ab0c4} /* (10, 17, 31) {real, imag} */,
  {32'h40e7f0f0, 32'hc1f28f61} /* (10, 17, 30) {real, imag} */,
  {32'hc04d92b2, 32'hc143598a} /* (10, 17, 29) {real, imag} */,
  {32'h4097fd34, 32'h4087a3de} /* (10, 17, 28) {real, imag} */,
  {32'hc1283058, 32'hc10cb17d} /* (10, 17, 27) {real, imag} */,
  {32'h407d34c0, 32'h40f23a7e} /* (10, 17, 26) {real, imag} */,
  {32'h4097a21a, 32'h413be796} /* (10, 17, 25) {real, imag} */,
  {32'h410b9965, 32'h41219c96} /* (10, 17, 24) {real, imag} */,
  {32'h41c3a501, 32'h3a496000} /* (10, 17, 23) {real, imag} */,
  {32'hc143e8e6, 32'hc0669f10} /* (10, 17, 22) {real, imag} */,
  {32'hbfb72755, 32'h3f89c330} /* (10, 17, 21) {real, imag} */,
  {32'h3e9c4c20, 32'h412341dc} /* (10, 17, 20) {real, imag} */,
  {32'h409d8868, 32'hc0eb0fa0} /* (10, 17, 19) {real, imag} */,
  {32'h402850f6, 32'hc0ac2784} /* (10, 17, 18) {real, imag} */,
  {32'hbc09d700, 32'h3ed073d8} /* (10, 17, 17) {real, imag} */,
  {32'hbf0fc3f8, 32'hbe3d7080} /* (10, 17, 16) {real, imag} */,
  {32'h408f3c18, 32'h3cbab580} /* (10, 17, 15) {real, imag} */,
  {32'h410a3788, 32'hbfa51ab0} /* (10, 17, 14) {real, imag} */,
  {32'h4012c526, 32'h40997cb2} /* (10, 17, 13) {real, imag} */,
  {32'hc095e1aa, 32'hbfcdc874} /* (10, 17, 12) {real, imag} */,
  {32'h40589c46, 32'h40cc273f} /* (10, 17, 11) {real, imag} */,
  {32'hc134e49a, 32'h40be73d4} /* (10, 17, 10) {real, imag} */,
  {32'h3fc1f130, 32'h40f96428} /* (10, 17, 9) {real, imag} */,
  {32'hbf997938, 32'hc18505fb} /* (10, 17, 8) {real, imag} */,
  {32'h402393b0, 32'hc095ad3c} /* (10, 17, 7) {real, imag} */,
  {32'hc089c5e8, 32'hc175cdd3} /* (10, 17, 6) {real, imag} */,
  {32'h403657c2, 32'hc115c76d} /* (10, 17, 5) {real, imag} */,
  {32'hc1b5a99e, 32'h41fcaf22} /* (10, 17, 4) {real, imag} */,
  {32'h4090e7a6, 32'h412e43ae} /* (10, 17, 3) {real, imag} */,
  {32'h3f5c3630, 32'hc1b93993} /* (10, 17, 2) {real, imag} */,
  {32'h40032fc3, 32'hbf93cbf2} /* (10, 17, 1) {real, imag} */,
  {32'h413de90c, 32'hc040fe68} /* (10, 17, 0) {real, imag} */,
  {32'hc1a5453d, 32'hc0ac8c80} /* (10, 16, 31) {real, imag} */,
  {32'h4009e580, 32'hc0aa6600} /* (10, 16, 30) {real, imag} */,
  {32'hc1aeefda, 32'hc0aaa78e} /* (10, 16, 29) {real, imag} */,
  {32'hc1dbafb6, 32'hc0bf50d1} /* (10, 16, 28) {real, imag} */,
  {32'hc1125f06, 32'h4164976e} /* (10, 16, 27) {real, imag} */,
  {32'h412b71b6, 32'hc10bbc37} /* (10, 16, 26) {real, imag} */,
  {32'h405816f7, 32'h42067e7f} /* (10, 16, 25) {real, imag} */,
  {32'hc0cebfc1, 32'hc01c4ee0} /* (10, 16, 24) {real, imag} */,
  {32'h4179b185, 32'hc106ae3e} /* (10, 16, 23) {real, imag} */,
  {32'hc09053fc, 32'h3e4510b8} /* (10, 16, 22) {real, imag} */,
  {32'hc10ef656, 32'hbe3320e0} /* (10, 16, 21) {real, imag} */,
  {32'hc11d1821, 32'h40b98ca4} /* (10, 16, 20) {real, imag} */,
  {32'h4048f4d5, 32'h408eaeee} /* (10, 16, 19) {real, imag} */,
  {32'h4067fb03, 32'hc085d71e} /* (10, 16, 18) {real, imag} */,
  {32'h403b3693, 32'h40a38305} /* (10, 16, 17) {real, imag} */,
  {32'hbfce95ec, 32'hbf9f1da4} /* (10, 16, 16) {real, imag} */,
  {32'h4040d3ab, 32'hc09d9b57} /* (10, 16, 15) {real, imag} */,
  {32'h40a00482, 32'h40a8780e} /* (10, 16, 14) {real, imag} */,
  {32'hc0c77be6, 32'h3fd3d458} /* (10, 16, 13) {real, imag} */,
  {32'h3ee9eea0, 32'h40704145} /* (10, 16, 12) {real, imag} */,
  {32'h3f09c568, 32'h40f117d1} /* (10, 16, 11) {real, imag} */,
  {32'h40003e33, 32'h3d0a94e0} /* (10, 16, 10) {real, imag} */,
  {32'h407c2e1c, 32'hc09838e8} /* (10, 16, 9) {real, imag} */,
  {32'hc12fa148, 32'h411e0ac6} /* (10, 16, 8) {real, imag} */,
  {32'hbe8ea178, 32'hbfdf18a8} /* (10, 16, 7) {real, imag} */,
  {32'hc0bc3174, 32'h40f54e17} /* (10, 16, 6) {real, imag} */,
  {32'h40c17c99, 32'hc157a39e} /* (10, 16, 5) {real, imag} */,
  {32'h41b357e2, 32'h412071cc} /* (10, 16, 4) {real, imag} */,
  {32'h41c75f52, 32'h418248b8} /* (10, 16, 3) {real, imag} */,
  {32'h41907af6, 32'hc10ec676} /* (10, 16, 2) {real, imag} */,
  {32'h41beff5f, 32'h41013de2} /* (10, 16, 1) {real, imag} */,
  {32'h418bcb55, 32'h40562c5a} /* (10, 16, 0) {real, imag} */,
  {32'hc0337599, 32'h4133453f} /* (10, 15, 31) {real, imag} */,
  {32'h416a758c, 32'h4122d10a} /* (10, 15, 30) {real, imag} */,
  {32'h415b2a12, 32'h419a80e8} /* (10, 15, 29) {real, imag} */,
  {32'hc0f3cc35, 32'hc0089e8f} /* (10, 15, 28) {real, imag} */,
  {32'hc1656444, 32'hbd689500} /* (10, 15, 27) {real, imag} */,
  {32'hc0d67327, 32'hc0926406} /* (10, 15, 26) {real, imag} */,
  {32'h41c6e286, 32'hc20f1630} /* (10, 15, 25) {real, imag} */,
  {32'hbf3b6d40, 32'h419dd63a} /* (10, 15, 24) {real, imag} */,
  {32'hc19702d2, 32'h41278fd5} /* (10, 15, 23) {real, imag} */,
  {32'h417d2cf1, 32'h40084da1} /* (10, 15, 22) {real, imag} */,
  {32'hc01da660, 32'h40b5e924} /* (10, 15, 21) {real, imag} */,
  {32'hbe91f6a0, 32'hc10db16a} /* (10, 15, 20) {real, imag} */,
  {32'h40901349, 32'h4179d812} /* (10, 15, 19) {real, imag} */,
  {32'h4035ade4, 32'hc08cda2f} /* (10, 15, 18) {real, imag} */,
  {32'hbf70398c, 32'hbffeba7e} /* (10, 15, 17) {real, imag} */,
  {32'h40310854, 32'h3fcabd30} /* (10, 15, 16) {real, imag} */,
  {32'hbf991cbe, 32'hc040acf7} /* (10, 15, 15) {real, imag} */,
  {32'hc0ad7c66, 32'h413726a6} /* (10, 15, 14) {real, imag} */,
  {32'hbfd67044, 32'hc1347b6a} /* (10, 15, 13) {real, imag} */,
  {32'hbfe80294, 32'h40a9e474} /* (10, 15, 12) {real, imag} */,
  {32'h40c347e0, 32'hc14a6ca6} /* (10, 15, 11) {real, imag} */,
  {32'hc07b304c, 32'h40bf2ce8} /* (10, 15, 10) {real, imag} */,
  {32'h4021c81c, 32'hc1857ff6} /* (10, 15, 9) {real, imag} */,
  {32'h40110e48, 32'h3f58e410} /* (10, 15, 8) {real, imag} */,
  {32'h40f2a822, 32'h419c5f3f} /* (10, 15, 7) {real, imag} */,
  {32'hc03f1122, 32'h4024f1dd} /* (10, 15, 6) {real, imag} */,
  {32'h41e24eb2, 32'h3fe2b648} /* (10, 15, 5) {real, imag} */,
  {32'h41137b40, 32'h3f77da05} /* (10, 15, 4) {real, imag} */,
  {32'h4059981a, 32'hc06ca6ee} /* (10, 15, 3) {real, imag} */,
  {32'h4036af38, 32'h40a3d715} /* (10, 15, 2) {real, imag} */,
  {32'hc04ab125, 32'hc0d41336} /* (10, 15, 1) {real, imag} */,
  {32'h3fa88f88, 32'h41dd0e40} /* (10, 15, 0) {real, imag} */,
  {32'h3ffa3d90, 32'h40749eb0} /* (10, 14, 31) {real, imag} */,
  {32'h41b5fe9c, 32'h4029252a} /* (10, 14, 30) {real, imag} */,
  {32'hc18ef8dc, 32'hc13987fd} /* (10, 14, 29) {real, imag} */,
  {32'h419385ba, 32'h4004878c} /* (10, 14, 28) {real, imag} */,
  {32'h3f0695b8, 32'h41aba2dc} /* (10, 14, 27) {real, imag} */,
  {32'h41205ea8, 32'hc184ace0} /* (10, 14, 26) {real, imag} */,
  {32'hc10d0705, 32'hc14068a0} /* (10, 14, 25) {real, imag} */,
  {32'h40701696, 32'hc09949da} /* (10, 14, 24) {real, imag} */,
  {32'h41144ff9, 32'hc17a80d2} /* (10, 14, 23) {real, imag} */,
  {32'h4166b0e8, 32'h400cae50} /* (10, 14, 22) {real, imag} */,
  {32'h412ac02f, 32'h40b6391c} /* (10, 14, 21) {real, imag} */,
  {32'h415a9fee, 32'h40881e53} /* (10, 14, 20) {real, imag} */,
  {32'hc0ea1976, 32'hbf5e2760} /* (10, 14, 19) {real, imag} */,
  {32'hc0d49248, 32'hbf184d68} /* (10, 14, 18) {real, imag} */,
  {32'hc05e035c, 32'hc14756af} /* (10, 14, 17) {real, imag} */,
  {32'h404a3f58, 32'hbf2ac338} /* (10, 14, 16) {real, imag} */,
  {32'hc083bc66, 32'h40d80182} /* (10, 14, 15) {real, imag} */,
  {32'hbfa4ae10, 32'h40ff98cd} /* (10, 14, 14) {real, imag} */,
  {32'hbebceaf8, 32'h3f640348} /* (10, 14, 13) {real, imag} */,
  {32'h40f2705c, 32'h40cde891} /* (10, 14, 12) {real, imag} */,
  {32'hc12fe7a9, 32'hc06d8158} /* (10, 14, 11) {real, imag} */,
  {32'h40123320, 32'hc1aea1db} /* (10, 14, 10) {real, imag} */,
  {32'hc1902a6c, 32'hc0c6d2fc} /* (10, 14, 9) {real, imag} */,
  {32'hbfb783ec, 32'hc0d2353c} /* (10, 14, 8) {real, imag} */,
  {32'h40935c66, 32'hc182a402} /* (10, 14, 7) {real, imag} */,
  {32'hc09ca25b, 32'hc1b16a7c} /* (10, 14, 6) {real, imag} */,
  {32'hc163cbfe, 32'hc167633b} /* (10, 14, 5) {real, imag} */,
  {32'h4009a3fc, 32'h41eb1616} /* (10, 14, 4) {real, imag} */,
  {32'h4197711e, 32'hbfb611d8} /* (10, 14, 3) {real, imag} */,
  {32'hc16c0720, 32'hbecea490} /* (10, 14, 2) {real, imag} */,
  {32'hc2093744, 32'h4227b199} /* (10, 14, 1) {real, imag} */,
  {32'hc16b68a6, 32'h4184c91a} /* (10, 14, 0) {real, imag} */,
  {32'h41d65675, 32'hc11ac424} /* (10, 13, 31) {real, imag} */,
  {32'h41a6b498, 32'hc0c74c0f} /* (10, 13, 30) {real, imag} */,
  {32'hc202a046, 32'hc132f8b8} /* (10, 13, 29) {real, imag} */,
  {32'hc18dd90b, 32'hc1a354ec} /* (10, 13, 28) {real, imag} */,
  {32'h41a89abf, 32'h40210344} /* (10, 13, 27) {real, imag} */,
  {32'h41113c64, 32'h415be47d} /* (10, 13, 26) {real, imag} */,
  {32'h412cabf8, 32'hc06aa304} /* (10, 13, 25) {real, imag} */,
  {32'hc14cbcf0, 32'hbcfa1100} /* (10, 13, 24) {real, imag} */,
  {32'h413eadde, 32'hc0a7c397} /* (10, 13, 23) {real, imag} */,
  {32'h3fba60c0, 32'h4079ce0c} /* (10, 13, 22) {real, imag} */,
  {32'hbe493690, 32'hbfa5abfa} /* (10, 13, 21) {real, imag} */,
  {32'hc140e8fe, 32'h418ee74a} /* (10, 13, 20) {real, imag} */,
  {32'h40ef03f9, 32'h40f90839} /* (10, 13, 19) {real, imag} */,
  {32'hc0e14a0c, 32'h415d7542} /* (10, 13, 18) {real, imag} */,
  {32'hbff0c7c4, 32'h400d9460} /* (10, 13, 17) {real, imag} */,
  {32'hc0746cb5, 32'hc158795e} /* (10, 13, 16) {real, imag} */,
  {32'h3ea7bcf0, 32'h4111d212} /* (10, 13, 15) {real, imag} */,
  {32'hc098c716, 32'hc07b2e4e} /* (10, 13, 14) {real, imag} */,
  {32'hc0e88c77, 32'hc0e1530f} /* (10, 13, 13) {real, imag} */,
  {32'h411d33de, 32'hbfa7e6a8} /* (10, 13, 12) {real, imag} */,
  {32'hc0ae4250, 32'h40e979a2} /* (10, 13, 11) {real, imag} */,
  {32'h418ce544, 32'hbf041d60} /* (10, 13, 10) {real, imag} */,
  {32'h3fd598a4, 32'h418578da} /* (10, 13, 9) {real, imag} */,
  {32'h40e79280, 32'hc086c6d7} /* (10, 13, 8) {real, imag} */,
  {32'h4149c79e, 32'h3ffeacc0} /* (10, 13, 7) {real, imag} */,
  {32'h4036cb72, 32'hbef69100} /* (10, 13, 6) {real, imag} */,
  {32'h41960cc5, 32'h416c1365} /* (10, 13, 5) {real, imag} */,
  {32'hc131a4a6, 32'h40700b64} /* (10, 13, 4) {real, imag} */,
  {32'h40e3026c, 32'h40fb14ef} /* (10, 13, 3) {real, imag} */,
  {32'h41426cc7, 32'hc056c966} /* (10, 13, 2) {real, imag} */,
  {32'hc11ebe8e, 32'hc1a5efdd} /* (10, 13, 1) {real, imag} */,
  {32'h4124906a, 32'h421b7734} /* (10, 13, 0) {real, imag} */,
  {32'h408662b8, 32'h420c5c7f} /* (10, 12, 31) {real, imag} */,
  {32'h420da722, 32'h4121d03c} /* (10, 12, 30) {real, imag} */,
  {32'h41ca170c, 32'h4129d38a} /* (10, 12, 29) {real, imag} */,
  {32'h4214a041, 32'hc0073d6f} /* (10, 12, 28) {real, imag} */,
  {32'hc192c47b, 32'h42376687} /* (10, 12, 27) {real, imag} */,
  {32'h414ae0e4, 32'hc122bd97} /* (10, 12, 26) {real, imag} */,
  {32'hc19ad65a, 32'h3da52700} /* (10, 12, 25) {real, imag} */,
  {32'hc1c22ed4, 32'hc202c722} /* (10, 12, 24) {real, imag} */,
  {32'h4124f23d, 32'h40b3e984} /* (10, 12, 23) {real, imag} */,
  {32'hc18335e7, 32'hbf57b110} /* (10, 12, 22) {real, imag} */,
  {32'hc1646191, 32'h40ead5f1} /* (10, 12, 21) {real, imag} */,
  {32'hbe9c2e00, 32'h40cb52da} /* (10, 12, 20) {real, imag} */,
  {32'h41481d85, 32'hc11e7d7a} /* (10, 12, 19) {real, imag} */,
  {32'h40996f1c, 32'h3dab5ac0} /* (10, 12, 18) {real, imag} */,
  {32'h3ef25de8, 32'hc09e926b} /* (10, 12, 17) {real, imag} */,
  {32'hc11848ee, 32'hbeb18c40} /* (10, 12, 16) {real, imag} */,
  {32'h3f177da4, 32'h414de58a} /* (10, 12, 15) {real, imag} */,
  {32'h4145bb6e, 32'hbfdb3db4} /* (10, 12, 14) {real, imag} */,
  {32'h412e09bb, 32'hc0cb0aaf} /* (10, 12, 13) {real, imag} */,
  {32'h40c30aec, 32'h3f3dee0c} /* (10, 12, 12) {real, imag} */,
  {32'h411af365, 32'hc06eaed2} /* (10, 12, 11) {real, imag} */,
  {32'h405a0180, 32'h41acbf78} /* (10, 12, 10) {real, imag} */,
  {32'h416023d3, 32'h41b5f409} /* (10, 12, 9) {real, imag} */,
  {32'h41170e2c, 32'hc204c510} /* (10, 12, 8) {real, imag} */,
  {32'h41d87586, 32'hc1ca890d} /* (10, 12, 7) {real, imag} */,
  {32'hc163add6, 32'h40c40ee2} /* (10, 12, 6) {real, imag} */,
  {32'hc263da6a, 32'h41bda6a2} /* (10, 12, 5) {real, imag} */,
  {32'hc130d02d, 32'hbca85b80} /* (10, 12, 4) {real, imag} */,
  {32'hc0904876, 32'h4108d8f0} /* (10, 12, 3) {real, imag} */,
  {32'h4202844e, 32'hc1223a8c} /* (10, 12, 2) {real, imag} */,
  {32'h402d642b, 32'hc2108dc7} /* (10, 12, 1) {real, imag} */,
  {32'hc23049f2, 32'h3e547e80} /* (10, 12, 0) {real, imag} */,
  {32'hbcff0080, 32'hc21d97e7} /* (10, 11, 31) {real, imag} */,
  {32'h3fe1e7f5, 32'hc26d233a} /* (10, 11, 30) {real, imag} */,
  {32'h42480be6, 32'h418f32e0} /* (10, 11, 29) {real, imag} */,
  {32'h400b6950, 32'hc25f0bf6} /* (10, 11, 28) {real, imag} */,
  {32'hc19c4626, 32'hc166a026} /* (10, 11, 27) {real, imag} */,
  {32'hc10b1c53, 32'h41fccad5} /* (10, 11, 26) {real, imag} */,
  {32'h4146973d, 32'h4099b56e} /* (10, 11, 25) {real, imag} */,
  {32'hc19166ba, 32'h422c6176} /* (10, 11, 24) {real, imag} */,
  {32'hc1a1e13c, 32'h414e305f} /* (10, 11, 23) {real, imag} */,
  {32'hc1f9a7e4, 32'h41c9b3f3} /* (10, 11, 22) {real, imag} */,
  {32'hc1ad1b2e, 32'hc18ddfed} /* (10, 11, 21) {real, imag} */,
  {32'h40031ba0, 32'hc1886313} /* (10, 11, 20) {real, imag} */,
  {32'h40f0928a, 32'hc08a5d80} /* (10, 11, 19) {real, imag} */,
  {32'hc0c5f3ae, 32'h413aaf0e} /* (10, 11, 18) {real, imag} */,
  {32'h40c50c58, 32'h408ad431} /* (10, 11, 17) {real, imag} */,
  {32'hc09bfff8, 32'hc124bf01} /* (10, 11, 16) {real, imag} */,
  {32'h4008e2e0, 32'hbfcb1724} /* (10, 11, 15) {real, imag} */,
  {32'hc0c3a4d6, 32'h3d28d600} /* (10, 11, 14) {real, imag} */,
  {32'h41334d0d, 32'hbf8e9cb6} /* (10, 11, 13) {real, imag} */,
  {32'h4055f040, 32'h4047a3d8} /* (10, 11, 12) {real, imag} */,
  {32'hc17ea705, 32'h41736052} /* (10, 11, 11) {real, imag} */,
  {32'hc128367b, 32'h40762538} /* (10, 11, 10) {real, imag} */,
  {32'hc179d600, 32'h412effbb} /* (10, 11, 9) {real, imag} */,
  {32'hc0a452f2, 32'h4275ec9e} /* (10, 11, 8) {real, imag} */,
  {32'hc0853b66, 32'hc20c39f7} /* (10, 11, 7) {real, imag} */,
  {32'h403c5c7c, 32'hc1d26c8b} /* (10, 11, 6) {real, imag} */,
  {32'hc00f8d2c, 32'h4231e0a4} /* (10, 11, 5) {real, imag} */,
  {32'hc2848b18, 32'hc0303238} /* (10, 11, 4) {real, imag} */,
  {32'hc252a1e0, 32'h40a3fa7e} /* (10, 11, 3) {real, imag} */,
  {32'h3faed53b, 32'h3ffdf630} /* (10, 11, 2) {real, imag} */,
  {32'hc007c589, 32'hc2121dad} /* (10, 11, 1) {real, imag} */,
  {32'hc1ebb2a8, 32'h411b2c15} /* (10, 11, 0) {real, imag} */,
  {32'h420427e9, 32'h41b81e56} /* (10, 10, 31) {real, imag} */,
  {32'h418e0c9a, 32'hc078dec0} /* (10, 10, 30) {real, imag} */,
  {32'h41ac73fb, 32'h418a376e} /* (10, 10, 29) {real, imag} */,
  {32'hc1b87ea4, 32'h41eb281c} /* (10, 10, 28) {real, imag} */,
  {32'h413012b8, 32'hc1eb84be} /* (10, 10, 27) {real, imag} */,
  {32'hc16b6f47, 32'hc1050dc2} /* (10, 10, 26) {real, imag} */,
  {32'h40b03890, 32'h40cd81b6} /* (10, 10, 25) {real, imag} */,
  {32'h41d6bf6c, 32'hc0a5bbce} /* (10, 10, 24) {real, imag} */,
  {32'h41e0e91b, 32'hc1eef1d6} /* (10, 10, 23) {real, imag} */,
  {32'h40439db4, 32'h4202d5e0} /* (10, 10, 22) {real, imag} */,
  {32'h41c4a43b, 32'h3ef90560} /* (10, 10, 21) {real, imag} */,
  {32'h4109c5f4, 32'hc13c7d89} /* (10, 10, 20) {real, imag} */,
  {32'h417cdb43, 32'h40f335f3} /* (10, 10, 19) {real, imag} */,
  {32'hc05a109e, 32'h41628796} /* (10, 10, 18) {real, imag} */,
  {32'h402630a6, 32'hc0d2848a} /* (10, 10, 17) {real, imag} */,
  {32'hc100e639, 32'hbf9672e0} /* (10, 10, 16) {real, imag} */,
  {32'h415dc0d2, 32'hc03b64d4} /* (10, 10, 15) {real, imag} */,
  {32'h3fbc4e9c, 32'h416a0c9a} /* (10, 10, 14) {real, imag} */,
  {32'h3f694830, 32'hc106cd80} /* (10, 10, 13) {real, imag} */,
  {32'h3f25f4fc, 32'hc126b9ed} /* (10, 10, 12) {real, imag} */,
  {32'h41c0c745, 32'hc16ec637} /* (10, 10, 11) {real, imag} */,
  {32'hc1dc55d4, 32'hc0b19d4a} /* (10, 10, 10) {real, imag} */,
  {32'hc1ca0c29, 32'hc15c6e19} /* (10, 10, 9) {real, imag} */,
  {32'hc02c20f0, 32'h41a8bc52} /* (10, 10, 8) {real, imag} */,
  {32'hc18f07e0, 32'hc1401637} /* (10, 10, 7) {real, imag} */,
  {32'h41c3dc9a, 32'h422fd7ae} /* (10, 10, 6) {real, imag} */,
  {32'hc0aee83c, 32'hc0f7817e} /* (10, 10, 5) {real, imag} */,
  {32'hc20f7d19, 32'hc266bfa6} /* (10, 10, 4) {real, imag} */,
  {32'h41d99759, 32'h40798e54} /* (10, 10, 3) {real, imag} */,
  {32'h41a9aea2, 32'hc1c20540} /* (10, 10, 2) {real, imag} */,
  {32'h4249f9b7, 32'hc1f54a88} /* (10, 10, 1) {real, imag} */,
  {32'hc174ec43, 32'h3f42f280} /* (10, 10, 0) {real, imag} */,
  {32'h4181205b, 32'h418c57de} /* (10, 9, 31) {real, imag} */,
  {32'hc211747e, 32'h41bcba78} /* (10, 9, 30) {real, imag} */,
  {32'h41119fda, 32'h4219c85b} /* (10, 9, 29) {real, imag} */,
  {32'hc12b9c7e, 32'h41525dcc} /* (10, 9, 28) {real, imag} */,
  {32'h41f343ab, 32'h4217cacf} /* (10, 9, 27) {real, imag} */,
  {32'hbf9c4840, 32'hc2053043} /* (10, 9, 26) {real, imag} */,
  {32'h40d02508, 32'hc0eb8fa8} /* (10, 9, 25) {real, imag} */,
  {32'h412644c6, 32'hbe53fc20} /* (10, 9, 24) {real, imag} */,
  {32'hc139f31a, 32'h41d448e0} /* (10, 9, 23) {real, imag} */,
  {32'hc1618dbb, 32'h420bbdd6} /* (10, 9, 22) {real, imag} */,
  {32'hc1856360, 32'hc0f953fb} /* (10, 9, 21) {real, imag} */,
  {32'hc1aa4c4f, 32'hc0fbe977} /* (10, 9, 20) {real, imag} */,
  {32'hc0ecd0a3, 32'h3fe4f91c} /* (10, 9, 19) {real, imag} */,
  {32'hc11e2a0f, 32'h404f8d90} /* (10, 9, 18) {real, imag} */,
  {32'hbf2c9590, 32'h4110eadc} /* (10, 9, 17) {real, imag} */,
  {32'hbf742bc8, 32'h412bf1ec} /* (10, 9, 16) {real, imag} */,
  {32'h40c4e116, 32'hbf1f86a0} /* (10, 9, 15) {real, imag} */,
  {32'hc0887236, 32'h3f8c3be0} /* (10, 9, 14) {real, imag} */,
  {32'hc1a8563d, 32'h4039f302} /* (10, 9, 13) {real, imag} */,
  {32'h4100f576, 32'h3f5c8dd8} /* (10, 9, 12) {real, imag} */,
  {32'h41030039, 32'hc16eac3e} /* (10, 9, 11) {real, imag} */,
  {32'h4136db93, 32'hc1e3bee8} /* (10, 9, 10) {real, imag} */,
  {32'h40280ea0, 32'h41f3e8a2} /* (10, 9, 9) {real, imag} */,
  {32'h424f4704, 32'h3fbdc564} /* (10, 9, 8) {real, imag} */,
  {32'h4223e2df, 32'h4244e624} /* (10, 9, 7) {real, imag} */,
  {32'h411af21a, 32'hc1855096} /* (10, 9, 6) {real, imag} */,
  {32'hc0f70274, 32'h41385918} /* (10, 9, 5) {real, imag} */,
  {32'h41c31cd7, 32'h41ad2412} /* (10, 9, 4) {real, imag} */,
  {32'h422ec116, 32'h41f3f9b1} /* (10, 9, 3) {real, imag} */,
  {32'hc09b86f4, 32'h42b132d8} /* (10, 9, 2) {real, imag} */,
  {32'hc2116038, 32'h4227f491} /* (10, 9, 1) {real, imag} */,
  {32'h3fee1034, 32'hc2429bde} /* (10, 9, 0) {real, imag} */,
  {32'hc106b42e, 32'h41558cdd} /* (10, 8, 31) {real, imag} */,
  {32'hc19d7a30, 32'h4203ec00} /* (10, 8, 30) {real, imag} */,
  {32'hc228e4a5, 32'h41a116b5} /* (10, 8, 29) {real, imag} */,
  {32'hc1fa7a53, 32'hc2236ca0} /* (10, 8, 28) {real, imag} */,
  {32'h4213f105, 32'hc100a5bb} /* (10, 8, 27) {real, imag} */,
  {32'hc26635fb, 32'hc191b4b9} /* (10, 8, 26) {real, imag} */,
  {32'hc2349aa7, 32'h40c9f7df} /* (10, 8, 25) {real, imag} */,
  {32'h41a2fa64, 32'h40565848} /* (10, 8, 24) {real, imag} */,
  {32'hc00e2b98, 32'h4110ff38} /* (10, 8, 23) {real, imag} */,
  {32'hc14caf3c, 32'hc0b816e6} /* (10, 8, 22) {real, imag} */,
  {32'h3f617b20, 32'h414759a1} /* (10, 8, 21) {real, imag} */,
  {32'hc1aafd3f, 32'h41819ec1} /* (10, 8, 20) {real, imag} */,
  {32'h3fadcf50, 32'hc1228071} /* (10, 8, 19) {real, imag} */,
  {32'h4129d326, 32'hc0a4edfc} /* (10, 8, 18) {real, imag} */,
  {32'h3f8a79c0, 32'hc14a68ee} /* (10, 8, 17) {real, imag} */,
  {32'h4145fd20, 32'h412cb7c2} /* (10, 8, 16) {real, imag} */,
  {32'h3fa93840, 32'h41049548} /* (10, 8, 15) {real, imag} */,
  {32'h41633baa, 32'hc18465c7} /* (10, 8, 14) {real, imag} */,
  {32'h4120d64e, 32'h4122e34f} /* (10, 8, 13) {real, imag} */,
  {32'hc1e4c20d, 32'h415613ce} /* (10, 8, 12) {real, imag} */,
  {32'h41e9962c, 32'hc04edc84} /* (10, 8, 11) {real, imag} */,
  {32'hbf88a95c, 32'hc08f9ed6} /* (10, 8, 10) {real, imag} */,
  {32'hc1f41b83, 32'hc184a1b3} /* (10, 8, 9) {real, imag} */,
  {32'hc0bc1fc8, 32'h423eec0c} /* (10, 8, 8) {real, imag} */,
  {32'h4287c4dc, 32'hc067d53a} /* (10, 8, 7) {real, imag} */,
  {32'h425d6051, 32'h41ccdb47} /* (10, 8, 6) {real, imag} */,
  {32'h41c447ee, 32'hc21426a3} /* (10, 8, 5) {real, imag} */,
  {32'h415ced36, 32'h4250f258} /* (10, 8, 4) {real, imag} */,
  {32'h427c06a7, 32'hc1c3508b} /* (10, 8, 3) {real, imag} */,
  {32'hc267cf06, 32'hc21714be} /* (10, 8, 2) {real, imag} */,
  {32'hc1977d43, 32'h41d895ce} /* (10, 8, 1) {real, imag} */,
  {32'h42aa4656, 32'hc1fb0e75} /* (10, 8, 0) {real, imag} */,
  {32'hc22280a4, 32'h42691d85} /* (10, 7, 31) {real, imag} */,
  {32'h41536437, 32'h42870005} /* (10, 7, 30) {real, imag} */,
  {32'hc20971e1, 32'h413f6956} /* (10, 7, 29) {real, imag} */,
  {32'h426e8b15, 32'h423a66e8} /* (10, 7, 28) {real, imag} */,
  {32'h421a6423, 32'h42484af1} /* (10, 7, 27) {real, imag} */,
  {32'h41615a82, 32'hc14a9b28} /* (10, 7, 26) {real, imag} */,
  {32'h42382fc4, 32'hc1c85fd2} /* (10, 7, 25) {real, imag} */,
  {32'h415addd7, 32'hc282ab1a} /* (10, 7, 24) {real, imag} */,
  {32'h41ab3bf7, 32'hc1f54726} /* (10, 7, 23) {real, imag} */,
  {32'h4003aaf4, 32'hc19fd4e8} /* (10, 7, 22) {real, imag} */,
  {32'hc0932dba, 32'hc1ba79ad} /* (10, 7, 21) {real, imag} */,
  {32'hc09f8a0c, 32'hc0f01ee5} /* (10, 7, 20) {real, imag} */,
  {32'hc0de0e68, 32'hc1c0e399} /* (10, 7, 19) {real, imag} */,
  {32'h40917570, 32'hc0145990} /* (10, 7, 18) {real, imag} */,
  {32'hc0a70490, 32'h41c02988} /* (10, 7, 17) {real, imag} */,
  {32'hc0545080, 32'hc1d8c94f} /* (10, 7, 16) {real, imag} */,
  {32'hc180f9ba, 32'h41095d58} /* (10, 7, 15) {real, imag} */,
  {32'h40436197, 32'hc1054784} /* (10, 7, 14) {real, imag} */,
  {32'h41d1deae, 32'hbdc70300} /* (10, 7, 13) {real, imag} */,
  {32'hc14bf5be, 32'h411365b4} /* (10, 7, 12) {real, imag} */,
  {32'h4165d371, 32'h412a6826} /* (10, 7, 11) {real, imag} */,
  {32'hc1d514c0, 32'hc247bc18} /* (10, 7, 10) {real, imag} */,
  {32'h41db64c7, 32'hc214caa3} /* (10, 7, 9) {real, imag} */,
  {32'hc188dd6a, 32'hc10a6770} /* (10, 7, 8) {real, imag} */,
  {32'hc1637b72, 32'h40ec7eda} /* (10, 7, 7) {real, imag} */,
  {32'h4192fa23, 32'hc250053a} /* (10, 7, 6) {real, imag} */,
  {32'h41821a78, 32'hc22367d3} /* (10, 7, 5) {real, imag} */,
  {32'h40f3f2f8, 32'hc1df32e5} /* (10, 7, 4) {real, imag} */,
  {32'hc15621a4, 32'h41f1f0d9} /* (10, 7, 3) {real, imag} */,
  {32'hc20fba36, 32'hc2a3d6ab} /* (10, 7, 2) {real, imag} */,
  {32'h410ecfe2, 32'hc29559f6} /* (10, 7, 1) {real, imag} */,
  {32'h422760ae, 32'hc23bd8f8} /* (10, 7, 0) {real, imag} */,
  {32'h42239bde, 32'hc1fa9943} /* (10, 6, 31) {real, imag} */,
  {32'h406b8e70, 32'h41f42eb8} /* (10, 6, 30) {real, imag} */,
  {32'hc2d90730, 32'hbf676b30} /* (10, 6, 29) {real, imag} */,
  {32'h429ad39d, 32'h40537b5c} /* (10, 6, 28) {real, imag} */,
  {32'hc0fbcaa0, 32'hc287a447} /* (10, 6, 27) {real, imag} */,
  {32'hc04cdb34, 32'hc10f85a2} /* (10, 6, 26) {real, imag} */,
  {32'h4092f6de, 32'hc11de7a4} /* (10, 6, 25) {real, imag} */,
  {32'h40b13e00, 32'h417d5120} /* (10, 6, 24) {real, imag} */,
  {32'h42370863, 32'hc212cd91} /* (10, 6, 23) {real, imag} */,
  {32'hc13ee720, 32'h427c5714} /* (10, 6, 22) {real, imag} */,
  {32'hbf91f4cc, 32'hc0c175e0} /* (10, 6, 21) {real, imag} */,
  {32'h41a15f80, 32'hbf8d39c8} /* (10, 6, 20) {real, imag} */,
  {32'hbfb538f8, 32'h419f7554} /* (10, 6, 19) {real, imag} */,
  {32'h3eb9b8c0, 32'hc1e5fcfa} /* (10, 6, 18) {real, imag} */,
  {32'hc0f05b14, 32'h4096e298} /* (10, 6, 17) {real, imag} */,
  {32'hc15ca9e6, 32'h402df9d0} /* (10, 6, 16) {real, imag} */,
  {32'hc1b07f57, 32'h4197784c} /* (10, 6, 15) {real, imag} */,
  {32'h3faa1110, 32'h4179907d} /* (10, 6, 14) {real, imag} */,
  {32'h40e4da32, 32'hc1b20aac} /* (10, 6, 13) {real, imag} */,
  {32'hbfe374f8, 32'h41944e68} /* (10, 6, 12) {real, imag} */,
  {32'hbf1a2058, 32'h4231cbbe} /* (10, 6, 11) {real, imag} */,
  {32'hc242fcb0, 32'hc1d18f4d} /* (10, 6, 10) {real, imag} */,
  {32'hc1b42806, 32'h3fc8ee20} /* (10, 6, 9) {real, imag} */,
  {32'h4293983f, 32'h41e4525a} /* (10, 6, 8) {real, imag} */,
  {32'h419b52cc, 32'hc25bf80d} /* (10, 6, 7) {real, imag} */,
  {32'h40e5309a, 32'h42103e16} /* (10, 6, 6) {real, imag} */,
  {32'hc1c011b6, 32'hc1d3b400} /* (10, 6, 5) {real, imag} */,
  {32'h40177be0, 32'h419297f0} /* (10, 6, 4) {real, imag} */,
  {32'h42429491, 32'h41f31ba6} /* (10, 6, 3) {real, imag} */,
  {32'hc2b6fe4c, 32'hc21750fc} /* (10, 6, 2) {real, imag} */,
  {32'h419ef180, 32'h42a3a889} /* (10, 6, 1) {real, imag} */,
  {32'hc28378f4, 32'hc2155d2e} /* (10, 6, 0) {real, imag} */,
  {32'hc2550e3e, 32'hc3087741} /* (10, 5, 31) {real, imag} */,
  {32'hc1882f77, 32'h426b7bf1} /* (10, 5, 30) {real, imag} */,
  {32'h4245214a, 32'h3f7a0440} /* (10, 5, 29) {real, imag} */,
  {32'hc17479dd, 32'hc1eadf90} /* (10, 5, 28) {real, imag} */,
  {32'hc281b62b, 32'hc1583bd9} /* (10, 5, 27) {real, imag} */,
  {32'h422b2aaf, 32'h424e778c} /* (10, 5, 26) {real, imag} */,
  {32'hbfdaf4a0, 32'hc12a619a} /* (10, 5, 25) {real, imag} */,
  {32'hc1e898e5, 32'hc1e068e9} /* (10, 5, 24) {real, imag} */,
  {32'h3dc35480, 32'h41c065cc} /* (10, 5, 23) {real, imag} */,
  {32'hc1b926d4, 32'h429e68fe} /* (10, 5, 22) {real, imag} */,
  {32'h4188cdd2, 32'hc14c2593} /* (10, 5, 21) {real, imag} */,
  {32'hbdf5e500, 32'h41620f92} /* (10, 5, 20) {real, imag} */,
  {32'hc0a1ddd8, 32'hc1855056} /* (10, 5, 19) {real, imag} */,
  {32'hc0992c3c, 32'hc185e202} /* (10, 5, 18) {real, imag} */,
  {32'h419371cb, 32'hc019a098} /* (10, 5, 17) {real, imag} */,
  {32'hc1445150, 32'hc037fe40} /* (10, 5, 16) {real, imag} */,
  {32'hc1764771, 32'h411bab2a} /* (10, 5, 15) {real, imag} */,
  {32'h41cf8022, 32'hc1537bdb} /* (10, 5, 14) {real, imag} */,
  {32'hc1b261f0, 32'hc1bc88f6} /* (10, 5, 13) {real, imag} */,
  {32'h4125ef1c, 32'h3f0d0ec0} /* (10, 5, 12) {real, imag} */,
  {32'hc129e554, 32'h42080e07} /* (10, 5, 11) {real, imag} */,
  {32'hc1bd15f4, 32'hc208eb68} /* (10, 5, 10) {real, imag} */,
  {32'h41c14280, 32'hbf68b0d0} /* (10, 5, 9) {real, imag} */,
  {32'hc09616fc, 32'hc1e5afb7} /* (10, 5, 8) {real, imag} */,
  {32'h429a1a78, 32'h40974130} /* (10, 5, 7) {real, imag} */,
  {32'hc22a8ed5, 32'h42615dcc} /* (10, 5, 6) {real, imag} */,
  {32'hc282dcf7, 32'h42293198} /* (10, 5, 5) {real, imag} */,
  {32'h42278745, 32'hc22278bc} /* (10, 5, 4) {real, imag} */,
  {32'h418dc034, 32'hc1ae18aa} /* (10, 5, 3) {real, imag} */,
  {32'h4034d640, 32'hc1eeb75a} /* (10, 5, 2) {real, imag} */,
  {32'h42613350, 32'h42b158f0} /* (10, 5, 1) {real, imag} */,
  {32'h42758348, 32'hc2a69388} /* (10, 5, 0) {real, imag} */,
  {32'h41454bb2, 32'hc0a29f20} /* (10, 4, 31) {real, imag} */,
  {32'h42b6b48c, 32'hc0336480} /* (10, 4, 30) {real, imag} */,
  {32'hc2b2c24d, 32'h42b1ba92} /* (10, 4, 29) {real, imag} */,
  {32'h42e15052, 32'h418f24e7} /* (10, 4, 28) {real, imag} */,
  {32'h41b9b61d, 32'h42052c3b} /* (10, 4, 27) {real, imag} */,
  {32'hc21d7e48, 32'h4239d4a8} /* (10, 4, 26) {real, imag} */,
  {32'h41e33702, 32'h41945709} /* (10, 4, 25) {real, imag} */,
  {32'hc1559636, 32'hc2b44b79} /* (10, 4, 24) {real, imag} */,
  {32'hc205f828, 32'hc22f2b8c} /* (10, 4, 23) {real, imag} */,
  {32'hc1d780ca, 32'hc26d0258} /* (10, 4, 22) {real, imag} */,
  {32'hc007c5b4, 32'hc11fc844} /* (10, 4, 21) {real, imag} */,
  {32'hc14dc63a, 32'h41c8881f} /* (10, 4, 20) {real, imag} */,
  {32'h4106f94a, 32'hc278084c} /* (10, 4, 19) {real, imag} */,
  {32'h41377230, 32'h41d0d431} /* (10, 4, 18) {real, imag} */,
  {32'h404a3ba8, 32'hc0145cf8} /* (10, 4, 17) {real, imag} */,
  {32'h400677c0, 32'hc06d4918} /* (10, 4, 16) {real, imag} */,
  {32'hc1cf5c5b, 32'h410a856e} /* (10, 4, 15) {real, imag} */,
  {32'h3f87b57c, 32'h41dad4a3} /* (10, 4, 14) {real, imag} */,
  {32'h4162ec06, 32'hc023ece0} /* (10, 4, 13) {real, imag} */,
  {32'hc09038dc, 32'h419a443f} /* (10, 4, 12) {real, imag} */,
  {32'hc1e66906, 32'h40c0a350} /* (10, 4, 11) {real, imag} */,
  {32'h415c9dd7, 32'h419c435b} /* (10, 4, 10) {real, imag} */,
  {32'hc07567b8, 32'hc25ee684} /* (10, 4, 9) {real, imag} */,
  {32'hc1af23b5, 32'hc1b6c24c} /* (10, 4, 8) {real, imag} */,
  {32'hc2b29ffe, 32'hc22a6db2} /* (10, 4, 7) {real, imag} */,
  {32'hc212f594, 32'h40bf120c} /* (10, 4, 6) {real, imag} */,
  {32'hc11dce5a, 32'hc2233435} /* (10, 4, 5) {real, imag} */,
  {32'hbfcbe620, 32'hc283a8aa} /* (10, 4, 4) {real, imag} */,
  {32'hc28a5d15, 32'h428f5e12} /* (10, 4, 3) {real, imag} */,
  {32'h42a52cbe, 32'h42331ebc} /* (10, 4, 2) {real, imag} */,
  {32'hc1f02df7, 32'hc302a482} /* (10, 4, 1) {real, imag} */,
  {32'hc2b27f32, 32'hc1cdc3bd} /* (10, 4, 0) {real, imag} */,
  {32'h425c489a, 32'h4274f3e6} /* (10, 3, 31) {real, imag} */,
  {32'h4315aa3e, 32'hbf00c4c0} /* (10, 3, 30) {real, imag} */,
  {32'h418168e1, 32'hc2a135f5} /* (10, 3, 29) {real, imag} */,
  {32'h4021b528, 32'h4210885d} /* (10, 3, 28) {real, imag} */,
  {32'h42846ba4, 32'hc26412c0} /* (10, 3, 27) {real, imag} */,
  {32'hc2192c0e, 32'h4280a9d5} /* (10, 3, 26) {real, imag} */,
  {32'h4181a697, 32'hc08b134e} /* (10, 3, 25) {real, imag} */,
  {32'h425089a7, 32'h42a0d266} /* (10, 3, 24) {real, imag} */,
  {32'hc1b290a9, 32'h42509d61} /* (10, 3, 23) {real, imag} */,
  {32'hc1ce76e4, 32'hc1095ebf} /* (10, 3, 22) {real, imag} */,
  {32'h40f676fa, 32'h400f1e20} /* (10, 3, 21) {real, imag} */,
  {32'hc22e5db8, 32'h4120ee5a} /* (10, 3, 20) {real, imag} */,
  {32'h416d8584, 32'h4206ef56} /* (10, 3, 19) {real, imag} */,
  {32'h4102062e, 32'h41d8a266} /* (10, 3, 18) {real, imag} */,
  {32'hc0bf3e58, 32'h3fd9d1c0} /* (10, 3, 17) {real, imag} */,
  {32'hc05ce8c8, 32'hc1483e6e} /* (10, 3, 16) {real, imag} */,
  {32'h3ff69a60, 32'hc10429f8} /* (10, 3, 15) {real, imag} */,
  {32'hc031f438, 32'h40d0cf70} /* (10, 3, 14) {real, imag} */,
  {32'hc16ef024, 32'hc1643f9e} /* (10, 3, 13) {real, imag} */,
  {32'h40bf46bc, 32'hc1226dee} /* (10, 3, 12) {real, imag} */,
  {32'h4186aeaa, 32'hc21a3a9c} /* (10, 3, 11) {real, imag} */,
  {32'hc1c328ce, 32'h41214275} /* (10, 3, 10) {real, imag} */,
  {32'hc18851f7, 32'hc20ff0c3} /* (10, 3, 9) {real, imag} */,
  {32'h41a9bc7a, 32'hc203e0e4} /* (10, 3, 8) {real, imag} */,
  {32'hc07a1098, 32'hc169a76b} /* (10, 3, 7) {real, imag} */,
  {32'h40eaaf6c, 32'hc22adc72} /* (10, 3, 6) {real, imag} */,
  {32'h4132e140, 32'h3e056e00} /* (10, 3, 5) {real, imag} */,
  {32'h41daf23d, 32'hc229383d} /* (10, 3, 4) {real, imag} */,
  {32'hc20df0be, 32'hc291166f} /* (10, 3, 3) {real, imag} */,
  {32'h42cf8d48, 32'h4273ff24} /* (10, 3, 2) {real, imag} */,
  {32'h41766df0, 32'h426fb12a} /* (10, 3, 1) {real, imag} */,
  {32'hc1cf0577, 32'hc11a2d76} /* (10, 3, 0) {real, imag} */,
  {32'h42fdb085, 32'h4156b2fc} /* (10, 2, 31) {real, imag} */,
  {32'hc31c4acf, 32'hc10cc4e2} /* (10, 2, 30) {real, imag} */,
  {32'hc2880bba, 32'hc2b8b4a8} /* (10, 2, 29) {real, imag} */,
  {32'h4260ba18, 32'hc250b834} /* (10, 2, 28) {real, imag} */,
  {32'hc1c36802, 32'h3f025230} /* (10, 2, 27) {real, imag} */,
  {32'hc1815051, 32'hc22b53b0} /* (10, 2, 26) {real, imag} */,
  {32'hc0a0d680, 32'hc0c991bc} /* (10, 2, 25) {real, imag} */,
  {32'h42f50c06, 32'hc23b3410} /* (10, 2, 24) {real, imag} */,
  {32'hc21b9f4a, 32'hc140a062} /* (10, 2, 23) {real, imag} */,
  {32'h428be256, 32'h422744c2} /* (10, 2, 22) {real, imag} */,
  {32'hbf3bf1a0, 32'hc0fcda50} /* (10, 2, 21) {real, imag} */,
  {32'hc1dc270c, 32'h417b77b4} /* (10, 2, 20) {real, imag} */,
  {32'hc1f3e268, 32'h41ea23e8} /* (10, 2, 19) {real, imag} */,
  {32'h419228b6, 32'hc1695271} /* (10, 2, 18) {real, imag} */,
  {32'hc2135aae, 32'hc053abb8} /* (10, 2, 17) {real, imag} */,
  {32'h41c45ad0, 32'hc012a208} /* (10, 2, 16) {real, imag} */,
  {32'h420d6406, 32'hc1d4abd3} /* (10, 2, 15) {real, imag} */,
  {32'hc2164c59, 32'h418250a2} /* (10, 2, 14) {real, imag} */,
  {32'hc0f42418, 32'h4232cb68} /* (10, 2, 13) {real, imag} */,
  {32'hc1470be1, 32'hc0e097f8} /* (10, 2, 12) {real, imag} */,
  {32'h4203aa3c, 32'hc2240c60} /* (10, 2, 11) {real, imag} */,
  {32'h418a5051, 32'h417179ce} /* (10, 2, 10) {real, imag} */,
  {32'hc1ec1908, 32'hc1b6d9f9} /* (10, 2, 9) {real, imag} */,
  {32'hc227cde4, 32'h42853e60} /* (10, 2, 8) {real, imag} */,
  {32'h426c5f0a, 32'hc21c05dc} /* (10, 2, 7) {real, imag} */,
  {32'h42595da2, 32'hc14cfa2a} /* (10, 2, 6) {real, imag} */,
  {32'hc287ec26, 32'h412e52a3} /* (10, 2, 5) {real, imag} */,
  {32'h402d23c0, 32'hc29c11ae} /* (10, 2, 4) {real, imag} */,
  {32'hc22eee2d, 32'h425692bc} /* (10, 2, 3) {real, imag} */,
  {32'hc2d83d7a, 32'hbfe02674} /* (10, 2, 2) {real, imag} */,
  {32'h429dd48d, 32'hc0a49e18} /* (10, 2, 1) {real, imag} */,
  {32'h42306348, 32'hc1519b82} /* (10, 2, 0) {real, imag} */,
  {32'hc2e15702, 32'h428210a5} /* (10, 1, 31) {real, imag} */,
  {32'h42a62adb, 32'h41a17841} /* (10, 1, 30) {real, imag} */,
  {32'h41ded948, 32'hc251b74e} /* (10, 1, 29) {real, imag} */,
  {32'hc1e5c135, 32'h42f88542} /* (10, 1, 28) {real, imag} */,
  {32'h42afb88a, 32'hc24c9250} /* (10, 1, 27) {real, imag} */,
  {32'h42cda2d8, 32'h42c31b7f} /* (10, 1, 26) {real, imag} */,
  {32'h4142e145, 32'hc199d975} /* (10, 1, 25) {real, imag} */,
  {32'h404d7658, 32'hc0fb3b14} /* (10, 1, 24) {real, imag} */,
  {32'hc0bbaa04, 32'h42049170} /* (10, 1, 23) {real, imag} */,
  {32'hc245066e, 32'h41c11247} /* (10, 1, 22) {real, imag} */,
  {32'h42453da6, 32'hc12022c2} /* (10, 1, 21) {real, imag} */,
  {32'h41870ba9, 32'h419b1774} /* (10, 1, 20) {real, imag} */,
  {32'h4187be62, 32'hbfb1ab40} /* (10, 1, 19) {real, imag} */,
  {32'hc00ba8f8, 32'hc0a37fa0} /* (10, 1, 18) {real, imag} */,
  {32'hc1c98537, 32'hc03372d8} /* (10, 1, 17) {real, imag} */,
  {32'hc1ac4fe1, 32'h41c6cf6f} /* (10, 1, 16) {real, imag} */,
  {32'h3f0443e0, 32'hc1dbb071} /* (10, 1, 15) {real, imag} */,
  {32'h40945a9c, 32'h42369011} /* (10, 1, 14) {real, imag} */,
  {32'hc120e439, 32'h3e77fe00} /* (10, 1, 13) {real, imag} */,
  {32'hc1952741, 32'h402faa60} /* (10, 1, 12) {real, imag} */,
  {32'h41dfce59, 32'h4248a61c} /* (10, 1, 11) {real, imag} */,
  {32'h3f630180, 32'h40d64d64} /* (10, 1, 10) {real, imag} */,
  {32'h42272078, 32'h419bdeed} /* (10, 1, 9) {real, imag} */,
  {32'hc212ba7a, 32'h407286e8} /* (10, 1, 8) {real, imag} */,
  {32'h41fb7ca8, 32'h41a43b1d} /* (10, 1, 7) {real, imag} */,
  {32'h4202f16f, 32'h422a7e2a} /* (10, 1, 6) {real, imag} */,
  {32'h41292ca4, 32'hc19961af} /* (10, 1, 5) {real, imag} */,
  {32'hc20cb128, 32'h421011a8} /* (10, 1, 4) {real, imag} */,
  {32'h425bbeb0, 32'h42a0d075} /* (10, 1, 3) {real, imag} */,
  {32'h42063bea, 32'hc2845d5a} /* (10, 1, 2) {real, imag} */,
  {32'hc32ee7ef, 32'hc25cd792} /* (10, 1, 1) {real, imag} */,
  {32'hc27fd99a, 32'h4241afb0} /* (10, 1, 0) {real, imag} */,
  {32'hc2264fce, 32'h41e251b4} /* (10, 0, 31) {real, imag} */,
  {32'hc0c18e54, 32'hc1d2c85d} /* (10, 0, 30) {real, imag} */,
  {32'hc29b8a06, 32'hc2521834} /* (10, 0, 29) {real, imag} */,
  {32'h42c040b0, 32'hc2e1f3ea} /* (10, 0, 28) {real, imag} */,
  {32'h432d08a2, 32'hc28add02} /* (10, 0, 27) {real, imag} */,
  {32'hc2671a2e, 32'hc2f255a4} /* (10, 0, 26) {real, imag} */,
  {32'h41d0ade6, 32'hc197bf08} /* (10, 0, 25) {real, imag} */,
  {32'hc17ffca0, 32'h41a35fee} /* (10, 0, 24) {real, imag} */,
  {32'h42bc53c4, 32'hc13c7650} /* (10, 0, 23) {real, imag} */,
  {32'hc16dab10, 32'h41ebb2a8} /* (10, 0, 22) {real, imag} */,
  {32'h42036ea2, 32'hc1b2d6fa} /* (10, 0, 21) {real, imag} */,
  {32'h420a140a, 32'h40d3bc64} /* (10, 0, 20) {real, imag} */,
  {32'hc1af0d72, 32'hc1e22765} /* (10, 0, 19) {real, imag} */,
  {32'hc10b6aa6, 32'hc0826d8c} /* (10, 0, 18) {real, imag} */,
  {32'h40d307f4, 32'hc1b31c8c} /* (10, 0, 17) {real, imag} */,
  {32'h41a17744, 32'h42255080} /* (10, 0, 16) {real, imag} */,
  {32'h413484f6, 32'h412d7a99} /* (10, 0, 15) {real, imag} */,
  {32'hc0ea7b9c, 32'hc19316d9} /* (10, 0, 14) {real, imag} */,
  {32'h408df0e6, 32'h4204f45e} /* (10, 0, 13) {real, imag} */,
  {32'h408af9cc, 32'hc19ba2e5} /* (10, 0, 12) {real, imag} */,
  {32'hc03e5118, 32'hc238861b} /* (10, 0, 11) {real, imag} */,
  {32'hc0baed68, 32'h40f1fe00} /* (10, 0, 10) {real, imag} */,
  {32'h4276b903, 32'h4268c0b0} /* (10, 0, 9) {real, imag} */,
  {32'hc2a0d834, 32'h422a0aea} /* (10, 0, 8) {real, imag} */,
  {32'hc23dd76f, 32'h42a52804} /* (10, 0, 7) {real, imag} */,
  {32'h4136cb56, 32'h40892ba0} /* (10, 0, 6) {real, imag} */,
  {32'hc1c942b4, 32'h42848356} /* (10, 0, 5) {real, imag} */,
  {32'hc124af6c, 32'h3f3be1c0} /* (10, 0, 4) {real, imag} */,
  {32'hc30bdca4, 32'hc10150be} /* (10, 0, 3) {real, imag} */,
  {32'h4245643a, 32'hc2a97762} /* (10, 0, 2) {real, imag} */,
  {32'hc2d0398b, 32'hc2cd5d5d} /* (10, 0, 1) {real, imag} */,
  {32'hc214a857, 32'hc212cb0c} /* (10, 0, 0) {real, imag} */,
  {32'hc2b98911, 32'h4338a2fc} /* (9, 31, 31) {real, imag} */,
  {32'hc1b55b5d, 32'hc2f72f4d} /* (9, 31, 30) {real, imag} */,
  {32'hc224c513, 32'h41111df0} /* (9, 31, 29) {real, imag} */,
  {32'hc1988370, 32'h4296735c} /* (9, 31, 28) {real, imag} */,
  {32'h42359c51, 32'h418d106a} /* (9, 31, 27) {real, imag} */,
  {32'hc2010847, 32'h41837184} /* (9, 31, 26) {real, imag} */,
  {32'h42528544, 32'hc1a4c572} /* (9, 31, 25) {real, imag} */,
  {32'hc1d997c0, 32'hc2b4196a} /* (9, 31, 24) {real, imag} */,
  {32'hc1695080, 32'h4291e97a} /* (9, 31, 23) {real, imag} */,
  {32'hc18f1224, 32'h4210b36e} /* (9, 31, 22) {real, imag} */,
  {32'h4224faaa, 32'hc2148a3c} /* (9, 31, 21) {real, imag} */,
  {32'h4128a015, 32'hc200716d} /* (9, 31, 20) {real, imag} */,
  {32'hc148344c, 32'h411e3da2} /* (9, 31, 19) {real, imag} */,
  {32'hc218a56d, 32'hc1c1dc4c} /* (9, 31, 18) {real, imag} */,
  {32'hbea6cb40, 32'hc0dcfdd2} /* (9, 31, 17) {real, imag} */,
  {32'h4202f15a, 32'h41b1b744} /* (9, 31, 16) {real, imag} */,
  {32'h41d88b71, 32'hc1ecb20c} /* (9, 31, 15) {real, imag} */,
  {32'h41918874, 32'hc15d5948} /* (9, 31, 14) {real, imag} */,
  {32'hc1c834fa, 32'hc1b04af7} /* (9, 31, 13) {real, imag} */,
  {32'h421eb594, 32'h40ac53c0} /* (9, 31, 12) {real, imag} */,
  {32'h427244b4, 32'h41947a1c} /* (9, 31, 11) {real, imag} */,
  {32'h413dd2f2, 32'h40968f54} /* (9, 31, 10) {real, imag} */,
  {32'h41ad5490, 32'hc22b3e9d} /* (9, 31, 9) {real, imag} */,
  {32'hc1e558d0, 32'hc1fe7ffa} /* (9, 31, 8) {real, imag} */,
  {32'h421c709c, 32'h422f771b} /* (9, 31, 7) {real, imag} */,
  {32'h415fa245, 32'hc01c27a2} /* (9, 31, 6) {real, imag} */,
  {32'h420ffc79, 32'hc22be735} /* (9, 31, 5) {real, imag} */,
  {32'hc2401b68, 32'h422333b4} /* (9, 31, 4) {real, imag} */,
  {32'h4296f5ba, 32'h428661b8} /* (9, 31, 3) {real, imag} */,
  {32'hc1451a0e, 32'h41ea00a4} /* (9, 31, 2) {real, imag} */,
  {32'hc299a83f, 32'h42d759fd} /* (9, 31, 1) {real, imag} */,
  {32'hc3016198, 32'h43068ac2} /* (9, 31, 0) {real, imag} */,
  {32'h42f3d57e, 32'h4286c258} /* (9, 30, 31) {real, imag} */,
  {32'hc250f278, 32'h4324d56e} /* (9, 30, 30) {real, imag} */,
  {32'h42105d86, 32'hc2bf6642} /* (9, 30, 29) {real, imag} */,
  {32'hc254e96e, 32'hc241d9e8} /* (9, 30, 28) {real, imag} */,
  {32'hc093b398, 32'hc2a75582} /* (9, 30, 27) {real, imag} */,
  {32'hc1af9100, 32'hc207bf7a} /* (9, 30, 26) {real, imag} */,
  {32'h4284728f, 32'hc1e1f310} /* (9, 30, 25) {real, imag} */,
  {32'h4208df36, 32'h42df697e} /* (9, 30, 24) {real, imag} */,
  {32'h420aeae9, 32'h41dfe238} /* (9, 30, 23) {real, imag} */,
  {32'hc20e0b4e, 32'h42190e6d} /* (9, 30, 22) {real, imag} */,
  {32'h415266f8, 32'h424ce4ab} /* (9, 30, 21) {real, imag} */,
  {32'h40439c0e, 32'h41e76a44} /* (9, 30, 20) {real, imag} */,
  {32'hc1cd3cb1, 32'hc1f8d4f4} /* (9, 30, 19) {real, imag} */,
  {32'hc11342fb, 32'hc10bc6aa} /* (9, 30, 18) {real, imag} */,
  {32'h414786f0, 32'h40f5cf9e} /* (9, 30, 17) {real, imag} */,
  {32'hc152d690, 32'hc0272ce0} /* (9, 30, 16) {real, imag} */,
  {32'h404f5e02, 32'hc1a9baac} /* (9, 30, 15) {real, imag} */,
  {32'hc0d3844a, 32'hc2039ad6} /* (9, 30, 14) {real, imag} */,
  {32'h4206c354, 32'h4029dea0} /* (9, 30, 13) {real, imag} */,
  {32'hc0302072, 32'h42277e64} /* (9, 30, 12) {real, imag} */,
  {32'hc127b754, 32'h428e8c93} /* (9, 30, 11) {real, imag} */,
  {32'h41e8bd14, 32'hc2682623} /* (9, 30, 10) {real, imag} */,
  {32'h41388534, 32'h41ea9f48} /* (9, 30, 9) {real, imag} */,
  {32'hc21cb670, 32'hc25f9877} /* (9, 30, 8) {real, imag} */,
  {32'h40e4e350, 32'hc2c26268} /* (9, 30, 7) {real, imag} */,
  {32'hc2f5b0e2, 32'h4266f61e} /* (9, 30, 6) {real, imag} */,
  {32'hc13eecd8, 32'hc234bad5} /* (9, 30, 5) {real, imag} */,
  {32'h42a41a1d, 32'h3f437b00} /* (9, 30, 4) {real, imag} */,
  {32'hc3099638, 32'h42767b21} /* (9, 30, 3) {real, imag} */,
  {32'hc2c55f78, 32'h42b5bc6b} /* (9, 30, 2) {real, imag} */,
  {32'h42fc1e3c, 32'hc2962f98} /* (9, 30, 1) {real, imag} */,
  {32'hc037fa00, 32'hc281ba82} /* (9, 30, 0) {real, imag} */,
  {32'hc1298a58, 32'h42c21fb0} /* (9, 29, 31) {real, imag} */,
  {32'hc309f91f, 32'hc308ffa8} /* (9, 29, 30) {real, imag} */,
  {32'h42a3012b, 32'h428e1ba2} /* (9, 29, 29) {real, imag} */,
  {32'h4041aee0, 32'h422d37e0} /* (9, 29, 28) {real, imag} */,
  {32'h41f901c2, 32'h428806d3} /* (9, 29, 27) {real, imag} */,
  {32'hc1ca6950, 32'h41d2a9df} /* (9, 29, 26) {real, imag} */,
  {32'h41f9445e, 32'h41c7b67a} /* (9, 29, 25) {real, imag} */,
  {32'hbea71100, 32'h424d8860} /* (9, 29, 24) {real, imag} */,
  {32'h41c20fe0, 32'h41f1319c} /* (9, 29, 23) {real, imag} */,
  {32'h421dabb0, 32'hc2031102} /* (9, 29, 22) {real, imag} */,
  {32'hc1f77378, 32'h42237a8a} /* (9, 29, 21) {real, imag} */,
  {32'hc1fe5622, 32'hc26bf5b3} /* (9, 29, 20) {real, imag} */,
  {32'hc1a27a06, 32'hc19a514b} /* (9, 29, 19) {real, imag} */,
  {32'h4111b210, 32'h41881cc2} /* (9, 29, 18) {real, imag} */,
  {32'hc0a12c06, 32'h411e077d} /* (9, 29, 17) {real, imag} */,
  {32'hc10dc17e, 32'hc04eb928} /* (9, 29, 16) {real, imag} */,
  {32'hc1e173a6, 32'hc16347eb} /* (9, 29, 15) {real, imag} */,
  {32'h41573b70, 32'h40c7b9f8} /* (9, 29, 14) {real, imag} */,
  {32'h4111c3b8, 32'h420407f6} /* (9, 29, 13) {real, imag} */,
  {32'h41c11508, 32'hc1fedbde} /* (9, 29, 12) {real, imag} */,
  {32'hc18f22a8, 32'h40426710} /* (9, 29, 11) {real, imag} */,
  {32'h427a3226, 32'h413ee1d4} /* (9, 29, 10) {real, imag} */,
  {32'hc15276d8, 32'hc1aab8d0} /* (9, 29, 9) {real, imag} */,
  {32'h42432f63, 32'hc255b97a} /* (9, 29, 8) {real, imag} */,
  {32'hc1950382, 32'h41c236f0} /* (9, 29, 7) {real, imag} */,
  {32'h412d0660, 32'h4222108c} /* (9, 29, 6) {real, imag} */,
  {32'h42a164ca, 32'h4278c792} /* (9, 29, 5) {real, imag} */,
  {32'hc295da43, 32'h41cf1944} /* (9, 29, 4) {real, imag} */,
  {32'hc0704160, 32'h41d15350} /* (9, 29, 3) {real, imag} */,
  {32'hc30ac511, 32'hc2abc953} /* (9, 29, 2) {real, imag} */,
  {32'hbf4a4b60, 32'hc301f7fe} /* (9, 29, 1) {real, imag} */,
  {32'hc01d2918, 32'h42862053} /* (9, 29, 0) {real, imag} */,
  {32'h42098e24, 32'hc24547c5} /* (9, 28, 31) {real, imag} */,
  {32'hc234dc7c, 32'h41f2b2f2} /* (9, 28, 30) {real, imag} */,
  {32'hc1638728, 32'h428485cf} /* (9, 28, 29) {real, imag} */,
  {32'h42647b98, 32'hc0bc3ff1} /* (9, 28, 28) {real, imag} */,
  {32'h42817acf, 32'hc27d665e} /* (9, 28, 27) {real, imag} */,
  {32'h4295df94, 32'hc2acf1ce} /* (9, 28, 26) {real, imag} */,
  {32'hc18fcb9a, 32'hc236a9d8} /* (9, 28, 25) {real, imag} */,
  {32'h4292f3e4, 32'hc22cfaea} /* (9, 28, 24) {real, imag} */,
  {32'h420194c1, 32'h41ff9d9f} /* (9, 28, 23) {real, imag} */,
  {32'h4203b9d1, 32'h40fddc6e} /* (9, 28, 22) {real, imag} */,
  {32'h400708a0, 32'hc1b3a2a6} /* (9, 28, 21) {real, imag} */,
  {32'h42346868, 32'h42074013} /* (9, 28, 20) {real, imag} */,
  {32'hc1b527e3, 32'h41c6e0fd} /* (9, 28, 19) {real, imag} */,
  {32'hc13ff77a, 32'h41d4d552} /* (9, 28, 18) {real, imag} */,
  {32'hc17fb606, 32'hc02386ec} /* (9, 28, 17) {real, imag} */,
  {32'h41991eff, 32'h41a9d768} /* (9, 28, 16) {real, imag} */,
  {32'h40813c8c, 32'hc192ebea} /* (9, 28, 15) {real, imag} */,
  {32'h41b1b88f, 32'h42226179} /* (9, 28, 14) {real, imag} */,
  {32'hc196aa4f, 32'hc1b40a83} /* (9, 28, 13) {real, imag} */,
  {32'hc0a29bb0, 32'hc0f51f9a} /* (9, 28, 12) {real, imag} */,
  {32'hc164e8c8, 32'h419b3af6} /* (9, 28, 11) {real, imag} */,
  {32'hc19a51f2, 32'hc1ffcc8e} /* (9, 28, 10) {real, imag} */,
  {32'hc20ac39b, 32'h416ad67a} /* (9, 28, 9) {real, imag} */,
  {32'hc304deb0, 32'hc218e6e6} /* (9, 28, 8) {real, imag} */,
  {32'h41a0c7ae, 32'hc20a5c70} /* (9, 28, 7) {real, imag} */,
  {32'h4208835b, 32'h41b7617a} /* (9, 28, 6) {real, imag} */,
  {32'hc1fc8599, 32'hc24b4a80} /* (9, 28, 5) {real, imag} */,
  {32'hc20f1f26, 32'h41196e5a} /* (9, 28, 4) {real, imag} */,
  {32'hc2742c4a, 32'h427d5122} /* (9, 28, 3) {real, imag} */,
  {32'hc23844d0, 32'hc2ae619e} /* (9, 28, 2) {real, imag} */,
  {32'h42582a12, 32'h42bd85e2} /* (9, 28, 1) {real, imag} */,
  {32'h41d3be15, 32'hc2bd329e} /* (9, 28, 0) {real, imag} */,
  {32'h427c5bfb, 32'hc2df11c0} /* (9, 27, 31) {real, imag} */,
  {32'hc27767c7, 32'h42510766} /* (9, 27, 30) {real, imag} */,
  {32'h428ba640, 32'hc1e0bbe1} /* (9, 27, 29) {real, imag} */,
  {32'h418d1405, 32'hc22f6dd0} /* (9, 27, 28) {real, imag} */,
  {32'h41e1306a, 32'h40d28e80} /* (9, 27, 27) {real, imag} */,
  {32'hc24fd236, 32'h4298151e} /* (9, 27, 26) {real, imag} */,
  {32'h424375ae, 32'hc2b5b906} /* (9, 27, 25) {real, imag} */,
  {32'hc19a9cc2, 32'hc2605998} /* (9, 27, 24) {real, imag} */,
  {32'hc1d8141e, 32'h428ca65a} /* (9, 27, 23) {real, imag} */,
  {32'h3f756680, 32'h428bef4e} /* (9, 27, 22) {real, imag} */,
  {32'h408ce71e, 32'h420f20f2} /* (9, 27, 21) {real, imag} */,
  {32'hc2526363, 32'hbf559440} /* (9, 27, 20) {real, imag} */,
  {32'h3f9a2d08, 32'h4144e99c} /* (9, 27, 19) {real, imag} */,
  {32'h3fdb8850, 32'hc12cdda3} /* (9, 27, 18) {real, imag} */,
  {32'h413e5e1d, 32'hc19bd404} /* (9, 27, 17) {real, imag} */,
  {32'hc17f35eb, 32'h417165fe} /* (9, 27, 16) {real, imag} */,
  {32'hbf549db0, 32'h4003b604} /* (9, 27, 15) {real, imag} */,
  {32'hc1af1419, 32'hc1d3205e} /* (9, 27, 14) {real, imag} */,
  {32'hc0dc147e, 32'hc166eed8} /* (9, 27, 13) {real, imag} */,
  {32'h416c8cfc, 32'hc0b685d0} /* (9, 27, 12) {real, imag} */,
  {32'hc1de654c, 32'hc102f82a} /* (9, 27, 11) {real, imag} */,
  {32'h41dc9e16, 32'hc281f12e} /* (9, 27, 10) {real, imag} */,
  {32'h42516011, 32'h4273fa24} /* (9, 27, 9) {real, imag} */,
  {32'h42867532, 32'h427392d0} /* (9, 27, 8) {real, imag} */,
  {32'h424d2168, 32'h4074fbc0} /* (9, 27, 7) {real, imag} */,
  {32'hc20e5be2, 32'h4290934e} /* (9, 27, 6) {real, imag} */,
  {32'h3f260630, 32'h4271aef8} /* (9, 27, 5) {real, imag} */,
  {32'hc11acf14, 32'hc1a5c4a0} /* (9, 27, 4) {real, imag} */,
  {32'hc2a61a4c, 32'h42265f88} /* (9, 27, 3) {real, imag} */,
  {32'h42523c29, 32'h425cb15e} /* (9, 27, 2) {real, imag} */,
  {32'hc205c89f, 32'hc22553df} /* (9, 27, 1) {real, imag} */,
  {32'h41c49a8a, 32'h421526b2} /* (9, 27, 0) {real, imag} */,
  {32'hc28b4a7f, 32'hc29ad133} /* (9, 26, 31) {real, imag} */,
  {32'h4240d117, 32'hc1acd8a0} /* (9, 26, 30) {real, imag} */,
  {32'h425fd3d3, 32'hc32b0b6c} /* (9, 26, 29) {real, imag} */,
  {32'h426da83f, 32'h409fc298} /* (9, 26, 28) {real, imag} */,
  {32'hc207552e, 32'h4178966e} /* (9, 26, 27) {real, imag} */,
  {32'h413e39fc, 32'hc1ca9e8a} /* (9, 26, 26) {real, imag} */,
  {32'h41ca9ac0, 32'hbf2f08e0} /* (9, 26, 25) {real, imag} */,
  {32'hc0f4738b, 32'h41dc300c} /* (9, 26, 24) {real, imag} */,
  {32'h423a447e, 32'h4202dee4} /* (9, 26, 23) {real, imag} */,
  {32'hbfedfa40, 32'hc206ee77} /* (9, 26, 22) {real, imag} */,
  {32'h408047da, 32'h425b990e} /* (9, 26, 21) {real, imag} */,
  {32'hc1a535cc, 32'hc214447c} /* (9, 26, 20) {real, imag} */,
  {32'hc10a3200, 32'hc114eaa0} /* (9, 26, 19) {real, imag} */,
  {32'hc1e2b7f6, 32'hc1bc3aee} /* (9, 26, 18) {real, imag} */,
  {32'hc194cc24, 32'h4008f960} /* (9, 26, 17) {real, imag} */,
  {32'hc14d876c, 32'hc192b09b} /* (9, 26, 16) {real, imag} */,
  {32'h42291546, 32'hc190718a} /* (9, 26, 15) {real, imag} */,
  {32'hc067b2b8, 32'hc10f7c81} /* (9, 26, 14) {real, imag} */,
  {32'hc0c3dcb1, 32'h4016b080} /* (9, 26, 13) {real, imag} */,
  {32'h418d2b6c, 32'h416e98c2} /* (9, 26, 12) {real, imag} */,
  {32'h4121f25b, 32'h41ef0a9d} /* (9, 26, 11) {real, imag} */,
  {32'hc261d9f6, 32'hc29c26ea} /* (9, 26, 10) {real, imag} */,
  {32'h41c3e03c, 32'h3e65cc80} /* (9, 26, 9) {real, imag} */,
  {32'hc132708e, 32'hc2537f5c} /* (9, 26, 8) {real, imag} */,
  {32'h413a48a1, 32'h423aac26} /* (9, 26, 7) {real, imag} */,
  {32'hc2457413, 32'h424cb13d} /* (9, 26, 6) {real, imag} */,
  {32'hc2acda34, 32'h4167050c} /* (9, 26, 5) {real, imag} */,
  {32'h4244bedd, 32'h4295fc38} /* (9, 26, 4) {real, imag} */,
  {32'hc29d4b2a, 32'hc1050ea0} /* (9, 26, 3) {real, imag} */,
  {32'hc1d49b7a, 32'h410900cd} /* (9, 26, 2) {real, imag} */,
  {32'h429cd4a9, 32'h418aa8a5} /* (9, 26, 1) {real, imag} */,
  {32'hc2620ed5, 32'hc11a268a} /* (9, 26, 0) {real, imag} */,
  {32'h4238df59, 32'hc1f28f0a} /* (9, 25, 31) {real, imag} */,
  {32'h40b6ee62, 32'hc2a65d63} /* (9, 25, 30) {real, imag} */,
  {32'hbfe3eca0, 32'h409f1168} /* (9, 25, 29) {real, imag} */,
  {32'h41b0b21b, 32'h41c4bdae} /* (9, 25, 28) {real, imag} */,
  {32'hc1f17a9c, 32'h427a9bed} /* (9, 25, 27) {real, imag} */,
  {32'hc27aea9e, 32'h41d729d5} /* (9, 25, 26) {real, imag} */,
  {32'hc1898508, 32'h41451207} /* (9, 25, 25) {real, imag} */,
  {32'h41f76c67, 32'hc15be764} /* (9, 25, 24) {real, imag} */,
  {32'hc1fd45c4, 32'h40a96c0c} /* (9, 25, 23) {real, imag} */,
  {32'hc21494bc, 32'h422e675b} /* (9, 25, 22) {real, imag} */,
  {32'hc1e92366, 32'hc202910d} /* (9, 25, 21) {real, imag} */,
  {32'hbe430440, 32'h3fa0e1b8} /* (9, 25, 20) {real, imag} */,
  {32'hc174df8f, 32'hc1e34990} /* (9, 25, 19) {real, imag} */,
  {32'h417ad4a5, 32'h40bd5cea} /* (9, 25, 18) {real, imag} */,
  {32'h419c9b71, 32'h4161d864} /* (9, 25, 17) {real, imag} */,
  {32'h4115631f, 32'hc156cf10} /* (9, 25, 16) {real, imag} */,
  {32'hc11cf8c6, 32'h40590510} /* (9, 25, 15) {real, imag} */,
  {32'h4091f086, 32'hc1527b75} /* (9, 25, 14) {real, imag} */,
  {32'h4076ff5c, 32'hc179881f} /* (9, 25, 13) {real, imag} */,
  {32'hc10ec02d, 32'hc0e445ce} /* (9, 25, 12) {real, imag} */,
  {32'hc1bc3ea0, 32'hc0a94338} /* (9, 25, 11) {real, imag} */,
  {32'hc23d3774, 32'h41f7bc75} /* (9, 25, 10) {real, imag} */,
  {32'hc1e263cc, 32'h41cfab30} /* (9, 25, 9) {real, imag} */,
  {32'h42142acb, 32'h42029231} /* (9, 25, 8) {real, imag} */,
  {32'h417b99c5, 32'h41e70f30} /* (9, 25, 7) {real, imag} */,
  {32'hc274880a, 32'h40488638} /* (9, 25, 6) {real, imag} */,
  {32'h42c73e97, 32'hc3060a73} /* (9, 25, 5) {real, imag} */,
  {32'h41e4cb45, 32'hc1d3a276} /* (9, 25, 4) {real, imag} */,
  {32'h4222a6e3, 32'hc22e5377} /* (9, 25, 3) {real, imag} */,
  {32'h4151a897, 32'hc20e3306} /* (9, 25, 2) {real, imag} */,
  {32'h420e93eb, 32'h42fc37da} /* (9, 25, 1) {real, imag} */,
  {32'h41ba8fbc, 32'hc16b8268} /* (9, 25, 0) {real, imag} */,
  {32'h401d9460, 32'h42774e02} /* (9, 24, 31) {real, imag} */,
  {32'hc222355e, 32'h41f744f7} /* (9, 24, 30) {real, imag} */,
  {32'hc1b1ee86, 32'hc1c9a136} /* (9, 24, 29) {real, imag} */,
  {32'hc1b2230e, 32'h421bccf0} /* (9, 24, 28) {real, imag} */,
  {32'h4204a51f, 32'hc29c4b86} /* (9, 24, 27) {real, imag} */,
  {32'hc20ab70c, 32'hc215abe6} /* (9, 24, 26) {real, imag} */,
  {32'hc1e92e5b, 32'h42269939} /* (9, 24, 25) {real, imag} */,
  {32'h42334e18, 32'hc11cbf17} /* (9, 24, 24) {real, imag} */,
  {32'hc16aac29, 32'hc13035b3} /* (9, 24, 23) {real, imag} */,
  {32'h40a643f4, 32'hc1eb8c39} /* (9, 24, 22) {real, imag} */,
  {32'h3fd46964, 32'hc0d906a8} /* (9, 24, 21) {real, imag} */,
  {32'hc00430d0, 32'h41e3e972} /* (9, 24, 20) {real, imag} */,
  {32'h4117afbf, 32'h41218854} /* (9, 24, 19) {real, imag} */,
  {32'h41cd3cfc, 32'hc088d2f5} /* (9, 24, 18) {real, imag} */,
  {32'hc0abe648, 32'hbe270140} /* (9, 24, 17) {real, imag} */,
  {32'hc0a8835a, 32'h41a308c4} /* (9, 24, 16) {real, imag} */,
  {32'hc0c591c4, 32'hc19d7acc} /* (9, 24, 15) {real, imag} */,
  {32'h415d27e3, 32'h40f0bbe5} /* (9, 24, 14) {real, imag} */,
  {32'h4173f5d9, 32'h420dee07} /* (9, 24, 13) {real, imag} */,
  {32'hbec2fa80, 32'hc20186a9} /* (9, 24, 12) {real, imag} */,
  {32'hbf01d208, 32'hc21a2a87} /* (9, 24, 11) {real, imag} */,
  {32'h4217218c, 32'hc097cbc4} /* (9, 24, 10) {real, imag} */,
  {32'h4196581e, 32'h41be7578} /* (9, 24, 9) {real, imag} */,
  {32'hc1ca3229, 32'h4214720e} /* (9, 24, 8) {real, imag} */,
  {32'hc0ac1214, 32'h419dc482} /* (9, 24, 7) {real, imag} */,
  {32'hc0b9a308, 32'h40959c34} /* (9, 24, 6) {real, imag} */,
  {32'h40f6cb00, 32'h4274442c} /* (9, 24, 5) {real, imag} */,
  {32'h42944bc0, 32'hc18f0918} /* (9, 24, 4) {real, imag} */,
  {32'hc1422650, 32'hc176c234} /* (9, 24, 3) {real, imag} */,
  {32'hc127df2d, 32'h425fd60e} /* (9, 24, 2) {real, imag} */,
  {32'h419f753d, 32'hc11ada96} /* (9, 24, 1) {real, imag} */,
  {32'hc1b74118, 32'hc28d3099} /* (9, 24, 0) {real, imag} */,
  {32'hc2817d8c, 32'hc2d67fe4} /* (9, 23, 31) {real, imag} */,
  {32'h41a955e4, 32'hc11cbd25} /* (9, 23, 30) {real, imag} */,
  {32'hc0afcd94, 32'hc19c62c7} /* (9, 23, 29) {real, imag} */,
  {32'h41ba2ea2, 32'h41a89343} /* (9, 23, 28) {real, imag} */,
  {32'hc1b79975, 32'hbf002d20} /* (9, 23, 27) {real, imag} */,
  {32'h4191aad7, 32'h422c126c} /* (9, 23, 26) {real, imag} */,
  {32'hc1f57ead, 32'h41b32fca} /* (9, 23, 25) {real, imag} */,
  {32'hc12a89d4, 32'hc117fb64} /* (9, 23, 24) {real, imag} */,
  {32'hc18fb27e, 32'h3fae95c8} /* (9, 23, 23) {real, imag} */,
  {32'hc140e380, 32'hc149942e} /* (9, 23, 22) {real, imag} */,
  {32'hc1b13a2f, 32'h41064b56} /* (9, 23, 21) {real, imag} */,
  {32'h414f1cb0, 32'hc16b9818} /* (9, 23, 20) {real, imag} */,
  {32'hc187e1c0, 32'h410d92eb} /* (9, 23, 19) {real, imag} */,
  {32'hc11e367b, 32'h405ca37c} /* (9, 23, 18) {real, imag} */,
  {32'h4168d9b4, 32'hc022f664} /* (9, 23, 17) {real, imag} */,
  {32'h40537136, 32'h40283700} /* (9, 23, 16) {real, imag} */,
  {32'hc0c2bd34, 32'hc0875402} /* (9, 23, 15) {real, imag} */,
  {32'hc123a95f, 32'h4056159c} /* (9, 23, 14) {real, imag} */,
  {32'h418b40fc, 32'hc110d9fd} /* (9, 23, 13) {real, imag} */,
  {32'hc1846c5b, 32'h40072c30} /* (9, 23, 12) {real, imag} */,
  {32'hc15fabc2, 32'h4125ea26} /* (9, 23, 11) {real, imag} */,
  {32'hc1a035f8, 32'h41aa2ca9} /* (9, 23, 10) {real, imag} */,
  {32'hc1e66fbc, 32'h40b24b42} /* (9, 23, 9) {real, imag} */,
  {32'h42ae1668, 32'hc130215c} /* (9, 23, 8) {real, imag} */,
  {32'h401774f8, 32'hc16d368f} /* (9, 23, 7) {real, imag} */,
  {32'h420e8eec, 32'h414878bd} /* (9, 23, 6) {real, imag} */,
  {32'h420fa1be, 32'h41c0e679} /* (9, 23, 5) {real, imag} */,
  {32'hc1d98cea, 32'h42a87f9f} /* (9, 23, 4) {real, imag} */,
  {32'h40da646c, 32'hc19ba2f1} /* (9, 23, 3) {real, imag} */,
  {32'hc1804e2e, 32'hc129b279} /* (9, 23, 2) {real, imag} */,
  {32'h41896506, 32'h425ed6c7} /* (9, 23, 1) {real, imag} */,
  {32'h41561a1a, 32'h412896bc} /* (9, 23, 0) {real, imag} */,
  {32'hc207c805, 32'h426171aa} /* (9, 22, 31) {real, imag} */,
  {32'hc0a98903, 32'hc29ac105} /* (9, 22, 30) {real, imag} */,
  {32'hc1b9063e, 32'h415b38b4} /* (9, 22, 29) {real, imag} */,
  {32'h409c52af, 32'h423dc0b0} /* (9, 22, 28) {real, imag} */,
  {32'h411481fe, 32'h41c02307} /* (9, 22, 27) {real, imag} */,
  {32'h4215b7fd, 32'hc0003790} /* (9, 22, 26) {real, imag} */,
  {32'hc26fc683, 32'h41da2904} /* (9, 22, 25) {real, imag} */,
  {32'hc1c93ca8, 32'h41952110} /* (9, 22, 24) {real, imag} */,
  {32'h4100b895, 32'hc1b00aef} /* (9, 22, 23) {real, imag} */,
  {32'h410a8986, 32'hc1050fb4} /* (9, 22, 22) {real, imag} */,
  {32'hc1139b3d, 32'hbf89aa30} /* (9, 22, 21) {real, imag} */,
  {32'h41e1d95d, 32'hc1638b8e} /* (9, 22, 20) {real, imag} */,
  {32'hbfcc1528, 32'hc17807f5} /* (9, 22, 19) {real, imag} */,
  {32'hc0bd1df5, 32'h40143d50} /* (9, 22, 18) {real, imag} */,
  {32'h3dfa3400, 32'hbd7b3380} /* (9, 22, 17) {real, imag} */,
  {32'h3d9e0a80, 32'h41526b2a} /* (9, 22, 16) {real, imag} */,
  {32'hc0535690, 32'h404a9ef2} /* (9, 22, 15) {real, imag} */,
  {32'h3f0c7d58, 32'hc0e11c30} /* (9, 22, 14) {real, imag} */,
  {32'hc0e8db5a, 32'hc1d9b0aa} /* (9, 22, 13) {real, imag} */,
  {32'h4151e7ae, 32'hc119f0c2} /* (9, 22, 12) {real, imag} */,
  {32'h41af6d94, 32'h417485d4} /* (9, 22, 11) {real, imag} */,
  {32'h4097d5dc, 32'hc1a67d44} /* (9, 22, 10) {real, imag} */,
  {32'h40cf5e62, 32'h41e17741} /* (9, 22, 9) {real, imag} */,
  {32'hc144da2f, 32'hc095d120} /* (9, 22, 8) {real, imag} */,
  {32'h417ba254, 32'hc08c83f6} /* (9, 22, 7) {real, imag} */,
  {32'h414743ff, 32'h42473cf0} /* (9, 22, 6) {real, imag} */,
  {32'h40333ece, 32'h41a67419} /* (9, 22, 5) {real, imag} */,
  {32'h410f2024, 32'hc29608ca} /* (9, 22, 4) {real, imag} */,
  {32'h4210f10f, 32'hbf70d560} /* (9, 22, 3) {real, imag} */,
  {32'h40a0648d, 32'h40aa73d0} /* (9, 22, 2) {real, imag} */,
  {32'h41fed8c6, 32'hc1f68e2c} /* (9, 22, 1) {real, imag} */,
  {32'h41584c6d, 32'h40439240} /* (9, 22, 0) {real, imag} */,
  {32'hc1ca62c0, 32'h4177f0b0} /* (9, 21, 31) {real, imag} */,
  {32'h41a3e4cd, 32'hc21f066b} /* (9, 21, 30) {real, imag} */,
  {32'hc12f00b4, 32'h421b303a} /* (9, 21, 29) {real, imag} */,
  {32'hc144e53a, 32'hc232d581} /* (9, 21, 28) {real, imag} */,
  {32'hc137b400, 32'h41f2b006} /* (9, 21, 27) {real, imag} */,
  {32'h426220fc, 32'hc2061bf9} /* (9, 21, 26) {real, imag} */,
  {32'h4213d34c, 32'h41745279} /* (9, 21, 25) {real, imag} */,
  {32'h3e532050, 32'h4141804a} /* (9, 21, 24) {real, imag} */,
  {32'hc0a0b818, 32'hc0857528} /* (9, 21, 23) {real, imag} */,
  {32'hbed7fce0, 32'h4155ec4c} /* (9, 21, 22) {real, imag} */,
  {32'hc0f8d2e0, 32'h40a96b36} /* (9, 21, 21) {real, imag} */,
  {32'hc11ff7c8, 32'h40601f53} /* (9, 21, 20) {real, imag} */,
  {32'hc0ab96f6, 32'h4181d58c} /* (9, 21, 19) {real, imag} */,
  {32'h4191c61f, 32'hc0a299e5} /* (9, 21, 18) {real, imag} */,
  {32'h40831dce, 32'h40d7a449} /* (9, 21, 17) {real, imag} */,
  {32'h3e277f80, 32'hc01d87f0} /* (9, 21, 16) {real, imag} */,
  {32'h3de5f160, 32'hc080f0ff} /* (9, 21, 15) {real, imag} */,
  {32'hc09b0ceb, 32'hbf874b14} /* (9, 21, 14) {real, imag} */,
  {32'hc057d628, 32'h3f617bf0} /* (9, 21, 13) {real, imag} */,
  {32'h41346020, 32'h40b9ea56} /* (9, 21, 12) {real, imag} */,
  {32'h41833766, 32'h413cad23} /* (9, 21, 11) {real, imag} */,
  {32'hc10bb725, 32'h4182b8c6} /* (9, 21, 10) {real, imag} */,
  {32'hc22edbca, 32'h401fa617} /* (9, 21, 9) {real, imag} */,
  {32'h40a00744, 32'h4187408f} /* (9, 21, 8) {real, imag} */,
  {32'h40f425d6, 32'hc1404ebd} /* (9, 21, 7) {real, imag} */,
  {32'h40e1709c, 32'hc236887f} /* (9, 21, 6) {real, imag} */,
  {32'h424be90d, 32'h40dc1e9a} /* (9, 21, 5) {real, imag} */,
  {32'hc22a08a4, 32'hc1ff76ea} /* (9, 21, 4) {real, imag} */,
  {32'hbfbf093c, 32'hc11339c8} /* (9, 21, 3) {real, imag} */,
  {32'h419d703b, 32'h41dc2bee} /* (9, 21, 2) {real, imag} */,
  {32'h4112e78b, 32'hc0cf12c7} /* (9, 21, 1) {real, imag} */,
  {32'h41907abd, 32'h41c25506} /* (9, 21, 0) {real, imag} */,
  {32'h4121a11e, 32'h40b65b04} /* (9, 20, 31) {real, imag} */,
  {32'h41b5a816, 32'h4141dc0e} /* (9, 20, 30) {real, imag} */,
  {32'h41aca749, 32'hc1518e78} /* (9, 20, 29) {real, imag} */,
  {32'h41863268, 32'h4162db8e} /* (9, 20, 28) {real, imag} */,
  {32'hc1e0e352, 32'hc06edb0e} /* (9, 20, 27) {real, imag} */,
  {32'h408d628f, 32'hc09e3398} /* (9, 20, 26) {real, imag} */,
  {32'h40e38722, 32'h422e3f24} /* (9, 20, 25) {real, imag} */,
  {32'hc18fdac4, 32'hbfef5724} /* (9, 20, 24) {real, imag} */,
  {32'hc20cf01f, 32'h405e95f8} /* (9, 20, 23) {real, imag} */,
  {32'hc0aa4182, 32'h40ade538} /* (9, 20, 22) {real, imag} */,
  {32'hc13ebf48, 32'hbdef7400} /* (9, 20, 21) {real, imag} */,
  {32'h411beb84, 32'hc1e4fc4a} /* (9, 20, 20) {real, imag} */,
  {32'h40878105, 32'h4170c754} /* (9, 20, 19) {real, imag} */,
  {32'h409c198c, 32'hc10cc531} /* (9, 20, 18) {real, imag} */,
  {32'h40210c8a, 32'h40562028} /* (9, 20, 17) {real, imag} */,
  {32'hbff71d20, 32'h40b5d6e1} /* (9, 20, 16) {real, imag} */,
  {32'hc05b1e5e, 32'h4050d0f8} /* (9, 20, 15) {real, imag} */,
  {32'hc0496668, 32'h4126b08f} /* (9, 20, 14) {real, imag} */,
  {32'h410a610e, 32'h3fc9e67c} /* (9, 20, 13) {real, imag} */,
  {32'hc058e316, 32'h40f8a5e8} /* (9, 20, 12) {real, imag} */,
  {32'hc1885942, 32'h41996d7c} /* (9, 20, 11) {real, imag} */,
  {32'h41603907, 32'hc1292a2c} /* (9, 20, 10) {real, imag} */,
  {32'hc18c83dc, 32'hc1495e5e} /* (9, 20, 9) {real, imag} */,
  {32'h41988f6c, 32'hc14468d4} /* (9, 20, 8) {real, imag} */,
  {32'hc1924782, 32'hc0edf8bc} /* (9, 20, 7) {real, imag} */,
  {32'h418315c2, 32'hc2020ab3} /* (9, 20, 6) {real, imag} */,
  {32'h409fb9f0, 32'h3f588f18} /* (9, 20, 5) {real, imag} */,
  {32'h4155ee32, 32'h418c8707} /* (9, 20, 4) {real, imag} */,
  {32'hc2047b78, 32'hc20b4c65} /* (9, 20, 3) {real, imag} */,
  {32'hc1ca7a1a, 32'hc15d3e12} /* (9, 20, 2) {real, imag} */,
  {32'h40b4f889, 32'hc1dad4f9} /* (9, 20, 1) {real, imag} */,
  {32'h41b4fe36, 32'h40753882} /* (9, 20, 0) {real, imag} */,
  {32'hbe4c3740, 32'hc1051722} /* (9, 19, 31) {real, imag} */,
  {32'hc149f5dc, 32'h40732ad8} /* (9, 19, 30) {real, imag} */,
  {32'h41445959, 32'hc1696240} /* (9, 19, 29) {real, imag} */,
  {32'hc1d3d4ac, 32'h40aff9a0} /* (9, 19, 28) {real, imag} */,
  {32'h413abd99, 32'h41e534f1} /* (9, 19, 27) {real, imag} */,
  {32'hbf3e1da0, 32'h40f9f576} /* (9, 19, 26) {real, imag} */,
  {32'h416e1213, 32'h40e69966} /* (9, 19, 25) {real, imag} */,
  {32'h41db150a, 32'h415a4897} /* (9, 19, 24) {real, imag} */,
  {32'hc08cdbb0, 32'hc106e4e8} /* (9, 19, 23) {real, imag} */,
  {32'hc15ddd80, 32'h402698bc} /* (9, 19, 22) {real, imag} */,
  {32'hc162e0a8, 32'h4008728c} /* (9, 19, 21) {real, imag} */,
  {32'h40fcdb4c, 32'hc1721faa} /* (9, 19, 20) {real, imag} */,
  {32'h40a8824a, 32'hc10e66a0} /* (9, 19, 19) {real, imag} */,
  {32'h40edddf4, 32'hc0883959} /* (9, 19, 18) {real, imag} */,
  {32'hc0f89216, 32'hc0d94786} /* (9, 19, 17) {real, imag} */,
  {32'h3f0784c0, 32'hbf8eca60} /* (9, 19, 16) {real, imag} */,
  {32'h4096895e, 32'h414b9a81} /* (9, 19, 15) {real, imag} */,
  {32'h406f6750, 32'h40d89a3d} /* (9, 19, 14) {real, imag} */,
  {32'h411c0f39, 32'h3f0ac9c8} /* (9, 19, 13) {real, imag} */,
  {32'hc05df290, 32'h40502a26} /* (9, 19, 12) {real, imag} */,
  {32'hc08fb16b, 32'hc18bd494} /* (9, 19, 11) {real, imag} */,
  {32'hc1becc92, 32'h3ff3db20} /* (9, 19, 10) {real, imag} */,
  {32'h40d13ee8, 32'hc088dbeb} /* (9, 19, 9) {real, imag} */,
  {32'hbfdaf060, 32'hc0c3ea02} /* (9, 19, 8) {real, imag} */,
  {32'hc06959c4, 32'h3f9ddb78} /* (9, 19, 7) {real, imag} */,
  {32'hc1adc0ad, 32'hc03eb268} /* (9, 19, 6) {real, imag} */,
  {32'hc0b7b98e, 32'h41963e6b} /* (9, 19, 5) {real, imag} */,
  {32'hc184c944, 32'hc238d4ff} /* (9, 19, 4) {real, imag} */,
  {32'h4155637d, 32'h41d3f00a} /* (9, 19, 3) {real, imag} */,
  {32'hc06e7828, 32'hc14e9b3c} /* (9, 19, 2) {real, imag} */,
  {32'h4105f17d, 32'hc1e106df} /* (9, 19, 1) {real, imag} */,
  {32'hc2084ef5, 32'hc2822d30} /* (9, 19, 0) {real, imag} */,
  {32'h40d97d86, 32'h41b50e72} /* (9, 18, 31) {real, imag} */,
  {32'h416f759e, 32'hc1f65c51} /* (9, 18, 30) {real, imag} */,
  {32'hc054e1d4, 32'h413dcbe6} /* (9, 18, 29) {real, imag} */,
  {32'hc140cece, 32'hc1867d4e} /* (9, 18, 28) {real, imag} */,
  {32'hc1acdd3e, 32'hc00ee108} /* (9, 18, 27) {real, imag} */,
  {32'h40a67c2b, 32'hc135aa98} /* (9, 18, 26) {real, imag} */,
  {32'h40dbf165, 32'h40f2fdba} /* (9, 18, 25) {real, imag} */,
  {32'hbfad53c0, 32'h406ed1c8} /* (9, 18, 24) {real, imag} */,
  {32'h404c1c62, 32'hbf86bc28} /* (9, 18, 23) {real, imag} */,
  {32'h418412c1, 32'h40955cea} /* (9, 18, 22) {real, imag} */,
  {32'h3e23b588, 32'hc1461d16} /* (9, 18, 21) {real, imag} */,
  {32'h412e828c, 32'h41a2bd85} /* (9, 18, 20) {real, imag} */,
  {32'hc037c673, 32'hc0672014} /* (9, 18, 19) {real, imag} */,
  {32'h4093a4df, 32'hbf7072b0} /* (9, 18, 18) {real, imag} */,
  {32'hc0bd8704, 32'h40572258} /* (9, 18, 17) {real, imag} */,
  {32'hc0051ca9, 32'hc04778e0} /* (9, 18, 16) {real, imag} */,
  {32'h40391b21, 32'hc0a2608c} /* (9, 18, 15) {real, imag} */,
  {32'h406386fa, 32'h4079861c} /* (9, 18, 14) {real, imag} */,
  {32'h409241d2, 32'hc0cda78a} /* (9, 18, 13) {real, imag} */,
  {32'h40f62384, 32'h3f88a230} /* (9, 18, 12) {real, imag} */,
  {32'hbf1b933e, 32'hc111ba7a} /* (9, 18, 11) {real, imag} */,
  {32'h4125b960, 32'hc0f8115a} /* (9, 18, 10) {real, imag} */,
  {32'hc08e08eb, 32'hc146daeb} /* (9, 18, 9) {real, imag} */,
  {32'hc1bbc7a2, 32'hc1938e71} /* (9, 18, 8) {real, imag} */,
  {32'hc1a46f40, 32'h3f8c3fb8} /* (9, 18, 7) {real, imag} */,
  {32'h417e2020, 32'h40d5ed6c} /* (9, 18, 6) {real, imag} */,
  {32'h4166fcc4, 32'h420bd2c0} /* (9, 18, 5) {real, imag} */,
  {32'hc16c2df8, 32'h416efa04} /* (9, 18, 4) {real, imag} */,
  {32'h419b47aa, 32'h4186fc7a} /* (9, 18, 3) {real, imag} */,
  {32'hc16facf2, 32'hc1b96ce5} /* (9, 18, 2) {real, imag} */,
  {32'hc0e5847e, 32'h414135e5} /* (9, 18, 1) {real, imag} */,
  {32'h4085f174, 32'hc116ce56} /* (9, 18, 0) {real, imag} */,
  {32'hc16971e6, 32'h41852323} /* (9, 17, 31) {real, imag} */,
  {32'h40315e4c, 32'hc1e7c3f8} /* (9, 17, 30) {real, imag} */,
  {32'h4182af92, 32'h411144de} /* (9, 17, 29) {real, imag} */,
  {32'hc1a97892, 32'hbfdcfebc} /* (9, 17, 28) {real, imag} */,
  {32'h40ac099b, 32'h41dd6b46} /* (9, 17, 27) {real, imag} */,
  {32'hc19c3f5f, 32'hc19c0084} /* (9, 17, 26) {real, imag} */,
  {32'h3f7039a4, 32'h4116da39} /* (9, 17, 25) {real, imag} */,
  {32'h4211e112, 32'h4171b084} /* (9, 17, 24) {real, imag} */,
  {32'h41861579, 32'h40e21e08} /* (9, 17, 23) {real, imag} */,
  {32'h4080174c, 32'h402cde7c} /* (9, 17, 22) {real, imag} */,
  {32'hc0ac629e, 32'h3ece2e80} /* (9, 17, 21) {real, imag} */,
  {32'h408f59b3, 32'h409a44f1} /* (9, 17, 20) {real, imag} */,
  {32'h40a0bda8, 32'h4068411e} /* (9, 17, 19) {real, imag} */,
  {32'h3f8157ad, 32'h4063dbb8} /* (9, 17, 18) {real, imag} */,
  {32'hc0892510, 32'hc0cfd3d6} /* (9, 17, 17) {real, imag} */,
  {32'hc0d46b38, 32'h3eae3920} /* (9, 17, 16) {real, imag} */,
  {32'hc0452817, 32'h3fed8bb8} /* (9, 17, 15) {real, imag} */,
  {32'hbfae87e7, 32'hc01d7690} /* (9, 17, 14) {real, imag} */,
  {32'hbf3d9bb4, 32'hc0e95507} /* (9, 17, 13) {real, imag} */,
  {32'h407c87d6, 32'h4117c780} /* (9, 17, 12) {real, imag} */,
  {32'hc0cea368, 32'hc1960dd8} /* (9, 17, 11) {real, imag} */,
  {32'h402b5f69, 32'h4124cdd1} /* (9, 17, 10) {real, imag} */,
  {32'h4197bb61, 32'h40625e99} /* (9, 17, 9) {real, imag} */,
  {32'hc0074008, 32'h4110421a} /* (9, 17, 8) {real, imag} */,
  {32'hc0a78f04, 32'h4119847d} /* (9, 17, 7) {real, imag} */,
  {32'hc13d28be, 32'hc1cdf444} /* (9, 17, 6) {real, imag} */,
  {32'hc095ebcd, 32'hbfc53100} /* (9, 17, 5) {real, imag} */,
  {32'h419836a8, 32'hc17472fc} /* (9, 17, 4) {real, imag} */,
  {32'hc05b7b12, 32'h4140a84c} /* (9, 17, 3) {real, imag} */,
  {32'hbd5af2a0, 32'hc1cb6e68} /* (9, 17, 2) {real, imag} */,
  {32'h41839134, 32'hc1229df0} /* (9, 17, 1) {real, imag} */,
  {32'h41dfac58, 32'hc026c54c} /* (9, 17, 0) {real, imag} */,
  {32'hc0f542bb, 32'h4126742d} /* (9, 16, 31) {real, imag} */,
  {32'h4143bd04, 32'hc076585c} /* (9, 16, 30) {real, imag} */,
  {32'h41046913, 32'hc13e2021} /* (9, 16, 29) {real, imag} */,
  {32'h4078be28, 32'h417e524e} /* (9, 16, 28) {real, imag} */,
  {32'h40556538, 32'h40a0fb20} /* (9, 16, 27) {real, imag} */,
  {32'h413e1a8e, 32'h4138b542} /* (9, 16, 26) {real, imag} */,
  {32'hc023aa18, 32'hc0e4eaf6} /* (9, 16, 25) {real, imag} */,
  {32'hc0d95689, 32'hc0cb59be} /* (9, 16, 24) {real, imag} */,
  {32'h40ffee8f, 32'h40f49720} /* (9, 16, 23) {real, imag} */,
  {32'h40279a5a, 32'h41182183} /* (9, 16, 22) {real, imag} */,
  {32'hbf79fca0, 32'hc0ff75fc} /* (9, 16, 21) {real, imag} */,
  {32'hc0e0623a, 32'h41847305} /* (9, 16, 20) {real, imag} */,
  {32'h40a07c27, 32'hbf2ba020} /* (9, 16, 19) {real, imag} */,
  {32'h3fcd9db8, 32'hbf3cf488} /* (9, 16, 18) {real, imag} */,
  {32'hc0ab4756, 32'hc0dd9e2f} /* (9, 16, 17) {real, imag} */,
  {32'hc039e0d6, 32'hc103c884} /* (9, 16, 16) {real, imag} */,
  {32'h40a6099a, 32'hc01547c2} /* (9, 16, 15) {real, imag} */,
  {32'hc0e4698a, 32'hbfa19b0e} /* (9, 16, 14) {real, imag} */,
  {32'hc124f9e8, 32'hc0929f92} /* (9, 16, 13) {real, imag} */,
  {32'hc0a7c4b8, 32'hc0ef5255} /* (9, 16, 12) {real, imag} */,
  {32'h403258e0, 32'h4140664a} /* (9, 16, 11) {real, imag} */,
  {32'h40168ed6, 32'h40841896} /* (9, 16, 10) {real, imag} */,
  {32'h3e8d6bf0, 32'hc0d52ef8} /* (9, 16, 9) {real, imag} */,
  {32'h40c2212f, 32'h417446e1} /* (9, 16, 8) {real, imag} */,
  {32'h410c2962, 32'h41682875} /* (9, 16, 7) {real, imag} */,
  {32'h3fce5ed4, 32'h41a192d8} /* (9, 16, 6) {real, imag} */,
  {32'h41bf7e16, 32'hc180f1b8} /* (9, 16, 5) {real, imag} */,
  {32'h4107c175, 32'hc1c860b3} /* (9, 16, 4) {real, imag} */,
  {32'hc1057d25, 32'h4104354b} /* (9, 16, 3) {real, imag} */,
  {32'hc0fefcd8, 32'hbffacce9} /* (9, 16, 2) {real, imag} */,
  {32'h4196cd39, 32'h41a8d8fc} /* (9, 16, 1) {real, imag} */,
  {32'h41284b8a, 32'hc1fac0d2} /* (9, 16, 0) {real, imag} */,
  {32'hc097d16c, 32'hbecbd7e0} /* (9, 15, 31) {real, imag} */,
  {32'h40649497, 32'h417217a8} /* (9, 15, 30) {real, imag} */,
  {32'h41c12d6c, 32'h41ca27d2} /* (9, 15, 29) {real, imag} */,
  {32'hc1513797, 32'hc1319bb0} /* (9, 15, 28) {real, imag} */,
  {32'h40e2181b, 32'h41ced1ec} /* (9, 15, 27) {real, imag} */,
  {32'h40b9609c, 32'h40219a3f} /* (9, 15, 26) {real, imag} */,
  {32'hc17c8e42, 32'hc11c7eb6} /* (9, 15, 25) {real, imag} */,
  {32'hc0e2ca0c, 32'hc0bad4fd} /* (9, 15, 24) {real, imag} */,
  {32'hc0cd4195, 32'hc05194fd} /* (9, 15, 23) {real, imag} */,
  {32'hc15b0018, 32'hc0cdc635} /* (9, 15, 22) {real, imag} */,
  {32'hbf9a68c0, 32'h40c56271} /* (9, 15, 21) {real, imag} */,
  {32'hbff5607e, 32'hc0f6a562} /* (9, 15, 20) {real, imag} */,
  {32'h40b0dfa7, 32'h4102a732} /* (9, 15, 19) {real, imag} */,
  {32'h3f545c0c, 32'h3fb6de70} /* (9, 15, 18) {real, imag} */,
  {32'h402718a8, 32'hbfd6b254} /* (9, 15, 17) {real, imag} */,
  {32'hc02038e6, 32'hc0401760} /* (9, 15, 16) {real, imag} */,
  {32'h411bea26, 32'h40835637} /* (9, 15, 15) {real, imag} */,
  {32'h40d89d92, 32'hc0c6ca24} /* (9, 15, 14) {real, imag} */,
  {32'h412c18b4, 32'hbfef70b2} /* (9, 15, 13) {real, imag} */,
  {32'hc0a836f4, 32'hc0d2ff22} /* (9, 15, 12) {real, imag} */,
  {32'hc12191fb, 32'h40a4736b} /* (9, 15, 11) {real, imag} */,
  {32'h411df8a0, 32'h41613a76} /* (9, 15, 10) {real, imag} */,
  {32'hc0515f86, 32'hc089b046} /* (9, 15, 9) {real, imag} */,
  {32'h41a5af42, 32'hc062ed9e} /* (9, 15, 8) {real, imag} */,
  {32'h40c1738c, 32'hc1171d8c} /* (9, 15, 7) {real, imag} */,
  {32'hc1aef25b, 32'h40ec4902} /* (9, 15, 6) {real, imag} */,
  {32'hc138493a, 32'hc0a024b6} /* (9, 15, 5) {real, imag} */,
  {32'hc1b2cc38, 32'hbfa37e8c} /* (9, 15, 4) {real, imag} */,
  {32'h406c1d00, 32'hc0f48078} /* (9, 15, 3) {real, imag} */,
  {32'hbf700fdc, 32'h41797fb8} /* (9, 15, 2) {real, imag} */,
  {32'hc1ca7449, 32'h41b32ab2} /* (9, 15, 1) {real, imag} */,
  {32'h413b6ac8, 32'hc100adc6} /* (9, 15, 0) {real, imag} */,
  {32'h4157a719, 32'h40f73310} /* (9, 14, 31) {real, imag} */,
  {32'hc1fad973, 32'hc10d8173} /* (9, 14, 30) {real, imag} */,
  {32'hc1f1ea8b, 32'h408f4a16} /* (9, 14, 29) {real, imag} */,
  {32'h418de397, 32'h4231c378} /* (9, 14, 28) {real, imag} */,
  {32'hbed76030, 32'hc1d478c7} /* (9, 14, 27) {real, imag} */,
  {32'hc155080e, 32'hc097c568} /* (9, 14, 26) {real, imag} */,
  {32'hc1b5fb48, 32'hc13fbf87} /* (9, 14, 25) {real, imag} */,
  {32'hc0e9ec70, 32'hbf6855a8} /* (9, 14, 24) {real, imag} */,
  {32'h3f07f510, 32'hc14ded48} /* (9, 14, 23) {real, imag} */,
  {32'h3fd85b36, 32'hc12babc4} /* (9, 14, 22) {real, imag} */,
  {32'hc0d8314a, 32'hc105c6f4} /* (9, 14, 21) {real, imag} */,
  {32'hc07f9036, 32'h40d65070} /* (9, 14, 20) {real, imag} */,
  {32'hc0caec28, 32'hc107d9c8} /* (9, 14, 19) {real, imag} */,
  {32'hbce7ea00, 32'h3fb17d56} /* (9, 14, 18) {real, imag} */,
  {32'h3fd56ed6, 32'hc0ca9dc3} /* (9, 14, 17) {real, imag} */,
  {32'hc0120ada, 32'h3ff708a8} /* (9, 14, 16) {real, imag} */,
  {32'hc0015a35, 32'hbe847bb0} /* (9, 14, 15) {real, imag} */,
  {32'hc01adc54, 32'hc04284f9} /* (9, 14, 14) {real, imag} */,
  {32'h3d90ea00, 32'h3fe1d02c} /* (9, 14, 13) {real, imag} */,
  {32'hc069ff0a, 32'hbea3f178} /* (9, 14, 12) {real, imag} */,
  {32'h40c3d99e, 32'h40eefca9} /* (9, 14, 11) {real, imag} */,
  {32'hc0480049, 32'h418d597a} /* (9, 14, 10) {real, imag} */,
  {32'hc13218f1, 32'h41083e06} /* (9, 14, 9) {real, imag} */,
  {32'h415bfce8, 32'hc1784d14} /* (9, 14, 8) {real, imag} */,
  {32'hc22cf9c2, 32'hc1374ae5} /* (9, 14, 7) {real, imag} */,
  {32'h3f8e5924, 32'h3ff0deff} /* (9, 14, 6) {real, imag} */,
  {32'h4154b3ba, 32'h40633ba8} /* (9, 14, 5) {real, imag} */,
  {32'h420c410c, 32'h4224f5c0} /* (9, 14, 4) {real, imag} */,
  {32'h40f74a3c, 32'h41b8d046} /* (9, 14, 3) {real, imag} */,
  {32'hc1a227ed, 32'h3faf4696} /* (9, 14, 2) {real, imag} */,
  {32'hc16736bf, 32'h41d2f166} /* (9, 14, 1) {real, imag} */,
  {32'hc0d10f5f, 32'h41ed053a} /* (9, 14, 0) {real, imag} */,
  {32'hc0cd3e7c, 32'hc1b788c2} /* (9, 13, 31) {real, imag} */,
  {32'h42003218, 32'hc094b316} /* (9, 13, 30) {real, imag} */,
  {32'h4001da8c, 32'h41acc3d4} /* (9, 13, 29) {real, imag} */,
  {32'h40f6f468, 32'hc2273f18} /* (9, 13, 28) {real, imag} */,
  {32'h40bb7404, 32'hc1191e78} /* (9, 13, 27) {real, imag} */,
  {32'hc193dce3, 32'hc127322f} /* (9, 13, 26) {real, imag} */,
  {32'h409cd22b, 32'h40d0ef9f} /* (9, 13, 25) {real, imag} */,
  {32'h41162a8c, 32'hc1d3a725} /* (9, 13, 24) {real, imag} */,
  {32'h40667184, 32'hc10dce4a} /* (9, 13, 23) {real, imag} */,
  {32'h4104aa32, 32'hc123bdc6} /* (9, 13, 22) {real, imag} */,
  {32'h3fc3eb38, 32'h406d6e97} /* (9, 13, 21) {real, imag} */,
  {32'hbf803a58, 32'hc14cb6a3} /* (9, 13, 20) {real, imag} */,
  {32'h40292645, 32'h417010e6} /* (9, 13, 19) {real, imag} */,
  {32'h3fd22d44, 32'hbf14e368} /* (9, 13, 18) {real, imag} */,
  {32'h40a3ccfa, 32'h40ac277e} /* (9, 13, 17) {real, imag} */,
  {32'hbf3ecf08, 32'h3ee26c10} /* (9, 13, 16) {real, imag} */,
  {32'hc06e1d4c, 32'hbfeecd56} /* (9, 13, 15) {real, imag} */,
  {32'h3f196908, 32'h40229c3e} /* (9, 13, 14) {real, imag} */,
  {32'h409d8b7a, 32'h4103a3ac} /* (9, 13, 13) {real, imag} */,
  {32'hbfeb0b78, 32'h417ab6a7} /* (9, 13, 12) {real, imag} */,
  {32'h41af6572, 32'hc11cd4f6} /* (9, 13, 11) {real, imag} */,
  {32'hc186a16b, 32'h4130c49a} /* (9, 13, 10) {real, imag} */,
  {32'hc1a9cac2, 32'h4178e696} /* (9, 13, 9) {real, imag} */,
  {32'hc16db2e4, 32'hc1108002} /* (9, 13, 8) {real, imag} */,
  {32'hbeafd790, 32'hbeb76070} /* (9, 13, 7) {real, imag} */,
  {32'h3f282e20, 32'h414bcbf1} /* (9, 13, 6) {real, imag} */,
  {32'hc22202dc, 32'h4190045c} /* (9, 13, 5) {real, imag} */,
  {32'h4230728b, 32'h41318b38} /* (9, 13, 4) {real, imag} */,
  {32'hc1198c5d, 32'hc20db04c} /* (9, 13, 3) {real, imag} */,
  {32'hc1456c06, 32'hc1bae1ec} /* (9, 13, 2) {real, imag} */,
  {32'hc2171710, 32'hc13a8fc8} /* (9, 13, 1) {real, imag} */,
  {32'hc02af172, 32'hc0eb78b1} /* (9, 13, 0) {real, imag} */,
  {32'h41ec5bdb, 32'h4227c8df} /* (9, 12, 31) {real, imag} */,
  {32'hc12a55e6, 32'h40ce15aa} /* (9, 12, 30) {real, imag} */,
  {32'hc2150edb, 32'h40a8368d} /* (9, 12, 29) {real, imag} */,
  {32'hc0539cf2, 32'h41cae3ea} /* (9, 12, 28) {real, imag} */,
  {32'hc13949e7, 32'hc1ee2075} /* (9, 12, 27) {real, imag} */,
  {32'hc2169408, 32'h42058bed} /* (9, 12, 26) {real, imag} */,
  {32'hc0eb5d0a, 32'hc1ac0d8f} /* (9, 12, 25) {real, imag} */,
  {32'h418056c3, 32'h4155b167} /* (9, 12, 24) {real, imag} */,
  {32'hc1258b4f, 32'h41db2949} /* (9, 12, 23) {real, imag} */,
  {32'hc12f7c48, 32'hc11a87f3} /* (9, 12, 22) {real, imag} */,
  {32'h41342bf8, 32'h41d73cec} /* (9, 12, 21) {real, imag} */,
  {32'h3ffa95e4, 32'h3efe04e0} /* (9, 12, 20) {real, imag} */,
  {32'h412d3dbb, 32'hc01b01d1} /* (9, 12, 19) {real, imag} */,
  {32'h41834268, 32'h4006e8d8} /* (9, 12, 18) {real, imag} */,
  {32'h4131fa0c, 32'h4045dfec} /* (9, 12, 17) {real, imag} */,
  {32'hc1312856, 32'hc07b9384} /* (9, 12, 16) {real, imag} */,
  {32'hbfbbefc0, 32'hc080bb8a} /* (9, 12, 15) {real, imag} */,
  {32'h401a26ac, 32'hc08c9aa4} /* (9, 12, 14) {real, imag} */,
  {32'h4113fa11, 32'h410c585c} /* (9, 12, 13) {real, imag} */,
  {32'h40e0c1d1, 32'hbf534880} /* (9, 12, 12) {real, imag} */,
  {32'h4131ba96, 32'hc0b458b2} /* (9, 12, 11) {real, imag} */,
  {32'hc0e273d0, 32'h415fea1b} /* (9, 12, 10) {real, imag} */,
  {32'h3db02680, 32'hc1aa969b} /* (9, 12, 9) {real, imag} */,
  {32'hbf0d69d8, 32'h41a60217} /* (9, 12, 8) {real, imag} */,
  {32'h419aa42c, 32'h407f28e8} /* (9, 12, 7) {real, imag} */,
  {32'h41106ce2, 32'h412d5f7b} /* (9, 12, 6) {real, imag} */,
  {32'h41846d40, 32'hc1c75f4f} /* (9, 12, 5) {real, imag} */,
  {32'h41083dee, 32'h40a3f550} /* (9, 12, 4) {real, imag} */,
  {32'hc1b14f5c, 32'h3f22e2f0} /* (9, 12, 3) {real, imag} */,
  {32'h420dbaee, 32'h40fe3526} /* (9, 12, 2) {real, imag} */,
  {32'h4217adde, 32'hc1bc2772} /* (9, 12, 1) {real, imag} */,
  {32'hc1cadcf1, 32'h410ba776} /* (9, 12, 0) {real, imag} */,
  {32'hc1440618, 32'hc15f7c22} /* (9, 11, 31) {real, imag} */,
  {32'hc0a2a3f6, 32'hc216bb10} /* (9, 11, 30) {real, imag} */,
  {32'hc22d6160, 32'hc16f4728} /* (9, 11, 29) {real, imag} */,
  {32'hc1c13bec, 32'hc0e7f0cd} /* (9, 11, 28) {real, imag} */,
  {32'hc2700c7e, 32'h419a344a} /* (9, 11, 27) {real, imag} */,
  {32'h418f9cb6, 32'h41f41f31} /* (9, 11, 26) {real, imag} */,
  {32'h424bc205, 32'h41e4afcd} /* (9, 11, 25) {real, imag} */,
  {32'h4216f8f4, 32'hc028e3e8} /* (9, 11, 24) {real, imag} */,
  {32'hc21b912e, 32'hc091254a} /* (9, 11, 23) {real, imag} */,
  {32'hbf2d2ae0, 32'h4176a6d2} /* (9, 11, 22) {real, imag} */,
  {32'hc1abfbb3, 32'hc1aedbe0} /* (9, 11, 21) {real, imag} */,
  {32'h40e2302e, 32'hc158cbe3} /* (9, 11, 20) {real, imag} */,
  {32'h412f2fb2, 32'hc0bde3be} /* (9, 11, 19) {real, imag} */,
  {32'hbf9ce3d8, 32'h411b6aae} /* (9, 11, 18) {real, imag} */,
  {32'h40d26758, 32'hc1554398} /* (9, 11, 17) {real, imag} */,
  {32'hbfd36880, 32'hc0bef81a} /* (9, 11, 16) {real, imag} */,
  {32'hc110f31a, 32'h40f0df89} /* (9, 11, 15) {real, imag} */,
  {32'h4115d313, 32'h405b5018} /* (9, 11, 14) {real, imag} */,
  {32'h3f9f4710, 32'h4124f199} /* (9, 11, 13) {real, imag} */,
  {32'h41124ca1, 32'h40fd9212} /* (9, 11, 12) {real, imag} */,
  {32'hc19cb933, 32'hbfc8cd08} /* (9, 11, 11) {real, imag} */,
  {32'h416987d8, 32'h4205d35e} /* (9, 11, 10) {real, imag} */,
  {32'h4203871e, 32'hbfb10f86} /* (9, 11, 9) {real, imag} */,
  {32'h41b67d04, 32'h41907434} /* (9, 11, 8) {real, imag} */,
  {32'h41e7625e, 32'h41a7476b} /* (9, 11, 7) {real, imag} */,
  {32'h41551cee, 32'h41f5976b} /* (9, 11, 6) {real, imag} */,
  {32'h4233f14a, 32'h4253038f} /* (9, 11, 5) {real, imag} */,
  {32'h41cb3b3c, 32'hc1a24d3a} /* (9, 11, 4) {real, imag} */,
  {32'hc1fb5d21, 32'h4285d6b2} /* (9, 11, 3) {real, imag} */,
  {32'hc07f8f63, 32'h41d69f64} /* (9, 11, 2) {real, imag} */,
  {32'h42313422, 32'h412e9ae6} /* (9, 11, 1) {real, imag} */,
  {32'hc23c5390, 32'h419743ca} /* (9, 11, 0) {real, imag} */,
  {32'h419823eb, 32'hc1c43a5a} /* (9, 10, 31) {real, imag} */,
  {32'hc24912a2, 32'hc1467b59} /* (9, 10, 30) {real, imag} */,
  {32'h40eeadf4, 32'hc19f3464} /* (9, 10, 29) {real, imag} */,
  {32'h404ab040, 32'h41229845} /* (9, 10, 28) {real, imag} */,
  {32'h4257bb85, 32'hc1d2625b} /* (9, 10, 27) {real, imag} */,
  {32'h419ea63f, 32'h42170218} /* (9, 10, 26) {real, imag} */,
  {32'h41edeaec, 32'h3c85fc00} /* (9, 10, 25) {real, imag} */,
  {32'hc12abe5b, 32'h41e8165b} /* (9, 10, 24) {real, imag} */,
  {32'h41e99050, 32'h41c53006} /* (9, 10, 23) {real, imag} */,
  {32'hc106da6a, 32'h4177ba16} /* (9, 10, 22) {real, imag} */,
  {32'h41a96541, 32'h403af756} /* (9, 10, 21) {real, imag} */,
  {32'hbfebca48, 32'hc201c921} /* (9, 10, 20) {real, imag} */,
  {32'hc1e0fb87, 32'hc15fa060} /* (9, 10, 19) {real, imag} */,
  {32'h40ee38ac, 32'hc18aee5a} /* (9, 10, 18) {real, imag} */,
  {32'h4114b340, 32'hc06f9bcc} /* (9, 10, 17) {real, imag} */,
  {32'h411864e1, 32'h417f419b} /* (9, 10, 16) {real, imag} */,
  {32'hc143d658, 32'hc14920b1} /* (9, 10, 15) {real, imag} */,
  {32'hbffca890, 32'hc1896992} /* (9, 10, 14) {real, imag} */,
  {32'hc036bd78, 32'hc118bb8c} /* (9, 10, 13) {real, imag} */,
  {32'h412af84d, 32'hc12b2208} /* (9, 10, 12) {real, imag} */,
  {32'h41b2dc4b, 32'h3f0ab918} /* (9, 10, 11) {real, imag} */,
  {32'hc0868c7d, 32'hc19694b1} /* (9, 10, 10) {real, imag} */,
  {32'h41220ea7, 32'h41321c1c} /* (9, 10, 9) {real, imag} */,
  {32'h411cdf3b, 32'hc18583c9} /* (9, 10, 8) {real, imag} */,
  {32'hc1d80aac, 32'hc134b619} /* (9, 10, 7) {real, imag} */,
  {32'hc0640058, 32'hc15117ba} /* (9, 10, 6) {real, imag} */,
  {32'h4145da5c, 32'h41b486d3} /* (9, 10, 5) {real, imag} */,
  {32'h3eeff074, 32'h419f51e4} /* (9, 10, 4) {real, imag} */,
  {32'hc242e442, 32'h4253824a} /* (9, 10, 3) {real, imag} */,
  {32'h42bb4483, 32'h40cc5106} /* (9, 10, 2) {real, imag} */,
  {32'hc11bc20e, 32'hbed0a120} /* (9, 10, 1) {real, imag} */,
  {32'hc1d5f358, 32'h4197d244} /* (9, 10, 0) {real, imag} */,
  {32'hc2595442, 32'h42100e2c} /* (9, 9, 31) {real, imag} */,
  {32'h424a2fb6, 32'hc21b5868} /* (9, 9, 30) {real, imag} */,
  {32'h4163ddae, 32'h412bd21a} /* (9, 9, 29) {real, imag} */,
  {32'h41fbca09, 32'h41e66966} /* (9, 9, 28) {real, imag} */,
  {32'hc17b0404, 32'hc106e38e} /* (9, 9, 27) {real, imag} */,
  {32'hc247a287, 32'hc21b5410} /* (9, 9, 26) {real, imag} */,
  {32'hc22b0036, 32'h42024028} /* (9, 9, 25) {real, imag} */,
  {32'h3fc3f610, 32'h4051793c} /* (9, 9, 24) {real, imag} */,
  {32'hbfd9d0a0, 32'h402ac1e0} /* (9, 9, 23) {real, imag} */,
  {32'h3fc01548, 32'hc23a6dff} /* (9, 9, 22) {real, imag} */,
  {32'h419ba6c3, 32'hc0cd347e} /* (9, 9, 21) {real, imag} */,
  {32'h4173ddd4, 32'h416b2694} /* (9, 9, 20) {real, imag} */,
  {32'h41a32468, 32'hc1a9c406} /* (9, 9, 19) {real, imag} */,
  {32'h3d322280, 32'h3fc0d980} /* (9, 9, 18) {real, imag} */,
  {32'hc0a2cd72, 32'hc1353414} /* (9, 9, 17) {real, imag} */,
  {32'h3f849d48, 32'hc16688fe} /* (9, 9, 16) {real, imag} */,
  {32'hc05a929c, 32'hc087934d} /* (9, 9, 15) {real, imag} */,
  {32'hc0ea2b85, 32'h41517c68} /* (9, 9, 14) {real, imag} */,
  {32'hc04d18d0, 32'h40181974} /* (9, 9, 13) {real, imag} */,
  {32'hc1aad1ec, 32'hc1f9dcee} /* (9, 9, 12) {real, imag} */,
  {32'hc1a92acf, 32'h41823ad4} /* (9, 9, 11) {real, imag} */,
  {32'h41a9ac44, 32'h42218165} /* (9, 9, 10) {real, imag} */,
  {32'hc1ca8a3c, 32'hc1b1570c} /* (9, 9, 9) {real, imag} */,
  {32'hc206d01e, 32'hc1934fe6} /* (9, 9, 8) {real, imag} */,
  {32'hc2573c8a, 32'hc1beff37} /* (9, 9, 7) {real, imag} */,
  {32'h414a57e4, 32'hc2187072} /* (9, 9, 6) {real, imag} */,
  {32'h421e8482, 32'h400edee0} /* (9, 9, 5) {real, imag} */,
  {32'h41785bb2, 32'hc249d2ab} /* (9, 9, 4) {real, imag} */,
  {32'h41f2be43, 32'h3faca280} /* (9, 9, 3) {real, imag} */,
  {32'h4217bdd0, 32'h41e91f33} /* (9, 9, 2) {real, imag} */,
  {32'hc20871b2, 32'hc1f8b241} /* (9, 9, 1) {real, imag} */,
  {32'hc1f6beaa, 32'h429ae8a4} /* (9, 9, 0) {real, imag} */,
  {32'hc2b716bc, 32'hc20770be} /* (9, 8, 31) {real, imag} */,
  {32'hc232c74a, 32'h4210011a} /* (9, 8, 30) {real, imag} */,
  {32'h417eb1e9, 32'h420ca02a} /* (9, 8, 29) {real, imag} */,
  {32'hc151e0f4, 32'hc23226d0} /* (9, 8, 28) {real, imag} */,
  {32'h40e6ea08, 32'hc15ff55e} /* (9, 8, 27) {real, imag} */,
  {32'h42d15e8a, 32'hc14b82e5} /* (9, 8, 26) {real, imag} */,
  {32'hc0b52374, 32'hc07becf8} /* (9, 8, 25) {real, imag} */,
  {32'hc18e88ac, 32'hc200f046} /* (9, 8, 24) {real, imag} */,
  {32'h3f345160, 32'h3f473ca0} /* (9, 8, 23) {real, imag} */,
  {32'h4146654b, 32'hc15e97b0} /* (9, 8, 22) {real, imag} */,
  {32'hc1ec8d94, 32'h417b3689} /* (9, 8, 21) {real, imag} */,
  {32'hc05498ec, 32'h40a14c34} /* (9, 8, 20) {real, imag} */,
  {32'hbf3e9da0, 32'h41e730b6} /* (9, 8, 19) {real, imag} */,
  {32'h40170504, 32'hc0cf53f8} /* (9, 8, 18) {real, imag} */,
  {32'hc1baa2da, 32'h401cf920} /* (9, 8, 17) {real, imag} */,
  {32'hc1045230, 32'hc1635639} /* (9, 8, 16) {real, imag} */,
  {32'hc1010c33, 32'hc1886980} /* (9, 8, 15) {real, imag} */,
  {32'h419c6dba, 32'h400a1918} /* (9, 8, 14) {real, imag} */,
  {32'hc181f876, 32'h3f91b2d8} /* (9, 8, 13) {real, imag} */,
  {32'hc14bb575, 32'h41a56bc1} /* (9, 8, 12) {real, imag} */,
  {32'h418d47ec, 32'h4133dd83} /* (9, 8, 11) {real, imag} */,
  {32'h40a55b76, 32'hc23bf026} /* (9, 8, 10) {real, imag} */,
  {32'hc0b4e4b8, 32'hc2741840} /* (9, 8, 9) {real, imag} */,
  {32'hc14b69f8, 32'h41b68da2} /* (9, 8, 8) {real, imag} */,
  {32'hc17a6b7c, 32'hc1aa3bd1} /* (9, 8, 7) {real, imag} */,
  {32'hc209d310, 32'h41102125} /* (9, 8, 6) {real, imag} */,
  {32'hc2c1353c, 32'h41f456e9} /* (9, 8, 5) {real, imag} */,
  {32'h41e2600e, 32'h42a95e2c} /* (9, 8, 4) {real, imag} */,
  {32'h41948684, 32'hc21ed154} /* (9, 8, 3) {real, imag} */,
  {32'h404ae808, 32'h40e88c42} /* (9, 8, 2) {real, imag} */,
  {32'h429de164, 32'hc1dd124c} /* (9, 8, 1) {real, imag} */,
  {32'h431ddfba, 32'hc160e175} /* (9, 8, 0) {real, imag} */,
  {32'hc193ed36, 32'h40d36f80} /* (9, 7, 31) {real, imag} */,
  {32'h424d8556, 32'h429d87ce} /* (9, 7, 30) {real, imag} */,
  {32'hc24ee99a, 32'hc20bbb94} /* (9, 7, 29) {real, imag} */,
  {32'h42e4a13f, 32'h41280b90} /* (9, 7, 28) {real, imag} */,
  {32'h417cc512, 32'hc26aae95} /* (9, 7, 27) {real, imag} */,
  {32'hc113b547, 32'hc2a44265} /* (9, 7, 26) {real, imag} */,
  {32'hc188038f, 32'hc0f3b4c9} /* (9, 7, 25) {real, imag} */,
  {32'hc2f0cfab, 32'h3ea09b00} /* (9, 7, 24) {real, imag} */,
  {32'h41fdbae0, 32'hc1301b7c} /* (9, 7, 23) {real, imag} */,
  {32'hc1722e64, 32'h4020530c} /* (9, 7, 22) {real, imag} */,
  {32'hc081278e, 32'hc13c1f8f} /* (9, 7, 21) {real, imag} */,
  {32'h41e76c28, 32'hc23b5ba2} /* (9, 7, 20) {real, imag} */,
  {32'hc17c7e19, 32'h41bb564a} /* (9, 7, 19) {real, imag} */,
  {32'h417c17b0, 32'hc177bc63} /* (9, 7, 18) {real, imag} */,
  {32'hc14dd36f, 32'h40c2fb90} /* (9, 7, 17) {real, imag} */,
  {32'hc17587a4, 32'h409736d4} /* (9, 7, 16) {real, imag} */,
  {32'hc17ed4d7, 32'h40aa5560} /* (9, 7, 15) {real, imag} */,
  {32'h410b9dc8, 32'h410c83ed} /* (9, 7, 14) {real, imag} */,
  {32'hc0c33b96, 32'h424b2a7f} /* (9, 7, 13) {real, imag} */,
  {32'hc1be0d3a, 32'h41eeb5fd} /* (9, 7, 12) {real, imag} */,
  {32'h4170e8b9, 32'h4106131b} /* (9, 7, 11) {real, imag} */,
  {32'hc1cd4f82, 32'hc1a03e9c} /* (9, 7, 10) {real, imag} */,
  {32'hc1ffa4e2, 32'h417d2ad4} /* (9, 7, 9) {real, imag} */,
  {32'hc1faeddc, 32'hc2a66952} /* (9, 7, 8) {real, imag} */,
  {32'hc2098c96, 32'h41979488} /* (9, 7, 7) {real, imag} */,
  {32'h418a022a, 32'h41687698} /* (9, 7, 6) {real, imag} */,
  {32'h40ac87b7, 32'hc1f50fe6} /* (9, 7, 5) {real, imag} */,
  {32'hc27e99ba, 32'h40fd8550} /* (9, 7, 4) {real, imag} */,
  {32'hc1d0761c, 32'h4264a232} /* (9, 7, 3) {real, imag} */,
  {32'hc2a4e0a9, 32'hc1975822} /* (9, 7, 2) {real, imag} */,
  {32'hc1b04b9a, 32'hc2d833c3} /* (9, 7, 1) {real, imag} */,
  {32'hc27e05fb, 32'h425bce54} /* (9, 7, 0) {real, imag} */,
  {32'h429a72ed, 32'hc1afb3ab} /* (9, 6, 31) {real, imag} */,
  {32'h428e0ca5, 32'h4256e73c} /* (9, 6, 30) {real, imag} */,
  {32'h40fa7a71, 32'h41300344} /* (9, 6, 29) {real, imag} */,
  {32'hc211b607, 32'hc20b5df0} /* (9, 6, 28) {real, imag} */,
  {32'h41188700, 32'hc18ee2f1} /* (9, 6, 27) {real, imag} */,
  {32'h422021e2, 32'h42e0b106} /* (9, 6, 26) {real, imag} */,
  {32'h4160ac1c, 32'hc114debc} /* (9, 6, 25) {real, imag} */,
  {32'h41b2a974, 32'h41709e50} /* (9, 6, 24) {real, imag} */,
  {32'h4281b360, 32'h4193e66a} /* (9, 6, 23) {real, imag} */,
  {32'h40ba1b82, 32'hbf7413e0} /* (9, 6, 22) {real, imag} */,
  {32'h40b14d3e, 32'hc0e0d034} /* (9, 6, 21) {real, imag} */,
  {32'hc19fa803, 32'h4210df88} /* (9, 6, 20) {real, imag} */,
  {32'h407f0252, 32'h40da27bd} /* (9, 6, 19) {real, imag} */,
  {32'hc1ac4b8f, 32'h41ab630c} /* (9, 6, 18) {real, imag} */,
  {32'hbf529608, 32'hc08ef32c} /* (9, 6, 17) {real, imag} */,
  {32'h4194424a, 32'hc11258a6} /* (9, 6, 16) {real, imag} */,
  {32'h40c99e11, 32'h4126cce2} /* (9, 6, 15) {real, imag} */,
  {32'hc17bae0a, 32'h41b66208} /* (9, 6, 14) {real, imag} */,
  {32'h4191722b, 32'hc13d35de} /* (9, 6, 13) {real, imag} */,
  {32'h4240a044, 32'h403615e8} /* (9, 6, 12) {real, imag} */,
  {32'hc11f9217, 32'hc24c80e6} /* (9, 6, 11) {real, imag} */,
  {32'h41b1528e, 32'hc111401e} /* (9, 6, 10) {real, imag} */,
  {32'h41450c60, 32'h40f27dff} /* (9, 6, 9) {real, imag} */,
  {32'h4219ff30, 32'hc1a777e0} /* (9, 6, 8) {real, imag} */,
  {32'h420bd38f, 32'hc1e85520} /* (9, 6, 7) {real, imag} */,
  {32'hc201664c, 32'hc262c454} /* (9, 6, 6) {real, imag} */,
  {32'hc2717628, 32'h4162771e} /* (9, 6, 5) {real, imag} */,
  {32'hc271d11d, 32'hc2914f9b} /* (9, 6, 4) {real, imag} */,
  {32'h4191052b, 32'h4109f474} /* (9, 6, 3) {real, imag} */,
  {32'h41f89cf7, 32'h43023edf} /* (9, 6, 2) {real, imag} */,
  {32'h4299f3f3, 32'hc1bcd3fb} /* (9, 6, 1) {real, imag} */,
  {32'hc2cab314, 32'h412172e2} /* (9, 6, 0) {real, imag} */,
  {32'hc0caabe4, 32'hc25da380} /* (9, 5, 31) {real, imag} */,
  {32'hc2ab153c, 32'h4257cf75} /* (9, 5, 30) {real, imag} */,
  {32'hc2729a6a, 32'hc2ac6598} /* (9, 5, 29) {real, imag} */,
  {32'h42417085, 32'hc215df06} /* (9, 5, 28) {real, imag} */,
  {32'h412266ec, 32'h425104d8} /* (9, 5, 27) {real, imag} */,
  {32'h420d033c, 32'hc0a68243} /* (9, 5, 26) {real, imag} */,
  {32'h404a13c8, 32'h4231d87f} /* (9, 5, 25) {real, imag} */,
  {32'hc2023793, 32'hc2cba612} /* (9, 5, 24) {real, imag} */,
  {32'hc1e18506, 32'hc258506e} /* (9, 5, 23) {real, imag} */,
  {32'h41ef8e53, 32'hc00e5bc6} /* (9, 5, 22) {real, imag} */,
  {32'hc1c9e2fe, 32'h412959d4} /* (9, 5, 21) {real, imag} */,
  {32'hbebce460, 32'h41bb6d71} /* (9, 5, 20) {real, imag} */,
  {32'h4272e794, 32'hc1e34290} /* (9, 5, 19) {real, imag} */,
  {32'h41bb0d8d, 32'hc04c8aa4} /* (9, 5, 18) {real, imag} */,
  {32'h40e1b5d2, 32'hc101d7fa} /* (9, 5, 17) {real, imag} */,
  {32'hc085bc28, 32'hc07beac0} /* (9, 5, 16) {real, imag} */,
  {32'h4185222a, 32'hc2198684} /* (9, 5, 15) {real, imag} */,
  {32'hc07337e8, 32'h41167b5f} /* (9, 5, 14) {real, imag} */,
  {32'h41d9f487, 32'hc167a7b0} /* (9, 5, 13) {real, imag} */,
  {32'h41b380b2, 32'h41224e6e} /* (9, 5, 12) {real, imag} */,
  {32'hc21aeb73, 32'hc2a334f4} /* (9, 5, 11) {real, imag} */,
  {32'hc08f75e4, 32'h40adce07} /* (9, 5, 10) {real, imag} */,
  {32'h424d7989, 32'hc21c80ee} /* (9, 5, 9) {real, imag} */,
  {32'h405c6a10, 32'hc196854a} /* (9, 5, 8) {real, imag} */,
  {32'h42830a6c, 32'hc089b938} /* (9, 5, 7) {real, imag} */,
  {32'hc2ae36c3, 32'hc0b8bb49} /* (9, 5, 6) {real, imag} */,
  {32'h4266d73b, 32'hc029ae98} /* (9, 5, 5) {real, imag} */,
  {32'hc21b24a3, 32'h427a6496} /* (9, 5, 4) {real, imag} */,
  {32'hc2a78a0b, 32'hc126c250} /* (9, 5, 3) {real, imag} */,
  {32'h42169584, 32'hc27fba59} /* (9, 5, 2) {real, imag} */,
  {32'h423bdf40, 32'hc19b5898} /* (9, 5, 1) {real, imag} */,
  {32'h42902cf0, 32'hc2a102b8} /* (9, 5, 0) {real, imag} */,
  {32'h42503bf2, 32'h41ed99df} /* (9, 4, 31) {real, imag} */,
  {32'h42398a27, 32'hc24d4b3e} /* (9, 4, 30) {real, imag} */,
  {32'h418a7f98, 32'h42eba3de} /* (9, 4, 29) {real, imag} */,
  {32'h4255c03e, 32'hc14895be} /* (9, 4, 28) {real, imag} */,
  {32'hc2c3b185, 32'h42f75bf0} /* (9, 4, 27) {real, imag} */,
  {32'h41a10216, 32'h42846dd7} /* (9, 4, 26) {real, imag} */,
  {32'h4306161d, 32'h41ce4a98} /* (9, 4, 25) {real, imag} */,
  {32'hc2470033, 32'h420af216} /* (9, 4, 24) {real, imag} */,
  {32'hc2129a89, 32'hc1ee60f6} /* (9, 4, 23) {real, imag} */,
  {32'hc276778a, 32'hc21dc06f} /* (9, 4, 22) {real, imag} */,
  {32'h41339f48, 32'hc1df8ebc} /* (9, 4, 21) {real, imag} */,
  {32'h410fd1fa, 32'h42044437} /* (9, 4, 20) {real, imag} */,
  {32'h3f73dac0, 32'h4203eb4a} /* (9, 4, 19) {real, imag} */,
  {32'h41726760, 32'h415e4694} /* (9, 4, 18) {real, imag} */,
  {32'hc1a176bb, 32'h410d8e30} /* (9, 4, 17) {real, imag} */,
  {32'hc0e879e0, 32'h41258d76} /* (9, 4, 16) {real, imag} */,
  {32'hc1f1089d, 32'h4163f134} /* (9, 4, 15) {real, imag} */,
  {32'h411c3204, 32'hc1454858} /* (9, 4, 14) {real, imag} */,
  {32'h4197d4b8, 32'h41a1aac0} /* (9, 4, 13) {real, imag} */,
  {32'hc0d7a2e7, 32'hc1d181a2} /* (9, 4, 12) {real, imag} */,
  {32'h42834e75, 32'hc1b86890} /* (9, 4, 11) {real, imag} */,
  {32'h41be7929, 32'hc21351d3} /* (9, 4, 10) {real, imag} */,
  {32'h42051adb, 32'h424e8b9f} /* (9, 4, 9) {real, imag} */,
  {32'hc1cdab5a, 32'hc1c3a06a} /* (9, 4, 8) {real, imag} */,
  {32'h419d9b58, 32'hc21441ea} /* (9, 4, 7) {real, imag} */,
  {32'hc2bf10cc, 32'h4275be8f} /* (9, 4, 6) {real, imag} */,
  {32'hc1d27da4, 32'hc195ebce} /* (9, 4, 5) {real, imag} */,
  {32'hc1cb5499, 32'h41e6011d} /* (9, 4, 4) {real, imag} */,
  {32'h42dee63e, 32'h40b5ecf0} /* (9, 4, 3) {real, imag} */,
  {32'hbfcdf680, 32'h41c5260c} /* (9, 4, 2) {real, imag} */,
  {32'hc0a9c914, 32'h421a78b0} /* (9, 4, 1) {real, imag} */,
  {32'h40a4cf58, 32'h41636e0a} /* (9, 4, 0) {real, imag} */,
  {32'hc04cfdc4, 32'h408dfca0} /* (9, 3, 31) {real, imag} */,
  {32'hc1122b38, 32'h4205ae60} /* (9, 3, 30) {real, imag} */,
  {32'h42cd0f2e, 32'h415bafac} /* (9, 3, 29) {real, imag} */,
  {32'hc01286a2, 32'h41d8efc0} /* (9, 3, 28) {real, imag} */,
  {32'h41ae67b6, 32'h41d5957c} /* (9, 3, 27) {real, imag} */,
  {32'h41d803a4, 32'hc281a2ec} /* (9, 3, 26) {real, imag} */,
  {32'h422113e7, 32'h42396f4f} /* (9, 3, 25) {real, imag} */,
  {32'hbe220e00, 32'h41467adc} /* (9, 3, 24) {real, imag} */,
  {32'hc1d9d8df, 32'hc2993b7c} /* (9, 3, 23) {real, imag} */,
  {32'hc25977b8, 32'h3fcd2790} /* (9, 3, 22) {real, imag} */,
  {32'h41115f24, 32'hc1981598} /* (9, 3, 21) {real, imag} */,
  {32'h40174db4, 32'h419aa43a} /* (9, 3, 20) {real, imag} */,
  {32'h420c92c4, 32'hc03e5fa0} /* (9, 3, 19) {real, imag} */,
  {32'hc20108b2, 32'h400dbbf0} /* (9, 3, 18) {real, imag} */,
  {32'h41e61d67, 32'hc0ec7df6} /* (9, 3, 17) {real, imag} */,
  {32'hc0945268, 32'h4130f8ae} /* (9, 3, 16) {real, imag} */,
  {32'hc115925a, 32'h41e2d80a} /* (9, 3, 15) {real, imag} */,
  {32'hc2145e06, 32'h414ebcbc} /* (9, 3, 14) {real, imag} */,
  {32'h41043e4f, 32'hc291026a} /* (9, 3, 13) {real, imag} */,
  {32'h41e71132, 32'hc1984cf4} /* (9, 3, 12) {real, imag} */,
  {32'hc142ba74, 32'h426ff774} /* (9, 3, 11) {real, imag} */,
  {32'hc05ba0a0, 32'h40affb1c} /* (9, 3, 10) {real, imag} */,
  {32'hc16886e2, 32'hbf9ce4a0} /* (9, 3, 9) {real, imag} */,
  {32'h42301fc2, 32'h413eadc4} /* (9, 3, 8) {real, imag} */,
  {32'hc247a229, 32'h423a0ff9} /* (9, 3, 7) {real, imag} */,
  {32'h42736f54, 32'hc2d8a940} /* (9, 3, 6) {real, imag} */,
  {32'h4294295e, 32'h41092591} /* (9, 3, 5) {real, imag} */,
  {32'hc13427aa, 32'h42b784da} /* (9, 3, 4) {real, imag} */,
  {32'h42aeea0c, 32'hc1e610f6} /* (9, 3, 3) {real, imag} */,
  {32'hc2b8755d, 32'hc324cae6} /* (9, 3, 2) {real, imag} */,
  {32'hc0f4c30e, 32'hc21d79d8} /* (9, 3, 1) {real, imag} */,
  {32'h42ad374a, 32'hc15184b8} /* (9, 3, 0) {real, imag} */,
  {32'h4201eff9, 32'hc2c2ab37} /* (9, 2, 31) {real, imag} */,
  {32'hc221ac6e, 32'h4326f769} /* (9, 2, 30) {real, imag} */,
  {32'hc3106e63, 32'h3dd41000} /* (9, 2, 29) {real, imag} */,
  {32'hc29a6a1b, 32'hc2e4c362} /* (9, 2, 28) {real, imag} */,
  {32'h3ff65e80, 32'h41ddc11d} /* (9, 2, 27) {real, imag} */,
  {32'h4219d92a, 32'h429d503c} /* (9, 2, 26) {real, imag} */,
  {32'h41847c64, 32'h4253d8ac} /* (9, 2, 25) {real, imag} */,
  {32'hc1e72e50, 32'hc17d52d8} /* (9, 2, 24) {real, imag} */,
  {32'hc1a81616, 32'hc19b6ce2} /* (9, 2, 23) {real, imag} */,
  {32'h42840df2, 32'h41c8eb4c} /* (9, 2, 22) {real, imag} */,
  {32'h41ecb7c8, 32'h416291ca} /* (9, 2, 21) {real, imag} */,
  {32'h40a9e132, 32'hc2147660} /* (9, 2, 20) {real, imag} */,
  {32'hc2398898, 32'h41a3ed42} /* (9, 2, 19) {real, imag} */,
  {32'h4187c3f5, 32'h42123996} /* (9, 2, 18) {real, imag} */,
  {32'hc0f4da68, 32'h408a36b4} /* (9, 2, 17) {real, imag} */,
  {32'h419e51ac, 32'hc0837470} /* (9, 2, 16) {real, imag} */,
  {32'h421d294a, 32'h42013f3c} /* (9, 2, 15) {real, imag} */,
  {32'h4207a9f0, 32'hc0e76ed4} /* (9, 2, 14) {real, imag} */,
  {32'hc1427b88, 32'hc181aefa} /* (9, 2, 13) {real, imag} */,
  {32'h41915308, 32'hc10cacba} /* (9, 2, 12) {real, imag} */,
  {32'hc252b3a4, 32'hc1cb7fa3} /* (9, 2, 11) {real, imag} */,
  {32'h424d0138, 32'h42391f38} /* (9, 2, 10) {real, imag} */,
  {32'hbfd72d00, 32'hc1ff1524} /* (9, 2, 9) {real, imag} */,
  {32'hc29cdff0, 32'h41cce74c} /* (9, 2, 8) {real, imag} */,
  {32'h42d03b41, 32'hc1b634c7} /* (9, 2, 7) {real, imag} */,
  {32'h42837eb1, 32'h42017d63} /* (9, 2, 6) {real, imag} */,
  {32'hc28fd89e, 32'hc1f0a673} /* (9, 2, 5) {real, imag} */,
  {32'h4250b09a, 32'hc2f63806} /* (9, 2, 4) {real, imag} */,
  {32'hc277e92b, 32'h42d2c36f} /* (9, 2, 3) {real, imag} */,
  {32'h4245b65c, 32'h4351139b} /* (9, 2, 2) {real, imag} */,
  {32'h42cf3a32, 32'hc2e4516d} /* (9, 2, 1) {real, imag} */,
  {32'h41b9cd2e, 32'hc2e7fe0b} /* (9, 2, 0) {real, imag} */,
  {32'hc202ab66, 32'h42f0fe5e} /* (9, 1, 31) {real, imag} */,
  {32'h428ed470, 32'hc2c1af67} /* (9, 1, 30) {real, imag} */,
  {32'h40a75892, 32'hc0114c20} /* (9, 1, 29) {real, imag} */,
  {32'hbf08e4f0, 32'h421c6b19} /* (9, 1, 28) {real, imag} */,
  {32'h41c3cf5a, 32'h4229bd0d} /* (9, 1, 27) {real, imag} */,
  {32'hc2d3856b, 32'h42988cf0} /* (9, 1, 26) {real, imag} */,
  {32'hc285fbd1, 32'h41efd61e} /* (9, 1, 25) {real, imag} */,
  {32'h418899ba, 32'hc1ecde22} /* (9, 1, 24) {real, imag} */,
  {32'h40d71210, 32'hc20002ef} /* (9, 1, 23) {real, imag} */,
  {32'h423bd214, 32'hc1d1b4ae} /* (9, 1, 22) {real, imag} */,
  {32'h41f7736d, 32'h4115ecaf} /* (9, 1, 21) {real, imag} */,
  {32'hc248cfa4, 32'hc133029d} /* (9, 1, 20) {real, imag} */,
  {32'h41b9b3d2, 32'hc1ce8b96} /* (9, 1, 19) {real, imag} */,
  {32'h4148d9ee, 32'hc14d3087} /* (9, 1, 18) {real, imag} */,
  {32'h4111e368, 32'h419ba860} /* (9, 1, 17) {real, imag} */,
  {32'h41276b58, 32'hc1e47d4e} /* (9, 1, 16) {real, imag} */,
  {32'h411af648, 32'hbfa21940} /* (9, 1, 15) {real, imag} */,
  {32'hc1a8b187, 32'hc1245951} /* (9, 1, 14) {real, imag} */,
  {32'hc0ad1ffa, 32'hc22957ff} /* (9, 1, 13) {real, imag} */,
  {32'hc1995747, 32'h40eabd6a} /* (9, 1, 12) {real, imag} */,
  {32'hc1cfbe1f, 32'hbf0a3150} /* (9, 1, 11) {real, imag} */,
  {32'hc1f64088, 32'h420ccac3} /* (9, 1, 10) {real, imag} */,
  {32'h41e99e8c, 32'h427af767} /* (9, 1, 9) {real, imag} */,
  {32'hc28bba62, 32'h430a86db} /* (9, 1, 8) {real, imag} */,
  {32'h4242625e, 32'h4224cee5} /* (9, 1, 7) {real, imag} */,
  {32'h422ef702, 32'hc2248e45} /* (9, 1, 6) {real, imag} */,
  {32'h42905610, 32'hc1550ecf} /* (9, 1, 5) {real, imag} */,
  {32'hc18780aa, 32'h4283491d} /* (9, 1, 4) {real, imag} */,
  {32'h413a2da7, 32'hc37a1e60} /* (9, 1, 3) {real, imag} */,
  {32'h43163f25, 32'hc2da83ad} /* (9, 1, 2) {real, imag} */,
  {32'hc320011c, 32'hc1373994} /* (9, 1, 1) {real, imag} */,
  {32'hc312e8dc, 32'hc2857d40} /* (9, 1, 0) {real, imag} */,
  {32'hc27b2318, 32'h42e71cb2} /* (9, 0, 31) {real, imag} */,
  {32'h41fae6d4, 32'hc1d20c4b} /* (9, 0, 30) {real, imag} */,
  {32'hc29bfccc, 32'h418a9164} /* (9, 0, 29) {real, imag} */,
  {32'h424e5482, 32'h411d796c} /* (9, 0, 28) {real, imag} */,
  {32'h424a25c1, 32'hc106bafe} /* (9, 0, 27) {real, imag} */,
  {32'hc28c67e7, 32'h4181a3d8} /* (9, 0, 26) {real, imag} */,
  {32'h4178c072, 32'h4203b7f8} /* (9, 0, 25) {real, imag} */,
  {32'hc298721b, 32'hc2aa85a8} /* (9, 0, 24) {real, imag} */,
  {32'h41a55593, 32'hc27ca8b9} /* (9, 0, 23) {real, imag} */,
  {32'h42bb3720, 32'hc18d606c} /* (9, 0, 22) {real, imag} */,
  {32'hc19f471a, 32'h403dedf8} /* (9, 0, 21) {real, imag} */,
  {32'h402ca36e, 32'hbf308b70} /* (9, 0, 20) {real, imag} */,
  {32'h421a8a1d, 32'hc11a283b} /* (9, 0, 19) {real, imag} */,
  {32'hc19f61b8, 32'hc16cabd1} /* (9, 0, 18) {real, imag} */,
  {32'hc104a436, 32'h4102a1ea} /* (9, 0, 17) {real, imag} */,
  {32'h40f3aeca, 32'hc1c0dff0} /* (9, 0, 16) {real, imag} */,
  {32'hc0702b48, 32'hc1252876} /* (9, 0, 15) {real, imag} */,
  {32'h419b6748, 32'h41d51116} /* (9, 0, 14) {real, imag} */,
  {32'hc1e9a5e6, 32'h4123d985} /* (9, 0, 13) {real, imag} */,
  {32'h40c1776f, 32'h418c4a10} /* (9, 0, 12) {real, imag} */,
  {32'hc16be6fc, 32'hc22f80c8} /* (9, 0, 11) {real, imag} */,
  {32'hc1f0ff1a, 32'h4225af46} /* (9, 0, 10) {real, imag} */,
  {32'h41eadff5, 32'hc0c4b7e8} /* (9, 0, 9) {real, imag} */,
  {32'h42a7e8cd, 32'h430b6576} /* (9, 0, 8) {real, imag} */,
  {32'hc2345e58, 32'h424c003a} /* (9, 0, 7) {real, imag} */,
  {32'hc17ece3e, 32'hc28f13c2} /* (9, 0, 6) {real, imag} */,
  {32'h4284656e, 32'hc22cb3f0} /* (9, 0, 5) {real, imag} */,
  {32'hc2958a7d, 32'h42815db2} /* (9, 0, 4) {real, imag} */,
  {32'h4319e11e, 32'hc16bf247} /* (9, 0, 3) {real, imag} */,
  {32'hc26499ea, 32'hc167d9aa} /* (9, 0, 2) {real, imag} */,
  {32'hc307a91e, 32'hc283d1b6} /* (9, 0, 1) {real, imag} */,
  {32'hc1a5d9aa, 32'h43401eb6} /* (9, 0, 0) {real, imag} */,
  {32'hc31ab97c, 32'h443b155e} /* (8, 31, 31) {real, imag} */,
  {32'hc25d46f4, 32'hc3f7ccaf} /* (8, 31, 30) {real, imag} */,
  {32'hc0c97524, 32'h419c4a48} /* (8, 31, 29) {real, imag} */,
  {32'h42bb06e9, 32'hc293abfe} /* (8, 31, 28) {real, imag} */,
  {32'h41c960d2, 32'hc3029a02} /* (8, 31, 27) {real, imag} */,
  {32'hc145625e, 32'h40bfcad4} /* (8, 31, 26) {real, imag} */,
  {32'hc20b76f8, 32'h40cbae50} /* (8, 31, 25) {real, imag} */,
  {32'hc2a5d7a2, 32'hc2df64de} /* (8, 31, 24) {real, imag} */,
  {32'hc29b417e, 32'hc1c8d134} /* (8, 31, 23) {real, imag} */,
  {32'h42935904, 32'h42664dac} /* (8, 31, 22) {real, imag} */,
  {32'h40aa6c6a, 32'hc297607b} /* (8, 31, 21) {real, imag} */,
  {32'hc232ed58, 32'hc0893718} /* (8, 31, 20) {real, imag} */,
  {32'hc05ec7d8, 32'h41b7875c} /* (8, 31, 19) {real, imag} */,
  {32'hc17f9a18, 32'h3e932500} /* (8, 31, 18) {real, imag} */,
  {32'h42a08d6a, 32'hbfbe8880} /* (8, 31, 17) {real, imag} */,
  {32'hc1a37950, 32'h41a82598} /* (8, 31, 16) {real, imag} */,
  {32'hc164f534, 32'hc1790630} /* (8, 31, 15) {real, imag} */,
  {32'h417eb598, 32'h427f34c6} /* (8, 31, 14) {real, imag} */,
  {32'h401b2dc0, 32'hc1ddd03c} /* (8, 31, 13) {real, imag} */,
  {32'h40a61de0, 32'h41b50eba} /* (8, 31, 12) {real, imag} */,
  {32'hc1a9a0aa, 32'h41e02abc} /* (8, 31, 11) {real, imag} */,
  {32'hc0ab4ac0, 32'h3ffae2b0} /* (8, 31, 10) {real, imag} */,
  {32'h418970c4, 32'hc2c5c97a} /* (8, 31, 9) {real, imag} */,
  {32'h4171a1f0, 32'h42291984} /* (8, 31, 8) {real, imag} */,
  {32'h42a00209, 32'h41634290} /* (8, 31, 7) {real, imag} */,
  {32'hc2799760, 32'hc1907299} /* (8, 31, 6) {real, imag} */,
  {32'h428b0384, 32'hc334eb20} /* (8, 31, 5) {real, imag} */,
  {32'h421c0c9e, 32'h42d48b9a} /* (8, 31, 4) {real, imag} */,
  {32'h41c0f28c, 32'hc1b6a390} /* (8, 31, 3) {real, imag} */,
  {32'h43561667, 32'hc3199e66} /* (8, 31, 2) {real, imag} */,
  {32'hc38e6341, 32'h4395bcc4} /* (8, 31, 1) {real, imag} */,
  {32'hc36ef09c, 32'h43e34c68} /* (8, 31, 0) {real, imag} */,
  {32'h439f9f65, 32'hc2071f3c} /* (8, 30, 31) {real, imag} */,
  {32'hc39d2d91, 32'h43c3518d} /* (8, 30, 30) {real, imag} */,
  {32'h42da04f0, 32'h4217dad0} /* (8, 30, 29) {real, imag} */,
  {32'h42e97562, 32'hc250f012} /* (8, 30, 28) {real, imag} */,
  {32'h42832198, 32'h43416ac8} /* (8, 30, 27) {real, imag} */,
  {32'h40ad6e90, 32'h4180a6e8} /* (8, 30, 26) {real, imag} */,
  {32'hc2148475, 32'h428d4496} /* (8, 30, 25) {real, imag} */,
  {32'hc1473310, 32'h42d1d10c} /* (8, 30, 24) {real, imag} */,
  {32'hbff704a0, 32'hc1bc109e} /* (8, 30, 23) {real, imag} */,
  {32'hc20dee6e, 32'h413163d8} /* (8, 30, 22) {real, imag} */,
  {32'h41a6ac77, 32'h410de65c} /* (8, 30, 21) {real, imag} */,
  {32'h423c9939, 32'hc23fba0e} /* (8, 30, 20) {real, imag} */,
  {32'h411d15f0, 32'hbf545020} /* (8, 30, 19) {real, imag} */,
  {32'hc09dee32, 32'hc0b49f00} /* (8, 30, 18) {real, imag} */,
  {32'hc12d5d0b, 32'h40996d00} /* (8, 30, 17) {real, imag} */,
  {32'h416d13b8, 32'hc19d37b0} /* (8, 30, 16) {real, imag} */,
  {32'hc0c6966a, 32'h3ea6ac00} /* (8, 30, 15) {real, imag} */,
  {32'h415567b9, 32'h41d92990} /* (8, 30, 14) {real, imag} */,
  {32'h42285d06, 32'h41eb853d} /* (8, 30, 13) {real, imag} */,
  {32'hc15ecdf4, 32'h4292de8f} /* (8, 30, 12) {real, imag} */,
  {32'h419a71ab, 32'hc197ed82} /* (8, 30, 11) {real, imag} */,
  {32'h41c748f4, 32'h41d59df4} /* (8, 30, 10) {real, imag} */,
  {32'hc1ec55f2, 32'hc1ca82e2} /* (8, 30, 9) {real, imag} */,
  {32'hc330fd1d, 32'h41d6d748} /* (8, 30, 8) {real, imag} */,
  {32'h4196f4a6, 32'hc0c22e98} /* (8, 30, 7) {real, imag} */,
  {32'h429e9253, 32'hc2fb174a} /* (8, 30, 6) {real, imag} */,
  {32'hc32ebb96, 32'h41b85d9c} /* (8, 30, 5) {real, imag} */,
  {32'h4242f6b3, 32'h424e8296} /* (8, 30, 4) {real, imag} */,
  {32'h42a78328, 32'hc2447754} /* (8, 30, 3) {real, imag} */,
  {32'hc3823403, 32'h42b4e650} /* (8, 30, 2) {real, imag} */,
  {32'h43888517, 32'hc3f40070} /* (8, 30, 1) {real, imag} */,
  {32'h42fc42b5, 32'hc38b19a9} /* (8, 30, 0) {real, imag} */,
  {32'hc213488d, 32'h4290a558} /* (8, 29, 31) {real, imag} */,
  {32'hc2845e41, 32'hc23364bd} /* (8, 29, 30) {real, imag} */,
  {32'h42d877de, 32'hc2cfc0d9} /* (8, 29, 29) {real, imag} */,
  {32'h42820570, 32'hc281e138} /* (8, 29, 28) {real, imag} */,
  {32'h416e6564, 32'h428fe0a8} /* (8, 29, 27) {real, imag} */,
  {32'hc252a4b3, 32'hc0da3848} /* (8, 29, 26) {real, imag} */,
  {32'hc24dac52, 32'h40d447ec} /* (8, 29, 25) {real, imag} */,
  {32'h422ccf68, 32'hc04b73b0} /* (8, 29, 24) {real, imag} */,
  {32'h412a857a, 32'h3fcd9e60} /* (8, 29, 23) {real, imag} */,
  {32'h41089b06, 32'h4153c0aa} /* (8, 29, 22) {real, imag} */,
  {32'hc12a61bc, 32'h418136d8} /* (8, 29, 21) {real, imag} */,
  {32'hc20fbf48, 32'hc258cd68} /* (8, 29, 20) {real, imag} */,
  {32'hc22a7df5, 32'hc1b44c9c} /* (8, 29, 19) {real, imag} */,
  {32'h40866b40, 32'h422c8c76} /* (8, 29, 18) {real, imag} */,
  {32'h419988c8, 32'hc225bc15} /* (8, 29, 17) {real, imag} */,
  {32'hc17474e4, 32'hc1292e52} /* (8, 29, 16) {real, imag} */,
  {32'h40028320, 32'hc199cea6} /* (8, 29, 15) {real, imag} */,
  {32'hc22e575b, 32'h41fac21f} /* (8, 29, 14) {real, imag} */,
  {32'hc1ccacfe, 32'h4134c978} /* (8, 29, 13) {real, imag} */,
  {32'hc0587b88, 32'hc20419a8} /* (8, 29, 12) {real, imag} */,
  {32'hc25662df, 32'h4221d8d2} /* (8, 29, 11) {real, imag} */,
  {32'h428ead30, 32'hbfb42ab0} /* (8, 29, 10) {real, imag} */,
  {32'h41a8b8af, 32'hc264496f} /* (8, 29, 9) {real, imag} */,
  {32'hc22e1450, 32'hc29ef616} /* (8, 29, 8) {real, imag} */,
  {32'hc237adf0, 32'hc1b0985a} /* (8, 29, 7) {real, imag} */,
  {32'h42cfefac, 32'h429edd44} /* (8, 29, 6) {real, imag} */,
  {32'h428f55ea, 32'h3f8d1cc0} /* (8, 29, 5) {real, imag} */,
  {32'h4222bfff, 32'h433c18ba} /* (8, 29, 4) {real, imag} */,
  {32'hc2a6f816, 32'hc346c4e4} /* (8, 29, 3) {real, imag} */,
  {32'hc270f4b2, 32'h425a3bc7} /* (8, 29, 2) {real, imag} */,
  {32'h43101fff, 32'h419d0d6e} /* (8, 29, 1) {real, imag} */,
  {32'h42859d64, 32'h41f37221} /* (8, 29, 0) {real, imag} */,
  {32'hc25a57ad, 32'h435baea4} /* (8, 28, 31) {real, imag} */,
  {32'hc2821360, 32'hc330f383} /* (8, 28, 30) {real, imag} */,
  {32'hc201e9d5, 32'h430e46a4} /* (8, 28, 29) {real, imag} */,
  {32'h42bc900c, 32'h42ed015a} /* (8, 28, 28) {real, imag} */,
  {32'h420e3495, 32'hc0fd4e50} /* (8, 28, 27) {real, imag} */,
  {32'h41633fe6, 32'h4164e30c} /* (8, 28, 26) {real, imag} */,
  {32'h419c011b, 32'h43037fdc} /* (8, 28, 25) {real, imag} */,
  {32'h4106a922, 32'hc09ab754} /* (8, 28, 24) {real, imag} */,
  {32'hc2d8f711, 32'hc22af942} /* (8, 28, 23) {real, imag} */,
  {32'h42002b24, 32'hc1326cbc} /* (8, 28, 22) {real, imag} */,
  {32'hc2818b92, 32'hc299272c} /* (8, 28, 21) {real, imag} */,
  {32'hc1865bf2, 32'h419d2302} /* (8, 28, 20) {real, imag} */,
  {32'h419366c8, 32'h41c886af} /* (8, 28, 19) {real, imag} */,
  {32'hc03b7150, 32'hc2124f36} /* (8, 28, 18) {real, imag} */,
  {32'h40c32c1e, 32'hc0edfd20} /* (8, 28, 17) {real, imag} */,
  {32'h408da71c, 32'h414063fe} /* (8, 28, 16) {real, imag} */,
  {32'hc11cceb9, 32'hc1bfdd70} /* (8, 28, 15) {real, imag} */,
  {32'hc1b25dfe, 32'hc1ea47a3} /* (8, 28, 14) {real, imag} */,
  {32'h412eae60, 32'h41690f32} /* (8, 28, 13) {real, imag} */,
  {32'hc11afb55, 32'hc1a907ba} /* (8, 28, 12) {real, imag} */,
  {32'hc167e050, 32'h4128e38c} /* (8, 28, 11) {real, imag} */,
  {32'h40f40074, 32'h4225a804} /* (8, 28, 10) {real, imag} */,
  {32'h41c761d4, 32'h41a15eb3} /* (8, 28, 9) {real, imag} */,
  {32'h4262a30c, 32'h41c807d1} /* (8, 28, 8) {real, imag} */,
  {32'h42066ff2, 32'hc02e94a0} /* (8, 28, 7) {real, imag} */,
  {32'h41dea777, 32'hc1704430} /* (8, 28, 6) {real, imag} */,
  {32'h411584d4, 32'h43363cf8} /* (8, 28, 5) {real, imag} */,
  {32'hc256a5fc, 32'h3ffd90e0} /* (8, 28, 4) {real, imag} */,
  {32'h421519bb, 32'h43111a58} /* (8, 28, 3) {real, imag} */,
  {32'h4210eeda, 32'hc32f9cbb} /* (8, 28, 2) {real, imag} */,
  {32'hc02d9b10, 32'h42951729} /* (8, 28, 1) {real, imag} */,
  {32'hc08d35bc, 32'h41d48d9d} /* (8, 28, 0) {real, imag} */,
  {32'hc2498d3e, 32'hc1d4dc76} /* (8, 27, 31) {real, imag} */,
  {32'h41fdf38c, 32'h42bc3380} /* (8, 27, 30) {real, imag} */,
  {32'h40a15212, 32'hbf0b3a00} /* (8, 27, 29) {real, imag} */,
  {32'h42a24525, 32'h42c69a94} /* (8, 27, 28) {real, imag} */,
  {32'h4202e055, 32'hc04cb670} /* (8, 27, 27) {real, imag} */,
  {32'h41bba392, 32'hc09e5190} /* (8, 27, 26) {real, imag} */,
  {32'hc28d5ad3, 32'hc20d851b} /* (8, 27, 25) {real, imag} */,
  {32'h42779066, 32'h42332e6d} /* (8, 27, 24) {real, imag} */,
  {32'h41688116, 32'hc1875d24} /* (8, 27, 23) {real, imag} */,
  {32'hc13893c7, 32'h3e8f9d70} /* (8, 27, 22) {real, imag} */,
  {32'h41aabec6, 32'h40f5ee30} /* (8, 27, 21) {real, imag} */,
  {32'h423ef5b4, 32'hc0ba8e10} /* (8, 27, 20) {real, imag} */,
  {32'hc2824a00, 32'h40b24264} /* (8, 27, 19) {real, imag} */,
  {32'hc18bd2cd, 32'hc1a1b507} /* (8, 27, 18) {real, imag} */,
  {32'hc0ee0ca9, 32'h41d3779f} /* (8, 27, 17) {real, imag} */,
  {32'h41c4836e, 32'hc256b5fa} /* (8, 27, 16) {real, imag} */,
  {32'hc0f541e9, 32'h4125b7aa} /* (8, 27, 15) {real, imag} */,
  {32'hc196f8a3, 32'hc1a6af55} /* (8, 27, 14) {real, imag} */,
  {32'hc0994038, 32'h411b4984} /* (8, 27, 13) {real, imag} */,
  {32'hc1b5a9f7, 32'hc1056e10} /* (8, 27, 12) {real, imag} */,
  {32'h41234873, 32'hc23372ee} /* (8, 27, 11) {real, imag} */,
  {32'hbf799470, 32'h40839e7d} /* (8, 27, 10) {real, imag} */,
  {32'h41462c66, 32'h3ff5edc8} /* (8, 27, 9) {real, imag} */,
  {32'hc1dbb600, 32'h41c00a36} /* (8, 27, 8) {real, imag} */,
  {32'h4270b5e3, 32'hc1c3fcb9} /* (8, 27, 7) {real, imag} */,
  {32'hc1ebacbe, 32'hc1ed3dd4} /* (8, 27, 6) {real, imag} */,
  {32'hc289fa0e, 32'hc20570e3} /* (8, 27, 5) {real, imag} */,
  {32'h424a3536, 32'h413c6a9c} /* (8, 27, 4) {real, imag} */,
  {32'h41b1f7b2, 32'hc1257f1e} /* (8, 27, 3) {real, imag} */,
  {32'hc253b0ca, 32'h42b26ddc} /* (8, 27, 2) {real, imag} */,
  {32'h42696196, 32'hc2b69e98} /* (8, 27, 1) {real, imag} */,
  {32'h41c1ab32, 32'hc2929991} /* (8, 27, 0) {real, imag} */,
  {32'h419d8c26, 32'h42a99431} /* (8, 26, 31) {real, imag} */,
  {32'h41b6bed3, 32'hc13cc094} /* (8, 26, 30) {real, imag} */,
  {32'h429b7592, 32'h41e017f9} /* (8, 26, 29) {real, imag} */,
  {32'h427a2418, 32'hc1904e32} /* (8, 26, 28) {real, imag} */,
  {32'h41008ce0, 32'h42d456ac} /* (8, 26, 27) {real, imag} */,
  {32'h41ce4340, 32'h421eb387} /* (8, 26, 26) {real, imag} */,
  {32'hbf8a6940, 32'hc2b27ad0} /* (8, 26, 25) {real, imag} */,
  {32'hc193adcd, 32'hc0264f18} /* (8, 26, 24) {real, imag} */,
  {32'h40901166, 32'hc16e5ca4} /* (8, 26, 23) {real, imag} */,
  {32'hc22a8e2e, 32'hc25a4c80} /* (8, 26, 22) {real, imag} */,
  {32'hc2854355, 32'hc1a35809} /* (8, 26, 21) {real, imag} */,
  {32'h416c6d22, 32'hc185cf78} /* (8, 26, 20) {real, imag} */,
  {32'h41ba1fd8, 32'h400dbe58} /* (8, 26, 19) {real, imag} */,
  {32'h415cbe66, 32'h3f0671c0} /* (8, 26, 18) {real, imag} */,
  {32'h4114d6de, 32'h41ad7bb1} /* (8, 26, 17) {real, imag} */,
  {32'hc01612b0, 32'h408feb3a} /* (8, 26, 16) {real, imag} */,
  {32'h412920b2, 32'hc09a6a14} /* (8, 26, 15) {real, imag} */,
  {32'hc1f1ebbf, 32'h418f998a} /* (8, 26, 14) {real, imag} */,
  {32'h424f5a3c, 32'hc21b3040} /* (8, 26, 13) {real, imag} */,
  {32'hc0e30984, 32'h41dda56c} /* (8, 26, 12) {real, imag} */,
  {32'h413cb83a, 32'h416efa4e} /* (8, 26, 11) {real, imag} */,
  {32'hc16b3910, 32'h422efd18} /* (8, 26, 10) {real, imag} */,
  {32'hc1f4b3d2, 32'h41ae4b26} /* (8, 26, 9) {real, imag} */,
  {32'hc25e7616, 32'h4212b9a2} /* (8, 26, 8) {real, imag} */,
  {32'hc19bc11b, 32'hc28e4dbc} /* (8, 26, 7) {real, imag} */,
  {32'hc298110f, 32'hc1ab0742} /* (8, 26, 6) {real, imag} */,
  {32'h42dcaf76, 32'hc1efcde0} /* (8, 26, 5) {real, imag} */,
  {32'h42c03230, 32'hc2fcbf34} /* (8, 26, 4) {real, imag} */,
  {32'h4258d32d, 32'h41e69999} /* (8, 26, 3) {real, imag} */,
  {32'hbf395c60, 32'hc307ecc8} /* (8, 26, 2) {real, imag} */,
  {32'hc2d156a4, 32'h42112804} /* (8, 26, 1) {real, imag} */,
  {32'hc28caeb0, 32'h410d48e9} /* (8, 26, 0) {real, imag} */,
  {32'h42257077, 32'hc00aba38} /* (8, 25, 31) {real, imag} */,
  {32'hc1bb003a, 32'h41b08edc} /* (8, 25, 30) {real, imag} */,
  {32'hc2cc5516, 32'hc0fa43f4} /* (8, 25, 29) {real, imag} */,
  {32'h419472d9, 32'hc1a5b038} /* (8, 25, 28) {real, imag} */,
  {32'h4226bce5, 32'hc2b7cdd3} /* (8, 25, 27) {real, imag} */,
  {32'hc2bfd08a, 32'h42315e5e} /* (8, 25, 26) {real, imag} */,
  {32'h41cc1a9f, 32'h40a1a4ec} /* (8, 25, 25) {real, imag} */,
  {32'hc19870c5, 32'hc20c10b2} /* (8, 25, 24) {real, imag} */,
  {32'hc1b9559e, 32'hc0ce2238} /* (8, 25, 23) {real, imag} */,
  {32'h4236f2d8, 32'h41eb0e28} /* (8, 25, 22) {real, imag} */,
  {32'h41094f69, 32'h41a55771} /* (8, 25, 21) {real, imag} */,
  {32'hc0c3d700, 32'hc141887c} /* (8, 25, 20) {real, imag} */,
  {32'hc14e3644, 32'h41cd2879} /* (8, 25, 19) {real, imag} */,
  {32'h41c291e4, 32'h4187569d} /* (8, 25, 18) {real, imag} */,
  {32'hc0af7d4c, 32'h40a8a514} /* (8, 25, 17) {real, imag} */,
  {32'h3f25fe20, 32'h41ade55e} /* (8, 25, 16) {real, imag} */,
  {32'hc13dc232, 32'hc10df0ec} /* (8, 25, 15) {real, imag} */,
  {32'hc0b04fbe, 32'hc0948e74} /* (8, 25, 14) {real, imag} */,
  {32'h4139572c, 32'h408ce9cc} /* (8, 25, 13) {real, imag} */,
  {32'hc1dd5002, 32'hc23daee9} /* (8, 25, 12) {real, imag} */,
  {32'hc18348cc, 32'h41193f92} /* (8, 25, 11) {real, imag} */,
  {32'hc12b41c6, 32'h424fc0fe} /* (8, 25, 10) {real, imag} */,
  {32'h423df1ad, 32'h41b3fb34} /* (8, 25, 9) {real, imag} */,
  {32'h4288010c, 32'hc1d1bdb9} /* (8, 25, 8) {real, imag} */,
  {32'h4276d96e, 32'hc281fd65} /* (8, 25, 7) {real, imag} */,
  {32'h41a5284a, 32'h42a9ccd5} /* (8, 25, 6) {real, imag} */,
  {32'hc1310274, 32'h42b22213} /* (8, 25, 5) {real, imag} */,
  {32'hc25d543c, 32'h428d45ec} /* (8, 25, 4) {real, imag} */,
  {32'h427059b8, 32'h4210220e} /* (8, 25, 3) {real, imag} */,
  {32'h4240a155, 32'hc2eb0cb7} /* (8, 25, 2) {real, imag} */,
  {32'hc23ee345, 32'hc1b28804} /* (8, 25, 1) {real, imag} */,
  {32'hc23a2ade, 32'h42f3bed4} /* (8, 25, 0) {real, imag} */,
  {32'h427e1188, 32'hc31da0a1} /* (8, 24, 31) {real, imag} */,
  {32'hc115f1c4, 32'h428e6564} /* (8, 24, 30) {real, imag} */,
  {32'hc2c04b40, 32'hc220f050} /* (8, 24, 29) {real, imag} */,
  {32'h42332f05, 32'h4194ec20} /* (8, 24, 28) {real, imag} */,
  {32'h40a6abd0, 32'h429e2490} /* (8, 24, 27) {real, imag} */,
  {32'h40b5cbe0, 32'h42270d86} /* (8, 24, 26) {real, imag} */,
  {32'hc2a99553, 32'hc0bc7d36} /* (8, 24, 25) {real, imag} */,
  {32'h420485c0, 32'hc1365f68} /* (8, 24, 24) {real, imag} */,
  {32'hc1af7f08, 32'hc23ce6aa} /* (8, 24, 23) {real, imag} */,
  {32'h41685a74, 32'h417dc720} /* (8, 24, 22) {real, imag} */,
  {32'h40f7f897, 32'hc1a6466f} /* (8, 24, 21) {real, imag} */,
  {32'h40f292b0, 32'hc144f32e} /* (8, 24, 20) {real, imag} */,
  {32'h41b0672c, 32'hc1edd74f} /* (8, 24, 19) {real, imag} */,
  {32'h4121bf6a, 32'hc1923866} /* (8, 24, 18) {real, imag} */,
  {32'hc074543c, 32'hc179a50a} /* (8, 24, 17) {real, imag} */,
  {32'hbea2f600, 32'h417dc31a} /* (8, 24, 16) {real, imag} */,
  {32'h412d183d, 32'hbffa7cac} /* (8, 24, 15) {real, imag} */,
  {32'h411ccf5e, 32'hc05d1eb0} /* (8, 24, 14) {real, imag} */,
  {32'hc12b8438, 32'h417a1912} /* (8, 24, 13) {real, imag} */,
  {32'h41998c81, 32'h4119e8c6} /* (8, 24, 12) {real, imag} */,
  {32'hc09d5c21, 32'hc0999134} /* (8, 24, 11) {real, imag} */,
  {32'hc1a0ab22, 32'hc163e99a} /* (8, 24, 10) {real, imag} */,
  {32'h414d02e0, 32'h3eb118c0} /* (8, 24, 9) {real, imag} */,
  {32'hc2a97062, 32'hc002b59a} /* (8, 24, 8) {real, imag} */,
  {32'hc27647ce, 32'hc141c431} /* (8, 24, 7) {real, imag} */,
  {32'h42208904, 32'h40804de0} /* (8, 24, 6) {real, imag} */,
  {32'hc2137dcd, 32'h42108789} /* (8, 24, 5) {real, imag} */,
  {32'h42306d2f, 32'h42e936fc} /* (8, 24, 4) {real, imag} */,
  {32'h428e993a, 32'hc2aa9d28} /* (8, 24, 3) {real, imag} */,
  {32'hc2cd8a2c, 32'h43160bc6} /* (8, 24, 2) {real, imag} */,
  {32'h400a16f8, 32'hc3294d79} /* (8, 24, 1) {real, imag} */,
  {32'h42883bf6, 32'hc1eb84f1} /* (8, 24, 0) {real, imag} */,
  {32'hc1d1aa47, 32'hc2ad844a} /* (8, 23, 31) {real, imag} */,
  {32'hc1bf2361, 32'hc29d4d69} /* (8, 23, 30) {real, imag} */,
  {32'h414221b8, 32'h424f2795} /* (8, 23, 29) {real, imag} */,
  {32'h422d04e8, 32'h4088b4e0} /* (8, 23, 28) {real, imag} */,
  {32'h4082bc10, 32'hc14f56b8} /* (8, 23, 27) {real, imag} */,
  {32'h417ba8a9, 32'hc141b4ca} /* (8, 23, 26) {real, imag} */,
  {32'h4200288a, 32'hc1b995c4} /* (8, 23, 25) {real, imag} */,
  {32'hc1118e6e, 32'hc10758a8} /* (8, 23, 24) {real, imag} */,
  {32'h40d812cc, 32'hc1ebe703} /* (8, 23, 23) {real, imag} */,
  {32'hc1560787, 32'h417c38b8} /* (8, 23, 22) {real, imag} */,
  {32'h40a621cc, 32'h4213137b} /* (8, 23, 21) {real, imag} */,
  {32'h4104fda4, 32'h41b9d412} /* (8, 23, 20) {real, imag} */,
  {32'hc24db555, 32'h413f1ce2} /* (8, 23, 19) {real, imag} */,
  {32'h41a9cbed, 32'h4095d290} /* (8, 23, 18) {real, imag} */,
  {32'hbf9c9bc0, 32'h4130cc5a} /* (8, 23, 17) {real, imag} */,
  {32'hc1598689, 32'h4025c5f0} /* (8, 23, 16) {real, imag} */,
  {32'hc0274878, 32'h41ed0923} /* (8, 23, 15) {real, imag} */,
  {32'hc1b3fee7, 32'hc2598a9e} /* (8, 23, 14) {real, imag} */,
  {32'hc1a3a69a, 32'h412e8856} /* (8, 23, 13) {real, imag} */,
  {32'h41d258ea, 32'h4194fd62} /* (8, 23, 12) {real, imag} */,
  {32'h410f1e36, 32'h41e9493a} /* (8, 23, 11) {real, imag} */,
  {32'hc0a8846e, 32'h416816c4} /* (8, 23, 10) {real, imag} */,
  {32'hc1fa917d, 32'hc175593a} /* (8, 23, 9) {real, imag} */,
  {32'hc1e2ada5, 32'hc1de6900} /* (8, 23, 8) {real, imag} */,
  {32'h4122a364, 32'h422d8d92} /* (8, 23, 7) {real, imag} */,
  {32'hc185bbdc, 32'hc187ef8f} /* (8, 23, 6) {real, imag} */,
  {32'hc22ebd77, 32'hc22dbb4a} /* (8, 23, 5) {real, imag} */,
  {32'h40b726f0, 32'h423df9be} /* (8, 23, 4) {real, imag} */,
  {32'hc1c86444, 32'h423709a9} /* (8, 23, 3) {real, imag} */,
  {32'h41c992d3, 32'h42bf68a9} /* (8, 23, 2) {real, imag} */,
  {32'h3f222060, 32'hc2101cd8} /* (8, 23, 1) {real, imag} */,
  {32'hc0c281ba, 32'h42c1d8a8} /* (8, 23, 0) {real, imag} */,
  {32'hc1ca73a4, 32'hc192aabe} /* (8, 22, 31) {real, imag} */,
  {32'h4226af7d, 32'h40868868} /* (8, 22, 30) {real, imag} */,
  {32'h4205d47c, 32'h40ca6260} /* (8, 22, 29) {real, imag} */,
  {32'h4286430c, 32'h41695e22} /* (8, 22, 28) {real, imag} */,
  {32'hc07232b0, 32'h42c63d7b} /* (8, 22, 27) {real, imag} */,
  {32'hc18f587e, 32'hc1787f55} /* (8, 22, 26) {real, imag} */,
  {32'hc18ac4ea, 32'hc1dcd86d} /* (8, 22, 25) {real, imag} */,
  {32'hc1838028, 32'hc0c17210} /* (8, 22, 24) {real, imag} */,
  {32'h4163e38b, 32'hc1247942} /* (8, 22, 23) {real, imag} */,
  {32'h4179c5d9, 32'h41a5dd0a} /* (8, 22, 22) {real, imag} */,
  {32'hbec03ec0, 32'hc0d0970f} /* (8, 22, 21) {real, imag} */,
  {32'h415e4724, 32'h41d15763} /* (8, 22, 20) {real, imag} */,
  {32'h40ccde8f, 32'h40f392aa} /* (8, 22, 19) {real, imag} */,
  {32'hc165cb9f, 32'h4012f760} /* (8, 22, 18) {real, imag} */,
  {32'h40e36254, 32'hc19af9e2} /* (8, 22, 17) {real, imag} */,
  {32'hc14588a8, 32'hc197b7e2} /* (8, 22, 16) {real, imag} */,
  {32'h3f7971e0, 32'hc14144ac} /* (8, 22, 15) {real, imag} */,
  {32'hc0e0690e, 32'hc094e560} /* (8, 22, 14) {real, imag} */,
  {32'hbfe6dfe4, 32'h3f8d6c98} /* (8, 22, 13) {real, imag} */,
  {32'h41bdc3c0, 32'h3f3c6ce0} /* (8, 22, 12) {real, imag} */,
  {32'h41aa6279, 32'hbf0523f8} /* (8, 22, 11) {real, imag} */,
  {32'hc1ee17fc, 32'hc2261f18} /* (8, 22, 10) {real, imag} */,
  {32'h4188950e, 32'h41a24b6f} /* (8, 22, 9) {real, imag} */,
  {32'h41ea5818, 32'h4033ae88} /* (8, 22, 8) {real, imag} */,
  {32'hc1ec384e, 32'h418ee337} /* (8, 22, 7) {real, imag} */,
  {32'hc210bda5, 32'hc17ebd69} /* (8, 22, 6) {real, imag} */,
  {32'hc1ab7e32, 32'hc2a41555} /* (8, 22, 5) {real, imag} */,
  {32'h424c77a8, 32'h4234e15e} /* (8, 22, 4) {real, imag} */,
  {32'hc249460c, 32'hc1a5b249} /* (8, 22, 3) {real, imag} */,
  {32'hc20fd719, 32'hc2b3bd62} /* (8, 22, 2) {real, imag} */,
  {32'h42cfaf59, 32'h41d4407a} /* (8, 22, 1) {real, imag} */,
  {32'hc23beeae, 32'h428c4c20} /* (8, 22, 0) {real, imag} */,
  {32'hc2037628, 32'hc1e6960d} /* (8, 21, 31) {real, imag} */,
  {32'h41f5ce3b, 32'h41a12178} /* (8, 21, 30) {real, imag} */,
  {32'h4238ccc1, 32'h40342c2d} /* (8, 21, 29) {real, imag} */,
  {32'hc28b21b5, 32'h42a060de} /* (8, 21, 28) {real, imag} */,
  {32'hc1bcd526, 32'hc19ebfd7} /* (8, 21, 27) {real, imag} */,
  {32'hc0a8008e, 32'h40f4bc14} /* (8, 21, 26) {real, imag} */,
  {32'h41a8a873, 32'hc1c6728f} /* (8, 21, 25) {real, imag} */,
  {32'hc004b076, 32'hc12d715a} /* (8, 21, 24) {real, imag} */,
  {32'h3f903270, 32'h41280104} /* (8, 21, 23) {real, imag} */,
  {32'hc11c9f9e, 32'hc1a0c3b8} /* (8, 21, 22) {real, imag} */,
  {32'h416568ad, 32'h3fa15d90} /* (8, 21, 21) {real, imag} */,
  {32'hc1c6ef2a, 32'h4138c5be} /* (8, 21, 20) {real, imag} */,
  {32'h40984b32, 32'h400784d2} /* (8, 21, 19) {real, imag} */,
  {32'h3fb95fac, 32'h3d486180} /* (8, 21, 18) {real, imag} */,
  {32'h40a2ac56, 32'h40a3ece5} /* (8, 21, 17) {real, imag} */,
  {32'h411ece31, 32'hbf978a0c} /* (8, 21, 16) {real, imag} */,
  {32'hbffe0f5a, 32'h40065b56} /* (8, 21, 15) {real, imag} */,
  {32'h3fed5cb4, 32'h3f9ca684} /* (8, 21, 14) {real, imag} */,
  {32'hc0dac656, 32'hc149b3d8} /* (8, 21, 13) {real, imag} */,
  {32'hc10f83e0, 32'h3f5fd1a0} /* (8, 21, 12) {real, imag} */,
  {32'h419a990e, 32'h42196bb4} /* (8, 21, 11) {real, imag} */,
  {32'h41266e6e, 32'hbf4d1cd0} /* (8, 21, 10) {real, imag} */,
  {32'h41cb2f3f, 32'hc0701562} /* (8, 21, 9) {real, imag} */,
  {32'hc18b5a4e, 32'hc18f6977} /* (8, 21, 8) {real, imag} */,
  {32'hc1f11dc1, 32'hc113ea3a} /* (8, 21, 7) {real, imag} */,
  {32'hc07f6e90, 32'h422e7e7a} /* (8, 21, 6) {real, imag} */,
  {32'h4152ea33, 32'hbf2f23a0} /* (8, 21, 5) {real, imag} */,
  {32'h3f99f5c0, 32'hc2204229} /* (8, 21, 4) {real, imag} */,
  {32'hc1aa676e, 32'hc0a6fdf8} /* (8, 21, 3) {real, imag} */,
  {32'h402d1858, 32'h41d2bbac} /* (8, 21, 2) {real, imag} */,
  {32'h41ed1330, 32'hc222bb48} /* (8, 21, 1) {real, imag} */,
  {32'hc11c1fd3, 32'hc02aedfa} /* (8, 21, 0) {real, imag} */,
  {32'h420b80dc, 32'hc1cd948e} /* (8, 20, 31) {real, imag} */,
  {32'h419a92d6, 32'hc20d3ba6} /* (8, 20, 30) {real, imag} */,
  {32'hc0c5a17c, 32'h41d9b3da} /* (8, 20, 29) {real, imag} */,
  {32'hc1d5dc1f, 32'hc1bcfd71} /* (8, 20, 28) {real, imag} */,
  {32'hc1b3ea0f, 32'h416ccb7d} /* (8, 20, 27) {real, imag} */,
  {32'h418b7903, 32'hc1152907} /* (8, 20, 26) {real, imag} */,
  {32'hc0b64dcc, 32'h422ce671} /* (8, 20, 25) {real, imag} */,
  {32'h412a10c8, 32'hc116bf3d} /* (8, 20, 24) {real, imag} */,
  {32'h412273ce, 32'hc1364586} /* (8, 20, 23) {real, imag} */,
  {32'h42083634, 32'h418975fe} /* (8, 20, 22) {real, imag} */,
  {32'hc03eb0e0, 32'h4133ae44} /* (8, 20, 21) {real, imag} */,
  {32'hc08c4234, 32'h40d53659} /* (8, 20, 20) {real, imag} */,
  {32'h4112e3d2, 32'hc0e0ea48} /* (8, 20, 19) {real, imag} */,
  {32'h418bb020, 32'hc0493570} /* (8, 20, 18) {real, imag} */,
  {32'hc0eef50a, 32'h410fc261} /* (8, 20, 17) {real, imag} */,
  {32'hc132bd45, 32'h40b4c28c} /* (8, 20, 16) {real, imag} */,
  {32'h3f01ad10, 32'h414e77ab} /* (8, 20, 15) {real, imag} */,
  {32'h4052bd2c, 32'hc1625476} /* (8, 20, 14) {real, imag} */,
  {32'h40474bd1, 32'hc1191b84} /* (8, 20, 13) {real, imag} */,
  {32'h40d8c79c, 32'hbfae9db4} /* (8, 20, 12) {real, imag} */,
  {32'hc164e9fa, 32'hc18951ff} /* (8, 20, 11) {real, imag} */,
  {32'hc0e243cc, 32'hc0bf5bc2} /* (8, 20, 10) {real, imag} */,
  {32'hbefb2850, 32'hc19de2cf} /* (8, 20, 9) {real, imag} */,
  {32'h414b4310, 32'hc21f4efc} /* (8, 20, 8) {real, imag} */,
  {32'h413c603a, 32'hc1769f2c} /* (8, 20, 7) {real, imag} */,
  {32'hc1837b13, 32'h42172fb7} /* (8, 20, 6) {real, imag} */,
  {32'hc1b0b77d, 32'hc1e9cc4a} /* (8, 20, 5) {real, imag} */,
  {32'hc1ac41f7, 32'hc22c708e} /* (8, 20, 4) {real, imag} */,
  {32'hc1bf319a, 32'h42242599} /* (8, 20, 3) {real, imag} */,
  {32'hc1be29e2, 32'h41387901} /* (8, 20, 2) {real, imag} */,
  {32'h3f4960a0, 32'hc058d224} /* (8, 20, 1) {real, imag} */,
  {32'hc1a8f996, 32'hc2436a96} /* (8, 20, 0) {real, imag} */,
  {32'hc1c2280a, 32'h424bb5ee} /* (8, 19, 31) {real, imag} */,
  {32'h41a920d2, 32'h3e692980} /* (8, 19, 30) {real, imag} */,
  {32'h41486506, 32'hc1b5cce9} /* (8, 19, 29) {real, imag} */,
  {32'h41f63d7b, 32'h415ed370} /* (8, 19, 28) {real, imag} */,
  {32'hc098218c, 32'h4085d2b6} /* (8, 19, 27) {real, imag} */,
  {32'hc1bdbb63, 32'h40958edc} /* (8, 19, 26) {real, imag} */,
  {32'h41a9f47e, 32'h41972a23} /* (8, 19, 25) {real, imag} */,
  {32'h41cde4cf, 32'hc0a8d67e} /* (8, 19, 24) {real, imag} */,
  {32'h40666696, 32'hc1107077} /* (8, 19, 23) {real, imag} */,
  {32'h3ffe3de8, 32'h40f42928} /* (8, 19, 22) {real, imag} */,
  {32'h41dea603, 32'h4019658c} /* (8, 19, 21) {real, imag} */,
  {32'h419008b4, 32'h41a4a892} /* (8, 19, 20) {real, imag} */,
  {32'h40a28c19, 32'hc16b8db4} /* (8, 19, 19) {real, imag} */,
  {32'hc0b14610, 32'h408e1473} /* (8, 19, 18) {real, imag} */,
  {32'hbe488810, 32'h40da474b} /* (8, 19, 17) {real, imag} */,
  {32'h40591664, 32'h407ff618} /* (8, 19, 16) {real, imag} */,
  {32'h3de2d620, 32'h40582426} /* (8, 19, 15) {real, imag} */,
  {32'hc0c4855c, 32'hc10209e4} /* (8, 19, 14) {real, imag} */,
  {32'h41a060f3, 32'h40f5c8ab} /* (8, 19, 13) {real, imag} */,
  {32'hc188e292, 32'hbff40620} /* (8, 19, 12) {real, imag} */,
  {32'hc1520a26, 32'hbf9f7a91} /* (8, 19, 11) {real, imag} */,
  {32'hc167c457, 32'h40ab68b0} /* (8, 19, 10) {real, imag} */,
  {32'hc0d2f225, 32'h40d41cda} /* (8, 19, 9) {real, imag} */,
  {32'hc114fa66, 32'hc1d5229a} /* (8, 19, 8) {real, imag} */,
  {32'hbff180a0, 32'h418ac6b1} /* (8, 19, 7) {real, imag} */,
  {32'h4158028e, 32'hc21252e4} /* (8, 19, 6) {real, imag} */,
  {32'h42201622, 32'hc0b54548} /* (8, 19, 5) {real, imag} */,
  {32'h40a8c084, 32'h41cde036} /* (8, 19, 4) {real, imag} */,
  {32'h40c437cf, 32'hc1691a96} /* (8, 19, 3) {real, imag} */,
  {32'h41d4654a, 32'hc200040a} /* (8, 19, 2) {real, imag} */,
  {32'hc1b0b318, 32'hc218c34e} /* (8, 19, 1) {real, imag} */,
  {32'h42006c71, 32'hc13709a5} /* (8, 19, 0) {real, imag} */,
  {32'hc18ab8bb, 32'h411969e5} /* (8, 18, 31) {real, imag} */,
  {32'h4156a0a4, 32'h41bb9cbc} /* (8, 18, 30) {real, imag} */,
  {32'hc118e334, 32'h4258facb} /* (8, 18, 29) {real, imag} */,
  {32'h404cd6a8, 32'h417fab6e} /* (8, 18, 28) {real, imag} */,
  {32'hc103763a, 32'hc12202d5} /* (8, 18, 27) {real, imag} */,
  {32'hc18cf122, 32'hc0157761} /* (8, 18, 26) {real, imag} */,
  {32'h41543c22, 32'h41e477b4} /* (8, 18, 25) {real, imag} */,
  {32'h41853804, 32'hbe3d0a40} /* (8, 18, 24) {real, imag} */,
  {32'h415bb775, 32'hc1c1f97e} /* (8, 18, 23) {real, imag} */,
  {32'hc14bc3a5, 32'h411526b4} /* (8, 18, 22) {real, imag} */,
  {32'h40e064fe, 32'hc174dbdf} /* (8, 18, 21) {real, imag} */,
  {32'h4151514e, 32'hc193030b} /* (8, 18, 20) {real, imag} */,
  {32'hbf8375b5, 32'hc0aaffca} /* (8, 18, 19) {real, imag} */,
  {32'h4012d046, 32'hbe8469d0} /* (8, 18, 18) {real, imag} */,
  {32'h3f4d9d38, 32'h3f345e70} /* (8, 18, 17) {real, imag} */,
  {32'h40f6b66c, 32'hc090de70} /* (8, 18, 16) {real, imag} */,
  {32'hc0cddbbd, 32'h4059533c} /* (8, 18, 15) {real, imag} */,
  {32'hc006208a, 32'hc115df52} /* (8, 18, 14) {real, imag} */,
  {32'hc03b07fa, 32'h4080ad46} /* (8, 18, 13) {real, imag} */,
  {32'h40f3b505, 32'h40e9a5c3} /* (8, 18, 12) {real, imag} */,
  {32'hc0f1fc50, 32'hc19d0d40} /* (8, 18, 11) {real, imag} */,
  {32'hbe7e7840, 32'hbedd3eb0} /* (8, 18, 10) {real, imag} */,
  {32'h42109259, 32'h408a7f08} /* (8, 18, 9) {real, imag} */,
  {32'h41d43ebe, 32'h4080adc2} /* (8, 18, 8) {real, imag} */,
  {32'h4105939e, 32'h418bae30} /* (8, 18, 7) {real, imag} */,
  {32'hc21c6187, 32'hbf932e86} /* (8, 18, 6) {real, imag} */,
  {32'hc14bcd0e, 32'hc12bcad3} /* (8, 18, 5) {real, imag} */,
  {32'h4209d4fc, 32'h41130592} /* (8, 18, 4) {real, imag} */,
  {32'hc1809946, 32'hc0cc47b8} /* (8, 18, 3) {real, imag} */,
  {32'h41066044, 32'hc0672d20} /* (8, 18, 2) {real, imag} */,
  {32'hc155ace6, 32'hc219da77} /* (8, 18, 1) {real, imag} */,
  {32'hc2125064, 32'hc10c4b1a} /* (8, 18, 0) {real, imag} */,
  {32'hc175211d, 32'hc1356120} /* (8, 17, 31) {real, imag} */,
  {32'hc0ad943c, 32'hc0e179cc} /* (8, 17, 30) {real, imag} */,
  {32'h40cce620, 32'hc1002af0} /* (8, 17, 29) {real, imag} */,
  {32'h3fd6f9a8, 32'h401c5178} /* (8, 17, 28) {real, imag} */,
  {32'h40a64806, 32'h420f1c74} /* (8, 17, 27) {real, imag} */,
  {32'hc181dd1f, 32'h421a823a} /* (8, 17, 26) {real, imag} */,
  {32'hc06976d8, 32'hc12fd4f0} /* (8, 17, 25) {real, imag} */,
  {32'h4037c1f2, 32'h41e69b56} /* (8, 17, 24) {real, imag} */,
  {32'hc09c779a, 32'h41de68a6} /* (8, 17, 23) {real, imag} */,
  {32'h40b78f7e, 32'h416b5c2c} /* (8, 17, 22) {real, imag} */,
  {32'hbf892684, 32'h40dda896} /* (8, 17, 21) {real, imag} */,
  {32'hc15c9e12, 32'hc0532c5a} /* (8, 17, 20) {real, imag} */,
  {32'h3fd0c0d4, 32'hc10ad0b0} /* (8, 17, 19) {real, imag} */,
  {32'h4062714c, 32'h40665429} /* (8, 17, 18) {real, imag} */,
  {32'h3d8ba980, 32'hbfd9bca4} /* (8, 17, 17) {real, imag} */,
  {32'hc006e07c, 32'hc039e62b} /* (8, 17, 16) {real, imag} */,
  {32'hbdf05c80, 32'hc116f39c} /* (8, 17, 15) {real, imag} */,
  {32'h3e4cafc0, 32'h3e8ea698} /* (8, 17, 14) {real, imag} */,
  {32'h40c1d0f1, 32'hc0468f68} /* (8, 17, 13) {real, imag} */,
  {32'h4091c62c, 32'hc0ac3b25} /* (8, 17, 12) {real, imag} */,
  {32'hc12be95e, 32'h40d7b906} /* (8, 17, 11) {real, imag} */,
  {32'h40f09aae, 32'h418e7886} /* (8, 17, 10) {real, imag} */,
  {32'h3f11b3bc, 32'hbecc9d60} /* (8, 17, 9) {real, imag} */,
  {32'hc1121a02, 32'hc1b7f29a} /* (8, 17, 8) {real, imag} */,
  {32'h419dc977, 32'hc0960203} /* (8, 17, 7) {real, imag} */,
  {32'h40fdc078, 32'h4160e626} /* (8, 17, 6) {real, imag} */,
  {32'h41d3601e, 32'hc1382dbd} /* (8, 17, 5) {real, imag} */,
  {32'hc0f11418, 32'h41fbcd3f} /* (8, 17, 4) {real, imag} */,
  {32'hc2135806, 32'hc17abb4e} /* (8, 17, 3) {real, imag} */,
  {32'hc1521a5c, 32'hc03ea4c5} /* (8, 17, 2) {real, imag} */,
  {32'h4227ae1a, 32'h40766cd3} /* (8, 17, 1) {real, imag} */,
  {32'hc0657634, 32'h411ba82d} /* (8, 17, 0) {real, imag} */,
  {32'hc240205c, 32'hc10d2635} /* (8, 16, 31) {real, imag} */,
  {32'hc19cc32a, 32'hc153f86c} /* (8, 16, 30) {real, imag} */,
  {32'hc1dd8a4d, 32'h417330c2} /* (8, 16, 29) {real, imag} */,
  {32'hc1c2d565, 32'h3fcd6960} /* (8, 16, 28) {real, imag} */,
  {32'hc197168c, 32'hc1b92494} /* (8, 16, 27) {real, imag} */,
  {32'h41be5b06, 32'hbff556f8} /* (8, 16, 26) {real, imag} */,
  {32'h41502127, 32'h41bb28d6} /* (8, 16, 25) {real, imag} */,
  {32'hc0fbbdc4, 32'hc175f4bd} /* (8, 16, 24) {real, imag} */,
  {32'hc0805cac, 32'h40e39349} /* (8, 16, 23) {real, imag} */,
  {32'hc0928cdc, 32'h3fd6aff8} /* (8, 16, 22) {real, imag} */,
  {32'hc09e7bbd, 32'h41339f6a} /* (8, 16, 21) {real, imag} */,
  {32'h40256686, 32'hc1204904} /* (8, 16, 20) {real, imag} */,
  {32'hbf2c37a0, 32'h40ad6d3d} /* (8, 16, 19) {real, imag} */,
  {32'hc167915e, 32'h4022ce3b} /* (8, 16, 18) {real, imag} */,
  {32'h4092b1d8, 32'h3f871208} /* (8, 16, 17) {real, imag} */,
  {32'h4101c616, 32'h402bde80} /* (8, 16, 16) {real, imag} */,
  {32'hbe845280, 32'hc015b99a} /* (8, 16, 15) {real, imag} */,
  {32'hbfa38060, 32'hbffaf5ae} /* (8, 16, 14) {real, imag} */,
  {32'h408c2f40, 32'h405c08de} /* (8, 16, 13) {real, imag} */,
  {32'h3fb3b61d, 32'h40bb79d0} /* (8, 16, 12) {real, imag} */,
  {32'hc08c106d, 32'hbfae2a78} /* (8, 16, 11) {real, imag} */,
  {32'hc180e715, 32'h401ababc} /* (8, 16, 10) {real, imag} */,
  {32'hbf7beafc, 32'hc0d818df} /* (8, 16, 9) {real, imag} */,
  {32'h41cf76bf, 32'h4119627b} /* (8, 16, 8) {real, imag} */,
  {32'h410c0b27, 32'h40c6f97a} /* (8, 16, 7) {real, imag} */,
  {32'hc1af3914, 32'h41d53874} /* (8, 16, 6) {real, imag} */,
  {32'h41db203a, 32'h411a41b8} /* (8, 16, 5) {real, imag} */,
  {32'h41aeeac7, 32'h41dacb80} /* (8, 16, 4) {real, imag} */,
  {32'h42040668, 32'h41e3452f} /* (8, 16, 3) {real, imag} */,
  {32'h416bba63, 32'hc13c9bcc} /* (8, 16, 2) {real, imag} */,
  {32'hc12471c8, 32'h4097550a} /* (8, 16, 1) {real, imag} */,
  {32'hc10c24ea, 32'hc259fe04} /* (8, 16, 0) {real, imag} */,
  {32'h3f3394b4, 32'hc20b3d4c} /* (8, 15, 31) {real, imag} */,
  {32'h41021c84, 32'h420d57fe} /* (8, 15, 30) {real, imag} */,
  {32'h4177e15f, 32'hbf903068} /* (8, 15, 29) {real, imag} */,
  {32'h4132d9bc, 32'h41727728} /* (8, 15, 28) {real, imag} */,
  {32'hc18d2795, 32'hc1453d6e} /* (8, 15, 27) {real, imag} */,
  {32'hbf4d7d18, 32'h414637ec} /* (8, 15, 26) {real, imag} */,
  {32'hc178eece, 32'hc1a87026} /* (8, 15, 25) {real, imag} */,
  {32'h40a855cc, 32'hc119cc5e} /* (8, 15, 24) {real, imag} */,
  {32'h3fcc31c8, 32'hc171da6c} /* (8, 15, 23) {real, imag} */,
  {32'hc1711fc4, 32'hc1243a27} /* (8, 15, 22) {real, imag} */,
  {32'hc00495f7, 32'hc086c153} /* (8, 15, 21) {real, imag} */,
  {32'h400cf738, 32'h3f61a720} /* (8, 15, 20) {real, imag} */,
  {32'hc052448f, 32'h3f4a04d8} /* (8, 15, 19) {real, imag} */,
  {32'hbfa16456, 32'h401cb6b8} /* (8, 15, 18) {real, imag} */,
  {32'hc08f3ed3, 32'h3f8fd7bc} /* (8, 15, 17) {real, imag} */,
  {32'hc06a3228, 32'h3faf57d0} /* (8, 15, 16) {real, imag} */,
  {32'hbfae6070, 32'h409ad7e7} /* (8, 15, 15) {real, imag} */,
  {32'hbf2820bc, 32'hc07db138} /* (8, 15, 14) {real, imag} */,
  {32'h401c4169, 32'h40597c12} /* (8, 15, 13) {real, imag} */,
  {32'hc152f9d7, 32'hc16eb843} /* (8, 15, 12) {real, imag} */,
  {32'h3fed3bee, 32'h3fdff588} /* (8, 15, 11) {real, imag} */,
  {32'hc0038f1e, 32'hc0a0a550} /* (8, 15, 10) {real, imag} */,
  {32'hc08b396f, 32'hc0b28ff5} /* (8, 15, 9) {real, imag} */,
  {32'hc13daf6a, 32'h40518c86} /* (8, 15, 8) {real, imag} */,
  {32'hc043f600, 32'hc04bf93c} /* (8, 15, 7) {real, imag} */,
  {32'h414d84d6, 32'h41459d94} /* (8, 15, 6) {real, imag} */,
  {32'hc18dee47, 32'h40ced654} /* (8, 15, 5) {real, imag} */,
  {32'hc15c6804, 32'h41cd6c62} /* (8, 15, 4) {real, imag} */,
  {32'hc0d4d636, 32'hc1e17f58} /* (8, 15, 3) {real, imag} */,
  {32'h405a7f66, 32'h41f1b20d} /* (8, 15, 2) {real, imag} */,
  {32'hc055f7c7, 32'h41146eaa} /* (8, 15, 1) {real, imag} */,
  {32'h413d8438, 32'hc21842f6} /* (8, 15, 0) {real, imag} */,
  {32'h3fa79be0, 32'h41b37e89} /* (8, 14, 31) {real, imag} */,
  {32'hc1b99da9, 32'h418ecf38} /* (8, 14, 30) {real, imag} */,
  {32'hc0c58366, 32'hc210eb5c} /* (8, 14, 29) {real, imag} */,
  {32'hc1496cc2, 32'hc24d0d5c} /* (8, 14, 28) {real, imag} */,
  {32'h41f76f53, 32'hc0dddf1f} /* (8, 14, 27) {real, imag} */,
  {32'hc1dd6808, 32'h4173ff7c} /* (8, 14, 26) {real, imag} */,
  {32'h415a5e08, 32'h41d6e2b2} /* (8, 14, 25) {real, imag} */,
  {32'h40d73c75, 32'h4134c7d2} /* (8, 14, 24) {real, imag} */,
  {32'h41839055, 32'h40d8446b} /* (8, 14, 23) {real, imag} */,
  {32'hc17821d3, 32'hc11023d2} /* (8, 14, 22) {real, imag} */,
  {32'h40d39037, 32'h412adca0} /* (8, 14, 21) {real, imag} */,
  {32'hc110e09c, 32'h41478326} /* (8, 14, 20) {real, imag} */,
  {32'hbf0d9378, 32'hc039bdc0} /* (8, 14, 19) {real, imag} */,
  {32'h40ca09c1, 32'hc16421bf} /* (8, 14, 18) {real, imag} */,
  {32'hc0f4bfa0, 32'h4114eca1} /* (8, 14, 17) {real, imag} */,
  {32'hc093f579, 32'hc1286e2a} /* (8, 14, 16) {real, imag} */,
  {32'hc097c7f4, 32'hc0bc556a} /* (8, 14, 15) {real, imag} */,
  {32'h409b80fb, 32'h4111e92b} /* (8, 14, 14) {real, imag} */,
  {32'h404eb26c, 32'hbfd9fbe0} /* (8, 14, 13) {real, imag} */,
  {32'h3fd9541c, 32'h40909f24} /* (8, 14, 12) {real, imag} */,
  {32'h3f29b718, 32'h417d5fdc} /* (8, 14, 11) {real, imag} */,
  {32'h40f0aa2a, 32'h40f071e7} /* (8, 14, 10) {real, imag} */,
  {32'hc0da3414, 32'hc1a0f259} /* (8, 14, 9) {real, imag} */,
  {32'hc1846240, 32'hc1d054fd} /* (8, 14, 8) {real, imag} */,
  {32'h4145a374, 32'hc1748a1c} /* (8, 14, 7) {real, imag} */,
  {32'hc07b7e04, 32'hc1f99b42} /* (8, 14, 6) {real, imag} */,
  {32'hbfc27310, 32'h41093ae4} /* (8, 14, 5) {real, imag} */,
  {32'h41d2c031, 32'h41477fea} /* (8, 14, 4) {real, imag} */,
  {32'hc061955d, 32'h410a0f84} /* (8, 14, 3) {real, imag} */,
  {32'hc0feb759, 32'hbfe07268} /* (8, 14, 2) {real, imag} */,
  {32'h41f3128d, 32'h41c4ee75} /* (8, 14, 1) {real, imag} */,
  {32'h41a308de, 32'h41582664} /* (8, 14, 0) {real, imag} */,
  {32'hc1d83a5a, 32'h4215055d} /* (8, 13, 31) {real, imag} */,
  {32'hc12e494e, 32'hc21750f6} /* (8, 13, 30) {real, imag} */,
  {32'h41d59035, 32'h41c557cc} /* (8, 13, 29) {real, imag} */,
  {32'h41af21ab, 32'h41854a5f} /* (8, 13, 28) {real, imag} */,
  {32'h4180902c, 32'h3fca81e0} /* (8, 13, 27) {real, imag} */,
  {32'h3e6c3e00, 32'h41839141} /* (8, 13, 26) {real, imag} */,
  {32'hc11edd2a, 32'h41d0e1c7} /* (8, 13, 25) {real, imag} */,
  {32'hc1b19cb6, 32'h407bed86} /* (8, 13, 24) {real, imag} */,
  {32'hc1b03ff9, 32'h41e5d0cc} /* (8, 13, 23) {real, imag} */,
  {32'hc093f70c, 32'hc169bcb0} /* (8, 13, 22) {real, imag} */,
  {32'h40d5362c, 32'hc19f7e34} /* (8, 13, 21) {real, imag} */,
  {32'h40e83df6, 32'hc1273106} /* (8, 13, 20) {real, imag} */,
  {32'hc0aa939e, 32'h414cdc7a} /* (8, 13, 19) {real, imag} */,
  {32'h4155e340, 32'hc00605c0} /* (8, 13, 18) {real, imag} */,
  {32'h41040869, 32'h3fc64790} /* (8, 13, 17) {real, imag} */,
  {32'hc11f0618, 32'h40b59704} /* (8, 13, 16) {real, imag} */,
  {32'h4002edef, 32'hc0f45a78} /* (8, 13, 15) {real, imag} */,
  {32'h3eba3eb0, 32'hc1027b3e} /* (8, 13, 14) {real, imag} */,
  {32'h3f418990, 32'hbfa5bcfc} /* (8, 13, 13) {real, imag} */,
  {32'h41453827, 32'hbf14c420} /* (8, 13, 12) {real, imag} */,
  {32'hc1d9fd8b, 32'hc1a1f9cc} /* (8, 13, 11) {real, imag} */,
  {32'h41275956, 32'hc0532b12} /* (8, 13, 10) {real, imag} */,
  {32'h41c8e5ff, 32'h40b14246} /* (8, 13, 9) {real, imag} */,
  {32'h41f7882c, 32'hc1117be8} /* (8, 13, 8) {real, imag} */,
  {32'h40a6aa29, 32'hc133ffc6} /* (8, 13, 7) {real, imag} */,
  {32'h4151b8f8, 32'h41c5a717} /* (8, 13, 6) {real, imag} */,
  {32'h4113554c, 32'h420b3c7b} /* (8, 13, 5) {real, imag} */,
  {32'hc086df60, 32'hc22a4926} /* (8, 13, 4) {real, imag} */,
  {32'hc1b079cb, 32'h41442bad} /* (8, 13, 3) {real, imag} */,
  {32'h3fda86c4, 32'hc1ba8134} /* (8, 13, 2) {real, imag} */,
  {32'hc162e619, 32'h42010d49} /* (8, 13, 1) {real, imag} */,
  {32'h3fbc0a20, 32'hc2224e86} /* (8, 13, 0) {real, imag} */,
  {32'hc14843c0, 32'h421a4967} /* (8, 12, 31) {real, imag} */,
  {32'hbcb99200, 32'hc23970a7} /* (8, 12, 30) {real, imag} */,
  {32'hc233bc92, 32'h41c22a4b} /* (8, 12, 29) {real, imag} */,
  {32'hc02f7040, 32'hc271c85c} /* (8, 12, 28) {real, imag} */,
  {32'h40c50e02, 32'hc1e9018c} /* (8, 12, 27) {real, imag} */,
  {32'hc1d7f7e4, 32'h419e31f4} /* (8, 12, 26) {real, imag} */,
  {32'hbe9a3f80, 32'hc125b840} /* (8, 12, 25) {real, imag} */,
  {32'h41e45c8a, 32'hc11ad8bc} /* (8, 12, 24) {real, imag} */,
  {32'hc151ea42, 32'hc0af584c} /* (8, 12, 23) {real, imag} */,
  {32'h413f6296, 32'hc19c8c09} /* (8, 12, 22) {real, imag} */,
  {32'hc16031f6, 32'hc1a9996b} /* (8, 12, 21) {real, imag} */,
  {32'hc063b189, 32'hc114f922} /* (8, 12, 20) {real, imag} */,
  {32'h417c1b13, 32'hc05e9780} /* (8, 12, 19) {real, imag} */,
  {32'hc1798f57, 32'hc10e90b8} /* (8, 12, 18) {real, imag} */,
  {32'h4101374a, 32'h40406880} /* (8, 12, 17) {real, imag} */,
  {32'h40edc20c, 32'h411b84b1} /* (8, 12, 16) {real, imag} */,
  {32'h3eff6ae0, 32'hc1cfdb9d} /* (8, 12, 15) {real, imag} */,
  {32'hc10a3fbf, 32'hc00d0968} /* (8, 12, 14) {real, imag} */,
  {32'hc0ce7142, 32'hc1447b40} /* (8, 12, 13) {real, imag} */,
  {32'h40824c0c, 32'h3f58ff60} /* (8, 12, 12) {real, imag} */,
  {32'hc0158832, 32'h413e71ca} /* (8, 12, 11) {real, imag} */,
  {32'hc1df7235, 32'h3fa37cc0} /* (8, 12, 10) {real, imag} */,
  {32'h40cfd2bf, 32'hc116b8b6} /* (8, 12, 9) {real, imag} */,
  {32'h40a22de8, 32'h42619ecd} /* (8, 12, 8) {real, imag} */,
  {32'h4216fa63, 32'h42312785} /* (8, 12, 7) {real, imag} */,
  {32'h40ca51b0, 32'hc18a8d50} /* (8, 12, 6) {real, imag} */,
  {32'h41cb7d0e, 32'hc20ff9a2} /* (8, 12, 5) {real, imag} */,
  {32'hc18a7f14, 32'h41d2f634} /* (8, 12, 4) {real, imag} */,
  {32'h3f241e60, 32'hc1ee5a05} /* (8, 12, 3) {real, imag} */,
  {32'hc1402fa5, 32'hc09a1ef8} /* (8, 12, 2) {real, imag} */,
  {32'hc1921fea, 32'hc0c421f8} /* (8, 12, 1) {real, imag} */,
  {32'hc099af14, 32'h41b00fc2} /* (8, 12, 0) {real, imag} */,
  {32'h429d84ea, 32'h420f4b96} /* (8, 11, 31) {real, imag} */,
  {32'h41880a27, 32'h41635e0c} /* (8, 11, 30) {real, imag} */,
  {32'h3eaf0cc0, 32'h418fc4f0} /* (8, 11, 29) {real, imag} */,
  {32'h4164fb11, 32'hc262c010} /* (8, 11, 28) {real, imag} */,
  {32'hc155e544, 32'hc24917fa} /* (8, 11, 27) {real, imag} */,
  {32'h41fa886b, 32'h41579606} /* (8, 11, 26) {real, imag} */,
  {32'hc1b328c5, 32'hc1991faa} /* (8, 11, 25) {real, imag} */,
  {32'h4012716c, 32'h41c6dfb7} /* (8, 11, 24) {real, imag} */,
  {32'hc0886ff4, 32'hc1716185} /* (8, 11, 23) {real, imag} */,
  {32'h418960eb, 32'h412231a2} /* (8, 11, 22) {real, imag} */,
  {32'hc025a0ce, 32'h414687b2} /* (8, 11, 21) {real, imag} */,
  {32'h404b911c, 32'h4187fb37} /* (8, 11, 20) {real, imag} */,
  {32'h40cee79c, 32'hc0b1d0ba} /* (8, 11, 19) {real, imag} */,
  {32'hc0864485, 32'h40ae282c} /* (8, 11, 18) {real, imag} */,
  {32'hc1239268, 32'h3fd372f8} /* (8, 11, 17) {real, imag} */,
  {32'h40341658, 32'h4079f678} /* (8, 11, 16) {real, imag} */,
  {32'h3f6c92c0, 32'h411c6d25} /* (8, 11, 15) {real, imag} */,
  {32'h409878db, 32'hc1a6fd97} /* (8, 11, 14) {real, imag} */,
  {32'hc19d83a1, 32'hc1316945} /* (8, 11, 13) {real, imag} */,
  {32'hc16ddf97, 32'hbf53f920} /* (8, 11, 12) {real, imag} */,
  {32'hc0cdff41, 32'h41c2d84b} /* (8, 11, 11) {real, imag} */,
  {32'hc21175c0, 32'h41cc521b} /* (8, 11, 10) {real, imag} */,
  {32'h419e3051, 32'hc1821352} /* (8, 11, 9) {real, imag} */,
  {32'hc1db142e, 32'hc1d0fafd} /* (8, 11, 8) {real, imag} */,
  {32'hc21d48c2, 32'h41a6cf54} /* (8, 11, 7) {real, imag} */,
  {32'h42020966, 32'hc1168eae} /* (8, 11, 6) {real, imag} */,
  {32'hc1f931a4, 32'h4137917a} /* (8, 11, 5) {real, imag} */,
  {32'h42063513, 32'hc1efebdf} /* (8, 11, 4) {real, imag} */,
  {32'h41bd987f, 32'hc22fa454} /* (8, 11, 3) {real, imag} */,
  {32'hc22713f8, 32'hc281d91e} /* (8, 11, 2) {real, imag} */,
  {32'h418703ff, 32'h41a1334a} /* (8, 11, 1) {real, imag} */,
  {32'h420471a4, 32'h426fcce2} /* (8, 11, 0) {real, imag} */,
  {32'hc27c76e2, 32'hc296ae3c} /* (8, 10, 31) {real, imag} */,
  {32'h40ba3b70, 32'h4229394e} /* (8, 10, 30) {real, imag} */,
  {32'h40e86664, 32'h40c110b4} /* (8, 10, 29) {real, imag} */,
  {32'hc1bbdc9d, 32'h41c3926c} /* (8, 10, 28) {real, imag} */,
  {32'h40899600, 32'hc1da3243} /* (8, 10, 27) {real, imag} */,
  {32'hc0877956, 32'h3f8ce5e0} /* (8, 10, 26) {real, imag} */,
  {32'hbf3e5950, 32'hc0671080} /* (8, 10, 25) {real, imag} */,
  {32'h4162b68c, 32'hc0b19a08} /* (8, 10, 24) {real, imag} */,
  {32'hc1dca146, 32'hc17a51de} /* (8, 10, 23) {real, imag} */,
  {32'h40714bf4, 32'hc0a9de56} /* (8, 10, 22) {real, imag} */,
  {32'h418b5ca8, 32'hc05a751c} /* (8, 10, 21) {real, imag} */,
  {32'hc0982cd4, 32'h4065fc7f} /* (8, 10, 20) {real, imag} */,
  {32'h41884b38, 32'h417f6ec4} /* (8, 10, 19) {real, imag} */,
  {32'h3f864080, 32'hc0c6701e} /* (8, 10, 18) {real, imag} */,
  {32'h40bf94b4, 32'hc0f39835} /* (8, 10, 17) {real, imag} */,
  {32'hbffc9b60, 32'hc02accf9} /* (8, 10, 16) {real, imag} */,
  {32'h413e805e, 32'hc0e54d9d} /* (8, 10, 15) {real, imag} */,
  {32'hc150f670, 32'h401ae49c} /* (8, 10, 14) {real, imag} */,
  {32'h3f8f9528, 32'h41a620e8} /* (8, 10, 13) {real, imag} */,
  {32'hc1543bca, 32'h3fb2a32e} /* (8, 10, 12) {real, imag} */,
  {32'h413a8d64, 32'hc0042ac4} /* (8, 10, 11) {real, imag} */,
  {32'h42070832, 32'hc1812024} /* (8, 10, 10) {real, imag} */,
  {32'h418e60d4, 32'h40375aba} /* (8, 10, 9) {real, imag} */,
  {32'hc1d5cddc, 32'h41328a00} /* (8, 10, 8) {real, imag} */,
  {32'hbf67f090, 32'hc1fbef28} /* (8, 10, 7) {real, imag} */,
  {32'hc1e232d8, 32'hc2133d87} /* (8, 10, 6) {real, imag} */,
  {32'h41585a60, 32'h40843a28} /* (8, 10, 5) {real, imag} */,
  {32'hc0e709d4, 32'hc07f4c74} /* (8, 10, 4) {real, imag} */,
  {32'hc25dba6a, 32'hc128c09e} /* (8, 10, 3) {real, imag} */,
  {32'h428d31e5, 32'hbeb72640} /* (8, 10, 2) {real, imag} */,
  {32'hc1aaa4cf, 32'h421718a4} /* (8, 10, 1) {real, imag} */,
  {32'hc22c02fe, 32'h3fe51cae} /* (8, 10, 0) {real, imag} */,
  {32'hc26f0cf7, 32'hc24c1c16} /* (8, 9, 31) {real, imag} */,
  {32'hc1256978, 32'hc29f1ed6} /* (8, 9, 30) {real, imag} */,
  {32'h41836ff4, 32'hc1f6c203} /* (8, 9, 29) {real, imag} */,
  {32'hc279e7af, 32'hc20475f8} /* (8, 9, 28) {real, imag} */,
  {32'h419ab56f, 32'h41f32cec} /* (8, 9, 27) {real, imag} */,
  {32'h417bcace, 32'h4245f398} /* (8, 9, 26) {real, imag} */,
  {32'h4148d430, 32'hc08c0b4f} /* (8, 9, 25) {real, imag} */,
  {32'hc0c19d2c, 32'h41d1a810} /* (8, 9, 24) {real, imag} */,
  {32'h41995e5b, 32'hc21a2e93} /* (8, 9, 23) {real, imag} */,
  {32'h409da6b4, 32'h40c719a4} /* (8, 9, 22) {real, imag} */,
  {32'hc193ca10, 32'hc12946f7} /* (8, 9, 21) {real, imag} */,
  {32'h411a7718, 32'h40c31374} /* (8, 9, 20) {real, imag} */,
  {32'h41bc2054, 32'h4215ddb2} /* (8, 9, 19) {real, imag} */,
  {32'hc196478f, 32'hbf9417b0} /* (8, 9, 18) {real, imag} */,
  {32'h41a2ab2a, 32'h40563c84} /* (8, 9, 17) {real, imag} */,
  {32'hc07bad50, 32'hc122a102} /* (8, 9, 16) {real, imag} */,
  {32'h4183c82e, 32'h41944432} /* (8, 9, 15) {real, imag} */,
  {32'h3e49b380, 32'hc09f9914} /* (8, 9, 14) {real, imag} */,
  {32'h41fdd08c, 32'hc00bfd38} /* (8, 9, 13) {real, imag} */,
  {32'h420410f1, 32'h419feadf} /* (8, 9, 12) {real, imag} */,
  {32'hc0a373a0, 32'hc1664917} /* (8, 9, 11) {real, imag} */,
  {32'h410ef536, 32'h41d20ff9} /* (8, 9, 10) {real, imag} */,
  {32'hc21fb036, 32'h41e62902} /* (8, 9, 9) {real, imag} */,
  {32'h418af769, 32'hc18da96e} /* (8, 9, 8) {real, imag} */,
  {32'hc084e101, 32'h4088aef9} /* (8, 9, 7) {real, imag} */,
  {32'hc1cf5313, 32'h4128f4f2} /* (8, 9, 6) {real, imag} */,
  {32'hc1823921, 32'hc189184e} /* (8, 9, 5) {real, imag} */,
  {32'hc21e7769, 32'h426a0318} /* (8, 9, 4) {real, imag} */,
  {32'h42802a0b, 32'hc2ac41ea} /* (8, 9, 3) {real, imag} */,
  {32'hc0f24de1, 32'h41146df4} /* (8, 9, 2) {real, imag} */,
  {32'hc214c43d, 32'hc08ea624} /* (8, 9, 1) {real, imag} */,
  {32'hc26bee84, 32'hc2084316} /* (8, 9, 0) {real, imag} */,
  {32'h429e88be, 32'hc1c8c846} /* (8, 8, 31) {real, imag} */,
  {32'h41f19fc4, 32'h423e492f} /* (8, 8, 30) {real, imag} */,
  {32'h4247e383, 32'hc2a5dad2} /* (8, 8, 29) {real, imag} */,
  {32'h42b7142b, 32'hc2a9aeb0} /* (8, 8, 28) {real, imag} */,
  {32'hc1add5de, 32'hc1839993} /* (8, 8, 27) {real, imag} */,
  {32'hc1b0eac9, 32'hc2527212} /* (8, 8, 26) {real, imag} */,
  {32'h3e586100, 32'hc2a30582} /* (8, 8, 25) {real, imag} */,
  {32'hc2085151, 32'hc1d6785c} /* (8, 8, 24) {real, imag} */,
  {32'hc1659144, 32'hc2477157} /* (8, 8, 23) {real, imag} */,
  {32'hc0a1585c, 32'h4265d3ca} /* (8, 8, 22) {real, imag} */,
  {32'h41e62d29, 32'h41f4a4db} /* (8, 8, 21) {real, imag} */,
  {32'hc147606e, 32'h40fa9cf2} /* (8, 8, 20) {real, imag} */,
  {32'hc0b2e290, 32'hc13863ee} /* (8, 8, 19) {real, imag} */,
  {32'h4108df88, 32'h40160a00} /* (8, 8, 18) {real, imag} */,
  {32'hc10fdf7e, 32'h3f8de700} /* (8, 8, 17) {real, imag} */,
  {32'h4173fc7c, 32'hc2088aca} /* (8, 8, 16) {real, imag} */,
  {32'h419e967b, 32'hbffc8080} /* (8, 8, 15) {real, imag} */,
  {32'hc1faa60c, 32'h42377312} /* (8, 8, 14) {real, imag} */,
  {32'hc15c4704, 32'hc09b75dc} /* (8, 8, 13) {real, imag} */,
  {32'h409777fc, 32'h4051ef9c} /* (8, 8, 12) {real, imag} */,
  {32'hc24d66f4, 32'hc0239e38} /* (8, 8, 11) {real, imag} */,
  {32'h42325bf2, 32'h422ef87a} /* (8, 8, 10) {real, imag} */,
  {32'h4294239a, 32'hc23de149} /* (8, 8, 9) {real, imag} */,
  {32'hc1a40a50, 32'hc24e9d0a} /* (8, 8, 8) {real, imag} */,
  {32'hc238652b, 32'h413db594} /* (8, 8, 7) {real, imag} */,
  {32'h421ff534, 32'hc2085d2a} /* (8, 8, 6) {real, imag} */,
  {32'h41fe6b80, 32'hc2046440} /* (8, 8, 5) {real, imag} */,
  {32'h42909f43, 32'hc311f9ca} /* (8, 8, 4) {real, imag} */,
  {32'hc0de06d0, 32'hc222d355} /* (8, 8, 3) {real, imag} */,
  {32'hc34cca1c, 32'h40ecca48} /* (8, 8, 2) {real, imag} */,
  {32'h41d0da43, 32'h420d6531} /* (8, 8, 1) {real, imag} */,
  {32'h426f2b45, 32'h4167523f} /* (8, 8, 0) {real, imag} */,
  {32'hc2e0d0ac, 32'hc23a4477} /* (8, 7, 31) {real, imag} */,
  {32'hc0cd717e, 32'hc1abf0a2} /* (8, 7, 30) {real, imag} */,
  {32'hc290b20f, 32'hc17d7c28} /* (8, 7, 29) {real, imag} */,
  {32'h41c22aac, 32'h4150d1b6} /* (8, 7, 28) {real, imag} */,
  {32'hc20cb2c1, 32'hc088a1f8} /* (8, 7, 27) {real, imag} */,
  {32'h41eb30e8, 32'hc2402643} /* (8, 7, 26) {real, imag} */,
  {32'h3fadb390, 32'h427a5ed4} /* (8, 7, 25) {real, imag} */,
  {32'hc1a990c0, 32'hc186e93c} /* (8, 7, 24) {real, imag} */,
  {32'hc10a1d6d, 32'hc0b3f560} /* (8, 7, 23) {real, imag} */,
  {32'h422f10c6, 32'hc13b7e06} /* (8, 7, 22) {real, imag} */,
  {32'hc2166b53, 32'h41f5dd58} /* (8, 7, 21) {real, imag} */,
  {32'h40fc1854, 32'hbf55b5e0} /* (8, 7, 20) {real, imag} */,
  {32'h402defc8, 32'h3dcbe500} /* (8, 7, 19) {real, imag} */,
  {32'h3ffb0c60, 32'hc1c31e02} /* (8, 7, 18) {real, imag} */,
  {32'h4113d6dc, 32'h419c1352} /* (8, 7, 17) {real, imag} */,
  {32'h40afa420, 32'h40a2dd88} /* (8, 7, 16) {real, imag} */,
  {32'hc028efd0, 32'hc0b98fa8} /* (8, 7, 15) {real, imag} */,
  {32'h41dea41e, 32'h418b848a} /* (8, 7, 14) {real, imag} */,
  {32'hc1ee42fd, 32'hc189774d} /* (8, 7, 13) {real, imag} */,
  {32'hc0bce188, 32'h40da6c8c} /* (8, 7, 12) {real, imag} */,
  {32'h424a3e95, 32'hc0efc252} /* (8, 7, 11) {real, imag} */,
  {32'h401ffe08, 32'h40d838fd} /* (8, 7, 10) {real, imag} */,
  {32'h41a1d4ec, 32'hc200bb78} /* (8, 7, 9) {real, imag} */,
  {32'h410c9297, 32'h42b7d7cf} /* (8, 7, 8) {real, imag} */,
  {32'hc2146562, 32'h42282370} /* (8, 7, 7) {real, imag} */,
  {32'hc24ef330, 32'h41597440} /* (8, 7, 6) {real, imag} */,
  {32'h42834172, 32'h4267f041} /* (8, 7, 5) {real, imag} */,
  {32'hc1c53914, 32'h426ac514} /* (8, 7, 4) {real, imag} */,
  {32'hc2bc07ad, 32'h42a0b01d} /* (8, 7, 3) {real, imag} */,
  {32'h3f003d80, 32'hc0b5d82a} /* (8, 7, 2) {real, imag} */,
  {32'h4232d6e3, 32'hc32115f5} /* (8, 7, 1) {real, imag} */,
  {32'h423ead20, 32'h42b1346e} /* (8, 7, 0) {real, imag} */,
  {32'h430454e9, 32'hc21d5d33} /* (8, 6, 31) {real, imag} */,
  {32'h42a7c062, 32'h4286cc9a} /* (8, 6, 30) {real, imag} */,
  {32'h42c46c78, 32'hc2b232b6} /* (8, 6, 29) {real, imag} */,
  {32'hc26a1e48, 32'h423f4ef0} /* (8, 6, 28) {real, imag} */,
  {32'hc25a0c09, 32'h4252e16e} /* (8, 6, 27) {real, imag} */,
  {32'hc1ecb41c, 32'hc2912e6c} /* (8, 6, 26) {real, imag} */,
  {32'h42b29774, 32'h41ffab29} /* (8, 6, 25) {real, imag} */,
  {32'h411f2506, 32'hc1da051a} /* (8, 6, 24) {real, imag} */,
  {32'h41967af4, 32'h41aa04aa} /* (8, 6, 23) {real, imag} */,
  {32'h418e9949, 32'h4198be8e} /* (8, 6, 22) {real, imag} */,
  {32'hc1319235, 32'hc0357ac8} /* (8, 6, 21) {real, imag} */,
  {32'h40aefd9c, 32'hc208796e} /* (8, 6, 20) {real, imag} */,
  {32'hc15aad03, 32'hc1504dd4} /* (8, 6, 19) {real, imag} */,
  {32'h4070ce9c, 32'hc1dc05a4} /* (8, 6, 18) {real, imag} */,
  {32'h4245dc67, 32'h419a6a68} /* (8, 6, 17) {real, imag} */,
  {32'hc162fe1b, 32'hc135b414} /* (8, 6, 16) {real, imag} */,
  {32'h40ec0508, 32'hc023d580} /* (8, 6, 15) {real, imag} */,
  {32'h404f2e84, 32'h3fefffb8} /* (8, 6, 14) {real, imag} */,
  {32'hc111f26b, 32'hc1b1e7c6} /* (8, 6, 13) {real, imag} */,
  {32'h41f04c91, 32'hc1a66fa6} /* (8, 6, 12) {real, imag} */,
  {32'h40a70466, 32'h41eb94e7} /* (8, 6, 11) {real, imag} */,
  {32'hc1e86803, 32'h412af14c} /* (8, 6, 10) {real, imag} */,
  {32'h40db210e, 32'hc2aaf63a} /* (8, 6, 9) {real, imag} */,
  {32'hc24e4518, 32'hc2a69b9a} /* (8, 6, 8) {real, imag} */,
  {32'hc26d95d8, 32'h422657a6} /* (8, 6, 7) {real, imag} */,
  {32'hc2449e06, 32'hc1aa8e3e} /* (8, 6, 6) {real, imag} */,
  {32'h4223f851, 32'hc216182e} /* (8, 6, 5) {real, imag} */,
  {32'h40554fe8, 32'hc15b733a} /* (8, 6, 4) {real, imag} */,
  {32'hc23e4158, 32'h42aea4d6} /* (8, 6, 3) {real, imag} */,
  {32'h41b80334, 32'hc18e5b32} /* (8, 6, 2) {real, imag} */,
  {32'h428f939a, 32'h4182bf92} /* (8, 6, 1) {real, imag} */,
  {32'hc13c72d9, 32'hc2997dd2} /* (8, 6, 0) {real, imag} */,
  {32'h42ee5e3b, 32'hc3390852} /* (8, 5, 31) {real, imag} */,
  {32'hc2bf1f12, 32'h4287b3e3} /* (8, 5, 30) {real, imag} */,
  {32'h41c046a9, 32'hc168c066} /* (8, 5, 29) {real, imag} */,
  {32'h42bcf31e, 32'h40bbb398} /* (8, 5, 28) {real, imag} */,
  {32'h421526bc, 32'h426bd36a} /* (8, 5, 27) {real, imag} */,
  {32'h421a3f53, 32'hc06a7894} /* (8, 5, 26) {real, imag} */,
  {32'h423c137c, 32'hc21bb7a4} /* (8, 5, 25) {real, imag} */,
  {32'h4208b99a, 32'hc1b97843} /* (8, 5, 24) {real, imag} */,
  {32'h41b45bac, 32'hbfd39b32} /* (8, 5, 23) {real, imag} */,
  {32'hc0b23544, 32'h4275521a} /* (8, 5, 22) {real, imag} */,
  {32'hc1b6bef6, 32'hc0a00c8a} /* (8, 5, 21) {real, imag} */,
  {32'hc15c88c3, 32'h414d045a} /* (8, 5, 20) {real, imag} */,
  {32'hc1555828, 32'h419a7fb0} /* (8, 5, 19) {real, imag} */,
  {32'h4140f5b8, 32'h414e38fa} /* (8, 5, 18) {real, imag} */,
  {32'hc1062daa, 32'hbfd6e380} /* (8, 5, 17) {real, imag} */,
  {32'h40fdcf70, 32'h414f4100} /* (8, 5, 16) {real, imag} */,
  {32'h4209ac5e, 32'h416189e0} /* (8, 5, 15) {real, imag} */,
  {32'hc13ae7e8, 32'hc21ba846} /* (8, 5, 14) {real, imag} */,
  {32'hc1b792a6, 32'hc21cb29f} /* (8, 5, 13) {real, imag} */,
  {32'h418239d2, 32'h40bee264} /* (8, 5, 12) {real, imag} */,
  {32'h426c5d1d, 32'hc2075eab} /* (8, 5, 11) {real, imag} */,
  {32'h41305d72, 32'hc19a795c} /* (8, 5, 10) {real, imag} */,
  {32'hc209780a, 32'h402b6217} /* (8, 5, 9) {real, imag} */,
  {32'hc1d4f721, 32'h41149f8a} /* (8, 5, 8) {real, imag} */,
  {32'h40fce990, 32'h420fd000} /* (8, 5, 7) {real, imag} */,
  {32'hc234e071, 32'h3ec280e0} /* (8, 5, 6) {real, imag} */,
  {32'h42be695a, 32'h42914fbd} /* (8, 5, 5) {real, imag} */,
  {32'h427fb484, 32'h42fdc3ea} /* (8, 5, 4) {real, imag} */,
  {32'h4261348c, 32'hc25c8906} /* (8, 5, 3) {real, imag} */,
  {32'hc28e355c, 32'hc28335f3} /* (8, 5, 2) {real, imag} */,
  {32'h429ff62f, 32'h4223f96a} /* (8, 5, 1) {real, imag} */,
  {32'h432e1eac, 32'hc2a147a2} /* (8, 5, 0) {real, imag} */,
  {32'hc2bcbd9f, 32'hc2b806ce} /* (8, 4, 31) {real, imag} */,
  {32'h4347cff7, 32'hc167bea4} /* (8, 4, 30) {real, imag} */,
  {32'h427994fb, 32'hc242dfcb} /* (8, 4, 29) {real, imag} */,
  {32'hc19bd3e8, 32'h41ed35d0} /* (8, 4, 28) {real, imag} */,
  {32'h41a24a4e, 32'hc02e3ada} /* (8, 4, 27) {real, imag} */,
  {32'hc22a9146, 32'hc29d1a73} /* (8, 4, 26) {real, imag} */,
  {32'h42a315c7, 32'hc2077653} /* (8, 4, 25) {real, imag} */,
  {32'h4231d532, 32'hc09d84c8} /* (8, 4, 24) {real, imag} */,
  {32'hc2159e20, 32'hc1a098b0} /* (8, 4, 23) {real, imag} */,
  {32'h40fa7cdc, 32'hc0f2d930} /* (8, 4, 22) {real, imag} */,
  {32'h422d980d, 32'h4161765e} /* (8, 4, 21) {real, imag} */,
  {32'hc16f0afd, 32'h3fd80d40} /* (8, 4, 20) {real, imag} */,
  {32'h41ac3504, 32'hc02bab88} /* (8, 4, 19) {real, imag} */,
  {32'h42242e99, 32'h41a9ff2e} /* (8, 4, 18) {real, imag} */,
  {32'hc14007a0, 32'h41c7bf45} /* (8, 4, 17) {real, imag} */,
  {32'h41fc2685, 32'hc13b59b6} /* (8, 4, 16) {real, imag} */,
  {32'hc0037800, 32'hc1720e66} /* (8, 4, 15) {real, imag} */,
  {32'hc1abead2, 32'h41a06d7a} /* (8, 4, 14) {real, imag} */,
  {32'hc246ccce, 32'h422317ea} /* (8, 4, 13) {real, imag} */,
  {32'h4064a024, 32'h421026d2} /* (8, 4, 12) {real, imag} */,
  {32'hc192852e, 32'hc22cb05c} /* (8, 4, 11) {real, imag} */,
  {32'h40ba8f9c, 32'hc2738494} /* (8, 4, 10) {real, imag} */,
  {32'hc26e023c, 32'h421b456d} /* (8, 4, 9) {real, imag} */,
  {32'h429a4c05, 32'hc2f6bff0} /* (8, 4, 8) {real, imag} */,
  {32'hc313c194, 32'h41a04418} /* (8, 4, 7) {real, imag} */,
  {32'h425920ba, 32'hc2bf7271} /* (8, 4, 6) {real, imag} */,
  {32'h42299cff, 32'h404cdf3e} /* (8, 4, 5) {real, imag} */,
  {32'hc27347f0, 32'hc33785ca} /* (8, 4, 4) {real, imag} */,
  {32'h41ebffde, 32'h425ebeab} /* (8, 4, 3) {real, imag} */,
  {32'h434b5179, 32'hc28137a6} /* (8, 4, 2) {real, imag} */,
  {32'hc357030a, 32'h42c03634} /* (8, 4, 1) {real, imag} */,
  {32'hc1b477cf, 32'hc19436ed} /* (8, 4, 0) {real, imag} */,
  {32'hc2883d50, 32'hc3227250} /* (8, 3, 31) {real, imag} */,
  {32'h4268dcd8, 32'h427af75e} /* (8, 3, 30) {real, imag} */,
  {32'h4301d463, 32'hc0c0294e} /* (8, 3, 29) {real, imag} */,
  {32'hc2ec0b64, 32'h423c5698} /* (8, 3, 28) {real, imag} */,
  {32'hc1eebb00, 32'hc1c1fdc7} /* (8, 3, 27) {real, imag} */,
  {32'hc21af31e, 32'h4291e48f} /* (8, 3, 26) {real, imag} */,
  {32'hc1f763fc, 32'h4235d019} /* (8, 3, 25) {real, imag} */,
  {32'hc1facf7a, 32'hc2ccd6ee} /* (8, 3, 24) {real, imag} */,
  {32'hc04da3a0, 32'h40f27100} /* (8, 3, 23) {real, imag} */,
  {32'h429abe98, 32'h41b17968} /* (8, 3, 22) {real, imag} */,
  {32'h420abe06, 32'h42017ebc} /* (8, 3, 21) {real, imag} */,
  {32'h4233fb08, 32'hc1c42d83} /* (8, 3, 20) {real, imag} */,
  {32'hc23ec5d6, 32'hc202b6a5} /* (8, 3, 19) {real, imag} */,
  {32'h3fb413d0, 32'h4224eec6} /* (8, 3, 18) {real, imag} */,
  {32'hc21ccd00, 32'hc114ad9a} /* (8, 3, 17) {real, imag} */,
  {32'h411d05ac, 32'h4217e272} /* (8, 3, 16) {real, imag} */,
  {32'hc0f603ce, 32'hc1ef5961} /* (8, 3, 15) {real, imag} */,
  {32'hc1add719, 32'hc0d40a90} /* (8, 3, 14) {real, imag} */,
  {32'hc1f2870c, 32'hc1a1cd8a} /* (8, 3, 13) {real, imag} */,
  {32'h41e84b5c, 32'hc1d5d845} /* (8, 3, 12) {real, imag} */,
  {32'h42169d26, 32'hc1c7cc70} /* (8, 3, 11) {real, imag} */,
  {32'h421c98df, 32'hc24872c4} /* (8, 3, 10) {real, imag} */,
  {32'hc2bb2927, 32'h42adc707} /* (8, 3, 9) {real, imag} */,
  {32'h42294e9f, 32'h42a30b08} /* (8, 3, 8) {real, imag} */,
  {32'hc1189e24, 32'hc2b58a0a} /* (8, 3, 7) {real, imag} */,
  {32'hc26bd1f4, 32'h422cfb82} /* (8, 3, 6) {real, imag} */,
  {32'h420e52dc, 32'h41bb442d} /* (8, 3, 5) {real, imag} */,
  {32'h42655dc1, 32'hc23038ac} /* (8, 3, 4) {real, imag} */,
  {32'h421abb78, 32'hc1760221} /* (8, 3, 3) {real, imag} */,
  {32'h431a5ab8, 32'h41c2288c} /* (8, 3, 2) {real, imag} */,
  {32'hc31b9b82, 32'h41d86e54} /* (8, 3, 1) {real, imag} */,
  {32'hc2843b3c, 32'hc278795a} /* (8, 3, 0) {real, imag} */,
  {32'h43ec60dd, 32'hc3a3915d} /* (8, 2, 31) {real, imag} */,
  {32'hc38b5d14, 32'h43a6623d} /* (8, 2, 30) {real, imag} */,
  {32'hc229269e, 32'hc2b1f4f1} /* (8, 2, 29) {real, imag} */,
  {32'hc206e064, 32'hc20fa7dc} /* (8, 2, 28) {real, imag} */,
  {32'hc18c42d4, 32'hc1425716} /* (8, 2, 27) {real, imag} */,
  {32'hc1ef4267, 32'h4256f146} /* (8, 2, 26) {real, imag} */,
  {32'h420e8564, 32'hc1e47d54} /* (8, 2, 25) {real, imag} */,
  {32'h3ea52b00, 32'h42eca7a3} /* (8, 2, 24) {real, imag} */,
  {32'h415485c2, 32'h41cc55cc} /* (8, 2, 23) {real, imag} */,
  {32'h41cac527, 32'hc0622378} /* (8, 2, 22) {real, imag} */,
  {32'h40113e50, 32'h412f9d40} /* (8, 2, 21) {real, imag} */,
  {32'h41835735, 32'hc1cfeb76} /* (8, 2, 20) {real, imag} */,
  {32'hc1b79892, 32'hc11ea2f3} /* (8, 2, 19) {real, imag} */,
  {32'hc0e3c328, 32'h40a10d90} /* (8, 2, 18) {real, imag} */,
  {32'hc21cb4aa, 32'h41358e42} /* (8, 2, 17) {real, imag} */,
  {32'hc19d1f50, 32'h3feef380} /* (8, 2, 16) {real, imag} */,
  {32'hbcab3000, 32'h421cd500} /* (8, 2, 15) {real, imag} */,
  {32'hc21b1bcb, 32'h418c7f6c} /* (8, 2, 14) {real, imag} */,
  {32'hc07baee0, 32'hc1e8c454} /* (8, 2, 13) {real, imag} */,
  {32'hc1b73dbb, 32'hc08970d8} /* (8, 2, 12) {real, imag} */,
  {32'hc297fb54, 32'hc2869a5e} /* (8, 2, 11) {real, imag} */,
  {32'hc19b4e91, 32'hc184dee9} /* (8, 2, 10) {real, imag} */,
  {32'hc25e4638, 32'h40fb36d0} /* (8, 2, 9) {real, imag} */,
  {32'hc302524c, 32'h41fffc14} /* (8, 2, 8) {real, imag} */,
  {32'h41c003d7, 32'hc1201158} /* (8, 2, 7) {real, imag} */,
  {32'h4294515e, 32'h41516a1a} /* (8, 2, 6) {real, imag} */,
  {32'hc31aaca2, 32'hc2514d8c} /* (8, 2, 5) {real, imag} */,
  {32'h431d287b, 32'hc31793b3} /* (8, 2, 4) {real, imag} */,
  {32'h4172692c, 32'hc2505156} /* (8, 2, 3) {real, imag} */,
  {32'hc295c910, 32'h43117414} /* (8, 2, 2) {real, imag} */,
  {32'h439cc651, 32'hc3a23a85} /* (8, 2, 1) {real, imag} */,
  {32'h439f12bb, 32'hc34ab2e5} /* (8, 2, 0) {real, imag} */,
  {32'hc3a97cdc, 32'h43ef71d8} /* (8, 1, 31) {real, imag} */,
  {32'hc1e35c30, 32'hc3487fc7} /* (8, 1, 30) {real, imag} */,
  {32'h40e25fcc, 32'h424f5e9d} /* (8, 1, 29) {real, imag} */,
  {32'hc2619988, 32'hc2488f35} /* (8, 1, 28) {real, imag} */,
  {32'h42c84090, 32'hc2f42c6f} /* (8, 1, 27) {real, imag} */,
  {32'hc2603869, 32'h4266a1e0} /* (8, 1, 26) {real, imag} */,
  {32'hc30e31fd, 32'h411eb520} /* (8, 1, 25) {real, imag} */,
  {32'hc1ccea3c, 32'hc2f46810} /* (8, 1, 24) {real, imag} */,
  {32'hc022dbb0, 32'h42549d80} /* (8, 1, 23) {real, imag} */,
  {32'hc24a442d, 32'h4158ba80} /* (8, 1, 22) {real, imag} */,
  {32'hc1c31106, 32'hc2d52058} /* (8, 1, 21) {real, imag} */,
  {32'hc2366bad, 32'hc2306e39} /* (8, 1, 20) {real, imag} */,
  {32'hc24a363c, 32'h409e383c} /* (8, 1, 19) {real, imag} */,
  {32'h41fa4d1c, 32'hc1715b24} /* (8, 1, 18) {real, imag} */,
  {32'h40f0be00, 32'h40e40e40} /* (8, 1, 17) {real, imag} */,
  {32'h40ab6220, 32'h3ff8b480} /* (8, 1, 16) {real, imag} */,
  {32'h4020b400, 32'h415a0b40} /* (8, 1, 15) {real, imag} */,
  {32'h41678a78, 32'h41719124} /* (8, 1, 14) {real, imag} */,
  {32'hc1b42600, 32'h409ecb4c} /* (8, 1, 13) {real, imag} */,
  {32'hc22706c3, 32'hc2a30ef6} /* (8, 1, 12) {real, imag} */,
  {32'h413f431c, 32'h41b422d2} /* (8, 1, 11) {real, imag} */,
  {32'hbf1b39c0, 32'h42592a1c} /* (8, 1, 10) {real, imag} */,
  {32'h3f997d60, 32'hc27b58d0} /* (8, 1, 9) {real, imag} */,
  {32'h42fbacfd, 32'h41466820} /* (8, 1, 8) {real, imag} */,
  {32'hc3215287, 32'hc1c1ac90} /* (8, 1, 7) {real, imag} */,
  {32'h4243b905, 32'h42248400} /* (8, 1, 6) {real, imag} */,
  {32'h434bd740, 32'hc19dcd9c} /* (8, 1, 5) {real, imag} */,
  {32'h4205f8fa, 32'hc3236678} /* (8, 1, 4) {real, imag} */,
  {32'h4234954a, 32'h4245f0d7} /* (8, 1, 3) {real, imag} */,
  {32'h43f48a1b, 32'hc282d6c2} /* (8, 1, 2) {real, imag} */,
  {32'hc4313580, 32'h43216347} /* (8, 1, 1) {real, imag} */,
  {32'hc3835188, 32'h43a391f8} /* (8, 1, 0) {real, imag} */,
  {32'hc33563f6, 32'h43ca9af3} /* (8, 0, 31) {real, imag} */,
  {32'hc20dcb76, 32'hc2b126bc} /* (8, 0, 30) {real, imag} */,
  {32'h428e316a, 32'h4250b6a8} /* (8, 0, 29) {real, imag} */,
  {32'hc2e37810, 32'hc19266bb} /* (8, 0, 28) {real, imag} */,
  {32'hc0da42e0, 32'hc2ec1c16} /* (8, 0, 27) {real, imag} */,
  {32'hc228f964, 32'hc294570a} /* (8, 0, 26) {real, imag} */,
  {32'h42ac9d5c, 32'h4288cbd3} /* (8, 0, 25) {real, imag} */,
  {32'hc2d38d82, 32'hc18c085a} /* (8, 0, 24) {real, imag} */,
  {32'h41f249ce, 32'h41d5c42c} /* (8, 0, 23) {real, imag} */,
  {32'hc0f76560, 32'hc14dca08} /* (8, 0, 22) {real, imag} */,
  {32'hc25b28a4, 32'hc1677b30} /* (8, 0, 21) {real, imag} */,
  {32'hc1cbcb25, 32'hc004cb18} /* (8, 0, 20) {real, imag} */,
  {32'h4022a6d0, 32'hc2026a1c} /* (8, 0, 19) {real, imag} */,
  {32'hc122d0aa, 32'h411f6fa0} /* (8, 0, 18) {real, imag} */,
  {32'hc189014a, 32'h40966ee0} /* (8, 0, 17) {real, imag} */,
  {32'hc192a52e, 32'h40b2b500} /* (8, 0, 16) {real, imag} */,
  {32'hc21c4bb3, 32'h422b2398} /* (8, 0, 15) {real, imag} */,
  {32'h42690062, 32'h426b3b2c} /* (8, 0, 14) {real, imag} */,
  {32'hc1a367e8, 32'hc1f07bd0} /* (8, 0, 13) {real, imag} */,
  {32'hc19833f9, 32'h41aa6b21} /* (8, 0, 12) {real, imag} */,
  {32'h420e4210, 32'hc18675f4} /* (8, 0, 11) {real, imag} */,
  {32'hc2af28b2, 32'hc2a4222b} /* (8, 0, 10) {real, imag} */,
  {32'h42046de9, 32'h420e0e5a} /* (8, 0, 9) {real, imag} */,
  {32'h42805624, 32'hc2692947} /* (8, 0, 8) {real, imag} */,
  {32'hc300ec64, 32'h42a60441} /* (8, 0, 7) {real, imag} */,
  {32'h42c0a852, 32'h42ab7964} /* (8, 0, 6) {real, imag} */,
  {32'h42e7a1b4, 32'hc279e395} /* (8, 0, 5) {real, imag} */,
  {32'hc12ac770, 32'h4204d0bc} /* (8, 0, 4) {real, imag} */,
  {32'h41dd4729, 32'hc301f19b} /* (8, 0, 3) {real, imag} */,
  {32'h42ffd7b3, 32'h42e10236} /* (8, 0, 2) {real, imag} */,
  {32'hc3ad76f9, 32'h42bc727c} /* (8, 0, 1) {real, imag} */,
  {32'hc30d681c, 32'h4348900f} /* (8, 0, 0) {real, imag} */,
  {32'h42b5c584, 32'hc31eda18} /* (7, 31, 31) {real, imag} */,
  {32'h42f87328, 32'h42a2f56c} /* (7, 31, 30) {real, imag} */,
  {32'hc363ad8c, 32'hc20570c0} /* (7, 31, 29) {real, imag} */,
  {32'h41825a50, 32'hc30a016b} /* (7, 31, 28) {real, imag} */,
  {32'h4272dda8, 32'h42ceb144} /* (7, 31, 27) {real, imag} */,
  {32'hc173b40e, 32'h42e5a7f4} /* (7, 31, 26) {real, imag} */,
  {32'hc130e090, 32'h4102357b} /* (7, 31, 25) {real, imag} */,
  {32'h4296102e, 32'hc1ea4e42} /* (7, 31, 24) {real, imag} */,
  {32'hc300646a, 32'hc0de7ad6} /* (7, 31, 23) {real, imag} */,
  {32'h426562bc, 32'hc10ef3d7} /* (7, 31, 22) {real, imag} */,
  {32'h4197413f, 32'h4175de9c} /* (7, 31, 21) {real, imag} */,
  {32'h40fb79d0, 32'h4215248c} /* (7, 31, 20) {real, imag} */,
  {32'h41e2a200, 32'hc1bc2a93} /* (7, 31, 19) {real, imag} */,
  {32'h41b5fa3c, 32'hc108c14c} /* (7, 31, 18) {real, imag} */,
  {32'h4155160c, 32'hc1789016} /* (7, 31, 17) {real, imag} */,
  {32'h4152a5cc, 32'hc0670cc0} /* (7, 31, 16) {real, imag} */,
  {32'h4141fbbc, 32'h403c1d68} /* (7, 31, 15) {real, imag} */,
  {32'h4208b74b, 32'h41c72c8e} /* (7, 31, 14) {real, imag} */,
  {32'h41a469f8, 32'h419ea475} /* (7, 31, 13) {real, imag} */,
  {32'hc1aeed44, 32'h410f0ae9} /* (7, 31, 12) {real, imag} */,
  {32'hc201637c, 32'h4228f2a6} /* (7, 31, 11) {real, imag} */,
  {32'hc25f00a4, 32'hc17cb691} /* (7, 31, 10) {real, imag} */,
  {32'h40cf1460, 32'h420bc873} /* (7, 31, 9) {real, imag} */,
  {32'hc17aa620, 32'h41de1d9a} /* (7, 31, 8) {real, imag} */,
  {32'hc28cd32c, 32'hc10cf255} /* (7, 31, 7) {real, imag} */,
  {32'h421d6edc, 32'h428cf708} /* (7, 31, 6) {real, imag} */,
  {32'hc2b453ba, 32'h41ace108} /* (7, 31, 5) {real, imag} */,
  {32'hc30c4383, 32'hc2fe5df2} /* (7, 31, 4) {real, imag} */,
  {32'hbe41a400, 32'hc277a3e8} /* (7, 31, 3) {real, imag} */,
  {32'h41e0acf0, 32'h43187d83} /* (7, 31, 2) {real, imag} */,
  {32'hc230f503, 32'h42826233} /* (7, 31, 1) {real, imag} */,
  {32'hc2b84076, 32'hc2a83466} /* (7, 31, 0) {real, imag} */,
  {32'hc238847a, 32'h41ea0a7c} /* (7, 30, 31) {real, imag} */,
  {32'hc1d1a5fa, 32'hc1170d60} /* (7, 30, 30) {real, imag} */,
  {32'h41df9a5e, 32'hc2e133ab} /* (7, 30, 29) {real, imag} */,
  {32'hc1f40e94, 32'hc2801cc9} /* (7, 30, 28) {real, imag} */,
  {32'h4241a6a2, 32'h4194124a} /* (7, 30, 27) {real, imag} */,
  {32'h42ce9746, 32'h410acb25} /* (7, 30, 26) {real, imag} */,
  {32'hc2f26f72, 32'hc298d1e2} /* (7, 30, 25) {real, imag} */,
  {32'h427be559, 32'hc21925dc} /* (7, 30, 24) {real, imag} */,
  {32'hc225a0f1, 32'hc28d376c} /* (7, 30, 23) {real, imag} */,
  {32'hc266c332, 32'h429aaa75} /* (7, 30, 22) {real, imag} */,
  {32'hc1a05e2d, 32'h42237fa7} /* (7, 30, 21) {real, imag} */,
  {32'hc189cd80, 32'h4295ae08} /* (7, 30, 20) {real, imag} */,
  {32'hc14c8b73, 32'h419d8cc0} /* (7, 30, 19) {real, imag} */,
  {32'hc1009174, 32'h40723658} /* (7, 30, 18) {real, imag} */,
  {32'h41d8d4b4, 32'hc1d63f87} /* (7, 30, 17) {real, imag} */,
  {32'h419f6ae8, 32'h41441bf8} /* (7, 30, 16) {real, imag} */,
  {32'h41a7a674, 32'h41ee0ad7} /* (7, 30, 15) {real, imag} */,
  {32'h426b3047, 32'h40f3842c} /* (7, 30, 14) {real, imag} */,
  {32'hc0bd04aa, 32'hbf867000} /* (7, 30, 13) {real, imag} */,
  {32'hc106cc9f, 32'hc0f10980} /* (7, 30, 12) {real, imag} */,
  {32'h3fffd500, 32'h4145317c} /* (7, 30, 11) {real, imag} */,
  {32'h4286b0c6, 32'hc26345cf} /* (7, 30, 10) {real, imag} */,
  {32'h41f3924e, 32'h4117a2dc} /* (7, 30, 9) {real, imag} */,
  {32'h41edcde6, 32'hc19cfd8f} /* (7, 30, 8) {real, imag} */,
  {32'hc2590a1c, 32'h4220e17f} /* (7, 30, 7) {real, imag} */,
  {32'hc3267c09, 32'h4043fa14} /* (7, 30, 6) {real, imag} */,
  {32'h41419120, 32'hc18057b0} /* (7, 30, 5) {real, imag} */,
  {32'hc2b23317, 32'hc3008d76} /* (7, 30, 4) {real, imag} */,
  {32'h42b6a7b6, 32'hc285fd2b} /* (7, 30, 3) {real, imag} */,
  {32'h41623297, 32'h43105f48} /* (7, 30, 2) {real, imag} */,
  {32'h42dcf233, 32'h42f28c85} /* (7, 30, 1) {real, imag} */,
  {32'hc2a16148, 32'h4354609c} /* (7, 30, 0) {real, imag} */,
  {32'h416bafb6, 32'h42371e30} /* (7, 29, 31) {real, imag} */,
  {32'hc305a3ec, 32'hc13fda7c} /* (7, 29, 30) {real, imag} */,
  {32'hc28fefb0, 32'hc1c6b946} /* (7, 29, 29) {real, imag} */,
  {32'hc269018a, 32'hc1ff5687} /* (7, 29, 28) {real, imag} */,
  {32'h430d5c06, 32'hc1a8d59c} /* (7, 29, 27) {real, imag} */,
  {32'h4142861a, 32'h42fe8193} /* (7, 29, 26) {real, imag} */,
  {32'hc2abbda9, 32'h4194f54c} /* (7, 29, 25) {real, imag} */,
  {32'h417702b2, 32'h3e8fd3c0} /* (7, 29, 24) {real, imag} */,
  {32'h42136ca8, 32'h4197544c} /* (7, 29, 23) {real, imag} */,
  {32'hc224beae, 32'hc2a31d1d} /* (7, 29, 22) {real, imag} */,
  {32'h40391620, 32'hc1408f40} /* (7, 29, 21) {real, imag} */,
  {32'hc128797e, 32'h3e073680} /* (7, 29, 20) {real, imag} */,
  {32'hc012bc4c, 32'h41dc3b72} /* (7, 29, 19) {real, imag} */,
  {32'hc16da4dc, 32'hc1bc094c} /* (7, 29, 18) {real, imag} */,
  {32'h4124b718, 32'h3fe6b870} /* (7, 29, 17) {real, imag} */,
  {32'h41ce1470, 32'h41375d30} /* (7, 29, 16) {real, imag} */,
  {32'hc1abdf74, 32'h41a54e5f} /* (7, 29, 15) {real, imag} */,
  {32'hbf8af560, 32'hc241f156} /* (7, 29, 14) {real, imag} */,
  {32'hc0c24206, 32'h41bf0f38} /* (7, 29, 13) {real, imag} */,
  {32'hc0da6a94, 32'h424148a0} /* (7, 29, 12) {real, imag} */,
  {32'hc1d4bb24, 32'h4243d6f3} /* (7, 29, 11) {real, imag} */,
  {32'hc0c124c4, 32'h41f5fb5c} /* (7, 29, 10) {real, imag} */,
  {32'hc2348ffc, 32'hc2721f52} /* (7, 29, 9) {real, imag} */,
  {32'h4207ff32, 32'h41d423bb} /* (7, 29, 8) {real, imag} */,
  {32'h42566eca, 32'h42b9e12f} /* (7, 29, 7) {real, imag} */,
  {32'hc29071e1, 32'hc0cb1190} /* (7, 29, 6) {real, imag} */,
  {32'hc1d6f958, 32'h4324e052} /* (7, 29, 5) {real, imag} */,
  {32'hc2822eea, 32'hc20c4ef4} /* (7, 29, 4) {real, imag} */,
  {32'h41d70a8a, 32'h3dfa7400} /* (7, 29, 3) {real, imag} */,
  {32'h41c08108, 32'hc217dfad} /* (7, 29, 2) {real, imag} */,
  {32'hc21aa320, 32'h41f0a477} /* (7, 29, 1) {real, imag} */,
  {32'hc311304e, 32'h427b8224} /* (7, 29, 0) {real, imag} */,
  {32'hc1d7a605, 32'h4297f762} /* (7, 28, 31) {real, imag} */,
  {32'hc1efba06, 32'h4237189d} /* (7, 28, 30) {real, imag} */,
  {32'h419ec4f5, 32'hc2c51aba} /* (7, 28, 29) {real, imag} */,
  {32'h4302fbd8, 32'hc08ec4ed} /* (7, 28, 28) {real, imag} */,
  {32'hc2b6c438, 32'hc0f5a364} /* (7, 28, 27) {real, imag} */,
  {32'hbf83d580, 32'h42bf9a90} /* (7, 28, 26) {real, imag} */,
  {32'h4194a884, 32'h426bf5b8} /* (7, 28, 25) {real, imag} */,
  {32'hc28568e7, 32'h42a05d36} /* (7, 28, 24) {real, imag} */,
  {32'h42621612, 32'hc0d7d64c} /* (7, 28, 23) {real, imag} */,
  {32'h42a5998a, 32'hc14ecbf8} /* (7, 28, 22) {real, imag} */,
  {32'hc250b300, 32'h4184f71a} /* (7, 28, 21) {real, imag} */,
  {32'hc2026253, 32'h416d58c8} /* (7, 28, 20) {real, imag} */,
  {32'h41b44b6c, 32'hc1c5b182} /* (7, 28, 19) {real, imag} */,
  {32'hc16e6ba4, 32'hc1846977} /* (7, 28, 18) {real, imag} */,
  {32'h41256228, 32'h4178d9c5} /* (7, 28, 17) {real, imag} */,
  {32'hc19b683d, 32'h42064a2f} /* (7, 28, 16) {real, imag} */,
  {32'hc0b5c55c, 32'h3fe8aa68} /* (7, 28, 15) {real, imag} */,
  {32'hc11f25c4, 32'h4106fb52} /* (7, 28, 14) {real, imag} */,
  {32'h40817ace, 32'h422c6fcb} /* (7, 28, 13) {real, imag} */,
  {32'hc0b139ea, 32'h415a33dc} /* (7, 28, 12) {real, imag} */,
  {32'h42538a42, 32'hc249b8a3} /* (7, 28, 11) {real, imag} */,
  {32'h41998901, 32'h423267f2} /* (7, 28, 10) {real, imag} */,
  {32'h42140cba, 32'hc2527130} /* (7, 28, 9) {real, imag} */,
  {32'hc20ba47a, 32'hc195a532} /* (7, 28, 8) {real, imag} */,
  {32'hc10bcf98, 32'hc120ff16} /* (7, 28, 7) {real, imag} */,
  {32'hc20a1dcd, 32'hc3129870} /* (7, 28, 6) {real, imag} */,
  {32'hc22e2681, 32'h425c61ea} /* (7, 28, 5) {real, imag} */,
  {32'h426be228, 32'hc0c927a5} /* (7, 28, 4) {real, imag} */,
  {32'h41abd557, 32'h42265b1b} /* (7, 28, 3) {real, imag} */,
  {32'h3ea56780, 32'hc2603a77} /* (7, 28, 2) {real, imag} */,
  {32'hc1ea1817, 32'hc2095a17} /* (7, 28, 1) {real, imag} */,
  {32'h41bbfffd, 32'hc300b0e1} /* (7, 28, 0) {real, imag} */,
  {32'hc2a4955d, 32'h42b88ce6} /* (7, 27, 31) {real, imag} */,
  {32'h41cfab74, 32'h424ec8b8} /* (7, 27, 30) {real, imag} */,
  {32'h42151427, 32'hc290869c} /* (7, 27, 29) {real, imag} */,
  {32'hc0f50088, 32'hc31f07f5} /* (7, 27, 28) {real, imag} */,
  {32'h411238c0, 32'h42762e4e} /* (7, 27, 27) {real, imag} */,
  {32'h40cdc388, 32'hc1887530} /* (7, 27, 26) {real, imag} */,
  {32'h413dc588, 32'h42398dfb} /* (7, 27, 25) {real, imag} */,
  {32'hc220fb88, 32'h40f09de0} /* (7, 27, 24) {real, imag} */,
  {32'h42061de4, 32'h42f06502} /* (7, 27, 23) {real, imag} */,
  {32'h3e93c1c0, 32'hc134f4f0} /* (7, 27, 22) {real, imag} */,
  {32'hc202909e, 32'hc1c0db73} /* (7, 27, 21) {real, imag} */,
  {32'hc1c9395e, 32'h41a67e4e} /* (7, 27, 20) {real, imag} */,
  {32'h411a0fa4, 32'hc14239da} /* (7, 27, 19) {real, imag} */,
  {32'h423194da, 32'hc0c49de6} /* (7, 27, 18) {real, imag} */,
  {32'hc048d2ae, 32'hbfedb66e} /* (7, 27, 17) {real, imag} */,
  {32'hc12b6be0, 32'hc12c3294} /* (7, 27, 16) {real, imag} */,
  {32'h410f59bc, 32'hc045de97} /* (7, 27, 15) {real, imag} */,
  {32'h3f4a2680, 32'hc025178c} /* (7, 27, 14) {real, imag} */,
  {32'hc1c4a5ba, 32'hc1768c32} /* (7, 27, 13) {real, imag} */,
  {32'hc1d75934, 32'h420e7bef} /* (7, 27, 12) {real, imag} */,
  {32'h42033086, 32'hc1921d41} /* (7, 27, 11) {real, imag} */,
  {32'hc268f056, 32'h423d28d4} /* (7, 27, 10) {real, imag} */,
  {32'h427f6004, 32'hc1a39232} /* (7, 27, 9) {real, imag} */,
  {32'hc0846494, 32'h428ed6a1} /* (7, 27, 8) {real, imag} */,
  {32'h418142f8, 32'h4233bf5b} /* (7, 27, 7) {real, imag} */,
  {32'h42dc0e4a, 32'hc30d2646} /* (7, 27, 6) {real, imag} */,
  {32'hc2822d1e, 32'h4131db3e} /* (7, 27, 5) {real, imag} */,
  {32'hc291bc22, 32'h43134a4b} /* (7, 27, 4) {real, imag} */,
  {32'hc126ab4c, 32'h428e5514} /* (7, 27, 3) {real, imag} */,
  {32'hc2da62d7, 32'hc28327c2} /* (7, 27, 2) {real, imag} */,
  {32'hc2cfc38b, 32'hc2abfb7e} /* (7, 27, 1) {real, imag} */,
  {32'h42cfe4fb, 32'h42d265b8} /* (7, 27, 0) {real, imag} */,
  {32'hc2a1af88, 32'h42bdc484} /* (7, 26, 31) {real, imag} */,
  {32'hc0f49bfc, 32'hc1c17162} /* (7, 26, 30) {real, imag} */,
  {32'h41dc204e, 32'h42208c7f} /* (7, 26, 29) {real, imag} */,
  {32'hc2a9d5e6, 32'hc11e60d8} /* (7, 26, 28) {real, imag} */,
  {32'hc2580094, 32'hc28eba4f} /* (7, 26, 27) {real, imag} */,
  {32'hc26fe55a, 32'hc24d8461} /* (7, 26, 26) {real, imag} */,
  {32'h4271fd86, 32'hc202f060} /* (7, 26, 25) {real, imag} */,
  {32'hc1def2a6, 32'h3e3b5080} /* (7, 26, 24) {real, imag} */,
  {32'h4082287c, 32'h41f51a9a} /* (7, 26, 23) {real, imag} */,
  {32'hc25ca0fe, 32'hc27232ce} /* (7, 26, 22) {real, imag} */,
  {32'hc0a5739a, 32'hc266bede} /* (7, 26, 21) {real, imag} */,
  {32'h42660b4d, 32'hc1aab17d} /* (7, 26, 20) {real, imag} */,
  {32'hc1d7bd56, 32'hbf886178} /* (7, 26, 19) {real, imag} */,
  {32'hc1b0d4eb, 32'h4201336e} /* (7, 26, 18) {real, imag} */,
  {32'h4076497c, 32'h41238cf8} /* (7, 26, 17) {real, imag} */,
  {32'hc1878b4f, 32'hc1abac9c} /* (7, 26, 16) {real, imag} */,
  {32'hc0e0b3de, 32'h40fbf010} /* (7, 26, 15) {real, imag} */,
  {32'h41f51d8f, 32'h41745dbe} /* (7, 26, 14) {real, imag} */,
  {32'h427330cf, 32'hc1a4d12c} /* (7, 26, 13) {real, imag} */,
  {32'hc1402b94, 32'hc22fc7c6} /* (7, 26, 12) {real, imag} */,
  {32'hc150162d, 32'h420d12b2} /* (7, 26, 11) {real, imag} */,
  {32'hbf25cfc0, 32'h41ae1cfc} /* (7, 26, 10) {real, imag} */,
  {32'hc27f006a, 32'hbfcc7968} /* (7, 26, 9) {real, imag} */,
  {32'h40aabe58, 32'h420a5222} /* (7, 26, 8) {real, imag} */,
  {32'hc2b54a0d, 32'h419cc3cc} /* (7, 26, 7) {real, imag} */,
  {32'h41df320b, 32'h4226fde3} /* (7, 26, 6) {real, imag} */,
  {32'h42816bda, 32'hbf8f9c40} /* (7, 26, 5) {real, imag} */,
  {32'hc1e75c92, 32'hc2e4088b} /* (7, 26, 4) {real, imag} */,
  {32'hc280c5b4, 32'h420db107} /* (7, 26, 3) {real, imag} */,
  {32'h4046c018, 32'h40d9cb12} /* (7, 26, 2) {real, imag} */,
  {32'hc19cbba0, 32'h4184ceee} /* (7, 26, 1) {real, imag} */,
  {32'hbf4b3fa0, 32'h414411b0} /* (7, 26, 0) {real, imag} */,
  {32'h42c43d52, 32'h422bf0ae} /* (7, 25, 31) {real, imag} */,
  {32'hc215e339, 32'h41ee9bce} /* (7, 25, 30) {real, imag} */,
  {32'h4223c2f3, 32'h420ad4c0} /* (7, 25, 29) {real, imag} */,
  {32'hc2bf39c3, 32'hc2a8b5ad} /* (7, 25, 28) {real, imag} */,
  {32'h3f8f0a40, 32'h4261e623} /* (7, 25, 27) {real, imag} */,
  {32'h42340359, 32'hc1f5e4bb} /* (7, 25, 26) {real, imag} */,
  {32'hc2306ade, 32'hc09eae44} /* (7, 25, 25) {real, imag} */,
  {32'hc203a5b2, 32'h421cd770} /* (7, 25, 24) {real, imag} */,
  {32'h419109e6, 32'hc21f407e} /* (7, 25, 23) {real, imag} */,
  {32'hc21af501, 32'hc132321c} /* (7, 25, 22) {real, imag} */,
  {32'h3f61a680, 32'h4027d27c} /* (7, 25, 21) {real, imag} */,
  {32'hc1ae0547, 32'hc19156b5} /* (7, 25, 20) {real, imag} */,
  {32'hc2356a36, 32'hc193d2da} /* (7, 25, 19) {real, imag} */,
  {32'h40b5ac6e, 32'hc207406f} /* (7, 25, 18) {real, imag} */,
  {32'hc1035790, 32'h41e032ca} /* (7, 25, 17) {real, imag} */,
  {32'h41edae04, 32'h413cf1da} /* (7, 25, 16) {real, imag} */,
  {32'h42005d48, 32'h40c38ae8} /* (7, 25, 15) {real, imag} */,
  {32'h40f26ba2, 32'h3ee16480} /* (7, 25, 14) {real, imag} */,
  {32'h416e76c5, 32'hc2089d01} /* (7, 25, 13) {real, imag} */,
  {32'h421bca2e, 32'h421cd278} /* (7, 25, 12) {real, imag} */,
  {32'hc206b1a4, 32'hc18276a0} /* (7, 25, 11) {real, imag} */,
  {32'h423d4089, 32'h424717d2} /* (7, 25, 10) {real, imag} */,
  {32'h415ae816, 32'h41936bde} /* (7, 25, 9) {real, imag} */,
  {32'hc1834ad8, 32'hc1fd22d3} /* (7, 25, 8) {real, imag} */,
  {32'hc15c1146, 32'h423cd596} /* (7, 25, 7) {real, imag} */,
  {32'h428fea0e, 32'h429a135d} /* (7, 25, 6) {real, imag} */,
  {32'hc29e2c88, 32'hc0645d50} /* (7, 25, 5) {real, imag} */,
  {32'h429f1629, 32'h42eb6efb} /* (7, 25, 4) {real, imag} */,
  {32'hc1556069, 32'h41ed471c} /* (7, 25, 3) {real, imag} */,
  {32'hc236cce5, 32'h4243c267} /* (7, 25, 2) {real, imag} */,
  {32'hc299cf30, 32'h4056cec8} /* (7, 25, 1) {real, imag} */,
  {32'h425a7054, 32'hc1b9784f} /* (7, 25, 0) {real, imag} */,
  {32'hc296c00e, 32'hc22d0075} /* (7, 24, 31) {real, imag} */,
  {32'h3f856060, 32'h42632b5c} /* (7, 24, 30) {real, imag} */,
  {32'h41982cc1, 32'h42959514} /* (7, 24, 29) {real, imag} */,
  {32'h425a8ee7, 32'hc0ab6b4c} /* (7, 24, 28) {real, imag} */,
  {32'h42aa5a32, 32'h428006c4} /* (7, 24, 27) {real, imag} */,
  {32'h4251bb2a, 32'hc1f05af8} /* (7, 24, 26) {real, imag} */,
  {32'h432a4379, 32'hc0e4bb80} /* (7, 24, 25) {real, imag} */,
  {32'hc1187ed8, 32'hc1a2b7e6} /* (7, 24, 24) {real, imag} */,
  {32'h40cae838, 32'hbf2ba2c0} /* (7, 24, 23) {real, imag} */,
  {32'hc205980e, 32'h41c12809} /* (7, 24, 22) {real, imag} */,
  {32'h3f796d00, 32'h40d9e252} /* (7, 24, 21) {real, imag} */,
  {32'h41041412, 32'h4202cb76} /* (7, 24, 20) {real, imag} */,
  {32'h410a1572, 32'h40906702} /* (7, 24, 19) {real, imag} */,
  {32'hbf4ddeb0, 32'hc21a2d9c} /* (7, 24, 18) {real, imag} */,
  {32'hc0e59f5c, 32'h4015dd50} /* (7, 24, 17) {real, imag} */,
  {32'h401dec7c, 32'h40579d10} /* (7, 24, 16) {real, imag} */,
  {32'h41395d76, 32'h41c56554} /* (7, 24, 15) {real, imag} */,
  {32'h3f3c3870, 32'h3ee79ec0} /* (7, 24, 14) {real, imag} */,
  {32'h419e365b, 32'hc18980e4} /* (7, 24, 13) {real, imag} */,
  {32'hc1513b32, 32'h42543b4a} /* (7, 24, 12) {real, imag} */,
  {32'h4099eb20, 32'hc1bd183c} /* (7, 24, 11) {real, imag} */,
  {32'hc26dad7a, 32'hc283cc07} /* (7, 24, 10) {real, imag} */,
  {32'hc270cc7b, 32'hc1927864} /* (7, 24, 9) {real, imag} */,
  {32'hc1f6decc, 32'hc1b4c59e} /* (7, 24, 8) {real, imag} */,
  {32'h42b37c96, 32'hc241bb7d} /* (7, 24, 7) {real, imag} */,
  {32'hc1c341e8, 32'h4232fcfe} /* (7, 24, 6) {real, imag} */,
  {32'hc24a916b, 32'h4122c0a4} /* (7, 24, 5) {real, imag} */,
  {32'hc24593dd, 32'h425c64e2} /* (7, 24, 4) {real, imag} */,
  {32'h42947456, 32'hc1e79b40} /* (7, 24, 3) {real, imag} */,
  {32'hc27fb875, 32'h410b3ec2} /* (7, 24, 2) {real, imag} */,
  {32'hc1eae67b, 32'h4237ca37} /* (7, 24, 1) {real, imag} */,
  {32'h40ef6634, 32'hc2d34e44} /* (7, 24, 0) {real, imag} */,
  {32'hc265ace8, 32'h428fe8c4} /* (7, 23, 31) {real, imag} */,
  {32'h42a02f5c, 32'hc229ce20} /* (7, 23, 30) {real, imag} */,
  {32'h3fb2e890, 32'hc2cf3024} /* (7, 23, 29) {real, imag} */,
  {32'h428b9538, 32'h4239c86d} /* (7, 23, 28) {real, imag} */,
  {32'hc26aa0b8, 32'h41f4b758} /* (7, 23, 27) {real, imag} */,
  {32'hc200d712, 32'hc28f58a0} /* (7, 23, 26) {real, imag} */,
  {32'h40077794, 32'hc1c4ee5e} /* (7, 23, 25) {real, imag} */,
  {32'h41afd0a8, 32'hc1a22fe2} /* (7, 23, 24) {real, imag} */,
  {32'hc285a116, 32'h420efad0} /* (7, 23, 23) {real, imag} */,
  {32'h427b5c34, 32'hc19d5bb4} /* (7, 23, 22) {real, imag} */,
  {32'hc05427f8, 32'h4163bbdd} /* (7, 23, 21) {real, imag} */,
  {32'hc18a0fc3, 32'hc0def6e4} /* (7, 23, 20) {real, imag} */,
  {32'h41f8dfda, 32'hc10d7c3c} /* (7, 23, 19) {real, imag} */,
  {32'h406ca8b0, 32'h41d61990} /* (7, 23, 18) {real, imag} */,
  {32'h411cbc1e, 32'h41b00191} /* (7, 23, 17) {real, imag} */,
  {32'h410b89ff, 32'hbfef0d10} /* (7, 23, 16) {real, imag} */,
  {32'h3fa17294, 32'hc03c59c8} /* (7, 23, 15) {real, imag} */,
  {32'hc11fb214, 32'hc118058f} /* (7, 23, 14) {real, imag} */,
  {32'hc2349329, 32'h3f5ef600} /* (7, 23, 13) {real, imag} */,
  {32'hc0abbfec, 32'h40601960} /* (7, 23, 12) {real, imag} */,
  {32'h4102469a, 32'h4178a527} /* (7, 23, 11) {real, imag} */,
  {32'hc12559a0, 32'h4184d80a} /* (7, 23, 10) {real, imag} */,
  {32'h40fba7f8, 32'h40a3e70a} /* (7, 23, 9) {real, imag} */,
  {32'h421de295, 32'h400d2f6c} /* (7, 23, 8) {real, imag} */,
  {32'hc0b0552e, 32'hc294778c} /* (7, 23, 7) {real, imag} */,
  {32'hc0eb92f2, 32'h419ed8e7} /* (7, 23, 6) {real, imag} */,
  {32'h41ead40b, 32'h41413283} /* (7, 23, 5) {real, imag} */,
  {32'hc199a36b, 32'hc0089cf0} /* (7, 23, 4) {real, imag} */,
  {32'hc1186be6, 32'hc01b5740} /* (7, 23, 3) {real, imag} */,
  {32'h420f2ce9, 32'h416e6737} /* (7, 23, 2) {real, imag} */,
  {32'h427d2728, 32'h42978a5a} /* (7, 23, 1) {real, imag} */,
  {32'hc176a613, 32'hc18fc4f7} /* (7, 23, 0) {real, imag} */,
  {32'h421f3f3e, 32'hc26ed494} /* (7, 22, 31) {real, imag} */,
  {32'h4216fea4, 32'hc2acad50} /* (7, 22, 30) {real, imag} */,
  {32'hc2855a22, 32'h427597e1} /* (7, 22, 29) {real, imag} */,
  {32'h4265006e, 32'h4231950f} /* (7, 22, 28) {real, imag} */,
  {32'hc22fb103, 32'h418806e2} /* (7, 22, 27) {real, imag} */,
  {32'hc24a98cd, 32'hc2237f2e} /* (7, 22, 26) {real, imag} */,
  {32'hbfd4ca58, 32'hc09cf54c} /* (7, 22, 25) {real, imag} */,
  {32'h4030f55c, 32'hc205d1bd} /* (7, 22, 24) {real, imag} */,
  {32'hc13232c6, 32'h4236c8e3} /* (7, 22, 23) {real, imag} */,
  {32'hc17104f6, 32'h41240c76} /* (7, 22, 22) {real, imag} */,
  {32'h412e3329, 32'hc1ded282} /* (7, 22, 21) {real, imag} */,
  {32'h415190d0, 32'h41df94ac} /* (7, 22, 20) {real, imag} */,
  {32'hc18872ea, 32'hc1d273e4} /* (7, 22, 19) {real, imag} */,
  {32'h405b7ee4, 32'h413075b9} /* (7, 22, 18) {real, imag} */,
  {32'hc101b3c9, 32'h408fb663} /* (7, 22, 17) {real, imag} */,
  {32'h4123e542, 32'h41b6a0f2} /* (7, 22, 16) {real, imag} */,
  {32'h4094a736, 32'h41027d02} /* (7, 22, 15) {real, imag} */,
  {32'hc186a09e, 32'h407b62a4} /* (7, 22, 14) {real, imag} */,
  {32'hc0e810d8, 32'h41a48c80} /* (7, 22, 13) {real, imag} */,
  {32'h4183a155, 32'h3e3d6940} /* (7, 22, 12) {real, imag} */,
  {32'hc0ac810a, 32'hc02d7188} /* (7, 22, 11) {real, imag} */,
  {32'hc243d6f2, 32'h419594f8} /* (7, 22, 10) {real, imag} */,
  {32'h42426510, 32'hc2667f5d} /* (7, 22, 9) {real, imag} */,
  {32'h3ffe81b8, 32'hc1660e61} /* (7, 22, 8) {real, imag} */,
  {32'h3ec05b20, 32'hc26f7462} /* (7, 22, 7) {real, imag} */,
  {32'h421f7257, 32'hc1ee52a3} /* (7, 22, 6) {real, imag} */,
  {32'hc02e6930, 32'hc199e17a} /* (7, 22, 5) {real, imag} */,
  {32'h41d462ac, 32'h428fa563} /* (7, 22, 4) {real, imag} */,
  {32'hc1498eb4, 32'h41de6402} /* (7, 22, 3) {real, imag} */,
  {32'h40503338, 32'h42f6855a} /* (7, 22, 2) {real, imag} */,
  {32'h401143f8, 32'h4183fc17} /* (7, 22, 1) {real, imag} */,
  {32'h40d33650, 32'hc1f09cea} /* (7, 22, 0) {real, imag} */,
  {32'h427bf42c, 32'hc2615415} /* (7, 21, 31) {real, imag} */,
  {32'hc1e02568, 32'hbf7cea08} /* (7, 21, 30) {real, imag} */,
  {32'hc16d7a7e, 32'hc21ab8a1} /* (7, 21, 29) {real, imag} */,
  {32'h41810960, 32'h422de64e} /* (7, 21, 28) {real, imag} */,
  {32'hc28d2ca1, 32'hbfedaab8} /* (7, 21, 27) {real, imag} */,
  {32'h41adffae, 32'hc0c86820} /* (7, 21, 26) {real, imag} */,
  {32'hc13c6b9f, 32'h41f8d717} /* (7, 21, 25) {real, imag} */,
  {32'hc2006ffa, 32'h41888868} /* (7, 21, 24) {real, imag} */,
  {32'h4186fa85, 32'hc2422324} /* (7, 21, 23) {real, imag} */,
  {32'h40606448, 32'h41c693c6} /* (7, 21, 22) {real, imag} */,
  {32'h4203e164, 32'h40af216d} /* (7, 21, 21) {real, imag} */,
  {32'hc1269b35, 32'hc1a355f7} /* (7, 21, 20) {real, imag} */,
  {32'h41731dea, 32'hc10c2253} /* (7, 21, 19) {real, imag} */,
  {32'h413043d8, 32'h4073704c} /* (7, 21, 18) {real, imag} */,
  {32'hc16c958a, 32'hc0549410} /* (7, 21, 17) {real, imag} */,
  {32'hc0cbf4ad, 32'hc148b5a6} /* (7, 21, 16) {real, imag} */,
  {32'hc025ff78, 32'h41b7fd0e} /* (7, 21, 15) {real, imag} */,
  {32'hc18bc499, 32'hc1a9aeb6} /* (7, 21, 14) {real, imag} */,
  {32'hc1211072, 32'hc0af68fa} /* (7, 21, 13) {real, imag} */,
  {32'hc1a05a5c, 32'h418387d3} /* (7, 21, 12) {real, imag} */,
  {32'hc1a4f2b5, 32'hc116265c} /* (7, 21, 11) {real, imag} */,
  {32'h40b2c3a8, 32'hc18ead9e} /* (7, 21, 10) {real, imag} */,
  {32'h422df75c, 32'h40970444} /* (7, 21, 9) {real, imag} */,
  {32'hc1d24664, 32'hc13e5e10} /* (7, 21, 8) {real, imag} */,
  {32'h422ef9db, 32'h409cd8ac} /* (7, 21, 7) {real, imag} */,
  {32'h4211bbfb, 32'hc1c02740} /* (7, 21, 6) {real, imag} */,
  {32'hc0784ce0, 32'hc1dcdf56} /* (7, 21, 5) {real, imag} */,
  {32'h421e94a9, 32'h40f163f8} /* (7, 21, 4) {real, imag} */,
  {32'hc24db34c, 32'hc05e71b0} /* (7, 21, 3) {real, imag} */,
  {32'h41d11d1c, 32'hc116652e} /* (7, 21, 2) {real, imag} */,
  {32'hc191ecc0, 32'hc152ac54} /* (7, 21, 1) {real, imag} */,
  {32'hc07693e6, 32'hc123c16e} /* (7, 21, 0) {real, imag} */,
  {32'h3fb45098, 32'hc0bf9ee0} /* (7, 20, 31) {real, imag} */,
  {32'hc0e53b70, 32'h416012ef} /* (7, 20, 30) {real, imag} */,
  {32'h41db934c, 32'h41a5bafc} /* (7, 20, 29) {real, imag} */,
  {32'h40223b87, 32'hc22c1cca} /* (7, 20, 28) {real, imag} */,
  {32'h41c898ac, 32'h4036c530} /* (7, 20, 27) {real, imag} */,
  {32'hc1b82773, 32'h4197b022} /* (7, 20, 26) {real, imag} */,
  {32'hc0b6f48a, 32'hc1521a50} /* (7, 20, 25) {real, imag} */,
  {32'h4121c44d, 32'h4256f7e6} /* (7, 20, 24) {real, imag} */,
  {32'h40355ddc, 32'hc0411b44} /* (7, 20, 23) {real, imag} */,
  {32'h4146250c, 32'h4211e0ae} /* (7, 20, 22) {real, imag} */,
  {32'h4135c048, 32'h3ef3fb80} /* (7, 20, 21) {real, imag} */,
  {32'hc1e75bf7, 32'h416993a8} /* (7, 20, 20) {real, imag} */,
  {32'h4063e8b2, 32'hbfb37864} /* (7, 20, 19) {real, imag} */,
  {32'hc003cafc, 32'h41947e8e} /* (7, 20, 18) {real, imag} */,
  {32'hc10d8517, 32'hc123b082} /* (7, 20, 17) {real, imag} */,
  {32'h41084df8, 32'h3f972d18} /* (7, 20, 16) {real, imag} */,
  {32'hbfbb182a, 32'hc0c8690c} /* (7, 20, 15) {real, imag} */,
  {32'hc045881c, 32'h40bac1fe} /* (7, 20, 14) {real, imag} */,
  {32'hc12c8284, 32'hc10fb72c} /* (7, 20, 13) {real, imag} */,
  {32'hc13ffbba, 32'hc21457f8} /* (7, 20, 12) {real, imag} */,
  {32'hc187e802, 32'h4142cdcc} /* (7, 20, 11) {real, imag} */,
  {32'hc0595f16, 32'h4159b743} /* (7, 20, 10) {real, imag} */,
  {32'hc20947c0, 32'h41e21120} /* (7, 20, 9) {real, imag} */,
  {32'hc2033bdf, 32'hc1028fa6} /* (7, 20, 8) {real, imag} */,
  {32'h41988034, 32'h4233ee16} /* (7, 20, 7) {real, imag} */,
  {32'hc23aff74, 32'hc064533c} /* (7, 20, 6) {real, imag} */,
  {32'h40c499a8, 32'hc1354124} /* (7, 20, 5) {real, imag} */,
  {32'h407a50c1, 32'hc23ecd2c} /* (7, 20, 4) {real, imag} */,
  {32'hc1b75b20, 32'hc07a0924} /* (7, 20, 3) {real, imag} */,
  {32'h424bf022, 32'h4169eaf1} /* (7, 20, 2) {real, imag} */,
  {32'hc1679247, 32'hc20c3ba4} /* (7, 20, 1) {real, imag} */,
  {32'h41bd79a6, 32'h41c422de} /* (7, 20, 0) {real, imag} */,
  {32'h41414b46, 32'hc20c11d3} /* (7, 19, 31) {real, imag} */,
  {32'h429642f4, 32'hc1962253} /* (7, 19, 30) {real, imag} */,
  {32'hc196a22b, 32'h41eaf3fb} /* (7, 19, 29) {real, imag} */,
  {32'hc129950f, 32'h41f39df1} /* (7, 19, 28) {real, imag} */,
  {32'hc108efcd, 32'hc119acbe} /* (7, 19, 27) {real, imag} */,
  {32'hc1308444, 32'hc123ae5a} /* (7, 19, 26) {real, imag} */,
  {32'hc205acbb, 32'h428d99c3} /* (7, 19, 25) {real, imag} */,
  {32'hbfb6c768, 32'hc0747f04} /* (7, 19, 24) {real, imag} */,
  {32'h41740484, 32'h4146f3b4} /* (7, 19, 23) {real, imag} */,
  {32'h41b9ca15, 32'h417ec4a2} /* (7, 19, 22) {real, imag} */,
  {32'hc0f638f9, 32'hc0867e48} /* (7, 19, 21) {real, imag} */,
  {32'hc02ad348, 32'hc12bbe82} /* (7, 19, 20) {real, imag} */,
  {32'hc0281d6f, 32'h3fa205e0} /* (7, 19, 19) {real, imag} */,
  {32'hc10b8159, 32'h3f2b8a80} /* (7, 19, 18) {real, imag} */,
  {32'hc0f5daaa, 32'h40f87738} /* (7, 19, 17) {real, imag} */,
  {32'h408acda9, 32'hc1418a22} /* (7, 19, 16) {real, imag} */,
  {32'hbf2f4a20, 32'hc1348e84} /* (7, 19, 15) {real, imag} */,
  {32'h3f6c77d0, 32'h3f8fc6a0} /* (7, 19, 14) {real, imag} */,
  {32'hc014c6c1, 32'h413b1b70} /* (7, 19, 13) {real, imag} */,
  {32'h42235bdc, 32'h3f812cec} /* (7, 19, 12) {real, imag} */,
  {32'h416520de, 32'h417e570c} /* (7, 19, 11) {real, imag} */,
  {32'h40aa2224, 32'h40b500dc} /* (7, 19, 10) {real, imag} */,
  {32'h402fd160, 32'hc09417f0} /* (7, 19, 9) {real, imag} */,
  {32'hc1303685, 32'hc0e322b8} /* (7, 19, 8) {real, imag} */,
  {32'h40cf8030, 32'h40d65270} /* (7, 19, 7) {real, imag} */,
  {32'h41050300, 32'h4204e286} /* (7, 19, 6) {real, imag} */,
  {32'hc1933174, 32'hc1061dc2} /* (7, 19, 5) {real, imag} */,
  {32'hc05f7d84, 32'h411b5e6e} /* (7, 19, 4) {real, imag} */,
  {32'hc19edd5b, 32'h41f3db93} /* (7, 19, 3) {real, imag} */,
  {32'h418841e6, 32'hc25ec246} /* (7, 19, 2) {real, imag} */,
  {32'h41bcdb89, 32'hc07735d0} /* (7, 19, 1) {real, imag} */,
  {32'h40d46383, 32'hc1022a6a} /* (7, 19, 0) {real, imag} */,
  {32'hc1af1ec9, 32'h41c0255a} /* (7, 18, 31) {real, imag} */,
  {32'hc22ae0da, 32'hc0f35afc} /* (7, 18, 30) {real, imag} */,
  {32'h41598294, 32'h41c68324} /* (7, 18, 29) {real, imag} */,
  {32'h41a947b6, 32'h419c2932} /* (7, 18, 28) {real, imag} */,
  {32'hc23faaf0, 32'h425a1ba8} /* (7, 18, 27) {real, imag} */,
  {32'hc1ffdc58, 32'hc018a818} /* (7, 18, 26) {real, imag} */,
  {32'h40c4a63d, 32'hbdf38d00} /* (7, 18, 25) {real, imag} */,
  {32'hc05d6616, 32'h41d576b0} /* (7, 18, 24) {real, imag} */,
  {32'hc10f17d4, 32'h4121df35} /* (7, 18, 23) {real, imag} */,
  {32'hbe9415a0, 32'hc2062254} /* (7, 18, 22) {real, imag} */,
  {32'h40c2c2f8, 32'h40bd9220} /* (7, 18, 21) {real, imag} */,
  {32'h3fe42df8, 32'hc047d40e} /* (7, 18, 20) {real, imag} */,
  {32'h40f81326, 32'hc0d7296e} /* (7, 18, 19) {real, imag} */,
  {32'h3f528d40, 32'h3fa7533e} /* (7, 18, 18) {real, imag} */,
  {32'hbfb434dc, 32'h40be55f3} /* (7, 18, 17) {real, imag} */,
  {32'hc0ac5870, 32'h4096e536} /* (7, 18, 16) {real, imag} */,
  {32'hc11c4bc4, 32'hc00a1302} /* (7, 18, 15) {real, imag} */,
  {32'h4197a04f, 32'h401e2b37} /* (7, 18, 14) {real, imag} */,
  {32'h4127e961, 32'hc0113914} /* (7, 18, 13) {real, imag} */,
  {32'h4126917d, 32'h40d7f5bb} /* (7, 18, 12) {real, imag} */,
  {32'h413b3802, 32'hc0554970} /* (7, 18, 11) {real, imag} */,
  {32'h412a14a3, 32'h411b51be} /* (7, 18, 10) {real, imag} */,
  {32'h41b7fda4, 32'hc0a65fb2} /* (7, 18, 9) {real, imag} */,
  {32'h4195979c, 32'h41b77cc4} /* (7, 18, 8) {real, imag} */,
  {32'h40295806, 32'h422278bc} /* (7, 18, 7) {real, imag} */,
  {32'hc1652818, 32'hc1b1cde7} /* (7, 18, 6) {real, imag} */,
  {32'hc025a000, 32'h405dddc0} /* (7, 18, 5) {real, imag} */,
  {32'hc1fb1faa, 32'hc1a8577a} /* (7, 18, 4) {real, imag} */,
  {32'hc22bc885, 32'hc0ab8bb2} /* (7, 18, 3) {real, imag} */,
  {32'h4102e660, 32'h41bb8cc6} /* (7, 18, 2) {real, imag} */,
  {32'hc18209a1, 32'h4108090b} /* (7, 18, 1) {real, imag} */,
  {32'h4202ef90, 32'h41510d35} /* (7, 18, 0) {real, imag} */,
  {32'h410b9d8d, 32'hc167df12} /* (7, 17, 31) {real, imag} */,
  {32'h404d5714, 32'hc043d5d0} /* (7, 17, 30) {real, imag} */,
  {32'hc149b631, 32'h40c9ff78} /* (7, 17, 29) {real, imag} */,
  {32'h40a6571c, 32'h413fc3ea} /* (7, 17, 28) {real, imag} */,
  {32'h408bfabd, 32'h3ff5de14} /* (7, 17, 27) {real, imag} */,
  {32'h41d63e51, 32'h41b6a2bf} /* (7, 17, 26) {real, imag} */,
  {32'h407a2283, 32'hc18f0d40} /* (7, 17, 25) {real, imag} */,
  {32'h412cec1e, 32'hc1be9519} /* (7, 17, 24) {real, imag} */,
  {32'hc0910012, 32'hc09c610a} /* (7, 17, 23) {real, imag} */,
  {32'hc0d832c7, 32'hc117d63e} /* (7, 17, 22) {real, imag} */,
  {32'hc1babd79, 32'hbdf79dc0} /* (7, 17, 21) {real, imag} */,
  {32'h4085c93e, 32'h404d0cc2} /* (7, 17, 20) {real, imag} */,
  {32'hc0ef5cb4, 32'h411d6c8c} /* (7, 17, 19) {real, imag} */,
  {32'h40d5e168, 32'h3e949dc0} /* (7, 17, 18) {real, imag} */,
  {32'hc02da927, 32'h4084df4a} /* (7, 17, 17) {real, imag} */,
  {32'h40df8410, 32'hc002c896} /* (7, 17, 16) {real, imag} */,
  {32'h40d6d114, 32'h4115b193} /* (7, 17, 15) {real, imag} */,
  {32'h40ac3c6a, 32'h4156353e} /* (7, 17, 14) {real, imag} */,
  {32'h418b1ba8, 32'hc11c67d6} /* (7, 17, 13) {real, imag} */,
  {32'hc0a18cce, 32'hc0447582} /* (7, 17, 12) {real, imag} */,
  {32'h3fdbc7d0, 32'hc10f9574} /* (7, 17, 11) {real, imag} */,
  {32'h3facade4, 32'h4092fc3b} /* (7, 17, 10) {real, imag} */,
  {32'hc0d204d6, 32'h41a1095c} /* (7, 17, 9) {real, imag} */,
  {32'hc0909acf, 32'h41241016} /* (7, 17, 8) {real, imag} */,
  {32'hc08521a4, 32'hc0dcee66} /* (7, 17, 7) {real, imag} */,
  {32'hc2041c38, 32'h41d95f1d} /* (7, 17, 6) {real, imag} */,
  {32'hc15b83e6, 32'h3ff4229c} /* (7, 17, 5) {real, imag} */,
  {32'hc159ef72, 32'hc0a165dc} /* (7, 17, 4) {real, imag} */,
  {32'h414ed295, 32'hc11240aa} /* (7, 17, 3) {real, imag} */,
  {32'h41374eaa, 32'hc2300c54} /* (7, 17, 2) {real, imag} */,
  {32'hbbe05800, 32'h4190e75f} /* (7, 17, 1) {real, imag} */,
  {32'hc257425c, 32'h416b1de2} /* (7, 17, 0) {real, imag} */,
  {32'h41c0646b, 32'h4197ea6d} /* (7, 16, 31) {real, imag} */,
  {32'hc1d802f9, 32'hc1c4a0c9} /* (7, 16, 30) {real, imag} */,
  {32'h41e0bd04, 32'hc196f108} /* (7, 16, 29) {real, imag} */,
  {32'h4230059c, 32'h3edaa3f0} /* (7, 16, 28) {real, imag} */,
  {32'hc123cb31, 32'hbf1ef800} /* (7, 16, 27) {real, imag} */,
  {32'hc1db20f8, 32'hc18308b9} /* (7, 16, 26) {real, imag} */,
  {32'h4106ceca, 32'hc12d097d} /* (7, 16, 25) {real, imag} */,
  {32'h41652113, 32'h4020a5da} /* (7, 16, 24) {real, imag} */,
  {32'hc0412746, 32'hc0be53b2} /* (7, 16, 23) {real, imag} */,
  {32'h40ad1108, 32'h4055b618} /* (7, 16, 22) {real, imag} */,
  {32'h40d8de7d, 32'h41031862} /* (7, 16, 21) {real, imag} */,
  {32'hc119c612, 32'hc0cf9697} /* (7, 16, 20) {real, imag} */,
  {32'h40d1ecb1, 32'hc14200c5} /* (7, 16, 19) {real, imag} */,
  {32'hc0b22a11, 32'hc0d0947c} /* (7, 16, 18) {real, imag} */,
  {32'hc1033058, 32'h3fc63230} /* (7, 16, 17) {real, imag} */,
  {32'hbfc845e4, 32'hc081be89} /* (7, 16, 16) {real, imag} */,
  {32'h4021af00, 32'hbf5a0760} /* (7, 16, 15) {real, imag} */,
  {32'hc01ffe86, 32'hc08abb2a} /* (7, 16, 14) {real, imag} */,
  {32'h3ec79a50, 32'hc1082e0f} /* (7, 16, 13) {real, imag} */,
  {32'h3fd67760, 32'h3fb69a2c} /* (7, 16, 12) {real, imag} */,
  {32'hc0974d89, 32'h417db782} /* (7, 16, 11) {real, imag} */,
  {32'hc10c9cfb, 32'hc19e4024} /* (7, 16, 10) {real, imag} */,
  {32'h3fce3244, 32'h41b60bca} /* (7, 16, 9) {real, imag} */,
  {32'h400e2e1c, 32'h418bdcbf} /* (7, 16, 8) {real, imag} */,
  {32'hc1f0ae1f, 32'h3dbca480} /* (7, 16, 7) {real, imag} */,
  {32'h40cdb740, 32'h41056348} /* (7, 16, 6) {real, imag} */,
  {32'h412776c3, 32'h4158a8a7} /* (7, 16, 5) {real, imag} */,
  {32'hc03d91e0, 32'h4151143e} /* (7, 16, 4) {real, imag} */,
  {32'h40990980, 32'hc11c1b51} /* (7, 16, 3) {real, imag} */,
  {32'hc200bf14, 32'hbf9f3090} /* (7, 16, 2) {real, imag} */,
  {32'hc21d34ec, 32'hc1af7c39} /* (7, 16, 1) {real, imag} */,
  {32'h40eb4281, 32'h3f1f9838} /* (7, 16, 0) {real, imag} */,
  {32'h41915150, 32'hc17fdabe} /* (7, 15, 31) {real, imag} */,
  {32'hc1c9ded2, 32'hc13d252c} /* (7, 15, 30) {real, imag} */,
  {32'hc090f35c, 32'h410ddba0} /* (7, 15, 29) {real, imag} */,
  {32'hc0449e66, 32'h41f8d28b} /* (7, 15, 28) {real, imag} */,
  {32'h3d5688c0, 32'h41be419a} /* (7, 15, 27) {real, imag} */,
  {32'hbf21dc74, 32'hc1a70ee8} /* (7, 15, 26) {real, imag} */,
  {32'h4229e9ea, 32'h40f4fca4} /* (7, 15, 25) {real, imag} */,
  {32'hc14e0228, 32'h41729f5d} /* (7, 15, 24) {real, imag} */,
  {32'h4124468a, 32'hc13b7f93} /* (7, 15, 23) {real, imag} */,
  {32'h40061aec, 32'h41961dd2} /* (7, 15, 22) {real, imag} */,
  {32'h417e1bcc, 32'hc1029608} /* (7, 15, 21) {real, imag} */,
  {32'hc07498de, 32'h4061fe1b} /* (7, 15, 20) {real, imag} */,
  {32'h40614ad5, 32'h3ea097b8} /* (7, 15, 19) {real, imag} */,
  {32'h40e83486, 32'h403c7d07} /* (7, 15, 18) {real, imag} */,
  {32'h40a87fe4, 32'hbfd77380} /* (7, 15, 17) {real, imag} */,
  {32'hbeccff00, 32'h3fc665cc} /* (7, 15, 16) {real, imag} */,
  {32'h40087c21, 32'hc016b3b0} /* (7, 15, 15) {real, imag} */,
  {32'hc1066d24, 32'hbd0d35c0} /* (7, 15, 14) {real, imag} */,
  {32'h3fb5a56a, 32'h40c4de1e} /* (7, 15, 13) {real, imag} */,
  {32'hc0c21327, 32'hc059148d} /* (7, 15, 12) {real, imag} */,
  {32'hc0066470, 32'h4117aec8} /* (7, 15, 11) {real, imag} */,
  {32'hc19ba644, 32'hc0c1f99d} /* (7, 15, 10) {real, imag} */,
  {32'h41470582, 32'h41941c50} /* (7, 15, 9) {real, imag} */,
  {32'hbf16d348, 32'hc1b7b59a} /* (7, 15, 8) {real, imag} */,
  {32'h41cf5895, 32'h41d433f7} /* (7, 15, 7) {real, imag} */,
  {32'hbfa17af2, 32'h41195baa} /* (7, 15, 6) {real, imag} */,
  {32'h407edaab, 32'h41eb28f2} /* (7, 15, 5) {real, imag} */,
  {32'h40ffb521, 32'hc20a7c80} /* (7, 15, 4) {real, imag} */,
  {32'h41531d94, 32'hc0c61a7f} /* (7, 15, 3) {real, imag} */,
  {32'h41225b68, 32'hc1aae998} /* (7, 15, 2) {real, imag} */,
  {32'h4097b2e2, 32'hc24448a0} /* (7, 15, 1) {real, imag} */,
  {32'hc242537e, 32'hc1506eac} /* (7, 15, 0) {real, imag} */,
  {32'hc0a15f08, 32'hc0291268} /* (7, 14, 31) {real, imag} */,
  {32'h40e75274, 32'h417f58d4} /* (7, 14, 30) {real, imag} */,
  {32'h41d8efae, 32'h419096ec} /* (7, 14, 29) {real, imag} */,
  {32'hc123bc98, 32'hc1e66a87} /* (7, 14, 28) {real, imag} */,
  {32'h41ebe758, 32'hc2690348} /* (7, 14, 27) {real, imag} */,
  {32'hc2203bb6, 32'h418f6946} /* (7, 14, 26) {real, imag} */,
  {32'h41a18061, 32'hc1a78726} /* (7, 14, 25) {real, imag} */,
  {32'hc08f6c55, 32'h4189893a} /* (7, 14, 24) {real, imag} */,
  {32'hc074d97a, 32'h40a73736} /* (7, 14, 23) {real, imag} */,
  {32'hc024dd30, 32'hc14cc514} /* (7, 14, 22) {real, imag} */,
  {32'hc0e748ef, 32'h414c7fb7} /* (7, 14, 21) {real, imag} */,
  {32'h4031a9e2, 32'hc103c4b3} /* (7, 14, 20) {real, imag} */,
  {32'h406a78de, 32'hc028b758} /* (7, 14, 19) {real, imag} */,
  {32'h4114781e, 32'h4071f0cc} /* (7, 14, 18) {real, imag} */,
  {32'h411c646d, 32'hbe1b2330} /* (7, 14, 17) {real, imag} */,
  {32'h404f32a8, 32'h3fc312be} /* (7, 14, 16) {real, imag} */,
  {32'hbf836628, 32'hc0d076fa} /* (7, 14, 15) {real, imag} */,
  {32'hc030ff27, 32'h40896d3e} /* (7, 14, 14) {real, imag} */,
  {32'hc0e1b57b, 32'h40cc6c00} /* (7, 14, 13) {real, imag} */,
  {32'h415595bc, 32'h40ae2c18} /* (7, 14, 12) {real, imag} */,
  {32'h409561fd, 32'hc0a8ddbe} /* (7, 14, 11) {real, imag} */,
  {32'h413a9d48, 32'hc146375a} /* (7, 14, 10) {real, imag} */,
  {32'hc0c08bb3, 32'hc13fb15d} /* (7, 14, 9) {real, imag} */,
  {32'hc151ada6, 32'hc08ab3ce} /* (7, 14, 8) {real, imag} */,
  {32'h4208560c, 32'hc10016d6} /* (7, 14, 7) {real, imag} */,
  {32'h42385d2a, 32'hc19c2af6} /* (7, 14, 6) {real, imag} */,
  {32'h403fcb94, 32'h409d404c} /* (7, 14, 5) {real, imag} */,
  {32'hc08d8e1d, 32'h41674fb2} /* (7, 14, 4) {real, imag} */,
  {32'h417bb0b4, 32'h404320c8} /* (7, 14, 3) {real, imag} */,
  {32'hc132fd1e, 32'h41ffebd2} /* (7, 14, 2) {real, imag} */,
  {32'hc22e08ed, 32'h4180c167} /* (7, 14, 1) {real, imag} */,
  {32'hc18343da, 32'h3fae7c96} /* (7, 14, 0) {real, imag} */,
  {32'hc058fa28, 32'h40f45ea1} /* (7, 13, 31) {real, imag} */,
  {32'h419b3421, 32'h41597868} /* (7, 13, 30) {real, imag} */,
  {32'hc239f36f, 32'hc22490c1} /* (7, 13, 29) {real, imag} */,
  {32'hc1f28e8c, 32'hc1902c30} /* (7, 13, 28) {real, imag} */,
  {32'h4212bdee, 32'h40dddebe} /* (7, 13, 27) {real, imag} */,
  {32'hc1a5f45c, 32'hc1696172} /* (7, 13, 26) {real, imag} */,
  {32'hc0df32f4, 32'h4033a518} /* (7, 13, 25) {real, imag} */,
  {32'h41f14d17, 32'hbf8d61e8} /* (7, 13, 24) {real, imag} */,
  {32'h3ebbd510, 32'h4121c649} /* (7, 13, 23) {real, imag} */,
  {32'h40b32e5c, 32'h415f6ea4} /* (7, 13, 22) {real, imag} */,
  {32'h400eb9ce, 32'hc198cc38} /* (7, 13, 21) {real, imag} */,
  {32'hc0f56f70, 32'h41aa9e37} /* (7, 13, 20) {real, imag} */,
  {32'hbf968858, 32'hc12be53f} /* (7, 13, 19) {real, imag} */,
  {32'hbfd237c8, 32'h418ec0e0} /* (7, 13, 18) {real, imag} */,
  {32'hc08e18ae, 32'h3f1f35e0} /* (7, 13, 17) {real, imag} */,
  {32'h416f8d12, 32'h404e5450} /* (7, 13, 16) {real, imag} */,
  {32'h3f175e30, 32'h41990c9d} /* (7, 13, 15) {real, imag} */,
  {32'hc11a9baf, 32'hc1840ce2} /* (7, 13, 14) {real, imag} */,
  {32'h410f7879, 32'hc133a649} /* (7, 13, 13) {real, imag} */,
  {32'h40a5b1f4, 32'h40c90ef1} /* (7, 13, 12) {real, imag} */,
  {32'h418b5156, 32'h4084f2a6} /* (7, 13, 11) {real, imag} */,
  {32'h412961e4, 32'h4130c468} /* (7, 13, 10) {real, imag} */,
  {32'h40a60f57, 32'h41d48ac8} /* (7, 13, 9) {real, imag} */,
  {32'hc112860a, 32'hbf94e868} /* (7, 13, 8) {real, imag} */,
  {32'hc1da2e8d, 32'h419a3778} /* (7, 13, 7) {real, imag} */,
  {32'hc1654d40, 32'hc2898520} /* (7, 13, 6) {real, imag} */,
  {32'h4191bd6d, 32'hbf743810} /* (7, 13, 5) {real, imag} */,
  {32'hc0f9cf4e, 32'h41ac378a} /* (7, 13, 4) {real, imag} */,
  {32'h3f2571c0, 32'hc0b210a8} /* (7, 13, 3) {real, imag} */,
  {32'h41a223df, 32'h411bd6d4} /* (7, 13, 2) {real, imag} */,
  {32'h42519686, 32'hc132c424} /* (7, 13, 1) {real, imag} */,
  {32'hc1f70753, 32'hc22c9a11} /* (7, 13, 0) {real, imag} */,
  {32'h406347d1, 32'hc20a4c24} /* (7, 12, 31) {real, imag} */,
  {32'hc12b2f51, 32'hc1a7233b} /* (7, 12, 30) {real, imag} */,
  {32'hc1350c9f, 32'h42338304} /* (7, 12, 29) {real, imag} */,
  {32'hbfa2dde8, 32'hc272c9d6} /* (7, 12, 28) {real, imag} */,
  {32'hc1a679fc, 32'h41a6285d} /* (7, 12, 27) {real, imag} */,
  {32'hc02be621, 32'hc29011e6} /* (7, 12, 26) {real, imag} */,
  {32'hc16921ab, 32'hc1aeab3b} /* (7, 12, 25) {real, imag} */,
  {32'hc1bf43fa, 32'h41a3e45f} /* (7, 12, 24) {real, imag} */,
  {32'h41c31cfa, 32'h3f096b40} /* (7, 12, 23) {real, imag} */,
  {32'h412208a8, 32'h40d65558} /* (7, 12, 22) {real, imag} */,
  {32'h41bb9888, 32'h422928ac} /* (7, 12, 21) {real, imag} */,
  {32'h4023482c, 32'hc0c1880c} /* (7, 12, 20) {real, imag} */,
  {32'h41b3a38a, 32'hc13a431e} /* (7, 12, 19) {real, imag} */,
  {32'h40b8b38f, 32'hc1504a16} /* (7, 12, 18) {real, imag} */,
  {32'hc11f7176, 32'hc1724445} /* (7, 12, 17) {real, imag} */,
  {32'hc088c7c9, 32'hc0b29969} /* (7, 12, 16) {real, imag} */,
  {32'h4038baa7, 32'hc11554b3} /* (7, 12, 15) {real, imag} */,
  {32'hc13a5c22, 32'hc10b8b6a} /* (7, 12, 14) {real, imag} */,
  {32'h40c4423a, 32'hc0ec548c} /* (7, 12, 13) {real, imag} */,
  {32'hc0ad03e7, 32'h415363c6} /* (7, 12, 12) {real, imag} */,
  {32'hbf2c3e30, 32'h40fe3314} /* (7, 12, 11) {real, imag} */,
  {32'hc18737f2, 32'h41247dba} /* (7, 12, 10) {real, imag} */,
  {32'h422341af, 32'h41ca6a0e} /* (7, 12, 9) {real, imag} */,
  {32'h408e0880, 32'hc253d7d0} /* (7, 12, 8) {real, imag} */,
  {32'hc1f558c6, 32'hc176552a} /* (7, 12, 7) {real, imag} */,
  {32'h403d907f, 32'hc106ec94} /* (7, 12, 6) {real, imag} */,
  {32'h424619f2, 32'h41f3df9d} /* (7, 12, 5) {real, imag} */,
  {32'hc1477f41, 32'hc0fa4344} /* (7, 12, 4) {real, imag} */,
  {32'h4097e842, 32'h409dd7a4} /* (7, 12, 3) {real, imag} */,
  {32'hc18685e2, 32'hc13f578e} /* (7, 12, 2) {real, imag} */,
  {32'hc132c174, 32'h41f35055} /* (7, 12, 1) {real, imag} */,
  {32'hc08d5fa9, 32'hc182a865} /* (7, 12, 0) {real, imag} */,
  {32'hc2106d0f, 32'h40973178} /* (7, 11, 31) {real, imag} */,
  {32'hc225b693, 32'hc2563358} /* (7, 11, 30) {real, imag} */,
  {32'hc253a9bc, 32'h4206cdd6} /* (7, 11, 29) {real, imag} */,
  {32'hc08ab05a, 32'h413c0940} /* (7, 11, 28) {real, imag} */,
  {32'h427facfe, 32'h428678a0} /* (7, 11, 27) {real, imag} */,
  {32'hc00d2d20, 32'hc1a22810} /* (7, 11, 26) {real, imag} */,
  {32'h41e34c9e, 32'hc2073c0e} /* (7, 11, 25) {real, imag} */,
  {32'hc0c15564, 32'hc2161ba8} /* (7, 11, 24) {real, imag} */,
  {32'hc15cbff7, 32'hc26039e0} /* (7, 11, 23) {real, imag} */,
  {32'h4149d95c, 32'hc0a23d40} /* (7, 11, 22) {real, imag} */,
  {32'h40ce0f8a, 32'hc00ce7ec} /* (7, 11, 21) {real, imag} */,
  {32'h408cbe81, 32'h419eb756} /* (7, 11, 20) {real, imag} */,
  {32'hc11c3938, 32'h41787e07} /* (7, 11, 19) {real, imag} */,
  {32'hc0d59bbe, 32'hc12a0768} /* (7, 11, 18) {real, imag} */,
  {32'hbf1507f0, 32'hbfd16780} /* (7, 11, 17) {real, imag} */,
  {32'h41535fb0, 32'hc1197b58} /* (7, 11, 16) {real, imag} */,
  {32'hc0a36d12, 32'h4183f6ac} /* (7, 11, 15) {real, imag} */,
  {32'h41ac02e0, 32'hbf860d24} /* (7, 11, 14) {real, imag} */,
  {32'h414929c4, 32'hc20758b6} /* (7, 11, 13) {real, imag} */,
  {32'h3ff9418c, 32'hc143cfbc} /* (7, 11, 12) {real, imag} */,
  {32'hc18af38e, 32'hc0e1466e} /* (7, 11, 11) {real, imag} */,
  {32'hc20a479b, 32'hc121e14a} /* (7, 11, 10) {real, imag} */,
  {32'hc20aa1cc, 32'h41653036} /* (7, 11, 9) {real, imag} */,
  {32'h41353d8a, 32'hbe8c5340} /* (7, 11, 8) {real, imag} */,
  {32'h42773daf, 32'h4105a6a2} /* (7, 11, 7) {real, imag} */,
  {32'hc21decbc, 32'h42165c94} /* (7, 11, 6) {real, imag} */,
  {32'hc0fe1ec0, 32'hc1985eb8} /* (7, 11, 5) {real, imag} */,
  {32'hc1b77c58, 32'hc13f2d26} /* (7, 11, 4) {real, imag} */,
  {32'hc1ae79d7, 32'h420513d0} /* (7, 11, 3) {real, imag} */,
  {32'h42832628, 32'hc203d6d8} /* (7, 11, 2) {real, imag} */,
  {32'hc29fe0a6, 32'hc250b715} /* (7, 11, 1) {real, imag} */,
  {32'hc1997b94, 32'hc1ca784a} /* (7, 11, 0) {real, imag} */,
  {32'h40a5aee5, 32'hc2021231} /* (7, 10, 31) {real, imag} */,
  {32'hc20bc30e, 32'hc28b9e77} /* (7, 10, 30) {real, imag} */,
  {32'hc1f677c4, 32'h42781b2c} /* (7, 10, 29) {real, imag} */,
  {32'hc2864941, 32'hc17d2920} /* (7, 10, 28) {real, imag} */,
  {32'h415a5624, 32'h422088ea} /* (7, 10, 27) {real, imag} */,
  {32'h41738338, 32'h4286653c} /* (7, 10, 26) {real, imag} */,
  {32'h420644bb, 32'hc243903a} /* (7, 10, 25) {real, imag} */,
  {32'h41ba5a0b, 32'h420baa91} /* (7, 10, 24) {real, imag} */,
  {32'hc12d5906, 32'hc22fd236} /* (7, 10, 23) {real, imag} */,
  {32'h421f5a86, 32'hc18e4fb4} /* (7, 10, 22) {real, imag} */,
  {32'hc1fda5f8, 32'h41a87907} /* (7, 10, 21) {real, imag} */,
  {32'hc1d8c330, 32'h40d941ee} /* (7, 10, 20) {real, imag} */,
  {32'hc21168a4, 32'h410147b9} /* (7, 10, 19) {real, imag} */,
  {32'h40822a82, 32'hc03eb824} /* (7, 10, 18) {real, imag} */,
  {32'hbef57d20, 32'hc1a23cb2} /* (7, 10, 17) {real, imag} */,
  {32'hbfc3f680, 32'hc010a4e8} /* (7, 10, 16) {real, imag} */,
  {32'hc112e8f6, 32'h408d8d1a} /* (7, 10, 15) {real, imag} */,
  {32'hc04a10dc, 32'hc12ec5b1} /* (7, 10, 14) {real, imag} */,
  {32'hc02d47d8, 32'h417400ed} /* (7, 10, 13) {real, imag} */,
  {32'h41e2f00a, 32'hc14cc1ab} /* (7, 10, 12) {real, imag} */,
  {32'hc0bddab8, 32'h401f5428} /* (7, 10, 11) {real, imag} */,
  {32'h40bdb44c, 32'hc1f397e8} /* (7, 10, 10) {real, imag} */,
  {32'hbfe71dac, 32'hc165e120} /* (7, 10, 9) {real, imag} */,
  {32'hc135ac8a, 32'h41a77e04} /* (7, 10, 8) {real, imag} */,
  {32'h41b7e89b, 32'h3e8e2200} /* (7, 10, 7) {real, imag} */,
  {32'hc1b66044, 32'h420a3632} /* (7, 10, 6) {real, imag} */,
  {32'hc1e6b2c4, 32'h41e7bd35} /* (7, 10, 5) {real, imag} */,
  {32'hc229186a, 32'hc11de6da} /* (7, 10, 4) {real, imag} */,
  {32'hc0f42ee6, 32'hc28b5120} /* (7, 10, 3) {real, imag} */,
  {32'h425648a0, 32'h42721f69} /* (7, 10, 2) {real, imag} */,
  {32'h41464c86, 32'hc1d1b83a} /* (7, 10, 1) {real, imag} */,
  {32'h4209ecc9, 32'h40d3563c} /* (7, 10, 0) {real, imag} */,
  {32'h41b07eb6, 32'hc2238d28} /* (7, 9, 31) {real, imag} */,
  {32'h420ebf6e, 32'h4137fa26} /* (7, 9, 30) {real, imag} */,
  {32'hc191d520, 32'h41eb6f4f} /* (7, 9, 29) {real, imag} */,
  {32'h424df3b6, 32'hc0c4ce78} /* (7, 9, 28) {real, imag} */,
  {32'hc1a39764, 32'hc22f0e74} /* (7, 9, 27) {real, imag} */,
  {32'hc204cbb8, 32'h40ebb6f8} /* (7, 9, 26) {real, imag} */,
  {32'h42919728, 32'h41668744} /* (7, 9, 25) {real, imag} */,
  {32'hbdc69700, 32'hc201620a} /* (7, 9, 24) {real, imag} */,
  {32'h4192d288, 32'hc0fd97f8} /* (7, 9, 23) {real, imag} */,
  {32'h422ee60a, 32'h420556fa} /* (7, 9, 22) {real, imag} */,
  {32'hc21fadc1, 32'h41628df9} /* (7, 9, 21) {real, imag} */,
  {32'hc14b462b, 32'h408bab3a} /* (7, 9, 20) {real, imag} */,
  {32'h41902bca, 32'hc18e58fb} /* (7, 9, 19) {real, imag} */,
  {32'h4108f466, 32'hc1958cdd} /* (7, 9, 18) {real, imag} */,
  {32'hc1109bfd, 32'h4191198c} /* (7, 9, 17) {real, imag} */,
  {32'h4090844e, 32'hc14320b6} /* (7, 9, 16) {real, imag} */,
  {32'h4088190a, 32'hc1213ed9} /* (7, 9, 15) {real, imag} */,
  {32'h40a1e674, 32'h4140654a} /* (7, 9, 14) {real, imag} */,
  {32'h41b48e4a, 32'hc0a6e8f7} /* (7, 9, 13) {real, imag} */,
  {32'h41561d57, 32'h409a434a} /* (7, 9, 12) {real, imag} */,
  {32'hc1ddeb6e, 32'hc14b1e71} /* (7, 9, 11) {real, imag} */,
  {32'h421fa698, 32'h4248883c} /* (7, 9, 10) {real, imag} */,
  {32'hc0f99b0e, 32'hc2732a5f} /* (7, 9, 9) {real, imag} */,
  {32'h4203f548, 32'h41ae53c3} /* (7, 9, 8) {real, imag} */,
  {32'hc22bc2da, 32'h42c96720} /* (7, 9, 7) {real, imag} */,
  {32'hc1dde8a4, 32'hc294ffb4} /* (7, 9, 6) {real, imag} */,
  {32'hc04abb94, 32'hc0de5dec} /* (7, 9, 5) {real, imag} */,
  {32'hc1bcd469, 32'h41db5a9e} /* (7, 9, 4) {real, imag} */,
  {32'h3fb493a8, 32'h41686ada} /* (7, 9, 3) {real, imag} */,
  {32'h4309ecae, 32'h410d9412} /* (7, 9, 2) {real, imag} */,
  {32'h421071f3, 32'h4206df18} /* (7, 9, 1) {real, imag} */,
  {32'hc1cc05fe, 32'h428e87bd} /* (7, 9, 0) {real, imag} */,
  {32'hc0d96468, 32'h41f39e8f} /* (7, 8, 31) {real, imag} */,
  {32'hc20e0fe0, 32'h41ad1850} /* (7, 8, 30) {real, imag} */,
  {32'h42c2a9c4, 32'hc0edf230} /* (7, 8, 29) {real, imag} */,
  {32'hc15d0036, 32'h42a4e5a2} /* (7, 8, 28) {real, imag} */,
  {32'h421e587a, 32'h428795e1} /* (7, 8, 27) {real, imag} */,
  {32'h41490317, 32'hc2b23c74} /* (7, 8, 26) {real, imag} */,
  {32'hc23c6546, 32'hc1195a2d} /* (7, 8, 25) {real, imag} */,
  {32'hc1e1205f, 32'h41679929} /* (7, 8, 24) {real, imag} */,
  {32'hc28dbcb1, 32'hc17e8498} /* (7, 8, 23) {real, imag} */,
  {32'hc1ccf904, 32'hc22194ce} /* (7, 8, 22) {real, imag} */,
  {32'hc1501102, 32'h404d86f8} /* (7, 8, 21) {real, imag} */,
  {32'h40c49170, 32'hc11e8159} /* (7, 8, 20) {real, imag} */,
  {32'h41a36af4, 32'h40bdb83a} /* (7, 8, 19) {real, imag} */,
  {32'hc0980da0, 32'hc11ef33e} /* (7, 8, 18) {real, imag} */,
  {32'hc1dab7a8, 32'h4091f1ac} /* (7, 8, 17) {real, imag} */,
  {32'hbf9ff068, 32'hc17f6078} /* (7, 8, 16) {real, imag} */,
  {32'hc0cbc1b2, 32'hc1dfff51} /* (7, 8, 15) {real, imag} */,
  {32'hc0bc2c00, 32'h4164a4ec} /* (7, 8, 14) {real, imag} */,
  {32'hc04ac420, 32'hc13944ad} /* (7, 8, 13) {real, imag} */,
  {32'hc2353cdf, 32'h40101984} /* (7, 8, 12) {real, imag} */,
  {32'h429716a8, 32'h40e6d094} /* (7, 8, 11) {real, imag} */,
  {32'h41bf8104, 32'hc209a6a6} /* (7, 8, 10) {real, imag} */,
  {32'h4270a90d, 32'h4251f2ac} /* (7, 8, 9) {real, imag} */,
  {32'h413b9776, 32'hc091299a} /* (7, 8, 8) {real, imag} */,
  {32'h42a4c1d5, 32'h414f3adb} /* (7, 8, 7) {real, imag} */,
  {32'h41fe6904, 32'h417803b0} /* (7, 8, 6) {real, imag} */,
  {32'hc2216e82, 32'h41cfe117} /* (7, 8, 5) {real, imag} */,
  {32'h427ae4b4, 32'h421683d8} /* (7, 8, 4) {real, imag} */,
  {32'hbee1ab80, 32'h40924bf0} /* (7, 8, 3) {real, imag} */,
  {32'hc1b16025, 32'hc26afe4a} /* (7, 8, 2) {real, imag} */,
  {32'hc26b92eb, 32'hc2939665} /* (7, 8, 1) {real, imag} */,
  {32'h41a40ae6, 32'h42d0a42f} /* (7, 8, 0) {real, imag} */,
  {32'h419f8a0f, 32'hc18baff2} /* (7, 7, 31) {real, imag} */,
  {32'h4241133b, 32'h42a99d5e} /* (7, 7, 30) {real, imag} */,
  {32'h4290d327, 32'h42a2cbdf} /* (7, 7, 29) {real, imag} */,
  {32'h41865250, 32'h419fd755} /* (7, 7, 28) {real, imag} */,
  {32'hc1d4d63f, 32'h41786768} /* (7, 7, 27) {real, imag} */,
  {32'hc260250e, 32'hbf9e5ab0} /* (7, 7, 26) {real, imag} */,
  {32'h40a086c0, 32'hc26dc29c} /* (7, 7, 25) {real, imag} */,
  {32'hc1169533, 32'hc10bb20e} /* (7, 7, 24) {real, imag} */,
  {32'h4109a35d, 32'h41dc2670} /* (7, 7, 23) {real, imag} */,
  {32'h421f2f5c, 32'hc1fc6e57} /* (7, 7, 22) {real, imag} */,
  {32'h41f25708, 32'h4238cf61} /* (7, 7, 21) {real, imag} */,
  {32'h42135472, 32'hc15cd62c} /* (7, 7, 20) {real, imag} */,
  {32'hc12127da, 32'hc0c90980} /* (7, 7, 19) {real, imag} */,
  {32'hc0730b3c, 32'h41dce655} /* (7, 7, 18) {real, imag} */,
  {32'h415651e9, 32'hc0ff13f0} /* (7, 7, 17) {real, imag} */,
  {32'h411b2104, 32'h3e2d2480} /* (7, 7, 16) {real, imag} */,
  {32'h416fd351, 32'h41844b7d} /* (7, 7, 15) {real, imag} */,
  {32'hbf9028a8, 32'hc136ab2a} /* (7, 7, 14) {real, imag} */,
  {32'h41b8cc51, 32'hc147207c} /* (7, 7, 13) {real, imag} */,
  {32'hc18d6ff6, 32'h40c42a1b} /* (7, 7, 12) {real, imag} */,
  {32'hbf820b48, 32'h415dde48} /* (7, 7, 11) {real, imag} */,
  {32'hc06f3960, 32'hc08f0e54} /* (7, 7, 10) {real, imag} */,
  {32'hc20bf601, 32'hc25cde86} /* (7, 7, 9) {real, imag} */,
  {32'h416b99c5, 32'hc2048056} /* (7, 7, 8) {real, imag} */,
  {32'h4239b460, 32'h3ffe3740} /* (7, 7, 7) {real, imag} */,
  {32'h406f2bc0, 32'h42517588} /* (7, 7, 6) {real, imag} */,
  {32'h412c1ada, 32'h42a2b879} /* (7, 7, 5) {real, imag} */,
  {32'hc1d655d2, 32'hc1cc4223} /* (7, 7, 4) {real, imag} */,
  {32'hc2a5015f, 32'h418069fc} /* (7, 7, 3) {real, imag} */,
  {32'h420c1205, 32'h421cf3ac} /* (7, 7, 2) {real, imag} */,
  {32'h427f4b9e, 32'hc1eed3ae} /* (7, 7, 1) {real, imag} */,
  {32'hc26c780b, 32'hc1ff7e4b} /* (7, 7, 0) {real, imag} */,
  {32'hc24d8314, 32'hc2552aee} /* (7, 6, 31) {real, imag} */,
  {32'h42eb1db2, 32'h41696b34} /* (7, 6, 30) {real, imag} */,
  {32'h417ac1a4, 32'h42af5495} /* (7, 6, 29) {real, imag} */,
  {32'h41333f76, 32'h422cba60} /* (7, 6, 28) {real, imag} */,
  {32'hc270be24, 32'h428fb517} /* (7, 6, 27) {real, imag} */,
  {32'hc228169c, 32'h3f3b9ad0} /* (7, 6, 26) {real, imag} */,
  {32'h428c2edb, 32'hc18c1e8c} /* (7, 6, 25) {real, imag} */,
  {32'hc1f40c7f, 32'h41a30c7a} /* (7, 6, 24) {real, imag} */,
  {32'h4233a1e8, 32'h3ec671c0} /* (7, 6, 23) {real, imag} */,
  {32'hc27f4c3c, 32'h41d438c8} /* (7, 6, 22) {real, imag} */,
  {32'h4229f85e, 32'h4245ca18} /* (7, 6, 21) {real, imag} */,
  {32'h4049a1e2, 32'hc1b2387c} /* (7, 6, 20) {real, imag} */,
  {32'hc1740330, 32'hc1f0bbb8} /* (7, 6, 19) {real, imag} */,
  {32'hc07f5098, 32'hc0ce5994} /* (7, 6, 18) {real, imag} */,
  {32'hc03f2688, 32'h41a5723f} /* (7, 6, 17) {real, imag} */,
  {32'h40906562, 32'hc1010908} /* (7, 6, 16) {real, imag} */,
  {32'h40c2a1bc, 32'h40cbe7e4} /* (7, 6, 15) {real, imag} */,
  {32'h41384b1a, 32'hc0b378dc} /* (7, 6, 14) {real, imag} */,
  {32'h40668f18, 32'h4239c0e8} /* (7, 6, 13) {real, imag} */,
  {32'h3e4336e0, 32'hc18abf6e} /* (7, 6, 12) {real, imag} */,
  {32'hbe469f00, 32'h42475580} /* (7, 6, 11) {real, imag} */,
  {32'h41694d62, 32'hc1287e03} /* (7, 6, 10) {real, imag} */,
  {32'h41d3dcf4, 32'hc24c4746} /* (7, 6, 9) {real, imag} */,
  {32'hc255f4c8, 32'h423d67af} /* (7, 6, 8) {real, imag} */,
  {32'hc16f5c30, 32'hc250142a} /* (7, 6, 7) {real, imag} */,
  {32'hc11be3b2, 32'hc1209d97} /* (7, 6, 6) {real, imag} */,
  {32'hc23ad454, 32'hc20b2df2} /* (7, 6, 5) {real, imag} */,
  {32'h4232be16, 32'h411eb7a4} /* (7, 6, 4) {real, imag} */,
  {32'hc0e85604, 32'hc1400248} /* (7, 6, 3) {real, imag} */,
  {32'hc2130494, 32'hc2acdcd0} /* (7, 6, 2) {real, imag} */,
  {32'h42e4fb1e, 32'h42518146} /* (7, 6, 1) {real, imag} */,
  {32'hc107f0f1, 32'hc1b4e87a} /* (7, 6, 0) {real, imag} */,
  {32'h422886c4, 32'h4214b73f} /* (7, 5, 31) {real, imag} */,
  {32'hc0b50ee8, 32'h43412296} /* (7, 5, 30) {real, imag} */,
  {32'h420ec3b9, 32'h414589c4} /* (7, 5, 29) {real, imag} */,
  {32'h41cda316, 32'hc246900c} /* (7, 5, 28) {real, imag} */,
  {32'h4302bb40, 32'hc29b068b} /* (7, 5, 27) {real, imag} */,
  {32'hc2bb0187, 32'h41882309} /* (7, 5, 26) {real, imag} */,
  {32'h4272f743, 32'h42f32c4c} /* (7, 5, 25) {real, imag} */,
  {32'hc09ce4dc, 32'hc1fc68d8} /* (7, 5, 24) {real, imag} */,
  {32'h428eddf4, 32'h42896408} /* (7, 5, 23) {real, imag} */,
  {32'h4158062f, 32'h40e599f8} /* (7, 5, 22) {real, imag} */,
  {32'hc211b5f2, 32'hc1895634} /* (7, 5, 21) {real, imag} */,
  {32'hc200db85, 32'hc1308654} /* (7, 5, 20) {real, imag} */,
  {32'hc285f885, 32'h411e6e5b} /* (7, 5, 19) {real, imag} */,
  {32'h42620042, 32'h41a895d4} /* (7, 5, 18) {real, imag} */,
  {32'h4049c6a0, 32'h416721e4} /* (7, 5, 17) {real, imag} */,
  {32'h41b24586, 32'h40333840} /* (7, 5, 16) {real, imag} */,
  {32'h41b023d6, 32'hc14f0be8} /* (7, 5, 15) {real, imag} */,
  {32'h4187ac8c, 32'h40b9ecd0} /* (7, 5, 14) {real, imag} */,
  {32'h418ada58, 32'hc1898e7a} /* (7, 5, 13) {real, imag} */,
  {32'h410d3fb4, 32'hc1ced78c} /* (7, 5, 12) {real, imag} */,
  {32'hbf78fe00, 32'hc23d919a} /* (7, 5, 11) {real, imag} */,
  {32'hc12d6317, 32'h42d46114} /* (7, 5, 10) {real, imag} */,
  {32'h4020e7d0, 32'h42910c2c} /* (7, 5, 9) {real, imag} */,
  {32'h418ed835, 32'h4220e866} /* (7, 5, 8) {real, imag} */,
  {32'h42806e24, 32'hc2987fd0} /* (7, 5, 7) {real, imag} */,
  {32'hc27e0bc2, 32'h41830c45} /* (7, 5, 6) {real, imag} */,
  {32'hc1c15832, 32'h4203d18a} /* (7, 5, 5) {real, imag} */,
  {32'h421b1c45, 32'h42524124} /* (7, 5, 4) {real, imag} */,
  {32'hc1e4439a, 32'hc2a45bb0} /* (7, 5, 3) {real, imag} */,
  {32'hc2a949ee, 32'h42a82804} /* (7, 5, 2) {real, imag} */,
  {32'hc257cfd4, 32'hc1c12c68} /* (7, 5, 1) {real, imag} */,
  {32'h42088cda, 32'hc32f2893} /* (7, 5, 0) {real, imag} */,
  {32'h423a873a, 32'hc252407e} /* (7, 4, 31) {real, imag} */,
  {32'h42bc43dc, 32'hc2f78532} /* (7, 4, 30) {real, imag} */,
  {32'hc1cbb34b, 32'hc28d1142} /* (7, 4, 29) {real, imag} */,
  {32'hc281663d, 32'h42b6e1fd} /* (7, 4, 28) {real, imag} */,
  {32'h42cfacde, 32'hc2a65582} /* (7, 4, 27) {real, imag} */,
  {32'hc22b3f4f, 32'h425f8920} /* (7, 4, 26) {real, imag} */,
  {32'h41bc0f8d, 32'h4245dfec} /* (7, 4, 25) {real, imag} */,
  {32'h428bc923, 32'h424f6af5} /* (7, 4, 24) {real, imag} */,
  {32'hbfb2c4d0, 32'h3ecb5b00} /* (7, 4, 23) {real, imag} */,
  {32'hc19e21d6, 32'h429b51f6} /* (7, 4, 22) {real, imag} */,
  {32'hc28f57b6, 32'hc21ecf2f} /* (7, 4, 21) {real, imag} */,
  {32'h41070858, 32'h40746d50} /* (7, 4, 20) {real, imag} */,
  {32'hc1ab9bbf, 32'hc030f5d0} /* (7, 4, 19) {real, imag} */,
  {32'hc16ee2ab, 32'h42598035} /* (7, 4, 18) {real, imag} */,
  {32'hc0830b72, 32'hc18f1e90} /* (7, 4, 17) {real, imag} */,
  {32'h40d56778, 32'h40edf990} /* (7, 4, 16) {real, imag} */,
  {32'h40af059e, 32'hbffd78b8} /* (7, 4, 15) {real, imag} */,
  {32'h40f4f8d6, 32'h42120ba5} /* (7, 4, 14) {real, imag} */,
  {32'hc284e363, 32'hc1824ace} /* (7, 4, 13) {real, imag} */,
  {32'h41c7de24, 32'hc203a2fd} /* (7, 4, 12) {real, imag} */,
  {32'h41b64fbc, 32'h424da62d} /* (7, 4, 11) {real, imag} */,
  {32'h40e2dc9a, 32'hc1ccdcca} /* (7, 4, 10) {real, imag} */,
  {32'hc21f7322, 32'hc24490d4} /* (7, 4, 9) {real, imag} */,
  {32'h4284a245, 32'h42809042} /* (7, 4, 8) {real, imag} */,
  {32'hc2a0453f, 32'hc20d4fa2} /* (7, 4, 7) {real, imag} */,
  {32'h4196a86e, 32'h426d9b96} /* (7, 4, 6) {real, imag} */,
  {32'h4205512d, 32'h4210005c} /* (7, 4, 5) {real, imag} */,
  {32'h43125308, 32'hbdf5f800} /* (7, 4, 4) {real, imag} */,
  {32'hc2a1a316, 32'h42adbab6} /* (7, 4, 3) {real, imag} */,
  {32'h42377488, 32'hc34348cd} /* (7, 4, 2) {real, imag} */,
  {32'hc1398d50, 32'h42845640} /* (7, 4, 1) {real, imag} */,
  {32'hc18193fa, 32'h42860847} /* (7, 4, 0) {real, imag} */,
  {32'hc3201888, 32'hc2f8eeee} /* (7, 3, 31) {real, imag} */,
  {32'h40b27b18, 32'h429ea427} /* (7, 3, 30) {real, imag} */,
  {32'hc05ba800, 32'h4329be72} /* (7, 3, 29) {real, imag} */,
  {32'hc151b128, 32'hc28d6148} /* (7, 3, 28) {real, imag} */,
  {32'h4048ad38, 32'hc24bc853} /* (7, 3, 27) {real, imag} */,
  {32'h42111a89, 32'hc2851798} /* (7, 3, 26) {real, imag} */,
  {32'h421a004b, 32'hc1ac9004} /* (7, 3, 25) {real, imag} */,
  {32'h423091da, 32'hc0f51d78} /* (7, 3, 24) {real, imag} */,
  {32'h41f59291, 32'h42ab50b3} /* (7, 3, 23) {real, imag} */,
  {32'hc16e62ae, 32'h421032db} /* (7, 3, 22) {real, imag} */,
  {32'hc0a66624, 32'hc1a67e48} /* (7, 3, 21) {real, imag} */,
  {32'h426d1722, 32'hc2b77543} /* (7, 3, 20) {real, imag} */,
  {32'hc136f168, 32'h4262535e} /* (7, 3, 19) {real, imag} */,
  {32'h417b285e, 32'hc129b086} /* (7, 3, 18) {real, imag} */,
  {32'hc126d720, 32'hc161a9ba} /* (7, 3, 17) {real, imag} */,
  {32'hc146bcb4, 32'hc10877e4} /* (7, 3, 16) {real, imag} */,
  {32'h418d29a0, 32'hc0be3104} /* (7, 3, 15) {real, imag} */,
  {32'hc29191ea, 32'hc1be09c5} /* (7, 3, 14) {real, imag} */,
  {32'hc0341bc0, 32'h40a1d470} /* (7, 3, 13) {real, imag} */,
  {32'h4194d8c8, 32'hc2444cd2} /* (7, 3, 12) {real, imag} */,
  {32'h4242b5d0, 32'hc0b7b212} /* (7, 3, 11) {real, imag} */,
  {32'h412e9182, 32'hc20e196f} /* (7, 3, 10) {real, imag} */,
  {32'h40fc1a6c, 32'hc2a45821} /* (7, 3, 9) {real, imag} */,
  {32'h410367c6, 32'h41d88aa6} /* (7, 3, 8) {real, imag} */,
  {32'hc2db5520, 32'h41721377} /* (7, 3, 7) {real, imag} */,
  {32'hc28e97ee, 32'h428995a0} /* (7, 3, 6) {real, imag} */,
  {32'hc27fd0fa, 32'hc2ded6f2} /* (7, 3, 5) {real, imag} */,
  {32'h42c9a06e, 32'hc05bfb30} /* (7, 3, 4) {real, imag} */,
  {32'h431b503a, 32'h40837770} /* (7, 3, 3) {real, imag} */,
  {32'h4224fc64, 32'hc22e8cd2} /* (7, 3, 2) {real, imag} */,
  {32'h42c4aa18, 32'h41b14728} /* (7, 3, 1) {real, imag} */,
  {32'h42d417a4, 32'h4143a364} /* (7, 3, 0) {real, imag} */,
  {32'hc2929622, 32'h4296d9d6} /* (7, 2, 31) {real, imag} */,
  {32'hc241b95e, 32'hc31b23dc} /* (7, 2, 30) {real, imag} */,
  {32'hc334bebd, 32'hc3105a04} /* (7, 2, 29) {real, imag} */,
  {32'h42d09552, 32'hc30b6f48} /* (7, 2, 28) {real, imag} */,
  {32'hc296a798, 32'h42507405} /* (7, 2, 27) {real, imag} */,
  {32'hc20e291c, 32'h41a8fb68} /* (7, 2, 26) {real, imag} */,
  {32'h410ec2df, 32'h42a3d740} /* (7, 2, 25) {real, imag} */,
  {32'h420d7d67, 32'hc2e409c4} /* (7, 2, 24) {real, imag} */,
  {32'h421dada7, 32'h416759f6} /* (7, 2, 23) {real, imag} */,
  {32'hc213f83b, 32'h41a25ab4} /* (7, 2, 22) {real, imag} */,
  {32'hc275f3da, 32'hc12258c2} /* (7, 2, 21) {real, imag} */,
  {32'h420adb56, 32'h41595080} /* (7, 2, 20) {real, imag} */,
  {32'hc0d34908, 32'h418e99e2} /* (7, 2, 19) {real, imag} */,
  {32'h40b57d54, 32'hc1df3f04} /* (7, 2, 18) {real, imag} */,
  {32'h4153272c, 32'h4259f6e0} /* (7, 2, 17) {real, imag} */,
  {32'h40ce8078, 32'hc1a397d6} /* (7, 2, 16) {real, imag} */,
  {32'hbfa204a0, 32'h406c4238} /* (7, 2, 15) {real, imag} */,
  {32'h41cfccf3, 32'h40a22870} /* (7, 2, 14) {real, imag} */,
  {32'hc0cdc688, 32'h4109f74c} /* (7, 2, 13) {real, imag} */,
  {32'h4200f1e0, 32'h41393ab8} /* (7, 2, 12) {real, imag} */,
  {32'hc2bf9607, 32'hc220dc4c} /* (7, 2, 11) {real, imag} */,
  {32'hc2958478, 32'hbf9ee308} /* (7, 2, 10) {real, imag} */,
  {32'h42b8c266, 32'h40ce0ed4} /* (7, 2, 9) {real, imag} */,
  {32'h4202cffd, 32'h3fb76c80} /* (7, 2, 8) {real, imag} */,
  {32'h41e3c286, 32'hc031fd80} /* (7, 2, 7) {real, imag} */,
  {32'hc2343a4c, 32'h420ce592} /* (7, 2, 6) {real, imag} */,
  {32'h42c5d0da, 32'hc227de53} /* (7, 2, 5) {real, imag} */,
  {32'h421fc913, 32'hc1e1c354} /* (7, 2, 4) {real, imag} */,
  {32'h42cd81c2, 32'hc100a6a8} /* (7, 2, 3) {real, imag} */,
  {32'hc2c99cb9, 32'hc28b8c5b} /* (7, 2, 2) {real, imag} */,
  {32'hc1bb9d90, 32'h4237db81} /* (7, 2, 1) {real, imag} */,
  {32'hc1ce5884, 32'h4296d556} /* (7, 2, 0) {real, imag} */,
  {32'h4034e640, 32'hc33ecf0a} /* (7, 1, 31) {real, imag} */,
  {32'hc31d11ac, 32'h42ea6605} /* (7, 1, 30) {real, imag} */,
  {32'h411ad04c, 32'h42547754} /* (7, 1, 29) {real, imag} */,
  {32'h42d027e4, 32'hc2071b6c} /* (7, 1, 28) {real, imag} */,
  {32'h42931f80, 32'h432b2d34} /* (7, 1, 27) {real, imag} */,
  {32'h41eb5192, 32'h41b31e20} /* (7, 1, 26) {real, imag} */,
  {32'h42407654, 32'h43062b76} /* (7, 1, 25) {real, imag} */,
  {32'h41a2d690, 32'hc23f3b32} /* (7, 1, 24) {real, imag} */,
  {32'h4219c5d6, 32'hc2e27a43} /* (7, 1, 23) {real, imag} */,
  {32'hc2ce2264, 32'h4200ba76} /* (7, 1, 22) {real, imag} */,
  {32'hc2220bea, 32'hc1fc9ccc} /* (7, 1, 21) {real, imag} */,
  {32'hc1f47c65, 32'h420c0adc} /* (7, 1, 20) {real, imag} */,
  {32'h41b77432, 32'hc222f05a} /* (7, 1, 19) {real, imag} */,
  {32'hc21dd2d8, 32'h4191527e} /* (7, 1, 18) {real, imag} */,
  {32'hc11750b0, 32'h41af309d} /* (7, 1, 17) {real, imag} */,
  {32'h41428859, 32'hc110be90} /* (7, 1, 16) {real, imag} */,
  {32'hc141eed4, 32'h415ea396} /* (7, 1, 15) {real, imag} */,
  {32'h402a5078, 32'hc1eea7ea} /* (7, 1, 14) {real, imag} */,
  {32'h41dab7ba, 32'h412684a7} /* (7, 1, 13) {real, imag} */,
  {32'h3f78e9a0, 32'h41ce10f1} /* (7, 1, 12) {real, imag} */,
  {32'hc1b01b7c, 32'hc274c4d6} /* (7, 1, 11) {real, imag} */,
  {32'hc29aed44, 32'hc1e7ce1c} /* (7, 1, 10) {real, imag} */,
  {32'h41483e92, 32'hc0025520} /* (7, 1, 9) {real, imag} */,
  {32'hc208bac0, 32'hc0f9aa44} /* (7, 1, 8) {real, imag} */,
  {32'h3f800a10, 32'h423c20ce} /* (7, 1, 7) {real, imag} */,
  {32'h42c3709e, 32'hc3353dff} /* (7, 1, 6) {real, imag} */,
  {32'hc1b061d8, 32'hc2117e2c} /* (7, 1, 5) {real, imag} */,
  {32'h3f9e3700, 32'h402f0630} /* (7, 1, 4) {real, imag} */,
  {32'hc02d1b90, 32'hc2fd06ee} /* (7, 1, 3) {real, imag} */,
  {32'hc2a0358f, 32'h4301b7aa} /* (7, 1, 2) {real, imag} */,
  {32'h42ec4ca6, 32'hc2c32d6d} /* (7, 1, 1) {real, imag} */,
  {32'h41b99dbc, 32'h42b71f40} /* (7, 1, 0) {real, imag} */,
  {32'hbe8f3380, 32'h42a86026} /* (7, 0, 31) {real, imag} */,
  {32'hc191f5cc, 32'h41fc1190} /* (7, 0, 30) {real, imag} */,
  {32'hc21b49ee, 32'h422476e2} /* (7, 0, 29) {real, imag} */,
  {32'hc23de0d1, 32'h4318a2ff} /* (7, 0, 28) {real, imag} */,
  {32'hc1c76b98, 32'h42c7ff14} /* (7, 0, 27) {real, imag} */,
  {32'h42f4548f, 32'hc22fb117} /* (7, 0, 26) {real, imag} */,
  {32'h4183d19c, 32'hbe4bf100} /* (7, 0, 25) {real, imag} */,
  {32'h4223400b, 32'h428f8840} /* (7, 0, 24) {real, imag} */,
  {32'hc204bddb, 32'hc1543624} /* (7, 0, 23) {real, imag} */,
  {32'hc2aa586f, 32'hbebfe9c0} /* (7, 0, 22) {real, imag} */,
  {32'h41ca0604, 32'hc1daec3d} /* (7, 0, 21) {real, imag} */,
  {32'h41fa7b08, 32'h41a7b956} /* (7, 0, 20) {real, imag} */,
  {32'h4201ffd5, 32'h400f7f30} /* (7, 0, 19) {real, imag} */,
  {32'hc0e631b8, 32'hc08de388} /* (7, 0, 18) {real, imag} */,
  {32'hc2089208, 32'h426f62b2} /* (7, 0, 17) {real, imag} */,
  {32'hc1afc62c, 32'hc1c81116} /* (7, 0, 16) {real, imag} */,
  {32'hc18bd962, 32'hc1e29123} /* (7, 0, 15) {real, imag} */,
  {32'h418a6950, 32'hc12bb3ec} /* (7, 0, 14) {real, imag} */,
  {32'hc1f1789a, 32'h425d05e1} /* (7, 0, 13) {real, imag} */,
  {32'h40b57ab0, 32'hc2a929be} /* (7, 0, 12) {real, imag} */,
  {32'hc261731e, 32'hc204d8b2} /* (7, 0, 11) {real, imag} */,
  {32'hc07023e0, 32'hc2075368} /* (7, 0, 10) {real, imag} */,
  {32'hc0fb13b8, 32'h42717f6b} /* (7, 0, 9) {real, imag} */,
  {32'h42549b79, 32'hc1e28376} /* (7, 0, 8) {real, imag} */,
  {32'hc1b3f908, 32'hc28b7d76} /* (7, 0, 7) {real, imag} */,
  {32'h42ba96ff, 32'hc192b732} /* (7, 0, 6) {real, imag} */,
  {32'hc2c6a598, 32'hc107117c} /* (7, 0, 5) {real, imag} */,
  {32'h42ff8c9c, 32'h42d8b34b} /* (7, 0, 4) {real, imag} */,
  {32'h42a7b584, 32'h4228b502} /* (7, 0, 3) {real, imag} */,
  {32'hc21f9641, 32'hc30aaf2c} /* (7, 0, 2) {real, imag} */,
  {32'h4279f326, 32'h42282e00} /* (7, 0, 1) {real, imag} */,
  {32'hc0f50dc8, 32'hc31453f1} /* (7, 0, 0) {real, imag} */,
  {32'hc2ba0944, 32'hc23ee0cc} /* (6, 31, 31) {real, imag} */,
  {32'hc1cd20b4, 32'hc2811892} /* (6, 31, 30) {real, imag} */,
  {32'h43894f81, 32'h421e08c4} /* (6, 31, 29) {real, imag} */,
  {32'hc1e3de64, 32'h43144d31} /* (6, 31, 28) {real, imag} */,
  {32'hc118ef4a, 32'h41c616cb} /* (6, 31, 27) {real, imag} */,
  {32'hc18df0c8, 32'hc2a58267} /* (6, 31, 26) {real, imag} */,
  {32'h42a5fbd2, 32'h4218b9a0} /* (6, 31, 25) {real, imag} */,
  {32'hc292d368, 32'hc25bf6e2} /* (6, 31, 24) {real, imag} */,
  {32'h4284c2c1, 32'hc0253b28} /* (6, 31, 23) {real, imag} */,
  {32'hc27e0c18, 32'h41be40d6} /* (6, 31, 22) {real, imag} */,
  {32'hc1c13c55, 32'h4200ae90} /* (6, 31, 21) {real, imag} */,
  {32'hc12ee552, 32'hc25e6bd7} /* (6, 31, 20) {real, imag} */,
  {32'h425f0898, 32'h427b5aa0} /* (6, 31, 19) {real, imag} */,
  {32'h408b75b0, 32'h40719e40} /* (6, 31, 18) {real, imag} */,
  {32'hc0f0e674, 32'hc23f0933} /* (6, 31, 17) {real, imag} */,
  {32'hc02dc500, 32'h40cf959c} /* (6, 31, 16) {real, imag} */,
  {32'h412d7dd2, 32'hc0369c30} /* (6, 31, 15) {real, imag} */,
  {32'h41afb06c, 32'hc1d6d750} /* (6, 31, 14) {real, imag} */,
  {32'hc19097d4, 32'h418e7a80} /* (6, 31, 13) {real, imag} */,
  {32'h4295daa0, 32'h423e729b} /* (6, 31, 12) {real, imag} */,
  {32'hc2809a5c, 32'h40256578} /* (6, 31, 11) {real, imag} */,
  {32'hc228b494, 32'h4153b20c} /* (6, 31, 10) {real, imag} */,
  {32'h42b4689b, 32'h424eab70} /* (6, 31, 9) {real, imag} */,
  {32'h41bfc8a0, 32'hc200fc9e} /* (6, 31, 8) {real, imag} */,
  {32'hc2628391, 32'h42a78f95} /* (6, 31, 7) {real, imag} */,
  {32'hc2939ef8, 32'hc2c4e475} /* (6, 31, 6) {real, imag} */,
  {32'h4219c744, 32'h4262d42a} /* (6, 31, 5) {real, imag} */,
  {32'hc308893e, 32'h4342d98b} /* (6, 31, 4) {real, imag} */,
  {32'h417d1ae0, 32'hc346ae4b} /* (6, 31, 3) {real, imag} */,
  {32'h4329e720, 32'h43048c46} /* (6, 31, 2) {real, imag} */,
  {32'hc11e9c5c, 32'hc21dae86} /* (6, 31, 1) {real, imag} */,
  {32'hc3445530, 32'hc1254cf2} /* (6, 31, 0) {real, imag} */,
  {32'h4343ff21, 32'h42165ac8} /* (6, 30, 31) {real, imag} */,
  {32'h43019375, 32'h41cbc0d0} /* (6, 30, 30) {real, imag} */,
  {32'h43011daa, 32'hc1f9ae84} /* (6, 30, 29) {real, imag} */,
  {32'hc28a67bc, 32'h42b98626} /* (6, 30, 28) {real, imag} */,
  {32'h413fa3e8, 32'hc1d0f7b0} /* (6, 30, 27) {real, imag} */,
  {32'hc25575f7, 32'hc1b103ea} /* (6, 30, 26) {real, imag} */,
  {32'hc1011cf2, 32'h413c8158} /* (6, 30, 25) {real, imag} */,
  {32'h4055b010, 32'h4280e5f5} /* (6, 30, 24) {real, imag} */,
  {32'hc2aac1f8, 32'hc20df8c7} /* (6, 30, 23) {real, imag} */,
  {32'hc26b8b98, 32'h3eb1b800} /* (6, 30, 22) {real, imag} */,
  {32'h3eb19cc0, 32'h41e9d8ec} /* (6, 30, 21) {real, imag} */,
  {32'hc2b33d81, 32'h42657099} /* (6, 30, 20) {real, imag} */,
  {32'h40f4e900, 32'hc23d9284} /* (6, 30, 19) {real, imag} */,
  {32'hc18a2c88, 32'hc0e42b00} /* (6, 30, 18) {real, imag} */,
  {32'hc1a6bd99, 32'hc106b126} /* (6, 30, 17) {real, imag} */,
  {32'hc142977c, 32'hc10f9ce5} /* (6, 30, 16) {real, imag} */,
  {32'hc207a8a4, 32'h41a0a31d} /* (6, 30, 15) {real, imag} */,
  {32'hbec337e0, 32'hc087b930} /* (6, 30, 14) {real, imag} */,
  {32'hc05b52e0, 32'h417439a6} /* (6, 30, 13) {real, imag} */,
  {32'h40d9d4b0, 32'hc248bc37} /* (6, 30, 12) {real, imag} */,
  {32'h41481a1e, 32'h4013c090} /* (6, 30, 11) {real, imag} */,
  {32'hc2d11bfc, 32'hc23123ee} /* (6, 30, 10) {real, imag} */,
  {32'h41be1ae8, 32'h3e88d080} /* (6, 30, 9) {real, imag} */,
  {32'h422fca05, 32'h428f1703} /* (6, 30, 8) {real, imag} */,
  {32'h4118ec0a, 32'hc11d7e22} /* (6, 30, 7) {real, imag} */,
  {32'h41ac2c82, 32'hc2dc7962} /* (6, 30, 6) {real, imag} */,
  {32'hc308ad48, 32'h42f6a060} /* (6, 30, 5) {real, imag} */,
  {32'h424ccdd4, 32'hc31abf3f} /* (6, 30, 4) {real, imag} */,
  {32'hc271957a, 32'h43271b62} /* (6, 30, 3) {real, imag} */,
  {32'h431c9cab, 32'hc3468f0c} /* (6, 30, 2) {real, imag} */,
  {32'hc303c69d, 32'h426fbfcc} /* (6, 30, 1) {real, imag} */,
  {32'hc2a9ccda, 32'hc1ffc3ac} /* (6, 30, 0) {real, imag} */,
  {32'hc1dd365a, 32'hc32ad81c} /* (6, 29, 31) {real, imag} */,
  {32'h4272ae35, 32'h4305d78c} /* (6, 29, 30) {real, imag} */,
  {32'h43137c73, 32'h41f2db98} /* (6, 29, 29) {real, imag} */,
  {32'hc2a104c9, 32'h41ff8df9} /* (6, 29, 28) {real, imag} */,
  {32'hc1596b68, 32'hc24ffc16} /* (6, 29, 27) {real, imag} */,
  {32'h413b0eb7, 32'h426a95e9} /* (6, 29, 26) {real, imag} */,
  {32'hc29da278, 32'h3eab6e80} /* (6, 29, 25) {real, imag} */,
  {32'hc196c656, 32'h4277e689} /* (6, 29, 24) {real, imag} */,
  {32'hc2a9c4c3, 32'hc298a246} /* (6, 29, 23) {real, imag} */,
  {32'hc1a804ca, 32'hc1e50a87} /* (6, 29, 22) {real, imag} */,
  {32'h42957154, 32'hc2adf11e} /* (6, 29, 21) {real, imag} */,
  {32'h40cf4e00, 32'h425224ee} /* (6, 29, 20) {real, imag} */,
  {32'h4280b83a, 32'h41dc0a11} /* (6, 29, 19) {real, imag} */,
  {32'h4236a2d9, 32'h414424ec} /* (6, 29, 18) {real, imag} */,
  {32'h41b50ec8, 32'hc1820322} /* (6, 29, 17) {real, imag} */,
  {32'h41981d48, 32'hc16e20c0} /* (6, 29, 16) {real, imag} */,
  {32'h4161ef60, 32'h418423c2} /* (6, 29, 15) {real, imag} */,
  {32'hc213b9e3, 32'h42462d6f} /* (6, 29, 14) {real, imag} */,
  {32'hc1d9206a, 32'h4195b173} /* (6, 29, 13) {real, imag} */,
  {32'h427175f0, 32'h41942454} /* (6, 29, 12) {real, imag} */,
  {32'h41ecc7f8, 32'hc2b3e3ee} /* (6, 29, 11) {real, imag} */,
  {32'hc21c87df, 32'h40c00d9c} /* (6, 29, 10) {real, imag} */,
  {32'h4190fd00, 32'hc218b7db} /* (6, 29, 9) {real, imag} */,
  {32'h430b83f1, 32'h4141393c} /* (6, 29, 8) {real, imag} */,
  {32'h4216b603, 32'hc20a58d7} /* (6, 29, 7) {real, imag} */,
  {32'h41cf05e8, 32'h423893eb} /* (6, 29, 6) {real, imag} */,
  {32'hc283e50d, 32'hc30eb8cc} /* (6, 29, 5) {real, imag} */,
  {32'hc29c1125, 32'hc11f9a06} /* (6, 29, 4) {real, imag} */,
  {32'h424e64fd, 32'h430b930d} /* (6, 29, 3) {real, imag} */,
  {32'hc27942cb, 32'h432b75f6} /* (6, 29, 2) {real, imag} */,
  {32'h4267e0bb, 32'h4116f520} /* (6, 29, 1) {real, imag} */,
  {32'h4326ee31, 32'hc381c499} /* (6, 29, 0) {real, imag} */,
  {32'hc2bc2d1a, 32'hc2d46abe} /* (6, 28, 31) {real, imag} */,
  {32'hc31603de, 32'h414fc6a8} /* (6, 28, 30) {real, imag} */,
  {32'h432e323b, 32'hc2dbbc22} /* (6, 28, 29) {real, imag} */,
  {32'h41bf32f4, 32'hc298c523} /* (6, 28, 28) {real, imag} */,
  {32'h42d41ead, 32'h428eb16a} /* (6, 28, 27) {real, imag} */,
  {32'hc3094143, 32'h419a9290} /* (6, 28, 26) {real, imag} */,
  {32'h42862526, 32'h427b3c7c} /* (6, 28, 25) {real, imag} */,
  {32'h42ad103f, 32'hc19cf149} /* (6, 28, 24) {real, imag} */,
  {32'hc14b9fa4, 32'hc1caaa41} /* (6, 28, 23) {real, imag} */,
  {32'h4089f588, 32'h418d73ab} /* (6, 28, 22) {real, imag} */,
  {32'hc0e070d0, 32'h42130ba5} /* (6, 28, 21) {real, imag} */,
  {32'h421a8aca, 32'hc1a418d5} /* (6, 28, 20) {real, imag} */,
  {32'hc27a62d8, 32'h41c585b2} /* (6, 28, 19) {real, imag} */,
  {32'h411502dc, 32'hc0c67ef0} /* (6, 28, 18) {real, imag} */,
  {32'hc1ee6b6c, 32'hc236ea68} /* (6, 28, 17) {real, imag} */,
  {32'hc162c786, 32'hc1a2825c} /* (6, 28, 16) {real, imag} */,
  {32'h41ec1d88, 32'hc0bd94b0} /* (6, 28, 15) {real, imag} */,
  {32'h41e74c3e, 32'hc0b81578} /* (6, 28, 14) {real, imag} */,
  {32'hc1fbb801, 32'hc2a5fa92} /* (6, 28, 13) {real, imag} */,
  {32'h425516f2, 32'hc2846188} /* (6, 28, 12) {real, imag} */,
  {32'hc25b5d1e, 32'h423fefcf} /* (6, 28, 11) {real, imag} */,
  {32'h4145462c, 32'h42339e90} /* (6, 28, 10) {real, imag} */,
  {32'h41a2a30e, 32'h4231c96c} /* (6, 28, 9) {real, imag} */,
  {32'h4282780d, 32'h412cf85a} /* (6, 28, 8) {real, imag} */,
  {32'h43179d7b, 32'hc1e1ddb0} /* (6, 28, 7) {real, imag} */,
  {32'hc219c3b7, 32'hc31c1902} /* (6, 28, 6) {real, imag} */,
  {32'h3e3afe00, 32'hc2b4ff5e} /* (6, 28, 5) {real, imag} */,
  {32'h42b28f7d, 32'h4254c42b} /* (6, 28, 4) {real, imag} */,
  {32'h42ebfbc2, 32'h423a55ef} /* (6, 28, 3) {real, imag} */,
  {32'h430227c8, 32'h42c2c969} /* (6, 28, 2) {real, imag} */,
  {32'hc2c8dad6, 32'h422437b3} /* (6, 28, 1) {real, imag} */,
  {32'h418ff82f, 32'h416d1a00} /* (6, 28, 0) {real, imag} */,
  {32'hc1c5ea26, 32'h425649e4} /* (6, 27, 31) {real, imag} */,
  {32'h4303b26a, 32'hc2883f88} /* (6, 27, 30) {real, imag} */,
  {32'hc11b62e0, 32'h4256204c} /* (6, 27, 29) {real, imag} */,
  {32'hc2e2e0ac, 32'hc1afaa8c} /* (6, 27, 28) {real, imag} */,
  {32'hc20b6906, 32'h4064e840} /* (6, 27, 27) {real, imag} */,
  {32'h40f337ce, 32'h4125f060} /* (6, 27, 26) {real, imag} */,
  {32'hc29e69a5, 32'h41d16dec} /* (6, 27, 25) {real, imag} */,
  {32'h42972646, 32'hc28b8f1e} /* (6, 27, 24) {real, imag} */,
  {32'h3fb7aa48, 32'h40a40e38} /* (6, 27, 23) {real, imag} */,
  {32'h427b2514, 32'h41f34150} /* (6, 27, 22) {real, imag} */,
  {32'hbffa6910, 32'hc0f12150} /* (6, 27, 21) {real, imag} */,
  {32'h41d413fb, 32'hc19726c8} /* (6, 27, 20) {real, imag} */,
  {32'h41c60ab0, 32'hc286e72b} /* (6, 27, 19) {real, imag} */,
  {32'h41228fa6, 32'h41984156} /* (6, 27, 18) {real, imag} */,
  {32'hc025a974, 32'h407ec15c} /* (6, 27, 17) {real, imag} */,
  {32'hc193ee7e, 32'hc1e43e68} /* (6, 27, 16) {real, imag} */,
  {32'hc12d7ad3, 32'h419ee658} /* (6, 27, 15) {real, imag} */,
  {32'h40642ce8, 32'h41a1822e} /* (6, 27, 14) {real, imag} */,
  {32'hc1c76df0, 32'hc19a16b9} /* (6, 27, 13) {real, imag} */,
  {32'h42aaa99b, 32'h41f30d90} /* (6, 27, 12) {real, imag} */,
  {32'h41fe7363, 32'h41864e74} /* (6, 27, 11) {real, imag} */,
  {32'hc28a68b6, 32'h41a591b6} /* (6, 27, 10) {real, imag} */,
  {32'h413d0f29, 32'hc25ccf55} /* (6, 27, 9) {real, imag} */,
  {32'hc0fc1cd8, 32'hc2804dea} /* (6, 27, 8) {real, imag} */,
  {32'h423822e2, 32'h40a5c04c} /* (6, 27, 7) {real, imag} */,
  {32'h411ce41f, 32'h410067bc} /* (6, 27, 6) {real, imag} */,
  {32'h40d6b1cc, 32'hc309dc09} /* (6, 27, 5) {real, imag} */,
  {32'hc275136c, 32'hc1c8c574} /* (6, 27, 4) {real, imag} */,
  {32'hc2187d72, 32'h41e07773} /* (6, 27, 3) {real, imag} */,
  {32'h41c75d9c, 32'h40b71fc8} /* (6, 27, 2) {real, imag} */,
  {32'hc2a0a33a, 32'hc276cb6e} /* (6, 27, 1) {real, imag} */,
  {32'h403e130c, 32'hc2ce318e} /* (6, 27, 0) {real, imag} */,
  {32'h42da9978, 32'hc2c265b2} /* (6, 26, 31) {real, imag} */,
  {32'hc17194e8, 32'h41c4dbda} /* (6, 26, 30) {real, imag} */,
  {32'hc1d2a23c, 32'h42da16d0} /* (6, 26, 29) {real, imag} */,
  {32'hc1159794, 32'hc2d03152} /* (6, 26, 28) {real, imag} */,
  {32'hc1b1a13e, 32'hc102ed64} /* (6, 26, 27) {real, imag} */,
  {32'h4190adfc, 32'h4209f1c4} /* (6, 26, 26) {real, imag} */,
  {32'h425ee2f9, 32'hc1d166f4} /* (6, 26, 25) {real, imag} */,
  {32'h40ea1318, 32'h42c128c0} /* (6, 26, 24) {real, imag} */,
  {32'h425657a6, 32'h4253df2a} /* (6, 26, 23) {real, imag} */,
  {32'hc252ec50, 32'h409da8de} /* (6, 26, 22) {real, imag} */,
  {32'hc0b10acc, 32'hc15d211c} /* (6, 26, 21) {real, imag} */,
  {32'h415d4c39, 32'hc195cbc4} /* (6, 26, 20) {real, imag} */,
  {32'hc1e04672, 32'h4283b14c} /* (6, 26, 19) {real, imag} */,
  {32'h412df428, 32'hc0c2056c} /* (6, 26, 18) {real, imag} */,
  {32'hc0bdb42c, 32'h418399e6} /* (6, 26, 17) {real, imag} */,
  {32'h41b8166a, 32'hbed4d300} /* (6, 26, 16) {real, imag} */,
  {32'hc12b63c2, 32'hbf164430} /* (6, 26, 15) {real, imag} */,
  {32'h40238b10, 32'hc1a74cc0} /* (6, 26, 14) {real, imag} */,
  {32'hc21843fb, 32'hc19d34a2} /* (6, 26, 13) {real, imag} */,
  {32'h411de987, 32'hc16aa8b8} /* (6, 26, 12) {real, imag} */,
  {32'h42042a32, 32'h41485b60} /* (6, 26, 11) {real, imag} */,
  {32'hc21eb608, 32'hc1659fb7} /* (6, 26, 10) {real, imag} */,
  {32'h3fe32f10, 32'h406a0388} /* (6, 26, 9) {real, imag} */,
  {32'hc20ec687, 32'hc191a1c6} /* (6, 26, 8) {real, imag} */,
  {32'hc2394ebf, 32'hc2ff4abf} /* (6, 26, 7) {real, imag} */,
  {32'h42d90949, 32'h428f9681} /* (6, 26, 6) {real, imag} */,
  {32'h42869f14, 32'h40fe4670} /* (6, 26, 5) {real, imag} */,
  {32'h420a23e3, 32'h42d8333a} /* (6, 26, 4) {real, imag} */,
  {32'h4324ddae, 32'hbff8b7e0} /* (6, 26, 3) {real, imag} */,
  {32'hc2b59c57, 32'h40f4acea} /* (6, 26, 2) {real, imag} */,
  {32'h427a3128, 32'hc2083bad} /* (6, 26, 1) {real, imag} */,
  {32'h41d6bc66, 32'h431b2bca} /* (6, 26, 0) {real, imag} */,
  {32'h42aa7709, 32'hc2c14bde} /* (6, 25, 31) {real, imag} */,
  {32'hc12390fc, 32'h41d26e05} /* (6, 25, 30) {real, imag} */,
  {32'h406976e9, 32'h4321862d} /* (6, 25, 29) {real, imag} */,
  {32'h41b22baa, 32'h41163c08} /* (6, 25, 28) {real, imag} */,
  {32'h41a224e4, 32'h4144f6e0} /* (6, 25, 27) {real, imag} */,
  {32'hc1dd482c, 32'hc29a0e5a} /* (6, 25, 26) {real, imag} */,
  {32'hc0fe183a, 32'hc267669b} /* (6, 25, 25) {real, imag} */,
  {32'h41afb220, 32'h4283e461} /* (6, 25, 24) {real, imag} */,
  {32'hc142bcce, 32'h41326232} /* (6, 25, 23) {real, imag} */,
  {32'hc21472d7, 32'h410423ff} /* (6, 25, 22) {real, imag} */,
  {32'h4202cb83, 32'h4184b4d4} /* (6, 25, 21) {real, imag} */,
  {32'h414d73e3, 32'hbf149fb0} /* (6, 25, 20) {real, imag} */,
  {32'hc127d15e, 32'hc0232a10} /* (6, 25, 19) {real, imag} */,
  {32'hbf963920, 32'hc21773c5} /* (6, 25, 18) {real, imag} */,
  {32'hc088d7c6, 32'hc22a8ef6} /* (6, 25, 17) {real, imag} */,
  {32'hc1a2fee8, 32'h41a637bc} /* (6, 25, 16) {real, imag} */,
  {32'h413ac133, 32'h41a44f58} /* (6, 25, 15) {real, imag} */,
  {32'hc1eebd94, 32'h41b37099} /* (6, 25, 14) {real, imag} */,
  {32'hc0ce3368, 32'hc1f320ba} /* (6, 25, 13) {real, imag} */,
  {32'hc1dae4e6, 32'h3f8c75e8} /* (6, 25, 12) {real, imag} */,
  {32'h4225e9dd, 32'hc252800e} /* (6, 25, 11) {real, imag} */,
  {32'hc0c7a228, 32'h42099ea9} /* (6, 25, 10) {real, imag} */,
  {32'h41240930, 32'hc0387ea8} /* (6, 25, 9) {real, imag} */,
  {32'hc2b2c89e, 32'hc1914844} /* (6, 25, 8) {real, imag} */,
  {32'h41c9045e, 32'h41d2925a} /* (6, 25, 7) {real, imag} */,
  {32'hc2015e6e, 32'hc23eebad} /* (6, 25, 6) {real, imag} */,
  {32'h40f98bae, 32'h4294cf7c} /* (6, 25, 5) {real, imag} */,
  {32'hc29730f2, 32'hc28ffcf7} /* (6, 25, 4) {real, imag} */,
  {32'h3f8f31be, 32'hc23315b1} /* (6, 25, 3) {real, imag} */,
  {32'hc22b36ca, 32'hc17a0c52} /* (6, 25, 2) {real, imag} */,
  {32'h4290dbe5, 32'hc2d4311a} /* (6, 25, 1) {real, imag} */,
  {32'hc23b07fc, 32'hc2a2e485} /* (6, 25, 0) {real, imag} */,
  {32'hc269a40f, 32'h4225184d} /* (6, 24, 31) {real, imag} */,
  {32'h4289f37d, 32'hc33115ec} /* (6, 24, 30) {real, imag} */,
  {32'hc02f21e4, 32'hc2968b92} /* (6, 24, 29) {real, imag} */,
  {32'h42803c72, 32'hc1c1b276} /* (6, 24, 28) {real, imag} */,
  {32'hc219819d, 32'h41253e8e} /* (6, 24, 27) {real, imag} */,
  {32'h416efac4, 32'hc0e01280} /* (6, 24, 26) {real, imag} */,
  {32'h42ca4292, 32'h41c1de4a} /* (6, 24, 25) {real, imag} */,
  {32'h41a8cf63, 32'h41deb2a0} /* (6, 24, 24) {real, imag} */,
  {32'h4262f0c0, 32'hc1f26245} /* (6, 24, 23) {real, imag} */,
  {32'hc16534a2, 32'hc26184c2} /* (6, 24, 22) {real, imag} */,
  {32'hc1af8542, 32'hc212fc30} /* (6, 24, 21) {real, imag} */,
  {32'hc1426ec8, 32'hc190c439} /* (6, 24, 20) {real, imag} */,
  {32'hc1f51bb6, 32'h41c0b3b6} /* (6, 24, 19) {real, imag} */,
  {32'h41f29448, 32'hc19947ee} /* (6, 24, 18) {real, imag} */,
  {32'hc160ed1e, 32'hc1adf7d4} /* (6, 24, 17) {real, imag} */,
  {32'hc16071a0, 32'h41b73d10} /* (6, 24, 16) {real, imag} */,
  {32'h40677198, 32'h412d9229} /* (6, 24, 15) {real, imag} */,
  {32'h40f85e40, 32'hc20a6f1b} /* (6, 24, 14) {real, imag} */,
  {32'hc0ca55fa, 32'h416de18b} /* (6, 24, 13) {real, imag} */,
  {32'h41f3c880, 32'hc166fca2} /* (6, 24, 12) {real, imag} */,
  {32'hc1f2d7ac, 32'hc2381544} /* (6, 24, 11) {real, imag} */,
  {32'h41f5fd79, 32'h41f8c743} /* (6, 24, 10) {real, imag} */,
  {32'h41418810, 32'hc1b55fe7} /* (6, 24, 9) {real, imag} */,
  {32'hc2a1b808, 32'hbff00528} /* (6, 24, 8) {real, imag} */,
  {32'h41136e60, 32'h401e5714} /* (6, 24, 7) {real, imag} */,
  {32'hc27a5b1b, 32'hc2b1e84c} /* (6, 24, 6) {real, imag} */,
  {32'hc170cd47, 32'h40b80fa3} /* (6, 24, 5) {real, imag} */,
  {32'h41d7bdde, 32'h4257a92d} /* (6, 24, 4) {real, imag} */,
  {32'hc0df9bae, 32'hc2aa83d6} /* (6, 24, 3) {real, imag} */,
  {32'hc2fc998d, 32'h4318ec84} /* (6, 24, 2) {real, imag} */,
  {32'hc1e7e766, 32'hc165aa3b} /* (6, 24, 1) {real, imag} */,
  {32'h42d9646a, 32'h421537ae} /* (6, 24, 0) {real, imag} */,
  {32'h4185f0a2, 32'hc172ae30} /* (6, 23, 31) {real, imag} */,
  {32'h42470d92, 32'hc1ef6203} /* (6, 23, 30) {real, imag} */,
  {32'h425579e8, 32'hc162adb0} /* (6, 23, 29) {real, imag} */,
  {32'h41d1ed85, 32'hc1eda8ae} /* (6, 23, 28) {real, imag} */,
  {32'h417e619a, 32'hc191177b} /* (6, 23, 27) {real, imag} */,
  {32'h40787598, 32'h428438eb} /* (6, 23, 26) {real, imag} */,
  {32'h4258e3ba, 32'hc05ada10} /* (6, 23, 25) {real, imag} */,
  {32'hc1229aa2, 32'hc1df03ba} /* (6, 23, 24) {real, imag} */,
  {32'h4288e649, 32'h415737b2} /* (6, 23, 23) {real, imag} */,
  {32'hc164e3d1, 32'h42402d41} /* (6, 23, 22) {real, imag} */,
  {32'h4159e161, 32'h420ec2f3} /* (6, 23, 21) {real, imag} */,
  {32'hc19e9d8e, 32'hc0f44fd4} /* (6, 23, 20) {real, imag} */,
  {32'hc04233c0, 32'hc1462a54} /* (6, 23, 19) {real, imag} */,
  {32'h418caf36, 32'h4175046e} /* (6, 23, 18) {real, imag} */,
  {32'hc1809284, 32'hc0d5942c} /* (6, 23, 17) {real, imag} */,
  {32'hc1f42998, 32'hc1e1f767} /* (6, 23, 16) {real, imag} */,
  {32'hc138cea5, 32'hc0d9f39c} /* (6, 23, 15) {real, imag} */,
  {32'hc14fe07d, 32'hc2125f5a} /* (6, 23, 14) {real, imag} */,
  {32'hc0fea95c, 32'h4112d3a2} /* (6, 23, 13) {real, imag} */,
  {32'h41b1cca2, 32'hc1a322a9} /* (6, 23, 12) {real, imag} */,
  {32'h41322559, 32'h4222aec9} /* (6, 23, 11) {real, imag} */,
  {32'h41b1d1d6, 32'hc23e7abd} /* (6, 23, 10) {real, imag} */,
  {32'hc11c9600, 32'hc1eda931} /* (6, 23, 9) {real, imag} */,
  {32'hc2178af0, 32'h41022b3f} /* (6, 23, 8) {real, imag} */,
  {32'h409eb520, 32'h422a549e} /* (6, 23, 7) {real, imag} */,
  {32'h420f9f26, 32'hc1683e12} /* (6, 23, 6) {real, imag} */,
  {32'h4212e484, 32'h42972ea4} /* (6, 23, 5) {real, imag} */,
  {32'hc262df7a, 32'h41dc433e} /* (6, 23, 4) {real, imag} */,
  {32'hbfea0980, 32'h4275c726} /* (6, 23, 3) {real, imag} */,
  {32'hc077e100, 32'hc2bb98c4} /* (6, 23, 2) {real, imag} */,
  {32'h413979d7, 32'h415f8708} /* (6, 23, 1) {real, imag} */,
  {32'h424c1824, 32'hc22ecf4f} /* (6, 23, 0) {real, imag} */,
  {32'h3e066a40, 32'hc0d8f8e4} /* (6, 22, 31) {real, imag} */,
  {32'hc19c66d4, 32'h41bafe50} /* (6, 22, 30) {real, imag} */,
  {32'h4287a710, 32'h424b4500} /* (6, 22, 29) {real, imag} */,
  {32'hc1a6fda8, 32'hc290dd06} /* (6, 22, 28) {real, imag} */,
  {32'h418711b7, 32'hc0117f70} /* (6, 22, 27) {real, imag} */,
  {32'h4299b7c0, 32'hc1802f6a} /* (6, 22, 26) {real, imag} */,
  {32'hbf107710, 32'hc18fe5a6} /* (6, 22, 25) {real, imag} */,
  {32'h42140b48, 32'h4281ae7c} /* (6, 22, 24) {real, imag} */,
  {32'hc0d01e12, 32'hc1b0fa8c} /* (6, 22, 23) {real, imag} */,
  {32'hc1b3f50c, 32'hc17bec4c} /* (6, 22, 22) {real, imag} */,
  {32'hc14b0a88, 32'h4110aea0} /* (6, 22, 21) {real, imag} */,
  {32'h4121b2fe, 32'hc0600d8c} /* (6, 22, 20) {real, imag} */,
  {32'hc138dc99, 32'hbfefbba8} /* (6, 22, 19) {real, imag} */,
  {32'h40b7caba, 32'h4181d5f3} /* (6, 22, 18) {real, imag} */,
  {32'hbfb1ea68, 32'h40341b70} /* (6, 22, 17) {real, imag} */,
  {32'h41c08d50, 32'h40d20cec} /* (6, 22, 16) {real, imag} */,
  {32'hbf289340, 32'hc2075783} /* (6, 22, 15) {real, imag} */,
  {32'h40cf952e, 32'hc0c9f704} /* (6, 22, 14) {real, imag} */,
  {32'hc14f513f, 32'hc083a01a} /* (6, 22, 13) {real, imag} */,
  {32'h41877c89, 32'hc01a9afc} /* (6, 22, 12) {real, imag} */,
  {32'hc11e4370, 32'hbfd9ca00} /* (6, 22, 11) {real, imag} */,
  {32'h40dd7920, 32'h4232c7ef} /* (6, 22, 10) {real, imag} */,
  {32'h41b4ca56, 32'h40e462a8} /* (6, 22, 9) {real, imag} */,
  {32'h42ac6fa0, 32'hc1ffcfe7} /* (6, 22, 8) {real, imag} */,
  {32'hc20233a1, 32'h42172bda} /* (6, 22, 7) {real, imag} */,
  {32'hc10d2e6c, 32'hc2adbade} /* (6, 22, 6) {real, imag} */,
  {32'hc1c8f7f3, 32'h4295019a} /* (6, 22, 5) {real, imag} */,
  {32'hc0bb991f, 32'h4186e5f0} /* (6, 22, 4) {real, imag} */,
  {32'h42a729f0, 32'h40369920} /* (6, 22, 3) {real, imag} */,
  {32'hc245e786, 32'h41c10a3e} /* (6, 22, 2) {real, imag} */,
  {32'hc15b1f3e, 32'h41ec4997} /* (6, 22, 1) {real, imag} */,
  {32'hc2779628, 32'hc206d598} /* (6, 22, 0) {real, imag} */,
  {32'h41f8cd3d, 32'h420d78b9} /* (6, 21, 31) {real, imag} */,
  {32'hc18a85c7, 32'hc1387600} /* (6, 21, 30) {real, imag} */,
  {32'hc29232b5, 32'h4168c1c8} /* (6, 21, 29) {real, imag} */,
  {32'h41834714, 32'hc2830d8d} /* (6, 21, 28) {real, imag} */,
  {32'hc0f7d478, 32'hc10141de} /* (6, 21, 27) {real, imag} */,
  {32'hc2293dc5, 32'h41cb339a} /* (6, 21, 26) {real, imag} */,
  {32'h4019be70, 32'h41c92498} /* (6, 21, 25) {real, imag} */,
  {32'h418d9d90, 32'hc20e6d0a} /* (6, 21, 24) {real, imag} */,
  {32'h418bf4c6, 32'hc27d8c55} /* (6, 21, 23) {real, imag} */,
  {32'hc129f2ec, 32'h4128bd1e} /* (6, 21, 22) {real, imag} */,
  {32'hc1837386, 32'h419eec9c} /* (6, 21, 21) {real, imag} */,
  {32'hc08e50e4, 32'hc1999b45} /* (6, 21, 20) {real, imag} */,
  {32'hc1705f64, 32'hc1d54e64} /* (6, 21, 19) {real, imag} */,
  {32'h40c3b2b8, 32'h3f39eee0} /* (6, 21, 18) {real, imag} */,
  {32'hc0e11018, 32'h41b00549} /* (6, 21, 17) {real, imag} */,
  {32'hc097c06e, 32'hc12c2a7e} /* (6, 21, 16) {real, imag} */,
  {32'h4112e040, 32'h40bba838} /* (6, 21, 15) {real, imag} */,
  {32'hc0fee6d0, 32'h416346a6} /* (6, 21, 14) {real, imag} */,
  {32'h4021568e, 32'hc1c46570} /* (6, 21, 13) {real, imag} */,
  {32'hc1cc63eb, 32'hc1a86d87} /* (6, 21, 12) {real, imag} */,
  {32'hc1659695, 32'h4170b3a8} /* (6, 21, 11) {real, imag} */,
  {32'h4091c660, 32'hc12257f8} /* (6, 21, 10) {real, imag} */,
  {32'h410c7567, 32'h41ba68e6} /* (6, 21, 9) {real, imag} */,
  {32'h41cb676c, 32'h40e1dacc} /* (6, 21, 8) {real, imag} */,
  {32'hc1f81566, 32'hc228bf94} /* (6, 21, 7) {real, imag} */,
  {32'hc1c415ee, 32'h40b9f336} /* (6, 21, 6) {real, imag} */,
  {32'hc2542c33, 32'h404e42b6} /* (6, 21, 5) {real, imag} */,
  {32'hc1ccbde0, 32'hc23ffe70} /* (6, 21, 4) {real, imag} */,
  {32'h42226d00, 32'hc1884b24} /* (6, 21, 3) {real, imag} */,
  {32'h4298f8f4, 32'hc1af4a50} /* (6, 21, 2) {real, imag} */,
  {32'hc2968d6b, 32'h41a8cfe2} /* (6, 21, 1) {real, imag} */,
  {32'h4208fc03, 32'hc0e202b4} /* (6, 21, 0) {real, imag} */,
  {32'hc2233f85, 32'h41b7ac02} /* (6, 20, 31) {real, imag} */,
  {32'h427271e7, 32'h42398b82} /* (6, 20, 30) {real, imag} */,
  {32'hc054a280, 32'hc2248600} /* (6, 20, 29) {real, imag} */,
  {32'hc0d304b8, 32'hc199be90} /* (6, 20, 28) {real, imag} */,
  {32'hc03dd4a0, 32'h41e4a9ac} /* (6, 20, 27) {real, imag} */,
  {32'h4128a822, 32'hc0a425f6} /* (6, 20, 26) {real, imag} */,
  {32'h3f39bf94, 32'h4118fe06} /* (6, 20, 25) {real, imag} */,
  {32'h41d71189, 32'hc25713d6} /* (6, 20, 24) {real, imag} */,
  {32'hc1ad2659, 32'h4195b48c} /* (6, 20, 23) {real, imag} */,
  {32'h41990576, 32'hc1de342a} /* (6, 20, 22) {real, imag} */,
  {32'hc1503954, 32'hc14a7b86} /* (6, 20, 21) {real, imag} */,
  {32'h41a41dc6, 32'h406ce4f8} /* (6, 20, 20) {real, imag} */,
  {32'h40bd49b4, 32'hc0f97f9e} /* (6, 20, 19) {real, imag} */,
  {32'hc02ab504, 32'h41a7c965} /* (6, 20, 18) {real, imag} */,
  {32'hbeacfba0, 32'h3ff91868} /* (6, 20, 17) {real, imag} */,
  {32'hc0ae2081, 32'h4185aff5} /* (6, 20, 16) {real, imag} */,
  {32'h4102d6a7, 32'h4184e030} /* (6, 20, 15) {real, imag} */,
  {32'hbf384df0, 32'h40faf81c} /* (6, 20, 14) {real, imag} */,
  {32'h41913f12, 32'hc085da36} /* (6, 20, 13) {real, imag} */,
  {32'hc1797c05, 32'hc133e90e} /* (6, 20, 12) {real, imag} */,
  {32'h41ab91ca, 32'h419293be} /* (6, 20, 11) {real, imag} */,
  {32'h416d3e10, 32'hc14d1dc1} /* (6, 20, 10) {real, imag} */,
  {32'h4187b037, 32'hc194f67c} /* (6, 20, 9) {real, imag} */,
  {32'hc202a464, 32'h412146d2} /* (6, 20, 8) {real, imag} */,
  {32'h3f79d7b4, 32'hc1895e89} /* (6, 20, 7) {real, imag} */,
  {32'hc2102dc8, 32'h4199e48a} /* (6, 20, 6) {real, imag} */,
  {32'hc1958a48, 32'hc215a820} /* (6, 20, 5) {real, imag} */,
  {32'hc207d209, 32'h421e093b} /* (6, 20, 4) {real, imag} */,
  {32'hc20de510, 32'h41f94920} /* (6, 20, 3) {real, imag} */,
  {32'h41cf7632, 32'h40c924e0} /* (6, 20, 2) {real, imag} */,
  {32'h411ee0b5, 32'hc1ab4a8a} /* (6, 20, 1) {real, imag} */,
  {32'h41577cce, 32'h4215fa5e} /* (6, 20, 0) {real, imag} */,
  {32'hc1a0fbba, 32'h4270d058} /* (6, 19, 31) {real, imag} */,
  {32'h41031037, 32'hc211440f} /* (6, 19, 30) {real, imag} */,
  {32'hc1a974ef, 32'h41665680} /* (6, 19, 29) {real, imag} */,
  {32'hc1a95114, 32'hc1c90d62} /* (6, 19, 28) {real, imag} */,
  {32'hc097f55e, 32'hc01a2ad2} /* (6, 19, 27) {real, imag} */,
  {32'hc1b7556e, 32'h413ed610} /* (6, 19, 26) {real, imag} */,
  {32'hc241c624, 32'hc0e8d12f} /* (6, 19, 25) {real, imag} */,
  {32'h41d076b6, 32'hc118d537} /* (6, 19, 24) {real, imag} */,
  {32'hc19357e3, 32'h40438646} /* (6, 19, 23) {real, imag} */,
  {32'hc098197c, 32'h4143c06e} /* (6, 19, 22) {real, imag} */,
  {32'h400eb97e, 32'hc17413cf} /* (6, 19, 21) {real, imag} */,
  {32'h4013e250, 32'hc16da261} /* (6, 19, 20) {real, imag} */,
  {32'h4118f005, 32'hc16fe5d2} /* (6, 19, 19) {real, imag} */,
  {32'hbf699bd8, 32'h4123805a} /* (6, 19, 18) {real, imag} */,
  {32'h40ce7c12, 32'h4042608c} /* (6, 19, 17) {real, imag} */,
  {32'h3fa2feb4, 32'h3fa66560} /* (6, 19, 16) {real, imag} */,
  {32'hc1470003, 32'hc0cbee2e} /* (6, 19, 15) {real, imag} */,
  {32'hc0de3ff3, 32'hc1748a00} /* (6, 19, 14) {real, imag} */,
  {32'hc10b9deb, 32'hc06a2fba} /* (6, 19, 13) {real, imag} */,
  {32'hc1b24be0, 32'hbe8a32e0} /* (6, 19, 12) {real, imag} */,
  {32'hc0b78f55, 32'h41645195} /* (6, 19, 11) {real, imag} */,
  {32'h41c1f9fb, 32'hc14715fe} /* (6, 19, 10) {real, imag} */,
  {32'h4215ad9a, 32'hc1400c4e} /* (6, 19, 9) {real, imag} */,
  {32'h41103959, 32'h41374d1d} /* (6, 19, 8) {real, imag} */,
  {32'hc14dc91a, 32'hc0d01877} /* (6, 19, 7) {real, imag} */,
  {32'hc1bf08b2, 32'h4132b384} /* (6, 19, 6) {real, imag} */,
  {32'h41cab528, 32'hc17cd26a} /* (6, 19, 5) {real, imag} */,
  {32'hc09d98e8, 32'hc1db4702} /* (6, 19, 4) {real, imag} */,
  {32'hc1df0e7d, 32'h4012b80e} /* (6, 19, 3) {real, imag} */,
  {32'h41bf82b4, 32'h41d7c55e} /* (6, 19, 2) {real, imag} */,
  {32'hc17230a4, 32'h3eca32c0} /* (6, 19, 1) {real, imag} */,
  {32'hc0fbe02b, 32'hc1e9a8fb} /* (6, 19, 0) {real, imag} */,
  {32'hc23c4a9a, 32'hc14d4a36} /* (6, 18, 31) {real, imag} */,
  {32'hc112a992, 32'h40c5103c} /* (6, 18, 30) {real, imag} */,
  {32'h41fbde78, 32'h424a1547} /* (6, 18, 29) {real, imag} */,
  {32'hc1f89222, 32'h41e0ef95} /* (6, 18, 28) {real, imag} */,
  {32'hbf548e10, 32'h40e23758} /* (6, 18, 27) {real, imag} */,
  {32'hc1dc80e7, 32'hc1c833d2} /* (6, 18, 26) {real, imag} */,
  {32'h405c4660, 32'h413bdbc2} /* (6, 18, 25) {real, imag} */,
  {32'h402c5493, 32'h40f26703} /* (6, 18, 24) {real, imag} */,
  {32'hc1fc4ea8, 32'hc021e0f0} /* (6, 18, 23) {real, imag} */,
  {32'h40d9dc32, 32'hc0f3d0ce} /* (6, 18, 22) {real, imag} */,
  {32'hc0ed9b5e, 32'h41032581} /* (6, 18, 21) {real, imag} */,
  {32'hc0946a59, 32'hc15047d0} /* (6, 18, 20) {real, imag} */,
  {32'h408d4446, 32'hc121f078} /* (6, 18, 19) {real, imag} */,
  {32'hc17d7b08, 32'hbf08bc58} /* (6, 18, 18) {real, imag} */,
  {32'hc0acc128, 32'hbfc54c64} /* (6, 18, 17) {real, imag} */,
  {32'hc0553879, 32'h3fc6a078} /* (6, 18, 16) {real, imag} */,
  {32'hc1460540, 32'h3f530638} /* (6, 18, 15) {real, imag} */,
  {32'h40ca4000, 32'h412a867e} /* (6, 18, 14) {real, imag} */,
  {32'h4011f3f4, 32'hc08b3437} /* (6, 18, 13) {real, imag} */,
  {32'hbfeb7e7c, 32'hc0805530} /* (6, 18, 12) {real, imag} */,
  {32'h40d705c2, 32'h3fc95a38} /* (6, 18, 11) {real, imag} */,
  {32'hc193392a, 32'h41c7005c} /* (6, 18, 10) {real, imag} */,
  {32'hc0858bae, 32'h418adbc2} /* (6, 18, 9) {real, imag} */,
  {32'h3e47d1b0, 32'h4197d943} /* (6, 18, 8) {real, imag} */,
  {32'h42137ffe, 32'h4142253e} /* (6, 18, 7) {real, imag} */,
  {32'h420784ea, 32'h41db4d76} /* (6, 18, 6) {real, imag} */,
  {32'hbfd70228, 32'h417286d2} /* (6, 18, 5) {real, imag} */,
  {32'hc261e6f3, 32'h40f5a56c} /* (6, 18, 4) {real, imag} */,
  {32'h418117b8, 32'hc26696b5} /* (6, 18, 3) {real, imag} */,
  {32'hc12143e6, 32'h40d6bc9a} /* (6, 18, 2) {real, imag} */,
  {32'h40c7ad68, 32'h41ff702d} /* (6, 18, 1) {real, imag} */,
  {32'h40125edb, 32'hc1731ee3} /* (6, 18, 0) {real, imag} */,
  {32'h415f48a4, 32'h40b19582} /* (6, 17, 31) {real, imag} */,
  {32'h42744d39, 32'h42226a93} /* (6, 17, 30) {real, imag} */,
  {32'hc113b21a, 32'h406c0548} /* (6, 17, 29) {real, imag} */,
  {32'hc1ca69f3, 32'h41b5eab9} /* (6, 17, 28) {real, imag} */,
  {32'hc18f0a32, 32'hc1ae0ce6} /* (6, 17, 27) {real, imag} */,
  {32'hc20e75b8, 32'hc18bde26} /* (6, 17, 26) {real, imag} */,
  {32'h40834240, 32'h41255ebd} /* (6, 17, 25) {real, imag} */,
  {32'h3f27dbd8, 32'h413f08cc} /* (6, 17, 24) {real, imag} */,
  {32'h41814287, 32'h40f92471} /* (6, 17, 23) {real, imag} */,
  {32'hc1041fc2, 32'hbc6d6c00} /* (6, 17, 22) {real, imag} */,
  {32'hc0a808a6, 32'h414e678d} /* (6, 17, 21) {real, imag} */,
  {32'h4101317c, 32'hc0ba55bf} /* (6, 17, 20) {real, imag} */,
  {32'hc0c7c5b2, 32'hc125c086} /* (6, 17, 19) {real, imag} */,
  {32'h3fcdde08, 32'h41419a84} /* (6, 17, 18) {real, imag} */,
  {32'hbfb5093c, 32'hc0e678e2} /* (6, 17, 17) {real, imag} */,
  {32'hc1922365, 32'h402e5bb8} /* (6, 17, 16) {real, imag} */,
  {32'h412e3afe, 32'hc05e903c} /* (6, 17, 15) {real, imag} */,
  {32'h41050039, 32'hc0475622} /* (6, 17, 14) {real, imag} */,
  {32'hc109b1c9, 32'hc0ff2e6c} /* (6, 17, 13) {real, imag} */,
  {32'hbfe3d600, 32'h40b8dddf} /* (6, 17, 12) {real, imag} */,
  {32'h3cf11680, 32'h3f9ea7f0} /* (6, 17, 11) {real, imag} */,
  {32'hc1bf2ffb, 32'hc19a68e0} /* (6, 17, 10) {real, imag} */,
  {32'h3f78e998, 32'hc0e25e4b} /* (6, 17, 9) {real, imag} */,
  {32'hc10a6b86, 32'hc1ad256c} /* (6, 17, 8) {real, imag} */,
  {32'hc19c85a0, 32'h41ac41d6} /* (6, 17, 7) {real, imag} */,
  {32'hc09eed94, 32'h4158bff6} /* (6, 17, 6) {real, imag} */,
  {32'hc1b95272, 32'hc158e390} /* (6, 17, 5) {real, imag} */,
  {32'h42001f9c, 32'hc0318b98} /* (6, 17, 4) {real, imag} */,
  {32'h41b878df, 32'h42191acc} /* (6, 17, 3) {real, imag} */,
  {32'hc2a9b2e7, 32'h4147a2c0} /* (6, 17, 2) {real, imag} */,
  {32'hc13b5b70, 32'h405611cc} /* (6, 17, 1) {real, imag} */,
  {32'hc219bc38, 32'hc087fb3e} /* (6, 17, 0) {real, imag} */,
  {32'h413bf624, 32'hc1674e94} /* (6, 16, 31) {real, imag} */,
  {32'h419166f2, 32'h411bff94} /* (6, 16, 30) {real, imag} */,
  {32'h41a8a990, 32'h410afacb} /* (6, 16, 29) {real, imag} */,
  {32'hc1706239, 32'hc00f233b} /* (6, 16, 28) {real, imag} */,
  {32'hc16248e3, 32'hc190443a} /* (6, 16, 27) {real, imag} */,
  {32'hc104e18a, 32'h41a078a6} /* (6, 16, 26) {real, imag} */,
  {32'h40826815, 32'hc115cde4} /* (6, 16, 25) {real, imag} */,
  {32'h413cddab, 32'hc1491a27} /* (6, 16, 24) {real, imag} */,
  {32'h403dfa79, 32'h3f1b2688} /* (6, 16, 23) {real, imag} */,
  {32'h40394bde, 32'h3eaeab60} /* (6, 16, 22) {real, imag} */,
  {32'h407386c6, 32'h41256ba0} /* (6, 16, 21) {real, imag} */,
  {32'h413ea319, 32'h3f9111a8} /* (6, 16, 20) {real, imag} */,
  {32'h40c95dcb, 32'h4005494a} /* (6, 16, 19) {real, imag} */,
  {32'h410a61c1, 32'hc121fee1} /* (6, 16, 18) {real, imag} */,
  {32'h413c23c3, 32'h40babb2d} /* (6, 16, 17) {real, imag} */,
  {32'h3faa1378, 32'hc0d4346c} /* (6, 16, 16) {real, imag} */,
  {32'hc00c13c8, 32'hc057b0a2} /* (6, 16, 15) {real, imag} */,
  {32'h40eb3790, 32'hc17b0781} /* (6, 16, 14) {real, imag} */,
  {32'h410af18a, 32'hc0a1df41} /* (6, 16, 13) {real, imag} */,
  {32'hc0fbb58a, 32'h411a90b1} /* (6, 16, 12) {real, imag} */,
  {32'h400c70aa, 32'h40709516} /* (6, 16, 11) {real, imag} */,
  {32'hbf8a0d58, 32'hc1961cce} /* (6, 16, 10) {real, imag} */,
  {32'hc1237472, 32'h4144038a} /* (6, 16, 9) {real, imag} */,
  {32'hc000e898, 32'hbff4ec40} /* (6, 16, 8) {real, imag} */,
  {32'h4012cb78, 32'hc0961285} /* (6, 16, 7) {real, imag} */,
  {32'hc0c97820, 32'hc181506a} /* (6, 16, 6) {real, imag} */,
  {32'hc184fc11, 32'h41d6ad2e} /* (6, 16, 5) {real, imag} */,
  {32'hc21c2c6a, 32'h3ff527f6} /* (6, 16, 4) {real, imag} */,
  {32'h4151f9e0, 32'hc13c0d61} /* (6, 16, 3) {real, imag} */,
  {32'h40123690, 32'h41a9e6fd} /* (6, 16, 2) {real, imag} */,
  {32'h3d413300, 32'hc1b9bdbe} /* (6, 16, 1) {real, imag} */,
  {32'h411a2890, 32'h41085827} /* (6, 16, 0) {real, imag} */,
  {32'h41a2c8dc, 32'hc1f8a322} /* (6, 15, 31) {real, imag} */,
  {32'h418d945c, 32'h41b1dda0} /* (6, 15, 30) {real, imag} */,
  {32'h408fd580, 32'hc22a151c} /* (6, 15, 29) {real, imag} */,
  {32'h4050f418, 32'h41b39769} /* (6, 15, 28) {real, imag} */,
  {32'hc1cc0352, 32'hc1e5b734} /* (6, 15, 27) {real, imag} */,
  {32'h41b741dd, 32'h41c07592} /* (6, 15, 26) {real, imag} */,
  {32'h4188da16, 32'hc1fef4d2} /* (6, 15, 25) {real, imag} */,
  {32'hc211f80b, 32'hc1d6a0ae} /* (6, 15, 24) {real, imag} */,
  {32'h40423790, 32'hc1010c8c} /* (6, 15, 23) {real, imag} */,
  {32'hc089c6d8, 32'hc1052632} /* (6, 15, 22) {real, imag} */,
  {32'hc1ad1484, 32'hc0366042} /* (6, 15, 21) {real, imag} */,
  {32'hbfd3e9ec, 32'h3ed97638} /* (6, 15, 20) {real, imag} */,
  {32'hbfda4b70, 32'h41543e1a} /* (6, 15, 19) {real, imag} */,
  {32'hc1418b27, 32'hc076bd75} /* (6, 15, 18) {real, imag} */,
  {32'hc0752ca4, 32'h3f96b1e8} /* (6, 15, 17) {real, imag} */,
  {32'h40ca4c90, 32'h40845dba} /* (6, 15, 16) {real, imag} */,
  {32'h3e3696c8, 32'hc0f0d662} /* (6, 15, 15) {real, imag} */,
  {32'hc069f374, 32'hc0a5ce86} /* (6, 15, 14) {real, imag} */,
  {32'h408a9780, 32'h40e810d4} /* (6, 15, 13) {real, imag} */,
  {32'h4007007a, 32'h3ef6ec48} /* (6, 15, 12) {real, imag} */,
  {32'hc17e2cc7, 32'h3f520568} /* (6, 15, 11) {real, imag} */,
  {32'h4166b148, 32'h41c13187} /* (6, 15, 10) {real, imag} */,
  {32'hc1e20432, 32'h41a6e910} /* (6, 15, 9) {real, imag} */,
  {32'hc18c7536, 32'hc18ad62c} /* (6, 15, 8) {real, imag} */,
  {32'h412913bc, 32'hc1db9d80} /* (6, 15, 7) {real, imag} */,
  {32'hbfbcc630, 32'h41304fd8} /* (6, 15, 6) {real, imag} */,
  {32'h3ece4060, 32'hc1d04560} /* (6, 15, 5) {real, imag} */,
  {32'hc200d902, 32'h41fba1b1} /* (6, 15, 4) {real, imag} */,
  {32'h4255bdae, 32'h3ffd8510} /* (6, 15, 3) {real, imag} */,
  {32'hbf82b4d8, 32'h40d98412} /* (6, 15, 2) {real, imag} */,
  {32'hc18befaa, 32'hc18a5b20} /* (6, 15, 1) {real, imag} */,
  {32'h424f5c0a, 32'h419a0b2c} /* (6, 15, 0) {real, imag} */,
  {32'hc2530567, 32'hc18f442b} /* (6, 14, 31) {real, imag} */,
  {32'hc082780e, 32'h421c8d8a} /* (6, 14, 30) {real, imag} */,
  {32'hc14755ad, 32'h40a182d8} /* (6, 14, 29) {real, imag} */,
  {32'hbf2b8338, 32'h418e1e4a} /* (6, 14, 28) {real, imag} */,
  {32'hc0c79162, 32'h4162a9a6} /* (6, 14, 27) {real, imag} */,
  {32'hbf168a80, 32'h424053fa} /* (6, 14, 26) {real, imag} */,
  {32'hc114a320, 32'hbff21718} /* (6, 14, 25) {real, imag} */,
  {32'hc20c1a88, 32'hc198bba6} /* (6, 14, 24) {real, imag} */,
  {32'h4142826a, 32'hc191674a} /* (6, 14, 23) {real, imag} */,
  {32'hc126de8a, 32'hc0ab65f4} /* (6, 14, 22) {real, imag} */,
  {32'h40966b12, 32'h41a49049} /* (6, 14, 21) {real, imag} */,
  {32'hc144604e, 32'hc11500d3} /* (6, 14, 20) {real, imag} */,
  {32'hc15545b7, 32'hc0fe6bd0} /* (6, 14, 19) {real, imag} */,
  {32'hc0f98a8e, 32'hc15d6c1e} /* (6, 14, 18) {real, imag} */,
  {32'h403b7110, 32'h40ca9773} /* (6, 14, 17) {real, imag} */,
  {32'hc086c878, 32'h40fde238} /* (6, 14, 16) {real, imag} */,
  {32'hbff103d0, 32'hc0b6cdaf} /* (6, 14, 15) {real, imag} */,
  {32'h413a2095, 32'h40af8b14} /* (6, 14, 14) {real, imag} */,
  {32'hc09780de, 32'h40a6246c} /* (6, 14, 13) {real, imag} */,
  {32'hc0cfca67, 32'h40d9b356} /* (6, 14, 12) {real, imag} */,
  {32'hc0e1c6f2, 32'h40e65a54} /* (6, 14, 11) {real, imag} */,
  {32'h412b32b6, 32'h416597f8} /* (6, 14, 10) {real, imag} */,
  {32'h4175c0a8, 32'h40de9e91} /* (6, 14, 9) {real, imag} */,
  {32'hc08b6284, 32'h4201d4fa} /* (6, 14, 8) {real, imag} */,
  {32'h41264102, 32'hc0eb842c} /* (6, 14, 7) {real, imag} */,
  {32'hc2289127, 32'h41496db8} /* (6, 14, 6) {real, imag} */,
  {32'h41ababf6, 32'h425036d2} /* (6, 14, 5) {real, imag} */,
  {32'hc148379e, 32'h4008b600} /* (6, 14, 4) {real, imag} */,
  {32'h416128bb, 32'hc0d71be4} /* (6, 14, 3) {real, imag} */,
  {32'h41ed8804, 32'h417c1898} /* (6, 14, 2) {real, imag} */,
  {32'hc119fa9c, 32'hc117ba4c} /* (6, 14, 1) {real, imag} */,
  {32'hc22f52d0, 32'h421b6ef3} /* (6, 14, 0) {real, imag} */,
  {32'h42480a73, 32'hc26a39cd} /* (6, 13, 31) {real, imag} */,
  {32'hc099c210, 32'h419d2b86} /* (6, 13, 30) {real, imag} */,
  {32'h4214fe54, 32'hbf9b84a0} /* (6, 13, 29) {real, imag} */,
  {32'h4042d200, 32'hc18364e6} /* (6, 13, 28) {real, imag} */,
  {32'h41a6ac1d, 32'hc1d89cad} /* (6, 13, 27) {real, imag} */,
  {32'hc223ed5e, 32'hc1ad90bc} /* (6, 13, 26) {real, imag} */,
  {32'hbe99ba40, 32'hc13d1eb4} /* (6, 13, 25) {real, imag} */,
  {32'h411249a5, 32'hbfdeb6d0} /* (6, 13, 24) {real, imag} */,
  {32'h40af1335, 32'hc1a47c80} /* (6, 13, 23) {real, imag} */,
  {32'hbf8b7aa0, 32'h4097f196} /* (6, 13, 22) {real, imag} */,
  {32'h41505c16, 32'h41912d59} /* (6, 13, 21) {real, imag} */,
  {32'h40a63700, 32'hc15583ec} /* (6, 13, 20) {real, imag} */,
  {32'hc1a2fb9e, 32'hc0ba56df} /* (6, 13, 19) {real, imag} */,
  {32'h410936e6, 32'h4050a428} /* (6, 13, 18) {real, imag} */,
  {32'h40658608, 32'h3f331ed8} /* (6, 13, 17) {real, imag} */,
  {32'hc0126594, 32'hc12f926c} /* (6, 13, 16) {real, imag} */,
  {32'h4087a8c0, 32'hc153534e} /* (6, 13, 15) {real, imag} */,
  {32'h4122f548, 32'h4210303a} /* (6, 13, 14) {real, imag} */,
  {32'h40d3f4a2, 32'hc12c7f70} /* (6, 13, 13) {real, imag} */,
  {32'hc183a5d3, 32'hc188a9a9} /* (6, 13, 12) {real, imag} */,
  {32'hc0f9cd83, 32'h3faf9830} /* (6, 13, 11) {real, imag} */,
  {32'hbfd68a60, 32'h4197cfca} /* (6, 13, 10) {real, imag} */,
  {32'h40c98e21, 32'hc01b17b0} /* (6, 13, 9) {real, imag} */,
  {32'h4104d511, 32'h41a1e879} /* (6, 13, 8) {real, imag} */,
  {32'hc21d6a50, 32'hc1ee3594} /* (6, 13, 7) {real, imag} */,
  {32'hc16358b6, 32'h420c171c} /* (6, 13, 6) {real, imag} */,
  {32'hc2445918, 32'hc1e7137b} /* (6, 13, 5) {real, imag} */,
  {32'h422d30c2, 32'h40e31ce2} /* (6, 13, 4) {real, imag} */,
  {32'hc21db5dc, 32'hc0c6c256} /* (6, 13, 3) {real, imag} */,
  {32'hc21b61be, 32'hc026cb60} /* (6, 13, 2) {real, imag} */,
  {32'h40c71b38, 32'hc240b519} /* (6, 13, 1) {real, imag} */,
  {32'hc05bdacc, 32'hc18f2b5a} /* (6, 13, 0) {real, imag} */,
  {32'hc201ae65, 32'h40e7e292} /* (6, 12, 31) {real, imag} */,
  {32'hc294b178, 32'hc20df868} /* (6, 12, 30) {real, imag} */,
  {32'hc197c00c, 32'hc08fc7d1} /* (6, 12, 29) {real, imag} */,
  {32'h40125490, 32'h41fa1f57} /* (6, 12, 28) {real, imag} */,
  {32'h41c204d9, 32'h418d0740} /* (6, 12, 27) {real, imag} */,
  {32'h417f7943, 32'hc2287cdd} /* (6, 12, 26) {real, imag} */,
  {32'h41bf89e5, 32'h424ea302} /* (6, 12, 25) {real, imag} */,
  {32'h41a71704, 32'hc1848805} /* (6, 12, 24) {real, imag} */,
  {32'h4199fc12, 32'hc023d712} /* (6, 12, 23) {real, imag} */,
  {32'h41f62828, 32'h415efbc4} /* (6, 12, 22) {real, imag} */,
  {32'hc111ea22, 32'hc05f1a62} /* (6, 12, 21) {real, imag} */,
  {32'h41134b02, 32'h40058276} /* (6, 12, 20) {real, imag} */,
  {32'h41a6c263, 32'h416d98b1} /* (6, 12, 19) {real, imag} */,
  {32'h41085110, 32'h4167cc37} /* (6, 12, 18) {real, imag} */,
  {32'hc0364d4a, 32'h41577c76} /* (6, 12, 17) {real, imag} */,
  {32'hc0ba3c00, 32'h3f548fb0} /* (6, 12, 16) {real, imag} */,
  {32'h3f119a28, 32'h409a3e6c} /* (6, 12, 15) {real, imag} */,
  {32'hc008f010, 32'h3efe9060} /* (6, 12, 14) {real, imag} */,
  {32'h41836dc1, 32'hc11238cf} /* (6, 12, 13) {real, imag} */,
  {32'hc0e4d248, 32'h4112580c} /* (6, 12, 12) {real, imag} */,
  {32'h417cb3fe, 32'h4162cdc0} /* (6, 12, 11) {real, imag} */,
  {32'h40b507be, 32'hc22b9231} /* (6, 12, 10) {real, imag} */,
  {32'h408e3309, 32'hc03e6c2e} /* (6, 12, 9) {real, imag} */,
  {32'hc1152b7c, 32'h3f1270e0} /* (6, 12, 8) {real, imag} */,
  {32'hc1019732, 32'h41fc381c} /* (6, 12, 7) {real, imag} */,
  {32'hc1c7436e, 32'hc1077f7c} /* (6, 12, 6) {real, imag} */,
  {32'h42573e90, 32'h40a3f87e} /* (6, 12, 5) {real, imag} */,
  {32'hc2229ce1, 32'hc1659d6a} /* (6, 12, 4) {real, imag} */,
  {32'hc00ca68c, 32'h3fea9ef4} /* (6, 12, 3) {real, imag} */,
  {32'h4186f4c8, 32'h4102cf7b} /* (6, 12, 2) {real, imag} */,
  {32'hc23da4af, 32'hc164b551} /* (6, 12, 1) {real, imag} */,
  {32'hc20c524c, 32'hc160aa61} /* (6, 12, 0) {real, imag} */,
  {32'h412c10ac, 32'hc2a3ac4a} /* (6, 11, 31) {real, imag} */,
  {32'h415990ee, 32'hc26c1a90} /* (6, 11, 30) {real, imag} */,
  {32'h40ef1ac8, 32'h3fc0e390} /* (6, 11, 29) {real, imag} */,
  {32'hc1807e04, 32'h41e15780} /* (6, 11, 28) {real, imag} */,
  {32'hc2a99b41, 32'hc1c32cfc} /* (6, 11, 27) {real, imag} */,
  {32'h41fac49f, 32'hc2a693f9} /* (6, 11, 26) {real, imag} */,
  {32'hc21a0703, 32'h4233c666} /* (6, 11, 25) {real, imag} */,
  {32'h41ea9d2a, 32'h41f6580e} /* (6, 11, 24) {real, imag} */,
  {32'h416eb5e0, 32'h41943fd0} /* (6, 11, 23) {real, imag} */,
  {32'h413d6020, 32'hc1f7d282} /* (6, 11, 22) {real, imag} */,
  {32'hc2010ecd, 32'hc16612a4} /* (6, 11, 21) {real, imag} */,
  {32'hc172f7a4, 32'h41870d34} /* (6, 11, 20) {real, imag} */,
  {32'h4128e212, 32'hc1004b3e} /* (6, 11, 19) {real, imag} */,
  {32'h40e1f08c, 32'h419c3d74} /* (6, 11, 18) {real, imag} */,
  {32'hc1076944, 32'hc19d52ec} /* (6, 11, 17) {real, imag} */,
  {32'hbff95ce0, 32'h418d1cbf} /* (6, 11, 16) {real, imag} */,
  {32'h41a775f0, 32'hbfa04438} /* (6, 11, 15) {real, imag} */,
  {32'hbf5d0960, 32'h413f1f2d} /* (6, 11, 14) {real, imag} */,
  {32'hc030255e, 32'h419142c9} /* (6, 11, 13) {real, imag} */,
  {32'h415fb4ca, 32'h417167ef} /* (6, 11, 12) {real, imag} */,
  {32'hc0656b20, 32'h4140796e} /* (6, 11, 11) {real, imag} */,
  {32'hc116dd80, 32'hc1855b18} /* (6, 11, 10) {real, imag} */,
  {32'h3fbce820, 32'hc145e589} /* (6, 11, 9) {real, imag} */,
  {32'hc16bc3d9, 32'h4122952d} /* (6, 11, 8) {real, imag} */,
  {32'hc24b8699, 32'hc20f4e66} /* (6, 11, 7) {real, imag} */,
  {32'h41771e02, 32'h41d944ed} /* (6, 11, 6) {real, imag} */,
  {32'h40ed4230, 32'h420da45a} /* (6, 11, 5) {real, imag} */,
  {32'hc2162de4, 32'h4184fd20} /* (6, 11, 4) {real, imag} */,
  {32'h41d893ba, 32'hc263c94c} /* (6, 11, 3) {real, imag} */,
  {32'h4293f748, 32'h4209ceec} /* (6, 11, 2) {real, imag} */,
  {32'hc13e2d48, 32'h4176331c} /* (6, 11, 1) {real, imag} */,
  {32'h422620e7, 32'h4246efc8} /* (6, 11, 0) {real, imag} */,
  {32'hc1d1bff3, 32'h4261965d} /* (6, 10, 31) {real, imag} */,
  {32'h4179cd7f, 32'h41925a4f} /* (6, 10, 30) {real, imag} */,
  {32'hc28cb46a, 32'h41a2f1b2} /* (6, 10, 29) {real, imag} */,
  {32'hc1d3e85c, 32'hc25dd996} /* (6, 10, 28) {real, imag} */,
  {32'hc1c4e156, 32'h426de349} /* (6, 10, 27) {real, imag} */,
  {32'hc209529d, 32'hc19e9736} /* (6, 10, 26) {real, imag} */,
  {32'hc2562338, 32'h41b0ba1b} /* (6, 10, 25) {real, imag} */,
  {32'h3e82ac20, 32'hc20e5d9c} /* (6, 10, 24) {real, imag} */,
  {32'h419eefd4, 32'h41d729a9} /* (6, 10, 23) {real, imag} */,
  {32'h41be711a, 32'h422fc3c4} /* (6, 10, 22) {real, imag} */,
  {32'hc1408108, 32'hc1b450ac} /* (6, 10, 21) {real, imag} */,
  {32'hc112c9b3, 32'hc1bc608c} /* (6, 10, 20) {real, imag} */,
  {32'hc0cd87b8, 32'hc1a019d8} /* (6, 10, 19) {real, imag} */,
  {32'h40d90170, 32'hbe6a7b00} /* (6, 10, 18) {real, imag} */,
  {32'h40f84749, 32'h4204ca97} /* (6, 10, 17) {real, imag} */,
  {32'h40eb98aa, 32'h3f5fbde0} /* (6, 10, 16) {real, imag} */,
  {32'hc04a096e, 32'hc0de6360} /* (6, 10, 15) {real, imag} */,
  {32'hc1d81998, 32'h41952004} /* (6, 10, 14) {real, imag} */,
  {32'h41e96710, 32'h4161270f} /* (6, 10, 13) {real, imag} */,
  {32'hc18f362a, 32'hc1c8c63e} /* (6, 10, 12) {real, imag} */,
  {32'hc237df3a, 32'h420090bf} /* (6, 10, 11) {real, imag} */,
  {32'h41047e84, 32'hc00d3380} /* (6, 10, 10) {real, imag} */,
  {32'hc1797458, 32'hc21bdf7c} /* (6, 10, 9) {real, imag} */,
  {32'h418e80f2, 32'h420a51fc} /* (6, 10, 8) {real, imag} */,
  {32'hc203ced0, 32'h41b511ab} /* (6, 10, 7) {real, imag} */,
  {32'h423c1cdf, 32'h42743f75} /* (6, 10, 6) {real, imag} */,
  {32'h41ab43d6, 32'hc285ec51} /* (6, 10, 5) {real, imag} */,
  {32'h42b8dde9, 32'h41a6b685} /* (6, 10, 4) {real, imag} */,
  {32'hbf42f200, 32'h41e41352} /* (6, 10, 3) {real, imag} */,
  {32'hc0fd86f2, 32'hc03ecd88} /* (6, 10, 2) {real, imag} */,
  {32'h413f051a, 32'h424865cb} /* (6, 10, 1) {real, imag} */,
  {32'h41b9564c, 32'hc24eb4ac} /* (6, 10, 0) {real, imag} */,
  {32'hc2013952, 32'h424eb2f1} /* (6, 9, 31) {real, imag} */,
  {32'hbfaa2900, 32'hc2db4d8a} /* (6, 9, 30) {real, imag} */,
  {32'hc2e81231, 32'h4256c047} /* (6, 9, 29) {real, imag} */,
  {32'hc1953b48, 32'h3ffbc018} /* (6, 9, 28) {real, imag} */,
  {32'h42997bbc, 32'h420fcbfe} /* (6, 9, 27) {real, imag} */,
  {32'h4186d1a8, 32'h4132337d} /* (6, 9, 26) {real, imag} */,
  {32'h4186dc30, 32'h42b06e72} /* (6, 9, 25) {real, imag} */,
  {32'h427475bb, 32'h407229d4} /* (6, 9, 24) {real, imag} */,
  {32'h41a17bc8, 32'hc0f30f50} /* (6, 9, 23) {real, imag} */,
  {32'hc2472b68, 32'hc1488658} /* (6, 9, 22) {real, imag} */,
  {32'h410e042a, 32'hc19af177} /* (6, 9, 21) {real, imag} */,
  {32'hc1aa6fb2, 32'h41d69c70} /* (6, 9, 20) {real, imag} */,
  {32'hc0f3e2eb, 32'hc1b3910c} /* (6, 9, 19) {real, imag} */,
  {32'h4098b2e0, 32'hc11cfbb2} /* (6, 9, 18) {real, imag} */,
  {32'h4131824e, 32'h4153d1fa} /* (6, 9, 17) {real, imag} */,
  {32'h40e27bc2, 32'h408a4090} /* (6, 9, 16) {real, imag} */,
  {32'h41bdb757, 32'h406c07b0} /* (6, 9, 15) {real, imag} */,
  {32'h3edb5300, 32'hc215726e} /* (6, 9, 14) {real, imag} */,
  {32'h41955121, 32'h416ef8e0} /* (6, 9, 13) {real, imag} */,
  {32'h41b400a8, 32'hc0238258} /* (6, 9, 12) {real, imag} */,
  {32'h3fef2eb0, 32'h41ce570b} /* (6, 9, 11) {real, imag} */,
  {32'hc080177c, 32'hc02d89b8} /* (6, 9, 10) {real, imag} */,
  {32'h42952965, 32'hc1c3be68} /* (6, 9, 9) {real, imag} */,
  {32'h41a7b55a, 32'h408e6db6} /* (6, 9, 8) {real, imag} */,
  {32'h42a0191d, 32'hc284e012} /* (6, 9, 7) {real, imag} */,
  {32'h415c0455, 32'h42128d59} /* (6, 9, 6) {real, imag} */,
  {32'h415f4492, 32'h420943a8} /* (6, 9, 5) {real, imag} */,
  {32'hc22905b7, 32'hc2048bff} /* (6, 9, 4) {real, imag} */,
  {32'h42c29c13, 32'h424c7a6f} /* (6, 9, 3) {real, imag} */,
  {32'h42b8a5b3, 32'h409bb5e8} /* (6, 9, 2) {real, imag} */,
  {32'hc183475f, 32'h409c6268} /* (6, 9, 1) {real, imag} */,
  {32'hc0fbbd82, 32'h43395994} /* (6, 9, 0) {real, imag} */,
  {32'h41097408, 32'h428de07e} /* (6, 8, 31) {real, imag} */,
  {32'h426ac824, 32'hc2174136} /* (6, 8, 30) {real, imag} */,
  {32'hc22af958, 32'h42ad91af} /* (6, 8, 29) {real, imag} */,
  {32'hc2963a28, 32'hc2a24dea} /* (6, 8, 28) {real, imag} */,
  {32'hc2b5375e, 32'hc256744e} /* (6, 8, 27) {real, imag} */,
  {32'hc22cb0f4, 32'h42d3964b} /* (6, 8, 26) {real, imag} */,
  {32'hc16f857c, 32'hc2327045} /* (6, 8, 25) {real, imag} */,
  {32'h414953f9, 32'h42572838} /* (6, 8, 24) {real, imag} */,
  {32'h4283870c, 32'hc2a6d8ac} /* (6, 8, 23) {real, imag} */,
  {32'hc1c68ca4, 32'h4202907c} /* (6, 8, 22) {real, imag} */,
  {32'hc19f6622, 32'hc11f5cde} /* (6, 8, 21) {real, imag} */,
  {32'hbfc33be0, 32'hc155d4fc} /* (6, 8, 20) {real, imag} */,
  {32'hc1da6072, 32'hc1df0fce} /* (6, 8, 19) {real, imag} */,
  {32'hc163d5c2, 32'hc0812b64} /* (6, 8, 18) {real, imag} */,
  {32'h412ac0a9, 32'h4125986a} /* (6, 8, 17) {real, imag} */,
  {32'h40a3f5f2, 32'hc11e5361} /* (6, 8, 16) {real, imag} */,
  {32'h3fb26478, 32'hc133f3a2} /* (6, 8, 15) {real, imag} */,
  {32'hc1c68f59, 32'h40397688} /* (6, 8, 14) {real, imag} */,
  {32'hc099d3ea, 32'h4265fe89} /* (6, 8, 13) {real, imag} */,
  {32'h4158dac4, 32'hc2469841} /* (6, 8, 12) {real, imag} */,
  {32'hc13e747b, 32'hc19b7443} /* (6, 8, 11) {real, imag} */,
  {32'hc20c5d71, 32'hc123b456} /* (6, 8, 10) {real, imag} */,
  {32'h41529356, 32'h421755cd} /* (6, 8, 9) {real, imag} */,
  {32'h422c8408, 32'hc24d9504} /* (6, 8, 8) {real, imag} */,
  {32'h425f49a1, 32'hc012c5b0} /* (6, 8, 7) {real, imag} */,
  {32'hc199189e, 32'h4253e1c2} /* (6, 8, 6) {real, imag} */,
  {32'hc281fe04, 32'hc07bac38} /* (6, 8, 5) {real, imag} */,
  {32'hc2e09564, 32'hc1fdcfd2} /* (6, 8, 4) {real, imag} */,
  {32'hc1fc565c, 32'hc28ab0ab} /* (6, 8, 3) {real, imag} */,
  {32'h40b4b8a4, 32'h421f11e6} /* (6, 8, 2) {real, imag} */,
  {32'hc214e660, 32'h42d48b86} /* (6, 8, 1) {real, imag} */,
  {32'h41289979, 32'hc1ad9432} /* (6, 8, 0) {real, imag} */,
  {32'h42284d05, 32'h4319927f} /* (6, 7, 31) {real, imag} */,
  {32'h42d2b656, 32'hc30fa3e3} /* (6, 7, 30) {real, imag} */,
  {32'h425040b6, 32'h4269904e} /* (6, 7, 29) {real, imag} */,
  {32'h42bfbf37, 32'hc1870928} /* (6, 7, 28) {real, imag} */,
  {32'hc2875496, 32'hc2941e70} /* (6, 7, 27) {real, imag} */,
  {32'h412ec9ee, 32'h42aab129} /* (6, 7, 26) {real, imag} */,
  {32'h42f3d8ad, 32'hc188ff2c} /* (6, 7, 25) {real, imag} */,
  {32'hc240aa32, 32'h40293890} /* (6, 7, 24) {real, imag} */,
  {32'hc21eae62, 32'hc0b2f81c} /* (6, 7, 23) {real, imag} */,
  {32'h42170309, 32'h40a8f324} /* (6, 7, 22) {real, imag} */,
  {32'h429055bf, 32'hc149890a} /* (6, 7, 21) {real, imag} */,
  {32'hc1cb8e45, 32'hc192904e} /* (6, 7, 20) {real, imag} */,
  {32'h414c7fd2, 32'h414fb80a} /* (6, 7, 19) {real, imag} */,
  {32'hbf75e780, 32'h4019ccb0} /* (6, 7, 18) {real, imag} */,
  {32'hc256b416, 32'h414376de} /* (6, 7, 17) {real, imag} */,
  {32'h41816112, 32'h41c87ed0} /* (6, 7, 16) {real, imag} */,
  {32'hc2087cb6, 32'hc1f5cd3d} /* (6, 7, 15) {real, imag} */,
  {32'hc1c1ffa4, 32'hc1e6e782} /* (6, 7, 14) {real, imag} */,
  {32'hc203ed54, 32'h3f8fa970} /* (6, 7, 13) {real, imag} */,
  {32'hc215ec18, 32'hc1a3238c} /* (6, 7, 12) {real, imag} */,
  {32'hc23d20d2, 32'hc0a3589c} /* (6, 7, 11) {real, imag} */,
  {32'h4280c76a, 32'hc21d68fa} /* (6, 7, 10) {real, imag} */,
  {32'h4248c47a, 32'hc11b41a6} /* (6, 7, 9) {real, imag} */,
  {32'hc225dd62, 32'hc1ec1a9a} /* (6, 7, 8) {real, imag} */,
  {32'hc04c7820, 32'h40087100} /* (6, 7, 7) {real, imag} */,
  {32'h40e5318c, 32'h41bd8107} /* (6, 7, 6) {real, imag} */,
  {32'hc27779f8, 32'h41455fbc} /* (6, 7, 5) {real, imag} */,
  {32'h433eb0f2, 32'hc20df073} /* (6, 7, 4) {real, imag} */,
  {32'h432ff37a, 32'h42361c5c} /* (6, 7, 3) {real, imag} */,
  {32'hc2ca080a, 32'h426d98b9} /* (6, 7, 2) {real, imag} */,
  {32'h4187725e, 32'hc23f52d4} /* (6, 7, 1) {real, imag} */,
  {32'hc27e4799, 32'hc320e77e} /* (6, 7, 0) {real, imag} */,
  {32'hc1c9df17, 32'hc1c353d1} /* (6, 6, 31) {real, imag} */,
  {32'hc31e4a78, 32'hc2893876} /* (6, 6, 30) {real, imag} */,
  {32'h424b6a2e, 32'hc1a44e2e} /* (6, 6, 29) {real, imag} */,
  {32'h42846d7f, 32'h42c51222} /* (6, 6, 28) {real, imag} */,
  {32'h4284b822, 32'hc29f5801} /* (6, 6, 27) {real, imag} */,
  {32'h417aa350, 32'hc1c292ad} /* (6, 6, 26) {real, imag} */,
  {32'h4256737f, 32'hc227b29c} /* (6, 6, 25) {real, imag} */,
  {32'h41db0eba, 32'h40cc79b8} /* (6, 6, 24) {real, imag} */,
  {32'hc2ab5b8e, 32'h4173e778} /* (6, 6, 23) {real, imag} */,
  {32'h4092b110, 32'h40cef738} /* (6, 6, 22) {real, imag} */,
  {32'h41f15bd2, 32'h41cd33ca} /* (6, 6, 21) {real, imag} */,
  {32'hc225396a, 32'hc280809e} /* (6, 6, 20) {real, imag} */,
  {32'hc07265a8, 32'hc1fae874} /* (6, 6, 19) {real, imag} */,
  {32'hc1120dce, 32'h42533594} /* (6, 6, 18) {real, imag} */,
  {32'h41c2e145, 32'hc12ec0c0} /* (6, 6, 17) {real, imag} */,
  {32'hc0996ee0, 32'h422c2606} /* (6, 6, 16) {real, imag} */,
  {32'hc1a07e4b, 32'h4199a21e} /* (6, 6, 15) {real, imag} */,
  {32'hc145f0fe, 32'h414faf9a} /* (6, 6, 14) {real, imag} */,
  {32'h41c476bf, 32'hc0abd580} /* (6, 6, 13) {real, imag} */,
  {32'h404a72c8, 32'hc14adc4e} /* (6, 6, 12) {real, imag} */,
  {32'hc200b5e7, 32'h409115e6} /* (6, 6, 11) {real, imag} */,
  {32'hc2c0e773, 32'h42b2d320} /* (6, 6, 10) {real, imag} */,
  {32'h42721b14, 32'hc2389764} /* (6, 6, 9) {real, imag} */,
  {32'hc28999fc, 32'hc1fbfb56} /* (6, 6, 8) {real, imag} */,
  {32'h42670961, 32'hc3316e6d} /* (6, 6, 7) {real, imag} */,
  {32'hc1c30c06, 32'h42237c70} /* (6, 6, 6) {real, imag} */,
  {32'hc2064e81, 32'h430739f8} /* (6, 6, 5) {real, imag} */,
  {32'hc25df43e, 32'hc286c054} /* (6, 6, 4) {real, imag} */,
  {32'h41c53223, 32'hc29e151c} /* (6, 6, 3) {real, imag} */,
  {32'h41a51704, 32'h4244e8b0} /* (6, 6, 2) {real, imag} */,
  {32'h42119b48, 32'h425bc8d4} /* (6, 6, 1) {real, imag} */,
  {32'hc1828be5, 32'hc2b96d73} /* (6, 6, 0) {real, imag} */,
  {32'h419b29a8, 32'h42098b82} /* (6, 5, 31) {real, imag} */,
  {32'h42e9e222, 32'h40514020} /* (6, 5, 30) {real, imag} */,
  {32'hc3163404, 32'h428809c8} /* (6, 5, 29) {real, imag} */,
  {32'h40b6f10c, 32'h435146d2} /* (6, 5, 28) {real, imag} */,
  {32'h42087ace, 32'hc2761671} /* (6, 5, 27) {real, imag} */,
  {32'hc242ce9a, 32'h40e1a486} /* (6, 5, 26) {real, imag} */,
  {32'hc2402c61, 32'hc22441e6} /* (6, 5, 25) {real, imag} */,
  {32'hc2a7d867, 32'hc1f1c5a1} /* (6, 5, 24) {real, imag} */,
  {32'hc1efff84, 32'hc2628746} /* (6, 5, 23) {real, imag} */,
  {32'h3de72a00, 32'hc20ca8f0} /* (6, 5, 22) {real, imag} */,
  {32'hc261e69f, 32'hc283a256} /* (6, 5, 21) {real, imag} */,
  {32'h41de92dd, 32'hc22aa107} /* (6, 5, 20) {real, imag} */,
  {32'h3f90d150, 32'hc1532609} /* (6, 5, 19) {real, imag} */,
  {32'h41ad58d7, 32'hc0a0a990} /* (6, 5, 18) {real, imag} */,
  {32'hc0e1bfd8, 32'hc227a95c} /* (6, 5, 17) {real, imag} */,
  {32'hc26ffccb, 32'hc1c2e535} /* (6, 5, 16) {real, imag} */,
  {32'hbe433100, 32'h420c8df0} /* (6, 5, 15) {real, imag} */,
  {32'h40676b38, 32'h41756850} /* (6, 5, 14) {real, imag} */,
  {32'h4234c79a, 32'h418db1dc} /* (6, 5, 13) {real, imag} */,
  {32'hc286df67, 32'hc09dfbb8} /* (6, 5, 12) {real, imag} */,
  {32'h421beab1, 32'h410ebf72} /* (6, 5, 11) {real, imag} */,
  {32'hc292584a, 32'h42295872} /* (6, 5, 10) {real, imag} */,
  {32'hc111ca10, 32'hc2cff635} /* (6, 5, 9) {real, imag} */,
  {32'hc1d8e977, 32'hc11c1c3a} /* (6, 5, 8) {real, imag} */,
  {32'h4243dd9d, 32'h42f12435} /* (6, 5, 7) {real, imag} */,
  {32'h41d6b857, 32'hc073f814} /* (6, 5, 6) {real, imag} */,
  {32'h41bd86ff, 32'hc1b4abe6} /* (6, 5, 5) {real, imag} */,
  {32'h426788e6, 32'h42290fe2} /* (6, 5, 4) {real, imag} */,
  {32'hc16481e8, 32'h3f9b7420} /* (6, 5, 3) {real, imag} */,
  {32'hc2205d04, 32'hc2e86110} /* (6, 5, 2) {real, imag} */,
  {32'h42bfeb8f, 32'hc2c29cdf} /* (6, 5, 1) {real, imag} */,
  {32'hc308eb55, 32'h426885aa} /* (6, 5, 0) {real, imag} */,
  {32'h40877600, 32'h42b81bc7} /* (6, 4, 31) {real, imag} */,
  {32'h400b7010, 32'hc162b146} /* (6, 4, 30) {real, imag} */,
  {32'h419294a8, 32'hc32c0177} /* (6, 4, 29) {real, imag} */,
  {32'hc30159db, 32'h42efa052} /* (6, 4, 28) {real, imag} */,
  {32'h4268e591, 32'hc277ea18} /* (6, 4, 27) {real, imag} */,
  {32'hbf4ce240, 32'hc2f7e02a} /* (6, 4, 26) {real, imag} */,
  {32'hc2b623b0, 32'h420b8f0c} /* (6, 4, 25) {real, imag} */,
  {32'h420ce118, 32'hc20b9304} /* (6, 4, 24) {real, imag} */,
  {32'hc23c6664, 32'h42c2c2ea} /* (6, 4, 23) {real, imag} */,
  {32'h4263207f, 32'h42376048} /* (6, 4, 22) {real, imag} */,
  {32'hc2627cc5, 32'h41c72b6d} /* (6, 4, 21) {real, imag} */,
  {32'h42407ba0, 32'h417f1209} /* (6, 4, 20) {real, imag} */,
  {32'h41ced14d, 32'h424b17da} /* (6, 4, 19) {real, imag} */,
  {32'h40678628, 32'hc05f3918} /* (6, 4, 18) {real, imag} */,
  {32'hc2155fae, 32'hbf766520} /* (6, 4, 17) {real, imag} */,
  {32'h41108dc0, 32'hc1db0863} /* (6, 4, 16) {real, imag} */,
  {32'h40e169d4, 32'h41404662} /* (6, 4, 15) {real, imag} */,
  {32'hbf7ce080, 32'h40174f28} /* (6, 4, 14) {real, imag} */,
  {32'hc1075ba6, 32'hc1064e4a} /* (6, 4, 13) {real, imag} */,
  {32'hc1b8ec48, 32'h40808ce2} /* (6, 4, 12) {real, imag} */,
  {32'h421351d7, 32'h41423576} /* (6, 4, 11) {real, imag} */,
  {32'h42589a55, 32'hc19d4a88} /* (6, 4, 10) {real, imag} */,
  {32'hc2e5606c, 32'h4257b180} /* (6, 4, 9) {real, imag} */,
  {32'hc285cb5a, 32'h411fda22} /* (6, 4, 8) {real, imag} */,
  {32'hc2a0f24e, 32'hc0079110} /* (6, 4, 7) {real, imag} */,
  {32'h41eac780, 32'hc241e630} /* (6, 4, 6) {real, imag} */,
  {32'h41c54052, 32'h425d93d8} /* (6, 4, 5) {real, imag} */,
  {32'h4239e960, 32'hc28ea0ea} /* (6, 4, 4) {real, imag} */,
  {32'hc2ab4e68, 32'hc331afff} /* (6, 4, 3) {real, imag} */,
  {32'hc22ac43d, 32'h42579d14} /* (6, 4, 2) {real, imag} */,
  {32'h42dd784e, 32'h42254986} /* (6, 4, 1) {real, imag} */,
  {32'h42c38022, 32'hc228419a} /* (6, 4, 0) {real, imag} */,
  {32'h42444c7b, 32'h43237084} /* (6, 3, 31) {real, imag} */,
  {32'h428e4d50, 32'hc28bd5e0} /* (6, 3, 30) {real, imag} */,
  {32'h41b41e92, 32'h41e243ef} /* (6, 3, 29) {real, imag} */,
  {32'h41c9e5ff, 32'h4218fe28} /* (6, 3, 28) {real, imag} */,
  {32'hc0f58ca4, 32'hc21440b0} /* (6, 3, 27) {real, imag} */,
  {32'h420c531e, 32'h42a6fc22} /* (6, 3, 26) {real, imag} */,
  {32'h41017fc0, 32'hc2c1df84} /* (6, 3, 25) {real, imag} */,
  {32'h411356de, 32'hc061f910} /* (6, 3, 24) {real, imag} */,
  {32'h420fba3e, 32'hc2833de6} /* (6, 3, 23) {real, imag} */,
  {32'h41228590, 32'hc2c42d18} /* (6, 3, 22) {real, imag} */,
  {32'h423e5436, 32'h42db04fa} /* (6, 3, 21) {real, imag} */,
  {32'hc20db5dc, 32'h4140d1e4} /* (6, 3, 20) {real, imag} */,
  {32'h41fcfa3e, 32'h41075b22} /* (6, 3, 19) {real, imag} */,
  {32'hc013fb68, 32'hc1eb94bd} /* (6, 3, 18) {real, imag} */,
  {32'h4111c86f, 32'h41a6aac6} /* (6, 3, 17) {real, imag} */,
  {32'h4229e246, 32'h41ec15e5} /* (6, 3, 16) {real, imag} */,
  {32'hbf3e6df0, 32'h41869516} /* (6, 3, 15) {real, imag} */,
  {32'h41682d7a, 32'hc261ff0e} /* (6, 3, 14) {real, imag} */,
  {32'h40082330, 32'hc16df6fa} /* (6, 3, 13) {real, imag} */,
  {32'hc226fb8c, 32'hc11103da} /* (6, 3, 12) {real, imag} */,
  {32'hbfb72950, 32'hc229f424} /* (6, 3, 11) {real, imag} */,
  {32'hbfdc4f5c, 32'hc1619944} /* (6, 3, 10) {real, imag} */,
  {32'hc1a38678, 32'hc18d467b} /* (6, 3, 9) {real, imag} */,
  {32'hc213ab2a, 32'hc1166848} /* (6, 3, 8) {real, imag} */,
  {32'hc213abc2, 32'hc1b5b836} /* (6, 3, 7) {real, imag} */,
  {32'hc22e6112, 32'h41690934} /* (6, 3, 6) {real, imag} */,
  {32'h41ac4fd3, 32'hc32ebce2} /* (6, 3, 5) {real, imag} */,
  {32'h426b347c, 32'hc19a20dd} /* (6, 3, 4) {real, imag} */,
  {32'hc309090d, 32'h4290bfdc} /* (6, 3, 3) {real, imag} */,
  {32'h42c676c8, 32'h40af4f60} /* (6, 3, 2) {real, imag} */,
  {32'h42ebc970, 32'hc2e98624} /* (6, 3, 1) {real, imag} */,
  {32'hc229a806, 32'h42b0b47b} /* (6, 3, 0) {real, imag} */,
  {32'h43af149e, 32'h418bba5a} /* (6, 2, 31) {real, imag} */,
  {32'h42540cc7, 32'hc1ab0530} /* (6, 2, 30) {real, imag} */,
  {32'hc2d45f46, 32'hc1d27284} /* (6, 2, 29) {real, imag} */,
  {32'hc2c387e4, 32'hc316fa48} /* (6, 2, 28) {real, imag} */,
  {32'hc25ee3ba, 32'h42afa5e0} /* (6, 2, 27) {real, imag} */,
  {32'hc2b5e7be, 32'h416ad552} /* (6, 2, 26) {real, imag} */,
  {32'h42f2b610, 32'hc196b6aa} /* (6, 2, 25) {real, imag} */,
  {32'hc2e3ccfb, 32'h42ccca32} /* (6, 2, 24) {real, imag} */,
  {32'hc0ec1490, 32'h42b8577a} /* (6, 2, 23) {real, imag} */,
  {32'h3f906708, 32'hc284a5ad} /* (6, 2, 22) {real, imag} */,
  {32'hc18c666b, 32'hc291750e} /* (6, 2, 21) {real, imag} */,
  {32'h40c59928, 32'h422d6ecc} /* (6, 2, 20) {real, imag} */,
  {32'h418ed2f0, 32'hc13ae314} /* (6, 2, 19) {real, imag} */,
  {32'hc08c10ae, 32'h4101c624} /* (6, 2, 18) {real, imag} */,
  {32'h413eaec8, 32'hc018e8bc} /* (6, 2, 17) {real, imag} */,
  {32'h41411802, 32'h4172c070} /* (6, 2, 16) {real, imag} */,
  {32'h3f8cde40, 32'h416c059f} /* (6, 2, 15) {real, imag} */,
  {32'h40429c24, 32'hc1eb8254} /* (6, 2, 14) {real, imag} */,
  {32'hc0e98a01, 32'h416e7bac} /* (6, 2, 13) {real, imag} */,
  {32'hc1d0bde6, 32'h423891a2} /* (6, 2, 12) {real, imag} */,
  {32'hbfb02790, 32'h4136d754} /* (6, 2, 11) {real, imag} */,
  {32'hc18f947c, 32'hc1a6a17d} /* (6, 2, 10) {real, imag} */,
  {32'hc2531c96, 32'hbf3db9c0} /* (6, 2, 9) {real, imag} */,
  {32'h42977da9, 32'h42246654} /* (6, 2, 8) {real, imag} */,
  {32'hc27dec04, 32'h4292f83c} /* (6, 2, 7) {real, imag} */,
  {32'h4281c4de, 32'h428a2b50} /* (6, 2, 6) {real, imag} */,
  {32'hc2cfb777, 32'h428e1df0} /* (6, 2, 5) {real, imag} */,
  {32'h419e7310, 32'h429ee298} /* (6, 2, 4) {real, imag} */,
  {32'h42dac500, 32'hc2e76ad3} /* (6, 2, 3) {real, imag} */,
  {32'hc26c4dd5, 32'hc2d1db66} /* (6, 2, 2) {real, imag} */,
  {32'hc2d26b99, 32'h423c7acf} /* (6, 2, 1) {real, imag} */,
  {32'hc28e0b78, 32'hc3175ed3} /* (6, 2, 0) {real, imag} */,
  {32'hc23ff09e, 32'hc22c33c1} /* (6, 1, 31) {real, imag} */,
  {32'hc1e23970, 32'hc26c1f83} /* (6, 1, 30) {real, imag} */,
  {32'hc214c978, 32'hc2eb21c4} /* (6, 1, 29) {real, imag} */,
  {32'h42f408bc, 32'h42e1420f} /* (6, 1, 28) {real, imag} */,
  {32'h417a47fd, 32'hc1110fbe} /* (6, 1, 27) {real, imag} */,
  {32'h42933236, 32'hc249d34d} /* (6, 1, 26) {real, imag} */,
  {32'hc1eef420, 32'hc0a76024} /* (6, 1, 25) {real, imag} */,
  {32'hc009d408, 32'hc2d2c038} /* (6, 1, 24) {real, imag} */,
  {32'hc2917c3c, 32'hc2853760} /* (6, 1, 23) {real, imag} */,
  {32'h42aad628, 32'h41caea08} /* (6, 1, 22) {real, imag} */,
  {32'hc26d79a0, 32'h4102faf6} /* (6, 1, 21) {real, imag} */,
  {32'h42311a0c, 32'h4297b78c} /* (6, 1, 20) {real, imag} */,
  {32'hc155981d, 32'h418289aa} /* (6, 1, 19) {real, imag} */,
  {32'h42852a29, 32'h41771c68} /* (6, 1, 18) {real, imag} */,
  {32'h418658ec, 32'h41098775} /* (6, 1, 17) {real, imag} */,
  {32'hc1d5eaa0, 32'h3daa9600} /* (6, 1, 16) {real, imag} */,
  {32'h41921392, 32'h414ed93d} /* (6, 1, 15) {real, imag} */,
  {32'h3ff499c0, 32'hc28fe486} /* (6, 1, 14) {real, imag} */,
  {32'hc1bde8de, 32'h42bb54ba} /* (6, 1, 13) {real, imag} */,
  {32'hc21d42c4, 32'hc2007c40} /* (6, 1, 12) {real, imag} */,
  {32'hc215eb68, 32'h41befa81} /* (6, 1, 11) {real, imag} */,
  {32'hc11ca024, 32'hc198d40c} /* (6, 1, 10) {real, imag} */,
  {32'h3fe99ca0, 32'h40d8961c} /* (6, 1, 9) {real, imag} */,
  {32'hc2416d4a, 32'h40475e70} /* (6, 1, 8) {real, imag} */,
  {32'hc272f64e, 32'hc16471c2} /* (6, 1, 7) {real, imag} */,
  {32'hc23c03d2, 32'hc1e5cf5e} /* (6, 1, 6) {real, imag} */,
  {32'h422c7d79, 32'h41aff4bb} /* (6, 1, 5) {real, imag} */,
  {32'h42aff948, 32'h413c3748} /* (6, 1, 4) {real, imag} */,
  {32'hc225668a, 32'h421376d9} /* (6, 1, 3) {real, imag} */,
  {32'hc2e3f0d6, 32'h42191e73} /* (6, 1, 2) {real, imag} */,
  {32'h4260623a, 32'h42447569} /* (6, 1, 1) {real, imag} */,
  {32'h43122fee, 32'hc2e849be} /* (6, 1, 0) {real, imag} */,
  {32'h41765170, 32'h43033c94} /* (6, 0, 31) {real, imag} */,
  {32'hc31994a6, 32'hc19f5cf8} /* (6, 0, 30) {real, imag} */,
  {32'h406c0b08, 32'h3fa35f10} /* (6, 0, 29) {real, imag} */,
  {32'hc1ede04a, 32'hc2cf0dfb} /* (6, 0, 28) {real, imag} */,
  {32'h42f2124e, 32'h43668418} /* (6, 0, 27) {real, imag} */,
  {32'h40ad4b82, 32'h4245f82a} /* (6, 0, 26) {real, imag} */,
  {32'h4216a6b1, 32'hc228c00e} /* (6, 0, 25) {real, imag} */,
  {32'hc1d6dc20, 32'hc3042b3b} /* (6, 0, 24) {real, imag} */,
  {32'hc23b7fa3, 32'h41bdcd57} /* (6, 0, 23) {real, imag} */,
  {32'h4238e124, 32'h422cb708} /* (6, 0, 22) {real, imag} */,
  {32'hc18fe117, 32'hc14143fc} /* (6, 0, 21) {real, imag} */,
  {32'h41ac2b19, 32'h40ec76c0} /* (6, 0, 20) {real, imag} */,
  {32'h41720f14, 32'h41e8650e} /* (6, 0, 19) {real, imag} */,
  {32'hc20b356e, 32'h4095610c} /* (6, 0, 18) {real, imag} */,
  {32'hc21ef45a, 32'h40b98b44} /* (6, 0, 17) {real, imag} */,
  {32'hc12f5960, 32'h42413338} /* (6, 0, 16) {real, imag} */,
  {32'hc13c41e9, 32'hc158cf82} /* (6, 0, 15) {real, imag} */,
  {32'h41eb8440, 32'h425a9b0a} /* (6, 0, 14) {real, imag} */,
  {32'hc28754ee, 32'hc21f5bf5} /* (6, 0, 13) {real, imag} */,
  {32'h411a783a, 32'hc21c3bf8} /* (6, 0, 12) {real, imag} */,
  {32'h417d39d2, 32'hc2992cf0} /* (6, 0, 11) {real, imag} */,
  {32'hc1edf7b0, 32'hc282d82a} /* (6, 0, 10) {real, imag} */,
  {32'hc1cdb552, 32'hc20ef86e} /* (6, 0, 9) {real, imag} */,
  {32'hc200407b, 32'hc1b1c3d6} /* (6, 0, 8) {real, imag} */,
  {32'h430f513c, 32'hc28418f9} /* (6, 0, 7) {real, imag} */,
  {32'hc16fcdc3, 32'h4237dc02} /* (6, 0, 6) {real, imag} */,
  {32'hc2206d6c, 32'hc2c191f8} /* (6, 0, 5) {real, imag} */,
  {32'hc28643ce, 32'hc2e9fe29} /* (6, 0, 4) {real, imag} */,
  {32'h40bb580c, 32'h4248509a} /* (6, 0, 3) {real, imag} */,
  {32'h43032f8c, 32'h43190e1a} /* (6, 0, 2) {real, imag} */,
  {32'h42a2d7b4, 32'h41da6e2c} /* (6, 0, 1) {real, imag} */,
  {32'h43269c08, 32'h43154c58} /* (6, 0, 0) {real, imag} */,
  {32'h416c05a0, 32'hc41e81ae} /* (5, 31, 31) {real, imag} */,
  {32'h43403fe4, 32'h43bd6940} /* (5, 31, 30) {real, imag} */,
  {32'hbf7aaca0, 32'h4362b010} /* (5, 31, 29) {real, imag} */,
  {32'hc1fcd254, 32'hc2b1f187} /* (5, 31, 28) {real, imag} */,
  {32'hc21abb4c, 32'h426dbd5b} /* (5, 31, 27) {real, imag} */,
  {32'h42b75f92, 32'h401f574a} /* (5, 31, 26) {real, imag} */,
  {32'h42bb9bb1, 32'hc2e08685} /* (5, 31, 25) {real, imag} */,
  {32'h420257e9, 32'h434eb418} /* (5, 31, 24) {real, imag} */,
  {32'hc1b1b013, 32'h4250c456} /* (5, 31, 23) {real, imag} */,
  {32'h40b726d6, 32'h41082ca2} /* (5, 31, 22) {real, imag} */,
  {32'hc11f606c, 32'h428f8c80} /* (5, 31, 21) {real, imag} */,
  {32'h41810b3e, 32'hc173e7e0} /* (5, 31, 20) {real, imag} */,
  {32'h421604a0, 32'hc2159cdc} /* (5, 31, 19) {real, imag} */,
  {32'h420f734e, 32'hc264c6da} /* (5, 31, 18) {real, imag} */,
  {32'hc1a7155c, 32'h422e4da2} /* (5, 31, 17) {real, imag} */,
  {32'h41bd6c58, 32'hc120dca0} /* (5, 31, 16) {real, imag} */,
  {32'h40820010, 32'h41f3b11c} /* (5, 31, 15) {real, imag} */,
  {32'h408597ac, 32'h4216732a} /* (5, 31, 14) {real, imag} */,
  {32'h41252162, 32'h41403bb0} /* (5, 31, 13) {real, imag} */,
  {32'hc174d0bc, 32'hc24da9c6} /* (5, 31, 12) {real, imag} */,
  {32'hc209fb35, 32'h4099c858} /* (5, 31, 11) {real, imag} */,
  {32'h418fc7e6, 32'hc117f8aa} /* (5, 31, 10) {real, imag} */,
  {32'hc19226db, 32'hc09ae570} /* (5, 31, 9) {real, imag} */,
  {32'hc2d25e04, 32'h425e7b18} /* (5, 31, 8) {real, imag} */,
  {32'hc1813d64, 32'hc33d4310} /* (5, 31, 7) {real, imag} */,
  {32'hc2378eed, 32'h3c58d600} /* (5, 31, 6) {real, imag} */,
  {32'hc3744681, 32'h43074182} /* (5, 31, 5) {real, imag} */,
  {32'h42dde68b, 32'hc095fb40} /* (5, 31, 4) {real, imag} */,
  {32'h425d397e, 32'hc22007ea} /* (5, 31, 3) {real, imag} */,
  {32'hc3086fde, 32'h430a2284} /* (5, 31, 2) {real, imag} */,
  {32'h43f060e9, 32'hc39f2673} /* (5, 31, 1) {real, imag} */,
  {32'h4324ff25, 32'hc405c81c} /* (5, 31, 0) {real, imag} */,
  {32'hc32cca40, 32'h43adf63e} /* (5, 30, 31) {real, imag} */,
  {32'h436d2e56, 32'hc3bd57a2} /* (5, 30, 30) {real, imag} */,
  {32'h41415538, 32'hc18b3b8a} /* (5, 30, 29) {real, imag} */,
  {32'hc25c2912, 32'h43036a50} /* (5, 30, 28) {real, imag} */,
  {32'hc2aa3c02, 32'hc3342666} /* (5, 30, 27) {real, imag} */,
  {32'h42ae94ba, 32'h429f0c2a} /* (5, 30, 26) {real, imag} */,
  {32'hc2904ed7, 32'h4245db4a} /* (5, 30, 25) {real, imag} */,
  {32'h417951a0, 32'h429701fa} /* (5, 30, 24) {real, imag} */,
  {32'hc224c0fa, 32'h41e36db2} /* (5, 30, 23) {real, imag} */,
  {32'h42017588, 32'h41ca96e2} /* (5, 30, 22) {real, imag} */,
  {32'hc101b790, 32'h3ff7e270} /* (5, 30, 21) {real, imag} */,
  {32'hbfb35b20, 32'h41822f56} /* (5, 30, 20) {real, imag} */,
  {32'hc201a987, 32'hc09c07dc} /* (5, 30, 19) {real, imag} */,
  {32'h423f1e55, 32'hc249b884} /* (5, 30, 18) {real, imag} */,
  {32'h415a2988, 32'h40cdeed0} /* (5, 30, 17) {real, imag} */,
  {32'h412b3344, 32'h41abb700} /* (5, 30, 16) {real, imag} */,
  {32'hc1822974, 32'hc216859a} /* (5, 30, 15) {real, imag} */,
  {32'h4192076e, 32'h4211aaf4} /* (5, 30, 14) {real, imag} */,
  {32'h40ce7328, 32'h421a37aa} /* (5, 30, 13) {real, imag} */,
  {32'h419586b6, 32'hc088a9b8} /* (5, 30, 12) {real, imag} */,
  {32'h420f8866, 32'h42516900} /* (5, 30, 11) {real, imag} */,
  {32'h41beff79, 32'h40ce1330} /* (5, 30, 10) {real, imag} */,
  {32'h42d92ae5, 32'h428c3b64} /* (5, 30, 9) {real, imag} */,
  {32'h43056d15, 32'h3fd109a0} /* (5, 30, 8) {real, imag} */,
  {32'hc32af61c, 32'hc2353dbc} /* (5, 30, 7) {real, imag} */,
  {32'h43249a2a, 32'hc1cc0767} /* (5, 30, 6) {real, imag} */,
  {32'h4288c4be, 32'hc1ec2dfc} /* (5, 30, 5) {real, imag} */,
  {32'hc336f44c, 32'h41fb52a2} /* (5, 30, 4) {real, imag} */,
  {32'hc33ce760, 32'h4306cc46} /* (5, 30, 3) {real, imag} */,
  {32'h433bdbe6, 32'hc387a5d4} /* (5, 30, 2) {real, imag} */,
  {32'hc3c6580c, 32'h43eb8fac} /* (5, 30, 1) {real, imag} */,
  {32'h42a57824, 32'h43f147f2} /* (5, 30, 0) {real, imag} */,
  {32'hc28aed16, 32'hc2f8f5f3} /* (5, 29, 31) {real, imag} */,
  {32'h43001353, 32'h42cf5c0d} /* (5, 29, 30) {real, imag} */,
  {32'h41262e60, 32'h4109d284} /* (5, 29, 29) {real, imag} */,
  {32'hc2a78ec3, 32'hc18d736a} /* (5, 29, 28) {real, imag} */,
  {32'hc1167d68, 32'hc2c09aa1} /* (5, 29, 27) {real, imag} */,
  {32'h43047121, 32'h430d7ca5} /* (5, 29, 26) {real, imag} */,
  {32'hc28990cb, 32'hc3205fca} /* (5, 29, 25) {real, imag} */,
  {32'hc24aef9c, 32'h428d20bb} /* (5, 29, 24) {real, imag} */,
  {32'hc0f7ada0, 32'h42da3f0a} /* (5, 29, 23) {real, imag} */,
  {32'hc20024a7, 32'h41a5c3f5} /* (5, 29, 22) {real, imag} */,
  {32'h410fe4d6, 32'hc1a07a6c} /* (5, 29, 21) {real, imag} */,
  {32'h41ebc1b8, 32'hc2a6b640} /* (5, 29, 20) {real, imag} */,
  {32'hbffe7aa8, 32'h420399d5} /* (5, 29, 19) {real, imag} */,
  {32'hc21daa88, 32'h4197254e} /* (5, 29, 18) {real, imag} */,
  {32'hc1e977a0, 32'h41d2c9a3} /* (5, 29, 17) {real, imag} */,
  {32'hc1534500, 32'hc1918a8c} /* (5, 29, 16) {real, imag} */,
  {32'h42084600, 32'hc106d35a} /* (5, 29, 15) {real, imag} */,
  {32'h4226dc80, 32'h41cd5ace} /* (5, 29, 14) {real, imag} */,
  {32'h41ef00fc, 32'hc2253cf1} /* (5, 29, 13) {real, imag} */,
  {32'hc22dbb70, 32'h41491614} /* (5, 29, 12) {real, imag} */,
  {32'h4029f148, 32'hc18cdc68} /* (5, 29, 11) {real, imag} */,
  {32'hc2b74aa4, 32'hc2390bd8} /* (5, 29, 10) {real, imag} */,
  {32'h42bd1a46, 32'hc16c2044} /* (5, 29, 9) {real, imag} */,
  {32'h42b3bb84, 32'h431b80f4} /* (5, 29, 8) {real, imag} */,
  {32'h422d30ba, 32'h4289c2c6} /* (5, 29, 7) {real, imag} */,
  {32'hc2c7d4fa, 32'hc228472c} /* (5, 29, 6) {real, imag} */,
  {32'hc2b02f43, 32'h42fb630f} /* (5, 29, 5) {real, imag} */,
  {32'h42d843f7, 32'hc2ed8a2c} /* (5, 29, 4) {real, imag} */,
  {32'h428aff1e, 32'h420bd3f9} /* (5, 29, 3) {real, imag} */,
  {32'h4360a5ef, 32'hc2dad565} /* (5, 29, 2) {real, imag} */,
  {32'hc3955e5a, 32'h427a46da} /* (5, 29, 1) {real, imag} */,
  {32'h42fe71f2, 32'hc3127e04} /* (5, 29, 0) {real, imag} */,
  {32'hc0151840, 32'hc38f4d38} /* (5, 28, 31) {real, imag} */,
  {32'hc303df64, 32'h4353003e} /* (5, 28, 30) {real, imag} */,
  {32'hc238f45e, 32'h42b3c671} /* (5, 28, 29) {real, imag} */,
  {32'hc0baa148, 32'hc21eed78} /* (5, 28, 28) {real, imag} */,
  {32'h426b421c, 32'h42688192} /* (5, 28, 27) {real, imag} */,
  {32'h418a7d73, 32'hc31bf20a} /* (5, 28, 26) {real, imag} */,
  {32'h41b9f53d, 32'h3f9ca760} /* (5, 28, 25) {real, imag} */,
  {32'h4167d100, 32'hc1e6e4c5} /* (5, 28, 24) {real, imag} */,
  {32'h42815194, 32'hc215cf26} /* (5, 28, 23) {real, imag} */,
  {32'hc27de46e, 32'h3fe13490} /* (5, 28, 22) {real, imag} */,
  {32'hc218b2ea, 32'hc1df2051} /* (5, 28, 21) {real, imag} */,
  {32'h3f8e2ab8, 32'hc1c2fdfe} /* (5, 28, 20) {real, imag} */,
  {32'h4180a853, 32'hbf9a40c0} /* (5, 28, 19) {real, imag} */,
  {32'hc106e7ac, 32'h425f0068} /* (5, 28, 18) {real, imag} */,
  {32'hc1868660, 32'h42192c00} /* (5, 28, 17) {real, imag} */,
  {32'h416e2d9c, 32'hc2218666} /* (5, 28, 16) {real, imag} */,
  {32'h422a10e8, 32'h3f456600} /* (5, 28, 15) {real, imag} */,
  {32'hc18fdad2, 32'hc13d3ee0} /* (5, 28, 14) {real, imag} */,
  {32'hc140ac96, 32'h4224a900} /* (5, 28, 13) {real, imag} */,
  {32'hc1f19ab0, 32'h418e5bc2} /* (5, 28, 12) {real, imag} */,
  {32'h3f9c7ae0, 32'hc0e11ae4} /* (5, 28, 11) {real, imag} */,
  {32'h4295c1fd, 32'hc21efad6} /* (5, 28, 10) {real, imag} */,
  {32'hc1b50152, 32'h4293be70} /* (5, 28, 9) {real, imag} */,
  {32'hc2a70200, 32'h429b1048} /* (5, 28, 8) {real, imag} */,
  {32'h41a06e97, 32'hc297e94a} /* (5, 28, 7) {real, imag} */,
  {32'hc284d238, 32'h42934035} /* (5, 28, 6) {real, imag} */,
  {32'hc1583ec2, 32'h42395a6e} /* (5, 28, 5) {real, imag} */,
  {32'hc28147fe, 32'hc31dcaba} /* (5, 28, 4) {real, imag} */,
  {32'h41d0a523, 32'h42e9ffbf} /* (5, 28, 3) {real, imag} */,
  {32'h42d3e678, 32'h42e34fec} /* (5, 28, 2) {real, imag} */,
  {32'hc340c2b3, 32'hc2e0cabd} /* (5, 28, 1) {real, imag} */,
  {32'h427d5679, 32'h4306af4e} /* (5, 28, 0) {real, imag} */,
  {32'hc370a6ff, 32'h43443386} /* (5, 27, 31) {real, imag} */,
  {32'hc1e5a9e8, 32'hc281f73a} /* (5, 27, 30) {real, imag} */,
  {32'h42137f6a, 32'h41a86d46} /* (5, 27, 29) {real, imag} */,
  {32'h41097efe, 32'h41940334} /* (5, 27, 28) {real, imag} */,
  {32'h42755a28, 32'hc2c39152} /* (5, 27, 27) {real, imag} */,
  {32'hc1689fc0, 32'hc2f63d12} /* (5, 27, 26) {real, imag} */,
  {32'h42398e6e, 32'h42591f58} /* (5, 27, 25) {real, imag} */,
  {32'hc16f0a8c, 32'h42c3169a} /* (5, 27, 24) {real, imag} */,
  {32'h41db6c82, 32'hc219163c} /* (5, 27, 23) {real, imag} */,
  {32'h423ccd13, 32'hc2933232} /* (5, 27, 22) {real, imag} */,
  {32'h412d6664, 32'hbce24c00} /* (5, 27, 21) {real, imag} */,
  {32'h424d52c2, 32'h428c7dce} /* (5, 27, 20) {real, imag} */,
  {32'h4080a13c, 32'hc20598ad} /* (5, 27, 19) {real, imag} */,
  {32'hc212cde6, 32'h40923948} /* (5, 27, 18) {real, imag} */,
  {32'hc1af52aa, 32'h3f58c7b8} /* (5, 27, 17) {real, imag} */,
  {32'h41f5e250, 32'h41a4bed0} /* (5, 27, 16) {real, imag} */,
  {32'h41828b46, 32'hc12c13cc} /* (5, 27, 15) {real, imag} */,
  {32'h41e1b198, 32'hc209cec5} /* (5, 27, 14) {real, imag} */,
  {32'h416b246e, 32'h40ec4c98} /* (5, 27, 13) {real, imag} */,
  {32'h420ca000, 32'h41823d8c} /* (5, 27, 12) {real, imag} */,
  {32'h41092884, 32'hc136533a} /* (5, 27, 11) {real, imag} */,
  {32'h4185b29c, 32'hc0eab918} /* (5, 27, 10) {real, imag} */,
  {32'hc27b881f, 32'hc1e98b43} /* (5, 27, 9) {real, imag} */,
  {32'hc1c10a2a, 32'h40660930} /* (5, 27, 8) {real, imag} */,
  {32'hc14cdc82, 32'h42a246dc} /* (5, 27, 7) {real, imag} */,
  {32'h4222bde3, 32'h425e7e1c} /* (5, 27, 6) {real, imag} */,
  {32'h430e3698, 32'h41c34550} /* (5, 27, 5) {real, imag} */,
  {32'hc124d726, 32'hc2619df8} /* (5, 27, 4) {real, imag} */,
  {32'hc3017d2a, 32'hc2e33386} /* (5, 27, 3) {real, imag} */,
  {32'h43320891, 32'hc320e1c0} /* (5, 27, 2) {real, imag} */,
  {32'h4287507e, 32'h4331a3aa} /* (5, 27, 1) {real, imag} */,
  {32'hc2e78040, 32'h42838146} /* (5, 27, 0) {real, imag} */,
  {32'hc30a64fb, 32'h423e21f4} /* (5, 26, 31) {real, imag} */,
  {32'h418609e2, 32'hbf1b73a0} /* (5, 26, 30) {real, imag} */,
  {32'h422ccc02, 32'hc2321e9c} /* (5, 26, 29) {real, imag} */,
  {32'hc2148a32, 32'h423693e0} /* (5, 26, 28) {real, imag} */,
  {32'h41aafabc, 32'h42e093ed} /* (5, 26, 27) {real, imag} */,
  {32'h4211c384, 32'h42bf80a0} /* (5, 26, 26) {real, imag} */,
  {32'hc1fb28aa, 32'h42879ca7} /* (5, 26, 25) {real, imag} */,
  {32'h42a86614, 32'hc3076c94} /* (5, 26, 24) {real, imag} */,
  {32'hc2c8b871, 32'hc0638dc8} /* (5, 26, 23) {real, imag} */,
  {32'hc0c8fbc0, 32'hc194f2e7} /* (5, 26, 22) {real, imag} */,
  {32'h424647ee, 32'hc1eca200} /* (5, 26, 21) {real, imag} */,
  {32'hc22e00b4, 32'h419d33f0} /* (5, 26, 20) {real, imag} */,
  {32'h3f5b19a0, 32'h417824da} /* (5, 26, 19) {real, imag} */,
  {32'hc1743bce, 32'h4253dd84} /* (5, 26, 18) {real, imag} */,
  {32'h41e4cd49, 32'hc1eaf739} /* (5, 26, 17) {real, imag} */,
  {32'h41303d9c, 32'h41384968} /* (5, 26, 16) {real, imag} */,
  {32'hc1c09ee9, 32'h41e251c1} /* (5, 26, 15) {real, imag} */,
  {32'hc0e09c94, 32'h4158bb20} /* (5, 26, 14) {real, imag} */,
  {32'h41965251, 32'h4192e5e1} /* (5, 26, 13) {real, imag} */,
  {32'h41a27b3c, 32'h40b2fb9f} /* (5, 26, 12) {real, imag} */,
  {32'hc1b4fb3c, 32'hc0137af0} /* (5, 26, 11) {real, imag} */,
  {32'h42b416d6, 32'hc1c1a6db} /* (5, 26, 10) {real, imag} */,
  {32'hc233db96, 32'hbff336f0} /* (5, 26, 9) {real, imag} */,
  {32'hc1cc40c6, 32'h41ce200e} /* (5, 26, 8) {real, imag} */,
  {32'h423342fd, 32'h42d536d7} /* (5, 26, 7) {real, imag} */,
  {32'h42a5fd80, 32'hc28cebd4} /* (5, 26, 6) {real, imag} */,
  {32'h433e7806, 32'hc1b52e24} /* (5, 26, 5) {real, imag} */,
  {32'h428f12d2, 32'h40f2e1c0} /* (5, 26, 4) {real, imag} */,
  {32'hc3001eaa, 32'h413a0ffa} /* (5, 26, 3) {real, imag} */,
  {32'hc291e5b2, 32'hc188b289} /* (5, 26, 2) {real, imag} */,
  {32'hc31b1ff5, 32'h42d742e8} /* (5, 26, 1) {real, imag} */,
  {32'h42004719, 32'h43166abc} /* (5, 26, 0) {real, imag} */,
  {32'hc228d8b8, 32'hc2e6b882} /* (5, 25, 31) {real, imag} */,
  {32'h430cea6a, 32'h42b22532} /* (5, 25, 30) {real, imag} */,
  {32'h424c9cdc, 32'hc29271d6} /* (5, 25, 29) {real, imag} */,
  {32'h42357c21, 32'h425c9e4e} /* (5, 25, 28) {real, imag} */,
  {32'h419452b7, 32'hc266e760} /* (5, 25, 27) {real, imag} */,
  {32'hc2100202, 32'h41324d8e} /* (5, 25, 26) {real, imag} */,
  {32'hc26e15f0, 32'h40563b5c} /* (5, 25, 25) {real, imag} */,
  {32'h41f3a273, 32'h41e7f7f3} /* (5, 25, 24) {real, imag} */,
  {32'h3e1347c0, 32'h40c16a76} /* (5, 25, 23) {real, imag} */,
  {32'hc16c7ef8, 32'h3f2a83a0} /* (5, 25, 22) {real, imag} */,
  {32'hc1432538, 32'h42347a9b} /* (5, 25, 21) {real, imag} */,
  {32'h41e09c88, 32'h41be8ee5} /* (5, 25, 20) {real, imag} */,
  {32'h41a9c2aa, 32'hc0443268} /* (5, 25, 19) {real, imag} */,
  {32'h41d18a32, 32'hc198470e} /* (5, 25, 18) {real, imag} */,
  {32'h41ab41db, 32'hc1e7dcb6} /* (5, 25, 17) {real, imag} */,
  {32'hc25c2296, 32'hc001b7c0} /* (5, 25, 16) {real, imag} */,
  {32'h3f405320, 32'hc20d756f} /* (5, 25, 15) {real, imag} */,
  {32'h405966f4, 32'h3e58a300} /* (5, 25, 14) {real, imag} */,
  {32'hc1a2ced2, 32'hc23b36fe} /* (5, 25, 13) {real, imag} */,
  {32'h4210ca0c, 32'hc20fe470} /* (5, 25, 12) {real, imag} */,
  {32'h4226787a, 32'h4272fb4b} /* (5, 25, 11) {real, imag} */,
  {32'hc112b758, 32'hc1dd2e79} /* (5, 25, 10) {real, imag} */,
  {32'h4197a494, 32'h41ff7110} /* (5, 25, 9) {real, imag} */,
  {32'h42989889, 32'h41b52b65} /* (5, 25, 8) {real, imag} */,
  {32'hc27efa9a, 32'h41af7956} /* (5, 25, 7) {real, imag} */,
  {32'hc25bd20e, 32'h40e0b2d4} /* (5, 25, 6) {real, imag} */,
  {32'hbe15d280, 32'h42641f60} /* (5, 25, 5) {real, imag} */,
  {32'hc1a3ad9a, 32'hc28afa08} /* (5, 25, 4) {real, imag} */,
  {32'h4283e204, 32'h4282c90a} /* (5, 25, 3) {real, imag} */,
  {32'h43155144, 32'h41666c74} /* (5, 25, 2) {real, imag} */,
  {32'h414cfe84, 32'h42a16e56} /* (5, 25, 1) {real, imag} */,
  {32'hc25ef592, 32'hc2dcaba8} /* (5, 25, 0) {real, imag} */,
  {32'hc0d6d278, 32'h40c7d1c0} /* (5, 24, 31) {real, imag} */,
  {32'h4241da96, 32'hc267b0cd} /* (5, 24, 30) {real, imag} */,
  {32'hc28c506e, 32'hc2b94b86} /* (5, 24, 29) {real, imag} */,
  {32'hc27b1a59, 32'h41d53a1e} /* (5, 24, 28) {real, imag} */,
  {32'hc1fcf01e, 32'h41918a88} /* (5, 24, 27) {real, imag} */,
  {32'h429fd6b6, 32'h42a558ac} /* (5, 24, 26) {real, imag} */,
  {32'hc288fa1f, 32'hbf76aa20} /* (5, 24, 25) {real, imag} */,
  {32'hc20ed91e, 32'hc1ac073d} /* (5, 24, 24) {real, imag} */,
  {32'hc2078337, 32'h4212c20b} /* (5, 24, 23) {real, imag} */,
  {32'hc2982b3e, 32'h4281ed6b} /* (5, 24, 22) {real, imag} */,
  {32'h42aa02fa, 32'hc1aade94} /* (5, 24, 21) {real, imag} */,
  {32'h420805b5, 32'h41f8ee35} /* (5, 24, 20) {real, imag} */,
  {32'h4117b219, 32'h411df366} /* (5, 24, 19) {real, imag} */,
  {32'hc0063386, 32'h40d44f1a} /* (5, 24, 18) {real, imag} */,
  {32'h41da320f, 32'h41140ed8} /* (5, 24, 17) {real, imag} */,
  {32'hc1c0bf92, 32'hc03b8520} /* (5, 24, 16) {real, imag} */,
  {32'hc175e20e, 32'hc0afdc20} /* (5, 24, 15) {real, imag} */,
  {32'hc0e64d93, 32'h411a9acb} /* (5, 24, 14) {real, imag} */,
  {32'h418b3e10, 32'hc188f1ed} /* (5, 24, 13) {real, imag} */,
  {32'hc2155c5f, 32'h4198f36b} /* (5, 24, 12) {real, imag} */,
  {32'hbfa7fce0, 32'h4135cbb5} /* (5, 24, 11) {real, imag} */,
  {32'hc0e83cc8, 32'hc1d6e28c} /* (5, 24, 10) {real, imag} */,
  {32'h4239ac79, 32'hc17a644f} /* (5, 24, 9) {real, imag} */,
  {32'h42d707e1, 32'hc2703d62} /* (5, 24, 8) {real, imag} */,
  {32'hc0bc94dc, 32'h420735da} /* (5, 24, 7) {real, imag} */,
  {32'hc1775a0c, 32'hc243788c} /* (5, 24, 6) {real, imag} */,
  {32'h42da7af8, 32'h41d93c40} /* (5, 24, 5) {real, imag} */,
  {32'hc2ad7dfc, 32'hc28fa744} /* (5, 24, 4) {real, imag} */,
  {32'h4312ab17, 32'hc1d46e00} /* (5, 24, 3) {real, imag} */,
  {32'hc1b265a1, 32'hc2aba9de} /* (5, 24, 2) {real, imag} */,
  {32'h421afb32, 32'h4344cd78} /* (5, 24, 1) {real, imag} */,
  {32'h4153d1f0, 32'h42da59b5} /* (5, 24, 0) {real, imag} */,
  {32'h41295400, 32'h3f3b6e40} /* (5, 23, 31) {real, imag} */,
  {32'hc1b15afe, 32'hc282eec6} /* (5, 23, 30) {real, imag} */,
  {32'hc1874c51, 32'h42d960be} /* (5, 23, 29) {real, imag} */,
  {32'hc2a38f21, 32'hc13768a8} /* (5, 23, 28) {real, imag} */,
  {32'h42d34d3c, 32'hc2893c01} /* (5, 23, 27) {real, imag} */,
  {32'h4190f4b9, 32'h423af000} /* (5, 23, 26) {real, imag} */,
  {32'hc2151514, 32'h41aacfac} /* (5, 23, 25) {real, imag} */,
  {32'hc1e4bd9b, 32'h417c9af6} /* (5, 23, 24) {real, imag} */,
  {32'hc1c449e6, 32'hc22cead6} /* (5, 23, 23) {real, imag} */,
  {32'hc0468c20, 32'h4176d026} /* (5, 23, 22) {real, imag} */,
  {32'hc0b69df8, 32'hc27e49c6} /* (5, 23, 21) {real, imag} */,
  {32'hc1a8c23a, 32'hc0c20d70} /* (5, 23, 20) {real, imag} */,
  {32'h41dc11be, 32'hc15e106a} /* (5, 23, 19) {real, imag} */,
  {32'h41a0f378, 32'h4104da26} /* (5, 23, 18) {real, imag} */,
  {32'hc0c16780, 32'h41b35102} /* (5, 23, 17) {real, imag} */,
  {32'hc2600372, 32'hc13695ee} /* (5, 23, 16) {real, imag} */,
  {32'h42500a7e, 32'hc140a10b} /* (5, 23, 15) {real, imag} */,
  {32'hc10cd778, 32'h40eef115} /* (5, 23, 14) {real, imag} */,
  {32'h4135a5a0, 32'hc171ee6a} /* (5, 23, 13) {real, imag} */,
  {32'h418177b6, 32'hc0e19748} /* (5, 23, 12) {real, imag} */,
  {32'hc23592da, 32'h41ea8a98} /* (5, 23, 11) {real, imag} */,
  {32'h4156cd5c, 32'hc089a28c} /* (5, 23, 10) {real, imag} */,
  {32'h424240bb, 32'hc1e430c4} /* (5, 23, 9) {real, imag} */,
  {32'h41bbff75, 32'h42228d56} /* (5, 23, 8) {real, imag} */,
  {32'h4251041a, 32'hc240c4c2} /* (5, 23, 7) {real, imag} */,
  {32'hc29965fc, 32'h42bfe2d4} /* (5, 23, 6) {real, imag} */,
  {32'hc1788e70, 32'h42a43a7b} /* (5, 23, 5) {real, imag} */,
  {32'hc2535846, 32'h42c884b1} /* (5, 23, 4) {real, imag} */,
  {32'h42814634, 32'hc0a02580} /* (5, 23, 3) {real, imag} */,
  {32'h42268b19, 32'hc2b31e5c} /* (5, 23, 2) {real, imag} */,
  {32'hc23fb772, 32'hc25dd7bb} /* (5, 23, 1) {real, imag} */,
  {32'hc18047cc, 32'hc1813c0b} /* (5, 23, 0) {real, imag} */,
  {32'h42c3a8e9, 32'hc29d4a72} /* (5, 22, 31) {real, imag} */,
  {32'hc29ec0b2, 32'h42a35c64} /* (5, 22, 30) {real, imag} */,
  {32'hc2a261e3, 32'hc2c7b439} /* (5, 22, 29) {real, imag} */,
  {32'hc195b5f2, 32'hc252f9e3} /* (5, 22, 28) {real, imag} */,
  {32'h41ac3770, 32'h418831ad} /* (5, 22, 27) {real, imag} */,
  {32'hc28f926c, 32'h4167ab24} /* (5, 22, 26) {real, imag} */,
  {32'h42a44b78, 32'hc216436c} /* (5, 22, 25) {real, imag} */,
  {32'hc12e06cf, 32'h4229de50} /* (5, 22, 24) {real, imag} */,
  {32'h41143e76, 32'hbfd1c660} /* (5, 22, 23) {real, imag} */,
  {32'hc067f488, 32'hc0d79028} /* (5, 22, 22) {real, imag} */,
  {32'h41d27a33, 32'h41872c4a} /* (5, 22, 21) {real, imag} */,
  {32'hc22bc93e, 32'h41085c10} /* (5, 22, 20) {real, imag} */,
  {32'h41a33a69, 32'h40cd5610} /* (5, 22, 19) {real, imag} */,
  {32'h40db2ce0, 32'hc04a6210} /* (5, 22, 18) {real, imag} */,
  {32'h3e03d000, 32'hc15ebe66} /* (5, 22, 17) {real, imag} */,
  {32'hbfb886f0, 32'hc098b3e0} /* (5, 22, 16) {real, imag} */,
  {32'h4137e060, 32'h41ed3151} /* (5, 22, 15) {real, imag} */,
  {32'hc0508ac0, 32'h408b00b0} /* (5, 22, 14) {real, imag} */,
  {32'h3fd4fcb0, 32'hc1526390} /* (5, 22, 13) {real, imag} */,
  {32'h41316b03, 32'hc138d334} /* (5, 22, 12) {real, imag} */,
  {32'hc012b140, 32'hc217fec2} /* (5, 22, 11) {real, imag} */,
  {32'h42258418, 32'h41f6ac0a} /* (5, 22, 10) {real, imag} */,
  {32'hc17d6b16, 32'hc20d9c0b} /* (5, 22, 9) {real, imag} */,
  {32'hc2158f5d, 32'hc1829078} /* (5, 22, 8) {real, imag} */,
  {32'h41f0b1c7, 32'h424c2358} /* (5, 22, 7) {real, imag} */,
  {32'hc1efcb06, 32'h4078b072} /* (5, 22, 6) {real, imag} */,
  {32'h4274999a, 32'h417ea65e} /* (5, 22, 5) {real, imag} */,
  {32'h4224ff5e, 32'h42063f81} /* (5, 22, 4) {real, imag} */,
  {32'hc22f0380, 32'h4184f5d0} /* (5, 22, 3) {real, imag} */,
  {32'hc08bc6f8, 32'h4219e14c} /* (5, 22, 2) {real, imag} */,
  {32'hc2a0e4b3, 32'hc22d7689} /* (5, 22, 1) {real, imag} */,
  {32'hc243d364, 32'hc287d7dd} /* (5, 22, 0) {real, imag} */,
  {32'h42034e15, 32'h4033d090} /* (5, 21, 31) {real, imag} */,
  {32'hc1d73ea6, 32'h42250068} /* (5, 21, 30) {real, imag} */,
  {32'h41cd5280, 32'h41f64f6d} /* (5, 21, 29) {real, imag} */,
  {32'h42dfb864, 32'h413596a8} /* (5, 21, 28) {real, imag} */,
  {32'hc2372034, 32'h4160bce0} /* (5, 21, 27) {real, imag} */,
  {32'h418e77f2, 32'hbf163d70} /* (5, 21, 26) {real, imag} */,
  {32'h4136632a, 32'h3fe86260} /* (5, 21, 25) {real, imag} */,
  {32'hc184f04e, 32'hc0d95326} /* (5, 21, 24) {real, imag} */,
  {32'h40b00e35, 32'h42222a24} /* (5, 21, 23) {real, imag} */,
  {32'hc22bb352, 32'h422dc3ba} /* (5, 21, 22) {real, imag} */,
  {32'h40b0a2b8, 32'h41e9f294} /* (5, 21, 21) {real, imag} */,
  {32'hc1c01e28, 32'hc00f1f9c} /* (5, 21, 20) {real, imag} */,
  {32'hc1327272, 32'h41c7516e} /* (5, 21, 19) {real, imag} */,
  {32'hc1131ae8, 32'hc1955686} /* (5, 21, 18) {real, imag} */,
  {32'hc0c48b3d, 32'hc19cb6da} /* (5, 21, 17) {real, imag} */,
  {32'hbf9d8d00, 32'h41b20dfa} /* (5, 21, 16) {real, imag} */,
  {32'hc11a0f62, 32'h3e9c7fe0} /* (5, 21, 15) {real, imag} */,
  {32'h41d16aec, 32'hc13148d4} /* (5, 21, 14) {real, imag} */,
  {32'h41d13bf3, 32'h417fd8dc} /* (5, 21, 13) {real, imag} */,
  {32'h409a71b2, 32'hbfbc46e8} /* (5, 21, 12) {real, imag} */,
  {32'h41378fcc, 32'hc1aa9380} /* (5, 21, 11) {real, imag} */,
  {32'hc110ea18, 32'hc0c1ecdc} /* (5, 21, 10) {real, imag} */,
  {32'h4171e8d0, 32'hc1cf5aeb} /* (5, 21, 9) {real, imag} */,
  {32'hbf973328, 32'hc20c67e1} /* (5, 21, 8) {real, imag} */,
  {32'h3f2c0288, 32'h42a6ce54} /* (5, 21, 7) {real, imag} */,
  {32'hc03642ec, 32'hc18095b8} /* (5, 21, 6) {real, imag} */,
  {32'hc1bdb58d, 32'hc2b170a3} /* (5, 21, 5) {real, imag} */,
  {32'hc1e77460, 32'h42682b8e} /* (5, 21, 4) {real, imag} */,
  {32'h41a4d93e, 32'h4106740e} /* (5, 21, 3) {real, imag} */,
  {32'hc1489a30, 32'h41e59765} /* (5, 21, 2) {real, imag} */,
  {32'hbf9efe60, 32'h429d6962} /* (5, 21, 1) {real, imag} */,
  {32'h41c8f1b3, 32'h42b0baaa} /* (5, 21, 0) {real, imag} */,
  {32'h422ac6d8, 32'hc22c003a} /* (5, 20, 31) {real, imag} */,
  {32'h4137ae95, 32'hc1fca544} /* (5, 20, 30) {real, imag} */,
  {32'hc1a9c614, 32'h4135fd83} /* (5, 20, 29) {real, imag} */,
  {32'h423f5e01, 32'hc2033124} /* (5, 20, 28) {real, imag} */,
  {32'hc25b8076, 32'hc23a1ef3} /* (5, 20, 27) {real, imag} */,
  {32'hc25f70d1, 32'h3d24f100} /* (5, 20, 26) {real, imag} */,
  {32'h3e9cdc20, 32'h40839458} /* (5, 20, 25) {real, imag} */,
  {32'h4182676a, 32'h4119ddfb} /* (5, 20, 24) {real, imag} */,
  {32'hc13cde58, 32'hc20f4c95} /* (5, 20, 23) {real, imag} */,
  {32'h411ee774, 32'hc20de55b} /* (5, 20, 22) {real, imag} */,
  {32'hc080d81a, 32'hc130f0fa} /* (5, 20, 21) {real, imag} */,
  {32'h412a01d3, 32'h41dcdc62} /* (5, 20, 20) {real, imag} */,
  {32'hc119c6c8, 32'hc00e3650} /* (5, 20, 19) {real, imag} */,
  {32'hc0279a3c, 32'h408e1fe2} /* (5, 20, 18) {real, imag} */,
  {32'h40791d36, 32'hc0a40d00} /* (5, 20, 17) {real, imag} */,
  {32'h409afc9c, 32'h40f323c4} /* (5, 20, 16) {real, imag} */,
  {32'hc12dad96, 32'hc11ad150} /* (5, 20, 15) {real, imag} */,
  {32'hc18654a4, 32'h40de997e} /* (5, 20, 14) {real, imag} */,
  {32'hc1976583, 32'hc08c4ea4} /* (5, 20, 13) {real, imag} */,
  {32'h401190cc, 32'h3e72b980} /* (5, 20, 12) {real, imag} */,
  {32'h418c88de, 32'hc19c4d8c} /* (5, 20, 11) {real, imag} */,
  {32'hc1703634, 32'hc18609d8} /* (5, 20, 10) {real, imag} */,
  {32'h42311b64, 32'hc19410ca} /* (5, 20, 9) {real, imag} */,
  {32'hc0c68c4a, 32'h410142cb} /* (5, 20, 8) {real, imag} */,
  {32'h40f02eee, 32'hc26de3d5} /* (5, 20, 7) {real, imag} */,
  {32'h422e4839, 32'h41672653} /* (5, 20, 6) {real, imag} */,
  {32'hc1980a6d, 32'hc215433d} /* (5, 20, 5) {real, imag} */,
  {32'hc29ff198, 32'h4267f0e4} /* (5, 20, 4) {real, imag} */,
  {32'h4222ef4a, 32'h41c0fd9a} /* (5, 20, 3) {real, imag} */,
  {32'hc0a03d16, 32'h40c57970} /* (5, 20, 2) {real, imag} */,
  {32'h41ab26b3, 32'hc22df8a6} /* (5, 20, 1) {real, imag} */,
  {32'h4239fd00, 32'hc1bfd97c} /* (5, 20, 0) {real, imag} */,
  {32'hc10b0af9, 32'hc0d25bf0} /* (5, 19, 31) {real, imag} */,
  {32'h418ebc06, 32'h41f4a9ea} /* (5, 19, 30) {real, imag} */,
  {32'hc2000af0, 32'hc1b8a0e5} /* (5, 19, 29) {real, imag} */,
  {32'hc20cca6e, 32'hc1015664} /* (5, 19, 28) {real, imag} */,
  {32'h41fa98e1, 32'hc1badc3e} /* (5, 19, 27) {real, imag} */,
  {32'hc1e4d8f7, 32'h419985b2} /* (5, 19, 26) {real, imag} */,
  {32'h423ea288, 32'hc21f04f5} /* (5, 19, 25) {real, imag} */,
  {32'h40d15ed0, 32'hbf300ec0} /* (5, 19, 24) {real, imag} */,
  {32'h417ec856, 32'hc2139c2e} /* (5, 19, 23) {real, imag} */,
  {32'h410d00be, 32'h4104f360} /* (5, 19, 22) {real, imag} */,
  {32'h41ccd305, 32'hc1934924} /* (5, 19, 21) {real, imag} */,
  {32'hc06aba3e, 32'hc009c59e} /* (5, 19, 20) {real, imag} */,
  {32'h4065a85c, 32'h4114474a} /* (5, 19, 19) {real, imag} */,
  {32'hc1120456, 32'h40396cee} /* (5, 19, 18) {real, imag} */,
  {32'hc06a4150, 32'h415ba4df} /* (5, 19, 17) {real, imag} */,
  {32'h4154af20, 32'hc0e4fac2} /* (5, 19, 16) {real, imag} */,
  {32'hc121ab96, 32'hc0be0252} /* (5, 19, 15) {real, imag} */,
  {32'h40436a5a, 32'h41227c04} /* (5, 19, 14) {real, imag} */,
  {32'h407d0bc4, 32'h419562d1} /* (5, 19, 13) {real, imag} */,
  {32'hc043e89e, 32'h4172e542} /* (5, 19, 12) {real, imag} */,
  {32'hc199ff5b, 32'h40302474} /* (5, 19, 11) {real, imag} */,
  {32'h41e4293b, 32'hc1678a76} /* (5, 19, 10) {real, imag} */,
  {32'hc1c0be85, 32'h41c1eaac} /* (5, 19, 9) {real, imag} */,
  {32'hc204192e, 32'hc141a90c} /* (5, 19, 8) {real, imag} */,
  {32'hc1467a1a, 32'h419c30ae} /* (5, 19, 7) {real, imag} */,
  {32'h40f2226c, 32'hc03d473c} /* (5, 19, 6) {real, imag} */,
  {32'hc2a36170, 32'hc1735890} /* (5, 19, 5) {real, imag} */,
  {32'h42696148, 32'h40e75d83} /* (5, 19, 4) {real, imag} */,
  {32'hc22229b8, 32'h407a81f8} /* (5, 19, 3) {real, imag} */,
  {32'h413fa9cd, 32'hc1729d78} /* (5, 19, 2) {real, imag} */,
  {32'h42080834, 32'hc1713f5a} /* (5, 19, 1) {real, imag} */,
  {32'hc234e37c, 32'hc04f699c} /* (5, 19, 0) {real, imag} */,
  {32'hc103a35c, 32'hc19d35d1} /* (5, 18, 31) {real, imag} */,
  {32'h3e96ab80, 32'h42961075} /* (5, 18, 30) {real, imag} */,
  {32'h41ce82e7, 32'hc284162e} /* (5, 18, 29) {real, imag} */,
  {32'hc11a7875, 32'hc1407624} /* (5, 18, 28) {real, imag} */,
  {32'h41fb5b2b, 32'hbe242720} /* (5, 18, 27) {real, imag} */,
  {32'h410074bd, 32'h40f1ee7c} /* (5, 18, 26) {real, imag} */,
  {32'h417ed071, 32'hc0cb7ac6} /* (5, 18, 25) {real, imag} */,
  {32'hc101cc2c, 32'h3f0cafb0} /* (5, 18, 24) {real, imag} */,
  {32'hc1f4c7fc, 32'h410e4a67} /* (5, 18, 23) {real, imag} */,
  {32'h42260c27, 32'hc1c5315d} /* (5, 18, 22) {real, imag} */,
  {32'h4168ef17, 32'h40e7bb01} /* (5, 18, 21) {real, imag} */,
  {32'h40d4a77c, 32'hc1d83d38} /* (5, 18, 20) {real, imag} */,
  {32'h4112b06e, 32'h409166ec} /* (5, 18, 19) {real, imag} */,
  {32'hc04918dc, 32'h40328958} /* (5, 18, 18) {real, imag} */,
  {32'h40f53763, 32'hc14e3cbc} /* (5, 18, 17) {real, imag} */,
  {32'hc0699f72, 32'hbfa4c778} /* (5, 18, 16) {real, imag} */,
  {32'h407a342e, 32'h40a08620} /* (5, 18, 15) {real, imag} */,
  {32'hc0f72706, 32'hc04ce638} /* (5, 18, 14) {real, imag} */,
  {32'h40f470a7, 32'hc1186616} /* (5, 18, 13) {real, imag} */,
  {32'h40a8ea5e, 32'hc1b11ece} /* (5, 18, 12) {real, imag} */,
  {32'h4131a0d1, 32'hbe2ff160} /* (5, 18, 11) {real, imag} */,
  {32'h41160a3c, 32'h421503bf} /* (5, 18, 10) {real, imag} */,
  {32'h410a6fd5, 32'h40f6ab62} /* (5, 18, 9) {real, imag} */,
  {32'hc1a51eac, 32'h41df73b4} /* (5, 18, 8) {real, imag} */,
  {32'hc2209ff9, 32'hc181354a} /* (5, 18, 7) {real, imag} */,
  {32'h421c1709, 32'hc22ea242} /* (5, 18, 6) {real, imag} */,
  {32'hc10eb16a, 32'hc0659e4a} /* (5, 18, 5) {real, imag} */,
  {32'hc1778a13, 32'hc27b9a17} /* (5, 18, 4) {real, imag} */,
  {32'h414c5552, 32'hc16a758e} /* (5, 18, 3) {real, imag} */,
  {32'hc19aa6bd, 32'hc20aa28e} /* (5, 18, 2) {real, imag} */,
  {32'hbf5f2358, 32'h428a24e4} /* (5, 18, 1) {real, imag} */,
  {32'h40d3c717, 32'h41bf5986} /* (5, 18, 0) {real, imag} */,
  {32'hbfc2b4e0, 32'hc238746a} /* (5, 17, 31) {real, imag} */,
  {32'hc144fa32, 32'hc2024792} /* (5, 17, 30) {real, imag} */,
  {32'h4119e4a5, 32'h3fec6e2a} /* (5, 17, 29) {real, imag} */,
  {32'hc1d85aca, 32'h41916f54} /* (5, 17, 28) {real, imag} */,
  {32'h42893b5c, 32'h40543f65} /* (5, 17, 27) {real, imag} */,
  {32'hc1acb186, 32'h42184b0e} /* (5, 17, 26) {real, imag} */,
  {32'hc1dd6cd8, 32'hc0dd4599} /* (5, 17, 25) {real, imag} */,
  {32'h41e40cb8, 32'hc107d9d8} /* (5, 17, 24) {real, imag} */,
  {32'hc10d2972, 32'h41399f30} /* (5, 17, 23) {real, imag} */,
  {32'h4124ce02, 32'hc0f60bec} /* (5, 17, 22) {real, imag} */,
  {32'h403084a0, 32'hc1b1e54a} /* (5, 17, 21) {real, imag} */,
  {32'hbf5b8078, 32'h40ff717e} /* (5, 17, 20) {real, imag} */,
  {32'h40bdda0c, 32'hbeb755c0} /* (5, 17, 19) {real, imag} */,
  {32'hc085b550, 32'h3dd7f380} /* (5, 17, 18) {real, imag} */,
  {32'hc02d9a4c, 32'hc0463598} /* (5, 17, 17) {real, imag} */,
  {32'h4118497a, 32'hc0dbc5d0} /* (5, 17, 16) {real, imag} */,
  {32'h3f8ce238, 32'h3eeba5c0} /* (5, 17, 15) {real, imag} */,
  {32'hc1477736, 32'h416a0e03} /* (5, 17, 14) {real, imag} */,
  {32'hc03d958d, 32'h412a5e7c} /* (5, 17, 13) {real, imag} */,
  {32'hc11b0c50, 32'h4087addc} /* (5, 17, 12) {real, imag} */,
  {32'h409817a8, 32'h3f386db0} /* (5, 17, 11) {real, imag} */,
  {32'hc15b06c4, 32'h411ae462} /* (5, 17, 10) {real, imag} */,
  {32'hc151f81e, 32'hc120b66c} /* (5, 17, 9) {real, imag} */,
  {32'h3e5afdc0, 32'h3f6d5460} /* (5, 17, 8) {real, imag} */,
  {32'hc1b88880, 32'hc11284cc} /* (5, 17, 7) {real, imag} */,
  {32'hc09c3052, 32'h41c72f6e} /* (5, 17, 6) {real, imag} */,
  {32'h3fe31780, 32'h408f0dc2} /* (5, 17, 5) {real, imag} */,
  {32'h40d01288, 32'hc1602bac} /* (5, 17, 4) {real, imag} */,
  {32'hc141c98b, 32'h410849e5} /* (5, 17, 3) {real, imag} */,
  {32'hc042ec1a, 32'h4183531a} /* (5, 17, 2) {real, imag} */,
  {32'hc2385235, 32'h408be574} /* (5, 17, 1) {real, imag} */,
  {32'h3f336c58, 32'hc1196b2a} /* (5, 17, 0) {real, imag} */,
  {32'h3fc732d8, 32'h416da2f2} /* (5, 16, 31) {real, imag} */,
  {32'h3ac3c000, 32'h403679c8} /* (5, 16, 30) {real, imag} */,
  {32'h40894628, 32'hc1ee4633} /* (5, 16, 29) {real, imag} */,
  {32'hc1849f0a, 32'h41e059b0} /* (5, 16, 28) {real, imag} */,
  {32'h3f95d467, 32'h41a87dc3} /* (5, 16, 27) {real, imag} */,
  {32'h4070f3fa, 32'hbfff73ca} /* (5, 16, 26) {real, imag} */,
  {32'h410b222c, 32'hc0576712} /* (5, 16, 25) {real, imag} */,
  {32'hc0146068, 32'h42237d60} /* (5, 16, 24) {real, imag} */,
  {32'hbf42dd60, 32'h3f925908} /* (5, 16, 23) {real, imag} */,
  {32'h4158893e, 32'hc14d014a} /* (5, 16, 22) {real, imag} */,
  {32'hc1088114, 32'hc10e9a0a} /* (5, 16, 21) {real, imag} */,
  {32'hc1f16725, 32'h4107737a} /* (5, 16, 20) {real, imag} */,
  {32'hc19668a2, 32'hbf8246c8} /* (5, 16, 19) {real, imag} */,
  {32'h4043b950, 32'h4032b9a4} /* (5, 16, 18) {real, imag} */,
  {32'h405f9a74, 32'h3e125da0} /* (5, 16, 17) {real, imag} */,
  {32'hc0ab79e8, 32'hc12f2dcd} /* (5, 16, 16) {real, imag} */,
  {32'hbe59b240, 32'hc0c3f829} /* (5, 16, 15) {real, imag} */,
  {32'hc09101fc, 32'h40fe2742} /* (5, 16, 14) {real, imag} */,
  {32'h40d2e928, 32'h4021528c} /* (5, 16, 13) {real, imag} */,
  {32'h40af7b6c, 32'h3f995a34} /* (5, 16, 12) {real, imag} */,
  {32'h4160a14c, 32'hc11af68e} /* (5, 16, 11) {real, imag} */,
  {32'hc0b96cf9, 32'hc171a1f8} /* (5, 16, 10) {real, imag} */,
  {32'h419f9ca3, 32'h41bdea5a} /* (5, 16, 9) {real, imag} */,
  {32'h41074b54, 32'hc11cc9b2} /* (5, 16, 8) {real, imag} */,
  {32'h414a93f0, 32'h41394ea6} /* (5, 16, 7) {real, imag} */,
  {32'hc170de74, 32'h405bfffd} /* (5, 16, 6) {real, imag} */,
  {32'hbfa1ebd9, 32'h407550c8} /* (5, 16, 5) {real, imag} */,
  {32'h40d374e2, 32'hc0f658e8} /* (5, 16, 4) {real, imag} */,
  {32'hc08ae172, 32'h42029d88} /* (5, 16, 3) {real, imag} */,
  {32'hc1b59cc8, 32'hc19d03d6} /* (5, 16, 2) {real, imag} */,
  {32'hc1be37e6, 32'h41a1c1cb} /* (5, 16, 1) {real, imag} */,
  {32'h417d0344, 32'h3dcb1c80} /* (5, 16, 0) {real, imag} */,
  {32'hc16017bc, 32'hc13022eb} /* (5, 15, 31) {real, imag} */,
  {32'hc0e3285e, 32'h4293c4a2} /* (5, 15, 30) {real, imag} */,
  {32'h3e8db3b0, 32'hc09eee26} /* (5, 15, 29) {real, imag} */,
  {32'hc10b8a43, 32'hc14ee416} /* (5, 15, 28) {real, imag} */,
  {32'hc224cf7a, 32'h41477ec0} /* (5, 15, 27) {real, imag} */,
  {32'hc07f051e, 32'h416f0443} /* (5, 15, 26) {real, imag} */,
  {32'hc1d33275, 32'hc0dca238} /* (5, 15, 25) {real, imag} */,
  {32'hc20a5fd8, 32'hc05752c8} /* (5, 15, 24) {real, imag} */,
  {32'h4135db4a, 32'h3fc34082} /* (5, 15, 23) {real, imag} */,
  {32'h416aec7e, 32'h418be0c6} /* (5, 15, 22) {real, imag} */,
  {32'h402f8754, 32'hc0765b92} /* (5, 15, 21) {real, imag} */,
  {32'h409bceb4, 32'hbf3875b0} /* (5, 15, 20) {real, imag} */,
  {32'hc1571246, 32'hc0cefd05} /* (5, 15, 19) {real, imag} */,
  {32'hc1253cfa, 32'hbf4fd5f0} /* (5, 15, 18) {real, imag} */,
  {32'h4116b1ff, 32'hc0f4090e} /* (5, 15, 17) {real, imag} */,
  {32'hc0f2cef8, 32'h4166e9f8} /* (5, 15, 16) {real, imag} */,
  {32'h409884aa, 32'h40a6dd98} /* (5, 15, 15) {real, imag} */,
  {32'h3fa56e80, 32'h4122d969} /* (5, 15, 14) {real, imag} */,
  {32'h40d1ea71, 32'h411e48ca} /* (5, 15, 13) {real, imag} */,
  {32'hc080f7e2, 32'h41ac8568} /* (5, 15, 12) {real, imag} */,
  {32'h406e78e4, 32'h41037866} /* (5, 15, 11) {real, imag} */,
  {32'h41df66a5, 32'hc19a8138} /* (5, 15, 10) {real, imag} */,
  {32'hc058ae27, 32'h4055ed03} /* (5, 15, 9) {real, imag} */,
  {32'hc212a1c2, 32'h3f0ab660} /* (5, 15, 8) {real, imag} */,
  {32'h40dfef6c, 32'hbdad6860} /* (5, 15, 7) {real, imag} */,
  {32'h3fff4e4c, 32'hc13fdc01} /* (5, 15, 6) {real, imag} */,
  {32'h40d2f6a0, 32'h414067fc} /* (5, 15, 5) {real, imag} */,
  {32'h4169e481, 32'h4097fd57} /* (5, 15, 4) {real, imag} */,
  {32'hc15ea388, 32'h3f811a10} /* (5, 15, 3) {real, imag} */,
  {32'hc1b2b146, 32'hc149bf5c} /* (5, 15, 2) {real, imag} */,
  {32'h41f730f2, 32'h414d3bcd} /* (5, 15, 1) {real, imag} */,
  {32'h4274ec83, 32'h42a1a6d9} /* (5, 15, 0) {real, imag} */,
  {32'hc1c945a5, 32'h40f29997} /* (5, 14, 31) {real, imag} */,
  {32'hc0eab31c, 32'h4120b72d} /* (5, 14, 30) {real, imag} */,
  {32'hc1f7a89b, 32'h41bc544c} /* (5, 14, 29) {real, imag} */,
  {32'hc198886d, 32'h40fd2e6e} /* (5, 14, 28) {real, imag} */,
  {32'hc26088a4, 32'hc10d6594} /* (5, 14, 27) {real, imag} */,
  {32'hc222cb11, 32'h4177a8c2} /* (5, 14, 26) {real, imag} */,
  {32'hc2281234, 32'hc221ae54} /* (5, 14, 25) {real, imag} */,
  {32'hc18dc809, 32'hc1adfaa6} /* (5, 14, 24) {real, imag} */,
  {32'h410989ee, 32'h41b07a2b} /* (5, 14, 23) {real, imag} */,
  {32'hc194f7c3, 32'h41129f3a} /* (5, 14, 22) {real, imag} */,
  {32'h419f7efb, 32'hc0c67806} /* (5, 14, 21) {real, imag} */,
  {32'h3eb651c0, 32'hc180d5e0} /* (5, 14, 20) {real, imag} */,
  {32'h3fe9c1c0, 32'hbff80b96} /* (5, 14, 19) {real, imag} */,
  {32'h4026e228, 32'hc127c0ce} /* (5, 14, 18) {real, imag} */,
  {32'h411c014a, 32'hc1837ca7} /* (5, 14, 17) {real, imag} */,
  {32'h409862bc, 32'h4125a508} /* (5, 14, 16) {real, imag} */,
  {32'hc0e9ba44, 32'hc07a02e2} /* (5, 14, 15) {real, imag} */,
  {32'h402f6868, 32'hc12972ec} /* (5, 14, 14) {real, imag} */,
  {32'h410275f8, 32'h411d6759} /* (5, 14, 13) {real, imag} */,
  {32'h41802c31, 32'hc134460e} /* (5, 14, 12) {real, imag} */,
  {32'hc1b973c1, 32'hc1b17ade} /* (5, 14, 11) {real, imag} */,
  {32'h41427e86, 32'h417ee842} /* (5, 14, 10) {real, imag} */,
  {32'hc085b06b, 32'h42075c86} /* (5, 14, 9) {real, imag} */,
  {32'h41bf3aed, 32'h41580c70} /* (5, 14, 8) {real, imag} */,
  {32'hc0af8c74, 32'h419b983e} /* (5, 14, 7) {real, imag} */,
  {32'h40aaa800, 32'h41ab5de5} /* (5, 14, 6) {real, imag} */,
  {32'h401a1428, 32'h422d1bc9} /* (5, 14, 5) {real, imag} */,
  {32'hc23595d8, 32'hc1b69a20} /* (5, 14, 4) {real, imag} */,
  {32'h417e169a, 32'hc0db7af8} /* (5, 14, 3) {real, imag} */,
  {32'h428ad44d, 32'h41c45782} /* (5, 14, 2) {real, imag} */,
  {32'hc271c8d4, 32'h41433f56} /* (5, 14, 1) {real, imag} */,
  {32'h41a88a61, 32'h4202ee7b} /* (5, 14, 0) {real, imag} */,
  {32'h40bf36d0, 32'hc2169cb4} /* (5, 13, 31) {real, imag} */,
  {32'hc07c7b2f, 32'h41fb40c6} /* (5, 13, 30) {real, imag} */,
  {32'h425b6cb7, 32'h41a11434} /* (5, 13, 29) {real, imag} */,
  {32'h4067799e, 32'hc1c5243a} /* (5, 13, 28) {real, imag} */,
  {32'hc23d7d10, 32'hc1e3ebda} /* (5, 13, 27) {real, imag} */,
  {32'h420fc01c, 32'h4106bf7c} /* (5, 13, 26) {real, imag} */,
  {32'h41d09fc8, 32'hc20a63b6} /* (5, 13, 25) {real, imag} */,
  {32'h41026563, 32'hc091f78c} /* (5, 13, 24) {real, imag} */,
  {32'hc1983655, 32'hc2236ce6} /* (5, 13, 23) {real, imag} */,
  {32'h419f075a, 32'h423bd273} /* (5, 13, 22) {real, imag} */,
  {32'hc1b08b15, 32'h41a3a3d0} /* (5, 13, 21) {real, imag} */,
  {32'h41637722, 32'hc080f538} /* (5, 13, 20) {real, imag} */,
  {32'hbeca2050, 32'hc0136e52} /* (5, 13, 19) {real, imag} */,
  {32'hc114ceb2, 32'h412ee45b} /* (5, 13, 18) {real, imag} */,
  {32'h40f6b2ae, 32'h400053be} /* (5, 13, 17) {real, imag} */,
  {32'h3f0dd680, 32'hc0442d40} /* (5, 13, 16) {real, imag} */,
  {32'h4060f484, 32'h40ef78fb} /* (5, 13, 15) {real, imag} */,
  {32'hc056fa21, 32'hc200a5bf} /* (5, 13, 14) {real, imag} */,
  {32'hc14b5cca, 32'hc1001794} /* (5, 13, 13) {real, imag} */,
  {32'hc05bb776, 32'h414c9842} /* (5, 13, 12) {real, imag} */,
  {32'h411e3590, 32'h40d09338} /* (5, 13, 11) {real, imag} */,
  {32'h3f1c3070, 32'hc13fbf48} /* (5, 13, 10) {real, imag} */,
  {32'h416720b2, 32'h40c201ec} /* (5, 13, 9) {real, imag} */,
  {32'h419b7c00, 32'hc217fb96} /* (5, 13, 8) {real, imag} */,
  {32'h41a78db4, 32'h404f9028} /* (5, 13, 7) {real, imag} */,
  {32'hc1cbe076, 32'h41e97f34} /* (5, 13, 6) {real, imag} */,
  {32'h41f5d285, 32'hc0347fc0} /* (5, 13, 5) {real, imag} */,
  {32'h40fcc967, 32'h41210f74} /* (5, 13, 4) {real, imag} */,
  {32'h423ddde5, 32'h419497e8} /* (5, 13, 3) {real, imag} */,
  {32'h40a4fc2c, 32'hc1d8c436} /* (5, 13, 2) {real, imag} */,
  {32'hc1eeb720, 32'h41d75d61} /* (5, 13, 1) {real, imag} */,
  {32'hc23d9c75, 32'h424cccd4} /* (5, 13, 0) {real, imag} */,
  {32'hc2063a4c, 32'hc1880942} /* (5, 12, 31) {real, imag} */,
  {32'hc2300b8c, 32'hc23d68f9} /* (5, 12, 30) {real, imag} */,
  {32'hc1967712, 32'hc21fa8eb} /* (5, 12, 29) {real, imag} */,
  {32'hc1b83ded, 32'hc1e98477} /* (5, 12, 28) {real, imag} */,
  {32'h42291522, 32'h41d25b3d} /* (5, 12, 27) {real, imag} */,
  {32'hc1b83d23, 32'h4208059c} /* (5, 12, 26) {real, imag} */,
  {32'h40c7da78, 32'h41cf477a} /* (5, 12, 25) {real, imag} */,
  {32'h4229003a, 32'h41c292c6} /* (5, 12, 24) {real, imag} */,
  {32'h41aca40e, 32'hc1d608f3} /* (5, 12, 23) {real, imag} */,
  {32'hc1a18a12, 32'hc0b74378} /* (5, 12, 22) {real, imag} */,
  {32'h403c6b18, 32'hc1c91b8f} /* (5, 12, 21) {real, imag} */,
  {32'h41150217, 32'h3efe9150} /* (5, 12, 20) {real, imag} */,
  {32'h40bf8916, 32'h40d161d6} /* (5, 12, 19) {real, imag} */,
  {32'hbfda39ac, 32'hc1017236} /* (5, 12, 18) {real, imag} */,
  {32'h40add3e1, 32'h41a05884} /* (5, 12, 17) {real, imag} */,
  {32'h403fdf88, 32'hc04865f4} /* (5, 12, 16) {real, imag} */,
  {32'h4075bd42, 32'h3f5e9170} /* (5, 12, 15) {real, imag} */,
  {32'h41471e86, 32'h418dd6e4} /* (5, 12, 14) {real, imag} */,
  {32'h3deafea0, 32'hc1604dcd} /* (5, 12, 13) {real, imag} */,
  {32'hc14ba351, 32'hbfea0ea4} /* (5, 12, 12) {real, imag} */,
  {32'hc204aeda, 32'h418968a3} /* (5, 12, 11) {real, imag} */,
  {32'h408af8c2, 32'hc0c408d0} /* (5, 12, 10) {real, imag} */,
  {32'h417e8c23, 32'h4136d282} /* (5, 12, 9) {real, imag} */,
  {32'h40ef5c94, 32'h4194d30e} /* (5, 12, 8) {real, imag} */,
  {32'h42414dd3, 32'h4208447c} /* (5, 12, 7) {real, imag} */,
  {32'hc21835e2, 32'hc09e26cc} /* (5, 12, 6) {real, imag} */,
  {32'hbfaa8e50, 32'hc2589cea} /* (5, 12, 5) {real, imag} */,
  {32'hc184258b, 32'hc18784bd} /* (5, 12, 4) {real, imag} */,
  {32'hc084d89c, 32'h4147d7fb} /* (5, 12, 3) {real, imag} */,
  {32'hc1a6ba6f, 32'h420b4443} /* (5, 12, 2) {real, imag} */,
  {32'h4209c586, 32'hc114b129} /* (5, 12, 1) {real, imag} */,
  {32'h426a3a66, 32'hc1dd8460} /* (5, 12, 0) {real, imag} */,
  {32'h42690c89, 32'h4116d3ec} /* (5, 11, 31) {real, imag} */,
  {32'h4217ff9e, 32'h42774973} /* (5, 11, 30) {real, imag} */,
  {32'hc113fadf, 32'hc204445a} /* (5, 11, 29) {real, imag} */,
  {32'hc21cde74, 32'h421d66db} /* (5, 11, 28) {real, imag} */,
  {32'h428546ef, 32'h3fcef328} /* (5, 11, 27) {real, imag} */,
  {32'hc17a4600, 32'hc20c0887} /* (5, 11, 26) {real, imag} */,
  {32'hc1fbbca9, 32'hc111271f} /* (5, 11, 25) {real, imag} */,
  {32'hc218dbb6, 32'hc05d8d78} /* (5, 11, 24) {real, imag} */,
  {32'h416e9592, 32'hc05c4970} /* (5, 11, 23) {real, imag} */,
  {32'h4148b4a0, 32'hc04bc518} /* (5, 11, 22) {real, imag} */,
  {32'h409cdaa0, 32'hc1bf4efc} /* (5, 11, 21) {real, imag} */,
  {32'h417fe532, 32'h4121f23a} /* (5, 11, 20) {real, imag} */,
  {32'h4182c355, 32'hbe29e060} /* (5, 11, 19) {real, imag} */,
  {32'hc1229ce1, 32'hc1a90c4a} /* (5, 11, 18) {real, imag} */,
  {32'h40ea0225, 32'h40d4f100} /* (5, 11, 17) {real, imag} */,
  {32'h41004d4e, 32'hc0453ae0} /* (5, 11, 16) {real, imag} */,
  {32'hc0fce7a3, 32'hc1c4b4de} /* (5, 11, 15) {real, imag} */,
  {32'h41168dcf, 32'h3f946800} /* (5, 11, 14) {real, imag} */,
  {32'h416d5484, 32'h40e8475b} /* (5, 11, 13) {real, imag} */,
  {32'h40f16e33, 32'hc01bf2d8} /* (5, 11, 12) {real, imag} */,
  {32'h41070a84, 32'h424fa8be} /* (5, 11, 11) {real, imag} */,
  {32'hc2264d5c, 32'hc132bfda} /* (5, 11, 10) {real, imag} */,
  {32'hbe57eb80, 32'hc292f808} /* (5, 11, 9) {real, imag} */,
  {32'h4031b338, 32'h415767fe} /* (5, 11, 8) {real, imag} */,
  {32'hc1b91051, 32'hc133d34f} /* (5, 11, 7) {real, imag} */,
  {32'h425b225a, 32'hc2382d75} /* (5, 11, 6) {real, imag} */,
  {32'h41d7193d, 32'h402fb1d4} /* (5, 11, 5) {real, imag} */,
  {32'hc0dcadbc, 32'h42294075} /* (5, 11, 4) {real, imag} */,
  {32'h3f1cfb50, 32'hbf7e8620} /* (5, 11, 3) {real, imag} */,
  {32'hc1de4097, 32'hc1c601fa} /* (5, 11, 2) {real, imag} */,
  {32'hc236c863, 32'hc22bf990} /* (5, 11, 1) {real, imag} */,
  {32'hc27a006c, 32'h42720b92} /* (5, 11, 0) {real, imag} */,
  {32'hc2aa4e50, 32'h4151e152} /* (5, 10, 31) {real, imag} */,
  {32'hc08401e8, 32'hc203eaa5} /* (5, 10, 30) {real, imag} */,
  {32'h41b1985f, 32'hc29aae78} /* (5, 10, 29) {real, imag} */,
  {32'h42791048, 32'h4259c0e2} /* (5, 10, 28) {real, imag} */,
  {32'hc120c952, 32'h415baa6c} /* (5, 10, 27) {real, imag} */,
  {32'hc06ebe80, 32'hc08c8750} /* (5, 10, 26) {real, imag} */,
  {32'h42121abe, 32'h40bc8cb0} /* (5, 10, 25) {real, imag} */,
  {32'hc0a07ec0, 32'hc215063c} /* (5, 10, 24) {real, imag} */,
  {32'hc10b234a, 32'h421e6b35} /* (5, 10, 23) {real, imag} */,
  {32'hc140f90c, 32'hc1247b48} /* (5, 10, 22) {real, imag} */,
  {32'h410cb52d, 32'h40561348} /* (5, 10, 21) {real, imag} */,
  {32'hc1cb4ab8, 32'hc00b14c0} /* (5, 10, 20) {real, imag} */,
  {32'h41885949, 32'h41c339e6} /* (5, 10, 19) {real, imag} */,
  {32'h41183eb9, 32'h409a298a} /* (5, 10, 18) {real, imag} */,
  {32'hc09438c3, 32'hbfc56630} /* (5, 10, 17) {real, imag} */,
  {32'h412a87f8, 32'hc206a288} /* (5, 10, 16) {real, imag} */,
  {32'hc024d786, 32'h41f7e79d} /* (5, 10, 15) {real, imag} */,
  {32'h405165cc, 32'hbe842ba0} /* (5, 10, 14) {real, imag} */,
  {32'hc1f45967, 32'h3fb98388} /* (5, 10, 13) {real, imag} */,
  {32'hc0e93548, 32'h4114f7fc} /* (5, 10, 12) {real, imag} */,
  {32'h41e6eed2, 32'hc188c17b} /* (5, 10, 11) {real, imag} */,
  {32'hc1c6ffd4, 32'hc22d9dee} /* (5, 10, 10) {real, imag} */,
  {32'hc23e3b68, 32'hc2261e6f} /* (5, 10, 9) {real, imag} */,
  {32'h4284a290, 32'h4195edee} /* (5, 10, 8) {real, imag} */,
  {32'hc17736c2, 32'h40a8f950} /* (5, 10, 7) {real, imag} */,
  {32'hc2265e07, 32'hc254b02e} /* (5, 10, 6) {real, imag} */,
  {32'h4115755c, 32'h427e9391} /* (5, 10, 5) {real, imag} */,
  {32'h41cb8478, 32'hc12d2eca} /* (5, 10, 4) {real, imag} */,
  {32'hc20247d3, 32'hc10eeb34} /* (5, 10, 3) {real, imag} */,
  {32'h422b4941, 32'h40690f30} /* (5, 10, 2) {real, imag} */,
  {32'h42abd910, 32'hc225679c} /* (5, 10, 1) {real, imag} */,
  {32'h43030176, 32'h42b92a64} /* (5, 10, 0) {real, imag} */,
  {32'h431189c3, 32'h4284f3e5} /* (5, 9, 31) {real, imag} */,
  {32'hc2b91e6a, 32'h41bdb18a} /* (5, 9, 30) {real, imag} */,
  {32'hc1393d3a, 32'h42054e12} /* (5, 9, 29) {real, imag} */,
  {32'hc11cde78, 32'hc2489b50} /* (5, 9, 28) {real, imag} */,
  {32'hc28b3866, 32'h425eb5f6} /* (5, 9, 27) {real, imag} */,
  {32'hc2b036df, 32'hc246ef6a} /* (5, 9, 26) {real, imag} */,
  {32'hc13db7e6, 32'hc13f4e4c} /* (5, 9, 25) {real, imag} */,
  {32'hc143f394, 32'h40ba8ca9} /* (5, 9, 24) {real, imag} */,
  {32'hc1b8742f, 32'h40af4728} /* (5, 9, 23) {real, imag} */,
  {32'h425f2208, 32'h420fa734} /* (5, 9, 22) {real, imag} */,
  {32'h42403b46, 32'h4203b502} /* (5, 9, 21) {real, imag} */,
  {32'hc1ff57b7, 32'h418ddc3a} /* (5, 9, 20) {real, imag} */,
  {32'h40db56d0, 32'h41b07989} /* (5, 9, 19) {real, imag} */,
  {32'hc0fb6978, 32'hc1cd6f72} /* (5, 9, 18) {real, imag} */,
  {32'hc1d52b76, 32'h416b72fc} /* (5, 9, 17) {real, imag} */,
  {32'h41b47e78, 32'h4166ccb0} /* (5, 9, 16) {real, imag} */,
  {32'hc1e610fe, 32'hc205860d} /* (5, 9, 15) {real, imag} */,
  {32'h41a17a12, 32'hc12b0134} /* (5, 9, 14) {real, imag} */,
  {32'hc1345e18, 32'hc15dab1e} /* (5, 9, 13) {real, imag} */,
  {32'h4189bda1, 32'h40971b28} /* (5, 9, 12) {real, imag} */,
  {32'h415c4f08, 32'hc11bb682} /* (5, 9, 11) {real, imag} */,
  {32'hc1c159b4, 32'hc0fb4dfc} /* (5, 9, 10) {real, imag} */,
  {32'h3fb9bdd0, 32'hc095846c} /* (5, 9, 9) {real, imag} */,
  {32'hc1695ad4, 32'hc11c2498} /* (5, 9, 8) {real, imag} */,
  {32'h428a8987, 32'h42302983} /* (5, 9, 7) {real, imag} */,
  {32'hc1a28200, 32'h4290e347} /* (5, 9, 6) {real, imag} */,
  {32'h4216bf28, 32'h409a33bc} /* (5, 9, 5) {real, imag} */,
  {32'h429aca3f, 32'hc1910ac0} /* (5, 9, 4) {real, imag} */,
  {32'h4223ac22, 32'hc2a3671f} /* (5, 9, 3) {real, imag} */,
  {32'h41ddc05a, 32'hc2a675be} /* (5, 9, 2) {real, imag} */,
  {32'hc22872c1, 32'h429fd4c3} /* (5, 9, 1) {real, imag} */,
  {32'hc298775e, 32'h41496648} /* (5, 9, 0) {real, imag} */,
  {32'hc24ddfec, 32'h430b1077} /* (5, 8, 31) {real, imag} */,
  {32'h4231ea65, 32'h411a6006} /* (5, 8, 30) {real, imag} */,
  {32'h41eb28d2, 32'hc23e4fde} /* (5, 8, 29) {real, imag} */,
  {32'hc22ab7ea, 32'h420dd6cf} /* (5, 8, 28) {real, imag} */,
  {32'h421a2c9e, 32'h41beb3bc} /* (5, 8, 27) {real, imag} */,
  {32'hc1e5b411, 32'hc2869efa} /* (5, 8, 26) {real, imag} */,
  {32'h42ce2114, 32'hc16badea} /* (5, 8, 25) {real, imag} */,
  {32'h42c23854, 32'hc2971b08} /* (5, 8, 24) {real, imag} */,
  {32'hc097c1c4, 32'hc222dfc8} /* (5, 8, 23) {real, imag} */,
  {32'hc277e2f0, 32'h4239d6f2} /* (5, 8, 22) {real, imag} */,
  {32'h41800e44, 32'hc254570a} /* (5, 8, 21) {real, imag} */,
  {32'h41c4a2eb, 32'h41cebc43} /* (5, 8, 20) {real, imag} */,
  {32'hc1477d3c, 32'h41a5cef0} /* (5, 8, 19) {real, imag} */,
  {32'hc1915f2c, 32'h41732926} /* (5, 8, 18) {real, imag} */,
  {32'hc129333e, 32'h41b9f8c4} /* (5, 8, 17) {real, imag} */,
  {32'h417237c8, 32'h41b3e313} /* (5, 8, 16) {real, imag} */,
  {32'h3fa6b0b0, 32'hbfc1be40} /* (5, 8, 15) {real, imag} */,
  {32'h4204d2f0, 32'hc01475f6} /* (5, 8, 14) {real, imag} */,
  {32'hc0a42aa8, 32'hc160487c} /* (5, 8, 13) {real, imag} */,
  {32'hc1ad59bb, 32'h407b1ad8} /* (5, 8, 12) {real, imag} */,
  {32'h418ce2ca, 32'hc224f210} /* (5, 8, 11) {real, imag} */,
  {32'hc1e2ad8d, 32'h41bc9e20} /* (5, 8, 10) {real, imag} */,
  {32'h4213ef06, 32'h4190864f} /* (5, 8, 9) {real, imag} */,
  {32'h40472380, 32'h41d72de8} /* (5, 8, 8) {real, imag} */,
  {32'h41f60890, 32'hc1c02e8d} /* (5, 8, 7) {real, imag} */,
  {32'hc283c939, 32'h4220553a} /* (5, 8, 6) {real, imag} */,
  {32'hc2099d42, 32'h410aa619} /* (5, 8, 5) {real, imag} */,
  {32'hc2b94d3b, 32'h4208eab5} /* (5, 8, 4) {real, imag} */,
  {32'h3fb5c7a0, 32'hc22525e2} /* (5, 8, 3) {real, imag} */,
  {32'hc282b0fa, 32'hc1da510b} /* (5, 8, 2) {real, imag} */,
  {32'hc287a8b9, 32'h4120d410} /* (5, 8, 1) {real, imag} */,
  {32'hc2b53461, 32'h411b7f82} /* (5, 8, 0) {real, imag} */,
  {32'hbfaef3c0, 32'hc2bf3525} /* (5, 7, 31) {real, imag} */,
  {32'hc1f78042, 32'hc1e6f84a} /* (5, 7, 30) {real, imag} */,
  {32'hc23d7d8b, 32'hc2b1539d} /* (5, 7, 29) {real, imag} */,
  {32'hc1a7726c, 32'h41e80466} /* (5, 7, 28) {real, imag} */,
  {32'h42d4ee56, 32'h406e9ca0} /* (5, 7, 27) {real, imag} */,
  {32'h421ae930, 32'h403ace00} /* (5, 7, 26) {real, imag} */,
  {32'h4311e7db, 32'h428fd714} /* (5, 7, 25) {real, imag} */,
  {32'h42d77162, 32'hc2ca7321} /* (5, 7, 24) {real, imag} */,
  {32'hc1a0f03b, 32'h42b3e79e} /* (5, 7, 23) {real, imag} */,
  {32'hc1c311d7, 32'h421ad2f5} /* (5, 7, 22) {real, imag} */,
  {32'hc2146361, 32'hc2390346} /* (5, 7, 21) {real, imag} */,
  {32'h4135ff6c, 32'h42214337} /* (5, 7, 20) {real, imag} */,
  {32'hc21d4748, 32'hc1a7591a} /* (5, 7, 19) {real, imag} */,
  {32'hc1d5d361, 32'h419fa4dc} /* (5, 7, 18) {real, imag} */,
  {32'h418dea1c, 32'h41dace3e} /* (5, 7, 17) {real, imag} */,
  {32'hc1e429d9, 32'hc115d6f8} /* (5, 7, 16) {real, imag} */,
  {32'h3f555380, 32'hc17e3bac} /* (5, 7, 15) {real, imag} */,
  {32'hbfe0c410, 32'hc1504639} /* (5, 7, 14) {real, imag} */,
  {32'h421eb368, 32'h416f5f74} /* (5, 7, 13) {real, imag} */,
  {32'h410e2e54, 32'hbfbea360} /* (5, 7, 12) {real, imag} */,
  {32'h411ea9b5, 32'h4291d3d6} /* (5, 7, 11) {real, imag} */,
  {32'h418f13e7, 32'hc151fb00} /* (5, 7, 10) {real, imag} */,
  {32'h4288fcd9, 32'hc1d805b4} /* (5, 7, 9) {real, imag} */,
  {32'hc28db922, 32'h4257d5a6} /* (5, 7, 8) {real, imag} */,
  {32'hc2d64901, 32'hc10e4604} /* (5, 7, 7) {real, imag} */,
  {32'h428df186, 32'h430bc5f5} /* (5, 7, 6) {real, imag} */,
  {32'hc22714bb, 32'hc26b8fec} /* (5, 7, 5) {real, imag} */,
  {32'hc1540939, 32'h42fdac48} /* (5, 7, 4) {real, imag} */,
  {32'h42943a46, 32'hc1d94b34} /* (5, 7, 3) {real, imag} */,
  {32'hc2ae4a4a, 32'h422f6797} /* (5, 7, 2) {real, imag} */,
  {32'h43435270, 32'hc2bdec69} /* (5, 7, 1) {real, imag} */,
  {32'hc288a5c1, 32'h41369a30} /* (5, 7, 0) {real, imag} */,
  {32'h418046b4, 32'h4314ce31} /* (5, 6, 31) {real, imag} */,
  {32'h421643f4, 32'hc2ad6d76} /* (5, 6, 30) {real, imag} */,
  {32'h40cb1f12, 32'hc1b23813} /* (5, 6, 29) {real, imag} */,
  {32'hc22c496f, 32'h42c412c7} /* (5, 6, 28) {real, imag} */,
  {32'h41a64e84, 32'hc14b69a3} /* (5, 6, 27) {real, imag} */,
  {32'hc1d12776, 32'hc163497c} /* (5, 6, 26) {real, imag} */,
  {32'hc2833c9e, 32'hbfc55ad8} /* (5, 6, 25) {real, imag} */,
  {32'h41d7caa2, 32'hc1a34e02} /* (5, 6, 24) {real, imag} */,
  {32'h421f5790, 32'hc17ac8e7} /* (5, 6, 23) {real, imag} */,
  {32'h4145cd8c, 32'hc1c08da8} /* (5, 6, 22) {real, imag} */,
  {32'h41f5aa1e, 32'hc1470f50} /* (5, 6, 21) {real, imag} */,
  {32'h41c45d23, 32'h41ef8d4f} /* (5, 6, 20) {real, imag} */,
  {32'hc18d8aa8, 32'hc0e5b824} /* (5, 6, 19) {real, imag} */,
  {32'hc24a6c0b, 32'hc00323f0} /* (5, 6, 18) {real, imag} */,
  {32'hc17a2536, 32'hc243cbab} /* (5, 6, 17) {real, imag} */,
  {32'h40bd364c, 32'h425d4a78} /* (5, 6, 16) {real, imag} */,
  {32'hc1a0b6af, 32'hc04c3d50} /* (5, 6, 15) {real, imag} */,
  {32'h411ff960, 32'hc0ce9cc8} /* (5, 6, 14) {real, imag} */,
  {32'hc19c07f4, 32'hc2133156} /* (5, 6, 13) {real, imag} */,
  {32'h4133cbda, 32'h41820551} /* (5, 6, 12) {real, imag} */,
  {32'hbfc87dc8, 32'hc28c3801} /* (5, 6, 11) {real, imag} */,
  {32'h42c4ba34, 32'hc21911ce} /* (5, 6, 10) {real, imag} */,
  {32'h41af0daa, 32'h40c8827a} /* (5, 6, 9) {real, imag} */,
  {32'h4296f84e, 32'h4276296f} /* (5, 6, 8) {real, imag} */,
  {32'hc23ab2dd, 32'hc0c5ffbe} /* (5, 6, 7) {real, imag} */,
  {32'h42b17f84, 32'hc29e6544} /* (5, 6, 6) {real, imag} */,
  {32'hc2a0f7b3, 32'h40b1cbf6} /* (5, 6, 5) {real, imag} */,
  {32'hc2299de3, 32'h4207c03a} /* (5, 6, 4) {real, imag} */,
  {32'hc11bfbed, 32'hc2a3ec3a} /* (5, 6, 3) {real, imag} */,
  {32'h429c4240, 32'h42279cd5} /* (5, 6, 2) {real, imag} */,
  {32'hc3189ef0, 32'hc132b830} /* (5, 6, 1) {real, imag} */,
  {32'h4184ae53, 32'hc21f18ce} /* (5, 6, 0) {real, imag} */,
  {32'hc281fdef, 32'h4263789c} /* (5, 5, 31) {real, imag} */,
  {32'h42857742, 32'hc0d88382} /* (5, 5, 30) {real, imag} */,
  {32'h42aa6349, 32'h4283ca92} /* (5, 5, 29) {real, imag} */,
  {32'hc2ac6e46, 32'h415a97c0} /* (5, 5, 28) {real, imag} */,
  {32'hc1674a76, 32'hc218a405} /* (5, 5, 27) {real, imag} */,
  {32'h4141e5f4, 32'h428ec96f} /* (5, 5, 26) {real, imag} */,
  {32'h4291f24d, 32'hc0f5cfb4} /* (5, 5, 25) {real, imag} */,
  {32'h42cbdf46, 32'hc2b1f924} /* (5, 5, 24) {real, imag} */,
  {32'h421d66e3, 32'h4277c35e} /* (5, 5, 23) {real, imag} */,
  {32'h424d72c9, 32'h420d2f55} /* (5, 5, 22) {real, imag} */,
  {32'hc10a30ee, 32'hc2274159} /* (5, 5, 21) {real, imag} */,
  {32'h40f00500, 32'hc1508fd6} /* (5, 5, 20) {real, imag} */,
  {32'h3e970bc0, 32'h41bc4e22} /* (5, 5, 19) {real, imag} */,
  {32'hc1bc1b75, 32'hbf034cc0} /* (5, 5, 18) {real, imag} */,
  {32'hc0e9adfc, 32'h411868a4} /* (5, 5, 17) {real, imag} */,
  {32'hc11f2270, 32'hc0efe100} /* (5, 5, 16) {real, imag} */,
  {32'h416a9ca6, 32'hc12ddc14} /* (5, 5, 15) {real, imag} */,
  {32'hc1d9fd5d, 32'h42342ced} /* (5, 5, 14) {real, imag} */,
  {32'hc1cbd79b, 32'h420f9955} /* (5, 5, 13) {real, imag} */,
  {32'hc1f4ff38, 32'hc0ef6fac} /* (5, 5, 12) {real, imag} */,
  {32'h422f3980, 32'h4151b87c} /* (5, 5, 11) {real, imag} */,
  {32'hc095d9d8, 32'h40bdbe4a} /* (5, 5, 10) {real, imag} */,
  {32'hc203d425, 32'hc0fb0ecc} /* (5, 5, 9) {real, imag} */,
  {32'hc13b32a4, 32'h403ce310} /* (5, 5, 8) {real, imag} */,
  {32'h42c2341f, 32'h4258c4be} /* (5, 5, 7) {real, imag} */,
  {32'h42c5e500, 32'hc0b7f790} /* (5, 5, 6) {real, imag} */,
  {32'h4248208e, 32'hc2849050} /* (5, 5, 5) {real, imag} */,
  {32'hbfbba5a0, 32'hc2fdd4cc} /* (5, 5, 4) {real, imag} */,
  {32'hc1a9f50c, 32'h41df377a} /* (5, 5, 3) {real, imag} */,
  {32'hc2e593d0, 32'h413fccb1} /* (5, 5, 2) {real, imag} */,
  {32'hc33e63ee, 32'h43169d31} /* (5, 5, 1) {real, imag} */,
  {32'hc361851f, 32'h42c1ffb6} /* (5, 5, 0) {real, imag} */,
  {32'h427b100a, 32'hc1214214} /* (5, 4, 31) {real, imag} */,
  {32'hc37ee45d, 32'hc33e6ad0} /* (5, 4, 30) {real, imag} */,
  {32'hc1b0ad47, 32'hc1a3fd99} /* (5, 4, 29) {real, imag} */,
  {32'h4302c0a7, 32'hc2f167f4} /* (5, 4, 28) {real, imag} */,
  {32'h42da8550, 32'hc23950e1} /* (5, 4, 27) {real, imag} */,
  {32'h418aa15c, 32'hc33592c5} /* (5, 4, 26) {real, imag} */,
  {32'h4288b46d, 32'h430cc50e} /* (5, 4, 25) {real, imag} */,
  {32'hc2497ae5, 32'h425b17e4} /* (5, 4, 24) {real, imag} */,
  {32'hc21a3bbe, 32'h41efd857} /* (5, 4, 23) {real, imag} */,
  {32'h40c74940, 32'hc1eff6f9} /* (5, 4, 22) {real, imag} */,
  {32'hc15def12, 32'h4237db26} /* (5, 4, 21) {real, imag} */,
  {32'hc10a5d80, 32'h41ae9722} /* (5, 4, 20) {real, imag} */,
  {32'h40083ec8, 32'h421d539c} /* (5, 4, 19) {real, imag} */,
  {32'hc0e505e0, 32'h40f8ab80} /* (5, 4, 18) {real, imag} */,
  {32'hc0fec0d8, 32'h4208da43} /* (5, 4, 17) {real, imag} */,
  {32'h406077c0, 32'hc183918a} /* (5, 4, 16) {real, imag} */,
  {32'hc0fad9f8, 32'hc18f55ea} /* (5, 4, 15) {real, imag} */,
  {32'hc2502c74, 32'h41c21798} /* (5, 4, 14) {real, imag} */,
  {32'h4261365c, 32'hc15cbfc8} /* (5, 4, 13) {real, imag} */,
  {32'h4131b618, 32'h41f64dae} /* (5, 4, 12) {real, imag} */,
  {32'h420c114c, 32'h4207003e} /* (5, 4, 11) {real, imag} */,
  {32'hc166d420, 32'hc1bee1f9} /* (5, 4, 10) {real, imag} */,
  {32'hc23f09b6, 32'hc286df63} /* (5, 4, 9) {real, imag} */,
  {32'hc2191f35, 32'h406276c0} /* (5, 4, 8) {real, imag} */,
  {32'h41ba3dfb, 32'hc1d6a434} /* (5, 4, 7) {real, imag} */,
  {32'hc30726f0, 32'h411995b0} /* (5, 4, 6) {real, imag} */,
  {32'hc1cb7f50, 32'h41b1c9fe} /* (5, 4, 5) {real, imag} */,
  {32'hc258118d, 32'h422398f0} /* (5, 4, 4) {real, imag} */,
  {32'h3ecc61c0, 32'h422af086} /* (5, 4, 3) {real, imag} */,
  {32'hc354d6e3, 32'h4256a8b4} /* (5, 4, 2) {real, imag} */,
  {32'h43157c1a, 32'hc24ff6f9} /* (5, 4, 1) {real, imag} */,
  {32'h4379e00b, 32'hc2801dfe} /* (5, 4, 0) {real, imag} */,
  {32'hc33eb8cf, 32'h41ac4df6} /* (5, 3, 31) {real, imag} */,
  {32'hc29b11af, 32'hc2987b23} /* (5, 3, 30) {real, imag} */,
  {32'h41af2f88, 32'h42dafb24} /* (5, 3, 29) {real, imag} */,
  {32'h422b9366, 32'hc19112ca} /* (5, 3, 28) {real, imag} */,
  {32'hc1702660, 32'h42e97d99} /* (5, 3, 27) {real, imag} */,
  {32'hc2929f59, 32'hc2997b10} /* (5, 3, 26) {real, imag} */,
  {32'h3f1ced40, 32'h42cb1523} /* (5, 3, 25) {real, imag} */,
  {32'hc2301685, 32'h426cb333} /* (5, 3, 24) {real, imag} */,
  {32'h42785a66, 32'h427e6784} /* (5, 3, 23) {real, imag} */,
  {32'h4201ac9c, 32'hc2437d77} /* (5, 3, 22) {real, imag} */,
  {32'h41dbcf98, 32'hc0d97908} /* (5, 3, 21) {real, imag} */,
  {32'hc07b9674, 32'hc22ba3ad} /* (5, 3, 20) {real, imag} */,
  {32'h41e27920, 32'hc1f7ac51} /* (5, 3, 19) {real, imag} */,
  {32'hc247b03e, 32'h3d9b7bc0} /* (5, 3, 18) {real, imag} */,
  {32'hc028abc0, 32'h41f64437} /* (5, 3, 17) {real, imag} */,
  {32'hc1d1ab22, 32'h4219d1ff} /* (5, 3, 16) {real, imag} */,
  {32'hc2059fac, 32'h4171782a} /* (5, 3, 15) {real, imag} */,
  {32'h425f345a, 32'h40658ebe} /* (5, 3, 14) {real, imag} */,
  {32'h41b566f8, 32'h4128627e} /* (5, 3, 13) {real, imag} */,
  {32'h420f51fa, 32'hc2a748da} /* (5, 3, 12) {real, imag} */,
  {32'h41aaaa2c, 32'hc1bedcf6} /* (5, 3, 11) {real, imag} */,
  {32'h424f3390, 32'hc16cb5dc} /* (5, 3, 10) {real, imag} */,
  {32'h40e5be54, 32'hc1009c88} /* (5, 3, 9) {real, imag} */,
  {32'h4285b44c, 32'hc1bc930e} /* (5, 3, 8) {real, imag} */,
  {32'hc1726298, 32'h40322440} /* (5, 3, 7) {real, imag} */,
  {32'h409ad4d0, 32'h42cb195c} /* (5, 3, 6) {real, imag} */,
  {32'h43227f8a, 32'hc281f623} /* (5, 3, 5) {real, imag} */,
  {32'h404cb7f8, 32'h42fb19e0} /* (5, 3, 4) {real, imag} */,
  {32'h42fefb3e, 32'hc114f4e0} /* (5, 3, 3) {real, imag} */,
  {32'hc304c7a4, 32'h429be739} /* (5, 3, 2) {real, imag} */,
  {32'h43d1102e, 32'hc1b7530c} /* (5, 3, 1) {real, imag} */,
  {32'hc2f20340, 32'h42837f8a} /* (5, 3, 0) {real, imag} */,
  {32'hc357ae3c, 32'h44143def} /* (5, 2, 31) {real, imag} */,
  {32'h42bcf0f3, 32'hc401952d} /* (5, 2, 30) {real, imag} */,
  {32'hc27abbe1, 32'h42e5bf2a} /* (5, 2, 29) {real, imag} */,
  {32'h43371c57, 32'h43139417} /* (5, 2, 28) {real, imag} */,
  {32'h42c14481, 32'hc3548160} /* (5, 2, 27) {real, imag} */,
  {32'h4195e634, 32'hc2c454b4} /* (5, 2, 26) {real, imag} */,
  {32'hc26976c3, 32'h426063f1} /* (5, 2, 25) {real, imag} */,
  {32'h409ffdec, 32'h42e022f4} /* (5, 2, 24) {real, imag} */,
  {32'h41f2d7ee, 32'hc27ec599} /* (5, 2, 23) {real, imag} */,
  {32'hc228baca, 32'hc2391302} /* (5, 2, 22) {real, imag} */,
  {32'h41e4a494, 32'h40539c60} /* (5, 2, 21) {real, imag} */,
  {32'hc1da6339, 32'hc28d242c} /* (5, 2, 20) {real, imag} */,
  {32'h407d83cc, 32'h41e0be71} /* (5, 2, 19) {real, imag} */,
  {32'hc1eedeef, 32'hc0cbe550} /* (5, 2, 18) {real, imag} */,
  {32'h4288a1a9, 32'hc172b570} /* (5, 2, 17) {real, imag} */,
  {32'hc1faa73a, 32'h4223a7bc} /* (5, 2, 16) {real, imag} */,
  {32'h40413420, 32'h3ea6be00} /* (5, 2, 15) {real, imag} */,
  {32'h4155fdde, 32'hc114db38} /* (5, 2, 14) {real, imag} */,
  {32'hc05c442c, 32'hbf70af20} /* (5, 2, 13) {real, imag} */,
  {32'hc166d6f2, 32'h411e1588} /* (5, 2, 12) {real, imag} */,
  {32'h420d6422, 32'hc218da4c} /* (5, 2, 11) {real, imag} */,
  {32'h4108ea48, 32'hc22afe2c} /* (5, 2, 10) {real, imag} */,
  {32'hc2638def, 32'hc2102053} /* (5, 2, 9) {real, imag} */,
  {32'h42866316, 32'hc2945528} /* (5, 2, 8) {real, imag} */,
  {32'h40681a30, 32'h42df5dc2} /* (5, 2, 7) {real, imag} */,
  {32'hc27d70ea, 32'h42a056c4} /* (5, 2, 6) {real, imag} */,
  {32'h434c4078, 32'hc1bb9c20} /* (5, 2, 5) {real, imag} */,
  {32'hc345f579, 32'h422f003d} /* (5, 2, 4) {real, imag} */,
  {32'hc2215075, 32'h43355913} /* (5, 2, 3) {real, imag} */,
  {32'h4281d011, 32'hc3c8341a} /* (5, 2, 2) {real, imag} */,
  {32'hc2adf6df, 32'h435bd8db} /* (5, 2, 1) {real, imag} */,
  {32'hc21ddad9, 32'h41f015d5} /* (5, 2, 0) {real, imag} */,
  {32'h4320da77, 32'hc3c1e99f} /* (5, 1, 31) {real, imag} */,
  {32'hc27eaecc, 32'h4240c3fe} /* (5, 1, 30) {real, imag} */,
  {32'h4224ff22, 32'h42a3cef2} /* (5, 1, 29) {real, imag} */,
  {32'h430bc1e0, 32'h41a06704} /* (5, 1, 28) {real, imag} */,
  {32'hc31c8194, 32'h42f1c7d9} /* (5, 1, 27) {real, imag} */,
  {32'hc22861da, 32'hc1a8f57a} /* (5, 1, 26) {real, imag} */,
  {32'hc23a5f53, 32'hc155821c} /* (5, 1, 25) {real, imag} */,
  {32'hc23ad242, 32'h429dedbd} /* (5, 1, 24) {real, imag} */,
  {32'h41bd035e, 32'hc226eed5} /* (5, 1, 23) {real, imag} */,
  {32'h42595bd2, 32'h42133520} /* (5, 1, 22) {real, imag} */,
  {32'h420d1c6b, 32'h423de90c} /* (5, 1, 21) {real, imag} */,
  {32'hc20ea159, 32'hc15769b8} /* (5, 1, 20) {real, imag} */,
  {32'hc122cc32, 32'hc094a6ee} /* (5, 1, 19) {real, imag} */,
  {32'h42d6c6d5, 32'hc1d2adc4} /* (5, 1, 18) {real, imag} */,
  {32'hc23af630, 32'h41763e7c} /* (5, 1, 17) {real, imag} */,
  {32'hc1c75d9c, 32'hc018c680} /* (5, 1, 16) {real, imag} */,
  {32'hbffa4f00, 32'hc17778bc} /* (5, 1, 15) {real, imag} */,
  {32'hc173c038, 32'hc1bbb46c} /* (5, 1, 14) {real, imag} */,
  {32'hc0ff7524, 32'h3f0a7610} /* (5, 1, 13) {real, imag} */,
  {32'h4048e3f0, 32'h4272b7bc} /* (5, 1, 12) {real, imag} */,
  {32'hc29d621e, 32'hc1aa5e41} /* (5, 1, 11) {real, imag} */,
  {32'h4259ef1e, 32'h414e307c} /* (5, 1, 10) {real, imag} */,
  {32'hc2aea70e, 32'hc1c6fc7e} /* (5, 1, 9) {real, imag} */,
  {32'hc2806f9f, 32'hc236711a} /* (5, 1, 8) {real, imag} */,
  {32'h41acc7a2, 32'h42a2aba2} /* (5, 1, 7) {real, imag} */,
  {32'h4257f1a2, 32'hc1a6c558} /* (5, 1, 6) {real, imag} */,
  {32'hc2ae8ca8, 32'h3ec75300} /* (5, 1, 5) {real, imag} */,
  {32'h425a5e39, 32'hc2c803c2} /* (5, 1, 4) {real, imag} */,
  {32'hc1e8e8c1, 32'hc286a82e} /* (5, 1, 3) {real, imag} */,
  {32'hc3e6bf56, 32'h4356dabe} /* (5, 1, 2) {real, imag} */,
  {32'h440461d6, 32'hc34e64b6} /* (5, 1, 1) {real, imag} */,
  {32'h4353ff34, 32'hc3a57171} /* (5, 1, 0) {real, imag} */,
  {32'h40cbd800, 32'hc3ec2d52} /* (5, 0, 31) {real, imag} */,
  {32'h42a3fd42, 32'h43082617} /* (5, 0, 30) {real, imag} */,
  {32'hc2c82050, 32'hc212d538} /* (5, 0, 29) {real, imag} */,
  {32'h41b36217, 32'h4302e6d2} /* (5, 0, 28) {real, imag} */,
  {32'h412ecb27, 32'h434b0f12} /* (5, 0, 27) {real, imag} */,
  {32'hc25651e8, 32'hc1fc5ebe} /* (5, 0, 26) {real, imag} */,
  {32'hc2289cf2, 32'hc276fb3e} /* (5, 0, 25) {real, imag} */,
  {32'h41ca093e, 32'hc3193bac} /* (5, 0, 24) {real, imag} */,
  {32'hc2e3fe1f, 32'hc11c4a18} /* (5, 0, 23) {real, imag} */,
  {32'hc2a21d07, 32'hc1bbd486} /* (5, 0, 22) {real, imag} */,
  {32'hc09fb744, 32'h4281ea35} /* (5, 0, 21) {real, imag} */,
  {32'hc0befcdc, 32'hc2b51744} /* (5, 0, 20) {real, imag} */,
  {32'h40e02348, 32'h41f92c35} /* (5, 0, 19) {real, imag} */,
  {32'h426e4290, 32'h4105bb2c} /* (5, 0, 18) {real, imag} */,
  {32'hc01bd8e0, 32'h41e37448} /* (5, 0, 17) {real, imag} */,
  {32'h427b7f55, 32'hc1885630} /* (5, 0, 16) {real, imag} */,
  {32'hc0623a20, 32'h4111a210} /* (5, 0, 15) {real, imag} */,
  {32'hc18c9a99, 32'h420cd645} /* (5, 0, 14) {real, imag} */,
  {32'h42541543, 32'hc2444b02} /* (5, 0, 13) {real, imag} */,
  {32'h4202f33e, 32'hc282a394} /* (5, 0, 12) {real, imag} */,
  {32'hc1beab88, 32'hc1804f14} /* (5, 0, 11) {real, imag} */,
  {32'hc2b985ef, 32'h40d78f7a} /* (5, 0, 10) {real, imag} */,
  {32'hc256ff66, 32'hc212a288} /* (5, 0, 9) {real, imag} */,
  {32'hc2cd4224, 32'h42687d7e} /* (5, 0, 8) {real, imag} */,
  {32'hc23e221a, 32'h42357c78} /* (5, 0, 7) {real, imag} */,
  {32'h42663ac0, 32'h41cc8226} /* (5, 0, 6) {real, imag} */,
  {32'h42245372, 32'h41c9b2ec} /* (5, 0, 5) {real, imag} */,
  {32'h419d89bd, 32'h410c4644} /* (5, 0, 4) {real, imag} */,
  {32'h423d9aa1, 32'h42fd8eae} /* (5, 0, 3) {real, imag} */,
  {32'hc376bdef, 32'h42a54a12} /* (5, 0, 2) {real, imag} */,
  {32'h43cd35fa, 32'hc27b25ec} /* (5, 0, 1) {real, imag} */,
  {32'h42339501, 32'hc3abdc1f} /* (5, 0, 0) {real, imag} */,
  {32'h42bcfbde, 32'h44bb28fa} /* (4, 31, 31) {real, imag} */,
  {32'hc3b38e34, 32'hc44d263e} /* (4, 31, 30) {real, imag} */,
  {32'h4281b961, 32'hc3062f9d} /* (4, 31, 29) {real, imag} */,
  {32'h42edb640, 32'h432257ff} /* (4, 31, 28) {real, imag} */,
  {32'h4113f2c0, 32'hc357d8f6} /* (4, 31, 27) {real, imag} */,
  {32'h4211754b, 32'hc2f5da0c} /* (4, 31, 26) {real, imag} */,
  {32'h42f6ba1f, 32'h429f12ff} /* (4, 31, 25) {real, imag} */,
  {32'hc31ba9a4, 32'hc2ed08fa} /* (4, 31, 24) {real, imag} */,
  {32'h42776204, 32'h42e8d155} /* (4, 31, 23) {real, imag} */,
  {32'hc1a3b448, 32'h410f9e08} /* (4, 31, 22) {real, imag} */,
  {32'hc2986a52, 32'hc1c60220} /* (4, 31, 21) {real, imag} */,
  {32'hc01f3560, 32'h4292c754} /* (4, 31, 20) {real, imag} */,
  {32'h40ddcc28, 32'h40963270} /* (4, 31, 19) {real, imag} */,
  {32'hc291813e, 32'h4192f1f4} /* (4, 31, 18) {real, imag} */,
  {32'hc140d650, 32'hc190ca90} /* (4, 31, 17) {real, imag} */,
  {32'hc22d8e4c, 32'hc147e880} /* (4, 31, 16) {real, imag} */,
  {32'hc20d08ec, 32'h3fc07500} /* (4, 31, 15) {real, imag} */,
  {32'h3e926600, 32'hc2bc7b95} /* (4, 31, 14) {real, imag} */,
  {32'h41d9c5a2, 32'hc22971b0} /* (4, 31, 13) {real, imag} */,
  {32'hc17c5010, 32'h42322201} /* (4, 31, 12) {real, imag} */,
  {32'h432b5207, 32'h41c9ac80} /* (4, 31, 11) {real, imag} */,
  {32'hc2daf00a, 32'h42ea97f7} /* (4, 31, 10) {real, imag} */,
  {32'h421267e4, 32'hc24f4ba2} /* (4, 31, 9) {real, imag} */,
  {32'h42e04cd0, 32'hc290370e} /* (4, 31, 8) {real, imag} */,
  {32'hc245e962, 32'hc2446086} /* (4, 31, 7) {real, imag} */,
  {32'hc08c6aa8, 32'hc2c3cefc} /* (4, 31, 6) {real, imag} */,
  {32'h439330a4, 32'hc3a0450b} /* (4, 31, 5) {real, imag} */,
  {32'hc29ba728, 32'h42dcff02} /* (4, 31, 4) {real, imag} */,
  {32'h428514ef, 32'h422b73c3} /* (4, 31, 3) {real, imag} */,
  {32'h41784f50, 32'hc3d81cb3} /* (4, 31, 2) {real, imag} */,
  {32'hc3cb1df0, 32'h44782d1c} /* (4, 31, 1) {real, imag} */,
  {32'hc39c767e, 32'h443b3ea5} /* (4, 31, 0) {real, imag} */,
  {32'h43432aff, 32'hc41c75af} /* (4, 30, 31) {real, imag} */,
  {32'hc32b445e, 32'h43afc3ae} /* (4, 30, 30) {real, imag} */,
  {32'hc2082f83, 32'h42660626} /* (4, 30, 29) {real, imag} */,
  {32'h43740485, 32'hc39364a7} /* (4, 30, 28) {real, imag} */,
  {32'hc0e3bce0, 32'h43a3ca80} /* (4, 30, 27) {real, imag} */,
  {32'h430475c6, 32'hc2144bbd} /* (4, 30, 26) {real, imag} */,
  {32'hc2ad75f8, 32'hc2a3fab6} /* (4, 30, 25) {real, imag} */,
  {32'hc0ac7a00, 32'h42ca5304} /* (4, 30, 24) {real, imag} */,
  {32'h42551531, 32'h41dfb258} /* (4, 30, 23) {real, imag} */,
  {32'h41b104c2, 32'h42145f23} /* (4, 30, 22) {real, imag} */,
  {32'h42636bff, 32'h42f16a3e} /* (4, 30, 21) {real, imag} */,
  {32'hc2003ec2, 32'h3f616320} /* (4, 30, 20) {real, imag} */,
  {32'h41b2888e, 32'hc1373fbe} /* (4, 30, 19) {real, imag} */,
  {32'h40407f80, 32'h4251f7d4} /* (4, 30, 18) {real, imag} */,
  {32'h4211dfe5, 32'hc1ec6444} /* (4, 30, 17) {real, imag} */,
  {32'hc2517374, 32'hc23f56f0} /* (4, 30, 16) {real, imag} */,
  {32'h40f4ed98, 32'h410e1a88} /* (4, 30, 15) {real, imag} */,
  {32'hc28388b0, 32'hc22625f4} /* (4, 30, 14) {real, imag} */,
  {32'h4222a99f, 32'h3f12a920} /* (4, 30, 13) {real, imag} */,
  {32'h41eac62c, 32'h41f772ef} /* (4, 30, 12) {real, imag} */,
  {32'hc2a064e4, 32'h424b3df4} /* (4, 30, 11) {real, imag} */,
  {32'h42b69c78, 32'h42682cad} /* (4, 30, 10) {real, imag} */,
  {32'h427af963, 32'hc2c90d8e} /* (4, 30, 9) {real, imag} */,
  {32'hc2eb876c, 32'h430021a8} /* (4, 30, 8) {real, imag} */,
  {32'hc1b4b366, 32'hc2a3aaba} /* (4, 30, 7) {real, imag} */,
  {32'h405f9280, 32'h40d557e8} /* (4, 30, 6) {real, imag} */,
  {32'hc210219a, 32'hc24e84f8} /* (4, 30, 5) {real, imag} */,
  {32'h4385d968, 32'hc32ceafa} /* (4, 30, 4) {real, imag} */,
  {32'h4288ccbc, 32'hc2d5c679} /* (4, 30, 3) {real, imag} */,
  {32'hc3c13411, 32'h443a9ae3} /* (4, 30, 2) {real, imag} */,
  {32'h4373e313, 32'hc48d7812} /* (4, 30, 1) {real, imag} */,
  {32'h42a873ca, 32'hc41b8361} /* (4, 30, 0) {real, imag} */,
  {32'h4332816c, 32'h43ff804d} /* (4, 29, 31) {real, imag} */,
  {32'hc3446ffa, 32'hc35276ca} /* (4, 29, 30) {real, imag} */,
  {32'h429929c6, 32'h43586d70} /* (4, 29, 29) {real, imag} */,
  {32'hc31b6fa6, 32'hc2c95cf0} /* (4, 29, 28) {real, imag} */,
  {32'hc2961198, 32'h42dd3458} /* (4, 29, 27) {real, imag} */,
  {32'hc2b7b41b, 32'hc2a7ffb8} /* (4, 29, 26) {real, imag} */,
  {32'hc33cf209, 32'h424f2ef6} /* (4, 29, 25) {real, imag} */,
  {32'h414b1530, 32'h42c74cf9} /* (4, 29, 24) {real, imag} */,
  {32'h40d78100, 32'hc2a93f6b} /* (4, 29, 23) {real, imag} */,
  {32'hc23dceee, 32'hc29ca1fb} /* (4, 29, 22) {real, imag} */,
  {32'h4269e49a, 32'h4096f9de} /* (4, 29, 21) {real, imag} */,
  {32'h40768790, 32'hc1aecaf5} /* (4, 29, 20) {real, imag} */,
  {32'hc0972e20, 32'h41d21fe2} /* (4, 29, 19) {real, imag} */,
  {32'h4061fe98, 32'h419c6e38} /* (4, 29, 18) {real, imag} */,
  {32'h408d0090, 32'hc1bfdd4c} /* (4, 29, 17) {real, imag} */,
  {32'hc1b62730, 32'hc0f2518e} /* (4, 29, 16) {real, imag} */,
  {32'h4281d867, 32'hc0af5030} /* (4, 29, 15) {real, imag} */,
  {32'h4125d8ba, 32'hc1af0b98} /* (4, 29, 14) {real, imag} */,
  {32'h423a48d8, 32'h41be3026} /* (4, 29, 13) {real, imag} */,
  {32'hc198d6ca, 32'h3ffda130} /* (4, 29, 12) {real, imag} */,
  {32'h4219ca86, 32'hc0a611e2} /* (4, 29, 11) {real, imag} */,
  {32'h40ef2e90, 32'h4115f158} /* (4, 29, 10) {real, imag} */,
  {32'hc2b16f2b, 32'hc13b5068} /* (4, 29, 9) {real, imag} */,
  {32'hc325f113, 32'hc2c0a2eb} /* (4, 29, 8) {real, imag} */,
  {32'hc2f56f56, 32'h42687492} /* (4, 29, 7) {real, imag} */,
  {32'hc2d664c7, 32'hc2a5ac4e} /* (4, 29, 6) {real, imag} */,
  {32'h429db742, 32'hc24c48df} /* (4, 29, 5) {real, imag} */,
  {32'hbfe73540, 32'h42819b4e} /* (4, 29, 4) {real, imag} */,
  {32'h431b7be8, 32'h402b47a0} /* (4, 29, 3) {real, imag} */,
  {32'hc39ba0b6, 32'hc0dba610} /* (4, 29, 2) {real, imag} */,
  {32'h43e1f68e, 32'hc33763de} /* (4, 29, 1) {real, imag} */,
  {32'h433b49b4, 32'h41de5d40} /* (4, 29, 0) {real, imag} */,
  {32'h42c9ca8e, 32'h43dc9988} /* (4, 28, 31) {real, imag} */,
  {32'hc39cdeb8, 32'hc3a45102} /* (4, 28, 30) {real, imag} */,
  {32'hc2881e6d, 32'hc26de8d8} /* (4, 28, 29) {real, imag} */,
  {32'hbf309880, 32'h41c50254} /* (4, 28, 28) {real, imag} */,
  {32'hc352178a, 32'hc1ddfa60} /* (4, 28, 27) {real, imag} */,
  {32'hc21b4e12, 32'h41680ec4} /* (4, 28, 26) {real, imag} */,
  {32'h4226ae7e, 32'h4202837b} /* (4, 28, 25) {real, imag} */,
  {32'hc12d8028, 32'hc208c266} /* (4, 28, 24) {real, imag} */,
  {32'hc0686298, 32'h3f301250} /* (4, 28, 23) {real, imag} */,
  {32'h4314f5f8, 32'hc1bd9372} /* (4, 28, 22) {real, imag} */,
  {32'h4229afe5, 32'h4190aaf2} /* (4, 28, 21) {real, imag} */,
  {32'h420c7af0, 32'h40e99160} /* (4, 28, 20) {real, imag} */,
  {32'hc27a9974, 32'hc2197b39} /* (4, 28, 19) {real, imag} */,
  {32'hc1c3b16e, 32'hc092e704} /* (4, 28, 18) {real, imag} */,
  {32'h41fdb649, 32'h405ccaa0} /* (4, 28, 17) {real, imag} */,
  {32'h411b8058, 32'hc148aeb0} /* (4, 28, 16) {real, imag} */,
  {32'h40647a38, 32'h424c7a16} /* (4, 28, 15) {real, imag} */,
  {32'h42b5fc4c, 32'h425f6674} /* (4, 28, 14) {real, imag} */,
  {32'hc1fdd090, 32'hc176d4fc} /* (4, 28, 13) {real, imag} */,
  {32'h3effea40, 32'hc01ff480} /* (4, 28, 12) {real, imag} */,
  {32'hc206815f, 32'hc2a5fba8} /* (4, 28, 11) {real, imag} */,
  {32'hc1d99a7e, 32'hc0d74e88} /* (4, 28, 10) {real, imag} */,
  {32'hc181d12b, 32'hc1ac50c2} /* (4, 28, 9) {real, imag} */,
  {32'h42ba5a9b, 32'h40f38fb0} /* (4, 28, 8) {real, imag} */,
  {32'hc18ae93d, 32'hc28066c6} /* (4, 28, 7) {real, imag} */,
  {32'h422993dc, 32'h420f6df9} /* (4, 28, 6) {real, imag} */,
  {32'h40b58230, 32'hc338bc7c} /* (4, 28, 5) {real, imag} */,
  {32'h4292d2dd, 32'h43865b51} /* (4, 28, 4) {real, imag} */,
  {32'h428ee2ef, 32'h43229676} /* (4, 28, 3) {real, imag} */,
  {32'hc29ab660, 32'hc3162c14} /* (4, 28, 2) {real, imag} */,
  {32'h42b24026, 32'h4361d018} /* (4, 28, 1) {real, imag} */,
  {32'h42c6aa05, 32'h439b0ace} /* (4, 28, 0) {real, imag} */,
  {32'hc3273919, 32'hc3d50744} /* (4, 27, 31) {real, imag} */,
  {32'h43178ee4, 32'h4333ba46} /* (4, 27, 30) {real, imag} */,
  {32'hc1af0b55, 32'h42e93b77} /* (4, 27, 29) {real, imag} */,
  {32'hc25ef40c, 32'hc2df9942} /* (4, 27, 28) {real, imag} */,
  {32'h42ceb339, 32'hc20cdd4b} /* (4, 27, 27) {real, imag} */,
  {32'h425a23f5, 32'h42e6e3d4} /* (4, 27, 26) {real, imag} */,
  {32'hc2cf902d, 32'hc181ab5c} /* (4, 27, 25) {real, imag} */,
  {32'h41d00de0, 32'hc126fd2c} /* (4, 27, 24) {real, imag} */,
  {32'hc2035136, 32'hc1995a1a} /* (4, 27, 23) {real, imag} */,
  {32'h3fcc9790, 32'h420a9feb} /* (4, 27, 22) {real, imag} */,
  {32'hc1b57205, 32'hc20c2c37} /* (4, 27, 21) {real, imag} */,
  {32'hc1eb5237, 32'hc22c107c} /* (4, 27, 20) {real, imag} */,
  {32'hc22f3ad7, 32'hc1f19f73} /* (4, 27, 19) {real, imag} */,
  {32'h403a6e38, 32'hc1448595} /* (4, 27, 18) {real, imag} */,
  {32'h41026610, 32'hc0178f48} /* (4, 27, 17) {real, imag} */,
  {32'h401a9888, 32'hc1990478} /* (4, 27, 16) {real, imag} */,
  {32'hc22410c4, 32'h4082d3a4} /* (4, 27, 15) {real, imag} */,
  {32'hc196a0d9, 32'h4185c7f2} /* (4, 27, 14) {real, imag} */,
  {32'h4219822d, 32'h41957af9} /* (4, 27, 13) {real, imag} */,
  {32'hc0d44234, 32'h413d89af} /* (4, 27, 12) {real, imag} */,
  {32'hc21a4f88, 32'h42a0e766} /* (4, 27, 11) {real, imag} */,
  {32'hbfd5ceb0, 32'h40b31bf8} /* (4, 27, 10) {real, imag} */,
  {32'hc1f83f24, 32'h42405159} /* (4, 27, 9) {real, imag} */,
  {32'h427cb314, 32'hc24b9c3f} /* (4, 27, 8) {real, imag} */,
  {32'hc2e753bb, 32'hc2653f26} /* (4, 27, 7) {real, imag} */,
  {32'h4206a2c7, 32'hc2f1ec7e} /* (4, 27, 6) {real, imag} */,
  {32'hc265fc1e, 32'h42b95de6} /* (4, 27, 5) {real, imag} */,
  {32'hc228ae92, 32'h422bbf90} /* (4, 27, 4) {real, imag} */,
  {32'h405af558, 32'hc294c7c9} /* (4, 27, 3) {real, imag} */,
  {32'hc259c804, 32'h4336cf6a} /* (4, 27, 2) {real, imag} */,
  {32'h43ce41d8, 32'hc3b4d8cc} /* (4, 27, 1) {real, imag} */,
  {32'hc24073f8, 32'hc38dfd5c} /* (4, 27, 0) {real, imag} */,
  {32'h42a0e1c2, 32'hc31f9cfa} /* (4, 26, 31) {real, imag} */,
  {32'h4253c317, 32'h4156a488} /* (4, 26, 30) {real, imag} */,
  {32'hc19b614a, 32'hc266197e} /* (4, 26, 29) {real, imag} */,
  {32'h42c3a942, 32'h41a1b694} /* (4, 26, 28) {real, imag} */,
  {32'h4269c1df, 32'hc296d57e} /* (4, 26, 27) {real, imag} */,
  {32'h41ee4528, 32'hc3143e2e} /* (4, 26, 26) {real, imag} */,
  {32'hbfc5d470, 32'hc1ddead0} /* (4, 26, 25) {real, imag} */,
  {32'h421334bc, 32'h42093238} /* (4, 26, 24) {real, imag} */,
  {32'h42d1f914, 32'h3e94fc80} /* (4, 26, 23) {real, imag} */,
  {32'hc1159660, 32'hc1c88e45} /* (4, 26, 22) {real, imag} */,
  {32'h4244950e, 32'hbf975880} /* (4, 26, 21) {real, imag} */,
  {32'hbeb190a0, 32'h3f843080} /* (4, 26, 20) {real, imag} */,
  {32'hc1b11aae, 32'h42499172} /* (4, 26, 19) {real, imag} */,
  {32'h420c9b02, 32'hc200760a} /* (4, 26, 18) {real, imag} */,
  {32'h41987420, 32'hc1000410} /* (4, 26, 17) {real, imag} */,
  {32'h40235d40, 32'hc146ef24} /* (4, 26, 16) {real, imag} */,
  {32'hc1c1ea18, 32'hc1e6fb50} /* (4, 26, 15) {real, imag} */,
  {32'h41483250, 32'h421092be} /* (4, 26, 14) {real, imag} */,
  {32'hc1b83df6, 32'hc1582e02} /* (4, 26, 13) {real, imag} */,
  {32'h3fc68b68, 32'hc1da01b8} /* (4, 26, 12) {real, imag} */,
  {32'h409c4360, 32'hc2a1b896} /* (4, 26, 11) {real, imag} */,
  {32'hc24fade6, 32'hc1ecd0db} /* (4, 26, 10) {real, imag} */,
  {32'hc2098e74, 32'hc1a1a230} /* (4, 26, 9) {real, imag} */,
  {32'h4153c086, 32'h42fe3c62} /* (4, 26, 8) {real, imag} */,
  {32'h42398278, 32'hc206b4e1} /* (4, 26, 7) {real, imag} */,
  {32'hc288be23, 32'hc3301496} /* (4, 26, 6) {real, imag} */,
  {32'h431805b6, 32'hc19c79b8} /* (4, 26, 5) {real, imag} */,
  {32'h422e3535, 32'hc3087a24} /* (4, 26, 4) {real, imag} */,
  {32'hc2a64d34, 32'h4211e968} /* (4, 26, 3) {real, imag} */,
  {32'hc32f2c4a, 32'h420caf86} /* (4, 26, 2) {real, imag} */,
  {32'h4303049c, 32'hc18e8568} /* (4, 26, 1) {real, imag} */,
  {32'hc2c4f972, 32'h42bb9902} /* (4, 26, 0) {real, imag} */,
  {32'hc228ecfb, 32'hc117ffab} /* (4, 25, 31) {real, imag} */,
  {32'hc323431a, 32'h43541684} /* (4, 25, 30) {real, imag} */,
  {32'hc20d1d39, 32'hc2adcdc0} /* (4, 25, 29) {real, imag} */,
  {32'h42ff0b43, 32'hc2850522} /* (4, 25, 28) {real, imag} */,
  {32'hc13a5468, 32'h42e10de4} /* (4, 25, 27) {real, imag} */,
  {32'hc2269843, 32'h414c2780} /* (4, 25, 26) {real, imag} */,
  {32'hc1b3fbf0, 32'h428d2a4b} /* (4, 25, 25) {real, imag} */,
  {32'hc1009df8, 32'hc20270ce} /* (4, 25, 24) {real, imag} */,
  {32'hc2523aa0, 32'hc23fe946} /* (4, 25, 23) {real, imag} */,
  {32'h41aa5edc, 32'h419ec5ce} /* (4, 25, 22) {real, imag} */,
  {32'h426cf6a8, 32'hc1a76526} /* (4, 25, 21) {real, imag} */,
  {32'hc1c0ab52, 32'hc16d6fc3} /* (4, 25, 20) {real, imag} */,
  {32'h421c7a89, 32'h40440310} /* (4, 25, 19) {real, imag} */,
  {32'h41fbb96d, 32'hc19ad70c} /* (4, 25, 18) {real, imag} */,
  {32'hc169ee65, 32'hc0ab893e} /* (4, 25, 17) {real, imag} */,
  {32'hc1cf3363, 32'h41a1f68e} /* (4, 25, 16) {real, imag} */,
  {32'h4169dd21, 32'h41e575d0} /* (4, 25, 15) {real, imag} */,
  {32'hc19fce6f, 32'h41ea2b3c} /* (4, 25, 14) {real, imag} */,
  {32'h4145b2ff, 32'h4207670f} /* (4, 25, 13) {real, imag} */,
  {32'hc271a2bb, 32'hc18be916} /* (4, 25, 12) {real, imag} */,
  {32'hc1fee72c, 32'h41360cbc} /* (4, 25, 11) {real, imag} */,
  {32'h3fa8fbb8, 32'hc1ad29c4} /* (4, 25, 10) {real, imag} */,
  {32'hc1be918c, 32'h422ef9ee} /* (4, 25, 9) {real, imag} */,
  {32'h430ff3c0, 32'h413b9f02} /* (4, 25, 8) {real, imag} */,
  {32'hc0c0cd3c, 32'h41daccb4} /* (4, 25, 7) {real, imag} */,
  {32'h42a59a06, 32'hc2490a1f} /* (4, 25, 6) {real, imag} */,
  {32'hc26943b4, 32'h416ec56c} /* (4, 25, 5) {real, imag} */,
  {32'hc283e131, 32'hc2fedf5c} /* (4, 25, 4) {real, imag} */,
  {32'hc1c280e4, 32'h41a5ce92} /* (4, 25, 3) {real, imag} */,
  {32'h42d5bbc0, 32'h41e5d76c} /* (4, 25, 2) {real, imag} */,
  {32'hc287ace6, 32'hc2138cf1} /* (4, 25, 1) {real, imag} */,
  {32'h41d42437, 32'h41a7e1b6} /* (4, 25, 0) {real, imag} */,
  {32'hc274d560, 32'hc360fa30} /* (4, 24, 31) {real, imag} */,
  {32'h42d50679, 32'h426886ca} /* (4, 24, 30) {real, imag} */,
  {32'hc2fb657a, 32'h41823571} /* (4, 24, 29) {real, imag} */,
  {32'hc19a78aa, 32'hc2694a9e} /* (4, 24, 28) {real, imag} */,
  {32'h422641c0, 32'hc2cb73ae} /* (4, 24, 27) {real, imag} */,
  {32'h41e7528d, 32'h4238c7da} /* (4, 24, 26) {real, imag} */,
  {32'h41f1b55c, 32'hc28d67fa} /* (4, 24, 25) {real, imag} */,
  {32'h41c1a968, 32'h42a96aad} /* (4, 24, 24) {real, imag} */,
  {32'h420f86ce, 32'hc1fdab14} /* (4, 24, 23) {real, imag} */,
  {32'h41d9b6d9, 32'hc1a1be3c} /* (4, 24, 22) {real, imag} */,
  {32'h404ff190, 32'hc068a700} /* (4, 24, 21) {real, imag} */,
  {32'hc040799c, 32'hc244d5f4} /* (4, 24, 20) {real, imag} */,
  {32'hc106ebea, 32'h413016ca} /* (4, 24, 19) {real, imag} */,
  {32'hc196f95e, 32'h414dc088} /* (4, 24, 18) {real, imag} */,
  {32'h40de2a27, 32'h41561e36} /* (4, 24, 17) {real, imag} */,
  {32'h411d78c0, 32'hc0668a60} /* (4, 24, 16) {real, imag} */,
  {32'h408f5d09, 32'h4140265a} /* (4, 24, 15) {real, imag} */,
  {32'hc184372a, 32'hc13c4c38} /* (4, 24, 14) {real, imag} */,
  {32'hc18b76bd, 32'hbf9c78d0} /* (4, 24, 13) {real, imag} */,
  {32'hc18978ea, 32'hc2bf2922} /* (4, 24, 12) {real, imag} */,
  {32'hc14af67c, 32'h41c0482c} /* (4, 24, 11) {real, imag} */,
  {32'h41c15c7d, 32'h42a9de3f} /* (4, 24, 10) {real, imag} */,
  {32'h423faf7a, 32'hc1aeda98} /* (4, 24, 9) {real, imag} */,
  {32'hc2c3a590, 32'h423c876e} /* (4, 24, 8) {real, imag} */,
  {32'h41331794, 32'hc1f4005e} /* (4, 24, 7) {real, imag} */,
  {32'hc29f4e7a, 32'h42c8aaf7} /* (4, 24, 6) {real, imag} */,
  {32'h4204296c, 32'h40ec8f70} /* (4, 24, 5) {real, imag} */,
  {32'hc0b2077e, 32'hc186f740} /* (4, 24, 4) {real, imag} */,
  {32'h41e50378, 32'h428ebdf2} /* (4, 24, 3) {real, imag} */,
  {32'hc2c484fb, 32'h4344d7f0} /* (4, 24, 2) {real, imag} */,
  {32'hc29bd6d8, 32'hc383e95e} /* (4, 24, 1) {real, imag} */,
  {32'hc2cba094, 32'hc36f9798} /* (4, 24, 0) {real, imag} */,
  {32'h422695b5, 32'h413bb026} /* (4, 23, 31) {real, imag} */,
  {32'hc23d0820, 32'hc3017c20} /* (4, 23, 30) {real, imag} */,
  {32'hc0f876b2, 32'hc0a07070} /* (4, 23, 29) {real, imag} */,
  {32'h429efbca, 32'h42164b17} /* (4, 23, 28) {real, imag} */,
  {32'hc289c221, 32'h42c5b894} /* (4, 23, 27) {real, imag} */,
  {32'hc1a4d14a, 32'hc1a7a880} /* (4, 23, 26) {real, imag} */,
  {32'hc2248615, 32'h41bc9d74} /* (4, 23, 25) {real, imag} */,
  {32'h424cb445, 32'h401f5c7c} /* (4, 23, 24) {real, imag} */,
  {32'h3fb4f0e8, 32'h422ab5d6} /* (4, 23, 23) {real, imag} */,
  {32'hc1ffe78e, 32'hc2156806} /* (4, 23, 22) {real, imag} */,
  {32'hc2056647, 32'h41a99456} /* (4, 23, 21) {real, imag} */,
  {32'h41572cd2, 32'h415ea8f6} /* (4, 23, 20) {real, imag} */,
  {32'h41fe2813, 32'hbe96bc00} /* (4, 23, 19) {real, imag} */,
  {32'hbf951ad0, 32'h416ad95c} /* (4, 23, 18) {real, imag} */,
  {32'hc11a236e, 32'h40b943ba} /* (4, 23, 17) {real, imag} */,
  {32'h407542e8, 32'hc16f97d0} /* (4, 23, 16) {real, imag} */,
  {32'hc105dcba, 32'hc1822020} /* (4, 23, 15) {real, imag} */,
  {32'hc03988b8, 32'hc1a7b4ce} /* (4, 23, 14) {real, imag} */,
  {32'hc12ef932, 32'h3fbbf9a0} /* (4, 23, 13) {real, imag} */,
  {32'h41268776, 32'h420fdc26} /* (4, 23, 12) {real, imag} */,
  {32'h41e9fbb3, 32'hc241b27d} /* (4, 23, 11) {real, imag} */,
  {32'h429f30f0, 32'hc1907dfc} /* (4, 23, 10) {real, imag} */,
  {32'hc1953d96, 32'h40739440} /* (4, 23, 9) {real, imag} */,
  {32'h412bf2c0, 32'h41891008} /* (4, 23, 8) {real, imag} */,
  {32'hc223309f, 32'h4291d9b8} /* (4, 23, 7) {real, imag} */,
  {32'h42789e1f, 32'h42a07470} /* (4, 23, 6) {real, imag} */,
  {32'h4243ab66, 32'hc2bdbd60} /* (4, 23, 5) {real, imag} */,
  {32'h42c776d6, 32'h42357a41} /* (4, 23, 4) {real, imag} */,
  {32'hc1fc65ce, 32'hc2b374cf} /* (4, 23, 3) {real, imag} */,
  {32'hc3226a58, 32'h41eef744} /* (4, 23, 2) {real, imag} */,
  {32'h42226929, 32'h426ab84a} /* (4, 23, 1) {real, imag} */,
  {32'h424592d8, 32'h425c403c} /* (4, 23, 0) {real, imag} */,
  {32'h418b3818, 32'h42d55529} /* (4, 22, 31) {real, imag} */,
  {32'hc27a8547, 32'hc28b1f18} /* (4, 22, 30) {real, imag} */,
  {32'hc05000a0, 32'hc202cafc} /* (4, 22, 29) {real, imag} */,
  {32'hc23d7614, 32'h421a4f13} /* (4, 22, 28) {real, imag} */,
  {32'hc23d1ad6, 32'hc1dc7101} /* (4, 22, 27) {real, imag} */,
  {32'h3f44a3e8, 32'hc26cc109} /* (4, 22, 26) {real, imag} */,
  {32'h428c022b, 32'h42561d96} /* (4, 22, 25) {real, imag} */,
  {32'hbff10bc0, 32'hbd81ed00} /* (4, 22, 24) {real, imag} */,
  {32'h418dae5e, 32'h42245d06} /* (4, 22, 23) {real, imag} */,
  {32'h4195a14a, 32'hc0779420} /* (4, 22, 22) {real, imag} */,
  {32'hc1b5a9b5, 32'h41fab617} /* (4, 22, 21) {real, imag} */,
  {32'h41f4c5b1, 32'hc10344c5} /* (4, 22, 20) {real, imag} */,
  {32'h4253918d, 32'h41876a83} /* (4, 22, 19) {real, imag} */,
  {32'hc14196b7, 32'hc148a786} /* (4, 22, 18) {real, imag} */,
  {32'hc10ea253, 32'h416121fa} /* (4, 22, 17) {real, imag} */,
  {32'hc181c392, 32'hc1a68d0e} /* (4, 22, 16) {real, imag} */,
  {32'hbf822258, 32'hc0fd5574} /* (4, 22, 15) {real, imag} */,
  {32'hc12ede21, 32'h4078a218} /* (4, 22, 14) {real, imag} */,
  {32'h411353bc, 32'h4113b242} /* (4, 22, 13) {real, imag} */,
  {32'h40187f38, 32'h41de2e0a} /* (4, 22, 12) {real, imag} */,
  {32'hc15bc12e, 32'hc0fcb0bc} /* (4, 22, 11) {real, imag} */,
  {32'hc175994c, 32'hbf5b5680} /* (4, 22, 10) {real, imag} */,
  {32'h41fb33c4, 32'h4213743c} /* (4, 22, 9) {real, imag} */,
  {32'hc1895b70, 32'h4140f97a} /* (4, 22, 8) {real, imag} */,
  {32'h41b4ac0b, 32'h41d714bf} /* (4, 22, 7) {real, imag} */,
  {32'hc1724fc0, 32'h413753dc} /* (4, 22, 6) {real, imag} */,
  {32'hc0f8a7e4, 32'h41175a5a} /* (4, 22, 5) {real, imag} */,
  {32'hc26be6b0, 32'h420871e9} /* (4, 22, 4) {real, imag} */,
  {32'hc2934b9f, 32'h428f9f5a} /* (4, 22, 3) {real, imag} */,
  {32'hc2640ef3, 32'hc2f5b14c} /* (4, 22, 2) {real, imag} */,
  {32'hc201589e, 32'h42563cf6} /* (4, 22, 1) {real, imag} */,
  {32'h42b30e7e, 32'hc2dfaae8} /* (4, 22, 0) {real, imag} */,
  {32'hc255d4f2, 32'hc191e996} /* (4, 21, 31) {real, imag} */,
  {32'h43189d6c, 32'h41fbbc26} /* (4, 21, 30) {real, imag} */,
  {32'hc29fb8a7, 32'h428d10e9} /* (4, 21, 29) {real, imag} */,
  {32'h4109132b, 32'hc2013432} /* (4, 21, 28) {real, imag} */,
  {32'h41e6b351, 32'h421cb460} /* (4, 21, 27) {real, imag} */,
  {32'h420ad97a, 32'hc1160b03} /* (4, 21, 26) {real, imag} */,
  {32'hc1cfc34c, 32'h420eb656} /* (4, 21, 25) {real, imag} */,
  {32'hc1d85dd6, 32'hc1f0b739} /* (4, 21, 24) {real, imag} */,
  {32'hc1605a04, 32'h406a90c8} /* (4, 21, 23) {real, imag} */,
  {32'hc2184bce, 32'hc1c76892} /* (4, 21, 22) {real, imag} */,
  {32'h41147e2c, 32'hc19d9009} /* (4, 21, 21) {real, imag} */,
  {32'h413a7344, 32'h411ee2c7} /* (4, 21, 20) {real, imag} */,
  {32'hbf78c720, 32'h41a41826} /* (4, 21, 19) {real, imag} */,
  {32'hc0b8a038, 32'hc002403c} /* (4, 21, 18) {real, imag} */,
  {32'h40e624a4, 32'hc0583d4c} /* (4, 21, 17) {real, imag} */,
  {32'h41a1ea46, 32'hc11f3cd4} /* (4, 21, 16) {real, imag} */,
  {32'hc10e0bb6, 32'hc0dbcb92} /* (4, 21, 15) {real, imag} */,
  {32'h413ce3ac, 32'hbf5786d0} /* (4, 21, 14) {real, imag} */,
  {32'hc1570cc2, 32'h408884b8} /* (4, 21, 13) {real, imag} */,
  {32'h40f88ec1, 32'hbf4ea8b0} /* (4, 21, 12) {real, imag} */,
  {32'h41185294, 32'h4166ec66} /* (4, 21, 11) {real, imag} */,
  {32'hc1ab1dd5, 32'hc1ee88fa} /* (4, 21, 10) {real, imag} */,
  {32'h41d6d7bc, 32'h41847f15} /* (4, 21, 9) {real, imag} */,
  {32'h41a494a2, 32'hc17a7876} /* (4, 21, 8) {real, imag} */,
  {32'hc18eae0a, 32'hc234d8f0} /* (4, 21, 7) {real, imag} */,
  {32'h423a3a0e, 32'h41b85cde} /* (4, 21, 6) {real, imag} */,
  {32'hc1a23467, 32'h42956090} /* (4, 21, 5) {real, imag} */,
  {32'h40fcfd4b, 32'hc12424f7} /* (4, 21, 4) {real, imag} */,
  {32'h41f2c277, 32'hc23b4a5e} /* (4, 21, 3) {real, imag} */,
  {32'h42e971b9, 32'h420eb975} /* (4, 21, 2) {real, imag} */,
  {32'h40e5028c, 32'hc28c3900} /* (4, 21, 1) {real, imag} */,
  {32'hc2cb9d0a, 32'hc2463f29} /* (4, 21, 0) {real, imag} */,
  {32'h422882d7, 32'h41baf9d6} /* (4, 20, 31) {real, imag} */,
  {32'h3fded940, 32'h3e32de70} /* (4, 20, 30) {real, imag} */,
  {32'hc2402bfb, 32'h41985ccf} /* (4, 20, 29) {real, imag} */,
  {32'hc0e3dbfb, 32'h41e777c8} /* (4, 20, 28) {real, imag} */,
  {32'h411dcef1, 32'hc249ddb8} /* (4, 20, 27) {real, imag} */,
  {32'h40d077fd, 32'h41494ba5} /* (4, 20, 26) {real, imag} */,
  {32'h41878914, 32'h4129b9fe} /* (4, 20, 25) {real, imag} */,
  {32'h420f2090, 32'hc1f8b868} /* (4, 20, 24) {real, imag} */,
  {32'hc015c80b, 32'h41e374ee} /* (4, 20, 23) {real, imag} */,
  {32'h40adc74d, 32'hc0d0b220} /* (4, 20, 22) {real, imag} */,
  {32'h411e010e, 32'hc0d2891c} /* (4, 20, 21) {real, imag} */,
  {32'hc0101ff8, 32'h4172fa44} /* (4, 20, 20) {real, imag} */,
  {32'hc19f6952, 32'h3f151d20} /* (4, 20, 19) {real, imag} */,
  {32'hc051dd90, 32'hc13080ae} /* (4, 20, 18) {real, imag} */,
  {32'hc0e8a2f4, 32'hc142592a} /* (4, 20, 17) {real, imag} */,
  {32'h3fc467e0, 32'h40c13ff8} /* (4, 20, 16) {real, imag} */,
  {32'hc1029be2, 32'h41871f2b} /* (4, 20, 15) {real, imag} */,
  {32'hc104b614, 32'hc167fe0a} /* (4, 20, 14) {real, imag} */,
  {32'h408a02d6, 32'hc127b1b6} /* (4, 20, 13) {real, imag} */,
  {32'hc0e0893e, 32'hc1837368} /* (4, 20, 12) {real, imag} */,
  {32'hc1419aec, 32'h42384e1a} /* (4, 20, 11) {real, imag} */,
  {32'h4015456e, 32'hc230ed9a} /* (4, 20, 10) {real, imag} */,
  {32'h4071a473, 32'hc1c5f7b0} /* (4, 20, 9) {real, imag} */,
  {32'hc24ec5aa, 32'h40edc880} /* (4, 20, 8) {real, imag} */,
  {32'h41b01484, 32'hc2047006} /* (4, 20, 7) {real, imag} */,
  {32'h419b597e, 32'h415bacdd} /* (4, 20, 6) {real, imag} */,
  {32'hc1f68674, 32'h42b45424} /* (4, 20, 5) {real, imag} */,
  {32'hc1aab72f, 32'h41321fdc} /* (4, 20, 4) {real, imag} */,
  {32'hc073f1f0, 32'h423019a4} /* (4, 20, 3) {real, imag} */,
  {32'h430d5c10, 32'h4079bdcd} /* (4, 20, 2) {real, imag} */,
  {32'hc2004123, 32'hc13b3934} /* (4, 20, 1) {real, imag} */,
  {32'h420bfdc7, 32'hc1b33d36} /* (4, 20, 0) {real, imag} */,
  {32'hc1337084, 32'h421453bb} /* (4, 19, 31) {real, imag} */,
  {32'hc24b999d, 32'h41834668} /* (4, 19, 30) {real, imag} */,
  {32'h4206eb2a, 32'hc1e45c0a} /* (4, 19, 29) {real, imag} */,
  {32'hc2395ece, 32'h4268e54c} /* (4, 19, 28) {real, imag} */,
  {32'hc08f9185, 32'hc25235de} /* (4, 19, 27) {real, imag} */,
  {32'h42120d58, 32'h4090f261} /* (4, 19, 26) {real, imag} */,
  {32'h40eb0031, 32'hc1c9082f} /* (4, 19, 25) {real, imag} */,
  {32'h421cabe7, 32'h41a35310} /* (4, 19, 24) {real, imag} */,
  {32'hc18d205a, 32'h402e136a} /* (4, 19, 23) {real, imag} */,
  {32'h41d118e7, 32'hc1f8ccc9} /* (4, 19, 22) {real, imag} */,
  {32'hc1290814, 32'hc0a8cffc} /* (4, 19, 21) {real, imag} */,
  {32'hc0f03c42, 32'hc1205d44} /* (4, 19, 20) {real, imag} */,
  {32'h40b92ff4, 32'h3fe7b114} /* (4, 19, 19) {real, imag} */,
  {32'hc08209d2, 32'h4086843c} /* (4, 19, 18) {real, imag} */,
  {32'h3e194bd0, 32'hc131b462} /* (4, 19, 17) {real, imag} */,
  {32'h4126a8f8, 32'h411b06d7} /* (4, 19, 16) {real, imag} */,
  {32'h40ae6b86, 32'hc1711fa6} /* (4, 19, 15) {real, imag} */,
  {32'hbe961460, 32'hc1a3f522} /* (4, 19, 14) {real, imag} */,
  {32'hc15f99d6, 32'hc171bbac} /* (4, 19, 13) {real, imag} */,
  {32'h40b5da12, 32'h413b02e8} /* (4, 19, 12) {real, imag} */,
  {32'hc1fd7c1e, 32'h415023d4} /* (4, 19, 11) {real, imag} */,
  {32'hc2214259, 32'hbfe0eb30} /* (4, 19, 10) {real, imag} */,
  {32'hc188e456, 32'h408758bb} /* (4, 19, 9) {real, imag} */,
  {32'h41619611, 32'hc0df9b08} /* (4, 19, 8) {real, imag} */,
  {32'hbfb1d7ec, 32'hc204b992} /* (4, 19, 7) {real, imag} */,
  {32'h40326250, 32'h4108f108} /* (4, 19, 6) {real, imag} */,
  {32'h41a01ff9, 32'hc13762b0} /* (4, 19, 5) {real, imag} */,
  {32'hc0d6e870, 32'h40104da8} /* (4, 19, 4) {real, imag} */,
  {32'h4246fa06, 32'hc02aeb1c} /* (4, 19, 3) {real, imag} */,
  {32'hc1f86896, 32'hc238eb5a} /* (4, 19, 2) {real, imag} */,
  {32'h41aa9332, 32'hc08b32b8} /* (4, 19, 1) {real, imag} */,
  {32'h424382bd, 32'h40e21602} /* (4, 19, 0) {real, imag} */,
  {32'h4212e12b, 32'hc209ead3} /* (4, 18, 31) {real, imag} */,
  {32'h41e8b6e4, 32'h42564630} /* (4, 18, 30) {real, imag} */,
  {32'h409eb44a, 32'h4194d078} /* (4, 18, 29) {real, imag} */,
  {32'h41e44f1a, 32'hc1e933a5} /* (4, 18, 28) {real, imag} */,
  {32'h41f48f75, 32'h4021e45d} /* (4, 18, 27) {real, imag} */,
  {32'h42135220, 32'h41955e4a} /* (4, 18, 26) {real, imag} */,
  {32'h41a750f4, 32'hc0f3aa25} /* (4, 18, 25) {real, imag} */,
  {32'hc1f81cac, 32'h41a10a3a} /* (4, 18, 24) {real, imag} */,
  {32'h401c9bd0, 32'h417b59b9} /* (4, 18, 23) {real, imag} */,
  {32'hc234699a, 32'h41b26794} /* (4, 18, 22) {real, imag} */,
  {32'h4149e050, 32'h409195a6} /* (4, 18, 21) {real, imag} */,
  {32'hc05f970e, 32'hbc90d300} /* (4, 18, 20) {real, imag} */,
  {32'hc0b86cea, 32'h3bb54400} /* (4, 18, 19) {real, imag} */,
  {32'h40182838, 32'hbfe049f0} /* (4, 18, 18) {real, imag} */,
  {32'hc13ab164, 32'h411cf10d} /* (4, 18, 17) {real, imag} */,
  {32'hc04f9d48, 32'hc09366b2} /* (4, 18, 16) {real, imag} */,
  {32'hc04f7c82, 32'hc0f6afa2} /* (4, 18, 15) {real, imag} */,
  {32'hc0b56c80, 32'hc1211f10} /* (4, 18, 14) {real, imag} */,
  {32'h411d3a4f, 32'h40a3ae9f} /* (4, 18, 13) {real, imag} */,
  {32'h412850f2, 32'hc101127e} /* (4, 18, 12) {real, imag} */,
  {32'hc10a6d14, 32'hc0eb4c34} /* (4, 18, 11) {real, imag} */,
  {32'h4112257c, 32'hc199eb18} /* (4, 18, 10) {real, imag} */,
  {32'h412e2cb6, 32'hc0f2d43e} /* (4, 18, 9) {real, imag} */,
  {32'hc1b941a2, 32'hc19d422e} /* (4, 18, 8) {real, imag} */,
  {32'hc2085c10, 32'h3ea2df90} /* (4, 18, 7) {real, imag} */,
  {32'h425fe590, 32'h423c1499} /* (4, 18, 6) {real, imag} */,
  {32'hc12e0e42, 32'hc06d72df} /* (4, 18, 5) {real, imag} */,
  {32'h41e4f0b6, 32'h410d15ea} /* (4, 18, 4) {real, imag} */,
  {32'h40f18352, 32'hc18a8004} /* (4, 18, 3) {real, imag} */,
  {32'h419882e0, 32'hc1438b20} /* (4, 18, 2) {real, imag} */,
  {32'hc288b9a8, 32'hc0b6c586} /* (4, 18, 1) {real, imag} */,
  {32'hc243eff4, 32'hc2043efe} /* (4, 18, 0) {real, imag} */,
  {32'h42141b30, 32'h421346f8} /* (4, 17, 31) {real, imag} */,
  {32'h40a0d90a, 32'hc0a878a7} /* (4, 17, 30) {real, imag} */,
  {32'hc1873f22, 32'hc2449480} /* (4, 17, 29) {real, imag} */,
  {32'h410dc397, 32'hc17df720} /* (4, 17, 28) {real, imag} */,
  {32'hc12ba6bd, 32'hc1d78fff} /* (4, 17, 27) {real, imag} */,
  {32'hc1947571, 32'hc12421ae} /* (4, 17, 26) {real, imag} */,
  {32'hc11c1abe, 32'hc20059d8} /* (4, 17, 25) {real, imag} */,
  {32'hc15e0af7, 32'h41de61a7} /* (4, 17, 24) {real, imag} */,
  {32'hc115b7eb, 32'h411569bb} /* (4, 17, 23) {real, imag} */,
  {32'hc0bf989e, 32'hbeb96a60} /* (4, 17, 22) {real, imag} */,
  {32'h41e0f5c4, 32'h413a5376} /* (4, 17, 21) {real, imag} */,
  {32'hc147f59e, 32'h4191e5ee} /* (4, 17, 20) {real, imag} */,
  {32'h41010a84, 32'hc0900d84} /* (4, 17, 19) {real, imag} */,
  {32'h4154ba55, 32'hbfc9d1f0} /* (4, 17, 18) {real, imag} */,
  {32'h40df1c8c, 32'h405de1b0} /* (4, 17, 17) {real, imag} */,
  {32'hc075b496, 32'h3f5edc80} /* (4, 17, 16) {real, imag} */,
  {32'h3f885f60, 32'h414c98b2} /* (4, 17, 15) {real, imag} */,
  {32'h40aeb2ea, 32'hc0d541ea} /* (4, 17, 14) {real, imag} */,
  {32'hc109d352, 32'hc1a2af53} /* (4, 17, 13) {real, imag} */,
  {32'h41bafeb5, 32'hc04deaf4} /* (4, 17, 12) {real, imag} */,
  {32'hc1146371, 32'h3de79880} /* (4, 17, 11) {real, imag} */,
  {32'hc0026d34, 32'h404f15fc} /* (4, 17, 10) {real, imag} */,
  {32'h402ebb25, 32'h4135c6ef} /* (4, 17, 9) {real, imag} */,
  {32'hc11e6645, 32'h41e8647d} /* (4, 17, 8) {real, imag} */,
  {32'hc0cb1b59, 32'hc18c32bc} /* (4, 17, 7) {real, imag} */,
  {32'h414a740c, 32'hc23ac4f4} /* (4, 17, 6) {real, imag} */,
  {32'h41f2bc76, 32'h405600f8} /* (4, 17, 5) {real, imag} */,
  {32'h41988a52, 32'hc14dcc02} /* (4, 17, 4) {real, imag} */,
  {32'h3fbbdecc, 32'h4283c130} /* (4, 17, 3) {real, imag} */,
  {32'h412951e5, 32'h413ce4f8} /* (4, 17, 2) {real, imag} */,
  {32'h40a52472, 32'h414aacef} /* (4, 17, 1) {real, imag} */,
  {32'hc150c096, 32'hc20dec9c} /* (4, 17, 0) {real, imag} */,
  {32'h41eae03b, 32'h40b18aa2} /* (4, 16, 31) {real, imag} */,
  {32'h4189ff48, 32'hc1b007eb} /* (4, 16, 30) {real, imag} */,
  {32'h418492bc, 32'h41e2cf56} /* (4, 16, 29) {real, imag} */,
  {32'hc0bd3bc4, 32'hc215f2c0} /* (4, 16, 28) {real, imag} */,
  {32'hc258f2c6, 32'hc03f4ab8} /* (4, 16, 27) {real, imag} */,
  {32'h40c3ba59, 32'h41bc9ed2} /* (4, 16, 26) {real, imag} */,
  {32'hc12bea6a, 32'h418b3990} /* (4, 16, 25) {real, imag} */,
  {32'hc0cc0988, 32'h41db2132} /* (4, 16, 24) {real, imag} */,
  {32'hc1b880b4, 32'h4127b853} /* (4, 16, 23) {real, imag} */,
  {32'hc10630a0, 32'h40cd8e90} /* (4, 16, 22) {real, imag} */,
  {32'h412e77b8, 32'h408680c4} /* (4, 16, 21) {real, imag} */,
  {32'h408336c4, 32'hc099201e} /* (4, 16, 20) {real, imag} */,
  {32'hc0c015a6, 32'h41445a24} /* (4, 16, 19) {real, imag} */,
  {32'hc0d17064, 32'h408a4414} /* (4, 16, 18) {real, imag} */,
  {32'hc0296902, 32'h405772cd} /* (4, 16, 17) {real, imag} */,
  {32'h414b95f8, 32'hbf880160} /* (4, 16, 16) {real, imag} */,
  {32'hc0d63fa3, 32'h4042e35f} /* (4, 16, 15) {real, imag} */,
  {32'hc04d1943, 32'h40dd7bf4} /* (4, 16, 14) {real, imag} */,
  {32'h41f43630, 32'h3eb01d40} /* (4, 16, 13) {real, imag} */,
  {32'hc1114f35, 32'hc0978e6a} /* (4, 16, 12) {real, imag} */,
  {32'hc048c4e2, 32'h415feb16} /* (4, 16, 11) {real, imag} */,
  {32'hc1684eea, 32'h3ed9d108} /* (4, 16, 10) {real, imag} */,
  {32'hc11c7eb1, 32'h40c372da} /* (4, 16, 9) {real, imag} */,
  {32'hc0c5f988, 32'hc11e7454} /* (4, 16, 8) {real, imag} */,
  {32'h418ca150, 32'hc10c4ecf} /* (4, 16, 7) {real, imag} */,
  {32'h4184f2a9, 32'hc2066b95} /* (4, 16, 6) {real, imag} */,
  {32'hc1d7413b, 32'h41b462c7} /* (4, 16, 5) {real, imag} */,
  {32'h41145f97, 32'hc231f3b8} /* (4, 16, 4) {real, imag} */,
  {32'hc215d25d, 32'hc02f2c28} /* (4, 16, 3) {real, imag} */,
  {32'h409f5fda, 32'h41d08f45} /* (4, 16, 2) {real, imag} */,
  {32'h41d840dd, 32'h402b7111} /* (4, 16, 1) {real, imag} */,
  {32'h4148e448, 32'h426c5683} /* (4, 16, 0) {real, imag} */,
  {32'hc1cd36ec, 32'h41404281} /* (4, 15, 31) {real, imag} */,
  {32'hbe279900, 32'h42219a16} /* (4, 15, 30) {real, imag} */,
  {32'hc23499d8, 32'hc18cd228} /* (4, 15, 29) {real, imag} */,
  {32'hc211a4cb, 32'hc1f35d76} /* (4, 15, 28) {real, imag} */,
  {32'hbfe86f20, 32'hc097b5a6} /* (4, 15, 27) {real, imag} */,
  {32'hc0ee8574, 32'h41ffe3e1} /* (4, 15, 26) {real, imag} */,
  {32'h4215e1ce, 32'h40e53a18} /* (4, 15, 25) {real, imag} */,
  {32'h41ef7a36, 32'hc2463678} /* (4, 15, 24) {real, imag} */,
  {32'h420730b9, 32'hc18ecd84} /* (4, 15, 23) {real, imag} */,
  {32'h41d5293c, 32'hc13905d5} /* (4, 15, 22) {real, imag} */,
  {32'hc1eac92a, 32'h405864fe} /* (4, 15, 21) {real, imag} */,
  {32'h4108599e, 32'hc033a55e} /* (4, 15, 20) {real, imag} */,
  {32'hc0d8cabf, 32'h40a83e98} /* (4, 15, 19) {real, imag} */,
  {32'hbfbe5c20, 32'h40a1de45} /* (4, 15, 18) {real, imag} */,
  {32'h409a3646, 32'hc070f963} /* (4, 15, 17) {real, imag} */,
  {32'h3f695a00, 32'h40c137ee} /* (4, 15, 16) {real, imag} */,
  {32'hc0051bac, 32'h3fb68f86} /* (4, 15, 15) {real, imag} */,
  {32'h40f60c0c, 32'h3f12c578} /* (4, 15, 14) {real, imag} */,
  {32'hbebc2210, 32'hbf869b30} /* (4, 15, 13) {real, imag} */,
  {32'hc110c6c6, 32'h4136043a} /* (4, 15, 12) {real, imag} */,
  {32'hc1d3849a, 32'h4104588e} /* (4, 15, 11) {real, imag} */,
  {32'h4098faa6, 32'h40e24f9e} /* (4, 15, 10) {real, imag} */,
  {32'h40e91896, 32'hc198c08e} /* (4, 15, 9) {real, imag} */,
  {32'h409209a6, 32'hc0e2d1dc} /* (4, 15, 8) {real, imag} */,
  {32'h3e98e140, 32'hc1e7d810} /* (4, 15, 7) {real, imag} */,
  {32'h41d1a697, 32'h4093d6ec} /* (4, 15, 6) {real, imag} */,
  {32'h4234854b, 32'hc18bfc5e} /* (4, 15, 5) {real, imag} */,
  {32'h40f1cbc6, 32'h421d48af} /* (4, 15, 4) {real, imag} */,
  {32'hc206d180, 32'h41e10f8c} /* (4, 15, 3) {real, imag} */,
  {32'h41f88291, 32'h416abbf8} /* (4, 15, 2) {real, imag} */,
  {32'hc27e1c20, 32'h41b7d518} /* (4, 15, 1) {real, imag} */,
  {32'hc18e07ce, 32'hc075556c} /* (4, 15, 0) {real, imag} */,
  {32'h42aa78b1, 32'hbf0c4480} /* (4, 14, 31) {real, imag} */,
  {32'h40e4ffec, 32'h411c618c} /* (4, 14, 30) {real, imag} */,
  {32'h4029f1b6, 32'hc12e54d8} /* (4, 14, 29) {real, imag} */,
  {32'h41785d5a, 32'hc1eae925} /* (4, 14, 28) {real, imag} */,
  {32'hc16b4bb4, 32'h41b9e8f4} /* (4, 14, 27) {real, imag} */,
  {32'h41a37259, 32'h4161ef0b} /* (4, 14, 26) {real, imag} */,
  {32'h41d8d510, 32'h41cd0771} /* (4, 14, 25) {real, imag} */,
  {32'h41eed788, 32'hc1b2c833} /* (4, 14, 24) {real, imag} */,
  {32'hbfe08756, 32'h414fb89a} /* (4, 14, 23) {real, imag} */,
  {32'hbf7bdc90, 32'hc1c35459} /* (4, 14, 22) {real, imag} */,
  {32'h3ff9a24c, 32'hc142dad4} /* (4, 14, 21) {real, imag} */,
  {32'hc19edacc, 32'hc063cfec} /* (4, 14, 20) {real, imag} */,
  {32'h408e093c, 32'hc1b71026} /* (4, 14, 19) {real, imag} */,
  {32'hc032db64, 32'h4183d7be} /* (4, 14, 18) {real, imag} */,
  {32'h40c1c102, 32'h40a10d9d} /* (4, 14, 17) {real, imag} */,
  {32'hbfc024e4, 32'h410743f1} /* (4, 14, 16) {real, imag} */,
  {32'hbf556610, 32'hc0f8d043} /* (4, 14, 15) {real, imag} */,
  {32'hc0e08806, 32'h4110a293} /* (4, 14, 14) {real, imag} */,
  {32'hbfd04fb8, 32'h3ff2c760} /* (4, 14, 13) {real, imag} */,
  {32'hbf197d90, 32'h411f3b4e} /* (4, 14, 12) {real, imag} */,
  {32'h4122b004, 32'hc159f99a} /* (4, 14, 11) {real, imag} */,
  {32'h40779cfc, 32'hbea15e80} /* (4, 14, 10) {real, imag} */,
  {32'hc0ac0f5a, 32'hc1a30709} /* (4, 14, 9) {real, imag} */,
  {32'h4125bd17, 32'h41d5ce8f} /* (4, 14, 8) {real, imag} */,
  {32'hc1a0dd64, 32'hc1bea639} /* (4, 14, 7) {real, imag} */,
  {32'h414800a6, 32'h41c66292} /* (4, 14, 6) {real, imag} */,
  {32'hc18e4bce, 32'hc0242894} /* (4, 14, 5) {real, imag} */,
  {32'h422bea1e, 32'hc10219a2} /* (4, 14, 4) {real, imag} */,
  {32'hc17e4aaa, 32'h4103a61c} /* (4, 14, 3) {real, imag} */,
  {32'hc210f74a, 32'hc2852984} /* (4, 14, 2) {real, imag} */,
  {32'h42542fee, 32'h41ddf8c0} /* (4, 14, 1) {real, imag} */,
  {32'h41601858, 32'h41bc2bb8} /* (4, 14, 0) {real, imag} */,
  {32'hc1a87538, 32'h4232f62f} /* (4, 13, 31) {real, imag} */,
  {32'hc1621ad9, 32'hc258a92b} /* (4, 13, 30) {real, imag} */,
  {32'hc15c857b, 32'h420b36d0} /* (4, 13, 29) {real, imag} */,
  {32'h41a44e0c, 32'h4245e86c} /* (4, 13, 28) {real, imag} */,
  {32'h42377ed7, 32'hbfcb9860} /* (4, 13, 27) {real, imag} */,
  {32'h42366ab3, 32'h4134a2a3} /* (4, 13, 26) {real, imag} */,
  {32'hc1b83b94, 32'h420b708c} /* (4, 13, 25) {real, imag} */,
  {32'hc1b22519, 32'h410f2562} /* (4, 13, 24) {real, imag} */,
  {32'h41b56de6, 32'hc17fa6b2} /* (4, 13, 23) {real, imag} */,
  {32'hc09ff11a, 32'h409eec46} /* (4, 13, 22) {real, imag} */,
  {32'h408fa300, 32'hc0ebd20c} /* (4, 13, 21) {real, imag} */,
  {32'h41402f1f, 32'h41a59862} /* (4, 13, 20) {real, imag} */,
  {32'h41bc0950, 32'h3fa35d58} /* (4, 13, 19) {real, imag} */,
  {32'hc14eadb9, 32'hc0c8ab7c} /* (4, 13, 18) {real, imag} */,
  {32'h410b33e2, 32'hc095e072} /* (4, 13, 17) {real, imag} */,
  {32'hc09dfff0, 32'h3f696e80} /* (4, 13, 16) {real, imag} */,
  {32'hbfdbc7e0, 32'hbfa11cf8} /* (4, 13, 15) {real, imag} */,
  {32'hc10c1c3d, 32'h410e365a} /* (4, 13, 14) {real, imag} */,
  {32'hc1ab32f0, 32'hc10afdeb} /* (4, 13, 13) {real, imag} */,
  {32'hc0916d0a, 32'hc07c1d70} /* (4, 13, 12) {real, imag} */,
  {32'hc044f5e0, 32'h418f237c} /* (4, 13, 11) {real, imag} */,
  {32'h41e5a762, 32'hc186f0d0} /* (4, 13, 10) {real, imag} */,
  {32'h414c0efb, 32'h41893ce7} /* (4, 13, 9) {real, imag} */,
  {32'h4104b47a, 32'hc2761f4c} /* (4, 13, 8) {real, imag} */,
  {32'h3f906948, 32'h41c7a6cd} /* (4, 13, 7) {real, imag} */,
  {32'h41151454, 32'h4228c8a4} /* (4, 13, 6) {real, imag} */,
  {32'h3ed73680, 32'hc2253773} /* (4, 13, 5) {real, imag} */,
  {32'hc195d6e6, 32'h41e71617} /* (4, 13, 4) {real, imag} */,
  {32'hc15e242d, 32'h41b1fa38} /* (4, 13, 3) {real, imag} */,
  {32'h42053c1a, 32'h420deb67} /* (4, 13, 2) {real, imag} */,
  {32'hc1507e0f, 32'h429913a3} /* (4, 13, 1) {real, imag} */,
  {32'hc28f88db, 32'hc22572f1} /* (4, 13, 0) {real, imag} */,
  {32'hc2406b13, 32'hc284a56e} /* (4, 12, 31) {real, imag} */,
  {32'h4138b9c4, 32'h41ca5db5} /* (4, 12, 30) {real, imag} */,
  {32'h418dba75, 32'h41be85c2} /* (4, 12, 29) {real, imag} */,
  {32'h41af7860, 32'h41194121} /* (4, 12, 28) {real, imag} */,
  {32'h41d9b28d, 32'hc284b788} /* (4, 12, 27) {real, imag} */,
  {32'h4296cbba, 32'hc22f654d} /* (4, 12, 26) {real, imag} */,
  {32'h408baf7c, 32'h41eda0b8} /* (4, 12, 25) {real, imag} */,
  {32'hc178f61f, 32'h408cbf60} /* (4, 12, 24) {real, imag} */,
  {32'hc1a79967, 32'h41c4fd78} /* (4, 12, 23) {real, imag} */,
  {32'h4128bde7, 32'h4241e6a8} /* (4, 12, 22) {real, imag} */,
  {32'h3d7f0a80, 32'h41d256b2} /* (4, 12, 21) {real, imag} */,
  {32'hc1003407, 32'hc1d3e6f2} /* (4, 12, 20) {real, imag} */,
  {32'hc006a634, 32'h411f7d80} /* (4, 12, 19) {real, imag} */,
  {32'h41e5678d, 32'hc1724e03} /* (4, 12, 18) {real, imag} */,
  {32'h40705870, 32'h3fe72508} /* (4, 12, 17) {real, imag} */,
  {32'hc02076a8, 32'h403fd65c} /* (4, 12, 16) {real, imag} */,
  {32'h40d695a4, 32'h40b13f36} /* (4, 12, 15) {real, imag} */,
  {32'h401d5798, 32'h411aaf2f} /* (4, 12, 14) {real, imag} */,
  {32'hc1eaf478, 32'h40811c2c} /* (4, 12, 13) {real, imag} */,
  {32'h416405ed, 32'hc10f672d} /* (4, 12, 12) {real, imag} */,
  {32'hc150d738, 32'hc1d315ca} /* (4, 12, 11) {real, imag} */,
  {32'hc19350e2, 32'hc0fe7a2c} /* (4, 12, 10) {real, imag} */,
  {32'hc2731cc2, 32'h3f86c658} /* (4, 12, 9) {real, imag} */,
  {32'hc2101e47, 32'hc225fba8} /* (4, 12, 8) {real, imag} */,
  {32'hc20da6d2, 32'h42406320} /* (4, 12, 7) {real, imag} */,
  {32'hbe680d00, 32'h421f3c63} /* (4, 12, 6) {real, imag} */,
  {32'hc1aebde7, 32'h3f3042c0} /* (4, 12, 5) {real, imag} */,
  {32'h421b8e9e, 32'h41ce89d4} /* (4, 12, 4) {real, imag} */,
  {32'hc1d23143, 32'hc1cf7982} /* (4, 12, 3) {real, imag} */,
  {32'h42098d7f, 32'hc268ec54} /* (4, 12, 2) {real, imag} */,
  {32'hc131b634, 32'hc1540cb4} /* (4, 12, 1) {real, imag} */,
  {32'hc206e686, 32'hc1a8e6b4} /* (4, 12, 0) {real, imag} */,
  {32'h4283bb7c, 32'hc1d5b101} /* (4, 11, 31) {real, imag} */,
  {32'hc2d435e9, 32'hc216f782} /* (4, 11, 30) {real, imag} */,
  {32'hc2009342, 32'h421c7290} /* (4, 11, 29) {real, imag} */,
  {32'h42238715, 32'hc09eef0e} /* (4, 11, 28) {real, imag} */,
  {32'h408e0db0, 32'hc1ad1626} /* (4, 11, 27) {real, imag} */,
  {32'h4232c6ce, 32'hc1a1320d} /* (4, 11, 26) {real, imag} */,
  {32'hc0c2ee5e, 32'hc2142022} /* (4, 11, 25) {real, imag} */,
  {32'h40f1fdaa, 32'h4238bd51} /* (4, 11, 24) {real, imag} */,
  {32'hc2008a9a, 32'h41921163} /* (4, 11, 23) {real, imag} */,
  {32'h422d1540, 32'hc128e39e} /* (4, 11, 22) {real, imag} */,
  {32'hc1b22704, 32'hc1064e55} /* (4, 11, 21) {real, imag} */,
  {32'hc1faf00c, 32'h423236ba} /* (4, 11, 20) {real, imag} */,
  {32'hc2007186, 32'hc19582de} /* (4, 11, 19) {real, imag} */,
  {32'h410e5edc, 32'h4162f55e} /* (4, 11, 18) {real, imag} */,
  {32'hc164df12, 32'hc0dd0df3} /* (4, 11, 17) {real, imag} */,
  {32'h412e8200, 32'hc13e5bbb} /* (4, 11, 16) {real, imag} */,
  {32'h40c08274, 32'h41a9633f} /* (4, 11, 15) {real, imag} */,
  {32'hc1a0b5a8, 32'hc154300e} /* (4, 11, 14) {real, imag} */,
  {32'hc1c817af, 32'h40cb48b2} /* (4, 11, 13) {real, imag} */,
  {32'h3e7e5840, 32'h3eb09ec0} /* (4, 11, 12) {real, imag} */,
  {32'h418fa62a, 32'hc09906da} /* (4, 11, 11) {real, imag} */,
  {32'hc11d3c06, 32'h4243c104} /* (4, 11, 10) {real, imag} */,
  {32'hc19f2d31, 32'h41ae3dff} /* (4, 11, 9) {real, imag} */,
  {32'hc1d42712, 32'h4185c662} /* (4, 11, 8) {real, imag} */,
  {32'hc1907aec, 32'hc15a62de} /* (4, 11, 7) {real, imag} */,
  {32'hc16f6492, 32'hc231f25c} /* (4, 11, 6) {real, imag} */,
  {32'hc2c7d1a3, 32'hc20dba6b} /* (4, 11, 5) {real, imag} */,
  {32'hc02c2870, 32'h41873b06} /* (4, 11, 4) {real, imag} */,
  {32'h42bab4df, 32'h4122b6f5} /* (4, 11, 3) {real, imag} */,
  {32'h4186f4e4, 32'hc2e556c3} /* (4, 11, 2) {real, imag} */,
  {32'h431e31ae, 32'hc1349cb6} /* (4, 11, 1) {real, imag} */,
  {32'h42379e16, 32'hc1a870ba} /* (4, 11, 0) {real, imag} */,
  {32'hc257de16, 32'hc2619c18} /* (4, 10, 31) {real, imag} */,
  {32'h4235c455, 32'h42eb84b0} /* (4, 10, 30) {real, imag} */,
  {32'h42779b88, 32'hc194ba08} /* (4, 10, 29) {real, imag} */,
  {32'hc15dbf3a, 32'h40a11f88} /* (4, 10, 28) {real, imag} */,
  {32'hc1dd4042, 32'h41a3569a} /* (4, 10, 27) {real, imag} */,
  {32'hc29661a0, 32'h427a6443} /* (4, 10, 26) {real, imag} */,
  {32'hc21f5925, 32'h4241eda9} /* (4, 10, 25) {real, imag} */,
  {32'h4164b454, 32'hc0046b90} /* (4, 10, 24) {real, imag} */,
  {32'h41d55c9e, 32'hc2cab916} /* (4, 10, 23) {real, imag} */,
  {32'hc0cc7a06, 32'hc04d5cbc} /* (4, 10, 22) {real, imag} */,
  {32'h421159a1, 32'hc1a8d722} /* (4, 10, 21) {real, imag} */,
  {32'h4152bfcc, 32'h41c87cbc} /* (4, 10, 20) {real, imag} */,
  {32'h4082d8d6, 32'h411d0b9e} /* (4, 10, 19) {real, imag} */,
  {32'hc0240bf0, 32'h414af578} /* (4, 10, 18) {real, imag} */,
  {32'h40d5e2e4, 32'h3edb1dc0} /* (4, 10, 17) {real, imag} */,
  {32'hc1084450, 32'hc151a6e0} /* (4, 10, 16) {real, imag} */,
  {32'hc1fd8eb5, 32'h402159e8} /* (4, 10, 15) {real, imag} */,
  {32'hc1203884, 32'hc1a4c168} /* (4, 10, 14) {real, imag} */,
  {32'hc00e278c, 32'h4169e5c4} /* (4, 10, 13) {real, imag} */,
  {32'hc1e550de, 32'h419c9728} /* (4, 10, 12) {real, imag} */,
  {32'hc1a4a1d6, 32'h40ebfbc6} /* (4, 10, 11) {real, imag} */,
  {32'hc1937b72, 32'hbf49ab10} /* (4, 10, 10) {real, imag} */,
  {32'h429f1636, 32'hc229b038} /* (4, 10, 9) {real, imag} */,
  {32'h4275dfd7, 32'hc27cae09} /* (4, 10, 8) {real, imag} */,
  {32'hc23658bb, 32'hc110c934} /* (4, 10, 7) {real, imag} */,
  {32'hc21e2d45, 32'h424bcc55} /* (4, 10, 6) {real, imag} */,
  {32'h421c5fcb, 32'h4219da17} /* (4, 10, 5) {real, imag} */,
  {32'h42285058, 32'hc281e748} /* (4, 10, 4) {real, imag} */,
  {32'h42917ebc, 32'hc23a0ff0} /* (4, 10, 3) {real, imag} */,
  {32'h43025771, 32'h4108a3d8} /* (4, 10, 2) {real, imag} */,
  {32'h410d952a, 32'h409b664c} /* (4, 10, 1) {real, imag} */,
  {32'hc2b398d0, 32'hc09a872c} /* (4, 10, 0) {real, imag} */,
  {32'h4200df26, 32'hc28a5565} /* (4, 9, 31) {real, imag} */,
  {32'h428158d7, 32'h428cd807} /* (4, 9, 30) {real, imag} */,
  {32'h41363098, 32'hc2270eb4} /* (4, 9, 29) {real, imag} */,
  {32'hc328a928, 32'h42a36873} /* (4, 9, 28) {real, imag} */,
  {32'h424cee6b, 32'hc22be578} /* (4, 9, 27) {real, imag} */,
  {32'hc1874724, 32'hc0e8df40} /* (4, 9, 26) {real, imag} */,
  {32'h422ee460, 32'hc2163e2b} /* (4, 9, 25) {real, imag} */,
  {32'h424ae03d, 32'hc17ac66c} /* (4, 9, 24) {real, imag} */,
  {32'h4214d184, 32'h3fe4e540} /* (4, 9, 23) {real, imag} */,
  {32'hc12bfd8e, 32'h41d120ab} /* (4, 9, 22) {real, imag} */,
  {32'h425e337a, 32'h40e392a4} /* (4, 9, 21) {real, imag} */,
  {32'hbf862a60, 32'h40c151c2} /* (4, 9, 20) {real, imag} */,
  {32'hc10aa946, 32'hc1043679} /* (4, 9, 19) {real, imag} */,
  {32'hc08c4532, 32'hc123d5dd} /* (4, 9, 18) {real, imag} */,
  {32'h40ee16ec, 32'hc18d4094} /* (4, 9, 17) {real, imag} */,
  {32'h41712584, 32'hc10cb538} /* (4, 9, 16) {real, imag} */,
  {32'h4182397f, 32'h4047fc24} /* (4, 9, 15) {real, imag} */,
  {32'hc146c3a7, 32'hc150492d} /* (4, 9, 14) {real, imag} */,
  {32'h419eea4b, 32'h415c881f} /* (4, 9, 13) {real, imag} */,
  {32'h415125bc, 32'h420f3090} /* (4, 9, 12) {real, imag} */,
  {32'h410780ae, 32'h417e4332} /* (4, 9, 11) {real, imag} */,
  {32'h422cc62a, 32'h418c1ebd} /* (4, 9, 10) {real, imag} */,
  {32'hc1ae5a1a, 32'h41f2c6e0} /* (4, 9, 9) {real, imag} */,
  {32'hc2a8d5c2, 32'h427a09af} /* (4, 9, 8) {real, imag} */,
  {32'hc0c58ee8, 32'h42985ea8} /* (4, 9, 7) {real, imag} */,
  {32'h430d5354, 32'hc2cbda98} /* (4, 9, 6) {real, imag} */,
  {32'hc19a46c2, 32'h41b28daf} /* (4, 9, 5) {real, imag} */,
  {32'hc209b9d6, 32'h4266601e} /* (4, 9, 4) {real, imag} */,
  {32'hc2e669b5, 32'h424ed022} /* (4, 9, 3) {real, imag} */,
  {32'h42760ab6, 32'hc20d5d08} /* (4, 9, 2) {real, imag} */,
  {32'hc32aab20, 32'hc20034d4} /* (4, 9, 1) {real, imag} */,
  {32'hc241c04d, 32'hc2625f0a} /* (4, 9, 0) {real, imag} */,
  {32'h43589cf6, 32'hc34ac724} /* (4, 8, 31) {real, imag} */,
  {32'hc2b44780, 32'h43001234} /* (4, 8, 30) {real, imag} */,
  {32'hc2e5a048, 32'h432e30d6} /* (4, 8, 29) {real, imag} */,
  {32'h42e1ab45, 32'hc2866790} /* (4, 8, 28) {real, imag} */,
  {32'h42a905fb, 32'h42f9fe90} /* (4, 8, 27) {real, imag} */,
  {32'h41038688, 32'h42706a4a} /* (4, 8, 26) {real, imag} */,
  {32'h428e2e12, 32'hc292bc18} /* (4, 8, 25) {real, imag} */,
  {32'h423d2c6c, 32'h40b22b48} /* (4, 8, 24) {real, imag} */,
  {32'h426429c5, 32'h423b7c14} /* (4, 8, 23) {real, imag} */,
  {32'h41be5ffc, 32'hc1d30b35} /* (4, 8, 22) {real, imag} */,
  {32'hc250756e, 32'h42658679} /* (4, 8, 21) {real, imag} */,
  {32'hc01c9d38, 32'h41f1ced6} /* (4, 8, 20) {real, imag} */,
  {32'hc1cf8500, 32'h41500814} /* (4, 8, 19) {real, imag} */,
  {32'hc16ad8ec, 32'hbf37ad90} /* (4, 8, 18) {real, imag} */,
  {32'hbf518b40, 32'h4001a570} /* (4, 8, 17) {real, imag} */,
  {32'hc080fddc, 32'hc1edf01a} /* (4, 8, 16) {real, imag} */,
  {32'h41f5275a, 32'hc0602830} /* (4, 8, 15) {real, imag} */,
  {32'h4222344d, 32'hc15dcd87} /* (4, 8, 14) {real, imag} */,
  {32'hc2030436, 32'h4143c17c} /* (4, 8, 13) {real, imag} */,
  {32'hc2020bec, 32'hc274b0d3} /* (4, 8, 12) {real, imag} */,
  {32'hc1a06aec, 32'h419a8202} /* (4, 8, 11) {real, imag} */,
  {32'hc207adaf, 32'h4119c556} /* (4, 8, 10) {real, imag} */,
  {32'h420f5203, 32'hc127e3f8} /* (4, 8, 9) {real, imag} */,
  {32'hc1536f94, 32'hc006c0d0} /* (4, 8, 8) {real, imag} */,
  {32'h42c36c0a, 32'h42a5fd58} /* (4, 8, 7) {real, imag} */,
  {32'hc2bbaa15, 32'hc20b434a} /* (4, 8, 6) {real, imag} */,
  {32'hc26e5782, 32'hc32d9a5a} /* (4, 8, 5) {real, imag} */,
  {32'h42f70dbb, 32'h4224669f} /* (4, 8, 4) {real, imag} */,
  {32'hc1bf5f6e, 32'h41d97164} /* (4, 8, 3) {real, imag} */,
  {32'hc2dd296c, 32'h431fc012} /* (4, 8, 2) {real, imag} */,
  {32'h439af01f, 32'hc2cf3f30} /* (4, 8, 1) {real, imag} */,
  {32'h4261f0f6, 32'hc1eaf0ce} /* (4, 8, 0) {real, imag} */,
  {32'h41f39528, 32'h430a9b04} /* (4, 7, 31) {real, imag} */,
  {32'h42782954, 32'hc2daf5ce} /* (4, 7, 30) {real, imag} */,
  {32'hc281e9be, 32'h4296d199} /* (4, 7, 29) {real, imag} */,
  {32'h4260141d, 32'h42a1dd69} /* (4, 7, 28) {real, imag} */,
  {32'hc1940c3e, 32'hc329599b} /* (4, 7, 27) {real, imag} */,
  {32'hc2939b44, 32'hc20f8e54} /* (4, 7, 26) {real, imag} */,
  {32'hc26da894, 32'hc287fc2a} /* (4, 7, 25) {real, imag} */,
  {32'hc1233be8, 32'hc1c59b88} /* (4, 7, 24) {real, imag} */,
  {32'h42acb57e, 32'h42599f78} /* (4, 7, 23) {real, imag} */,
  {32'hc127a66c, 32'hc0e0a1b0} /* (4, 7, 22) {real, imag} */,
  {32'hc1006864, 32'hc0e42a24} /* (4, 7, 21) {real, imag} */,
  {32'h4215b438, 32'h4217359f} /* (4, 7, 20) {real, imag} */,
  {32'hc0e688c8, 32'hc26bd32e} /* (4, 7, 19) {real, imag} */,
  {32'hc1aa7d3f, 32'h3f3e0100} /* (4, 7, 18) {real, imag} */,
  {32'h41c126fc, 32'hc166606a} /* (4, 7, 17) {real, imag} */,
  {32'h420a683f, 32'hc19dc170} /* (4, 7, 16) {real, imag} */,
  {32'hc197ca50, 32'hc1962801} /* (4, 7, 15) {real, imag} */,
  {32'h420d2124, 32'h41cdf778} /* (4, 7, 14) {real, imag} */,
  {32'h41d1828e, 32'hbf4c77e0} /* (4, 7, 13) {real, imag} */,
  {32'hc162c673, 32'hc19f06b6} /* (4, 7, 12) {real, imag} */,
  {32'h422a2a2a, 32'hc22fd104} /* (4, 7, 11) {real, imag} */,
  {32'hc29db9b0, 32'h42732022} /* (4, 7, 10) {real, imag} */,
  {32'h41f2e272, 32'hc13dfefe} /* (4, 7, 9) {real, imag} */,
  {32'hc0137cc0, 32'h423766b0} /* (4, 7, 8) {real, imag} */,
  {32'h4305089d, 32'hc2621c4c} /* (4, 7, 7) {real, imag} */,
  {32'hc30e4d3c, 32'h428562d6} /* (4, 7, 6) {real, imag} */,
  {32'hc2245b4e, 32'h43081135} /* (4, 7, 5) {real, imag} */,
  {32'hc1757094, 32'hc28a2517} /* (4, 7, 4) {real, imag} */,
  {32'hc297e01a, 32'hc247858e} /* (4, 7, 3) {real, imag} */,
  {32'h4316ec3e, 32'h41025e60} /* (4, 7, 2) {real, imag} */,
  {32'hc36aa675, 32'hc1be47cc} /* (4, 7, 1) {real, imag} */,
  {32'hc29a4abe, 32'h42b7b3c5} /* (4, 7, 0) {real, imag} */,
  {32'hc2d55c7b, 32'h400a9750} /* (4, 6, 31) {real, imag} */,
  {32'hc31e71ee, 32'h42b8b38b} /* (4, 6, 30) {real, imag} */,
  {32'hc16f7136, 32'hc26558a7} /* (4, 6, 29) {real, imag} */,
  {32'hc27eb666, 32'h42a4f044} /* (4, 6, 28) {real, imag} */,
  {32'hc2a0cc4a, 32'hc190c484} /* (4, 6, 27) {real, imag} */,
  {32'hc2577456, 32'h4229c3a2} /* (4, 6, 26) {real, imag} */,
  {32'hc0fa15a4, 32'h4294c585} /* (4, 6, 25) {real, imag} */,
  {32'h42c1b707, 32'hc1f8391a} /* (4, 6, 24) {real, imag} */,
  {32'h428f11fe, 32'hc17275e6} /* (4, 6, 23) {real, imag} */,
  {32'hc1fdeb46, 32'hc2cba27a} /* (4, 6, 22) {real, imag} */,
  {32'h424be4e2, 32'hc20c0734} /* (4, 6, 21) {real, imag} */,
  {32'h40381078, 32'hc2b81b75} /* (4, 6, 20) {real, imag} */,
  {32'h4197c325, 32'hc1ecbc2e} /* (4, 6, 19) {real, imag} */,
  {32'h413d102c, 32'h40806566} /* (4, 6, 18) {real, imag} */,
  {32'h41b2d392, 32'h40e59752} /* (4, 6, 17) {real, imag} */,
  {32'h411f34d2, 32'h3ef64100} /* (4, 6, 16) {real, imag} */,
  {32'h3e9f1700, 32'h418e8912} /* (4, 6, 15) {real, imag} */,
  {32'hc1b657f6, 32'h41890cb6} /* (4, 6, 14) {real, imag} */,
  {32'hc137a7be, 32'hc1fa011e} /* (4, 6, 13) {real, imag} */,
  {32'hc1ec4be3, 32'h421be1aa} /* (4, 6, 12) {real, imag} */,
  {32'hc24a516c, 32'hc1925cee} /* (4, 6, 11) {real, imag} */,
  {32'hc1618134, 32'h423f84bf} /* (4, 6, 10) {real, imag} */,
  {32'h42781e54, 32'hc2129546} /* (4, 6, 9) {real, imag} */,
  {32'h41fbd9c4, 32'h42470b49} /* (4, 6, 8) {real, imag} */,
  {32'hbfd1d7d0, 32'hc231bc1a} /* (4, 6, 7) {real, imag} */,
  {32'hc0adf3e0, 32'hc2d7f3ed} /* (4, 6, 6) {real, imag} */,
  {32'h42477ec8, 32'h421f8df9} /* (4, 6, 5) {real, imag} */,
  {32'h423e2fba, 32'hc15b5630} /* (4, 6, 4) {real, imag} */,
  {32'h411bd762, 32'h422cf3f3} /* (4, 6, 3) {real, imag} */,
  {32'hc2adf448, 32'hc2f36825} /* (4, 6, 2) {real, imag} */,
  {32'hc1d52714, 32'hc2944c32} /* (4, 6, 1) {real, imag} */,
  {32'hc25f8326, 32'hc2f3a05f} /* (4, 6, 0) {real, imag} */,
  {32'h425783fc, 32'hc336db67} /* (4, 5, 31) {real, imag} */,
  {32'hc133e8fc, 32'h427b6a22} /* (4, 5, 30) {real, imag} */,
  {32'h426f58ec, 32'hc186933a} /* (4, 5, 29) {real, imag} */,
  {32'h4319bfa6, 32'hc280b2c4} /* (4, 5, 28) {real, imag} */,
  {32'hc25b46a0, 32'h43001300} /* (4, 5, 27) {real, imag} */,
  {32'hc15eb798, 32'hc06fb080} /* (4, 5, 26) {real, imag} */,
  {32'hc2d18537, 32'hc2f23c86} /* (4, 5, 25) {real, imag} */,
  {32'hc1cf3ff0, 32'hc247541b} /* (4, 5, 24) {real, imag} */,
  {32'h422b8d42, 32'hc1d0d9ae} /* (4, 5, 23) {real, imag} */,
  {32'hc167a3e7, 32'hc17a58b0} /* (4, 5, 22) {real, imag} */,
  {32'hc1cdb396, 32'h424dd29e} /* (4, 5, 21) {real, imag} */,
  {32'h400446b8, 32'hc24f8c76} /* (4, 5, 20) {real, imag} */,
  {32'h42a84158, 32'hc1854ff6} /* (4, 5, 19) {real, imag} */,
  {32'h418da94a, 32'h41cba59b} /* (4, 5, 18) {real, imag} */,
  {32'hc1561608, 32'h3eb9acc0} /* (4, 5, 17) {real, imag} */,
  {32'h419ed534, 32'hc10bb9b8} /* (4, 5, 16) {real, imag} */,
  {32'h4109b428, 32'hc08ed78c} /* (4, 5, 15) {real, imag} */,
  {32'h41290abc, 32'hc0d3fcec} /* (4, 5, 14) {real, imag} */,
  {32'h4215e6c7, 32'hc0b1aa4a} /* (4, 5, 13) {real, imag} */,
  {32'h40c8a97c, 32'h409d3a18} /* (4, 5, 12) {real, imag} */,
  {32'hc20deb09, 32'h413c62d2} /* (4, 5, 11) {real, imag} */,
  {32'h412e98e9, 32'hc2d17d84} /* (4, 5, 10) {real, imag} */,
  {32'hc28f2edc, 32'hc0ecf378} /* (4, 5, 9) {real, imag} */,
  {32'h4189fe78, 32'hc29ccfb2} /* (4, 5, 8) {real, imag} */,
  {32'h4218aeea, 32'hc1049670} /* (4, 5, 7) {real, imag} */,
  {32'hc227c962, 32'h434f2845} /* (4, 5, 6) {real, imag} */,
  {32'h3f33a880, 32'h419b8ee6} /* (4, 5, 5) {real, imag} */,
  {32'hc29623ad, 32'h420d019c} /* (4, 5, 4) {real, imag} */,
  {32'hc2bc84de, 32'h41a7aad2} /* (4, 5, 3) {real, imag} */,
  {32'hc2db163e, 32'h42cf12ff} /* (4, 5, 2) {real, imag} */,
  {32'h438ab83c, 32'hc2fc39d6} /* (4, 5, 1) {real, imag} */,
  {32'h431c8412, 32'hc308ac3a} /* (4, 5, 0) {real, imag} */,
  {32'hc399286f, 32'h43598428} /* (4, 4, 31) {real, imag} */,
  {32'h4385594a, 32'h42703c55} /* (4, 4, 30) {real, imag} */,
  {32'hc29059ab, 32'hc2e1e375} /* (4, 4, 29) {real, imag} */,
  {32'hc3971dfc, 32'h432bed84} /* (4, 4, 28) {real, imag} */,
  {32'hc0d48644, 32'hc3020d26} /* (4, 4, 27) {real, imag} */,
  {32'h428959f0, 32'h4294aaaa} /* (4, 4, 26) {real, imag} */,
  {32'hc2d7fd16, 32'hc08284b8} /* (4, 4, 25) {real, imag} */,
  {32'hc1c737c0, 32'hc1eda3b6} /* (4, 4, 24) {real, imag} */,
  {32'h42bd93b8, 32'hc236749e} /* (4, 4, 23) {real, imag} */,
  {32'hc1e8ff88, 32'h41e2df88} /* (4, 4, 22) {real, imag} */,
  {32'h421955d6, 32'hc243cc94} /* (4, 4, 21) {real, imag} */,
  {32'h3d0ea800, 32'h41978172} /* (4, 4, 20) {real, imag} */,
  {32'hc2048fbe, 32'h4276738b} /* (4, 4, 19) {real, imag} */,
  {32'hc12498e8, 32'h416fbd1c} /* (4, 4, 18) {real, imag} */,
  {32'hc1c74447, 32'hc0e89c90} /* (4, 4, 17) {real, imag} */,
  {32'h41279da8, 32'hc139a79c} /* (4, 4, 16) {real, imag} */,
  {32'h41489a6e, 32'hbf384580} /* (4, 4, 15) {real, imag} */,
  {32'h41854db4, 32'hc1a27f84} /* (4, 4, 14) {real, imag} */,
  {32'h429c8fd1, 32'h41a127b6} /* (4, 4, 13) {real, imag} */,
  {32'hc147e068, 32'hc12f92e4} /* (4, 4, 12) {real, imag} */,
  {32'h42359af6, 32'h417a0752} /* (4, 4, 11) {real, imag} */,
  {32'h419d79c4, 32'hc223ae70} /* (4, 4, 10) {real, imag} */,
  {32'h42a8b910, 32'h429d0343} /* (4, 4, 9) {real, imag} */,
  {32'h427a8e60, 32'hc04e67f0} /* (4, 4, 8) {real, imag} */,
  {32'hc2a9a5e2, 32'h41e9115c} /* (4, 4, 7) {real, imag} */,
  {32'h42a9e92c, 32'hc2c4f558} /* (4, 4, 6) {real, imag} */,
  {32'h4044aea8, 32'hc196d934} /* (4, 4, 5) {real, imag} */,
  {32'hc2d345e9, 32'hc1ec51c4} /* (4, 4, 4) {real, imag} */,
  {32'hc26352aa, 32'h42d0f913} /* (4, 4, 3) {real, imag} */,
  {32'h439e3b3e, 32'hc2ac0b71} /* (4, 4, 2) {real, imag} */,
  {32'hc39f7cc5, 32'h43f6cfa4} /* (4, 4, 1) {real, imag} */,
  {32'hc306c1a6, 32'h428ad316} /* (4, 4, 0) {real, imag} */,
  {32'h41ec92b0, 32'hc3a0893f} /* (4, 3, 31) {real, imag} */,
  {32'h437fe440, 32'h433d60c8} /* (4, 3, 30) {real, imag} */,
  {32'h42167406, 32'h42cf41fe} /* (4, 3, 29) {real, imag} */,
  {32'hc280f7d0, 32'hc295e026} /* (4, 3, 28) {real, imag} */,
  {32'h4287aa9a, 32'h42da851c} /* (4, 3, 27) {real, imag} */,
  {32'h3fb42200, 32'hc21a6814} /* (4, 3, 26) {real, imag} */,
  {32'h42564e04, 32'hc2657b43} /* (4, 3, 25) {real, imag} */,
  {32'h41ac8d74, 32'h422ec4f6} /* (4, 3, 24) {real, imag} */,
  {32'hc2ef3c6c, 32'h40e227d0} /* (4, 3, 23) {real, imag} */,
  {32'hc1dd359e, 32'h42631d4e} /* (4, 3, 22) {real, imag} */,
  {32'h42122ca4, 32'hc2affebe} /* (4, 3, 21) {real, imag} */,
  {32'hc2ad3ee4, 32'h4243f376} /* (4, 3, 20) {real, imag} */,
  {32'h4234c688, 32'h41a5a17b} /* (4, 3, 19) {real, imag} */,
  {32'h41fa612f, 32'h42073940} /* (4, 3, 18) {real, imag} */,
  {32'hc21474e9, 32'hc2798708} /* (4, 3, 17) {real, imag} */,
  {32'hc0dc4390, 32'h4249baad} /* (4, 3, 16) {real, imag} */,
  {32'hc113e884, 32'h40f01be0} /* (4, 3, 15) {real, imag} */,
  {32'hc149de1e, 32'h42043e8c} /* (4, 3, 14) {real, imag} */,
  {32'hc263e17a, 32'h4166ba3a} /* (4, 3, 13) {real, imag} */,
  {32'h400e5930, 32'hc26928f6} /* (4, 3, 12) {real, imag} */,
  {32'h40478b68, 32'h4228211f} /* (4, 3, 11) {real, imag} */,
  {32'hc1c21d7e, 32'hc2a6689b} /* (4, 3, 10) {real, imag} */,
  {32'h424013b4, 32'hc2621aec} /* (4, 3, 9) {real, imag} */,
  {32'h40e33f68, 32'hc0fd9b1c} /* (4, 3, 8) {real, imag} */,
  {32'hc318712c, 32'h43105535} /* (4, 3, 7) {real, imag} */,
  {32'h41f1c324, 32'h43117148} /* (4, 3, 6) {real, imag} */,
  {32'h422d7c0f, 32'h42ba5224} /* (4, 3, 5) {real, imag} */,
  {32'h426def32, 32'hc13ddf32} /* (4, 3, 4) {real, imag} */,
  {32'hc30ff4fc, 32'h4090f940} /* (4, 3, 3) {real, imag} */,
  {32'h43260ce4, 32'hc1b18c98} /* (4, 3, 2) {real, imag} */,
  {32'hc384a7bc, 32'hc1c1d010} /* (4, 3, 1) {real, imag} */,
  {32'h41ef2aaa, 32'hc193afc6} /* (4, 3, 0) {real, imag} */,
  {32'h43f08c8a, 32'hc48965da} /* (4, 2, 31) {real, imag} */,
  {32'hc33ec105, 32'h44495bc2} /* (4, 2, 30) {real, imag} */,
  {32'h42821580, 32'hc32da934} /* (4, 2, 29) {real, imag} */,
  {32'hc2b91d45, 32'hc38a876f} /* (4, 2, 28) {real, imag} */,
  {32'h42986463, 32'h434622dc} /* (4, 2, 27) {real, imag} */,
  {32'hc28ab4f8, 32'hc2918d04} /* (4, 2, 26) {real, imag} */,
  {32'h41a5f234, 32'hc26c1119} /* (4, 2, 25) {real, imag} */,
  {32'h423ef19b, 32'h435ab78a} /* (4, 2, 24) {real, imag} */,
  {32'h426dfbaa, 32'h41e0ed6a} /* (4, 2, 23) {real, imag} */,
  {32'hc2eb4c5e, 32'h419deb00} /* (4, 2, 22) {real, imag} */,
  {32'h42b59bdb, 32'h428f6174} /* (4, 2, 21) {real, imag} */,
  {32'hc2125cf0, 32'hc1d237ea} /* (4, 2, 20) {real, imag} */,
  {32'h408f6f9c, 32'h40eded76} /* (4, 2, 19) {real, imag} */,
  {32'h4170319c, 32'hc0c3af98} /* (4, 2, 18) {real, imag} */,
  {32'hc0f61ca0, 32'hbc22a000} /* (4, 2, 17) {real, imag} */,
  {32'hc223f8d4, 32'h41e3caa0} /* (4, 2, 16) {real, imag} */,
  {32'hc1bcb0d8, 32'hc1c08c0c} /* (4, 2, 15) {real, imag} */,
  {32'hc22e2507, 32'h428269a2} /* (4, 2, 14) {real, imag} */,
  {32'h41181756, 32'hc1b076fe} /* (4, 2, 13) {real, imag} */,
  {32'h40b3865c, 32'hc24f6d0b} /* (4, 2, 12) {real, imag} */,
  {32'hc28c1c13, 32'h40abad80} /* (4, 2, 11) {real, imag} */,
  {32'h3f6bdf80, 32'hc2666b70} /* (4, 2, 10) {real, imag} */,
  {32'hc2a4985f, 32'h41c35f9a} /* (4, 2, 9) {real, imag} */,
  {32'hc2b9f1ce, 32'h432b0f20} /* (4, 2, 8) {real, imag} */,
  {32'h42b66e31, 32'hc183c5d2} /* (4, 2, 7) {real, imag} */,
  {32'hc28f3f24, 32'hc1e6b50e} /* (4, 2, 6) {real, imag} */,
  {32'hc333c5dc, 32'h43402cb6} /* (4, 2, 5) {real, imag} */,
  {32'hc2202d16, 32'hc347adf6} /* (4, 2, 4) {real, imag} */,
  {32'h426704e9, 32'hc2ee9807} /* (4, 2, 3) {real, imag} */,
  {32'hc0d94ba0, 32'h440b0116} /* (4, 2, 2) {real, imag} */,
  {32'h42ded3d6, 32'hc4219004} /* (4, 2, 1) {real, imag} */,
  {32'h439cd4c0, 32'hc40c71b3} /* (4, 2, 0) {real, imag} */,
  {32'hc21772e0, 32'h4458d853} /* (4, 1, 31) {real, imag} */,
  {32'h432f9d72, 32'hc3cf50f3} /* (4, 1, 30) {real, imag} */,
  {32'hc171be28, 32'h4302885f} /* (4, 1, 29) {real, imag} */,
  {32'hc260ad09, 32'h437f9fd8} /* (4, 1, 28) {real, imag} */,
  {32'h4331077c, 32'hc3e08325} /* (4, 1, 27) {real, imag} */,
  {32'hc2dbaf48, 32'h42a3e556} /* (4, 1, 26) {real, imag} */,
  {32'h4300b8bc, 32'h41b01ae5} /* (4, 1, 25) {real, imag} */,
  {32'hc2b01946, 32'hc33bfc2a} /* (4, 1, 24) {real, imag} */,
  {32'h4105c998, 32'h41541c58} /* (4, 1, 23) {real, imag} */,
  {32'h41686ba0, 32'h4236185d} /* (4, 1, 22) {real, imag} */,
  {32'hc364b8de, 32'hc3129b63} /* (4, 1, 21) {real, imag} */,
  {32'h42e1514a, 32'h4203cac8} /* (4, 1, 20) {real, imag} */,
  {32'hc21824d6, 32'h4173f114} /* (4, 1, 19) {real, imag} */,
  {32'hc2a6409a, 32'h40c98150} /* (4, 1, 18) {real, imag} */,
  {32'hc18d8c20, 32'hc10868f8} /* (4, 1, 17) {real, imag} */,
  {32'h424af840, 32'h41b6bf80} /* (4, 1, 16) {real, imag} */,
  {32'hc22ec200, 32'hc21d2702} /* (4, 1, 15) {real, imag} */,
  {32'h40ac85e0, 32'h4208e3d6} /* (4, 1, 14) {real, imag} */,
  {32'hc1981388, 32'hc154f7dc} /* (4, 1, 13) {real, imag} */,
  {32'hbf9bd7e0, 32'hc27854dc} /* (4, 1, 12) {real, imag} */,
  {32'h42897bf3, 32'hc1a34d00} /* (4, 1, 11) {real, imag} */,
  {32'hc23af6c4, 32'hc268f83d} /* (4, 1, 10) {real, imag} */,
  {32'h428076e7, 32'h42a40421} /* (4, 1, 9) {real, imag} */,
  {32'h433c3915, 32'hc10f8560} /* (4, 1, 8) {real, imag} */,
  {32'hc1c76b14, 32'hc0e401d4} /* (4, 1, 7) {real, imag} */,
  {32'h42f6f576, 32'h429b6962} /* (4, 1, 6) {real, imag} */,
  {32'h4380b248, 32'hc3208d62} /* (4, 1, 5) {real, imag} */,
  {32'hc221809b, 32'hc16d77c8} /* (4, 1, 4) {real, imag} */,
  {32'hc213a924, 32'hc32c0029} /* (4, 1, 3) {real, imag} */,
  {32'h445fd3a6, 32'hc368218a} /* (4, 1, 2) {real, imag} */,
  {32'hc48513ed, 32'h4451fb6d} /* (4, 1, 1) {real, imag} */,
  {32'hc4187fe4, 32'h44335fe0} /* (4, 1, 0) {real, imag} */,
  {32'h436f90fe, 32'h4440bafc} /* (4, 0, 31) {real, imag} */,
  {32'hc364ea90, 32'hc236a84a} /* (4, 0, 30) {real, imag} */,
  {32'h41984c66, 32'h42bcfcfa} /* (4, 0, 29) {real, imag} */,
  {32'hc274b3bf, 32'hc2cde885} /* (4, 0, 28) {real, imag} */,
  {32'h4326fd99, 32'hc33667ff} /* (4, 0, 27) {real, imag} */,
  {32'h42ab15ba, 32'h3f8befe0} /* (4, 0, 26) {real, imag} */,
  {32'h430e97b6, 32'h42ab2bc3} /* (4, 0, 25) {real, imag} */,
  {32'hc247e0dc, 32'hc2a2d840} /* (4, 0, 24) {real, imag} */,
  {32'hc300b2a8, 32'hc3253aa0} /* (4, 0, 23) {real, imag} */,
  {32'h42a47e98, 32'hc1c650e6} /* (4, 0, 22) {real, imag} */,
  {32'h4155b9cc, 32'hc2f4933e} /* (4, 0, 21) {real, imag} */,
  {32'h41a397ed, 32'hc096216b} /* (4, 0, 20) {real, imag} */,
  {32'hc0e360a8, 32'h4091b990} /* (4, 0, 19) {real, imag} */,
  {32'hc2c221a6, 32'hc1d5fd12} /* (4, 0, 18) {real, imag} */,
  {32'hc21c7caa, 32'h4183608c} /* (4, 0, 17) {real, imag} */,
  {32'h420191b2, 32'hc14d3fd0} /* (4, 0, 16) {real, imag} */,
  {32'h41aa29bc, 32'hc137d618} /* (4, 0, 15) {real, imag} */,
  {32'h421b0ebc, 32'hc127d330} /* (4, 0, 14) {real, imag} */,
  {32'hc0f1b178, 32'hc28c06a6} /* (4, 0, 13) {real, imag} */,
  {32'hc08333dc, 32'hc1316e76} /* (4, 0, 12) {real, imag} */,
  {32'h42770dd3, 32'hc20fc4d3} /* (4, 0, 11) {real, imag} */,
  {32'hbccb5000, 32'hc2cc627c} /* (4, 0, 10) {real, imag} */,
  {32'h430b83f2, 32'h4299802f} /* (4, 0, 9) {real, imag} */,
  {32'h42ea2170, 32'hc17f0be0} /* (4, 0, 8) {real, imag} */,
  {32'hc30e61f0, 32'hc23353b6} /* (4, 0, 7) {real, imag} */,
  {32'hc222c951, 32'hc29fb892} /* (4, 0, 6) {real, imag} */,
  {32'h41329750, 32'hc3187eb1} /* (4, 0, 5) {real, imag} */,
  {32'h42754747, 32'h42b13347} /* (4, 0, 4) {real, imag} */,
  {32'h429d0aa4, 32'hc322791b} /* (4, 0, 3) {real, imag} */,
  {32'h437725c6, 32'h41c318cb} /* (4, 0, 2) {real, imag} */,
  {32'hc42bf624, 32'h43ccd967} /* (4, 0, 1) {real, imag} */,
  {32'hc38faec1, 32'h43fc1558} /* (4, 0, 0) {real, imag} */,
  {32'h438b212e, 32'h44ca2031} /* (3, 31, 31) {real, imag} */,
  {32'hc3c5f1ad, 32'hc444bcfa} /* (3, 31, 30) {real, imag} */,
  {32'h437d3044, 32'hc379e8f7} /* (3, 31, 29) {real, imag} */,
  {32'hc29b7a82, 32'h437ebbff} /* (3, 31, 28) {real, imag} */,
  {32'hc33a1b36, 32'hc3b8baaa} /* (3, 31, 27) {real, imag} */,
  {32'h42955a09, 32'hc2c55144} /* (3, 31, 26) {real, imag} */,
  {32'h42454553, 32'h42b71530} /* (3, 31, 25) {real, imag} */,
  {32'hc3102c5c, 32'h401ab560} /* (3, 31, 24) {real, imag} */,
  {32'h428ca284, 32'hc1847ca0} /* (3, 31, 23) {real, imag} */,
  {32'h414395b0, 32'h3fc13540} /* (3, 31, 22) {real, imag} */,
  {32'hc1e0473c, 32'hc21af7f2} /* (3, 31, 21) {real, imag} */,
  {32'h41eedfc1, 32'hc1efbf23} /* (3, 31, 20) {real, imag} */,
  {32'h417e001e, 32'hc15c94bc} /* (3, 31, 19) {real, imag} */,
  {32'hc2c587d5, 32'hc1bb3c98} /* (3, 31, 18) {real, imag} */,
  {32'h42452447, 32'hc0882d00} /* (3, 31, 17) {real, imag} */,
  {32'h41715e44, 32'hc23f3618} /* (3, 31, 16) {real, imag} */,
  {32'h41700bfc, 32'h41625b80} /* (3, 31, 15) {real, imag} */,
  {32'h42b71b25, 32'hc2475e64} /* (3, 31, 14) {real, imag} */,
  {32'hc157b482, 32'h421169f7} /* (3, 31, 13) {real, imag} */,
  {32'hc143ca46, 32'h419624f3} /* (3, 31, 12) {real, imag} */,
  {32'h4300eb3a, 32'hc336d1ee} /* (3, 31, 11) {real, imag} */,
  {32'h4287fa64, 32'hc20096ba} /* (3, 31, 10) {real, imag} */,
  {32'h40a00cb8, 32'h42ef47f0} /* (3, 31, 9) {real, imag} */,
  {32'h4299005c, 32'hc2dbc563} /* (3, 31, 8) {real, imag} */,
  {32'hc1f0d0fa, 32'h4345a00c} /* (3, 31, 7) {real, imag} */,
  {32'hc08bdd50, 32'hc2a0a354} /* (3, 31, 6) {real, imag} */,
  {32'h4362772c, 32'hc389fb8a} /* (3, 31, 5) {real, imag} */,
  {32'h426cf194, 32'h43484a69} /* (3, 31, 4) {real, imag} */,
  {32'hc2f741e3, 32'hc27883e4} /* (3, 31, 3) {real, imag} */,
  {32'h42c41024, 32'hc3d490cc} /* (3, 31, 2) {real, imag} */,
  {32'hc413db37, 32'h442fc8ba} /* (3, 31, 1) {real, imag} */,
  {32'hc307e6ed, 32'h447244dc} /* (3, 31, 0) {real, imag} */,
  {32'h4386b62e, 32'hc438dfd0} /* (3, 30, 31) {real, imag} */,
  {32'hc3b92a70, 32'h441b7155} /* (3, 30, 30) {real, imag} */,
  {32'h426abfa6, 32'h4283af30} /* (3, 30, 29) {real, imag} */,
  {32'h4224eae2, 32'hc3ebc390} /* (3, 30, 28) {real, imag} */,
  {32'hc3266219, 32'h434c42a7} /* (3, 30, 27) {real, imag} */,
  {32'hc211aa9c, 32'h42a510d0} /* (3, 30, 26) {real, imag} */,
  {32'hc3173322, 32'hc2d54875} /* (3, 30, 25) {real, imag} */,
  {32'hc32c5786, 32'h430d74c8} /* (3, 30, 24) {real, imag} */,
  {32'h42bcfbff, 32'h42fd7860} /* (3, 30, 23) {real, imag} */,
  {32'hc1b1f798, 32'hc29febae} /* (3, 30, 22) {real, imag} */,
  {32'h42758d28, 32'h42cf9f8c} /* (3, 30, 21) {real, imag} */,
  {32'h4121cdda, 32'hc20125aa} /* (3, 30, 20) {real, imag} */,
  {32'hc1a62403, 32'hc168924a} /* (3, 30, 19) {real, imag} */,
  {32'h41c5d356, 32'hc24aac54} /* (3, 30, 18) {real, imag} */,
  {32'h4019f838, 32'hc0e441d0} /* (3, 30, 17) {real, imag} */,
  {32'h4002aa00, 32'hbd0c0000} /* (3, 30, 16) {real, imag} */,
  {32'hc1955c67, 32'h424c5c7a} /* (3, 30, 15) {real, imag} */,
  {32'hc28c216e, 32'h419fc5e8} /* (3, 30, 14) {real, imag} */,
  {32'hc1ea09f3, 32'h4147619e} /* (3, 30, 13) {real, imag} */,
  {32'hc19cf575, 32'hc194ad04} /* (3, 30, 12) {real, imag} */,
  {32'hc20305b8, 32'hc1637f0c} /* (3, 30, 11) {real, imag} */,
  {32'hc1866ff0, 32'hc17cff40} /* (3, 30, 10) {real, imag} */,
  {32'hc22e67a2, 32'h42099ebb} /* (3, 30, 9) {real, imag} */,
  {32'hc2bb9e2c, 32'h433cf2d6} /* (3, 30, 8) {real, imag} */,
  {32'hc1f2596c, 32'h42e34d2f} /* (3, 30, 7) {real, imag} */,
  {32'h4248bff0, 32'h431a2b39} /* (3, 30, 6) {real, imag} */,
  {32'hc2c12646, 32'h4328baad} /* (3, 30, 5) {real, imag} */,
  {32'h433c83a0, 32'hc19fef78} /* (3, 30, 4) {real, imag} */,
  {32'h42ce2aab, 32'h414ad61c} /* (3, 30, 3) {real, imag} */,
  {32'hc40083f8, 32'h44090cbf} /* (3, 30, 2) {real, imag} */,
  {32'h4346b570, 32'hc4994ca2} /* (3, 30, 1) {real, imag} */,
  {32'hc24383b0, 32'hc44000c4} /* (3, 30, 0) {real, imag} */,
  {32'h4113e8a8, 32'h439e6f1d} /* (3, 29, 31) {real, imag} */,
  {32'hc3e09e62, 32'h4121c110} /* (3, 29, 30) {real, imag} */,
  {32'h42543ba2, 32'h42d3e996} /* (3, 29, 29) {real, imag} */,
  {32'h431c5d4a, 32'hc1a923d0} /* (3, 29, 28) {real, imag} */,
  {32'hc3102551, 32'h41ccfea8} /* (3, 29, 27) {real, imag} */,
  {32'hc0130960, 32'hc2908352} /* (3, 29, 26) {real, imag} */,
  {32'h430edcd8, 32'hbf14bc40} /* (3, 29, 25) {real, imag} */,
  {32'hc28d34ab, 32'hc2fabd4c} /* (3, 29, 24) {real, imag} */,
  {32'h41efd600, 32'h4282d1f0} /* (3, 29, 23) {real, imag} */,
  {32'h423a4e4a, 32'hc2b3f0ac} /* (3, 29, 22) {real, imag} */,
  {32'hc09bea18, 32'hc237e99a} /* (3, 29, 21) {real, imag} */,
  {32'h424acd2b, 32'hc2b0fbe4} /* (3, 29, 20) {real, imag} */,
  {32'hc21b9c84, 32'hc1ac4697} /* (3, 29, 19) {real, imag} */,
  {32'hc23426b4, 32'h41d4392d} /* (3, 29, 18) {real, imag} */,
  {32'h419e39e6, 32'h418c56b8} /* (3, 29, 17) {real, imag} */,
  {32'h41e3fcbc, 32'hc1d0fbf4} /* (3, 29, 16) {real, imag} */,
  {32'hc23bd913, 32'h41a5a6f8} /* (3, 29, 15) {real, imag} */,
  {32'h415caf12, 32'h408f064c} /* (3, 29, 14) {real, imag} */,
  {32'h42018940, 32'hbf704320} /* (3, 29, 13) {real, imag} */,
  {32'hc1e5aac6, 32'h41ab65c4} /* (3, 29, 12) {real, imag} */,
  {32'h4291561a, 32'hc23518c0} /* (3, 29, 11) {real, imag} */,
  {32'hc30f0812, 32'h4206334f} /* (3, 29, 10) {real, imag} */,
  {32'h4291523a, 32'h42d9491c} /* (3, 29, 9) {real, imag} */,
  {32'hc264ae9a, 32'hc2d04b00} /* (3, 29, 8) {real, imag} */,
  {32'h431f8208, 32'hc1328a3c} /* (3, 29, 7) {real, imag} */,
  {32'h421e944e, 32'h41a0a336} /* (3, 29, 6) {real, imag} */,
  {32'hc33963ab, 32'hc34f28cb} /* (3, 29, 5) {real, imag} */,
  {32'h41af8a44, 32'h42ca7ff7} /* (3, 29, 4) {real, imag} */,
  {32'h416457d8, 32'h41808490} /* (3, 29, 3) {real, imag} */,
  {32'hc39deaa4, 32'h42efafe8} /* (3, 29, 2) {real, imag} */,
  {32'h433b0260, 32'hc3b692bb} /* (3, 29, 1) {real, imag} */,
  {32'hc235478a, 32'hc2926d07} /* (3, 29, 0) {real, imag} */,
  {32'h435e155f, 32'h44036c94} /* (3, 28, 31) {real, imag} */,
  {32'hc3120686, 32'hc3af3ed8} /* (3, 28, 30) {real, imag} */,
  {32'hc2237bb6, 32'hc2e855ba} /* (3, 28, 29) {real, imag} */,
  {32'h42b2074c, 32'h405a21f8} /* (3, 28, 28) {real, imag} */,
  {32'h42c67148, 32'h424d7946} /* (3, 28, 27) {real, imag} */,
  {32'h4290c6d7, 32'h42e99742} /* (3, 28, 26) {real, imag} */,
  {32'hc1124630, 32'h433c76e4} /* (3, 28, 25) {real, imag} */,
  {32'hc243e51b, 32'h427804ad} /* (3, 28, 24) {real, imag} */,
  {32'hc210a5ec, 32'hc219c7fc} /* (3, 28, 23) {real, imag} */,
  {32'hc18d24ee, 32'hc2dd50ba} /* (3, 28, 22) {real, imag} */,
  {32'hc275defd, 32'h41bc7584} /* (3, 28, 21) {real, imag} */,
  {32'hc151b681, 32'hc0980f0c} /* (3, 28, 20) {real, imag} */,
  {32'hc1562f1e, 32'h42619bbe} /* (3, 28, 19) {real, imag} */,
  {32'h42200990, 32'hc118001c} /* (3, 28, 18) {real, imag} */,
  {32'h420246c6, 32'h41211c80} /* (3, 28, 17) {real, imag} */,
  {32'h3e516000, 32'hc1c1b8c2} /* (3, 28, 16) {real, imag} */,
  {32'hc154865a, 32'hc138f4e0} /* (3, 28, 15) {real, imag} */,
  {32'hc1a77410, 32'hc28350d4} /* (3, 28, 14) {real, imag} */,
  {32'h41c760df, 32'h419bacd7} /* (3, 28, 13) {real, imag} */,
  {32'hc14fa033, 32'h41df1f25} /* (3, 28, 12) {real, imag} */,
  {32'hc24cfbdb, 32'hc265a594} /* (3, 28, 11) {real, imag} */,
  {32'hc273b3eb, 32'h429fc476} /* (3, 28, 10) {real, imag} */,
  {32'h428ec202, 32'h4294b460} /* (3, 28, 9) {real, imag} */,
  {32'hc118fdc0, 32'hc28242da} /* (3, 28, 8) {real, imag} */,
  {32'h42b069d2, 32'h42591b66} /* (3, 28, 7) {real, imag} */,
  {32'h43062036, 32'h413f47ec} /* (3, 28, 6) {real, imag} */,
  {32'hc28ad0b4, 32'h41bdbd94} /* (3, 28, 5) {real, imag} */,
  {32'h423c5c40, 32'h4244a3d0} /* (3, 28, 4) {real, imag} */,
  {32'h40a10dc4, 32'hbf119940} /* (3, 28, 3) {real, imag} */,
  {32'hc37a30ec, 32'hc3acdede} /* (3, 28, 2) {real, imag} */,
  {32'h435352d9, 32'h42ed73e2} /* (3, 28, 1) {real, imag} */,
  {32'h4332c5c4, 32'h42b27564} /* (3, 28, 0) {real, imag} */,
  {32'hc34570e8, 32'hc32fae1f} /* (3, 27, 31) {real, imag} */,
  {32'h426d1aa1, 32'h42de933e} /* (3, 27, 30) {real, imag} */,
  {32'hc1190572, 32'hc259c45e} /* (3, 27, 29) {real, imag} */,
  {32'hc29efca4, 32'hc2c6cf33} /* (3, 27, 28) {real, imag} */,
  {32'h4365269f, 32'h42cfc9a4} /* (3, 27, 27) {real, imag} */,
  {32'hc2567fa4, 32'h41e2442a} /* (3, 27, 26) {real, imag} */,
  {32'h42771937, 32'h42e4046c} /* (3, 27, 25) {real, imag} */,
  {32'hc1802457, 32'hc135ed80} /* (3, 27, 24) {real, imag} */,
  {32'h410f9626, 32'hc25c5db4} /* (3, 27, 23) {real, imag} */,
  {32'hc184c455, 32'hc2758861} /* (3, 27, 22) {real, imag} */,
  {32'hc20c0560, 32'h41762245} /* (3, 27, 21) {real, imag} */,
  {32'hc1b20d1c, 32'hc1be2121} /* (3, 27, 20) {real, imag} */,
  {32'h4250f690, 32'h41196b7a} /* (3, 27, 19) {real, imag} */,
  {32'h4194f382, 32'hc0c26768} /* (3, 27, 18) {real, imag} */,
  {32'h40e11f18, 32'h4217c565} /* (3, 27, 17) {real, imag} */,
  {32'hc175cf30, 32'hc0e8dee0} /* (3, 27, 16) {real, imag} */,
  {32'h41a0bed6, 32'h41a7a2a6} /* (3, 27, 15) {real, imag} */,
  {32'hc1b5c9c6, 32'hc1fccbf2} /* (3, 27, 14) {real, imag} */,
  {32'h41a80868, 32'hc1c3eabd} /* (3, 27, 13) {real, imag} */,
  {32'hc1af5c54, 32'hc136ecd6} /* (3, 27, 12) {real, imag} */,
  {32'hc11ffb60, 32'h4210ff11} /* (3, 27, 11) {real, imag} */,
  {32'hc2499cf6, 32'h413c8a24} /* (3, 27, 10) {real, imag} */,
  {32'h41f7c75f, 32'hc1a86f83} /* (3, 27, 9) {real, imag} */,
  {32'h4282201a, 32'h42b57d50} /* (3, 27, 8) {real, imag} */,
  {32'h42c6438e, 32'hc1c362ae} /* (3, 27, 7) {real, imag} */,
  {32'h42108d38, 32'hc2087de9} /* (3, 27, 6) {real, imag} */,
  {32'hc30234f3, 32'h4324c7c0} /* (3, 27, 5) {real, imag} */,
  {32'h42964e42, 32'hc2d16195} /* (3, 27, 4) {real, imag} */,
  {32'hc1933b19, 32'h41f1b0dc} /* (3, 27, 3) {real, imag} */,
  {32'hc33421ab, 32'h43124807} /* (3, 27, 2) {real, imag} */,
  {32'hc1d5ee20, 32'hc390bc77} /* (3, 27, 1) {real, imag} */,
  {32'h42c5d6b2, 32'hc3b26d66} /* (3, 27, 0) {real, imag} */,
  {32'hc09be3f0, 32'hc2bf61cc} /* (3, 26, 31) {real, imag} */,
  {32'hc25f40d4, 32'hc25d5d05} /* (3, 26, 30) {real, imag} */,
  {32'h4215a302, 32'h40edc3b8} /* (3, 26, 29) {real, imag} */,
  {32'h42bc13b7, 32'h4227448a} /* (3, 26, 28) {real, imag} */,
  {32'h4251464b, 32'h41b57e25} /* (3, 26, 27) {real, imag} */,
  {32'h4265c9d8, 32'h431af928} /* (3, 26, 26) {real, imag} */,
  {32'hc2c62343, 32'h42d63e79} /* (3, 26, 25) {real, imag} */,
  {32'h42d37c60, 32'h4210501c} /* (3, 26, 24) {real, imag} */,
  {32'hc2e350d3, 32'hc2ad6267} /* (3, 26, 23) {real, imag} */,
  {32'h412f3f10, 32'hc03f29f0} /* (3, 26, 22) {real, imag} */,
  {32'hc230158c, 32'h42b29ab7} /* (3, 26, 21) {real, imag} */,
  {32'h40e172f4, 32'h408188e6} /* (3, 26, 20) {real, imag} */,
  {32'hc20969b1, 32'hc0b7be58} /* (3, 26, 19) {real, imag} */,
  {32'hc1d9731d, 32'hc1da4a30} /* (3, 26, 18) {real, imag} */,
  {32'h3fd42400, 32'hc18d86db} /* (3, 26, 17) {real, imag} */,
  {32'hc0ef9ea8, 32'hc156ffd0} /* (3, 26, 16) {real, imag} */,
  {32'h42093aa3, 32'hc1866961} /* (3, 26, 15) {real, imag} */,
  {32'h41d4e705, 32'hc1096a5d} /* (3, 26, 14) {real, imag} */,
  {32'hc232d10f, 32'hc2774e1b} /* (3, 26, 13) {real, imag} */,
  {32'hc197c56d, 32'hc1d7df98} /* (3, 26, 12) {real, imag} */,
  {32'h4120ab62, 32'h415c8748} /* (3, 26, 11) {real, imag} */,
  {32'hc05981f2, 32'h42ae0626} /* (3, 26, 10) {real, imag} */,
  {32'hc1af90d4, 32'hc1256f98} /* (3, 26, 9) {real, imag} */,
  {32'hc214b644, 32'hc198993b} /* (3, 26, 8) {real, imag} */,
  {32'h428587df, 32'h430383bb} /* (3, 26, 7) {real, imag} */,
  {32'hc21f225c, 32'h4113d9f0} /* (3, 26, 6) {real, imag} */,
  {32'h42731ee9, 32'h41f67b6b} /* (3, 26, 5) {real, imag} */,
  {32'h425f7566, 32'h42c1bc8b} /* (3, 26, 4) {real, imag} */,
  {32'h42cad4e3, 32'hc2044557} /* (3, 26, 3) {real, imag} */,
  {32'h41fbbe17, 32'hc1b28af6} /* (3, 26, 2) {real, imag} */,
  {32'h420cee83, 32'hc1c69302} /* (3, 26, 1) {real, imag} */,
  {32'h427a2d6d, 32'hc2cda874} /* (3, 26, 0) {real, imag} */,
  {32'h42f87b13, 32'h43330bb2} /* (3, 25, 31) {real, imag} */,
  {32'hc323fd6e, 32'h428ab052} /* (3, 25, 30) {real, imag} */,
  {32'h41fb7850, 32'hc2702370} /* (3, 25, 29) {real, imag} */,
  {32'h426199da, 32'h42ad6164} /* (3, 25, 28) {real, imag} */,
  {32'hc2b011ea, 32'h4230ef1a} /* (3, 25, 27) {real, imag} */,
  {32'hc29e5214, 32'h4254c0d6} /* (3, 25, 26) {real, imag} */,
  {32'hc20930ea, 32'hc181bfb0} /* (3, 25, 25) {real, imag} */,
  {32'h41b3f990, 32'hc3152804} /* (3, 25, 24) {real, imag} */,
  {32'h421fffe0, 32'h4233d37e} /* (3, 25, 23) {real, imag} */,
  {32'hc25d0e95, 32'h424815d9} /* (3, 25, 22) {real, imag} */,
  {32'h42065ef2, 32'hc18ba666} /* (3, 25, 21) {real, imag} */,
  {32'hc1a084bb, 32'h41da4da6} /* (3, 25, 20) {real, imag} */,
  {32'h41354234, 32'hc2086c03} /* (3, 25, 19) {real, imag} */,
  {32'hc0faef70, 32'hc0f654bc} /* (3, 25, 18) {real, imag} */,
  {32'h417f7af0, 32'hc1bf5091} /* (3, 25, 17) {real, imag} */,
  {32'hc21510c5, 32'h418836d0} /* (3, 25, 16) {real, imag} */,
  {32'hc0b14560, 32'hc2422016} /* (3, 25, 15) {real, imag} */,
  {32'hc1a43fc4, 32'h41ad5425} /* (3, 25, 14) {real, imag} */,
  {32'h41ae0fb2, 32'h411e18cc} /* (3, 25, 13) {real, imag} */,
  {32'h40287778, 32'hc2819a86} /* (3, 25, 12) {real, imag} */,
  {32'h41dbefbc, 32'h423da241} /* (3, 25, 11) {real, imag} */,
  {32'hc22f05ad, 32'hc1ac0b42} /* (3, 25, 10) {real, imag} */,
  {32'hc1d08f05, 32'h41d67b6c} /* (3, 25, 9) {real, imag} */,
  {32'hc13b918f, 32'hc20cc103} /* (3, 25, 8) {real, imag} */,
  {32'h4158a14e, 32'hc31122f2} /* (3, 25, 7) {real, imag} */,
  {32'h41bf36a4, 32'hc2223e90} /* (3, 25, 6) {real, imag} */,
  {32'hc2639814, 32'h423f6420} /* (3, 25, 5) {real, imag} */,
  {32'h430aed18, 32'hc2d6cd04} /* (3, 25, 4) {real, imag} */,
  {32'h42e4fcf0, 32'hc2a13a6c} /* (3, 25, 3) {real, imag} */,
  {32'h4059aba0, 32'h422159bb} /* (3, 25, 2) {real, imag} */,
  {32'h41e4c4c4, 32'h42decd05} /* (3, 25, 1) {real, imag} */,
  {32'h42444c45, 32'h4344d689} /* (3, 25, 0) {real, imag} */,
  {32'hc3128969, 32'hc30a31a7} /* (3, 24, 31) {real, imag} */,
  {32'h42b02dba, 32'hc26bdbd4} /* (3, 24, 30) {real, imag} */,
  {32'h428dd0b8, 32'h42cb8a1c} /* (3, 24, 29) {real, imag} */,
  {32'hc1d981c1, 32'h420cc7f4} /* (3, 24, 28) {real, imag} */,
  {32'h41331e4e, 32'h43139231} /* (3, 24, 27) {real, imag} */,
  {32'h42b5dad0, 32'hc20d4bfe} /* (3, 24, 26) {real, imag} */,
  {32'h42b74bbe, 32'hc23288d4} /* (3, 24, 25) {real, imag} */,
  {32'h4230a6bf, 32'hc23a5244} /* (3, 24, 24) {real, imag} */,
  {32'hc28a41fd, 32'h4214b17b} /* (3, 24, 23) {real, imag} */,
  {32'hc1463556, 32'hc2c42f08} /* (3, 24, 22) {real, imag} */,
  {32'h42bb758e, 32'h41a6649c} /* (3, 24, 21) {real, imag} */,
  {32'hbfdbb580, 32'h4203720d} /* (3, 24, 20) {real, imag} */,
  {32'hc215f490, 32'h410874d1} /* (3, 24, 19) {real, imag} */,
  {32'h4159a48a, 32'h419185d6} /* (3, 24, 18) {real, imag} */,
  {32'hc24bbbda, 32'hc0a8d478} /* (3, 24, 17) {real, imag} */,
  {32'hc0ddf216, 32'h409873b8} /* (3, 24, 16) {real, imag} */,
  {32'h41caac78, 32'hc0e43ec8} /* (3, 24, 15) {real, imag} */,
  {32'h40c53c54, 32'h4145cd1c} /* (3, 24, 14) {real, imag} */,
  {32'h417a5bf8, 32'h41c4ac58} /* (3, 24, 13) {real, imag} */,
  {32'hc1abd35e, 32'hc14f728b} /* (3, 24, 12) {real, imag} */,
  {32'hc14a178c, 32'hc22ca752} /* (3, 24, 11) {real, imag} */,
  {32'h420b67e4, 32'h41429254} /* (3, 24, 10) {real, imag} */,
  {32'h41aeff89, 32'hc2e89dc2} /* (3, 24, 9) {real, imag} */,
  {32'hc27cb637, 32'hc14aeeae} /* (3, 24, 8) {real, imag} */,
  {32'h4184e67a, 32'hc285a0af} /* (3, 24, 7) {real, imag} */,
  {32'hc12b25b0, 32'hc202ade4} /* (3, 24, 6) {real, imag} */,
  {32'hc2625e7e, 32'hc2b82c5e} /* (3, 24, 5) {real, imag} */,
  {32'h42b4b4a2, 32'hc247a290} /* (3, 24, 4) {real, imag} */,
  {32'hc33af478, 32'h41bd16fe} /* (3, 24, 3) {real, imag} */,
  {32'h418df328, 32'h43666a17} /* (3, 24, 2) {real, imag} */,
  {32'h418d1e08, 32'hc38ab418} /* (3, 24, 1) {real, imag} */,
  {32'hbf8267b8, 32'hc2d93bd0} /* (3, 24, 0) {real, imag} */,
  {32'hc297e79a, 32'h42a59518} /* (3, 23, 31) {real, imag} */,
  {32'hbfac9b80, 32'hc2857be4} /* (3, 23, 30) {real, imag} */,
  {32'hc10562c8, 32'h3f0fccd0} /* (3, 23, 29) {real, imag} */,
  {32'hc240add6, 32'hc191f6cc} /* (3, 23, 28) {real, imag} */,
  {32'h42578040, 32'h4132cd32} /* (3, 23, 27) {real, imag} */,
  {32'hc27e768d, 32'h413dca92} /* (3, 23, 26) {real, imag} */,
  {32'hc1d013f0, 32'h428df7a0} /* (3, 23, 25) {real, imag} */,
  {32'hc2644dc6, 32'hc20fefb0} /* (3, 23, 24) {real, imag} */,
  {32'h40ea1370, 32'h3f51edb0} /* (3, 23, 23) {real, imag} */,
  {32'h420a9b88, 32'hc1d610bf} /* (3, 23, 22) {real, imag} */,
  {32'hc1214a9c, 32'h420e380c} /* (3, 23, 21) {real, imag} */,
  {32'h3e64adc0, 32'h4217f69c} /* (3, 23, 20) {real, imag} */,
  {32'hc1d4bf80, 32'h41720502} /* (3, 23, 19) {real, imag} */,
  {32'h413ed22e, 32'h41acef00} /* (3, 23, 18) {real, imag} */,
  {32'h420a37da, 32'h40fa0df0} /* (3, 23, 17) {real, imag} */,
  {32'h40802860, 32'h419c67ee} /* (3, 23, 16) {real, imag} */,
  {32'h414c947a, 32'h422308e2} /* (3, 23, 15) {real, imag} */,
  {32'hc0dd0820, 32'hc15677b4} /* (3, 23, 14) {real, imag} */,
  {32'h425de838, 32'hc1d0cecf} /* (3, 23, 13) {real, imag} */,
  {32'hbf9dcd68, 32'h424335f8} /* (3, 23, 12) {real, imag} */,
  {32'hc204fa0d, 32'hc1a342cb} /* (3, 23, 11) {real, imag} */,
  {32'hc1be23cc, 32'hc092a084} /* (3, 23, 10) {real, imag} */,
  {32'h425035ee, 32'hc12b1165} /* (3, 23, 9) {real, imag} */,
  {32'hc22bd04e, 32'h40061c90} /* (3, 23, 8) {real, imag} */,
  {32'h40166744, 32'hc0cb49e8} /* (3, 23, 7) {real, imag} */,
  {32'h41848122, 32'hc23ccd06} /* (3, 23, 6) {real, imag} */,
  {32'hc2e693d0, 32'hc24a8502} /* (3, 23, 5) {real, imag} */,
  {32'h426d8282, 32'hc2185003} /* (3, 23, 4) {real, imag} */,
  {32'h4237e092, 32'h4183dd1c} /* (3, 23, 3) {real, imag} */,
  {32'hc24a2376, 32'hc205b718} /* (3, 23, 2) {real, imag} */,
  {32'h43388caf, 32'hc29c9c56} /* (3, 23, 1) {real, imag} */,
  {32'h42258dbf, 32'h425fe889} /* (3, 23, 0) {real, imag} */,
  {32'hc232449c, 32'hc0f6292c} /* (3, 22, 31) {real, imag} */,
  {32'h42b70c3c, 32'hc0a186d0} /* (3, 22, 30) {real, imag} */,
  {32'h43193ed6, 32'hc2c2956e} /* (3, 22, 29) {real, imag} */,
  {32'hc165ca9e, 32'hc2eafa26} /* (3, 22, 28) {real, imag} */,
  {32'hc26fcb39, 32'hc2622a63} /* (3, 22, 27) {real, imag} */,
  {32'hc24e9e8b, 32'h40dbfeac} /* (3, 22, 26) {real, imag} */,
  {32'hc2910626, 32'hc19fb762} /* (3, 22, 25) {real, imag} */,
  {32'h41067ca8, 32'h42046cd7} /* (3, 22, 24) {real, imag} */,
  {32'h420e9fcf, 32'hc270bd0c} /* (3, 22, 23) {real, imag} */,
  {32'h41d7238e, 32'hc04a8508} /* (3, 22, 22) {real, imag} */,
  {32'hc1039e86, 32'h41ecb538} /* (3, 22, 21) {real, imag} */,
  {32'hc0b4d242, 32'h41b12439} /* (3, 22, 20) {real, imag} */,
  {32'h420a354c, 32'hc24c9b4e} /* (3, 22, 19) {real, imag} */,
  {32'h417d609c, 32'h41915d0f} /* (3, 22, 18) {real, imag} */,
  {32'hc11b3326, 32'hc10f4595} /* (3, 22, 17) {real, imag} */,
  {32'hc1897b5c, 32'h4068cd00} /* (3, 22, 16) {real, imag} */,
  {32'hc1054ade, 32'hbfdde958} /* (3, 22, 15) {real, imag} */,
  {32'hc20cc029, 32'h419fa615} /* (3, 22, 14) {real, imag} */,
  {32'hc15b5dfe, 32'hbe233180} /* (3, 22, 13) {real, imag} */,
  {32'hbff07ad8, 32'h41a66749} /* (3, 22, 12) {real, imag} */,
  {32'h424fba9a, 32'hc1931ffc} /* (3, 22, 11) {real, imag} */,
  {32'hc116a544, 32'h41b643f5} /* (3, 22, 10) {real, imag} */,
  {32'hc1b9da56, 32'hc115c860} /* (3, 22, 9) {real, imag} */,
  {32'h424bd0aa, 32'hc16ea763} /* (3, 22, 8) {real, imag} */,
  {32'hc2db9f34, 32'h40db5ea6} /* (3, 22, 7) {real, imag} */,
  {32'hc0bb8568, 32'hc143454e} /* (3, 22, 6) {real, imag} */,
  {32'hc2ac7088, 32'h41b7fd9a} /* (3, 22, 5) {real, imag} */,
  {32'h4235e2de, 32'h43235727} /* (3, 22, 4) {real, imag} */,
  {32'hbf584d80, 32'h429075dc} /* (3, 22, 3) {real, imag} */,
  {32'hc31ec78c, 32'hc2fbe1ff} /* (3, 22, 2) {real, imag} */,
  {32'h42c817ba, 32'h423a4dc8} /* (3, 22, 1) {real, imag} */,
  {32'h42849f61, 32'h4278072a} /* (3, 22, 0) {real, imag} */,
  {32'hc2b8e774, 32'hc23f7807} /* (3, 21, 31) {real, imag} */,
  {32'h42950fb2, 32'h42068f4e} /* (3, 21, 30) {real, imag} */,
  {32'h42b4224c, 32'h4102b159} /* (3, 21, 29) {real, imag} */,
  {32'h4287bb99, 32'h40d5f778} /* (3, 21, 28) {real, imag} */,
  {32'hc210d74a, 32'hc20b5067} /* (3, 21, 27) {real, imag} */,
  {32'h425c4067, 32'h42861f04} /* (3, 21, 26) {real, imag} */,
  {32'hc06b9e70, 32'hc151321b} /* (3, 21, 25) {real, imag} */,
  {32'hbf1e3700, 32'hc0fde0dc} /* (3, 21, 24) {real, imag} */,
  {32'h4129fa38, 32'h41b35a3c} /* (3, 21, 23) {real, imag} */,
  {32'h42080c22, 32'h40996903} /* (3, 21, 22) {real, imag} */,
  {32'hc1d52a7d, 32'h3ff7f640} /* (3, 21, 21) {real, imag} */,
  {32'hc08ddfe1, 32'hc1f884e9} /* (3, 21, 20) {real, imag} */,
  {32'h419ae9fb, 32'hc0aba20a} /* (3, 21, 19) {real, imag} */,
  {32'hc204bfde, 32'hc1a6a20b} /* (3, 21, 18) {real, imag} */,
  {32'hc0ec3d20, 32'h416de1ae} /* (3, 21, 17) {real, imag} */,
  {32'h3f9de3e0, 32'h3ee62900} /* (3, 21, 16) {real, imag} */,
  {32'h412d5b48, 32'hc1919e0f} /* (3, 21, 15) {real, imag} */,
  {32'hc1c82bd0, 32'h40cd52dc} /* (3, 21, 14) {real, imag} */,
  {32'hc16a7b7a, 32'h40925aea} /* (3, 21, 13) {real, imag} */,
  {32'h412e2100, 32'h412afede} /* (3, 21, 12) {real, imag} */,
  {32'hc129a446, 32'h4212d836} /* (3, 21, 11) {real, imag} */,
  {32'h417859ce, 32'hc15237ea} /* (3, 21, 10) {real, imag} */,
  {32'h40704060, 32'hc21106ba} /* (3, 21, 9) {real, imag} */,
  {32'h4238f2d2, 32'hc2604cc0} /* (3, 21, 8) {real, imag} */,
  {32'hc25d5aa3, 32'hc22c7b75} /* (3, 21, 7) {real, imag} */,
  {32'hc1eff2ea, 32'hc23d41b4} /* (3, 21, 6) {real, imag} */,
  {32'h4256309a, 32'hc2149e23} /* (3, 21, 5) {real, imag} */,
  {32'hc29b5269, 32'h429318c2} /* (3, 21, 4) {real, imag} */,
  {32'h40f84228, 32'h41b9b21c} /* (3, 21, 3) {real, imag} */,
  {32'h42634094, 32'h42f53af5} /* (3, 21, 2) {real, imag} */,
  {32'hc1ee0242, 32'hc218340d} /* (3, 21, 1) {real, imag} */,
  {32'hc2b762d6, 32'hc25f2424} /* (3, 21, 0) {real, imag} */,
  {32'h415f142c, 32'h41da0870} /* (3, 20, 31) {real, imag} */,
  {32'h411cf7e4, 32'hc24fb951} /* (3, 20, 30) {real, imag} */,
  {32'hbe635e00, 32'h4174aa9a} /* (3, 20, 29) {real, imag} */,
  {32'h4141555f, 32'h419a2bc2} /* (3, 20, 28) {real, imag} */,
  {32'h420bb7e3, 32'hc15c4991} /* (3, 20, 27) {real, imag} */,
  {32'h41cb6b9e, 32'h4117bdac} /* (3, 20, 26) {real, imag} */,
  {32'hc2d8ca08, 32'hc2495334} /* (3, 20, 25) {real, imag} */,
  {32'h42417d35, 32'h40292ebc} /* (3, 20, 24) {real, imag} */,
  {32'h3f2c1e20, 32'h3f1ca020} /* (3, 20, 23) {real, imag} */,
  {32'h41f453cb, 32'hbfd9dd04} /* (3, 20, 22) {real, imag} */,
  {32'hc19bbc1c, 32'hc04ed0bc} /* (3, 20, 21) {real, imag} */,
  {32'h4178b58d, 32'hc1c53978} /* (3, 20, 20) {real, imag} */,
  {32'hc11cbc82, 32'hc18fb57a} /* (3, 20, 19) {real, imag} */,
  {32'h40748478, 32'hc159223a} /* (3, 20, 18) {real, imag} */,
  {32'h3f74aed0, 32'h419e8ed8} /* (3, 20, 17) {real, imag} */,
  {32'h3f2994a0, 32'hc01d9470} /* (3, 20, 16) {real, imag} */,
  {32'h3fc41ee8, 32'h412d4dfe} /* (3, 20, 15) {real, imag} */,
  {32'h40b6adb4, 32'h40d589d5} /* (3, 20, 14) {real, imag} */,
  {32'hc1d9960f, 32'hc1ad5c78} /* (3, 20, 13) {real, imag} */,
  {32'h40956592, 32'hc00aed1c} /* (3, 20, 12) {real, imag} */,
  {32'h4159db49, 32'hc192ba30} /* (3, 20, 11) {real, imag} */,
  {32'hbf6c63c0, 32'hc10e7468} /* (3, 20, 10) {real, imag} */,
  {32'h41249dfa, 32'hc24daae6} /* (3, 20, 9) {real, imag} */,
  {32'h3f1fc740, 32'h411ac4d3} /* (3, 20, 8) {real, imag} */,
  {32'h4287c204, 32'hc1e62e40} /* (3, 20, 7) {real, imag} */,
  {32'hc0f5f32a, 32'hc155240e} /* (3, 20, 6) {real, imag} */,
  {32'hbe166f00, 32'hc0f3433e} /* (3, 20, 5) {real, imag} */,
  {32'h4152f407, 32'hc1042d13} /* (3, 20, 4) {real, imag} */,
  {32'h42cbb245, 32'hc2299bc2} /* (3, 20, 3) {real, imag} */,
  {32'hc2679357, 32'h42160d4b} /* (3, 20, 2) {real, imag} */,
  {32'hc275ba97, 32'h4282e989} /* (3, 20, 1) {real, imag} */,
  {32'h423c8df4, 32'hc2140b69} /* (3, 20, 0) {real, imag} */,
  {32'hc0aee6d8, 32'hc095839c} /* (3, 19, 31) {real, imag} */,
  {32'hc28caf72, 32'hc1954501} /* (3, 19, 30) {real, imag} */,
  {32'hc1b08511, 32'h423a78f5} /* (3, 19, 29) {real, imag} */,
  {32'hc18ebc2c, 32'h40842240} /* (3, 19, 28) {real, imag} */,
  {32'hc18de877, 32'h40e7bb96} /* (3, 19, 27) {real, imag} */,
  {32'h41573000, 32'h41bcb2bb} /* (3, 19, 26) {real, imag} */,
  {32'h40b4b850, 32'hc19694b2} /* (3, 19, 25) {real, imag} */,
  {32'hc22cc102, 32'h42606242} /* (3, 19, 24) {real, imag} */,
  {32'h41d2703e, 32'hc20fc7c1} /* (3, 19, 23) {real, imag} */,
  {32'hc138b466, 32'h411a1ff6} /* (3, 19, 22) {real, imag} */,
  {32'hbf01bcf8, 32'hbfd34230} /* (3, 19, 21) {real, imag} */,
  {32'hc17de3f4, 32'h3fdfb93a} /* (3, 19, 20) {real, imag} */,
  {32'hc0105586, 32'h416a14c6} /* (3, 19, 19) {real, imag} */,
  {32'hc0b9f1de, 32'h40728a08} /* (3, 19, 18) {real, imag} */,
  {32'hc0f41ebc, 32'h4093ef56} /* (3, 19, 17) {real, imag} */,
  {32'hbf19d340, 32'h413a8abe} /* (3, 19, 16) {real, imag} */,
  {32'hbfd2abd0, 32'h4069dc7c} /* (3, 19, 15) {real, imag} */,
  {32'h40d9bfea, 32'h40317d1c} /* (3, 19, 14) {real, imag} */,
  {32'hc0726c8e, 32'h41a13f5b} /* (3, 19, 13) {real, imag} */,
  {32'hc12e40b4, 32'hc0830360} /* (3, 19, 12) {real, imag} */,
  {32'hc12c6a38, 32'h41c04750} /* (3, 19, 11) {real, imag} */,
  {32'hc1a60419, 32'hc112f10a} /* (3, 19, 10) {real, imag} */,
  {32'h42561cfd, 32'h42095707} /* (3, 19, 9) {real, imag} */,
  {32'hbff03200, 32'hc19b8eeb} /* (3, 19, 8) {real, imag} */,
  {32'hc18a5c5a, 32'hc164b474} /* (3, 19, 7) {real, imag} */,
  {32'hc1817b96, 32'h41f4c927} /* (3, 19, 6) {real, imag} */,
  {32'hc0b7e9b4, 32'h41ebdb76} /* (3, 19, 5) {real, imag} */,
  {32'hc20550ac, 32'hc1747700} /* (3, 19, 4) {real, imag} */,
  {32'h4210456b, 32'hc1c0fdfe} /* (3, 19, 3) {real, imag} */,
  {32'h40b77220, 32'hc1880d4b} /* (3, 19, 2) {real, imag} */,
  {32'h42a66380, 32'h423b228e} /* (3, 19, 1) {real, imag} */,
  {32'hc1aa9dca, 32'h4209b4c2} /* (3, 19, 0) {real, imag} */,
  {32'hc2592f62, 32'h414525b0} /* (3, 18, 31) {real, imag} */,
  {32'hc1060c31, 32'h4213f6f2} /* (3, 18, 30) {real, imag} */,
  {32'hc11af6f4, 32'hc187687d} /* (3, 18, 29) {real, imag} */,
  {32'hc1dcd7e9, 32'hc08277b8} /* (3, 18, 28) {real, imag} */,
  {32'h420c26c6, 32'hbfd8433c} /* (3, 18, 27) {real, imag} */,
  {32'hc0d6acbd, 32'hc11db2c6} /* (3, 18, 26) {real, imag} */,
  {32'h41901fbb, 32'hc11ac518} /* (3, 18, 25) {real, imag} */,
  {32'h421ffa6e, 32'h410d7e40} /* (3, 18, 24) {real, imag} */,
  {32'hc24a3b22, 32'hc151a126} /* (3, 18, 23) {real, imag} */,
  {32'h418a5067, 32'hc1e6c589} /* (3, 18, 22) {real, imag} */,
  {32'h40da0040, 32'hc1f6ff7c} /* (3, 18, 21) {real, imag} */,
  {32'h413c64ec, 32'h4109d70a} /* (3, 18, 20) {real, imag} */,
  {32'h414c26d4, 32'hc129770d} /* (3, 18, 19) {real, imag} */,
  {32'hc10f1944, 32'h411a1a36} /* (3, 18, 18) {real, imag} */,
  {32'hc0b80e40, 32'hc0b6b443} /* (3, 18, 17) {real, imag} */,
  {32'h413edba2, 32'hbffc3de8} /* (3, 18, 16) {real, imag} */,
  {32'h40053f00, 32'hc0b6b553} /* (3, 18, 15) {real, imag} */,
  {32'hc09bcb85, 32'hc11176da} /* (3, 18, 14) {real, imag} */,
  {32'h41299ee2, 32'hc126a845} /* (3, 18, 13) {real, imag} */,
  {32'hc0090b70, 32'hc0a9df88} /* (3, 18, 12) {real, imag} */,
  {32'hc20ae42e, 32'hc08f1050} /* (3, 18, 11) {real, imag} */,
  {32'h4116a772, 32'hc19dfb7b} /* (3, 18, 10) {real, imag} */,
  {32'h40f83344, 32'hc1828025} /* (3, 18, 9) {real, imag} */,
  {32'hc170f6b2, 32'h4246ecd2} /* (3, 18, 8) {real, imag} */,
  {32'h421feaac, 32'h4175da48} /* (3, 18, 7) {real, imag} */,
  {32'hc1b13a19, 32'h4028782a} /* (3, 18, 6) {real, imag} */,
  {32'hbf141120, 32'h40052af6} /* (3, 18, 5) {real, imag} */,
  {32'hc0841acc, 32'hc1dbcd59} /* (3, 18, 4) {real, imag} */,
  {32'hc215aad1, 32'hc159017d} /* (3, 18, 3) {real, imag} */,
  {32'hc0dd0cc3, 32'h42843c23} /* (3, 18, 2) {real, imag} */,
  {32'hc29e17f7, 32'hc2428931} /* (3, 18, 1) {real, imag} */,
  {32'hc28da347, 32'h41964cbe} /* (3, 18, 0) {real, imag} */,
  {32'h4182b63e, 32'h41926500} /* (3, 17, 31) {real, imag} */,
  {32'hc189cdca, 32'h413bd64e} /* (3, 17, 30) {real, imag} */,
  {32'hc17a73ae, 32'h41275e32} /* (3, 17, 29) {real, imag} */,
  {32'hc0950918, 32'hc21799a4} /* (3, 17, 28) {real, imag} */,
  {32'h4196c9f7, 32'h41a85aa9} /* (3, 17, 27) {real, imag} */,
  {32'hc1001d20, 32'hc17f6dbc} /* (3, 17, 26) {real, imag} */,
  {32'h418d532c, 32'hc12d16ea} /* (3, 17, 25) {real, imag} */,
  {32'hc15cde8a, 32'hc19dec32} /* (3, 17, 24) {real, imag} */,
  {32'h405702ae, 32'hc1872b81} /* (3, 17, 23) {real, imag} */,
  {32'hc1822c33, 32'h416544aa} /* (3, 17, 22) {real, imag} */,
  {32'hbce35200, 32'hbfb9c150} /* (3, 17, 21) {real, imag} */,
  {32'hc0caa182, 32'hc0a21812} /* (3, 17, 20) {real, imag} */,
  {32'h3f2f2a00, 32'h4037837a} /* (3, 17, 19) {real, imag} */,
  {32'hbcf44300, 32'hc1904980} /* (3, 17, 18) {real, imag} */,
  {32'hc064c2f8, 32'h3fb26c18} /* (3, 17, 17) {real, imag} */,
  {32'hc158cf85, 32'h3fc61e60} /* (3, 17, 16) {real, imag} */,
  {32'h40a68d4c, 32'h40bb8be6} /* (3, 17, 15) {real, imag} */,
  {32'hc11b413a, 32'h41013485} /* (3, 17, 14) {real, imag} */,
  {32'hc1547d2c, 32'h418ef485} /* (3, 17, 13) {real, imag} */,
  {32'hc1381afd, 32'h4196bb42} /* (3, 17, 12) {real, imag} */,
  {32'hc12c9d4b, 32'hc1a118b5} /* (3, 17, 11) {real, imag} */,
  {32'h4173307e, 32'hc148ef36} /* (3, 17, 10) {real, imag} */,
  {32'h417e315c, 32'hc08134fc} /* (3, 17, 9) {real, imag} */,
  {32'h419acc97, 32'h3f9c1128} /* (3, 17, 8) {real, imag} */,
  {32'h41accfe0, 32'hbfcddd10} /* (3, 17, 7) {real, imag} */,
  {32'h41943d4e, 32'hc0061612} /* (3, 17, 6) {real, imag} */,
  {32'h41edb577, 32'hbfb3cbb0} /* (3, 17, 5) {real, imag} */,
  {32'hc16145fe, 32'hc0dc6f14} /* (3, 17, 4) {real, imag} */,
  {32'hc2808cc0, 32'h41cee3a7} /* (3, 17, 3) {real, imag} */,
  {32'hc194af8a, 32'h411fccb0} /* (3, 17, 2) {real, imag} */,
  {32'h42a17b80, 32'hc2277b2c} /* (3, 17, 1) {real, imag} */,
  {32'hc2337e84, 32'h41b18582} /* (3, 17, 0) {real, imag} */,
  {32'hc0af30b4, 32'hc03c0a68} /* (3, 16, 31) {real, imag} */,
  {32'h40d90fac, 32'hbf128988} /* (3, 16, 30) {real, imag} */,
  {32'h41eb0303, 32'h422e40de} /* (3, 16, 29) {real, imag} */,
  {32'h411c1ec0, 32'hc00c4d38} /* (3, 16, 28) {real, imag} */,
  {32'h414fe293, 32'hc16d7850} /* (3, 16, 27) {real, imag} */,
  {32'h4072a92a, 32'hc178a9f9} /* (3, 16, 26) {real, imag} */,
  {32'hc1aebb2a, 32'h41b31b3b} /* (3, 16, 25) {real, imag} */,
  {32'h41fba7bf, 32'hc1be59d0} /* (3, 16, 24) {real, imag} */,
  {32'h40886756, 32'h40cb3669} /* (3, 16, 23) {real, imag} */,
  {32'hc125e91a, 32'h41a2c417} /* (3, 16, 22) {real, imag} */,
  {32'hc0e6fa9a, 32'hc111ab0c} /* (3, 16, 21) {real, imag} */,
  {32'hc0856fe5, 32'h4129079e} /* (3, 16, 20) {real, imag} */,
  {32'h40333a05, 32'h40ba6856} /* (3, 16, 19) {real, imag} */,
  {32'h4122937e, 32'h40ae75e4} /* (3, 16, 18) {real, imag} */,
  {32'hbffacd48, 32'hc03ed0c0} /* (3, 16, 17) {real, imag} */,
  {32'h3fd1a9c8, 32'hc05c7700} /* (3, 16, 16) {real, imag} */,
  {32'h413ffe27, 32'hbfd35518} /* (3, 16, 15) {real, imag} */,
  {32'h40f5b383, 32'hc11ea877} /* (3, 16, 14) {real, imag} */,
  {32'hc0d158ba, 32'h40d528c2} /* (3, 16, 13) {real, imag} */,
  {32'hc139331e, 32'h4081cc74} /* (3, 16, 12) {real, imag} */,
  {32'hc1eeed08, 32'h408856d8} /* (3, 16, 11) {real, imag} */,
  {32'hbf086600, 32'hc0481378} /* (3, 16, 10) {real, imag} */,
  {32'h403f123f, 32'hc007e4d2} /* (3, 16, 9) {real, imag} */,
  {32'h416bbcce, 32'hc1538ad8} /* (3, 16, 8) {real, imag} */,
  {32'hc17075b8, 32'hc0fc8bc4} /* (3, 16, 7) {real, imag} */,
  {32'h402f0676, 32'h4184355a} /* (3, 16, 6) {real, imag} */,
  {32'h40b545aa, 32'h417ac034} /* (3, 16, 5) {real, imag} */,
  {32'hc1e98968, 32'hc21179a6} /* (3, 16, 4) {real, imag} */,
  {32'hc20e4236, 32'h414a1a5d} /* (3, 16, 3) {real, imag} */,
  {32'h419d2c51, 32'hc122a35e} /* (3, 16, 2) {real, imag} */,
  {32'hc0b43ffc, 32'hc1c12f97} /* (3, 16, 1) {real, imag} */,
  {32'h41b74be6, 32'hc23e92b2} /* (3, 16, 0) {real, imag} */,
  {32'hc205c3d2, 32'h419d4324} /* (3, 15, 31) {real, imag} */,
  {32'h428296a8, 32'h41868343} /* (3, 15, 30) {real, imag} */,
  {32'hc1ba49de, 32'h419c4b9f} /* (3, 15, 29) {real, imag} */,
  {32'hc18e27d9, 32'h41061f1e} /* (3, 15, 28) {real, imag} */,
  {32'h401c06c8, 32'h3fcee030} /* (3, 15, 27) {real, imag} */,
  {32'hc1daa758, 32'hc19a75af} /* (3, 15, 26) {real, imag} */,
  {32'hc04aad64, 32'h41cdfab9} /* (3, 15, 25) {real, imag} */,
  {32'hc1a5128c, 32'h4118aa35} /* (3, 15, 24) {real, imag} */,
  {32'h40cda0d1, 32'hc1280d06} /* (3, 15, 23) {real, imag} */,
  {32'hc2376fa4, 32'hc1dac151} /* (3, 15, 22) {real, imag} */,
  {32'h41a4fefc, 32'hc07934d8} /* (3, 15, 21) {real, imag} */,
  {32'hc0aad153, 32'hc173c3ae} /* (3, 15, 20) {real, imag} */,
  {32'hc12112b7, 32'h3fc5ae18} /* (3, 15, 19) {real, imag} */,
  {32'hc03e6330, 32'h41187eea} /* (3, 15, 18) {real, imag} */,
  {32'h40e70ac3, 32'h4077a49f} /* (3, 15, 17) {real, imag} */,
  {32'hc117df17, 32'h40434fa4} /* (3, 15, 16) {real, imag} */,
  {32'h4037888a, 32'hc01b6bef} /* (3, 15, 15) {real, imag} */,
  {32'h3f5cc040, 32'h412472a0} /* (3, 15, 14) {real, imag} */,
  {32'h411581d7, 32'hc11bb4a1} /* (3, 15, 13) {real, imag} */,
  {32'h40d870d1, 32'hbf93ccb4} /* (3, 15, 12) {real, imag} */,
  {32'h3fa28b28, 32'h41f11a5b} /* (3, 15, 11) {real, imag} */,
  {32'hc119e5e2, 32'hc0af48ac} /* (3, 15, 10) {real, imag} */,
  {32'h408459ad, 32'h41965a47} /* (3, 15, 9) {real, imag} */,
  {32'hc189de38, 32'h3fefaa58} /* (3, 15, 8) {real, imag} */,
  {32'hc14f053f, 32'hc14ab3ca} /* (3, 15, 7) {real, imag} */,
  {32'h4193803a, 32'hc02bc7e8} /* (3, 15, 6) {real, imag} */,
  {32'hc21e3a2e, 32'h41d8efd7} /* (3, 15, 5) {real, imag} */,
  {32'hc1370e89, 32'hc1fba4ad} /* (3, 15, 4) {real, imag} */,
  {32'h3f085870, 32'h41c00865} /* (3, 15, 3) {real, imag} */,
  {32'h42cc239c, 32'h41ba47f5} /* (3, 15, 2) {real, imag} */,
  {32'hc21bc6f6, 32'h41e22126} /* (3, 15, 1) {real, imag} */,
  {32'hbf902698, 32'h41600a85} /* (3, 15, 0) {real, imag} */,
  {32'h426bf1d0, 32'h4194f8ff} /* (3, 14, 31) {real, imag} */,
  {32'hc235f922, 32'h41c70217} /* (3, 14, 30) {real, imag} */,
  {32'hc0ccb23c, 32'hc106d499} /* (3, 14, 29) {real, imag} */,
  {32'h418eb679, 32'hc181c231} /* (3, 14, 28) {real, imag} */,
  {32'hc21e942c, 32'h41799248} /* (3, 14, 27) {real, imag} */,
  {32'h4148ac15, 32'hc18adb1e} /* (3, 14, 26) {real, imag} */,
  {32'h41cba67c, 32'h40eee748} /* (3, 14, 25) {real, imag} */,
  {32'h41e07071, 32'h4143ad2d} /* (3, 14, 24) {real, imag} */,
  {32'hc19bf01a, 32'h41b0f807} /* (3, 14, 23) {real, imag} */,
  {32'h41c3de0a, 32'h41063547} /* (3, 14, 22) {real, imag} */,
  {32'hbe1a6660, 32'h41cb4818} /* (3, 14, 21) {real, imag} */,
  {32'h41705754, 32'hbf4ba3f8} /* (3, 14, 20) {real, imag} */,
  {32'hc17edb84, 32'h417b0a23} /* (3, 14, 19) {real, imag} */,
  {32'hbff5a840, 32'hc02a98a7} /* (3, 14, 18) {real, imag} */,
  {32'hc171396e, 32'hc14bd9fe} /* (3, 14, 17) {real, imag} */,
  {32'hc012eb52, 32'hc09798ae} /* (3, 14, 16) {real, imag} */,
  {32'h40924bbc, 32'h4073414e} /* (3, 14, 15) {real, imag} */,
  {32'hc0ca0260, 32'hbfb6cf82} /* (3, 14, 14) {real, imag} */,
  {32'hc180ad16, 32'h411f6a11} /* (3, 14, 13) {real, imag} */,
  {32'h400ace90, 32'hc15e8bea} /* (3, 14, 12) {real, imag} */,
  {32'hc0180bfa, 32'hc14af27c} /* (3, 14, 11) {real, imag} */,
  {32'hbf861578, 32'h41ef5290} /* (3, 14, 10) {real, imag} */,
  {32'h41910ed2, 32'hc0c75538} /* (3, 14, 9) {real, imag} */,
  {32'hc1456db2, 32'h404add64} /* (3, 14, 8) {real, imag} */,
  {32'hc10a7a09, 32'h4227c2cf} /* (3, 14, 7) {real, imag} */,
  {32'hc1376ab7, 32'hc236e5cf} /* (3, 14, 6) {real, imag} */,
  {32'hc251d2d0, 32'hc20810b7} /* (3, 14, 5) {real, imag} */,
  {32'h41ae4b4b, 32'hc225ab92} /* (3, 14, 4) {real, imag} */,
  {32'hc116552a, 32'hc1bd0678} /* (3, 14, 3) {real, imag} */,
  {32'hc28b8a44, 32'h417c47fa} /* (3, 14, 2) {real, imag} */,
  {32'h41b0cf88, 32'h416be52e} /* (3, 14, 1) {real, imag} */,
  {32'h412e4c7e, 32'hc1754f6b} /* (3, 14, 0) {real, imag} */,
  {32'h41331ed4, 32'hc100da8d} /* (3, 13, 31) {real, imag} */,
  {32'hc297a6c2, 32'h4127e60c} /* (3, 13, 30) {real, imag} */,
  {32'hc2023a9c, 32'h3fb8abf8} /* (3, 13, 29) {real, imag} */,
  {32'h4177eac5, 32'hc18f5a0a} /* (3, 13, 28) {real, imag} */,
  {32'h40680950, 32'hc0dc75ec} /* (3, 13, 27) {real, imag} */,
  {32'h425169ec, 32'hc17c86ae} /* (3, 13, 26) {real, imag} */,
  {32'h41d626a3, 32'h41511935} /* (3, 13, 25) {real, imag} */,
  {32'h41c45df1, 32'hc10e4149} /* (3, 13, 24) {real, imag} */,
  {32'hc118861d, 32'h4196ab48} /* (3, 13, 23) {real, imag} */,
  {32'h4124e390, 32'hbfc19058} /* (3, 13, 22) {real, imag} */,
  {32'h418d752f, 32'h40c1b39c} /* (3, 13, 21) {real, imag} */,
  {32'hc162b714, 32'hc132f456} /* (3, 13, 20) {real, imag} */,
  {32'hc176916b, 32'h41a90857} /* (3, 13, 19) {real, imag} */,
  {32'hc09527ea, 32'hc0034e04} /* (3, 13, 18) {real, imag} */,
  {32'h40d5701c, 32'hc10e5495} /* (3, 13, 17) {real, imag} */,
  {32'h40f0db4a, 32'h41310cb4} /* (3, 13, 16) {real, imag} */,
  {32'hc056f0bc, 32'h41596335} /* (3, 13, 15) {real, imag} */,
  {32'h40d9d916, 32'h4053573c} /* (3, 13, 14) {real, imag} */,
  {32'h40ced592, 32'h40e55c5d} /* (3, 13, 13) {real, imag} */,
  {32'hc1afcb6c, 32'hc0c25a14} /* (3, 13, 12) {real, imag} */,
  {32'hc1de2da7, 32'hc1fcc16f} /* (3, 13, 11) {real, imag} */,
  {32'h41c246f8, 32'h414c586f} /* (3, 13, 10) {real, imag} */,
  {32'h40afec92, 32'hc00b10a4} /* (3, 13, 9) {real, imag} */,
  {32'hc156f8d2, 32'hc12c62ff} /* (3, 13, 8) {real, imag} */,
  {32'h41695c86, 32'h419a929e} /* (3, 13, 7) {real, imag} */,
  {32'hc1b7b730, 32'h4238687a} /* (3, 13, 6) {real, imag} */,
  {32'h41bab1ac, 32'hc2304fca} /* (3, 13, 5) {real, imag} */,
  {32'h41a1edb8, 32'h423a414b} /* (3, 13, 4) {real, imag} */,
  {32'hc0b47044, 32'hbfebd670} /* (3, 13, 3) {real, imag} */,
  {32'h428462ae, 32'hc1eebb38} /* (3, 13, 2) {real, imag} */,
  {32'hc16f4dbc, 32'hc1ebe85a} /* (3, 13, 1) {real, imag} */,
  {32'hc1a83052, 32'h4212207f} /* (3, 13, 0) {real, imag} */,
  {32'hbeb512f0, 32'h41dcc26b} /* (3, 12, 31) {real, imag} */,
  {32'h4243148a, 32'hc2035dee} /* (3, 12, 30) {real, imag} */,
  {32'hc22c2f9a, 32'hc1c74696} /* (3, 12, 29) {real, imag} */,
  {32'hc1f1e924, 32'h41ab2e68} /* (3, 12, 28) {real, imag} */,
  {32'hc20d7132, 32'hc268b61a} /* (3, 12, 27) {real, imag} */,
  {32'h3ea43b80, 32'h426dbe92} /* (3, 12, 26) {real, imag} */,
  {32'h40641cf2, 32'hc13e7d90} /* (3, 12, 25) {real, imag} */,
  {32'hc219ee7b, 32'hc1b2fbcb} /* (3, 12, 24) {real, imag} */,
  {32'h411f6c2e, 32'h41a91ce6} /* (3, 12, 23) {real, imag} */,
  {32'hc10740f6, 32'h40eb1c94} /* (3, 12, 22) {real, imag} */,
  {32'h411bdf58, 32'h41a1a365} /* (3, 12, 21) {real, imag} */,
  {32'h415cc6a4, 32'hc10441c0} /* (3, 12, 20) {real, imag} */,
  {32'hc09b78f2, 32'hc213d1be} /* (3, 12, 19) {real, imag} */,
  {32'h40080dba, 32'hc060b44c} /* (3, 12, 18) {real, imag} */,
  {32'h417dedf6, 32'h41cb082a} /* (3, 12, 17) {real, imag} */,
  {32'h410c0ca4, 32'hc15a8026} /* (3, 12, 16) {real, imag} */,
  {32'hc10bf942, 32'hbfcc3a78} /* (3, 12, 15) {real, imag} */,
  {32'h410b398a, 32'h3c752400} /* (3, 12, 14) {real, imag} */,
  {32'h4003612c, 32'h41469a32} /* (3, 12, 13) {real, imag} */,
  {32'h40228de0, 32'h4238334c} /* (3, 12, 12) {real, imag} */,
  {32'hc0ee0060, 32'h417f0772} /* (3, 12, 11) {real, imag} */,
  {32'h419981ef, 32'hc14a317e} /* (3, 12, 10) {real, imag} */,
  {32'h4023c2ce, 32'h41c6adc6} /* (3, 12, 9) {real, imag} */,
  {32'hc1c703ae, 32'hc1bad1b5} /* (3, 12, 8) {real, imag} */,
  {32'h4190e3af, 32'hc231611e} /* (3, 12, 7) {real, imag} */,
  {32'h3fbd9838, 32'h3f64c720} /* (3, 12, 6) {real, imag} */,
  {32'hc286917c, 32'h421f8de0} /* (3, 12, 5) {real, imag} */,
  {32'h42c8eef3, 32'h404de800} /* (3, 12, 4) {real, imag} */,
  {32'h40120fa8, 32'hc235a489} /* (3, 12, 3) {real, imag} */,
  {32'h41e83531, 32'hc0338438} /* (3, 12, 2) {real, imag} */,
  {32'h41396734, 32'hc25e7596} /* (3, 12, 1) {real, imag} */,
  {32'h40b96967, 32'h411d3bc8} /* (3, 12, 0) {real, imag} */,
  {32'h42fa12d6, 32'hc12b5500} /* (3, 11, 31) {real, imag} */,
  {32'hc24e8c76, 32'h424334b3} /* (3, 11, 30) {real, imag} */,
  {32'hc23bf26b, 32'h42a4e481} /* (3, 11, 29) {real, imag} */,
  {32'hc2150224, 32'hc155491c} /* (3, 11, 28) {real, imag} */,
  {32'hc15761bf, 32'h40a98410} /* (3, 11, 27) {real, imag} */,
  {32'hc24097d4, 32'hc1958af6} /* (3, 11, 26) {real, imag} */,
  {32'hc2a63933, 32'h416a0c95} /* (3, 11, 25) {real, imag} */,
  {32'hc12fec94, 32'hc267af67} /* (3, 11, 24) {real, imag} */,
  {32'hc0a4fc58, 32'hc1ffaeca} /* (3, 11, 23) {real, imag} */,
  {32'hc0b834b4, 32'hc21c5c4b} /* (3, 11, 22) {real, imag} */,
  {32'h42653e83, 32'h41701b66} /* (3, 11, 21) {real, imag} */,
  {32'h40cfb02c, 32'h40cf08c6} /* (3, 11, 20) {real, imag} */,
  {32'hbf3f9810, 32'h4142a686} /* (3, 11, 19) {real, imag} */,
  {32'h41dedd20, 32'h41f0a776} /* (3, 11, 18) {real, imag} */,
  {32'hbf4bcce0, 32'hbfa80d74} /* (3, 11, 17) {real, imag} */,
  {32'hbf903880, 32'hbfbcc784} /* (3, 11, 16) {real, imag} */,
  {32'hc11ad89a, 32'hc0effd99} /* (3, 11, 15) {real, imag} */,
  {32'h40546434, 32'hc1a272ce} /* (3, 11, 14) {real, imag} */,
  {32'h419881f2, 32'hc1ad29dd} /* (3, 11, 13) {real, imag} */,
  {32'hc15f32b2, 32'h3fb9fb48} /* (3, 11, 12) {real, imag} */,
  {32'hc21ac305, 32'hc089e864} /* (3, 11, 11) {real, imag} */,
  {32'hc21df5aa, 32'h420c093f} /* (3, 11, 10) {real, imag} */,
  {32'hc15c4fe4, 32'hc18f7b70} /* (3, 11, 9) {real, imag} */,
  {32'hc0639286, 32'hc1a6c752} /* (3, 11, 8) {real, imag} */,
  {32'h42856eb1, 32'h41e8ee68} /* (3, 11, 7) {real, imag} */,
  {32'hc19d6f14, 32'hc270f351} /* (3, 11, 6) {real, imag} */,
  {32'hc08fab06, 32'h41dc678a} /* (3, 11, 5) {real, imag} */,
  {32'h41c8cf8c, 32'hc24da9f9} /* (3, 11, 4) {real, imag} */,
  {32'h41e6e7ba, 32'hc1ae5c0b} /* (3, 11, 3) {real, imag} */,
  {32'hc2d5d38d, 32'h41b33722} /* (3, 11, 2) {real, imag} */,
  {32'h42cd8756, 32'h4225e6c8} /* (3, 11, 1) {real, imag} */,
  {32'h4211b222, 32'hc171d7c0} /* (3, 11, 0) {real, imag} */,
  {32'hc06ffc70, 32'h417452f9} /* (3, 10, 31) {real, imag} */,
  {32'h42a544ce, 32'h429ceb6a} /* (3, 10, 30) {real, imag} */,
  {32'hc1fd9537, 32'h4196a8f3} /* (3, 10, 29) {real, imag} */,
  {32'hc1977f49, 32'h41b37f46} /* (3, 10, 28) {real, imag} */,
  {32'h41d927f0, 32'h41d0c061} /* (3, 10, 27) {real, imag} */,
  {32'hc18a8b13, 32'hc0cfc7b0} /* (3, 10, 26) {real, imag} */,
  {32'h40eeecce, 32'hbfd13bd0} /* (3, 10, 25) {real, imag} */,
  {32'h42e001b1, 32'h41103712} /* (3, 10, 24) {real, imag} */,
  {32'hc1ab540c, 32'hc286bf25} /* (3, 10, 23) {real, imag} */,
  {32'h420c61c8, 32'hc22c5cf8} /* (3, 10, 22) {real, imag} */,
  {32'hc244b1c8, 32'h426334c8} /* (3, 10, 21) {real, imag} */,
  {32'h40667548, 32'h4255fb72} /* (3, 10, 20) {real, imag} */,
  {32'hc1953b51, 32'hc17005ee} /* (3, 10, 19) {real, imag} */,
  {32'h4092b83a, 32'h4087bc42} /* (3, 10, 18) {real, imag} */,
  {32'hc14707f6, 32'hc10c7012} /* (3, 10, 17) {real, imag} */,
  {32'h40e29554, 32'hc130e058} /* (3, 10, 16) {real, imag} */,
  {32'h41b2c20f, 32'h41456150} /* (3, 10, 15) {real, imag} */,
  {32'hc12ebe65, 32'hc0a2c992} /* (3, 10, 14) {real, imag} */,
  {32'hc1025e0a, 32'h421b5d9a} /* (3, 10, 13) {real, imag} */,
  {32'hc1eec019, 32'h3fc6f190} /* (3, 10, 12) {real, imag} */,
  {32'hbf0cf880, 32'hc141f05e} /* (3, 10, 11) {real, imag} */,
  {32'hc1bad715, 32'hc22013f4} /* (3, 10, 10) {real, imag} */,
  {32'h4194554e, 32'hc149a738} /* (3, 10, 9) {real, imag} */,
  {32'hc251cbbe, 32'hc016e708} /* (3, 10, 8) {real, imag} */,
  {32'h4166134f, 32'hc21f5bae} /* (3, 10, 7) {real, imag} */,
  {32'h42083e74, 32'hc2dd4fa1} /* (3, 10, 6) {real, imag} */,
  {32'h4180d284, 32'hc2a307a4} /* (3, 10, 5) {real, imag} */,
  {32'h3f83c350, 32'h4048e4fc} /* (3, 10, 4) {real, imag} */,
  {32'h42a6c17b, 32'hc2529d9c} /* (3, 10, 3) {real, imag} */,
  {32'h429f5756, 32'h427b698b} /* (3, 10, 2) {real, imag} */,
  {32'hc2d3e324, 32'h41897a88} /* (3, 10, 1) {real, imag} */,
  {32'hc287fa7f, 32'hc33ea4c6} /* (3, 10, 0) {real, imag} */,
  {32'hc27795e8, 32'hc2ed6d13} /* (3, 9, 31) {real, imag} */,
  {32'h42a7e9ab, 32'h41b47d80} /* (3, 9, 30) {real, imag} */,
  {32'hc3087acc, 32'h4226fbfa} /* (3, 9, 29) {real, imag} */,
  {32'h4238b899, 32'hc31aa75f} /* (3, 9, 28) {real, imag} */,
  {32'h42a4cbc4, 32'hc29d598e} /* (3, 9, 27) {real, imag} */,
  {32'hc1e75c84, 32'hc2a3f96a} /* (3, 9, 26) {real, imag} */,
  {32'hc254eafd, 32'hc1528f79} /* (3, 9, 25) {real, imag} */,
  {32'hc15bbcbc, 32'h41844f28} /* (3, 9, 24) {real, imag} */,
  {32'h41ad8804, 32'hc1d3a513} /* (3, 9, 23) {real, imag} */,
  {32'h41d9940a, 32'h420d2a07} /* (3, 9, 22) {real, imag} */,
  {32'hc1d3e2b4, 32'h4205e877} /* (3, 9, 21) {real, imag} */,
  {32'h41456739, 32'hc2181171} /* (3, 9, 20) {real, imag} */,
  {32'hc1853528, 32'hc26465c2} /* (3, 9, 19) {real, imag} */,
  {32'h41cd9e79, 32'h4123f46c} /* (3, 9, 18) {real, imag} */,
  {32'hc1121583, 32'hbf49c540} /* (3, 9, 17) {real, imag} */,
  {32'hc0dde594, 32'h40d32aec} /* (3, 9, 16) {real, imag} */,
  {32'hc073f594, 32'h4097f1d8} /* (3, 9, 15) {real, imag} */,
  {32'hc1b41663, 32'hc0c85a80} /* (3, 9, 14) {real, imag} */,
  {32'hc1b03020, 32'hc16ef376} /* (3, 9, 13) {real, imag} */,
  {32'h412f173d, 32'hc0d687b8} /* (3, 9, 12) {real, imag} */,
  {32'h41c46804, 32'h4103f459} /* (3, 9, 11) {real, imag} */,
  {32'h4205812a, 32'h4243e931} /* (3, 9, 10) {real, imag} */,
  {32'h410a7659, 32'hc222197c} /* (3, 9, 9) {real, imag} */,
  {32'h411f3d84, 32'h41ede882} /* (3, 9, 8) {real, imag} */,
  {32'h421173f5, 32'hc165eae5} /* (3, 9, 7) {real, imag} */,
  {32'hc24603f8, 32'hc20e3438} /* (3, 9, 6) {real, imag} */,
  {32'hc2ddd7c6, 32'hc2154068} /* (3, 9, 5) {real, imag} */,
  {32'hc19bf0e6, 32'h425ecc94} /* (3, 9, 4) {real, imag} */,
  {32'h41b84d18, 32'hc23e9d6e} /* (3, 9, 3) {real, imag} */,
  {32'hc2665a42, 32'hc181fe32} /* (3, 9, 2) {real, imag} */,
  {32'hc1a28894, 32'h433f06c8} /* (3, 9, 1) {real, imag} */,
  {32'h4234a610, 32'hc20ac6de} /* (3, 9, 0) {real, imag} */,
  {32'h42cf3762, 32'hc322f266} /* (3, 8, 31) {real, imag} */,
  {32'hc0105558, 32'h43124676} /* (3, 8, 30) {real, imag} */,
  {32'hc233f0ed, 32'hc2289476} /* (3, 8, 29) {real, imag} */,
  {32'hc1bce2d3, 32'h42019e9e} /* (3, 8, 28) {real, imag} */,
  {32'hc10c9246, 32'hc187d8fe} /* (3, 8, 27) {real, imag} */,
  {32'h42ca45dd, 32'hc1da6bbc} /* (3, 8, 26) {real, imag} */,
  {32'h42e48f04, 32'hc24fa266} /* (3, 8, 25) {real, imag} */,
  {32'h41fe9020, 32'hc179c12c} /* (3, 8, 24) {real, imag} */,
  {32'h41f6db09, 32'h3f2d2460} /* (3, 8, 23) {real, imag} */,
  {32'hc0c157d4, 32'h4211af98} /* (3, 8, 22) {real, imag} */,
  {32'hc2306cc4, 32'hc1e50fca} /* (3, 8, 21) {real, imag} */,
  {32'hc0d10834, 32'h40d67b40} /* (3, 8, 20) {real, imag} */,
  {32'h41eab061, 32'h4139719c} /* (3, 8, 19) {real, imag} */,
  {32'h413f6402, 32'hc14bce21} /* (3, 8, 18) {real, imag} */,
  {32'h4081045e, 32'hc1d57d22} /* (3, 8, 17) {real, imag} */,
  {32'hc1972066, 32'h3ffe8b00} /* (3, 8, 16) {real, imag} */,
  {32'h4003f905, 32'hc12c3c2c} /* (3, 8, 15) {real, imag} */,
  {32'h403d8e10, 32'hc12b3e47} /* (3, 8, 14) {real, imag} */,
  {32'hc1dc8429, 32'h402f686e} /* (3, 8, 13) {real, imag} */,
  {32'h4199747c, 32'hc1b9a9c0} /* (3, 8, 12) {real, imag} */,
  {32'hc2b4911c, 32'hc288fe0c} /* (3, 8, 11) {real, imag} */,
  {32'hc0df400c, 32'h42ca7580} /* (3, 8, 10) {real, imag} */,
  {32'h41af1869, 32'hc26d7f2e} /* (3, 8, 9) {real, imag} */,
  {32'hc2e1ea56, 32'hc1ba126a} /* (3, 8, 8) {real, imag} */,
  {32'hc2a9ebe8, 32'hc139d652} /* (3, 8, 7) {real, imag} */,
  {32'h3fca9440, 32'h423b81b2} /* (3, 8, 6) {real, imag} */,
  {32'hc1954455, 32'hc294b6ba} /* (3, 8, 5) {real, imag} */,
  {32'h420619a0, 32'h42e4b3a3} /* (3, 8, 4) {real, imag} */,
  {32'hc2f808f4, 32'hc2a44dbc} /* (3, 8, 3) {real, imag} */,
  {32'hc1af1fa2, 32'h42be3ce8} /* (3, 8, 2) {real, imag} */,
  {32'h42e7b9a8, 32'hc1132ad8} /* (3, 8, 1) {real, imag} */,
  {32'h4295147a, 32'hc2ea27f6} /* (3, 8, 0) {real, imag} */,
  {32'h423076bc, 32'hc232ca43} /* (3, 7, 31) {real, imag} */,
  {32'h3fed8a60, 32'hc03b2208} /* (3, 7, 30) {real, imag} */,
  {32'h41deff9a, 32'h427546aa} /* (3, 7, 29) {real, imag} */,
  {32'h42856c24, 32'h42b1b920} /* (3, 7, 28) {real, imag} */,
  {32'h4182bcda, 32'hc1fed316} /* (3, 7, 27) {real, imag} */,
  {32'h41681952, 32'h42caecca} /* (3, 7, 26) {real, imag} */,
  {32'h422f0cc8, 32'hc200c0b2} /* (3, 7, 25) {real, imag} */,
  {32'hc2050816, 32'h41cf8699} /* (3, 7, 24) {real, imag} */,
  {32'h40c2a9a8, 32'hc233d7a6} /* (3, 7, 23) {real, imag} */,
  {32'hc229c60e, 32'h3e0be000} /* (3, 7, 22) {real, imag} */,
  {32'hc24061f4, 32'h409a3a4a} /* (3, 7, 21) {real, imag} */,
  {32'hc242e009, 32'hc1f10370} /* (3, 7, 20) {real, imag} */,
  {32'h41ae2193, 32'h42880cb5} /* (3, 7, 19) {real, imag} */,
  {32'h4129e350, 32'h424a54da} /* (3, 7, 18) {real, imag} */,
  {32'h41fa1d60, 32'hc181b31e} /* (3, 7, 17) {real, imag} */,
  {32'h408d7c2a, 32'h413217b8} /* (3, 7, 16) {real, imag} */,
  {32'h420bd6d2, 32'h400b0c24} /* (3, 7, 15) {real, imag} */,
  {32'hc2100f70, 32'h4106978a} /* (3, 7, 14) {real, imag} */,
  {32'h42145ac8, 32'hc1257040} /* (3, 7, 13) {real, imag} */,
  {32'h41a59d9e, 32'hc0f521c2} /* (3, 7, 12) {real, imag} */,
  {32'hc13af7e6, 32'h41b63460} /* (3, 7, 11) {real, imag} */,
  {32'h42d30b97, 32'h41bf68be} /* (3, 7, 10) {real, imag} */,
  {32'hc2803f6e, 32'hbf030f60} /* (3, 7, 9) {real, imag} */,
  {32'h417e47f8, 32'hc1d88c33} /* (3, 7, 8) {real, imag} */,
  {32'hc2262d40, 32'hc1e06cf5} /* (3, 7, 7) {real, imag} */,
  {32'h41a91c79, 32'h41e92690} /* (3, 7, 6) {real, imag} */,
  {32'h42bfc94c, 32'h429479b0} /* (3, 7, 5) {real, imag} */,
  {32'hc2da0f3e, 32'h42bba650} /* (3, 7, 4) {real, imag} */,
  {32'h42ade4d2, 32'h421fbdd8} /* (3, 7, 3) {real, imag} */,
  {32'h428712e4, 32'hc23f3df0} /* (3, 7, 2) {real, imag} */,
  {32'hc0e8fd34, 32'h4207fff5} /* (3, 7, 1) {real, imag} */,
  {32'h418387a8, 32'h42eb6a65} /* (3, 7, 0) {real, imag} */,
  {32'hc29e4cf5, 32'hc286638e} /* (3, 6, 31) {real, imag} */,
  {32'h423c4596, 32'hc29bf081} /* (3, 6, 30) {real, imag} */,
  {32'hc1a02d23, 32'hc1374dde} /* (3, 6, 29) {real, imag} */,
  {32'hc0a660d4, 32'hc1e978d7} /* (3, 6, 28) {real, imag} */,
  {32'h42029042, 32'hc2fd7113} /* (3, 6, 27) {real, imag} */,
  {32'h428d53ff, 32'h42e6ffca} /* (3, 6, 26) {real, imag} */,
  {32'hc29a75da, 32'hc224d705} /* (3, 6, 25) {real, imag} */,
  {32'h408d6e9c, 32'hc178f8e8} /* (3, 6, 24) {real, imag} */,
  {32'hc001a938, 32'h4325ee80} /* (3, 6, 23) {real, imag} */,
  {32'h414e4240, 32'hc2a5b3d6} /* (3, 6, 22) {real, imag} */,
  {32'h41bdaebc, 32'h41c4bbce} /* (3, 6, 21) {real, imag} */,
  {32'h4252bbe4, 32'hc1c50423} /* (3, 6, 20) {real, imag} */,
  {32'h4229b7dc, 32'h4189972f} /* (3, 6, 19) {real, imag} */,
  {32'hc248af90, 32'h41767674} /* (3, 6, 18) {real, imag} */,
  {32'h41605295, 32'hc1ae6192} /* (3, 6, 17) {real, imag} */,
  {32'hc1ead7be, 32'hc189763a} /* (3, 6, 16) {real, imag} */,
  {32'hc15ba5e5, 32'hc1f70bee} /* (3, 6, 15) {real, imag} */,
  {32'h4136db84, 32'hc055d9d0} /* (3, 6, 14) {real, imag} */,
  {32'hc1bb5419, 32'h411315fa} /* (3, 6, 13) {real, imag} */,
  {32'hc28946a7, 32'h41b56639} /* (3, 6, 12) {real, imag} */,
  {32'hc1bd3dc2, 32'h41b17498} /* (3, 6, 11) {real, imag} */,
  {32'hc18fca36, 32'hc2030b17} /* (3, 6, 10) {real, imag} */,
  {32'hc1b46039, 32'hc09d0640} /* (3, 6, 9) {real, imag} */,
  {32'h42037188, 32'hc26a7fcc} /* (3, 6, 8) {real, imag} */,
  {32'hc350e1a3, 32'h42ee1f9e} /* (3, 6, 7) {real, imag} */,
  {32'hc28d582f, 32'h41d92ee2} /* (3, 6, 6) {real, imag} */,
  {32'hc25a6d3e, 32'hc0aed530} /* (3, 6, 5) {real, imag} */,
  {32'hc1fd37b9, 32'h414c6382} /* (3, 6, 4) {real, imag} */,
  {32'h42a00ccf, 32'hc1da2589} /* (3, 6, 3) {real, imag} */,
  {32'h423434a6, 32'hc320df64} /* (3, 6, 2) {real, imag} */,
  {32'hc08bc390, 32'hc308a489} /* (3, 6, 1) {real, imag} */,
  {32'h422f9e37, 32'h42b04e70} /* (3, 6, 0) {real, imag} */,
  {32'h4306491a, 32'hc3eace32} /* (3, 5, 31) {real, imag} */,
  {32'hc294e3e9, 32'h43652a78} /* (3, 5, 30) {real, imag} */,
  {32'hc16a5314, 32'h42f876e0} /* (3, 5, 29) {real, imag} */,
  {32'h41871689, 32'hc25cf160} /* (3, 5, 28) {real, imag} */,
  {32'hc21f8ef4, 32'h4335da33} /* (3, 5, 27) {real, imag} */,
  {32'hc2af94e0, 32'hc2288bce} /* (3, 5, 26) {real, imag} */,
  {32'hc31764a0, 32'hc252af56} /* (3, 5, 25) {real, imag} */,
  {32'h42c3d770, 32'hc2909d12} /* (3, 5, 24) {real, imag} */,
  {32'h4221601f, 32'hc1d69cbb} /* (3, 5, 23) {real, imag} */,
  {32'hc21e19a6, 32'hc0b0a254} /* (3, 5, 22) {real, imag} */,
  {32'h421624b0, 32'h421a92bd} /* (3, 5, 21) {real, imag} */,
  {32'h4213a2d3, 32'hc18206e4} /* (3, 5, 20) {real, imag} */,
  {32'h427bd61b, 32'hc0cdde00} /* (3, 5, 19) {real, imag} */,
  {32'hc1f29a8d, 32'h41c3e0b8} /* (3, 5, 18) {real, imag} */,
  {32'hbf81fb40, 32'h41afa890} /* (3, 5, 17) {real, imag} */,
  {32'hc18bc1c4, 32'h42529c88} /* (3, 5, 16) {real, imag} */,
  {32'hc1329818, 32'h410828a0} /* (3, 5, 15) {real, imag} */,
  {32'hc23b65da, 32'hc06dce04} /* (3, 5, 14) {real, imag} */,
  {32'h40b65128, 32'hc032d840} /* (3, 5, 13) {real, imag} */,
  {32'h41e7aa32, 32'h424fdc4c} /* (3, 5, 12) {real, imag} */,
  {32'h410b4320, 32'hc2609603} /* (3, 5, 11) {real, imag} */,
  {32'hc2664c4e, 32'h42733bba} /* (3, 5, 10) {real, imag} */,
  {32'h428ad328, 32'h424e2b04} /* (3, 5, 9) {real, imag} */,
  {32'hc2085e88, 32'h4271071b} /* (3, 5, 8) {real, imag} */,
  {32'h42f039ec, 32'h414ec69e} /* (3, 5, 7) {real, imag} */,
  {32'h42239d58, 32'h4294977b} /* (3, 5, 6) {real, imag} */,
  {32'hc32e4aa7, 32'hc2dc03ee} /* (3, 5, 5) {real, imag} */,
  {32'hc1cc8edb, 32'hc201246a} /* (3, 5, 4) {real, imag} */,
  {32'hc2bafe02, 32'hc1a51018} /* (3, 5, 3) {real, imag} */,
  {32'hc1f7e393, 32'h431ea27c} /* (3, 5, 2) {real, imag} */,
  {32'h43d2f20f, 32'hc3268130} /* (3, 5, 1) {real, imag} */,
  {32'h430edccc, 32'hc3705470} /* (3, 5, 0) {real, imag} */,
  {32'hc396a54a, 32'h43319041} /* (3, 4, 31) {real, imag} */,
  {32'h43803921, 32'hc34ba7fc} /* (3, 4, 30) {real, imag} */,
  {32'hc2c27495, 32'h4208deef} /* (3, 4, 29) {real, imag} */,
  {32'hbf9838c0, 32'h42f03fbf} /* (3, 4, 28) {real, imag} */,
  {32'h40ebaf40, 32'hc32cc5a6} /* (3, 4, 27) {real, imag} */,
  {32'hc21004c2, 32'hc2e1b6cb} /* (3, 4, 26) {real, imag} */,
  {32'h4295983a, 32'hc235f9b4} /* (3, 4, 25) {real, imag} */,
  {32'h427166da, 32'hc17c37c0} /* (3, 4, 24) {real, imag} */,
  {32'hc05011c0, 32'hc22848f2} /* (3, 4, 23) {real, imag} */,
  {32'hc2248982, 32'h4264840d} /* (3, 4, 22) {real, imag} */,
  {32'hc1ba3ca0, 32'hc24b4d88} /* (3, 4, 21) {real, imag} */,
  {32'h41c5716a, 32'h42060a1b} /* (3, 4, 20) {real, imag} */,
  {32'h409acb20, 32'h4181f396} /* (3, 4, 19) {real, imag} */,
  {32'h4142c1d4, 32'hc18c8040} /* (3, 4, 18) {real, imag} */,
  {32'h41894563, 32'h41a377c6} /* (3, 4, 17) {real, imag} */,
  {32'h4076f4a0, 32'h3ff64100} /* (3, 4, 16) {real, imag} */,
  {32'h415c511a, 32'hc25ca3e3} /* (3, 4, 15) {real, imag} */,
  {32'h423607bb, 32'hc1e93018} /* (3, 4, 14) {real, imag} */,
  {32'h415b9b70, 32'hc11d67b4} /* (3, 4, 13) {real, imag} */,
  {32'hbf5cf840, 32'hc1c08c5e} /* (3, 4, 12) {real, imag} */,
  {32'h42583bbc, 32'h42087adc} /* (3, 4, 11) {real, imag} */,
  {32'hc2a2b46d, 32'h41b98a3e} /* (3, 4, 10) {real, imag} */,
  {32'h429d16a2, 32'hc169d1fe} /* (3, 4, 9) {real, imag} */,
  {32'h42a1d7cd, 32'hc2ba1026} /* (3, 4, 8) {real, imag} */,
  {32'h42bad0a2, 32'hbfa167d0} /* (3, 4, 7) {real, imag} */,
  {32'hc04da6a0, 32'h428fc411} /* (3, 4, 6) {real, imag} */,
  {32'h43202c9e, 32'hc215bdda} /* (3, 4, 5) {real, imag} */,
  {32'hc35ca69c, 32'h42ff1557} /* (3, 4, 4) {real, imag} */,
  {32'h4301aa1c, 32'hc288865a} /* (3, 4, 3) {real, imag} */,
  {32'h43b6d26d, 32'hc31d9ee4} /* (3, 4, 2) {real, imag} */,
  {32'hc3739e1b, 32'h4398bea1} /* (3, 4, 1) {real, imag} */,
  {32'hc2962749, 32'h43c7cf61} /* (3, 4, 0) {real, imag} */,
  {32'hc26fe028, 32'hc39a68c2} /* (3, 3, 31) {real, imag} */,
  {32'h418c6614, 32'h43244571} /* (3, 3, 30) {real, imag} */,
  {32'hc0c1033c, 32'hc0ead730} /* (3, 3, 29) {real, imag} */,
  {32'hc2b75bd8, 32'h40dc1cc0} /* (3, 3, 28) {real, imag} */,
  {32'h429910a4, 32'hc24c3bd0} /* (3, 3, 27) {real, imag} */,
  {32'h431681a7, 32'h3f12b5c0} /* (3, 3, 26) {real, imag} */,
  {32'hc280eaf8, 32'hc339c366} /* (3, 3, 25) {real, imag} */,
  {32'h438ed91b, 32'h4248351e} /* (3, 3, 24) {real, imag} */,
  {32'hc2e99b35, 32'h41987b9d} /* (3, 3, 23) {real, imag} */,
  {32'hc2269809, 32'hc2823fdf} /* (3, 3, 22) {real, imag} */,
  {32'h40d198ec, 32'hc0af4acc} /* (3, 3, 21) {real, imag} */,
  {32'h41e5fa20, 32'h417d17ec} /* (3, 3, 20) {real, imag} */,
  {32'hc2dfa02b, 32'h41951d61} /* (3, 3, 19) {real, imag} */,
  {32'h425b19ea, 32'h41bee993} /* (3, 3, 18) {real, imag} */,
  {32'h4249aeb8, 32'h41d495b8} /* (3, 3, 17) {real, imag} */,
  {32'h424e0df4, 32'hc214de02} /* (3, 3, 16) {real, imag} */,
  {32'hc21fb1be, 32'hc190bba0} /* (3, 3, 15) {real, imag} */,
  {32'h4131e518, 32'hc201cb2e} /* (3, 3, 14) {real, imag} */,
  {32'h41a80afc, 32'h42155288} /* (3, 3, 13) {real, imag} */,
  {32'h426be6b6, 32'h42753fc5} /* (3, 3, 12) {real, imag} */,
  {32'h40a12cec, 32'h4248b006} /* (3, 3, 11) {real, imag} */,
  {32'h4269b175, 32'h4231e282} /* (3, 3, 10) {real, imag} */,
  {32'hc2e8a09f, 32'hc0f6d5f4} /* (3, 3, 9) {real, imag} */,
  {32'h4151bf80, 32'h42906aff} /* (3, 3, 8) {real, imag} */,
  {32'hc2d79894, 32'hc287ec15} /* (3, 3, 7) {real, imag} */,
  {32'h42f12712, 32'h4277e2be} /* (3, 3, 6) {real, imag} */,
  {32'hc27635fc, 32'h431150e8} /* (3, 3, 5) {real, imag} */,
  {32'hc2b4845c, 32'hc38e6b02} /* (3, 3, 4) {real, imag} */,
  {32'hc20bbf00, 32'h430e3076} /* (3, 3, 3) {real, imag} */,
  {32'h4348cdb4, 32'h4342bc9b} /* (3, 3, 2) {real, imag} */,
  {32'hc34535c4, 32'h421a0770} /* (3, 3, 1) {real, imag} */,
  {32'hc22ca1ac, 32'hc33e3ef8} /* (3, 3, 0) {real, imag} */,
  {32'h43f1cfbd, 32'hc4a748c3} /* (3, 2, 31) {real, imag} */,
  {32'hc2fe8570, 32'h445151ab} /* (3, 2, 30) {real, imag} */,
  {32'h411cc4d8, 32'hc2f3afae} /* (3, 2, 29) {real, imag} */,
  {32'hc35ca5ea, 32'hc2b56009} /* (3, 2, 28) {real, imag} */,
  {32'h42f3d155, 32'h43565b26} /* (3, 2, 27) {real, imag} */,
  {32'h4232621e, 32'h4238be28} /* (3, 2, 26) {real, imag} */,
  {32'h4117a2e4, 32'h4079e800} /* (3, 2, 25) {real, imag} */,
  {32'h4256f266, 32'h43216a1a} /* (3, 2, 24) {real, imag} */,
  {32'hc275f065, 32'h425e5328} /* (3, 2, 23) {real, imag} */,
  {32'hc314726c, 32'hc1982ca4} /* (3, 2, 22) {real, imag} */,
  {32'h42881bb5, 32'hc2862667} /* (3, 2, 21) {real, imag} */,
  {32'hc1bc2c1b, 32'h42693b0e} /* (3, 2, 20) {real, imag} */,
  {32'h425e6a05, 32'h4196e3ed} /* (3, 2, 19) {real, imag} */,
  {32'h4132b4b0, 32'hc1478200} /* (3, 2, 18) {real, imag} */,
  {32'hc201c7b6, 32'hc0f61460} /* (3, 2, 17) {real, imag} */,
  {32'h3f724500, 32'h421c49ac} /* (3, 2, 16) {real, imag} */,
  {32'hbff716c0, 32'hc21abf14} /* (3, 2, 15) {real, imag} */,
  {32'hc03c48a0, 32'hc1aa31c0} /* (3, 2, 14) {real, imag} */,
  {32'hc068e3f0, 32'h417b29b6} /* (3, 2, 13) {real, imag} */,
  {32'h42726f92, 32'hc2423112} /* (3, 2, 12) {real, imag} */,
  {32'hc2364a56, 32'h4192abd4} /* (3, 2, 11) {real, imag} */,
  {32'h42836c33, 32'hc27597c8} /* (3, 2, 10) {real, imag} */,
  {32'hc290b252, 32'h41e40b90} /* (3, 2, 9) {real, imag} */,
  {32'hc0d1b190, 32'hbffe5240} /* (3, 2, 8) {real, imag} */,
  {32'h42bb17dc, 32'hc23e1ef0} /* (3, 2, 7) {real, imag} */,
  {32'h417f00da, 32'hc2028cfe} /* (3, 2, 6) {real, imag} */,
  {32'hc2cd7983, 32'h4331b72a} /* (3, 2, 5) {real, imag} */,
  {32'h4323a17e, 32'hc309011a} /* (3, 2, 4) {real, imag} */,
  {32'hc294d17f, 32'hc29d4716} /* (3, 2, 3) {real, imag} */,
  {32'hc11aed1c, 32'h440fadbf} /* (3, 2, 2) {real, imag} */,
  {32'h3fbed500, 32'hc4269688} /* (3, 2, 1) {real, imag} */,
  {32'h4393e7b0, 32'hc3da52de} /* (3, 2, 0) {real, imag} */,
  {32'hc2e9c6c8, 32'h449561f5} /* (3, 1, 31) {real, imag} */,
  {32'h435cca18, 32'hc39c594f} /* (3, 1, 30) {real, imag} */,
  {32'hc27a1988, 32'hc375788c} /* (3, 1, 29) {real, imag} */,
  {32'hc38630c0, 32'h4386405f} /* (3, 1, 28) {real, imag} */,
  {32'h4317f194, 32'hc3d51bf3} /* (3, 1, 27) {real, imag} */,
  {32'hc20418dc, 32'hc2a38482} /* (3, 1, 26) {real, imag} */,
  {32'h4343b622, 32'h4246308e} /* (3, 1, 25) {real, imag} */,
  {32'hc2ad06e4, 32'hc3227cf8} /* (3, 1, 24) {real, imag} */,
  {32'h421398f6, 32'hc1d6e6bc} /* (3, 1, 23) {real, imag} */,
  {32'h4260c774, 32'h428d70ef} /* (3, 1, 22) {real, imag} */,
  {32'hc14fa2b0, 32'hc2cd8983} /* (3, 1, 21) {real, imag} */,
  {32'hc24d66e1, 32'h4253515c} /* (3, 1, 20) {real, imag} */,
  {32'hc24cd8fc, 32'h412a8b44} /* (3, 1, 19) {real, imag} */,
  {32'hc2904f90, 32'hc0b4e5d8} /* (3, 1, 18) {real, imag} */,
  {32'hc1966280, 32'hc20fadfc} /* (3, 1, 17) {real, imag} */,
  {32'h4232219c, 32'h41efc280} /* (3, 1, 16) {real, imag} */,
  {32'hc0c5df00, 32'hc20106c4} /* (3, 1, 15) {real, imag} */,
  {32'h4203b3a8, 32'h4276ad63} /* (3, 1, 14) {real, imag} */,
  {32'hc2decf02, 32'hc20c1d73} /* (3, 1, 13) {real, imag} */,
  {32'h420290c7, 32'h420fa2c4} /* (3, 1, 12) {real, imag} */,
  {32'h430c5e51, 32'hc1d67054} /* (3, 1, 11) {real, imag} */,
  {32'hc22eff9c, 32'hc312eb82} /* (3, 1, 10) {real, imag} */,
  {32'h4311f08c, 32'h4185475c} /* (3, 1, 9) {real, imag} */,
  {32'h4327304c, 32'hc16b47f8} /* (3, 1, 8) {real, imag} */,
  {32'hc2b4bb4c, 32'hc31d7d20} /* (3, 1, 7) {real, imag} */,
  {32'hc30eebc3, 32'hc2ca7150} /* (3, 1, 6) {real, imag} */,
  {32'h4335198a, 32'hc3905df3} /* (3, 1, 5) {real, imag} */,
  {32'h41c73958, 32'h431cecfa} /* (3, 1, 4) {real, imag} */,
  {32'h437c33fa, 32'h42ecd2e0} /* (3, 1, 3) {real, imag} */,
  {32'h443d8d10, 32'hc3f3f585} /* (3, 1, 2) {real, imag} */,
  {32'hc490dbee, 32'h449f9f39} /* (3, 1, 1) {real, imag} */,
  {32'hc3b9ef3e, 32'h446e4f86} /* (3, 1, 0) {real, imag} */,
  {32'h43ea177a, 32'h442cf7a2} /* (3, 0, 31) {real, imag} */,
  {32'hc364a3a4, 32'hc3612c2f} /* (3, 0, 30) {real, imag} */,
  {32'hc33eb7a6, 32'hc1e8afc0} /* (3, 0, 29) {real, imag} */,
  {32'hc37d26c0, 32'hc1919b99} /* (3, 0, 28) {real, imag} */,
  {32'h42bb0b1e, 32'hc38131fd} /* (3, 0, 27) {real, imag} */,
  {32'hc2cfc59c, 32'hc277bc00} /* (3, 0, 26) {real, imag} */,
  {32'h42da2024, 32'h428ea669} /* (3, 0, 25) {real, imag} */,
  {32'hc2e257d6, 32'h428073c2} /* (3, 0, 24) {real, imag} */,
  {32'h41c4c22d, 32'h42b3fec3} /* (3, 0, 23) {real, imag} */,
  {32'h42162baa, 32'h42846b08} /* (3, 0, 22) {real, imag} */,
  {32'hc1155080, 32'hc28487f6} /* (3, 0, 21) {real, imag} */,
  {32'h424214b6, 32'h42725419} /* (3, 0, 20) {real, imag} */,
  {32'hc0cb6f38, 32'hc195d12c} /* (3, 0, 19) {real, imag} */,
  {32'h40f00918, 32'hc23c0ce8} /* (3, 0, 18) {real, imag} */,
  {32'hc1690f1c, 32'hc201531a} /* (3, 0, 17) {real, imag} */,
  {32'hc13646c8, 32'hc21b86b4} /* (3, 0, 16) {real, imag} */,
  {32'hc2280867, 32'h41629ea6} /* (3, 0, 15) {real, imag} */,
  {32'h422c18a3, 32'h42a6ac24} /* (3, 0, 14) {real, imag} */,
  {32'hc181a72a, 32'h429dc86d} /* (3, 0, 13) {real, imag} */,
  {32'hc2d18f99, 32'h408b0f18} /* (3, 0, 12) {real, imag} */,
  {32'h4277e490, 32'h41ee88e6} /* (3, 0, 11) {real, imag} */,
  {32'h4301800e, 32'h429d42b4} /* (3, 0, 10) {real, imag} */,
  {32'h41d12fd5, 32'hc22c796e} /* (3, 0, 9) {real, imag} */,
  {32'h42e56964, 32'hc1e0a3d8} /* (3, 0, 8) {real, imag} */,
  {32'hc31ec62a, 32'hc332fd1a} /* (3, 0, 7) {real, imag} */,
  {32'hc3547680, 32'h42681938} /* (3, 0, 6) {real, imag} */,
  {32'h4395434c, 32'hc364d05f} /* (3, 0, 5) {real, imag} */,
  {32'h43372f4a, 32'hc1fc1c81} /* (3, 0, 4) {real, imag} */,
  {32'hc311781a, 32'hc3792164} /* (3, 0, 3) {real, imag} */,
  {32'h434e934c, 32'hc2071224} /* (3, 0, 2) {real, imag} */,
  {32'hc40eb485, 32'h4409e052} /* (3, 0, 1) {real, imag} */,
  {32'hc35da878, 32'h43e39f5c} /* (3, 0, 0) {real, imag} */,
  {32'h449a8ca6, 32'h457e51cd} /* (2, 31, 31) {real, imag} */,
  {32'hc49c278f, 32'hc4efe52a} /* (2, 31, 30) {real, imag} */,
  {32'h423fa34a, 32'hc36f7131} /* (2, 31, 29) {real, imag} */,
  {32'h43749288, 32'h42077330} /* (2, 31, 28) {real, imag} */,
  {32'hc33815ed, 32'hc417d19a} /* (2, 31, 27) {real, imag} */,
  {32'h41502990, 32'hc2845b7a} /* (2, 31, 26) {real, imag} */,
  {32'h43281887, 32'h43087eff} /* (2, 31, 25) {real, imag} */,
  {32'hc3d7245c, 32'hc392be8c} /* (2, 31, 24) {real, imag} */,
  {32'hc229f10c, 32'hc198cb18} /* (2, 31, 23) {real, imag} */,
  {32'h420eca06, 32'hc2e146ee} /* (2, 31, 22) {real, imag} */,
  {32'hc2db0e2e, 32'hc312e070} /* (2, 31, 21) {real, imag} */,
  {32'hc14d603a, 32'h422f69b4} /* (2, 31, 20) {real, imag} */,
  {32'h4171fb38, 32'h4207b4f1} /* (2, 31, 19) {real, imag} */,
  {32'hc300f966, 32'h4233731c} /* (2, 31, 18) {real, imag} */,
  {32'h427a7804, 32'hc2042ef0} /* (2, 31, 17) {real, imag} */,
  {32'h4176d240, 32'h41d4e740} /* (2, 31, 16) {real, imag} */,
  {32'hbf84d780, 32'hc108b740} /* (2, 31, 15) {real, imag} */,
  {32'h42e67c74, 32'h41cecd08} /* (2, 31, 14) {real, imag} */,
  {32'h40479920, 32'hc2a78be6} /* (2, 31, 13) {real, imag} */,
  {32'hc154eca6, 32'hc17c7af0} /* (2, 31, 12) {real, imag} */,
  {32'h4386d478, 32'hc31a1dd8} /* (2, 31, 11) {real, imag} */,
  {32'h41700fb8, 32'h411b6ff0} /* (2, 31, 10) {real, imag} */,
  {32'hc149fc2e, 32'hc2cb6b52} /* (2, 31, 9) {real, imag} */,
  {32'h438f7ca2, 32'hc31630d8} /* (2, 31, 8) {real, imag} */,
  {32'hc3043199, 32'h42eb5eba} /* (2, 31, 7) {real, imag} */,
  {32'h43880448, 32'hc30680db} /* (2, 31, 6) {real, imag} */,
  {32'h439993ea, 32'hc48fe4ac} /* (2, 31, 5) {real, imag} */,
  {32'h43b1f020, 32'h443d8e3f} /* (2, 31, 4) {real, imag} */,
  {32'h42f2449b, 32'hc35fe64b} /* (2, 31, 3) {real, imag} */,
  {32'h4339b1d8, 32'hc477a464} /* (2, 31, 2) {real, imag} */,
  {32'hc48f9594, 32'h45214223} /* (2, 31, 1) {real, imag} */,
  {32'hc3baea6e, 32'h451dc3f4} /* (2, 31, 0) {real, imag} */,
  {32'h44236615, 32'hc4de493e} /* (2, 30, 31) {real, imag} */,
  {32'hc465d2b1, 32'h44a671e6} /* (2, 30, 30) {real, imag} */,
  {32'h42295796, 32'h421cfb63} /* (2, 30, 29) {real, imag} */,
  {32'h426db4a8, 32'hc41b221f} /* (2, 30, 28) {real, imag} */,
  {32'h440d4af3, 32'h44111fd5} /* (2, 30, 27) {real, imag} */,
  {32'h3f2b0f80, 32'hc2c493aa} /* (2, 30, 26) {real, imag} */,
  {32'h4261e91e, 32'hc2bdbe9f} /* (2, 30, 25) {real, imag} */,
  {32'h43653395, 32'h43c3db1c} /* (2, 30, 24) {real, imag} */,
  {32'hc29f9407, 32'hc23fc222} /* (2, 30, 23) {real, imag} */,
  {32'hc2ba0d4b, 32'hc3156a19} /* (2, 30, 22) {real, imag} */,
  {32'h4322cd9c, 32'h429e6a47} /* (2, 30, 21) {real, imag} */,
  {32'h40af64c0, 32'hc21d5574} /* (2, 30, 20) {real, imag} */,
  {32'hc1307838, 32'hc1dd66ea} /* (2, 30, 19) {real, imag} */,
  {32'h430765d0, 32'h4226bd2c} /* (2, 30, 18) {real, imag} */,
  {32'hc1c13a28, 32'hc232bfe0} /* (2, 30, 17) {real, imag} */,
  {32'h4214d1ac, 32'h427691b0} /* (2, 30, 16) {real, imag} */,
  {32'h42de1f3a, 32'h414b7180} /* (2, 30, 15) {real, imag} */,
  {32'hc29567f0, 32'h4259a154} /* (2, 30, 14) {real, imag} */,
  {32'hbfb487c0, 32'h41902582} /* (2, 30, 13) {real, imag} */,
  {32'hc1027f60, 32'hc2c591ae} /* (2, 30, 12) {real, imag} */,
  {32'hc3805cd5, 32'h41b88854} /* (2, 30, 11) {real, imag} */,
  {32'h42652a7e, 32'h40db2100} /* (2, 30, 10) {real, imag} */,
  {32'hc1c3dc54, 32'h4271ac7e} /* (2, 30, 9) {real, imag} */,
  {32'hc41e7e61, 32'h439704fc} /* (2, 30, 8) {real, imag} */,
  {32'h4399a97f, 32'hc24fcd1e} /* (2, 30, 7) {real, imag} */,
  {32'hc280071b, 32'h42f4a9bc} /* (2, 30, 6) {real, imag} */,
  {32'hc3fe4407, 32'h43872992} /* (2, 30, 5) {real, imag} */,
  {32'h44192852, 32'hc3926a80} /* (2, 30, 4) {real, imag} */,
  {32'h42dffc3b, 32'hc1b87a0e} /* (2, 30, 3) {real, imag} */,
  {32'hc48f84e8, 32'h44ffa782} /* (2, 30, 2) {real, imag} */,
  {32'h4420accb, 32'hc54a49df} /* (2, 30, 1) {real, imag} */,
  {32'h423a738c, 32'hc4cde068} /* (2, 30, 0) {real, imag} */,
  {32'h43bf7302, 32'h4439e2e8} /* (2, 29, 31) {real, imag} */,
  {32'hc420e53a, 32'hc321ac7e} /* (2, 29, 30) {real, imag} */,
  {32'h435501b9, 32'h42906d1b} /* (2, 29, 29) {real, imag} */,
  {32'h435a40d6, 32'hc3b03350} /* (2, 29, 28) {real, imag} */,
  {32'h414c7078, 32'hc2620af7} /* (2, 29, 27) {real, imag} */,
  {32'h426f982f, 32'hc0a2c878} /* (2, 29, 26) {real, imag} */,
  {32'h43146677, 32'h428d3ada} /* (2, 29, 25) {real, imag} */,
  {32'hc124a1e8, 32'h42eb6388} /* (2, 29, 24) {real, imag} */,
  {32'h4135396c, 32'h40e5d0bc} /* (2, 29, 23) {real, imag} */,
  {32'h4172a660, 32'hc0ce0308} /* (2, 29, 22) {real, imag} */,
  {32'h422cb8da, 32'h42898de2} /* (2, 29, 21) {real, imag} */,
  {32'hc1a3c080, 32'hc25f870c} /* (2, 29, 20) {real, imag} */,
  {32'hc1c28a98, 32'h40efafc0} /* (2, 29, 19) {real, imag} */,
  {32'hc26f3b1f, 32'hc1ecd2d0} /* (2, 29, 18) {real, imag} */,
  {32'h4139fff0, 32'h421fd0c9} /* (2, 29, 17) {real, imag} */,
  {32'hc1d7a2be, 32'hbfd33a80} /* (2, 29, 16) {real, imag} */,
  {32'h415f5bd0, 32'h411b8064} /* (2, 29, 15) {real, imag} */,
  {32'hc2588b41, 32'h41c6f5b0} /* (2, 29, 14) {real, imag} */,
  {32'hc2d6742c, 32'hc1dbaf80} /* (2, 29, 13) {real, imag} */,
  {32'hc212a288, 32'hc29596f2} /* (2, 29, 12) {real, imag} */,
  {32'hc0cf8e34, 32'hbfbb3640} /* (2, 29, 11) {real, imag} */,
  {32'h4316d8fe, 32'h4252c26f} /* (2, 29, 10) {real, imag} */,
  {32'h42513125, 32'h40aeb01c} /* (2, 29, 9) {real, imag} */,
  {32'hc33712ea, 32'hc2f4e2b8} /* (2, 29, 8) {real, imag} */,
  {32'hbfd97380, 32'h41fa0100} /* (2, 29, 7) {real, imag} */,
  {32'h42dc9fd8, 32'h42d1fd88} /* (2, 29, 6) {real, imag} */,
  {32'h42bbe6eb, 32'hc31587f0} /* (2, 29, 5) {real, imag} */,
  {32'h43166d0a, 32'h4376549f} /* (2, 29, 4) {real, imag} */,
  {32'h41ce3310, 32'h4254dfda} /* (2, 29, 3) {real, imag} */,
  {32'hc41fb1a4, 32'h431f25cc} /* (2, 29, 2) {real, imag} */,
  {32'h44129068, 32'hc417f8ec} /* (2, 29, 1) {real, imag} */,
  {32'hc2de3172, 32'hc165d790} /* (2, 29, 0) {real, imag} */,
  {32'h43618f6e, 32'h4497ddf0} /* (2, 28, 31) {real, imag} */,
  {32'hc3e2ee3b, 32'hc4515d55} /* (2, 28, 30) {real, imag} */,
  {32'h426e939f, 32'h4258aef8} /* (2, 28, 29) {real, imag} */,
  {32'h41abbfb1, 32'hc28d0c11} /* (2, 28, 28) {real, imag} */,
  {32'hc3949ecf, 32'hc2851b33} /* (2, 28, 27) {real, imag} */,
  {32'h4161ad30, 32'hc1f1f322} /* (2, 28, 26) {real, imag} */,
  {32'h427c0ff6, 32'h42b17366} /* (2, 28, 25) {real, imag} */,
  {32'hc2eeb37e, 32'hc321debf} /* (2, 28, 24) {real, imag} */,
  {32'h427ab29a, 32'hc213988b} /* (2, 28, 23) {real, imag} */,
  {32'h43096fe9, 32'hc2520a3b} /* (2, 28, 22) {real, imag} */,
  {32'hc2141ca9, 32'h41695b28} /* (2, 28, 21) {real, imag} */,
  {32'h412c6b20, 32'h422f2003} /* (2, 28, 20) {real, imag} */,
  {32'h410048fa, 32'hc05dedc0} /* (2, 28, 19) {real, imag} */,
  {32'hc2b0e644, 32'hc202989e} /* (2, 28, 18) {real, imag} */,
  {32'h427f1042, 32'hc1aac720} /* (2, 28, 17) {real, imag} */,
  {32'hc0bf27cc, 32'h421a8148} /* (2, 28, 16) {real, imag} */,
  {32'hc15e0c08, 32'h42501f30} /* (2, 28, 15) {real, imag} */,
  {32'hbffdb2e0, 32'hc2a729c9} /* (2, 28, 14) {real, imag} */,
  {32'hc155b052, 32'h418c3480} /* (2, 28, 13) {real, imag} */,
  {32'hc2d6df8c, 32'h42a31e0c} /* (2, 28, 12) {real, imag} */,
  {32'h42d02030, 32'hc30049b4} /* (2, 28, 11) {real, imag} */,
  {32'hc220723c, 32'h4171a05c} /* (2, 28, 10) {real, imag} */,
  {32'hc3017fec, 32'h42507801} /* (2, 28, 9) {real, imag} */,
  {32'hc2293fc4, 32'hc25f7698} /* (2, 28, 8) {real, imag} */,
  {32'hc25711ee, 32'hc074e910} /* (2, 28, 7) {real, imag} */,
  {32'h431df7ef, 32'h420878b5} /* (2, 28, 6) {real, imag} */,
  {32'h42c443d0, 32'hc39627c9} /* (2, 28, 5) {real, imag} */,
  {32'h4229d978, 32'h4370ce9c} /* (2, 28, 4) {real, imag} */,
  {32'hc1af5a6a, 32'hc1f39108} /* (2, 28, 3) {real, imag} */,
  {32'hc401cb0d, 32'hc4280d93} /* (2, 28, 2) {real, imag} */,
  {32'h441a08e0, 32'h43fddd74} /* (2, 28, 1) {real, imag} */,
  {32'h40c9c47c, 32'h43d13c11} /* (2, 28, 0) {real, imag} */,
  {32'hc4270033, 32'hc4410574} /* (2, 27, 31) {real, imag} */,
  {32'h4365869a, 32'h4356c668} /* (2, 27, 30) {real, imag} */,
  {32'hc2c96c14, 32'hc2dd4f9f} /* (2, 27, 29) {real, imag} */,
  {32'hc29caacc, 32'h4242db99} /* (2, 27, 28) {real, imag} */,
  {32'hc1b1b1c0, 32'h4358fed4} /* (2, 27, 27) {real, imag} */,
  {32'h42cba9b0, 32'h42609924} /* (2, 27, 26) {real, imag} */,
  {32'hc240ba0a, 32'hc27752bf} /* (2, 27, 25) {real, imag} */,
  {32'h4154f618, 32'hc286b4dd} /* (2, 27, 24) {real, imag} */,
  {32'h421342ce, 32'h4190a70c} /* (2, 27, 23) {real, imag} */,
  {32'hc1d39fd6, 32'hc1804570} /* (2, 27, 22) {real, imag} */,
  {32'h42c33362, 32'hc1d034f2} /* (2, 27, 21) {real, imag} */,
  {32'h41f2074a, 32'h41dcde56} /* (2, 27, 20) {real, imag} */,
  {32'h4218609f, 32'hc2356125} /* (2, 27, 19) {real, imag} */,
  {32'h427ca22e, 32'hc1901886} /* (2, 27, 18) {real, imag} */,
  {32'h42424610, 32'h4090c038} /* (2, 27, 17) {real, imag} */,
  {32'hc2643512, 32'hc1c21e70} /* (2, 27, 16) {real, imag} */,
  {32'hc10b2960, 32'hc082c438} /* (2, 27, 15) {real, imag} */,
  {32'hc21087de, 32'hc200e9dd} /* (2, 27, 14) {real, imag} */,
  {32'h41ce867a, 32'h422f5cfb} /* (2, 27, 13) {real, imag} */,
  {32'hc191c01e, 32'h41847e2e} /* (2, 27, 12) {real, imag} */,
  {32'hc2b563e2, 32'h41da194a} /* (2, 27, 11) {real, imag} */,
  {32'hc182a872, 32'h43199ff4} /* (2, 27, 10) {real, imag} */,
  {32'h41601158, 32'hc0185800} /* (2, 27, 9) {real, imag} */,
  {32'hc2d56597, 32'h422e74b2} /* (2, 27, 8) {real, imag} */,
  {32'hc2aaad71, 32'hc2b666a4} /* (2, 27, 7) {real, imag} */,
  {32'hc2ba3fe0, 32'h429e51e2} /* (2, 27, 6) {real, imag} */,
  {32'h434db3ea, 32'h435e4b48} /* (2, 27, 5) {real, imag} */,
  {32'h4375339a, 32'hc1f20a46} /* (2, 27, 4) {real, imag} */,
  {32'hc2b0f36e, 32'hc27d6582} /* (2, 27, 3) {real, imag} */,
  {32'hc30643fa, 32'h43942bea} /* (2, 27, 2) {real, imag} */,
  {32'hc1d5a9a0, 32'hc46606d8} /* (2, 27, 1) {real, imag} */,
  {32'hc3258e78, 32'hc41f9ef6} /* (2, 27, 0) {real, imag} */,
  {32'hc2049112, 32'hc18215a0} /* (2, 26, 31) {real, imag} */,
  {32'h424c1c4e, 32'h432332a8} /* (2, 26, 30) {real, imag} */,
  {32'h42fd0614, 32'hc2547d8c} /* (2, 26, 29) {real, imag} */,
  {32'hc2840037, 32'hc285a730} /* (2, 26, 28) {real, imag} */,
  {32'hc26ee071, 32'h4325f949} /* (2, 26, 27) {real, imag} */,
  {32'hc24f8864, 32'h3fb97c40} /* (2, 26, 26) {real, imag} */,
  {32'h41ed6965, 32'h4172c4f6} /* (2, 26, 25) {real, imag} */,
  {32'hc2116c64, 32'h42af178a} /* (2, 26, 24) {real, imag} */,
  {32'hc295bed5, 32'hc27aa33a} /* (2, 26, 23) {real, imag} */,
  {32'hc1dda1d8, 32'hc116cdc2} /* (2, 26, 22) {real, imag} */,
  {32'h41c2b8a8, 32'h4252ba5b} /* (2, 26, 21) {real, imag} */,
  {32'h41cff8f1, 32'h4044d490} /* (2, 26, 20) {real, imag} */,
  {32'h416102dc, 32'h41b04966} /* (2, 26, 19) {real, imag} */,
  {32'hc19e8340, 32'h4116e484} /* (2, 26, 18) {real, imag} */,
  {32'hc1aee871, 32'h414c7b80} /* (2, 26, 17) {real, imag} */,
  {32'h424725c8, 32'hc1666cc6} /* (2, 26, 16) {real, imag} */,
  {32'h419fe181, 32'h41672778} /* (2, 26, 15) {real, imag} */,
  {32'hbf5d3ab0, 32'h420cc0e1} /* (2, 26, 14) {real, imag} */,
  {32'hc1502b44, 32'h421b272d} /* (2, 26, 13) {real, imag} */,
  {32'hc2132704, 32'hc2177e49} /* (2, 26, 12) {real, imag} */,
  {32'h41fe3364, 32'h425dd87f} /* (2, 26, 11) {real, imag} */,
  {32'h419677dc, 32'h41746fa2} /* (2, 26, 10) {real, imag} */,
  {32'hc195a43c, 32'h42d9de23} /* (2, 26, 9) {real, imag} */,
  {32'h42b24902, 32'h41e92cf6} /* (2, 26, 8) {real, imag} */,
  {32'h41415fea, 32'h41d2075b} /* (2, 26, 7) {real, imag} */,
  {32'h433ffe4d, 32'h429069ef} /* (2, 26, 6) {real, imag} */,
  {32'h40a30c48, 32'h42473f44} /* (2, 26, 5) {real, imag} */,
  {32'hc35b0684, 32'hc1cdde0a} /* (2, 26, 4) {real, imag} */,
  {32'hc20987f5, 32'h42e1909e} /* (2, 26, 3) {real, imag} */,
  {32'hc12cebbe, 32'h42b8c494} /* (2, 26, 2) {real, imag} */,
  {32'hc2f1fd13, 32'hc312a7d0} /* (2, 26, 1) {real, imag} */,
  {32'h42474ea4, 32'h425e7f2a} /* (2, 26, 0) {real, imag} */,
  {32'h436f5f45, 32'h42f9ba94} /* (2, 25, 31) {real, imag} */,
  {32'hc24876a5, 32'h40e384d0} /* (2, 25, 30) {real, imag} */,
  {32'hc1faec9b, 32'h42a42d6b} /* (2, 25, 29) {real, imag} */,
  {32'hc0f19b70, 32'hc25ab0ea} /* (2, 25, 28) {real, imag} */,
  {32'hc2f13c02, 32'hc2bee870} /* (2, 25, 27) {real, imag} */,
  {32'hc3091135, 32'h424048a9} /* (2, 25, 26) {real, imag} */,
  {32'hc1a6753a, 32'h4099a804} /* (2, 25, 25) {real, imag} */,
  {32'hc2839ef4, 32'h4293757c} /* (2, 25, 24) {real, imag} */,
  {32'hc275dbf1, 32'hc19c3e0f} /* (2, 25, 23) {real, imag} */,
  {32'h40d32048, 32'hc2253a7a} /* (2, 25, 22) {real, imag} */,
  {32'h4087179c, 32'h42348296} /* (2, 25, 21) {real, imag} */,
  {32'h413d4598, 32'hc09ae8dc} /* (2, 25, 20) {real, imag} */,
  {32'hc2447e66, 32'h40620b70} /* (2, 25, 19) {real, imag} */,
  {32'h411d9759, 32'h41a08ad0} /* (2, 25, 18) {real, imag} */,
  {32'hc1135e08, 32'h41b9ec84} /* (2, 25, 17) {real, imag} */,
  {32'h427ddeaa, 32'hc20601bf} /* (2, 25, 16) {real, imag} */,
  {32'hc18025dc, 32'hc22601c8} /* (2, 25, 15) {real, imag} */,
  {32'h41b6ff48, 32'hc2491d60} /* (2, 25, 14) {real, imag} */,
  {32'h42024f1e, 32'h42cf2e90} /* (2, 25, 13) {real, imag} */,
  {32'hc10efc10, 32'h418f10c3} /* (2, 25, 12) {real, imag} */,
  {32'hc0cdb394, 32'hc0dfcd3c} /* (2, 25, 11) {real, imag} */,
  {32'h41ec98f6, 32'h420313f4} /* (2, 25, 10) {real, imag} */,
  {32'hc248cda5, 32'hc1f5b2b7} /* (2, 25, 9) {real, imag} */,
  {32'hc214511c, 32'hc2968686} /* (2, 25, 8) {real, imag} */,
  {32'hc0fa38e6, 32'h422d3d58} /* (2, 25, 7) {real, imag} */,
  {32'h422f275c, 32'h41955306} /* (2, 25, 6) {real, imag} */,
  {32'h41c185d8, 32'hc1f29f7e} /* (2, 25, 5) {real, imag} */,
  {32'hc22a150e, 32'hc2b7d37b} /* (2, 25, 4) {real, imag} */,
  {32'hc1935713, 32'h424247da} /* (2, 25, 3) {real, imag} */,
  {32'hc20f083d, 32'hc202339a} /* (2, 25, 2) {real, imag} */,
  {32'h42fa430e, 32'h42bd8edc} /* (2, 25, 1) {real, imag} */,
  {32'h434c8c52, 32'h42c257c0} /* (2, 25, 0) {real, imag} */,
  {32'hc361340c, 32'hc3af5316} /* (2, 24, 31) {real, imag} */,
  {32'h42e7b864, 32'h432540ea} /* (2, 24, 30) {real, imag} */,
  {32'h41a9e904, 32'hc16add20} /* (2, 24, 29) {real, imag} */,
  {32'hc26726cb, 32'hc32a4501} /* (2, 24, 28) {real, imag} */,
  {32'h4332a462, 32'h430ae316} /* (2, 24, 27) {real, imag} */,
  {32'h4212a4b4, 32'h42ab2067} /* (2, 24, 26) {real, imag} */,
  {32'hc2aa0286, 32'h41caab05} /* (2, 24, 25) {real, imag} */,
  {32'h4256f98b, 32'h425e71c3} /* (2, 24, 24) {real, imag} */,
  {32'hc148a6a5, 32'hbff7dee0} /* (2, 24, 23) {real, imag} */,
  {32'hc293459f, 32'h3eaced00} /* (2, 24, 22) {real, imag} */,
  {32'h4218a4ae, 32'h41f05804} /* (2, 24, 21) {real, imag} */,
  {32'h41fdf99e, 32'hc1aa7214} /* (2, 24, 20) {real, imag} */,
  {32'h41725f5c, 32'hc0525830} /* (2, 24, 19) {real, imag} */,
  {32'h40935fd2, 32'hbe328a00} /* (2, 24, 18) {real, imag} */,
  {32'hc0c43f54, 32'hc013cfa0} /* (2, 24, 17) {real, imag} */,
  {32'hc145a060, 32'hc020f100} /* (2, 24, 16) {real, imag} */,
  {32'h41e0f3a5, 32'h414ee5a8} /* (2, 24, 15) {real, imag} */,
  {32'h4164f979, 32'h3fc24240} /* (2, 24, 14) {real, imag} */,
  {32'h415ebbec, 32'h3eb65e00} /* (2, 24, 13) {real, imag} */,
  {32'hbf6fb240, 32'h423f5f1c} /* (2, 24, 12) {real, imag} */,
  {32'hc15c77f8, 32'h428ab257} /* (2, 24, 11) {real, imag} */,
  {32'h3e193600, 32'h430b2cdc} /* (2, 24, 10) {real, imag} */,
  {32'hbf0e9e30, 32'hc28c7a80} /* (2, 24, 9) {real, imag} */,
  {32'hc22042e1, 32'h4207c3c1} /* (2, 24, 8) {real, imag} */,
  {32'hc2d5479e, 32'hc22af68c} /* (2, 24, 7) {real, imag} */,
  {32'h402d6048, 32'hc2dbba0d} /* (2, 24, 6) {real, imag} */,
  {32'h42916811, 32'h42654c6e} /* (2, 24, 5) {real, imag} */,
  {32'hc27457e3, 32'hc1dafaa8} /* (2, 24, 4) {real, imag} */,
  {32'hc3173aea, 32'h420fb1c7} /* (2, 24, 3) {real, imag} */,
  {32'hc2a8daf2, 32'h43b09143} /* (2, 24, 2) {real, imag} */,
  {32'hc3adac72, 32'hc43359a1} /* (2, 24, 1) {real, imag} */,
  {32'hc27c6876, 32'hc3b86c38} /* (2, 24, 0) {real, imag} */,
  {32'h43402ff3, 32'h43398617} /* (2, 23, 31) {real, imag} */,
  {32'hc3266e86, 32'hc12b2ce8} /* (2, 23, 30) {real, imag} */,
  {32'hc350f001, 32'hc25e35ca} /* (2, 23, 29) {real, imag} */,
  {32'h431b6ff6, 32'hc105b984} /* (2, 23, 28) {real, imag} */,
  {32'h42a42bba, 32'h42836dae} /* (2, 23, 27) {real, imag} */,
  {32'h417b3df4, 32'h423c593c} /* (2, 23, 26) {real, imag} */,
  {32'h4207d026, 32'h3fd47a40} /* (2, 23, 25) {real, imag} */,
  {32'hc2f2c975, 32'hc182410d} /* (2, 23, 24) {real, imag} */,
  {32'h42162f83, 32'h41a86cda} /* (2, 23, 23) {real, imag} */,
  {32'hc1b291ab, 32'hc28198ce} /* (2, 23, 22) {real, imag} */,
  {32'hc2526777, 32'h40713f78} /* (2, 23, 21) {real, imag} */,
  {32'hc0f55a40, 32'h41779a9a} /* (2, 23, 20) {real, imag} */,
  {32'h42172379, 32'hc21467e4} /* (2, 23, 19) {real, imag} */,
  {32'hc105f056, 32'h41bcd1c0} /* (2, 23, 18) {real, imag} */,
  {32'hc1978bf9, 32'hc17a209e} /* (2, 23, 17) {real, imag} */,
  {32'h41cf1294, 32'hc1114541} /* (2, 23, 16) {real, imag} */,
  {32'h41a7e769, 32'h40bc1703} /* (2, 23, 15) {real, imag} */,
  {32'h414e6516, 32'h4204d180} /* (2, 23, 14) {real, imag} */,
  {32'hc14cdf2c, 32'h4261574e} /* (2, 23, 13) {real, imag} */,
  {32'hc2531de0, 32'h4229bd88} /* (2, 23, 12) {real, imag} */,
  {32'h41d18cd2, 32'hc24118a4} /* (2, 23, 11) {real, imag} */,
  {32'hc220cbe4, 32'hc29713d2} /* (2, 23, 10) {real, imag} */,
  {32'h421f2a15, 32'h41f1d3fc} /* (2, 23, 9) {real, imag} */,
  {32'hc1d87504, 32'hc1ef0aff} /* (2, 23, 8) {real, imag} */,
  {32'h41a8918c, 32'h4196a786} /* (2, 23, 7) {real, imag} */,
  {32'h42c49fbe, 32'hc25751aa} /* (2, 23, 6) {real, imag} */,
  {32'hc23003e5, 32'hc0db97c4} /* (2, 23, 5) {real, imag} */,
  {32'h4248504a, 32'h427e38a7} /* (2, 23, 4) {real, imag} */,
  {32'h42a9d896, 32'h409676bc} /* (2, 23, 3) {real, imag} */,
  {32'hc348f286, 32'hc202ccce} /* (2, 23, 2) {real, imag} */,
  {32'h42a5c1ce, 32'hc33e0d4f} /* (2, 23, 1) {real, imag} */,
  {32'h41e289de, 32'h3dfce180} /* (2, 23, 0) {real, imag} */,
  {32'h428bfc50, 32'h43192d8e} /* (2, 22, 31) {real, imag} */,
  {32'hc2b6092d, 32'hc32dc03f} /* (2, 22, 30) {real, imag} */,
  {32'h4204d820, 32'h41eb3554} /* (2, 22, 29) {real, imag} */,
  {32'h428fcb8b, 32'h425086ec} /* (2, 22, 28) {real, imag} */,
  {32'hc11d1f29, 32'h4282f3ca} /* (2, 22, 27) {real, imag} */,
  {32'hc0fe8f1a, 32'h42cee914} /* (2, 22, 26) {real, imag} */,
  {32'hc1b9911d, 32'h417d8608} /* (2, 22, 25) {real, imag} */,
  {32'hc24d0a5a, 32'hc1ffae8f} /* (2, 22, 24) {real, imag} */,
  {32'hbfa6c240, 32'h421d8bec} /* (2, 22, 23) {real, imag} */,
  {32'h421c3f11, 32'hc203d51d} /* (2, 22, 22) {real, imag} */,
  {32'h416ea898, 32'hc1fb4316} /* (2, 22, 21) {real, imag} */,
  {32'hc2080f6d, 32'hc1575e80} /* (2, 22, 20) {real, imag} */,
  {32'hc17fcb80, 32'h41ecd942} /* (2, 22, 19) {real, imag} */,
  {32'hc1b3c318, 32'h40ab4514} /* (2, 22, 18) {real, imag} */,
  {32'h40c40ea0, 32'hc10f308e} /* (2, 22, 17) {real, imag} */,
  {32'h41b7dceb, 32'hc1d5859f} /* (2, 22, 16) {real, imag} */,
  {32'h41304c20, 32'h41a27551} /* (2, 22, 15) {real, imag} */,
  {32'h41b16540, 32'h414af992} /* (2, 22, 14) {real, imag} */,
  {32'h41f8c024, 32'h40e8b832} /* (2, 22, 13) {real, imag} */,
  {32'hc1080a50, 32'hc08e4ea5} /* (2, 22, 12) {real, imag} */,
  {32'hc258beb4, 32'h41c6c376} /* (2, 22, 11) {real, imag} */,
  {32'hc1bb6622, 32'h41e0f066} /* (2, 22, 10) {real, imag} */,
  {32'h3fdde7e0, 32'hbfaa0c00} /* (2, 22, 9) {real, imag} */,
  {32'hc1d0fd6b, 32'hc2727656} /* (2, 22, 8) {real, imag} */,
  {32'h4235fd8e, 32'hc242482a} /* (2, 22, 7) {real, imag} */,
  {32'hc17247a5, 32'hc266b4ff} /* (2, 22, 6) {real, imag} */,
  {32'hc18f940c, 32'hc2b27dfe} /* (2, 22, 5) {real, imag} */,
  {32'hc23568ae, 32'h4155ab3a} /* (2, 22, 4) {real, imag} */,
  {32'h42a4ca0b, 32'h4227fb86} /* (2, 22, 3) {real, imag} */,
  {32'hc19e5354, 32'h428a12b2} /* (2, 22, 2) {real, imag} */,
  {32'h434faa34, 32'hc27ca70c} /* (2, 22, 1) {real, imag} */,
  {32'h428a570d, 32'h413ebb66} /* (2, 22, 0) {real, imag} */,
  {32'hc37ec771, 32'hc30da39e} /* (2, 21, 31) {real, imag} */,
  {32'h4319306d, 32'h41b24cba} /* (2, 21, 30) {real, imag} */,
  {32'hc18e8312, 32'h426bfa12} /* (2, 21, 29) {real, imag} */,
  {32'hc2124734, 32'h42150820} /* (2, 21, 28) {real, imag} */,
  {32'h42d6ce88, 32'h4248f7a9} /* (2, 21, 27) {real, imag} */,
  {32'h4220c4ce, 32'hc244c9ef} /* (2, 21, 26) {real, imag} */,
  {32'hc11f140a, 32'h42386918} /* (2, 21, 25) {real, imag} */,
  {32'h42896e33, 32'h40b4d2f0} /* (2, 21, 24) {real, imag} */,
  {32'hc1cf93db, 32'h4208396a} /* (2, 21, 23) {real, imag} */,
  {32'h42519d12, 32'h42bbb0d4} /* (2, 21, 22) {real, imag} */,
  {32'h41d0bc03, 32'h41d12ecb} /* (2, 21, 21) {real, imag} */,
  {32'hc233fed2, 32'h3df79380} /* (2, 21, 20) {real, imag} */,
  {32'h41391205, 32'hbf151410} /* (2, 21, 19) {real, imag} */,
  {32'hc0ddc4f4, 32'hc120ba79} /* (2, 21, 18) {real, imag} */,
  {32'hc0520d40, 32'h408332cc} /* (2, 21, 17) {real, imag} */,
  {32'hc1eedc6a, 32'hc1791388} /* (2, 21, 16) {real, imag} */,
  {32'h41cca3a8, 32'hc09bd22c} /* (2, 21, 15) {real, imag} */,
  {32'h402daac8, 32'h40169d84} /* (2, 21, 14) {real, imag} */,
  {32'hc0fa2496, 32'h404118c4} /* (2, 21, 13) {real, imag} */,
  {32'hc168fe80, 32'hc195082a} /* (2, 21, 12) {real, imag} */,
  {32'h41426aaa, 32'h423d529e} /* (2, 21, 11) {real, imag} */,
  {32'h41c8f378, 32'hc1a618fa} /* (2, 21, 10) {real, imag} */,
  {32'h41630ade, 32'h41b0570f} /* (2, 21, 9) {real, imag} */,
  {32'hc032d8e0, 32'h4290e87e} /* (2, 21, 8) {real, imag} */,
  {32'hc1f734af, 32'h416060ba} /* (2, 21, 7) {real, imag} */,
  {32'h41d95e28, 32'hc2849fb6} /* (2, 21, 6) {real, imag} */,
  {32'h426a9e68, 32'h42931dde} /* (2, 21, 5) {real, imag} */,
  {32'h42a62c8b, 32'hbf7b5de0} /* (2, 21, 4) {real, imag} */,
  {32'hc22009f9, 32'h42d2d85d} /* (2, 21, 3) {real, imag} */,
  {32'h427b62cc, 32'h42565ff9} /* (2, 21, 2) {real, imag} */,
  {32'hc337664b, 32'hc356faf2} /* (2, 21, 1) {real, imag} */,
  {32'hc2e75818, 32'hc37c5288} /* (2, 21, 0) {real, imag} */,
  {32'h41d62370, 32'hc1ba7dc9} /* (2, 20, 31) {real, imag} */,
  {32'hc240137a, 32'h40b48c66} /* (2, 20, 30) {real, imag} */,
  {32'h424e30c0, 32'h4226b801} /* (2, 20, 29) {real, imag} */,
  {32'hc1f2b55e, 32'h4212961c} /* (2, 20, 28) {real, imag} */,
  {32'h3f9b2a58, 32'h42017c31} /* (2, 20, 27) {real, imag} */,
  {32'h40058e7c, 32'h4259df1e} /* (2, 20, 26) {real, imag} */,
  {32'hc1b844b6, 32'hc1572328} /* (2, 20, 25) {real, imag} */,
  {32'h411eb543, 32'h414ede7c} /* (2, 20, 24) {real, imag} */,
  {32'hc112c2d6, 32'hc2ac6ac2} /* (2, 20, 23) {real, imag} */,
  {32'h41580539, 32'h4214cb81} /* (2, 20, 22) {real, imag} */,
  {32'h41468e33, 32'h417bdaa6} /* (2, 20, 21) {real, imag} */,
  {32'hc1cee3a3, 32'hc149987c} /* (2, 20, 20) {real, imag} */,
  {32'hc18e2508, 32'h418972b7} /* (2, 20, 19) {real, imag} */,
  {32'hc0ac70eb, 32'hc1d7f7ac} /* (2, 20, 18) {real, imag} */,
  {32'h3fd2e160, 32'h400af3c4} /* (2, 20, 17) {real, imag} */,
  {32'hc042deb8, 32'hbf052280} /* (2, 20, 16) {real, imag} */,
  {32'hc1a9709e, 32'hc1223beb} /* (2, 20, 15) {real, imag} */,
  {32'hc0706066, 32'hc184bdc0} /* (2, 20, 14) {real, imag} */,
  {32'h411abc1b, 32'h405fb568} /* (2, 20, 13) {real, imag} */,
  {32'h4105b682, 32'hc209bc0b} /* (2, 20, 12) {real, imag} */,
  {32'h3f8957c8, 32'hc01cae78} /* (2, 20, 11) {real, imag} */,
  {32'hc129badf, 32'h412c0cd8} /* (2, 20, 10) {real, imag} */,
  {32'hc23b9a10, 32'hc1e64ff6} /* (2, 20, 9) {real, imag} */,
  {32'h42226ba8, 32'hc1a238c8} /* (2, 20, 8) {real, imag} */,
  {32'hc044c48c, 32'h40198a20} /* (2, 20, 7) {real, imag} */,
  {32'hc1e182d4, 32'h41e744bd} /* (2, 20, 6) {real, imag} */,
  {32'h418f1630, 32'hc2179563} /* (2, 20, 5) {real, imag} */,
  {32'hc15346e7, 32'h411ac8f0} /* (2, 20, 4) {real, imag} */,
  {32'hc029a338, 32'hc16139e8} /* (2, 20, 3) {real, imag} */,
  {32'h4266d1a6, 32'h40a5cf8a} /* (2, 20, 2) {real, imag} */,
  {32'h429e6c41, 32'hc1a1a41b} /* (2, 20, 1) {real, imag} */,
  {32'hc27a99f8, 32'h4299642f} /* (2, 20, 0) {real, imag} */,
  {32'h42852174, 32'h42e13528} /* (2, 19, 31) {real, imag} */,
  {32'hc09dc0d1, 32'hc1d03f37} /* (2, 19, 30) {real, imag} */,
  {32'hc166517e, 32'hc13fa0da} /* (2, 19, 29) {real, imag} */,
  {32'h41f93d06, 32'h425e2a38} /* (2, 19, 28) {real, imag} */,
  {32'hc173cf1b, 32'hc242feb0} /* (2, 19, 27) {real, imag} */,
  {32'hc1cbf1b2, 32'hc220b54a} /* (2, 19, 26) {real, imag} */,
  {32'hc1ade94e, 32'h42916be0} /* (2, 19, 25) {real, imag} */,
  {32'hc2043d48, 32'hc0dab934} /* (2, 19, 24) {real, imag} */,
  {32'h419c0716, 32'hc165da26} /* (2, 19, 23) {real, imag} */,
  {32'hc10265eb, 32'hbf184260} /* (2, 19, 22) {real, imag} */,
  {32'hc120c750, 32'hc0ddda3c} /* (2, 19, 21) {real, imag} */,
  {32'hc1864210, 32'h411dadd4} /* (2, 19, 20) {real, imag} */,
  {32'h4006fafe, 32'h40c5ac1d} /* (2, 19, 19) {real, imag} */,
  {32'hc101dde6, 32'h41cf9884} /* (2, 19, 18) {real, imag} */,
  {32'h40edcf4a, 32'h4017d888} /* (2, 19, 17) {real, imag} */,
  {32'h41919657, 32'h3c12c000} /* (2, 19, 16) {real, imag} */,
  {32'hbfa035e8, 32'hc0d37944} /* (2, 19, 15) {real, imag} */,
  {32'h418e1739, 32'hc13f5a68} /* (2, 19, 14) {real, imag} */,
  {32'h3f8cc4a4, 32'hc018e2be} /* (2, 19, 13) {real, imag} */,
  {32'h41a7ac6c, 32'h3fa927fc} /* (2, 19, 12) {real, imag} */,
  {32'h3dc54cc0, 32'hc16c31d6} /* (2, 19, 11) {real, imag} */,
  {32'h41282283, 32'h41ecb167} /* (2, 19, 10) {real, imag} */,
  {32'h41a40452, 32'h4182777f} /* (2, 19, 9) {real, imag} */,
  {32'hc176a6f8, 32'hc18d64d5} /* (2, 19, 8) {real, imag} */,
  {32'hc21337bd, 32'h3f92ce80} /* (2, 19, 7) {real, imag} */,
  {32'hc28fcadc, 32'h4294cd69} /* (2, 19, 6) {real, imag} */,
  {32'h411176f5, 32'h424d6826} /* (2, 19, 5) {real, imag} */,
  {32'h41e08c9e, 32'h42954a4e} /* (2, 19, 4) {real, imag} */,
  {32'hc1d56011, 32'h40e8b270} /* (2, 19, 3) {real, imag} */,
  {32'h3e912b90, 32'h415aeada} /* (2, 19, 2) {real, imag} */,
  {32'h416edcd8, 32'h41be4fd0} /* (2, 19, 1) {real, imag} */,
  {32'h4283b25b, 32'h41b4f546} /* (2, 19, 0) {real, imag} */,
  {32'hc2936cda, 32'h4215fa9e} /* (2, 18, 31) {real, imag} */,
  {32'h414058ae, 32'hc1ee52e4} /* (2, 18, 30) {real, imag} */,
  {32'h41871741, 32'h406e0244} /* (2, 18, 29) {real, imag} */,
  {32'h3f204700, 32'hc20764cc} /* (2, 18, 28) {real, imag} */,
  {32'h41f5e5bd, 32'hc20eee69} /* (2, 18, 27) {real, imag} */,
  {32'h4234eb86, 32'h419b0419} /* (2, 18, 26) {real, imag} */,
  {32'h419ab10b, 32'h40a0bd0b} /* (2, 18, 25) {real, imag} */,
  {32'h41822b3c, 32'h411f6dd0} /* (2, 18, 24) {real, imag} */,
  {32'h401de938, 32'h420a4cba} /* (2, 18, 23) {real, imag} */,
  {32'hc16209c6, 32'h41f479ba} /* (2, 18, 22) {real, imag} */,
  {32'h4145b670, 32'hc05ef24e} /* (2, 18, 21) {real, imag} */,
  {32'h4180b1be, 32'hc1632266} /* (2, 18, 20) {real, imag} */,
  {32'hc18d1994, 32'h3f1d4970} /* (2, 18, 19) {real, imag} */,
  {32'h411525c0, 32'h410ca1ad} /* (2, 18, 18) {real, imag} */,
  {32'hbfac7a54, 32'hc0ed19d4} /* (2, 18, 17) {real, imag} */,
  {32'hc146f328, 32'h40277508} /* (2, 18, 16) {real, imag} */,
  {32'h40b6b285, 32'h40ff774c} /* (2, 18, 15) {real, imag} */,
  {32'h4136a9ba, 32'hc0420b1c} /* (2, 18, 14) {real, imag} */,
  {32'h413fa720, 32'hc17fbf85} /* (2, 18, 13) {real, imag} */,
  {32'hc12bd637, 32'hbfcf9010} /* (2, 18, 12) {real, imag} */,
  {32'hbed7f310, 32'h40b868f9} /* (2, 18, 11) {real, imag} */,
  {32'h409f489c, 32'h412d9404} /* (2, 18, 10) {real, imag} */,
  {32'h3fdda870, 32'hc1506888} /* (2, 18, 9) {real, imag} */,
  {32'h41ca4710, 32'h4259325e} /* (2, 18, 8) {real, imag} */,
  {32'hc175f5c2, 32'h3fa0016c} /* (2, 18, 7) {real, imag} */,
  {32'h41a51003, 32'h41aa4b07} /* (2, 18, 6) {real, imag} */,
  {32'hc0896a54, 32'h4211a8ed} /* (2, 18, 5) {real, imag} */,
  {32'hc2900790, 32'hc2f746ce} /* (2, 18, 4) {real, imag} */,
  {32'h423d1730, 32'hc1d9de6e} /* (2, 18, 3) {real, imag} */,
  {32'h42198180, 32'h42a04db1} /* (2, 18, 2) {real, imag} */,
  {32'hc2cd7b7e, 32'hc2eabfd3} /* (2, 18, 1) {real, imag} */,
  {32'hc2a77c88, 32'h4228e8aa} /* (2, 18, 0) {real, imag} */,
  {32'h4245332e, 32'h41e047ba} /* (2, 17, 31) {real, imag} */,
  {32'hc27f8f5f, 32'h416a21e7} /* (2, 17, 30) {real, imag} */,
  {32'hc11ab296, 32'hc03e9374} /* (2, 17, 29) {real, imag} */,
  {32'h4202c30a, 32'hc243aa60} /* (2, 17, 28) {real, imag} */,
  {32'hc16c4280, 32'h41b40e34} /* (2, 17, 27) {real, imag} */,
  {32'h4201d340, 32'hc20abd32} /* (2, 17, 26) {real, imag} */,
  {32'h3d6dd380, 32'h424dc8c6} /* (2, 17, 25) {real, imag} */,
  {32'hc164169c, 32'h416ec949} /* (2, 17, 24) {real, imag} */,
  {32'h41b616d6, 32'h4020d5dc} /* (2, 17, 23) {real, imag} */,
  {32'h4196a946, 32'hc188e540} /* (2, 17, 22) {real, imag} */,
  {32'h4082ebeb, 32'h41a2fd2f} /* (2, 17, 21) {real, imag} */,
  {32'hc0ce7006, 32'hc1921c9b} /* (2, 17, 20) {real, imag} */,
  {32'h3fb63008, 32'h3f03d4a0} /* (2, 17, 19) {real, imag} */,
  {32'hc1c0e9ca, 32'h40c40ba4} /* (2, 17, 18) {real, imag} */,
  {32'hc1077516, 32'hbecd0760} /* (2, 17, 17) {real, imag} */,
  {32'h40041880, 32'hc12855ce} /* (2, 17, 16) {real, imag} */,
  {32'hc0e5b774, 32'h41877c16} /* (2, 17, 15) {real, imag} */,
  {32'h404cf680, 32'hc1953856} /* (2, 17, 14) {real, imag} */,
  {32'hc037e660, 32'h3fcf16d0} /* (2, 17, 13) {real, imag} */,
  {32'hc043176c, 32'h3f751ce0} /* (2, 17, 12) {real, imag} */,
  {32'hc0c64fd5, 32'h410e91ee} /* (2, 17, 11) {real, imag} */,
  {32'h41aaa4a6, 32'hc0bd627a} /* (2, 17, 10) {real, imag} */,
  {32'hc119a460, 32'hc0c3a456} /* (2, 17, 9) {real, imag} */,
  {32'h4183d676, 32'h411eef2d} /* (2, 17, 8) {real, imag} */,
  {32'hc06d9d22, 32'hc1a1f54d} /* (2, 17, 7) {real, imag} */,
  {32'h41b499ad, 32'h41c2db41} /* (2, 17, 6) {real, imag} */,
  {32'h41d506d2, 32'h3ec4bc00} /* (2, 17, 5) {real, imag} */,
  {32'hc0a83a2e, 32'h4259a864} /* (2, 17, 4) {real, imag} */,
  {32'h3f55eed0, 32'h41ae4512} /* (2, 17, 3) {real, imag} */,
  {32'hc2969dc8, 32'hc0a64de6} /* (2, 17, 2) {real, imag} */,
  {32'h42d8b7bb, 32'hc208a035} /* (2, 17, 1) {real, imag} */,
  {32'h429e1a9c, 32'hc22872dc} /* (2, 17, 0) {real, imag} */,
  {32'hc2334536, 32'hc2268e82} /* (2, 16, 31) {real, imag} */,
  {32'hc10c637a, 32'h3e944aa0} /* (2, 16, 30) {real, imag} */,
  {32'h41b78b31, 32'hc08c2cc4} /* (2, 16, 29) {real, imag} */,
  {32'h401aa1c0, 32'h40d89d80} /* (2, 16, 28) {real, imag} */,
  {32'hc1a67f1f, 32'h41da9012} /* (2, 16, 27) {real, imag} */,
  {32'hc21d8f6c, 32'h412f8e7a} /* (2, 16, 26) {real, imag} */,
  {32'hc142ea0a, 32'h41867e0a} /* (2, 16, 25) {real, imag} */,
  {32'h41efe47c, 32'hc18c5e67} /* (2, 16, 24) {real, imag} */,
  {32'h4144a3e1, 32'hc0f0e445} /* (2, 16, 23) {real, imag} */,
  {32'hbf03c5e0, 32'h421b2b71} /* (2, 16, 22) {real, imag} */,
  {32'h4177ff2e, 32'h4132d880} /* (2, 16, 21) {real, imag} */,
  {32'hc08fda7c, 32'h403d1a24} /* (2, 16, 20) {real, imag} */,
  {32'hc11fb016, 32'hbf9a7120} /* (2, 16, 19) {real, imag} */,
  {32'h410c6980, 32'h40cbd145} /* (2, 16, 18) {real, imag} */,
  {32'hc08d928e, 32'h40f72d5a} /* (2, 16, 17) {real, imag} */,
  {32'hc037c0c0, 32'h40e494ad} /* (2, 16, 16) {real, imag} */,
  {32'hc139d611, 32'h417d8d87} /* (2, 16, 15) {real, imag} */,
  {32'h3f95ae14, 32'h3fd9919c} /* (2, 16, 14) {real, imag} */,
  {32'hc12a5e32, 32'hc1c1c261} /* (2, 16, 13) {real, imag} */,
  {32'hbee650c0, 32'hc1555d4b} /* (2, 16, 12) {real, imag} */,
  {32'hc14d2b06, 32'h405605aa} /* (2, 16, 11) {real, imag} */,
  {32'h41b94db1, 32'h410198d4} /* (2, 16, 10) {real, imag} */,
  {32'h4133885d, 32'h4182e297} /* (2, 16, 9) {real, imag} */,
  {32'hc0ea404e, 32'h41858af1} /* (2, 16, 8) {real, imag} */,
  {32'hc08f0be0, 32'hc004e262} /* (2, 16, 7) {real, imag} */,
  {32'h419dce61, 32'hc16ad602} /* (2, 16, 6) {real, imag} */,
  {32'h41eb2fb7, 32'h40cbc738} /* (2, 16, 5) {real, imag} */,
  {32'h422bbcf2, 32'h424741fe} /* (2, 16, 4) {real, imag} */,
  {32'hc1cf7133, 32'h419dbc54} /* (2, 16, 3) {real, imag} */,
  {32'hc2076392, 32'hc19de3d2} /* (2, 16, 2) {real, imag} */,
  {32'h3f9e5810, 32'h418130c1} /* (2, 16, 1) {real, imag} */,
  {32'hc2314a74, 32'hc192931c} /* (2, 16, 0) {real, imag} */,
  {32'hc1e19cca, 32'hc2202236} /* (2, 15, 31) {real, imag} */,
  {32'h41a3a000, 32'hc2178ab5} /* (2, 15, 30) {real, imag} */,
  {32'h41fa42b6, 32'h42883d44} /* (2, 15, 29) {real, imag} */,
  {32'hc0df42c0, 32'h416e89d1} /* (2, 15, 28) {real, imag} */,
  {32'h41aa9ea2, 32'hc1126878} /* (2, 15, 27) {real, imag} */,
  {32'hc24d2cc7, 32'h4113145f} /* (2, 15, 26) {real, imag} */,
  {32'h401fbeb0, 32'h410ab948} /* (2, 15, 25) {real, imag} */,
  {32'h41879a94, 32'h41269452} /* (2, 15, 24) {real, imag} */,
  {32'h41b6fad8, 32'h41d95a70} /* (2, 15, 23) {real, imag} */,
  {32'h41af9a6d, 32'h418f97ae} /* (2, 15, 22) {real, imag} */,
  {32'h41336541, 32'h3ffc9c38} /* (2, 15, 21) {real, imag} */,
  {32'h40e76244, 32'hc02cce56} /* (2, 15, 20) {real, imag} */,
  {32'hc0a8be09, 32'hc1186840} /* (2, 15, 19) {real, imag} */,
  {32'hc0916bbd, 32'h404225d7} /* (2, 15, 18) {real, imag} */,
  {32'h3fcbda30, 32'h402c4b48} /* (2, 15, 17) {real, imag} */,
  {32'hc02cbaa0, 32'hc091286b} /* (2, 15, 16) {real, imag} */,
  {32'h410a6e46, 32'hc0b992d4} /* (2, 15, 15) {real, imag} */,
  {32'hc0a266bf, 32'h408fd91c} /* (2, 15, 14) {real, imag} */,
  {32'h4041344e, 32'hc0baf1c8} /* (2, 15, 13) {real, imag} */,
  {32'h419cac00, 32'h4076f37a} /* (2, 15, 12) {real, imag} */,
  {32'h41674185, 32'h416dc099} /* (2, 15, 11) {real, imag} */,
  {32'hbf7ddfa0, 32'hc19a7406} /* (2, 15, 10) {real, imag} */,
  {32'h4153e97c, 32'hc0ad8238} /* (2, 15, 9) {real, imag} */,
  {32'hc19cef42, 32'h40d87504} /* (2, 15, 8) {real, imag} */,
  {32'h423a2378, 32'hc1d861be} /* (2, 15, 7) {real, imag} */,
  {32'hc2ad099e, 32'hc0936fd2} /* (2, 15, 6) {real, imag} */,
  {32'hc0c4d4e2, 32'h418c5fdf} /* (2, 15, 5) {real, imag} */,
  {32'h424a6ea4, 32'hc12c7503} /* (2, 15, 4) {real, imag} */,
  {32'hc110e744, 32'h420c909d} /* (2, 15, 3) {real, imag} */,
  {32'h424e3094, 32'hc22ded53} /* (2, 15, 2) {real, imag} */,
  {32'hc28b13d8, 32'hc2686974} /* (2, 15, 1) {real, imag} */,
  {32'hc231333e, 32'hc192da69} /* (2, 15, 0) {real, imag} */,
  {32'h42ed5e2c, 32'hc29de420} /* (2, 14, 31) {real, imag} */,
  {32'hc2cf0be4, 32'h42309d06} /* (2, 14, 30) {real, imag} */,
  {32'hc1fa3f1a, 32'hc245ef33} /* (2, 14, 29) {real, imag} */,
  {32'h424b4d3a, 32'h415665b0} /* (2, 14, 28) {real, imag} */,
  {32'hc241a103, 32'h40923ade} /* (2, 14, 27) {real, imag} */,
  {32'h42b231e0, 32'hc11bb2a4} /* (2, 14, 26) {real, imag} */,
  {32'h3fddb050, 32'h41d165dd} /* (2, 14, 25) {real, imag} */,
  {32'h4083a498, 32'h41a3313c} /* (2, 14, 24) {real, imag} */,
  {32'h4141b3fe, 32'hc100a0e2} /* (2, 14, 23) {real, imag} */,
  {32'hc13b8522, 32'hc06f69d9} /* (2, 14, 22) {real, imag} */,
  {32'h40a84b76, 32'hc126893a} /* (2, 14, 21) {real, imag} */,
  {32'h41a1d6a8, 32'hc09a8f90} /* (2, 14, 20) {real, imag} */,
  {32'h411acfe8, 32'h41abdf00} /* (2, 14, 19) {real, imag} */,
  {32'hc0c93737, 32'h3f31b760} /* (2, 14, 18) {real, imag} */,
  {32'h40c15c00, 32'h41400aba} /* (2, 14, 17) {real, imag} */,
  {32'h40b77698, 32'h41017d10} /* (2, 14, 16) {real, imag} */,
  {32'h41108258, 32'hc11f102a} /* (2, 14, 15) {real, imag} */,
  {32'h410aabbc, 32'hc08925b8} /* (2, 14, 14) {real, imag} */,
  {32'h40f15a48, 32'hbfa214f8} /* (2, 14, 13) {real, imag} */,
  {32'h40cd082a, 32'h3f88d3c0} /* (2, 14, 12) {real, imag} */,
  {32'h417de461, 32'hc1d5c64f} /* (2, 14, 11) {real, imag} */,
  {32'h3e27c280, 32'hc08c1b3a} /* (2, 14, 10) {real, imag} */,
  {32'hc12f97a2, 32'hc12f915e} /* (2, 14, 9) {real, imag} */,
  {32'hc162c96c, 32'hc13b8c77} /* (2, 14, 8) {real, imag} */,
  {32'h423b57ea, 32'hc10bbe92} /* (2, 14, 7) {real, imag} */,
  {32'hc1d81212, 32'h402d2b4a} /* (2, 14, 6) {real, imag} */,
  {32'hc1b537e2, 32'hc0ba9aea} /* (2, 14, 5) {real, imag} */,
  {32'h42a251fd, 32'hc2b12ff6} /* (2, 14, 4) {real, imag} */,
  {32'hc1d74ed8, 32'hc01a21d0} /* (2, 14, 3) {real, imag} */,
  {32'hc2b727d4, 32'h40d7ee10} /* (2, 14, 2) {real, imag} */,
  {32'h42bf9ba8, 32'h41988f2a} /* (2, 14, 1) {real, imag} */,
  {32'h42b8ee80, 32'h416ab05a} /* (2, 14, 0) {real, imag} */,
  {32'h3fd7c3a0, 32'hc1ebf86a} /* (2, 13, 31) {real, imag} */,
  {32'h4269bf58, 32'h4229cfc1} /* (2, 13, 30) {real, imag} */,
  {32'hc1af012f, 32'h3fdb01f4} /* (2, 13, 29) {real, imag} */,
  {32'h4124dbf4, 32'h418e3978} /* (2, 13, 28) {real, imag} */,
  {32'hc1c52af1, 32'hc156f4d8} /* (2, 13, 27) {real, imag} */,
  {32'hc147d7c5, 32'h40a5688a} /* (2, 13, 26) {real, imag} */,
  {32'h420976df, 32'hc1968840} /* (2, 13, 25) {real, imag} */,
  {32'hc11bfbee, 32'h418b2236} /* (2, 13, 24) {real, imag} */,
  {32'hc19d8fe6, 32'hbf925a28} /* (2, 13, 23) {real, imag} */,
  {32'hc084d18c, 32'hc182db12} /* (2, 13, 22) {real, imag} */,
  {32'hbecd9cc0, 32'h3fdec99c} /* (2, 13, 21) {real, imag} */,
  {32'h40c73917, 32'h40b01e1a} /* (2, 13, 20) {real, imag} */,
  {32'hc08ba44a, 32'hc0b181ff} /* (2, 13, 19) {real, imag} */,
  {32'hbf04cf80, 32'hc134fb20} /* (2, 13, 18) {real, imag} */,
  {32'hc0190918, 32'h411f43dc} /* (2, 13, 17) {real, imag} */,
  {32'h40a59fea, 32'h4032be80} /* (2, 13, 16) {real, imag} */,
  {32'h405abb88, 32'hc02d98d4} /* (2, 13, 15) {real, imag} */,
  {32'hc02baa00, 32'h41ce3f2c} /* (2, 13, 14) {real, imag} */,
  {32'hc047586c, 32'h412ea9fa} /* (2, 13, 13) {real, imag} */,
  {32'h3fe0b58c, 32'hc1d4fb50} /* (2, 13, 12) {real, imag} */,
  {32'h4118ac56, 32'h412867be} /* (2, 13, 11) {real, imag} */,
  {32'hc0819c50, 32'h40af7925} /* (2, 13, 10) {real, imag} */,
  {32'h40c1d43a, 32'hc01d8de4} /* (2, 13, 9) {real, imag} */,
  {32'h40ad8211, 32'hc1cc66da} /* (2, 13, 8) {real, imag} */,
  {32'hbff48120, 32'h428a2cf8} /* (2, 13, 7) {real, imag} */,
  {32'h41b14bf2, 32'hc1afa850} /* (2, 13, 6) {real, imag} */,
  {32'hc23a846c, 32'hc00dae3e} /* (2, 13, 5) {real, imag} */,
  {32'hc1d5883a, 32'hc21ecb61} /* (2, 13, 4) {real, imag} */,
  {32'hbfac7780, 32'hc1502be0} /* (2, 13, 3) {real, imag} */,
  {32'hc20e4f1e, 32'hc167abe4} /* (2, 13, 2) {real, imag} */,
  {32'hc21c7d97, 32'hc113550c} /* (2, 13, 1) {real, imag} */,
  {32'h41027bfb, 32'h4225661a} /* (2, 13, 0) {real, imag} */,
  {32'hc1ab62a4, 32'h42213c8a} /* (2, 12, 31) {real, imag} */,
  {32'h41b40982, 32'h427805bf} /* (2, 12, 30) {real, imag} */,
  {32'h42204db8, 32'hc2cb0d8d} /* (2, 12, 29) {real, imag} */,
  {32'hc0ca665e, 32'hc1889a34} /* (2, 12, 28) {real, imag} */,
  {32'hc1daf9d8, 32'h4224ce90} /* (2, 12, 27) {real, imag} */,
  {32'h421db3c1, 32'hc2806a92} /* (2, 12, 26) {real, imag} */,
  {32'hc21d679e, 32'hc1a80a1c} /* (2, 12, 25) {real, imag} */,
  {32'h422e814e, 32'h4080e754} /* (2, 12, 24) {real, imag} */,
  {32'h40c84b5c, 32'h3eb72958} /* (2, 12, 23) {real, imag} */,
  {32'hc18a4af6, 32'h41c51ec2} /* (2, 12, 22) {real, imag} */,
  {32'h40ef1290, 32'hc1373b0a} /* (2, 12, 21) {real, imag} */,
  {32'hc13541c5, 32'hbfe96030} /* (2, 12, 20) {real, imag} */,
  {32'hc1a30b8a, 32'hbedf8640} /* (2, 12, 19) {real, imag} */,
  {32'hbe506700, 32'h4188490a} /* (2, 12, 18) {real, imag} */,
  {32'hc14593a3, 32'hc16812a2} /* (2, 12, 17) {real, imag} */,
  {32'hbee326a0, 32'h4108a782} /* (2, 12, 16) {real, imag} */,
  {32'hc091b126, 32'hc0fca8c5} /* (2, 12, 15) {real, imag} */,
  {32'hc1005a66, 32'hc18b997e} /* (2, 12, 14) {real, imag} */,
  {32'h4193eb3e, 32'h413aedce} /* (2, 12, 13) {real, imag} */,
  {32'hc19e9020, 32'hc173ed3c} /* (2, 12, 12) {real, imag} */,
  {32'h4128b3b2, 32'h41746ab6} /* (2, 12, 11) {real, imag} */,
  {32'hc15cc9ad, 32'h42277931} /* (2, 12, 10) {real, imag} */,
  {32'h416fa592, 32'hc0cb4ac0} /* (2, 12, 9) {real, imag} */,
  {32'h425d92be, 32'hc267b706} /* (2, 12, 8) {real, imag} */,
  {32'hc050fca8, 32'hbfedfb68} /* (2, 12, 7) {real, imag} */,
  {32'h421f481d, 32'hc1fbad7e} /* (2, 12, 6) {real, imag} */,
  {32'hc185177c, 32'hc2873e2c} /* (2, 12, 5) {real, imag} */,
  {32'hc1782abd, 32'hc2292714} /* (2, 12, 4) {real, imag} */,
  {32'hc22447cc, 32'h42b9c513} /* (2, 12, 3) {real, imag} */,
  {32'hc168bfc4, 32'hc20b29d9} /* (2, 12, 2) {real, imag} */,
  {32'h418dbb10, 32'h424edcce} /* (2, 12, 1) {real, imag} */,
  {32'hc1cefb2e, 32'h40c52ea4} /* (2, 12, 0) {real, imag} */,
  {32'h43142643, 32'hc2fd49c0} /* (2, 11, 31) {real, imag} */,
  {32'hc2fe1270, 32'h431ed873} /* (2, 11, 30) {real, imag} */,
  {32'h4023e340, 32'h4277a786} /* (2, 11, 29) {real, imag} */,
  {32'hc23f1ee5, 32'h421c0493} /* (2, 11, 28) {real, imag} */,
  {32'hc15a71d2, 32'hc18c84fc} /* (2, 11, 27) {real, imag} */,
  {32'h42813fec, 32'h42427f08} /* (2, 11, 26) {real, imag} */,
  {32'h42103c38, 32'h40ea89a0} /* (2, 11, 25) {real, imag} */,
  {32'hc08def00, 32'hc1910a5c} /* (2, 11, 24) {real, imag} */,
  {32'h42305ead, 32'hc229fd46} /* (2, 11, 23) {real, imag} */,
  {32'h419161e5, 32'hc169e697} /* (2, 11, 22) {real, imag} */,
  {32'hc102d655, 32'h4210971c} /* (2, 11, 21) {real, imag} */,
  {32'hc1c39266, 32'h414c57b0} /* (2, 11, 20) {real, imag} */,
  {32'hc1b2fa69, 32'hc1976b8d} /* (2, 11, 19) {real, imag} */,
  {32'h41943a03, 32'hc1b19f74} /* (2, 11, 18) {real, imag} */,
  {32'h3fa159d0, 32'h4062bc10} /* (2, 11, 17) {real, imag} */,
  {32'hc0e8ae80, 32'hc14c01e0} /* (2, 11, 16) {real, imag} */,
  {32'h414e8726, 32'h40c2d7d8} /* (2, 11, 15) {real, imag} */,
  {32'h402c17e8, 32'h41f8d454} /* (2, 11, 14) {real, imag} */,
  {32'h411a6802, 32'hc165c86e} /* (2, 11, 13) {real, imag} */,
  {32'hc1b214c2, 32'h41c69456} /* (2, 11, 12) {real, imag} */,
  {32'hc1bcbc84, 32'hc2680c92} /* (2, 11, 11) {real, imag} */,
  {32'h42289506, 32'h3d11a500} /* (2, 11, 10) {real, imag} */,
  {32'hc217dfa5, 32'h42911108} /* (2, 11, 9) {real, imag} */,
  {32'h40ff78c0, 32'h41d1d204} /* (2, 11, 8) {real, imag} */,
  {32'h4067e5c0, 32'hc22691ce} /* (2, 11, 7) {real, imag} */,
  {32'h42087ba0, 32'hc18d4d40} /* (2, 11, 6) {real, imag} */,
  {32'hc21a4298, 32'hc10ac690} /* (2, 11, 5) {real, imag} */,
  {32'hc18591ee, 32'hc1f35683} /* (2, 11, 4) {real, imag} */,
  {32'hc2b1fdbe, 32'h426f4b50} /* (2, 11, 3) {real, imag} */,
  {32'hc35abadc, 32'hc2d3deda} /* (2, 11, 2) {real, imag} */,
  {32'h437f268b, 32'hc0d725a8} /* (2, 11, 1) {real, imag} */,
  {32'h4389ce5d, 32'hc3778516} /* (2, 11, 0) {real, imag} */,
  {32'hc34aff5e, 32'h4281f45c} /* (2, 10, 31) {real, imag} */,
  {32'h42f391fb, 32'hc15bc58b} /* (2, 10, 30) {real, imag} */,
  {32'hc1e0982b, 32'h42e47be9} /* (2, 10, 29) {real, imag} */,
  {32'h41d3c7de, 32'h4246efe6} /* (2, 10, 28) {real, imag} */,
  {32'h41869264, 32'hc2a18892} /* (2, 10, 27) {real, imag} */,
  {32'h41fdd627, 32'h426013e4} /* (2, 10, 26) {real, imag} */,
  {32'hbf8ef1ac, 32'hc159de60} /* (2, 10, 25) {real, imag} */,
  {32'h4255b0d7, 32'hc1954fd2} /* (2, 10, 24) {real, imag} */,
  {32'hc260d6da, 32'h4220df5a} /* (2, 10, 23) {real, imag} */,
  {32'hbfea4c20, 32'h424c9420} /* (2, 10, 22) {real, imag} */,
  {32'hc216e702, 32'hc1a2d40e} /* (2, 10, 21) {real, imag} */,
  {32'hc19af9fa, 32'hc1d53585} /* (2, 10, 20) {real, imag} */,
  {32'h41c8d53f, 32'hc1d11e9c} /* (2, 10, 19) {real, imag} */,
  {32'h41c0c61b, 32'hc12032ca} /* (2, 10, 18) {real, imag} */,
  {32'hc1bdc029, 32'h419d826d} /* (2, 10, 17) {real, imag} */,
  {32'hc1aec4c2, 32'h3f444240} /* (2, 10, 16) {real, imag} */,
  {32'hc1e9fdbf, 32'hc1769b22} /* (2, 10, 15) {real, imag} */,
  {32'h41073b3a, 32'hc092f108} /* (2, 10, 14) {real, imag} */,
  {32'h41ecc631, 32'hc1b38fcc} /* (2, 10, 13) {real, imag} */,
  {32'hc24553db, 32'h40e65624} /* (2, 10, 12) {real, imag} */,
  {32'h4024c698, 32'h42100391} /* (2, 10, 11) {real, imag} */,
  {32'h42aa2bec, 32'hc2018c54} /* (2, 10, 10) {real, imag} */,
  {32'h42350a76, 32'h427b559a} /* (2, 10, 9) {real, imag} */,
  {32'hc24a2445, 32'h421760e7} /* (2, 10, 8) {real, imag} */,
  {32'h415bbe62, 32'h42ddf52c} /* (2, 10, 7) {real, imag} */,
  {32'h422292d6, 32'hc266c934} /* (2, 10, 6) {real, imag} */,
  {32'h3e391ac0, 32'h41cd0e9e} /* (2, 10, 5) {real, imag} */,
  {32'hc2ba2af8, 32'hc23be002} /* (2, 10, 4) {real, imag} */,
  {32'hc0b536f4, 32'hc24c774e} /* (2, 10, 3) {real, imag} */,
  {32'h432f0482, 32'hc1daf4d2} /* (2, 10, 2) {real, imag} */,
  {32'hc2baa7d5, 32'h4327cda6} /* (2, 10, 1) {real, imag} */,
  {32'hc20f9265, 32'h425f01b5} /* (2, 10, 0) {real, imag} */,
  {32'hc2f8a35a, 32'hc35f6d6a} /* (2, 9, 31) {real, imag} */,
  {32'h433fd624, 32'h432a173e} /* (2, 9, 30) {real, imag} */,
  {32'hc29015e6, 32'h42ab9c58} /* (2, 9, 29) {real, imag} */,
  {32'hc21c96d7, 32'h41bdd2e2} /* (2, 9, 28) {real, imag} */,
  {32'h4199915c, 32'hc3359284} /* (2, 9, 27) {real, imag} */,
  {32'h426bfe36, 32'h41d8d551} /* (2, 9, 26) {real, imag} */,
  {32'h41ce223e, 32'h4217bfcc} /* (2, 9, 25) {real, imag} */,
  {32'h4241bf96, 32'hc26776c6} /* (2, 9, 24) {real, imag} */,
  {32'hc24c4c6f, 32'h424c36e2} /* (2, 9, 23) {real, imag} */,
  {32'hc1100568, 32'hc16480a2} /* (2, 9, 22) {real, imag} */,
  {32'h409fd91e, 32'hc1e670be} /* (2, 9, 21) {real, imag} */,
  {32'h4172a2c0, 32'hc2175f02} /* (2, 9, 20) {real, imag} */,
  {32'hc07f0694, 32'h421ae0b2} /* (2, 9, 19) {real, imag} */,
  {32'h422d80e2, 32'hc1a1496e} /* (2, 9, 18) {real, imag} */,
  {32'h416ff52b, 32'hc2005432} /* (2, 9, 17) {real, imag} */,
  {32'hc1730038, 32'h41672c50} /* (2, 9, 16) {real, imag} */,
  {32'h410ecd4d, 32'h410bf496} /* (2, 9, 15) {real, imag} */,
  {32'hc20c1f7e, 32'h40e1d778} /* (2, 9, 14) {real, imag} */,
  {32'h41c3632e, 32'h41699866} /* (2, 9, 13) {real, imag} */,
  {32'hc199486c, 32'hc019d0c8} /* (2, 9, 12) {real, imag} */,
  {32'hc1c7aa18, 32'h417ab444} /* (2, 9, 11) {real, imag} */,
  {32'hc28e002f, 32'hc25c61a8} /* (2, 9, 10) {real, imag} */,
  {32'h426f050b, 32'hc1d67fb1} /* (2, 9, 9) {real, imag} */,
  {32'hc15aed62, 32'h41140442} /* (2, 9, 8) {real, imag} */,
  {32'hc20a5f27, 32'hc24c0c1a} /* (2, 9, 7) {real, imag} */,
  {32'h4178b5e8, 32'hc1592062} /* (2, 9, 6) {real, imag} */,
  {32'hc2abb5f9, 32'hc2237ff0} /* (2, 9, 5) {real, imag} */,
  {32'hc2873486, 32'hc2170552} /* (2, 9, 4) {real, imag} */,
  {32'hc20fb737, 32'hc1e857b9} /* (2, 9, 3) {real, imag} */,
  {32'h42ad8888, 32'h42e01ff8} /* (2, 9, 2) {real, imag} */,
  {32'hc29451ae, 32'h433904e8} /* (2, 9, 1) {real, imag} */,
  {32'h424aa00c, 32'hc20d744b} /* (2, 9, 0) {real, imag} */,
  {32'h43b5c157, 32'hc4112adc} /* (2, 8, 31) {real, imag} */,
  {32'hc33f0c4f, 32'h43d06838} /* (2, 8, 30) {real, imag} */,
  {32'h4253555f, 32'hc2d7e9f8} /* (2, 8, 29) {real, imag} */,
  {32'h3fd68a80, 32'h41c91c40} /* (2, 8, 28) {real, imag} */,
  {32'hc1f8c5b4, 32'h42870e92} /* (2, 8, 27) {real, imag} */,
  {32'hc2ea0d5d, 32'h41bdcb7a} /* (2, 8, 26) {real, imag} */,
  {32'h42ff5bea, 32'h41902a48} /* (2, 8, 25) {real, imag} */,
  {32'hc2ab5d06, 32'h43101e94} /* (2, 8, 24) {real, imag} */,
  {32'h4284f416, 32'h41a8a870} /* (2, 8, 23) {real, imag} */,
  {32'hc22c508c, 32'hc18f452a} /* (2, 8, 22) {real, imag} */,
  {32'h41ee1014, 32'h4227141c} /* (2, 8, 21) {real, imag} */,
  {32'hc2075e9c, 32'h41c401de} /* (2, 8, 20) {real, imag} */,
  {32'h40a198ea, 32'hc1bff2a4} /* (2, 8, 19) {real, imag} */,
  {32'h41d07c40, 32'h414c796c} /* (2, 8, 18) {real, imag} */,
  {32'hbf307700, 32'h413181b0} /* (2, 8, 17) {real, imag} */,
  {32'hc1feae98, 32'h41cd6df6} /* (2, 8, 16) {real, imag} */,
  {32'h4186fbd8, 32'hc1c53c18} /* (2, 8, 15) {real, imag} */,
  {32'h4121f701, 32'h4155b7d4} /* (2, 8, 14) {real, imag} */,
  {32'hc16a6c9b, 32'h3f5db2f0} /* (2, 8, 13) {real, imag} */,
  {32'hc1e0cc30, 32'h40c0fdf8} /* (2, 8, 12) {real, imag} */,
  {32'hc231212e, 32'h4168aaa7} /* (2, 8, 11) {real, imag} */,
  {32'hc0d429a0, 32'h4155b45c} /* (2, 8, 10) {real, imag} */,
  {32'h426798c5, 32'hc1e44078} /* (2, 8, 9) {real, imag} */,
  {32'h42a58fd0, 32'h40dd5e80} /* (2, 8, 8) {real, imag} */,
  {32'hc2eb7692, 32'h4266dbe0} /* (2, 8, 7) {real, imag} */,
  {32'h3e520e00, 32'hc0c633b8} /* (2, 8, 6) {real, imag} */,
  {32'hc2576e3e, 32'h4315dee9} /* (2, 8, 5) {real, imag} */,
  {32'h42accfc2, 32'hc3273daa} /* (2, 8, 4) {real, imag} */,
  {32'hc2eebe20, 32'h428f2050} /* (2, 8, 3) {real, imag} */,
  {32'hc3152f81, 32'h4351d054} /* (2, 8, 2) {real, imag} */,
  {32'h43901023, 32'hc3243157} /* (2, 8, 1) {real, imag} */,
  {32'h433dd339, 32'hc30f6562} /* (2, 8, 0) {real, imag} */,
  {32'hc18db408, 32'h432b26e5} /* (2, 7, 31) {real, imag} */,
  {32'h42e81867, 32'hc2ba0e5a} /* (2, 7, 30) {real, imag} */,
  {32'hc228be51, 32'h3e802000} /* (2, 7, 29) {real, imag} */,
  {32'hc1ed21cf, 32'hc1141120} /* (2, 7, 28) {real, imag} */,
  {32'h4219960b, 32'hc29064a5} /* (2, 7, 27) {real, imag} */,
  {32'h41612a03, 32'hc1c7ca80} /* (2, 7, 26) {real, imag} */,
  {32'hc26e6242, 32'hc11d2530} /* (2, 7, 25) {real, imag} */,
  {32'h425e6638, 32'hc0e42340} /* (2, 7, 24) {real, imag} */,
  {32'h42c6f857, 32'h4178de30} /* (2, 7, 23) {real, imag} */,
  {32'hc0f37354, 32'hc1c0124e} /* (2, 7, 22) {real, imag} */,
  {32'h41e8bc02, 32'h42bbabb6} /* (2, 7, 21) {real, imag} */,
  {32'hc207c762, 32'hc1189ea6} /* (2, 7, 20) {real, imag} */,
  {32'hc009e154, 32'h41e5af00} /* (2, 7, 19) {real, imag} */,
  {32'hc24bebae, 32'hc15dc0aa} /* (2, 7, 18) {real, imag} */,
  {32'h3fb90060, 32'hc1555f3c} /* (2, 7, 17) {real, imag} */,
  {32'hc0a4c510, 32'h411eb480} /* (2, 7, 16) {real, imag} */,
  {32'h41d01222, 32'h4175274c} /* (2, 7, 15) {real, imag} */,
  {32'hbf6d9400, 32'h41dbe4c7} /* (2, 7, 14) {real, imag} */,
  {32'h4060bb3c, 32'hc168b740} /* (2, 7, 13) {real, imag} */,
  {32'h41c1445a, 32'h41b16f34} /* (2, 7, 12) {real, imag} */,
  {32'h425457e3, 32'h4286bd30} /* (2, 7, 11) {real, imag} */,
  {32'h41866b04, 32'h41bde736} /* (2, 7, 10) {real, imag} */,
  {32'hc1a827f4, 32'hc280c9ae} /* (2, 7, 9) {real, imag} */,
  {32'h415594f0, 32'hc284e04c} /* (2, 7, 8) {real, imag} */,
  {32'hc1284eb8, 32'h43325ac3} /* (2, 7, 7) {real, imag} */,
  {32'hc22d6c51, 32'hc155f5e7} /* (2, 7, 6) {real, imag} */,
  {32'h428c1f8c, 32'hc2ae5ab1} /* (2, 7, 5) {real, imag} */,
  {32'hc2700f04, 32'hc0630dc6} /* (2, 7, 4) {real, imag} */,
  {32'h4298b422, 32'hc3550ebe} /* (2, 7, 3) {real, imag} */,
  {32'h4287b135, 32'hc1ab2952} /* (2, 7, 2) {real, imag} */,
  {32'hc36fd513, 32'h4302e5ff} /* (2, 7, 1) {real, imag} */,
  {32'hc2e43bf9, 32'h432e1050} /* (2, 7, 0) {real, imag} */,
  {32'h428fd7fc, 32'h426c843d} /* (2, 6, 31) {real, imag} */,
  {32'hc2995c37, 32'h42ec7520} /* (2, 6, 30) {real, imag} */,
  {32'h41ac1bce, 32'hc2684065} /* (2, 6, 29) {real, imag} */,
  {32'hc2746029, 32'h4265aafd} /* (2, 6, 28) {real, imag} */,
  {32'hc284ce94, 32'hc27cf65a} /* (2, 6, 27) {real, imag} */,
  {32'hc2716d2a, 32'h41770220} /* (2, 6, 26) {real, imag} */,
  {32'hc155c86a, 32'hc21b2191} /* (2, 6, 25) {real, imag} */,
  {32'hc2a1a9c2, 32'h4230456c} /* (2, 6, 24) {real, imag} */,
  {32'hc15a81ee, 32'h404eac50} /* (2, 6, 23) {real, imag} */,
  {32'h40deb9fc, 32'h41af409c} /* (2, 6, 22) {real, imag} */,
  {32'hc23fa2d1, 32'h425273bc} /* (2, 6, 21) {real, imag} */,
  {32'hc1460155, 32'h41fccf56} /* (2, 6, 20) {real, imag} */,
  {32'h41e620cb, 32'hc0905a47} /* (2, 6, 19) {real, imag} */,
  {32'h40d320e2, 32'hc0809e1a} /* (2, 6, 18) {real, imag} */,
  {32'h40923857, 32'hc14fc5cc} /* (2, 6, 17) {real, imag} */,
  {32'hc19adb9e, 32'h410dd4fc} /* (2, 6, 16) {real, imag} */,
  {32'h413c6d3c, 32'h40a11078} /* (2, 6, 15) {real, imag} */,
  {32'h414b11b9, 32'hc2080739} /* (2, 6, 14) {real, imag} */,
  {32'hc265ba30, 32'h419dc17a} /* (2, 6, 13) {real, imag} */,
  {32'h416e8b67, 32'hc1d35656} /* (2, 6, 12) {real, imag} */,
  {32'hc185d116, 32'h423171f8} /* (2, 6, 11) {real, imag} */,
  {32'h40f0e514, 32'hc2c39b07} /* (2, 6, 10) {real, imag} */,
  {32'h426cb950, 32'h42305eb5} /* (2, 6, 9) {real, imag} */,
  {32'hc23ea4b8, 32'h42caf836} /* (2, 6, 8) {real, imag} */,
  {32'h4257e242, 32'hc1d5bb02} /* (2, 6, 7) {real, imag} */,
  {32'hc291d2e7, 32'h429c6dfa} /* (2, 6, 6) {real, imag} */,
  {32'h420778c7, 32'h424cce52} /* (2, 6, 5) {real, imag} */,
  {32'h41aa2fde, 32'h422c441f} /* (2, 6, 4) {real, imag} */,
  {32'hc2c53ab4, 32'h42841f25} /* (2, 6, 3) {real, imag} */,
  {32'h42e4231d, 32'h433dd510} /* (2, 6, 2) {real, imag} */,
  {32'h4266f9b8, 32'hc29fe056} /* (2, 6, 1) {real, imag} */,
  {32'hc29dea26, 32'hc28c6068} /* (2, 6, 0) {real, imag} */,
  {32'h439c9aa8, 32'hc44bda3a} /* (2, 5, 31) {real, imag} */,
  {32'hc29e0562, 32'h439b9fa6} /* (2, 5, 30) {real, imag} */,
  {32'hc1a9bbf8, 32'h42dd3276} /* (2, 5, 29) {real, imag} */,
  {32'hc31f9d65, 32'hc2edf1db} /* (2, 5, 28) {real, imag} */,
  {32'h42e0f64a, 32'h438c2b24} /* (2, 5, 27) {real, imag} */,
  {32'h428932ca, 32'h42077585} /* (2, 5, 26) {real, imag} */,
  {32'hc212f7f6, 32'hc04bfca8} /* (2, 5, 25) {real, imag} */,
  {32'h42672788, 32'h42f41657} /* (2, 5, 24) {real, imag} */,
  {32'hc25e3f3a, 32'hc186429b} /* (2, 5, 23) {real, imag} */,
  {32'h4218b85e, 32'h42acb31a} /* (2, 5, 22) {real, imag} */,
  {32'h41b72698, 32'h431ad7da} /* (2, 5, 21) {real, imag} */,
  {32'hc1fe53be, 32'h40337970} /* (2, 5, 20) {real, imag} */,
  {32'hc2120d2e, 32'hc13361f0} /* (2, 5, 19) {real, imag} */,
  {32'h426a980e, 32'h42460022} /* (2, 5, 18) {real, imag} */,
  {32'h423659b8, 32'h411533f8} /* (2, 5, 17) {real, imag} */,
  {32'h411c84f0, 32'h40c7ad40} /* (2, 5, 16) {real, imag} */,
  {32'hc2050210, 32'hc201c9be} /* (2, 5, 15) {real, imag} */,
  {32'hc1d8253c, 32'hc23a27f6} /* (2, 5, 14) {real, imag} */,
  {32'h41e24444, 32'hc1c47288} /* (2, 5, 13) {real, imag} */,
  {32'hc20d1eef, 32'h42838256} /* (2, 5, 12) {real, imag} */,
  {32'hc2e95f5e, 32'h41b4b37c} /* (2, 5, 11) {real, imag} */,
  {32'hc0d461d8, 32'hc29c1cd8} /* (2, 5, 10) {real, imag} */,
  {32'h419b2f0c, 32'h4265f546} /* (2, 5, 9) {real, imag} */,
  {32'hc308d338, 32'h42a0bc11} /* (2, 5, 8) {real, imag} */,
  {32'h42872f95, 32'h4080750c} /* (2, 5, 7) {real, imag} */,
  {32'hc2abd1c8, 32'hc2e3a448} /* (2, 5, 6) {real, imag} */,
  {32'hc3c4e768, 32'h43a726d8} /* (2, 5, 5) {real, imag} */,
  {32'h431a14bd, 32'hc2e80a69} /* (2, 5, 4) {real, imag} */,
  {32'h42ad02e2, 32'hc20044f4} /* (2, 5, 3) {real, imag} */,
  {32'hc324119d, 32'h4290588e} /* (2, 5, 2) {real, imag} */,
  {32'h44073fac, 32'hc3fd65db} /* (2, 5, 1) {real, imag} */,
  {32'h43b3e0ba, 32'hc40d0ebe} /* (2, 5, 0) {real, imag} */,
  {32'hc4142e20, 32'h43478754} /* (2, 4, 31) {real, imag} */,
  {32'h44075289, 32'hc3d781f0} /* (2, 4, 30) {real, imag} */,
  {32'h41238644, 32'hc1e94cc4} /* (2, 4, 29) {real, imag} */,
  {32'hc2b81cbb, 32'h43b18e05} /* (2, 4, 28) {real, imag} */,
  {32'hc2902c7b, 32'hc34257ba} /* (2, 4, 27) {real, imag} */,
  {32'hc30e7f8e, 32'h42b71bd9} /* (2, 4, 26) {real, imag} */,
  {32'hc28ecc47, 32'h40b5bd00} /* (2, 4, 25) {real, imag} */,
  {32'hc0d46fa0, 32'hc30187a7} /* (2, 4, 24) {real, imag} */,
  {32'hc2a80881, 32'h42969d7c} /* (2, 4, 23) {real, imag} */,
  {32'h4224a7d6, 32'h42ccc689} /* (2, 4, 22) {real, imag} */,
  {32'hc2aadc0e, 32'hc33571c0} /* (2, 4, 21) {real, imag} */,
  {32'h422fdbb0, 32'hc14d24f8} /* (2, 4, 20) {real, imag} */,
  {32'h3f267730, 32'hc009e340} /* (2, 4, 19) {real, imag} */,
  {32'h415a3cdc, 32'hc14915ec} /* (2, 4, 18) {real, imag} */,
  {32'hc283681b, 32'h40fd2080} /* (2, 4, 17) {real, imag} */,
  {32'h41b8f010, 32'hc1c0fc28} /* (2, 4, 16) {real, imag} */,
  {32'h41c00a6c, 32'hc20ce950} /* (2, 4, 15) {real, imag} */,
  {32'h422c9ae9, 32'h40859458} /* (2, 4, 14) {real, imag} */,
  {32'h40cd5ada, 32'h421455c8} /* (2, 4, 13) {real, imag} */,
  {32'h42b9fad0, 32'hc244051a} /* (2, 4, 12) {real, imag} */,
  {32'hc0426530, 32'hc08e0bb0} /* (2, 4, 11) {real, imag} */,
  {32'hc28aa077, 32'hc2391356} /* (2, 4, 10) {real, imag} */,
  {32'h41f3947c, 32'h412eb710} /* (2, 4, 9) {real, imag} */,
  {32'h4324bb09, 32'h407beed0} /* (2, 4, 8) {real, imag} */,
  {32'hc10807ba, 32'h42bbc9fa} /* (2, 4, 7) {real, imag} */,
  {32'h406d4e20, 32'hc28c759b} /* (2, 4, 6) {real, imag} */,
  {32'h4336ef7a, 32'h4279dcce} /* (2, 4, 5) {real, imag} */,
  {32'hc372ce66, 32'h4300ffd4} /* (2, 4, 4) {real, imag} */,
  {32'hc236d12d, 32'h42f166d7} /* (2, 4, 3) {real, imag} */,
  {32'h44263759, 32'hc3e8793e} /* (2, 4, 2) {real, imag} */,
  {32'hc3f06a2b, 32'h4480ec20} /* (2, 4, 1) {real, imag} */,
  {32'hc2ccc3d9, 32'h434b0f31} /* (2, 4, 0) {real, imag} */,
  {32'hc335e400, 32'hc4344a9b} /* (2, 3, 31) {real, imag} */,
  {32'h440b30b7, 32'h443bec5e} /* (2, 3, 30) {real, imag} */,
  {32'hc2a96350, 32'hc0c90cd0} /* (2, 3, 29) {real, imag} */,
  {32'hc38652ad, 32'h438ee5df} /* (2, 3, 28) {real, imag} */,
  {32'h425be0f6, 32'hc37cc279} /* (2, 3, 27) {real, imag} */,
  {32'hc2e6903b, 32'h41a7a94a} /* (2, 3, 26) {real, imag} */,
  {32'hc047e840, 32'h4306bf7d} /* (2, 3, 25) {real, imag} */,
  {32'h43148a29, 32'h401ff6c0} /* (2, 3, 24) {real, imag} */,
  {32'hc314d4f1, 32'h427311a9} /* (2, 3, 23) {real, imag} */,
  {32'hc31025b4, 32'h4277ac0b} /* (2, 3, 22) {real, imag} */,
  {32'hc2239768, 32'hc2c2bb68} /* (2, 3, 21) {real, imag} */,
  {32'hc1935bd4, 32'hc16cab7c} /* (2, 3, 20) {real, imag} */,
  {32'hc108beee, 32'hc246e10e} /* (2, 3, 19) {real, imag} */,
  {32'hc0f16c38, 32'h40835300} /* (2, 3, 18) {real, imag} */,
  {32'hbf8dd180, 32'hc186e470} /* (2, 3, 17) {real, imag} */,
  {32'hc2777611, 32'h4093b554} /* (2, 3, 16) {real, imag} */,
  {32'h40e9bca0, 32'hc05fb680} /* (2, 3, 15) {real, imag} */,
  {32'h428cf004, 32'h4153c000} /* (2, 3, 14) {real, imag} */,
  {32'h41f78b43, 32'h417896a8} /* (2, 3, 13) {real, imag} */,
  {32'h41934b14, 32'h415f4074} /* (2, 3, 12) {real, imag} */,
  {32'hc238b2a0, 32'h42edc01c} /* (2, 3, 11) {real, imag} */,
  {32'h428d4bef, 32'hc2efb46c} /* (2, 3, 10) {real, imag} */,
  {32'hc2180585, 32'hc287be34} /* (2, 3, 9) {real, imag} */,
  {32'h4318fe81, 32'hc1c77a6a} /* (2, 3, 8) {real, imag} */,
  {32'hc2605cc2, 32'h42848912} /* (2, 3, 7) {real, imag} */,
  {32'hc2b355fb, 32'hc3030ae2} /* (2, 3, 6) {real, imag} */,
  {32'hc3218b7a, 32'h4364fb5d} /* (2, 3, 5) {real, imag} */,
  {32'hc2161dc2, 32'hc26bed58} /* (2, 3, 4) {real, imag} */,
  {32'hc1db2dc5, 32'hc2e4cca9} /* (2, 3, 3) {real, imag} */,
  {32'h44352fb9, 32'h413b9de0} /* (2, 3, 2) {real, imag} */,
  {32'hc3f400a4, 32'h439df32a} /* (2, 3, 1) {real, imag} */,
  {32'hc2829084, 32'hc2084102} /* (2, 3, 0) {real, imag} */,
  {32'h44504766, 32'hc552372c} /* (2, 2, 31) {real, imag} */,
  {32'h434e8cc1, 32'h4507abd6} /* (2, 2, 30) {real, imag} */,
  {32'h43111e9e, 32'hc208e9f5} /* (2, 2, 29) {real, imag} */,
  {32'hc4166c53, 32'hc3a100cd} /* (2, 2, 28) {real, imag} */,
  {32'h433b54cc, 32'h4436aff8} /* (2, 2, 27) {real, imag} */,
  {32'h4251e8b6, 32'h4344ec63} /* (2, 2, 26) {real, imag} */,
  {32'hc384c80a, 32'hc39a4332} /* (2, 2, 25) {real, imag} */,
  {32'h438674f9, 32'h43504f33} /* (2, 2, 24) {real, imag} */,
  {32'hc2c692e9, 32'h428a3f12} /* (2, 2, 23) {real, imag} */,
  {32'hc21ab112, 32'h4097bb28} /* (2, 2, 22) {real, imag} */,
  {32'h43347ee8, 32'h432d5de8} /* (2, 2, 21) {real, imag} */,
  {32'hc28cc899, 32'hc29e415d} /* (2, 2, 20) {real, imag} */,
  {32'hc1fe1406, 32'h40aa9ec8} /* (2, 2, 19) {real, imag} */,
  {32'h429da34d, 32'h428e0c74} /* (2, 2, 18) {real, imag} */,
  {32'hc28a6250, 32'h3f837700} /* (2, 2, 17) {real, imag} */,
  {32'h416c4f00, 32'hc2104af0} /* (2, 2, 16) {real, imag} */,
  {32'hc113da80, 32'hc289f61c} /* (2, 2, 15) {real, imag} */,
  {32'hc2c516ff, 32'h414ef660} /* (2, 2, 14) {real, imag} */,
  {32'h40cf13b8, 32'h3fc3a6e0} /* (2, 2, 13) {real, imag} */,
  {32'h41897b3c, 32'h41aae894} /* (2, 2, 12) {real, imag} */,
  {32'hc34c73bc, 32'h4249b7f0} /* (2, 2, 11) {real, imag} */,
  {32'h4260e2c8, 32'hc2df0af2} /* (2, 2, 10) {real, imag} */,
  {32'hc1d374dc, 32'hc299c1c2} /* (2, 2, 9) {real, imag} */,
  {32'hc35437c8, 32'h432472d9} /* (2, 2, 8) {real, imag} */,
  {32'h417d2340, 32'hc2d3eac6} /* (2, 2, 7) {real, imag} */,
  {32'hc229c644, 32'h42cef88a} /* (2, 2, 6) {real, imag} */,
  {32'hc42d0160, 32'h43a7ebff} /* (2, 2, 5) {real, imag} */,
  {32'h440941cd, 32'hc44371a2} /* (2, 2, 4) {real, imag} */,
  {32'h427f2855, 32'hc26102bb} /* (2, 2, 3) {real, imag} */,
  {32'h42f4924e, 32'h44d88acc} /* (2, 2, 2) {real, imag} */,
  {32'hc1d752c0, 32'hc502118c} /* (2, 2, 1) {real, imag} */,
  {32'h440b7060, 32'hc4a7e604} /* (2, 2, 0) {real, imag} */,
  {32'h42f86750, 32'h4529b903} /* (2, 1, 31) {real, imag} */,
  {32'h42ee0e68, 32'hc4aaae7a} /* (2, 1, 30) {real, imag} */,
  {32'hc33a276d, 32'h40a08ef0} /* (2, 1, 29) {real, imag} */,
  {32'hc3dc86e2, 32'h4398e014} /* (2, 1, 28) {real, imag} */,
  {32'h4363816a, 32'hc4718c38} /* (2, 1, 27) {real, imag} */,
  {32'h43112d04, 32'hc374f8a7} /* (2, 1, 26) {real, imag} */,
  {32'h42939891, 32'h43478352} /* (2, 1, 25) {real, imag} */,
  {32'hc30f74cd, 32'hc3558e1b} /* (2, 1, 24) {real, imag} */,
  {32'hc336faf0, 32'hc30dc6d2} /* (2, 1, 23) {real, imag} */,
  {32'hc2d77f44, 32'h42a65fbe} /* (2, 1, 22) {real, imag} */,
  {32'hc283d576, 32'hc38f4012} /* (2, 1, 21) {real, imag} */,
  {32'hc1ecedd8, 32'h40f741c0} /* (2, 1, 20) {real, imag} */,
  {32'hc1dffb5c, 32'h4234aa0a} /* (2, 1, 19) {real, imag} */,
  {32'hc2c8dfec, 32'hbf3cdfc0} /* (2, 1, 18) {real, imag} */,
  {32'hbeed0800, 32'hc1183ac0} /* (2, 1, 17) {real, imag} */,
  {32'hc1f495a0, 32'hbeb71000} /* (2, 1, 16) {real, imag} */,
  {32'hc12599c0, 32'hc214ded0} /* (2, 1, 15) {real, imag} */,
  {32'h42daa5dc, 32'h42880f20} /* (2, 1, 14) {real, imag} */,
  {32'hc24a1bc6, 32'h42e92971} /* (2, 1, 13) {real, imag} */,
  {32'h4285ba76, 32'h40122200} /* (2, 1, 12) {real, imag} */,
  {32'h43348aa9, 32'hc1935440} /* (2, 1, 11) {real, imag} */,
  {32'h4303e908, 32'hc2ba4ae6} /* (2, 1, 10) {real, imag} */,
  {32'h40f683f0, 32'h4190f330} /* (2, 1, 9) {real, imag} */,
  {32'h44000f56, 32'hc28d6e6a} /* (2, 1, 8) {real, imag} */,
  {32'hc35cb168, 32'h42b74614} /* (2, 1, 7) {real, imag} */,
  {32'h42ff04f4, 32'hc149e850} /* (2, 1, 6) {real, imag} */,
  {32'h44034d8e, 32'hc40bc240} /* (2, 1, 5) {real, imag} */,
  {32'hc3e05324, 32'h435ea849} /* (2, 1, 4) {real, imag} */,
  {32'hc314915b, 32'hc313d34a} /* (2, 1, 3) {real, imag} */,
  {32'h44ea9d8c, 32'hc4a27ae8} /* (2, 1, 2) {real, imag} */,
  {32'hc535cd5e, 32'h4550e473} /* (2, 1, 1) {real, imag} */,
  {32'hc444fd2f, 32'h45165d50} /* (2, 1, 0) {real, imag} */,
  {32'h4470e104, 32'h44ec0e8e} /* (2, 0, 31) {real, imag} */,
  {32'hc435d57c, 32'hc4207178} /* (2, 0, 30) {real, imag} */,
  {32'h41155278, 32'hc32e916b} /* (2, 0, 29) {real, imag} */,
  {32'hc3e057a2, 32'h41c906de} /* (2, 0, 28) {real, imag} */,
  {32'h42bef660, 32'hc4027b6e} /* (2, 0, 27) {real, imag} */,
  {32'hc1cc0ed0, 32'hc2fda7a9} /* (2, 0, 26) {real, imag} */,
  {32'h429edf80, 32'h4279e11a} /* (2, 0, 25) {real, imag} */,
  {32'hc3636826, 32'hc16d7678} /* (2, 0, 24) {real, imag} */,
  {32'h4108f680, 32'hc2b9d653} /* (2, 0, 23) {real, imag} */,
  {32'hc2180096, 32'hc2b3be15} /* (2, 0, 22) {real, imag} */,
  {32'hc1ac7e70, 32'hc2bac327} /* (2, 0, 21) {real, imag} */,
  {32'h42c660fc, 32'h42f57d49} /* (2, 0, 20) {real, imag} */,
  {32'h424340a5, 32'hc1c16e8c} /* (2, 0, 19) {real, imag} */,
  {32'hc1bf586c, 32'hc092fd90} /* (2, 0, 18) {real, imag} */,
  {32'h41ffb550, 32'h4239dfd8} /* (2, 0, 17) {real, imag} */,
  {32'hc1989560, 32'hc1cb7780} /* (2, 0, 16) {real, imag} */,
  {32'h418f8c50, 32'h40e49340} /* (2, 0, 15) {real, imag} */,
  {32'hc1a7126c, 32'h417d1f48} /* (2, 0, 14) {real, imag} */,
  {32'hc2782e0f, 32'hc26edb9a} /* (2, 0, 13) {real, imag} */,
  {32'h426a2688, 32'hc2084516} /* (2, 0, 12) {real, imag} */,
  {32'h42b0cc68, 32'h40de7b70} /* (2, 0, 11) {real, imag} */,
  {32'h428c045b, 32'h427bd012} /* (2, 0, 10) {real, imag} */,
  {32'h423864c0, 32'hc2eac555} /* (2, 0, 9) {real, imag} */,
  {32'h43acbdad, 32'h4276a2ae} /* (2, 0, 8) {real, imag} */,
  {32'hc3cae62c, 32'hc29552c5} /* (2, 0, 7) {real, imag} */,
  {32'hc2cfe556, 32'hc27a6036} /* (2, 0, 6) {real, imag} */,
  {32'h42c38d3c, 32'hc3f507e0} /* (2, 0, 5) {real, imag} */,
  {32'h433dad19, 32'hc1b42216} /* (2, 0, 4) {real, imag} */,
  {32'h430c00ce, 32'hc341eae5} /* (2, 0, 3) {real, imag} */,
  {32'h444404b0, 32'hc38b545d} /* (2, 0, 2) {real, imag} */,
  {32'hc4cff07a, 32'h44b2125a} /* (2, 0, 1) {real, imag} */,
  {32'hc3b53fda, 32'h44cad3ee} /* (2, 0, 0) {real, imag} */,
  {32'hc45e807f, 32'hc5051eba} /* (1, 31, 31) {real, imag} */,
  {32'h44437dd2, 32'h448d7892} /* (1, 31, 30) {real, imag} */,
  {32'h432748c3, 32'h42aabca4} /* (1, 31, 29) {real, imag} */,
  {32'h42452ff0, 32'hc295e8bc} /* (1, 31, 28) {real, imag} */,
  {32'h42cb8555, 32'h43d10912} /* (1, 31, 27) {real, imag} */,
  {32'h4273d8a0, 32'h42916576} /* (1, 31, 26) {real, imag} */,
  {32'hc33da750, 32'hc35765a7} /* (1, 31, 25) {real, imag} */,
  {32'h4383edb8, 32'h433e16fb} /* (1, 31, 24) {real, imag} */,
  {32'hc2db9d9d, 32'h425e3d44} /* (1, 31, 23) {real, imag} */,
  {32'h41f0fa80, 32'h3f5b2a00} /* (1, 31, 22) {real, imag} */,
  {32'h432ba468, 32'h42c51618} /* (1, 31, 21) {real, imag} */,
  {32'h42bd88cd, 32'hc2393048} /* (1, 31, 20) {real, imag} */,
  {32'h41ad7a16, 32'hc1680adc} /* (1, 31, 19) {real, imag} */,
  {32'h42620168, 32'h42455168} /* (1, 31, 18) {real, imag} */,
  {32'hc1c66fc0, 32'hc1b2c118} /* (1, 31, 17) {real, imag} */,
  {32'hc2282a3b, 32'hc1106080} /* (1, 31, 16) {real, imag} */,
  {32'hc093d580, 32'h41165ab0} /* (1, 31, 15) {real, imag} */,
  {32'hc2fbf214, 32'h428b41ac} /* (1, 31, 14) {real, imag} */,
  {32'hc1dfe9fe, 32'h423eafaf} /* (1, 31, 13) {real, imag} */,
  {32'h4291d4af, 32'hc264fe8c} /* (1, 31, 12) {real, imag} */,
  {32'hc2b83ee4, 32'h431b97a4} /* (1, 31, 11) {real, imag} */,
  {32'hc3320274, 32'h403c0a80} /* (1, 31, 10) {real, imag} */,
  {32'hc1c4b314, 32'h42b93c22} /* (1, 31, 9) {real, imag} */,
  {32'h40341800, 32'h42f7fdda} /* (1, 31, 8) {real, imag} */,
  {32'h4185dfa4, 32'h42c8961a} /* (1, 31, 7) {real, imag} */,
  {32'hc35f0ca4, 32'hc23f58fc} /* (1, 31, 6) {real, imag} */,
  {32'hc2876293, 32'h4400fa9b} /* (1, 31, 5) {real, imag} */,
  {32'hc382ae50, 32'hc3e83337} /* (1, 31, 4) {real, imag} */,
  {32'h422ca10b, 32'h42856d84} /* (1, 31, 3) {real, imag} */,
  {32'hc2443648, 32'h4410fd6c} /* (1, 31, 2) {real, imag} */,
  {32'h4400b8d5, 32'hc4b1e7e4} /* (1, 31, 1) {real, imag} */,
  {32'hc232040d, 32'hc4c01c98} /* (1, 31, 0) {real, imag} */,
  {32'hc3b431c0, 32'h44702c3c} /* (1, 30, 31) {real, imag} */,
  {32'h4387c93c, 32'hc45c1cbe} /* (1, 30, 30) {real, imag} */,
  {32'hc36e81e8, 32'h42808aa8} /* (1, 30, 29) {real, imag} */,
  {32'h428d391a, 32'h438655b2} /* (1, 30, 28) {real, imag} */,
  {32'hc359c9a3, 32'hc3c7f1c0} /* (1, 30, 27) {real, imag} */,
  {32'hc249f078, 32'h427a8add} /* (1, 30, 26) {real, imag} */,
  {32'h42f8d7ac, 32'h42ad9a66} /* (1, 30, 25) {real, imag} */,
  {32'hc328047d, 32'hc37c12e7} /* (1, 30, 24) {real, imag} */,
  {32'hc19a9206, 32'h4186b240} /* (1, 30, 23) {real, imag} */,
  {32'h41d3e0f2, 32'h424e64f7} /* (1, 30, 22) {real, imag} */,
  {32'hc2f1186c, 32'hc284745c} /* (1, 30, 21) {real, imag} */,
  {32'h408d67e8, 32'hc1bfac0c} /* (1, 30, 20) {real, imag} */,
  {32'hc0e7e6e0, 32'h426a6ec9} /* (1, 30, 19) {real, imag} */,
  {32'hc0a274d8, 32'h412c7268} /* (1, 30, 18) {real, imag} */,
  {32'h41872d36, 32'h41d0c4f0} /* (1, 30, 17) {real, imag} */,
  {32'h41b892d8, 32'hc1ca4ef0} /* (1, 30, 16) {real, imag} */,
  {32'h40aa0c68, 32'hc1e5e2b0} /* (1, 30, 15) {real, imag} */,
  {32'h4255873b, 32'h4188cc8c} /* (1, 30, 14) {real, imag} */,
  {32'h426850f8, 32'h41f70c96} /* (1, 30, 13) {real, imag} */,
  {32'h412c6a84, 32'hc268c50e} /* (1, 30, 12) {real, imag} */,
  {32'h41657cd4, 32'h4207e688} /* (1, 30, 11) {real, imag} */,
  {32'hc0a8fc08, 32'h41d53f6e} /* (1, 30, 10) {real, imag} */,
  {32'h413723f4, 32'h4303d722} /* (1, 30, 9) {real, imag} */,
  {32'h4338413d, 32'hc35cd90d} /* (1, 30, 8) {real, imag} */,
  {32'h42079018, 32'hc1fca166} /* (1, 30, 7) {real, imag} */,
  {32'h42a30198, 32'hc2ba99ae} /* (1, 30, 6) {real, imag} */,
  {32'h43421415, 32'hc3a61052} /* (1, 30, 5) {real, imag} */,
  {32'hc38f5bca, 32'h4214d0ac} /* (1, 30, 4) {real, imag} */,
  {32'hc36e31a8, 32'h42af3322} /* (1, 30, 3) {real, imag} */,
  {32'h44094b88, 32'hc493f951} /* (1, 30, 2) {real, imag} */,
  {32'hc30413af, 32'h44efbcfe} /* (1, 30, 1) {real, imag} */,
  {32'h420c97bf, 32'h4470c0fc} /* (1, 30, 0) {real, imag} */,
  {32'hc389bc6c, 32'hc405a2e2} /* (1, 29, 31) {real, imag} */,
  {32'h434c77df, 32'hc06b6af0} /* (1, 29, 30) {real, imag} */,
  {32'hc2960c13, 32'h432bfd65} /* (1, 29, 29) {real, imag} */,
  {32'hc28bc006, 32'h432874b8} /* (1, 29, 28) {real, imag} */,
  {32'hc3018fcd, 32'hc21f6c28} /* (1, 29, 27) {real, imag} */,
  {32'hc29afc8a, 32'h4144b580} /* (1, 29, 26) {real, imag} */,
  {32'h42ab5c71, 32'h42897640} /* (1, 29, 25) {real, imag} */,
  {32'hc26f8b98, 32'hc2184463} /* (1, 29, 24) {real, imag} */,
  {32'h42abe8a6, 32'hc2d2517a} /* (1, 29, 23) {real, imag} */,
  {32'hc1cc66b6, 32'h427662ec} /* (1, 29, 22) {real, imag} */,
  {32'hc196b940, 32'h423dc13a} /* (1, 29, 21) {real, imag} */,
  {32'h41c53394, 32'hc0cff450} /* (1, 29, 20) {real, imag} */,
  {32'hc105f5fe, 32'h4128dc70} /* (1, 29, 19) {real, imag} */,
  {32'h423fc7ec, 32'hc3007baa} /* (1, 29, 18) {real, imag} */,
  {32'hc0f1af42, 32'h41c178c0} /* (1, 29, 17) {real, imag} */,
  {32'hc177bcea, 32'h42781438} /* (1, 29, 16) {real, imag} */,
  {32'hc029237c, 32'h40d10fc0} /* (1, 29, 15) {real, imag} */,
  {32'h41a0d6e8, 32'h424e14a2} /* (1, 29, 14) {real, imag} */,
  {32'hc17adffe, 32'hc25015dc} /* (1, 29, 13) {real, imag} */,
  {32'hc2565714, 32'hc03581a0} /* (1, 29, 12) {real, imag} */,
  {32'hc2019c1d, 32'hc0e47f00} /* (1, 29, 11) {real, imag} */,
  {32'h429fe398, 32'hc29ba928} /* (1, 29, 10) {real, imag} */,
  {32'h42370d09, 32'h41ce1170} /* (1, 29, 9) {real, imag} */,
  {32'h41d9430b, 32'hc2e78a1e} /* (1, 29, 8) {real, imag} */,
  {32'hc23a3d3e, 32'h41fe7e48} /* (1, 29, 7) {real, imag} */,
  {32'hc17dc2fc, 32'h42609c94} /* (1, 29, 6) {real, imag} */,
  {32'hc1a1f8c0, 32'h435f28d8} /* (1, 29, 5) {real, imag} */,
  {32'hc307109f, 32'hc3752fe8} /* (1, 29, 4) {real, imag} */,
  {32'h429b1453, 32'h420e843c} /* (1, 29, 3) {real, imag} */,
  {32'h43ee3068, 32'hc0599970} /* (1, 29, 2) {real, imag} */,
  {32'hc3705718, 32'h437e304e} /* (1, 29, 1) {real, imag} */,
  {32'h4210eb4c, 32'h42cb9d44} /* (1, 29, 0) {real, imag} */,
  {32'hc38635c2, 32'hc426166c} /* (1, 28, 31) {real, imag} */,
  {32'h43508add, 32'h43d3efe8} /* (1, 28, 30) {real, imag} */,
  {32'hc301b1c4, 32'hbf38d000} /* (1, 28, 29) {real, imag} */,
  {32'hc37eb99f, 32'h42ef367e} /* (1, 28, 28) {real, imag} */,
  {32'h4376bdd8, 32'h429fc6ec} /* (1, 28, 27) {real, imag} */,
  {32'h42d70632, 32'hc2a180fa} /* (1, 28, 26) {real, imag} */,
  {32'h428dcc60, 32'hc2c59324} /* (1, 28, 25) {real, imag} */,
  {32'h429b8570, 32'hc0fcd1a0} /* (1, 28, 24) {real, imag} */,
  {32'hbf980070, 32'hc1c3d660} /* (1, 28, 23) {real, imag} */,
  {32'hc1ac448a, 32'h416daace} /* (1, 28, 22) {real, imag} */,
  {32'h42ff44fe, 32'hc2acdc58} /* (1, 28, 21) {real, imag} */,
  {32'hc29ad8fa, 32'h4221abac} /* (1, 28, 20) {real, imag} */,
  {32'h420df3d3, 32'h41a9c358} /* (1, 28, 19) {real, imag} */,
  {32'h42479c3a, 32'hc28e29fc} /* (1, 28, 18) {real, imag} */,
  {32'hc23f732d, 32'h404cc5a0} /* (1, 28, 17) {real, imag} */,
  {32'hbf94b4c0, 32'hc101a990} /* (1, 28, 16) {real, imag} */,
  {32'h41abef1a, 32'h4031e3e0} /* (1, 28, 15) {real, imag} */,
  {32'h418d1c6c, 32'h41effc70} /* (1, 28, 14) {real, imag} */,
  {32'hc0b3b008, 32'hbfdbf580} /* (1, 28, 13) {real, imag} */,
  {32'hc1c87f26, 32'hc0becc7c} /* (1, 28, 12) {real, imag} */,
  {32'h42948f26, 32'hc21c2af0} /* (1, 28, 11) {real, imag} */,
  {32'h42b23f76, 32'h4189654f} /* (1, 28, 10) {real, imag} */,
  {32'hc2244a6c, 32'hc2b0b00f} /* (1, 28, 9) {real, imag} */,
  {32'hc1376340, 32'h42ac4057} /* (1, 28, 8) {real, imag} */,
  {32'hc1a58870, 32'h4278cb67} /* (1, 28, 7) {real, imag} */,
  {32'h410a0094, 32'h42d7b0b4} /* (1, 28, 6) {real, imag} */,
  {32'hc290a30c, 32'h42806744} /* (1, 28, 5) {real, imag} */,
  {32'hc1b93db8, 32'hc334def1} /* (1, 28, 4) {real, imag} */,
  {32'hc1889cd4, 32'hc2dcf5dc} /* (1, 28, 3) {real, imag} */,
  {32'h438a39aa, 32'h438c2e9e} /* (1, 28, 2) {real, imag} */,
  {32'hc3d15336, 32'hc37d8492} /* (1, 28, 1) {real, imag} */,
  {32'h4329cbe2, 32'hc39ae198} /* (1, 28, 0) {real, imag} */,
  {32'h43c530a8, 32'h43806910} /* (1, 27, 31) {real, imag} */,
  {32'hc36da8df, 32'hc34d9682} /* (1, 27, 30) {real, imag} */,
  {32'hc2c8c026, 32'h42c37758} /* (1, 27, 29) {real, imag} */,
  {32'h42b183da, 32'h416ac69c} /* (1, 27, 28) {real, imag} */,
  {32'hc286b98b, 32'hc231356a} /* (1, 27, 27) {real, imag} */,
  {32'hc227042c, 32'h3d302800} /* (1, 27, 26) {real, imag} */,
  {32'h41ddec30, 32'h4326c512} /* (1, 27, 25) {real, imag} */,
  {32'hc27355cb, 32'h4237f4f7} /* (1, 27, 24) {real, imag} */,
  {32'hc23eb896, 32'hc2af7f2b} /* (1, 27, 23) {real, imag} */,
  {32'hc286184e, 32'h415de598} /* (1, 27, 22) {real, imag} */,
  {32'hc2cd146f, 32'hc1e60dad} /* (1, 27, 21) {real, imag} */,
  {32'hc22aee67, 32'hc28d0122} /* (1, 27, 20) {real, imag} */,
  {32'h411844c5, 32'hc2157db8} /* (1, 27, 19) {real, imag} */,
  {32'hc1edcbec, 32'h41eacc3d} /* (1, 27, 18) {real, imag} */,
  {32'h3f773ac0, 32'hc0d45a40} /* (1, 27, 17) {real, imag} */,
  {32'hbd77e000, 32'hc157c280} /* (1, 27, 16) {real, imag} */,
  {32'hc2264529, 32'h3de0b000} /* (1, 27, 15) {real, imag} */,
  {32'h414f8038, 32'h41c396f3} /* (1, 27, 14) {real, imag} */,
  {32'h411899db, 32'h41335440} /* (1, 27, 13) {real, imag} */,
  {32'h4224acd9, 32'h429caf10} /* (1, 27, 12) {real, imag} */,
  {32'hc1338068, 32'hc2425166} /* (1, 27, 11) {real, imag} */,
  {32'h415122d4, 32'hc105a8a0} /* (1, 27, 10) {real, imag} */,
  {32'hc1aed074, 32'h421908a2} /* (1, 27, 9) {real, imag} */,
  {32'h42e38956, 32'hc2e62af0} /* (1, 27, 8) {real, imag} */,
  {32'hc280c89a, 32'hc1f0b104} /* (1, 27, 7) {real, imag} */,
  {32'hc119c9b6, 32'h42a7f44a} /* (1, 27, 6) {real, imag} */,
  {32'hc21ce07a, 32'hc286928d} /* (1, 27, 5) {real, imag} */,
  {32'h420e68d3, 32'h42bc327c} /* (1, 27, 4) {real, imag} */,
  {32'hc2c9ab72, 32'h43533d66} /* (1, 27, 3) {real, imag} */,
  {32'h42220ec4, 32'hc310471c} /* (1, 27, 2) {real, imag} */,
  {32'hc2edad1a, 32'h4417e4f2} /* (1, 27, 1) {real, imag} */,
  {32'h438ec484, 32'h439e1a86} /* (1, 27, 0) {real, imag} */,
  {32'hc2b87dbb, 32'hc1aa8d80} /* (1, 26, 31) {real, imag} */,
  {32'hc28683fe, 32'h4350a5a6} /* (1, 26, 30) {real, imag} */,
  {32'hc315cf1e, 32'h42f6145d} /* (1, 26, 29) {real, imag} */,
  {32'h4298287b, 32'h42c5b1f5} /* (1, 26, 28) {real, imag} */,
  {32'h42a02943, 32'hc2c079d0} /* (1, 26, 27) {real, imag} */,
  {32'hc3273dcc, 32'hc290a679} /* (1, 26, 26) {real, imag} */,
  {32'h417beff4, 32'hc2d6dac6} /* (1, 26, 25) {real, imag} */,
  {32'h427f8872, 32'hc24fa0d0} /* (1, 26, 24) {real, imag} */,
  {32'h420a3330, 32'h4254ef42} /* (1, 26, 23) {real, imag} */,
  {32'h42d28e27, 32'hc215409d} /* (1, 26, 22) {real, imag} */,
  {32'h41827b46, 32'hc22ef4f5} /* (1, 26, 21) {real, imag} */,
  {32'hc2611ded, 32'h40ca9ace} /* (1, 26, 20) {real, imag} */,
  {32'hc1cbbdc2, 32'hc19a98fa} /* (1, 26, 19) {real, imag} */,
  {32'hc197cf66, 32'hc202393a} /* (1, 26, 18) {real, imag} */,
  {32'hc090536c, 32'h40a2d018} /* (1, 26, 17) {real, imag} */,
  {32'h41f8f9e1, 32'h42709563} /* (1, 26, 16) {real, imag} */,
  {32'hc103930a, 32'h41a094da} /* (1, 26, 15) {real, imag} */,
  {32'h419987ae, 32'hc206dec2} /* (1, 26, 14) {real, imag} */,
  {32'hc2a28fbc, 32'h41b3100a} /* (1, 26, 13) {real, imag} */,
  {32'hc0c84a90, 32'h41b45f6c} /* (1, 26, 12) {real, imag} */,
  {32'hc19959f2, 32'h4162bbc4} /* (1, 26, 11) {real, imag} */,
  {32'hc1873e14, 32'hc21008d1} /* (1, 26, 10) {real, imag} */,
  {32'hc2444cd8, 32'h41d1a445} /* (1, 26, 9) {real, imag} */,
  {32'h420b55e6, 32'hc2539e9a} /* (1, 26, 8) {real, imag} */,
  {32'h42b68656, 32'hc2b64d0c} /* (1, 26, 7) {real, imag} */,
  {32'h3f189d80, 32'hc2bd28cb} /* (1, 26, 6) {real, imag} */,
  {32'hc1b7dbc4, 32'hc28fe52c} /* (1, 26, 5) {real, imag} */,
  {32'h41b1a7cd, 32'h4298fcf5} /* (1, 26, 4) {real, imag} */,
  {32'h42f6a4f0, 32'hc27c3286} /* (1, 26, 3) {real, imag} */,
  {32'h417db064, 32'hc30b50dc} /* (1, 26, 2) {real, imag} */,
  {32'hc26c9f9a, 32'hc33a6544} /* (1, 26, 1) {real, imag} */,
  {32'h42356e10, 32'h42520e2b} /* (1, 26, 0) {real, imag} */,
  {32'hc2d1b5e7, 32'h430dfefb} /* (1, 25, 31) {real, imag} */,
  {32'h42ec2e76, 32'h423cb59c} /* (1, 25, 30) {real, imag} */,
  {32'h420a4be4, 32'h42d96061} /* (1, 25, 29) {real, imag} */,
  {32'hc30a1869, 32'h43216f03} /* (1, 25, 28) {real, imag} */,
  {32'h424e39a6, 32'hc2f25e30} /* (1, 25, 27) {real, imag} */,
  {32'h4220ac2e, 32'hc2b65131} /* (1, 25, 26) {real, imag} */,
  {32'hc15e9dc8, 32'hc1f10092} /* (1, 25, 25) {real, imag} */,
  {32'h4211c8a7, 32'hc207c3cb} /* (1, 25, 24) {real, imag} */,
  {32'h41c918d9, 32'hc2193770} /* (1, 25, 23) {real, imag} */,
  {32'h40cd6864, 32'hc2ca2050} /* (1, 25, 22) {real, imag} */,
  {32'hc1bdbded, 32'hc2805545} /* (1, 25, 21) {real, imag} */,
  {32'h41fbb48b, 32'h425c8d32} /* (1, 25, 20) {real, imag} */,
  {32'hc186ad71, 32'hc099cf4e} /* (1, 25, 19) {real, imag} */,
  {32'h41a3d794, 32'h4216facc} /* (1, 25, 18) {real, imag} */,
  {32'h420372ce, 32'h41c615df} /* (1, 25, 17) {real, imag} */,
  {32'hc1d26e54, 32'h4219d9da} /* (1, 25, 16) {real, imag} */,
  {32'hc1dd60c5, 32'hc1779052} /* (1, 25, 15) {real, imag} */,
  {32'h40ea08f0, 32'hc1c3fe17} /* (1, 25, 14) {real, imag} */,
  {32'hc205f04a, 32'hc18b5588} /* (1, 25, 13) {real, imag} */,
  {32'h40791388, 32'hc18e11b0} /* (1, 25, 12) {real, imag} */,
  {32'hc244f6ba, 32'hc2199404} /* (1, 25, 11) {real, imag} */,
  {32'hc283a886, 32'hc01db4d0} /* (1, 25, 10) {real, imag} */,
  {32'h4202508c, 32'h4301773e} /* (1, 25, 9) {real, imag} */,
  {32'h42884408, 32'h4249310f} /* (1, 25, 8) {real, imag} */,
  {32'h4279ad66, 32'hc2c38d46} /* (1, 25, 7) {real, imag} */,
  {32'h42a26a91, 32'hc2365b0e} /* (1, 25, 6) {real, imag} */,
  {32'h41192e74, 32'hc1b50ef0} /* (1, 25, 5) {real, imag} */,
  {32'hc2a39e7e, 32'h42cde196} /* (1, 25, 4) {real, imag} */,
  {32'hc271b020, 32'h42ab7657} /* (1, 25, 3) {real, imag} */,
  {32'hc258d57d, 32'hc2af4ae6} /* (1, 25, 2) {real, imag} */,
  {32'hc305a924, 32'hc37a1d6d} /* (1, 25, 1) {real, imag} */,
  {32'h404b4720, 32'h4191c2c4} /* (1, 25, 0) {real, imag} */,
  {32'h42f439ae, 32'h438bafb7} /* (1, 24, 31) {real, imag} */,
  {32'hc13cf956, 32'hc3a35b55} /* (1, 24, 30) {real, imag} */,
  {32'h41006e6c, 32'hc1c3b9d8} /* (1, 24, 29) {real, imag} */,
  {32'h42dd95d9, 32'h4288f362} /* (1, 24, 28) {real, imag} */,
  {32'hc004270c, 32'hc29e8b02} /* (1, 24, 27) {real, imag} */,
  {32'hc2ad6cd3, 32'h4171be52} /* (1, 24, 26) {real, imag} */,
  {32'hc279b0c0, 32'h42d77ba9} /* (1, 24, 25) {real, imag} */,
  {32'hc270fbc2, 32'hc28973c2} /* (1, 24, 24) {real, imag} */,
  {32'hc27298d2, 32'h407e6f78} /* (1, 24, 23) {real, imag} */,
  {32'h4245b411, 32'hc11ff71a} /* (1, 24, 22) {real, imag} */,
  {32'hc21999f8, 32'h41dec7e0} /* (1, 24, 21) {real, imag} */,
  {32'hc1f49af8, 32'hc1a96622} /* (1, 24, 20) {real, imag} */,
  {32'h4200cf0b, 32'h41d7af76} /* (1, 24, 19) {real, imag} */,
  {32'hc1810001, 32'hc0f935f0} /* (1, 24, 18) {real, imag} */,
  {32'h4184ae63, 32'hc0c854f0} /* (1, 24, 17) {real, imag} */,
  {32'hc222c1c8, 32'h4168e528} /* (1, 24, 16) {real, imag} */,
  {32'h4204c90e, 32'hc15f0748} /* (1, 24, 15) {real, imag} */,
  {32'h4061ead8, 32'hc1bea27c} /* (1, 24, 14) {real, imag} */,
  {32'h3fd6ffe8, 32'hc133180f} /* (1, 24, 13) {real, imag} */,
  {32'hc0c4af90, 32'h421946a0} /* (1, 24, 12) {real, imag} */,
  {32'hc149df06, 32'h4157c460} /* (1, 24, 11) {real, imag} */,
  {32'hc2018337, 32'h428348c5} /* (1, 24, 10) {real, imag} */,
  {32'h426daa82, 32'h41f8d261} /* (1, 24, 9) {real, imag} */,
  {32'h4188680b, 32'hc2c7f908} /* (1, 24, 8) {real, imag} */,
  {32'hc25f742c, 32'h3f60d780} /* (1, 24, 7) {real, imag} */,
  {32'hbf013980, 32'hc24930a8} /* (1, 24, 6) {real, imag} */,
  {32'h414e5ebd, 32'hc3867352} /* (1, 24, 5) {real, imag} */,
  {32'hc2cbd00f, 32'hc1258e8c} /* (1, 24, 4) {real, imag} */,
  {32'hc234e7b9, 32'h415a2b83} /* (1, 24, 3) {real, imag} */,
  {32'hc1b675db, 32'hc3267cfa} /* (1, 24, 2) {real, imag} */,
  {32'h4351bf0d, 32'h43d6be97} /* (1, 24, 1) {real, imag} */,
  {32'h42581380, 32'h42bd6e45} /* (1, 24, 0) {real, imag} */,
  {32'hc31104d1, 32'hc245e2fc} /* (1, 23, 31) {real, imag} */,
  {32'h42e8eb63, 32'h42dbc34a} /* (1, 23, 30) {real, imag} */,
  {32'hc33ee058, 32'hc302d1be} /* (1, 23, 29) {real, imag} */,
  {32'h42a7f8fb, 32'h4285a7ed} /* (1, 23, 28) {real, imag} */,
  {32'h42f9e722, 32'h42271212} /* (1, 23, 27) {real, imag} */,
  {32'hc1abecb7, 32'hc1ea45b0} /* (1, 23, 26) {real, imag} */,
  {32'hc1cf393d, 32'h426a14a7} /* (1, 23, 25) {real, imag} */,
  {32'h4288e82e, 32'h42a20eb7} /* (1, 23, 24) {real, imag} */,
  {32'hc2c8a6cc, 32'h422c60b6} /* (1, 23, 23) {real, imag} */,
  {32'h423eea94, 32'h3fc36a40} /* (1, 23, 22) {real, imag} */,
  {32'h417947c2, 32'h414bcae7} /* (1, 23, 21) {real, imag} */,
  {32'h4207d7f9, 32'hbee0f600} /* (1, 23, 20) {real, imag} */,
  {32'h418fd55f, 32'h3fa24870} /* (1, 23, 19) {real, imag} */,
  {32'hc19cac8b, 32'hc12eac5a} /* (1, 23, 18) {real, imag} */,
  {32'hc20f37a3, 32'h41b172c7} /* (1, 23, 17) {real, imag} */,
  {32'h419e53ee, 32'hbe0e5880} /* (1, 23, 16) {real, imag} */,
  {32'hc1b63bba, 32'h420382c4} /* (1, 23, 15) {real, imag} */,
  {32'h41cf82f3, 32'hc1ad1621} /* (1, 23, 14) {real, imag} */,
  {32'hc2266924, 32'hc0240468} /* (1, 23, 13) {real, imag} */,
  {32'hc211c1f1, 32'h41889200} /* (1, 23, 12) {real, imag} */,
  {32'h4224f42e, 32'h41724685} /* (1, 23, 11) {real, imag} */,
  {32'h418f8000, 32'hc1c2f098} /* (1, 23, 10) {real, imag} */,
  {32'h410c5f44, 32'h428447de} /* (1, 23, 9) {real, imag} */,
  {32'hc19b4f68, 32'h42bf81fd} /* (1, 23, 8) {real, imag} */,
  {32'hc03452c8, 32'h41f7c38e} /* (1, 23, 7) {real, imag} */,
  {32'h42a9e53c, 32'hc2bd0633} /* (1, 23, 6) {real, imag} */,
  {32'h3e070100, 32'h40aef894} /* (1, 23, 5) {real, imag} */,
  {32'h4268751a, 32'hc29abc69} /* (1, 23, 4) {real, imag} */,
  {32'hc3192ebc, 32'h41672720} /* (1, 23, 3) {real, imag} */,
  {32'h4376e0f2, 32'hc2478e0c} /* (1, 23, 2) {real, imag} */,
  {32'hc2a0c426, 32'h42ab26da} /* (1, 23, 1) {real, imag} */,
  {32'hc29f7c78, 32'h41756dc2} /* (1, 23, 0) {real, imag} */,
  {32'hc29a212a, 32'hc2a3bd0a} /* (1, 22, 31) {real, imag} */,
  {32'h4122f028, 32'hc2accc35} /* (1, 22, 30) {real, imag} */,
  {32'h41d9ee4a, 32'hc1c6b9b6} /* (1, 22, 29) {real, imag} */,
  {32'hc221dd6a, 32'hc27e94ef} /* (1, 22, 28) {real, imag} */,
  {32'h422dc173, 32'hc2ab2c3d} /* (1, 22, 27) {real, imag} */,
  {32'hbffe5970, 32'h41b84388} /* (1, 22, 26) {real, imag} */,
  {32'h41d50370, 32'h410024f4} /* (1, 22, 25) {real, imag} */,
  {32'h4134666e, 32'h425eddc1} /* (1, 22, 24) {real, imag} */,
  {32'h410c06f5, 32'hc28c37f0} /* (1, 22, 23) {real, imag} */,
  {32'h4127d2b2, 32'h41c5cf92} /* (1, 22, 22) {real, imag} */,
  {32'hc0ec2190, 32'hc0d0ae84} /* (1, 22, 21) {real, imag} */,
  {32'h417f8d1d, 32'hc0586bbc} /* (1, 22, 20) {real, imag} */,
  {32'h41856903, 32'h40b9be58} /* (1, 22, 19) {real, imag} */,
  {32'h41838c15, 32'h4042c7a0} /* (1, 22, 18) {real, imag} */,
  {32'h410c61c0, 32'hc05c9af0} /* (1, 22, 17) {real, imag} */,
  {32'h411d6070, 32'h40a12488} /* (1, 22, 16) {real, imag} */,
  {32'h403f4d22, 32'hc1144c4c} /* (1, 22, 15) {real, imag} */,
  {32'h4181a6dd, 32'h41aa68f6} /* (1, 22, 14) {real, imag} */,
  {32'h40d55749, 32'h418b1b98} /* (1, 22, 13) {real, imag} */,
  {32'hc0d3590e, 32'hc1fdd004} /* (1, 22, 12) {real, imag} */,
  {32'hc1f4f380, 32'h41346e72} /* (1, 22, 11) {real, imag} */,
  {32'hc1d02841, 32'hc1135367} /* (1, 22, 10) {real, imag} */,
  {32'h414dfbf5, 32'h41233f5c} /* (1, 22, 9) {real, imag} */,
  {32'hc24bba98, 32'h41bfc872} /* (1, 22, 8) {real, imag} */,
  {32'hc1d23304, 32'h4281202c} /* (1, 22, 7) {real, imag} */,
  {32'h40672078, 32'h3f8f9f18} /* (1, 22, 6) {real, imag} */,
  {32'hc08d4008, 32'h407c8ba0} /* (1, 22, 5) {real, imag} */,
  {32'hc09d5d6c, 32'hc1fb0986} /* (1, 22, 4) {real, imag} */,
  {32'hc0a9ac52, 32'hc2202885} /* (1, 22, 3) {real, imag} */,
  {32'h42f41fe5, 32'h42134612} /* (1, 22, 2) {real, imag} */,
  {32'hc2c259d2, 32'hc0a70a08} /* (1, 22, 1) {real, imag} */,
  {32'hc2b2e1b0, 32'h42a043ea} /* (1, 22, 0) {real, imag} */,
  {32'h4323de24, 32'h422fce6f} /* (1, 21, 31) {real, imag} */,
  {32'hc2e8f8aa, 32'hc1964e22} /* (1, 21, 30) {real, imag} */,
  {32'h4166200e, 32'hc21f1c78} /* (1, 21, 29) {real, imag} */,
  {32'h42abc068, 32'hc1265388} /* (1, 21, 28) {real, imag} */,
  {32'hc1c9ba3e, 32'hc176e724} /* (1, 21, 27) {real, imag} */,
  {32'hc0eaab3e, 32'hc285965c} /* (1, 21, 26) {real, imag} */,
  {32'h4180aecd, 32'h421b8f00} /* (1, 21, 25) {real, imag} */,
  {32'hc0e89990, 32'h40c06070} /* (1, 21, 24) {real, imag} */,
  {32'h42325744, 32'hc1655f67} /* (1, 21, 23) {real, imag} */,
  {32'hc1f7cdf0, 32'h40ebc124} /* (1, 21, 22) {real, imag} */,
  {32'h41355a2d, 32'hbf71b090} /* (1, 21, 21) {real, imag} */,
  {32'h4232e298, 32'h41d49cbb} /* (1, 21, 20) {real, imag} */,
  {32'hc14989d2, 32'hc086ba02} /* (1, 21, 19) {real, imag} */,
  {32'h412277d8, 32'h3ec13430} /* (1, 21, 18) {real, imag} */,
  {32'hbf850998, 32'hbfcc8a58} /* (1, 21, 17) {real, imag} */,
  {32'h4118115c, 32'hc19a32ae} /* (1, 21, 16) {real, imag} */,
  {32'h411e5df3, 32'h41208dff} /* (1, 21, 15) {real, imag} */,
  {32'hc1e80dcc, 32'h4008884a} /* (1, 21, 14) {real, imag} */,
  {32'h3fc70094, 32'h40af245a} /* (1, 21, 13) {real, imag} */,
  {32'hc04d8f18, 32'hc1a038e3} /* (1, 21, 12) {real, imag} */,
  {32'hc0948dba, 32'h3ebf8320} /* (1, 21, 11) {real, imag} */,
  {32'hc126bfcf, 32'hc1c5841d} /* (1, 21, 10) {real, imag} */,
  {32'hc1948c71, 32'hc1bacfde} /* (1, 21, 9) {real, imag} */,
  {32'h41a3f5e6, 32'hc28d63d2} /* (1, 21, 8) {real, imag} */,
  {32'h4198998b, 32'hbf557520} /* (1, 21, 7) {real, imag} */,
  {32'hc13fcf11, 32'hc2e98ab8} /* (1, 21, 6) {real, imag} */,
  {32'hc29d399c, 32'hc299e792} /* (1, 21, 5) {real, imag} */,
  {32'hc03fa890, 32'h409299ea} /* (1, 21, 4) {real, imag} */,
  {32'hc236db60, 32'h41a0b2bf} /* (1, 21, 3) {real, imag} */,
  {32'hc2997f3a, 32'hc24b5417} /* (1, 21, 2) {real, imag} */,
  {32'h430d4d46, 32'h42abe816} /* (1, 21, 1) {real, imag} */,
  {32'h42c9d5c6, 32'h42b62806} /* (1, 21, 0) {real, imag} */,
  {32'h42324109, 32'hc198b334} /* (1, 20, 31) {real, imag} */,
  {32'hc24085c8, 32'hc115f4fd} /* (1, 20, 30) {real, imag} */,
  {32'h42734650, 32'h40dca54b} /* (1, 20, 29) {real, imag} */,
  {32'hc141be9f, 32'hc25c059c} /* (1, 20, 28) {real, imag} */,
  {32'h423fe2fa, 32'h3ffc48a0} /* (1, 20, 27) {real, imag} */,
  {32'h410e817c, 32'hc1ab12e2} /* (1, 20, 26) {real, imag} */,
  {32'hc1605df8, 32'hc1a0daf6} /* (1, 20, 25) {real, imag} */,
  {32'hc1a4ec99, 32'hc2053b22} /* (1, 20, 24) {real, imag} */,
  {32'hbf697240, 32'h41b534f7} /* (1, 20, 23) {real, imag} */,
  {32'hc1a36bb4, 32'h421a8b10} /* (1, 20, 22) {real, imag} */,
  {32'h3f35b5f0, 32'h418ca44e} /* (1, 20, 21) {real, imag} */,
  {32'hc0ee6734, 32'hc194cecc} /* (1, 20, 20) {real, imag} */,
  {32'h40c10178, 32'h40defbdf} /* (1, 20, 19) {real, imag} */,
  {32'hc1113626, 32'h40fb7c56} /* (1, 20, 18) {real, imag} */,
  {32'h40390b00, 32'hc045e794} /* (1, 20, 17) {real, imag} */,
  {32'hbfb5f100, 32'hc196331a} /* (1, 20, 16) {real, imag} */,
  {32'h41051c90, 32'hc167fe7f} /* (1, 20, 15) {real, imag} */,
  {32'hc1bd529d, 32'hc103340f} /* (1, 20, 14) {real, imag} */,
  {32'hc131b6d4, 32'h4124ab6e} /* (1, 20, 13) {real, imag} */,
  {32'h41a316fe, 32'hc1df073c} /* (1, 20, 12) {real, imag} */,
  {32'h41fdc0a6, 32'hc1fba5a2} /* (1, 20, 11) {real, imag} */,
  {32'h41d5f800, 32'h41801114} /* (1, 20, 10) {real, imag} */,
  {32'h403afe10, 32'h41a57411} /* (1, 20, 9) {real, imag} */,
  {32'h41b58b15, 32'h41be5198} /* (1, 20, 8) {real, imag} */,
  {32'h402c5fe0, 32'h3feb2ab8} /* (1, 20, 7) {real, imag} */,
  {32'h3fa2166c, 32'h42a25958} /* (1, 20, 6) {real, imag} */,
  {32'h41112b06, 32'hc28b6376} /* (1, 20, 5) {real, imag} */,
  {32'hc1acd018, 32'hc2140de8} /* (1, 20, 4) {real, imag} */,
  {32'hc1dd4110, 32'h41244324} /* (1, 20, 3) {real, imag} */,
  {32'h40113c88, 32'hc0d8a20e} /* (1, 20, 2) {real, imag} */,
  {32'h42ca29b6, 32'hc218dc6d} /* (1, 20, 1) {real, imag} */,
  {32'hc3030c94, 32'h42b3813a} /* (1, 20, 0) {real, imag} */,
  {32'h428dd743, 32'hc28ef763} /* (1, 19, 31) {real, imag} */,
  {32'hc006cdb8, 32'hc1c5d4b2} /* (1, 19, 30) {real, imag} */,
  {32'h42011367, 32'h421d3626} /* (1, 19, 29) {real, imag} */,
  {32'hc2805749, 32'h4104308f} /* (1, 19, 28) {real, imag} */,
  {32'hc21b6b67, 32'hc275d11c} /* (1, 19, 27) {real, imag} */,
  {32'h414a7fde, 32'h41700fa8} /* (1, 19, 26) {real, imag} */,
  {32'h405b5458, 32'h411c4c70} /* (1, 19, 25) {real, imag} */,
  {32'hc100a85d, 32'h416915e8} /* (1, 19, 24) {real, imag} */,
  {32'h41d5119d, 32'h4209b39c} /* (1, 19, 23) {real, imag} */,
  {32'hc1a1407f, 32'h41b821db} /* (1, 19, 22) {real, imag} */,
  {32'h40cb2416, 32'hc1b15d90} /* (1, 19, 21) {real, imag} */,
  {32'h41472753, 32'hc129a27a} /* (1, 19, 20) {real, imag} */,
  {32'hc1c6f232, 32'hc10cae89} /* (1, 19, 19) {real, imag} */,
  {32'hc123d96a, 32'hbeec4ba0} /* (1, 19, 18) {real, imag} */,
  {32'h41343bd6, 32'h40d1e390} /* (1, 19, 17) {real, imag} */,
  {32'hc0639600, 32'h40de10ca} /* (1, 19, 16) {real, imag} */,
  {32'hc02fd34a, 32'h41404c78} /* (1, 19, 15) {real, imag} */,
  {32'hc103dc36, 32'h41686a0d} /* (1, 19, 14) {real, imag} */,
  {32'hc0bc6e92, 32'h3ea3e460} /* (1, 19, 13) {real, imag} */,
  {32'hc14081e7, 32'h4041b49f} /* (1, 19, 12) {real, imag} */,
  {32'hc01f1304, 32'hc038cf0c} /* (1, 19, 11) {real, imag} */,
  {32'h41af7133, 32'h41f1999f} /* (1, 19, 10) {real, imag} */,
  {32'hc178b59e, 32'h41886482} /* (1, 19, 9) {real, imag} */,
  {32'h4143b79d, 32'hc1f06712} /* (1, 19, 8) {real, imag} */,
  {32'h42120d7c, 32'hc29831c2} /* (1, 19, 7) {real, imag} */,
  {32'h4293169d, 32'h41c7ba9a} /* (1, 19, 6) {real, imag} */,
  {32'h410d0ad5, 32'h41992611} /* (1, 19, 5) {real, imag} */,
  {32'hc0db5110, 32'h414e75b5} /* (1, 19, 4) {real, imag} */,
  {32'hc198cdd4, 32'hc1ac950a} /* (1, 19, 3) {real, imag} */,
  {32'hc1bb3779, 32'hc1eab69e} /* (1, 19, 2) {real, imag} */,
  {32'hc26401bd, 32'h42933a7f} /* (1, 19, 1) {real, imag} */,
  {32'hc2436a57, 32'h41083867} /* (1, 19, 0) {real, imag} */,
  {32'h42c4b779, 32'hc20fe765} /* (1, 18, 31) {real, imag} */,
  {32'hc15d3084, 32'hc1cdb03a} /* (1, 18, 30) {real, imag} */,
  {32'h421b9850, 32'h3f9bb590} /* (1, 18, 29) {real, imag} */,
  {32'hc23d840e, 32'hc1763211} /* (1, 18, 28) {real, imag} */,
  {32'hc218cbb4, 32'h416fadd7} /* (1, 18, 27) {real, imag} */,
  {32'hc122da1f, 32'hc1ef14b8} /* (1, 18, 26) {real, imag} */,
  {32'hc1b82442, 32'hc2037826} /* (1, 18, 25) {real, imag} */,
  {32'hc08ff580, 32'h414e2dbc} /* (1, 18, 24) {real, imag} */,
  {32'h420e531b, 32'hbf4338d0} /* (1, 18, 23) {real, imag} */,
  {32'hc1a544be, 32'h3e33c2c0} /* (1, 18, 22) {real, imag} */,
  {32'hc045394e, 32'h41c94fb0} /* (1, 18, 21) {real, imag} */,
  {32'hc178110c, 32'hc02e68cc} /* (1, 18, 20) {real, imag} */,
  {32'h41367d5d, 32'hc09a9158} /* (1, 18, 19) {real, imag} */,
  {32'hc11ea98a, 32'h417f9220} /* (1, 18, 18) {real, imag} */,
  {32'hc02945f4, 32'hc104fdea} /* (1, 18, 17) {real, imag} */,
  {32'h40e99c08, 32'h41432fe6} /* (1, 18, 16) {real, imag} */,
  {32'hc1814ffa, 32'h3fa45c0c} /* (1, 18, 15) {real, imag} */,
  {32'h3f8aa420, 32'h3f35f7f8} /* (1, 18, 14) {real, imag} */,
  {32'h41719f6d, 32'hc059c710} /* (1, 18, 13) {real, imag} */,
  {32'h3ce8a900, 32'h41748f6d} /* (1, 18, 12) {real, imag} */,
  {32'h402e05ee, 32'hc1b96590} /* (1, 18, 11) {real, imag} */,
  {32'h3f7e3f30, 32'h40895292} /* (1, 18, 10) {real, imag} */,
  {32'hc21650d9, 32'h4179350f} /* (1, 18, 9) {real, imag} */,
  {32'h41f89aca, 32'hc24a80cf} /* (1, 18, 8) {real, imag} */,
  {32'h41983a2e, 32'hc081111c} /* (1, 18, 7) {real, imag} */,
  {32'hc1e540e4, 32'h3fea04f8} /* (1, 18, 6) {real, imag} */,
  {32'hc19cfd9f, 32'hc096e4c6} /* (1, 18, 5) {real, imag} */,
  {32'hc09546a0, 32'h4228358e} /* (1, 18, 4) {real, imag} */,
  {32'hc13cf097, 32'h4248bc6c} /* (1, 18, 3) {real, imag} */,
  {32'hc1b6d492, 32'hc1ecca9e} /* (1, 18, 2) {real, imag} */,
  {32'h428be489, 32'h42516ef3} /* (1, 18, 1) {real, imag} */,
  {32'h42747193, 32'h41ffb631} /* (1, 18, 0) {real, imag} */,
  {32'hc125ef08, 32'hc16780f5} /* (1, 17, 31) {real, imag} */,
  {32'hc0eafcfa, 32'hc11c0698} /* (1, 17, 30) {real, imag} */,
  {32'hc1961288, 32'hc11295f2} /* (1, 17, 29) {real, imag} */,
  {32'h41901655, 32'h41483510} /* (1, 17, 28) {real, imag} */,
  {32'hc21b85d8, 32'h40dc5198} /* (1, 17, 27) {real, imag} */,
  {32'h4008c140, 32'hc194b2ac} /* (1, 17, 26) {real, imag} */,
  {32'h4101a2c8, 32'h41921534} /* (1, 17, 25) {real, imag} */,
  {32'hc1d680bf, 32'h4224106e} /* (1, 17, 24) {real, imag} */,
  {32'hc10976b9, 32'hc1a6338a} /* (1, 17, 23) {real, imag} */,
  {32'h40f924de, 32'h4064fd74} /* (1, 17, 22) {real, imag} */,
  {32'h413bad0a, 32'h417b1543} /* (1, 17, 21) {real, imag} */,
  {32'hc1340926, 32'hc057d0c4} /* (1, 17, 20) {real, imag} */,
  {32'h3f892e78, 32'hc11c9a8e} /* (1, 17, 19) {real, imag} */,
  {32'hc15efb1b, 32'hc1055e4a} /* (1, 17, 18) {real, imag} */,
  {32'hbfbd3690, 32'hc00d141c} /* (1, 17, 17) {real, imag} */,
  {32'hc02ce960, 32'h40b7e2b4} /* (1, 17, 16) {real, imag} */,
  {32'hbe734580, 32'hbf960ff8} /* (1, 17, 15) {real, imag} */,
  {32'hc0a1b1ce, 32'h40e75863} /* (1, 17, 14) {real, imag} */,
  {32'h40eed376, 32'h4141fb16} /* (1, 17, 13) {real, imag} */,
  {32'h3f84e1f4, 32'hc11666d4} /* (1, 17, 12) {real, imag} */,
  {32'h40b32f48, 32'h413c36ff} /* (1, 17, 11) {real, imag} */,
  {32'h41b91b34, 32'hc15f459b} /* (1, 17, 10) {real, imag} */,
  {32'hc11f0d53, 32'h420a1459} /* (1, 17, 9) {real, imag} */,
  {32'h421f596e, 32'hbfd63e30} /* (1, 17, 8) {real, imag} */,
  {32'hc138aa56, 32'h41827fb8} /* (1, 17, 7) {real, imag} */,
  {32'h4279d792, 32'hc1a54b50} /* (1, 17, 6) {real, imag} */,
  {32'h41accb58, 32'h41086622} /* (1, 17, 5) {real, imag} */,
  {32'hc2220670, 32'hc1832d86} /* (1, 17, 4) {real, imag} */,
  {32'h41a4fc56, 32'h3f4532f8} /* (1, 17, 3) {real, imag} */,
  {32'h4182232a, 32'h40fce43f} /* (1, 17, 2) {real, imag} */,
  {32'hc257d086, 32'h422109b9} /* (1, 17, 1) {real, imag} */,
  {32'hc284ef19, 32'h412aa3ba} /* (1, 17, 0) {real, imag} */,
  {32'h41f6979e, 32'h416c7048} /* (1, 16, 31) {real, imag} */,
  {32'h41b91719, 32'h4299ace6} /* (1, 16, 30) {real, imag} */,
  {32'h424061b0, 32'h419a23d2} /* (1, 16, 29) {real, imag} */,
  {32'h410ecb32, 32'h405b263c} /* (1, 16, 28) {real, imag} */,
  {32'h407b8358, 32'hc0e9cee5} /* (1, 16, 27) {real, imag} */,
  {32'h4219db56, 32'h41b547ba} /* (1, 16, 26) {real, imag} */,
  {32'hc1597bb1, 32'hc1cc31ac} /* (1, 16, 25) {real, imag} */,
  {32'hc069e614, 32'h4208feb1} /* (1, 16, 24) {real, imag} */,
  {32'hc1ae8e87, 32'h3fa570a0} /* (1, 16, 23) {real, imag} */,
  {32'h3d3c3e40, 32'hc190d0fa} /* (1, 16, 22) {real, imag} */,
  {32'hc169687d, 32'h412d999b} /* (1, 16, 21) {real, imag} */,
  {32'h41590dac, 32'h3eb331f0} /* (1, 16, 20) {real, imag} */,
  {32'hc14e43da, 32'hc0e1be20} /* (1, 16, 19) {real, imag} */,
  {32'hc0eea78e, 32'h416f3338} /* (1, 16, 18) {real, imag} */,
  {32'hbf04c250, 32'hc10960a8} /* (1, 16, 17) {real, imag} */,
  {32'h40973015, 32'hc05d47f2} /* (1, 16, 16) {real, imag} */,
  {32'hc184b0e6, 32'hc16d9278} /* (1, 16, 15) {real, imag} */,
  {32'h410c3e05, 32'h401f78e0} /* (1, 16, 14) {real, imag} */,
  {32'h41235176, 32'hc0fdea08} /* (1, 16, 13) {real, imag} */,
  {32'hc0b9e43b, 32'hc14e9974} /* (1, 16, 12) {real, imag} */,
  {32'h418bbbb5, 32'hc12e4bb9} /* (1, 16, 11) {real, imag} */,
  {32'hbe825a38, 32'h40d1df1e} /* (1, 16, 10) {real, imag} */,
  {32'h41cd6721, 32'h3fd34a70} /* (1, 16, 9) {real, imag} */,
  {32'h41c1283c, 32'hc1a2f2af} /* (1, 16, 8) {real, imag} */,
  {32'hc0820f8e, 32'hc15cd2b7} /* (1, 16, 7) {real, imag} */,
  {32'hc1c22903, 32'hc022d85c} /* (1, 16, 6) {real, imag} */,
  {32'hc1aa7b26, 32'hc1219f2c} /* (1, 16, 5) {real, imag} */,
  {32'hc17a58c8, 32'h419d1d48} /* (1, 16, 4) {real, imag} */,
  {32'hc1d39fab, 32'h4120bec3} /* (1, 16, 3) {real, imag} */,
  {32'hc1a3d771, 32'hc18770ee} /* (1, 16, 2) {real, imag} */,
  {32'h42098b9d, 32'h4149784c} /* (1, 16, 1) {real, imag} */,
  {32'hc0efd7e7, 32'hc122cc3e} /* (1, 16, 0) {real, imag} */,
  {32'h40a44d70, 32'hc1b6d400} /* (1, 15, 31) {real, imag} */,
  {32'hc19b260b, 32'hc013c058} /* (1, 15, 30) {real, imag} */,
  {32'hc0d2cf34, 32'hc20a933c} /* (1, 15, 29) {real, imag} */,
  {32'h417b565d, 32'hc2405243} /* (1, 15, 28) {real, imag} */,
  {32'h4208a31f, 32'hc235e92c} /* (1, 15, 27) {real, imag} */,
  {32'h41ea49fc, 32'hc0303fe0} /* (1, 15, 26) {real, imag} */,
  {32'h3fccbed8, 32'h42248f7b} /* (1, 15, 25) {real, imag} */,
  {32'hc03f78c0, 32'h3fed7940} /* (1, 15, 24) {real, imag} */,
  {32'hbfd2a920, 32'h40ba87d2} /* (1, 15, 23) {real, imag} */,
  {32'hc1a64b0a, 32'h4221c772} /* (1, 15, 22) {real, imag} */,
  {32'h41e5df86, 32'h41f12692} /* (1, 15, 21) {real, imag} */,
  {32'h4095aa5c, 32'h418e2483} /* (1, 15, 20) {real, imag} */,
  {32'hc1103ca9, 32'hc11e5e0a} /* (1, 15, 19) {real, imag} */,
  {32'h3fca4330, 32'hc0833d12} /* (1, 15, 18) {real, imag} */,
  {32'hc037f29c, 32'h3f8786e8} /* (1, 15, 17) {real, imag} */,
  {32'h413d7e54, 32'hc0c15354} /* (1, 15, 16) {real, imag} */,
  {32'hbf4dd690, 32'h40d946c6} /* (1, 15, 15) {real, imag} */,
  {32'hc0204738, 32'h4062f9c0} /* (1, 15, 14) {real, imag} */,
  {32'hc151767d, 32'hc118cc7a} /* (1, 15, 13) {real, imag} */,
  {32'hbf4194c4, 32'hc098517f} /* (1, 15, 12) {real, imag} */,
  {32'h3f17f270, 32'hc04637c0} /* (1, 15, 11) {real, imag} */,
  {32'hbe4e1c40, 32'hc166a1c7} /* (1, 15, 10) {real, imag} */,
  {32'hc19fd84e, 32'hc133413f} /* (1, 15, 9) {real, imag} */,
  {32'hc1d3c668, 32'hc1a6f96a} /* (1, 15, 8) {real, imag} */,
  {32'h41249155, 32'h4190ee16} /* (1, 15, 7) {real, imag} */,
  {32'h41705ed8, 32'h412f18a6} /* (1, 15, 6) {real, imag} */,
  {32'hc160c559, 32'h4187aa36} /* (1, 15, 5) {real, imag} */,
  {32'h41b4da1a, 32'h4131fb9c} /* (1, 15, 4) {real, imag} */,
  {32'hc1a72d96, 32'hc2513974} /* (1, 15, 3) {real, imag} */,
  {32'hc22ac71a, 32'h41f4a56f} /* (1, 15, 2) {real, imag} */,
  {32'h4277127e, 32'h40c93f96} /* (1, 15, 1) {real, imag} */,
  {32'h4176f21c, 32'hc1db9551} /* (1, 15, 0) {real, imag} */,
  {32'hc2e2a071, 32'hc20fd614} /* (1, 14, 31) {real, imag} */,
  {32'h3ff2d938, 32'hc2019d40} /* (1, 14, 30) {real, imag} */,
  {32'h4191496b, 32'hc0dd68fc} /* (1, 14, 29) {real, imag} */,
  {32'h4178b0cd, 32'h4209a0ef} /* (1, 14, 28) {real, imag} */,
  {32'h41b26e32, 32'h4202c892} /* (1, 14, 27) {real, imag} */,
  {32'hc0ed7900, 32'hc19ec8eb} /* (1, 14, 26) {real, imag} */,
  {32'hc187d04d, 32'h4016baec} /* (1, 14, 25) {real, imag} */,
  {32'h3f35d060, 32'hc139117d} /* (1, 14, 24) {real, imag} */,
  {32'hc1ba4c99, 32'h4181545c} /* (1, 14, 23) {real, imag} */,
  {32'h401771b8, 32'h406be576} /* (1, 14, 22) {real, imag} */,
  {32'h4114668f, 32'hc18b524b} /* (1, 14, 21) {real, imag} */,
  {32'hbf31d620, 32'hc1a909c6} /* (1, 14, 20) {real, imag} */,
  {32'hc0f6bfec, 32'hc10d1a0e} /* (1, 14, 19) {real, imag} */,
  {32'hc0c5e6be, 32'h4117935e} /* (1, 14, 18) {real, imag} */,
  {32'hbff8dd14, 32'h40581d42} /* (1, 14, 17) {real, imag} */,
  {32'h409253cc, 32'h3ff2faa0} /* (1, 14, 16) {real, imag} */,
  {32'h411f791a, 32'hbefa0a10} /* (1, 14, 15) {real, imag} */,
  {32'h4189f15c, 32'hbfd02bd0} /* (1, 14, 14) {real, imag} */,
  {32'hc12c196a, 32'h40421708} /* (1, 14, 13) {real, imag} */,
  {32'h4028de50, 32'h40fe8608} /* (1, 14, 12) {real, imag} */,
  {32'h4075da64, 32'h416f9b2e} /* (1, 14, 11) {real, imag} */,
  {32'hc1b21411, 32'h40b1dafb} /* (1, 14, 10) {real, imag} */,
  {32'h40047168, 32'h411eeba1} /* (1, 14, 9) {real, imag} */,
  {32'hc13eee4a, 32'h4089bd9a} /* (1, 14, 8) {real, imag} */,
  {32'hc22b065c, 32'h417748c3} /* (1, 14, 7) {real, imag} */,
  {32'h423ad4d2, 32'h4241957e} /* (1, 14, 6) {real, imag} */,
  {32'h42919716, 32'hc017a030} /* (1, 14, 5) {real, imag} */,
  {32'hc215f331, 32'h418eeaca} /* (1, 14, 4) {real, imag} */,
  {32'hc15d4d72, 32'h42480060} /* (1, 14, 3) {real, imag} */,
  {32'h41b11154, 32'hc121aa1c} /* (1, 14, 2) {real, imag} */,
  {32'hc2c7efb7, 32'hc24420fa} /* (1, 14, 1) {real, imag} */,
  {32'hc28496a8, 32'hc29175da} /* (1, 14, 0) {real, imag} */,
  {32'hc2f2207f, 32'hc24b6ed2} /* (1, 13, 31) {real, imag} */,
  {32'h42b4bc7c, 32'hc26cfcd7} /* (1, 13, 30) {real, imag} */,
  {32'h42111167, 32'h40a708ac} /* (1, 13, 29) {real, imag} */,
  {32'h422cca1a, 32'hc14da4ee} /* (1, 13, 28) {real, imag} */,
  {32'hc1ddfae1, 32'h428794a8} /* (1, 13, 27) {real, imag} */,
  {32'h4279b68c, 32'hc1bd6c24} /* (1, 13, 26) {real, imag} */,
  {32'hc2024fe1, 32'hc13d6834} /* (1, 13, 25) {real, imag} */,
  {32'h41311b70, 32'hbf967930} /* (1, 13, 24) {real, imag} */,
  {32'hc0ed28a6, 32'h424aa31b} /* (1, 13, 23) {real, imag} */,
  {32'hc181a8d4, 32'hc1a3fbee} /* (1, 13, 22) {real, imag} */,
  {32'hc189d3ba, 32'h407505e8} /* (1, 13, 21) {real, imag} */,
  {32'hc18f2c7c, 32'h41ce15c2} /* (1, 13, 20) {real, imag} */,
  {32'hc11338a5, 32'hc0ff35d8} /* (1, 13, 19) {real, imag} */,
  {32'h4035b89c, 32'h3fbcf35c} /* (1, 13, 18) {real, imag} */,
  {32'hc0694eec, 32'hc0de5447} /* (1, 13, 17) {real, imag} */,
  {32'h3eeac6c0, 32'h415afd30} /* (1, 13, 16) {real, imag} */,
  {32'hc14b414b, 32'hc156573c} /* (1, 13, 15) {real, imag} */,
  {32'h4190b7a2, 32'h41859dce} /* (1, 13, 14) {real, imag} */,
  {32'h41aef196, 32'hc15c3bc0} /* (1, 13, 13) {real, imag} */,
  {32'h4098f4c6, 32'h40fd4136} /* (1, 13, 12) {real, imag} */,
  {32'h40c4dd14, 32'h409b92cc} /* (1, 13, 11) {real, imag} */,
  {32'hc145d67b, 32'h40fad942} /* (1, 13, 10) {real, imag} */,
  {32'hc196b422, 32'h400df850} /* (1, 13, 9) {real, imag} */,
  {32'hc253a692, 32'h420a8ef8} /* (1, 13, 8) {real, imag} */,
  {32'hc0c9928a, 32'h420ac519} /* (1, 13, 7) {real, imag} */,
  {32'hc26c52d4, 32'hc22c5876} /* (1, 13, 6) {real, imag} */,
  {32'hc0593d80, 32'h40e18578} /* (1, 13, 5) {real, imag} */,
  {32'hc0dec014, 32'h40132782} /* (1, 13, 4) {real, imag} */,
  {32'h41c0eedd, 32'h421ef386} /* (1, 13, 3) {real, imag} */,
  {32'hc12ea184, 32'hc2550303} /* (1, 13, 2) {real, imag} */,
  {32'h42d60461, 32'hc252522a} /* (1, 13, 1) {real, imag} */,
  {32'h422de2fc, 32'h41c37504} /* (1, 13, 0) {real, imag} */,
  {32'h428eb778, 32'hc2b68df2} /* (1, 12, 31) {real, imag} */,
  {32'hc0293c60, 32'h4145c6c3} /* (1, 12, 30) {real, imag} */,
  {32'h411cdab6, 32'hc255f2c5} /* (1, 12, 29) {real, imag} */,
  {32'h4028b070, 32'h41bb93f0} /* (1, 12, 28) {real, imag} */,
  {32'h41f6b204, 32'h420a5836} /* (1, 12, 27) {real, imag} */,
  {32'hc180bab6, 32'h4016d16c} /* (1, 12, 26) {real, imag} */,
  {32'hc2698472, 32'hc270a582} /* (1, 12, 25) {real, imag} */,
  {32'hc2433869, 32'hc1851ece} /* (1, 12, 24) {real, imag} */,
  {32'h412d854e, 32'h423afbce} /* (1, 12, 23) {real, imag} */,
  {32'h41ec31d7, 32'hc085ee4c} /* (1, 12, 22) {real, imag} */,
  {32'h41a0b3a0, 32'h405c677e} /* (1, 12, 21) {real, imag} */,
  {32'hc18b05e8, 32'h40de5688} /* (1, 12, 20) {real, imag} */,
  {32'hc0958a32, 32'h40d23f3a} /* (1, 12, 19) {real, imag} */,
  {32'h40ceaeca, 32'hc1147098} /* (1, 12, 18) {real, imag} */,
  {32'hc1146eda, 32'h417824b7} /* (1, 12, 17) {real, imag} */,
  {32'hc0dabad4, 32'hbe913760} /* (1, 12, 16) {real, imag} */,
  {32'hc0b7f6b4, 32'h41511771} /* (1, 12, 15) {real, imag} */,
  {32'h3ff0b960, 32'h40a3a71b} /* (1, 12, 14) {real, imag} */,
  {32'hbfe47798, 32'h4186fce6} /* (1, 12, 13) {real, imag} */,
  {32'hc0c375b8, 32'h40e12750} /* (1, 12, 12) {real, imag} */,
  {32'hc1da9f96, 32'hc181605a} /* (1, 12, 11) {real, imag} */,
  {32'hc0a6bbfc, 32'hc231d5a4} /* (1, 12, 10) {real, imag} */,
  {32'h421adf06, 32'hc287c9b9} /* (1, 12, 9) {real, imag} */,
  {32'hc22db9e7, 32'h3f23fbc8} /* (1, 12, 8) {real, imag} */,
  {32'hc181c80f, 32'h420d510a} /* (1, 12, 7) {real, imag} */,
  {32'h41bda31c, 32'h3f4dac10} /* (1, 12, 6) {real, imag} */,
  {32'hbfade358, 32'hc26175e6} /* (1, 12, 5) {real, imag} */,
  {32'hc1b2b2a8, 32'h41007c9c} /* (1, 12, 4) {real, imag} */,
  {32'h410590aa, 32'h427ffcb9} /* (1, 12, 3) {real, imag} */,
  {32'h41b3c308, 32'hc1e31ed0} /* (1, 12, 2) {real, imag} */,
  {32'hc28b8a2c, 32'hc22640cb} /* (1, 12, 1) {real, imag} */,
  {32'h4241e4cc, 32'h41870442} /* (1, 12, 0) {real, imag} */,
  {32'hc19646e0, 32'h430e093a} /* (1, 11, 31) {real, imag} */,
  {32'h42cdcf1d, 32'hc2c3f802} /* (1, 11, 30) {real, imag} */,
  {32'h40b354fc, 32'h42862c54} /* (1, 11, 29) {real, imag} */,
  {32'h41ba1ae2, 32'hc110126f} /* (1, 11, 28) {real, imag} */,
  {32'hc0881754, 32'hc2a7b84e} /* (1, 11, 27) {real, imag} */,
  {32'h41ae376f, 32'h40e97dac} /* (1, 11, 26) {real, imag} */,
  {32'hc14b00fa, 32'h42a9f242} /* (1, 11, 25) {real, imag} */,
  {32'hc0ecbdb3, 32'hc0d71a68} /* (1, 11, 24) {real, imag} */,
  {32'hc04a0130, 32'h4210e139} /* (1, 11, 23) {real, imag} */,
  {32'hc213e61b, 32'h418f1fbd} /* (1, 11, 22) {real, imag} */,
  {32'h41644246, 32'hc1df5f68} /* (1, 11, 21) {real, imag} */,
  {32'h41441d6a, 32'hc1278238} /* (1, 11, 20) {real, imag} */,
  {32'hc0ff13e3, 32'h40441dd4} /* (1, 11, 19) {real, imag} */,
  {32'hc0c4ac32, 32'hbeac0020} /* (1, 11, 18) {real, imag} */,
  {32'h40a82e30, 32'hc1231d44} /* (1, 11, 17) {real, imag} */,
  {32'h413e3f90, 32'hbec713f0} /* (1, 11, 16) {real, imag} */,
  {32'hc108b458, 32'hc173777c} /* (1, 11, 15) {real, imag} */,
  {32'h410ed309, 32'hc0bc9cf2} /* (1, 11, 14) {real, imag} */,
  {32'hc190e9f7, 32'hc08ecd62} /* (1, 11, 13) {real, imag} */,
  {32'hbfafb5a0, 32'hbf9ba914} /* (1, 11, 12) {real, imag} */,
  {32'hc124eefe, 32'h4207eb66} /* (1, 11, 11) {real, imag} */,
  {32'hc1a1b892, 32'h4236bc46} /* (1, 11, 10) {real, imag} */,
  {32'hc19de350, 32'hc13a3f43} /* (1, 11, 9) {real, imag} */,
  {32'h409ed5d3, 32'hc2019452} /* (1, 11, 8) {real, imag} */,
  {32'hbfd48870, 32'hc1966c2a} /* (1, 11, 7) {real, imag} */,
  {32'hc1cd4165, 32'hc22fc008} /* (1, 11, 6) {real, imag} */,
  {32'h42074e18, 32'h419d220e} /* (1, 11, 5) {real, imag} */,
  {32'hc253304d, 32'hc1d2de78} /* (1, 11, 4) {real, imag} */,
  {32'h41ee98a9, 32'h41d9adca} /* (1, 11, 3) {real, imag} */,
  {32'h42a43401, 32'h4277ad3b} /* (1, 11, 2) {real, imag} */,
  {32'hc304efa7, 32'h424b3317} /* (1, 11, 1) {real, imag} */,
  {32'hc2e00824, 32'h40e2f4ef} /* (1, 11, 0) {real, imag} */,
  {32'h42a1f924, 32'hc255dd35} /* (1, 10, 31) {real, imag} */,
  {32'hc2d87b5b, 32'h42d562ca} /* (1, 10, 30) {real, imag} */,
  {32'h421f50ab, 32'h42a0e393} /* (1, 10, 29) {real, imag} */,
  {32'h42636854, 32'hc28ee754} /* (1, 10, 28) {real, imag} */,
  {32'h42d69fea, 32'hc13b80d4} /* (1, 10, 27) {real, imag} */,
  {32'h424c6d40, 32'hc2862900} /* (1, 10, 26) {real, imag} */,
  {32'h41af071e, 32'hc131bc86} /* (1, 10, 25) {real, imag} */,
  {32'h412f56e4, 32'hc19eabdd} /* (1, 10, 24) {real, imag} */,
  {32'hc2402403, 32'hc221be2d} /* (1, 10, 23) {real, imag} */,
  {32'h42000927, 32'h408d4248} /* (1, 10, 22) {real, imag} */,
  {32'hc24215eb, 32'hc1fa71e7} /* (1, 10, 21) {real, imag} */,
  {32'hc0d28038, 32'h423d0f89} /* (1, 10, 20) {real, imag} */,
  {32'h420de142, 32'h4182fa3a} /* (1, 10, 19) {real, imag} */,
  {32'hc10128bd, 32'h40cd123c} /* (1, 10, 18) {real, imag} */,
  {32'hc15f9ed6, 32'hc19e2d30} /* (1, 10, 17) {real, imag} */,
  {32'h41467746, 32'h4117d14d} /* (1, 10, 16) {real, imag} */,
  {32'h41fa5521, 32'hc102a849} /* (1, 10, 15) {real, imag} */,
  {32'h40a3a82a, 32'h40e9046c} /* (1, 10, 14) {real, imag} */,
  {32'h4024b0e0, 32'h40c474de} /* (1, 10, 13) {real, imag} */,
  {32'h3fddf8a0, 32'hc1da2302} /* (1, 10, 12) {real, imag} */,
  {32'hc1eba776, 32'hc22074ae} /* (1, 10, 11) {real, imag} */,
  {32'hc1be5216, 32'h421a2037} /* (1, 10, 10) {real, imag} */,
  {32'h4186dca2, 32'h3d11a400} /* (1, 10, 9) {real, imag} */,
  {32'h4085ca34, 32'hc23ae7aa} /* (1, 10, 8) {real, imag} */,
  {32'h4267590b, 32'h3fafa060} /* (1, 10, 7) {real, imag} */,
  {32'h42303f0c, 32'hc1f29432} /* (1, 10, 6) {real, imag} */,
  {32'hc2c22bee, 32'hc2b42088} /* (1, 10, 5) {real, imag} */,
  {32'h42a85f56, 32'h41dd0c14} /* (1, 10, 4) {real, imag} */,
  {32'h42487475, 32'h3e834500} /* (1, 10, 3) {real, imag} */,
  {32'hc2f2b96d, 32'hc1817f56} /* (1, 10, 2) {real, imag} */,
  {32'h425a6777, 32'hc2ba254a} /* (1, 10, 1) {real, imag} */,
  {32'h41ef7455, 32'hc1d97a7e} /* (1, 10, 0) {real, imag} */,
  {32'h424e4433, 32'h42bb9f4a} /* (1, 9, 31) {real, imag} */,
  {32'hc1c3468d, 32'hc06de730} /* (1, 9, 30) {real, imag} */,
  {32'hc2b00d74, 32'hc0937d34} /* (1, 9, 29) {real, imag} */,
  {32'hc188c80a, 32'hc1e37712} /* (1, 9, 28) {real, imag} */,
  {32'h4207a0fe, 32'h42c3eb28} /* (1, 9, 27) {real, imag} */,
  {32'hc1f09665, 32'hc2ddc9cd} /* (1, 9, 26) {real, imag} */,
  {32'hc1448d64, 32'h40a78bea} /* (1, 9, 25) {real, imag} */,
  {32'hc223bda6, 32'hc208c2cc} /* (1, 9, 24) {real, imag} */,
  {32'hc1d50526, 32'hc24145b0} /* (1, 9, 23) {real, imag} */,
  {32'hc1a002a6, 32'hc1885af4} /* (1, 9, 22) {real, imag} */,
  {32'h407e1b50, 32'hc1b3e658} /* (1, 9, 21) {real, imag} */,
  {32'h41da9b23, 32'hc13a7cca} /* (1, 9, 20) {real, imag} */,
  {32'hc21200f2, 32'h41a13c92} /* (1, 9, 19) {real, imag} */,
  {32'hc082d1c8, 32'h41b76ea5} /* (1, 9, 18) {real, imag} */,
  {32'h42123726, 32'hc19c849b} /* (1, 9, 17) {real, imag} */,
  {32'h42414cfe, 32'hc0736ee0} /* (1, 9, 16) {real, imag} */,
  {32'hc0deee40, 32'h422bcfd4} /* (1, 9, 15) {real, imag} */,
  {32'hc200eb3a, 32'h416faa3e} /* (1, 9, 14) {real, imag} */,
  {32'hbe16b380, 32'hc179b3bc} /* (1, 9, 13) {real, imag} */,
  {32'h410e7bae, 32'h418a5c59} /* (1, 9, 12) {real, imag} */,
  {32'hc21df98b, 32'hc12b5e18} /* (1, 9, 11) {real, imag} */,
  {32'hc17de771, 32'hc1b44600} /* (1, 9, 10) {real, imag} */,
  {32'h410f0604, 32'h4121119e} /* (1, 9, 9) {real, imag} */,
  {32'h41e0365c, 32'h40115278} /* (1, 9, 8) {real, imag} */,
  {32'h4296ab8e, 32'hc1b04e34} /* (1, 9, 7) {real, imag} */,
  {32'h40ce164c, 32'h42c697a3} /* (1, 9, 6) {real, imag} */,
  {32'hc2c14421, 32'h42a77ef0} /* (1, 9, 5) {real, imag} */,
  {32'h42a46d48, 32'h41ca7db0} /* (1, 9, 4) {real, imag} */,
  {32'h4120e8bc, 32'hc1e28043} /* (1, 9, 3) {real, imag} */,
  {32'hc28ee069, 32'hc2f40aae} /* (1, 9, 2) {real, imag} */,
  {32'h4300b88f, 32'hc26ee25d} /* (1, 9, 1) {real, imag} */,
  {32'hc3452506, 32'h429a2a7b} /* (1, 9, 0) {real, imag} */,
  {32'hc341e188, 32'h4388f062} /* (1, 8, 31) {real, imag} */,
  {32'h42319f12, 32'hc3140f39} /* (1, 8, 30) {real, imag} */,
  {32'h41ee5f69, 32'h422e453f} /* (1, 8, 29) {real, imag} */,
  {32'h422d8761, 32'hc22c64a4} /* (1, 8, 28) {real, imag} */,
  {32'hc27133ec, 32'hc38fe8f2} /* (1, 8, 27) {real, imag} */,
  {32'h428718a4, 32'hc1fd1de6} /* (1, 8, 26) {real, imag} */,
  {32'h427440bb, 32'h4290e3a9} /* (1, 8, 25) {real, imag} */,
  {32'hc15d1198, 32'h42a72a15} /* (1, 8, 24) {real, imag} */,
  {32'hc154f35a, 32'hc20b6ace} /* (1, 8, 23) {real, imag} */,
  {32'h420785ed, 32'hc21e6c16} /* (1, 8, 22) {real, imag} */,
  {32'h41d5578e, 32'hc117bd44} /* (1, 8, 21) {real, imag} */,
  {32'h40341030, 32'hc1de7a08} /* (1, 8, 20) {real, imag} */,
  {32'h408cad2c, 32'h4165c9d3} /* (1, 8, 19) {real, imag} */,
  {32'hbfb6a734, 32'hc244c38a} /* (1, 8, 18) {real, imag} */,
  {32'h41645777, 32'h420c1152} /* (1, 8, 17) {real, imag} */,
  {32'h41a432fc, 32'hc1cf8da0} /* (1, 8, 16) {real, imag} */,
  {32'h4192a7f4, 32'h41cbb3c5} /* (1, 8, 15) {real, imag} */,
  {32'hc08badd3, 32'h3fb8a840} /* (1, 8, 14) {real, imag} */,
  {32'h4227db64, 32'h41637ecd} /* (1, 8, 13) {real, imag} */,
  {32'hc14460a4, 32'hc1ef9dc4} /* (1, 8, 12) {real, imag} */,
  {32'hc208a511, 32'h41f810ba} /* (1, 8, 11) {real, imag} */,
  {32'h41a7b7a6, 32'hc21e1118} /* (1, 8, 10) {real, imag} */,
  {32'h42355328, 32'h41f9132d} /* (1, 8, 9) {real, imag} */,
  {32'h42ac586f, 32'hc29f9ebb} /* (1, 8, 8) {real, imag} */,
  {32'h429efa44, 32'h4219b3fe} /* (1, 8, 7) {real, imag} */,
  {32'hc2e57110, 32'h422cbbb5} /* (1, 8, 6) {real, imag} */,
  {32'h42c3dd96, 32'hc1fa3858} /* (1, 8, 5) {real, imag} */,
  {32'hc307f4ef, 32'h433296ab} /* (1, 8, 4) {real, imag} */,
  {32'hc14025ca, 32'h40f4f228} /* (1, 8, 3) {real, imag} */,
  {32'h429bee5f, 32'hc360a0c1} /* (1, 8, 2) {real, imag} */,
  {32'hc31045fa, 32'h43087120} /* (1, 8, 1) {real, imag} */,
  {32'hc2eba7dd, 32'h42ee221e} /* (1, 8, 0) {real, imag} */,
  {32'h41a3916c, 32'hc2f64628} /* (1, 7, 31) {real, imag} */,
  {32'hc31c3aa2, 32'h431d68a2} /* (1, 7, 30) {real, imag} */,
  {32'h41e47f5c, 32'h42bf1342} /* (1, 7, 29) {real, imag} */,
  {32'hc2a6bcdc, 32'h41b1b8eb} /* (1, 7, 28) {real, imag} */,
  {32'h41180928, 32'hc142b73e} /* (1, 7, 27) {real, imag} */,
  {32'h42497c81, 32'h4130da7c} /* (1, 7, 26) {real, imag} */,
  {32'hc1eda525, 32'hc1de9bd9} /* (1, 7, 25) {real, imag} */,
  {32'hc1b7bfe5, 32'h41ea80b8} /* (1, 7, 24) {real, imag} */,
  {32'hc28f01cd, 32'h43083f10} /* (1, 7, 23) {real, imag} */,
  {32'h42053ccb, 32'hc228d0c5} /* (1, 7, 22) {real, imag} */,
  {32'h4134756c, 32'h41a73cf8} /* (1, 7, 21) {real, imag} */,
  {32'hc1a4d03c, 32'hc1c5a7b1} /* (1, 7, 20) {real, imag} */,
  {32'h418f3ebb, 32'hc0d23174} /* (1, 7, 19) {real, imag} */,
  {32'hc19df544, 32'hc1a2f7f8} /* (1, 7, 18) {real, imag} */,
  {32'h416d6560, 32'h412cb390} /* (1, 7, 17) {real, imag} */,
  {32'h41cb9550, 32'h4123cc70} /* (1, 7, 16) {real, imag} */,
  {32'h406a60c0, 32'h4000f2c2} /* (1, 7, 15) {real, imag} */,
  {32'hc1223dd9, 32'hc1ded4e0} /* (1, 7, 14) {real, imag} */,
  {32'hc08822a4, 32'h426aba3e} /* (1, 7, 13) {real, imag} */,
  {32'hc22c496e, 32'h411b638e} /* (1, 7, 12) {real, imag} */,
  {32'hc1a8bec0, 32'hc25b007c} /* (1, 7, 11) {real, imag} */,
  {32'h42320cdd, 32'hc2b160b4} /* (1, 7, 10) {real, imag} */,
  {32'h430e6762, 32'h41fa55ec} /* (1, 7, 9) {real, imag} */,
  {32'h41c22c35, 32'h4228dfb0} /* (1, 7, 8) {real, imag} */,
  {32'h427dbfb6, 32'hc2443134} /* (1, 7, 7) {real, imag} */,
  {32'hc2392445, 32'h4247d89d} /* (1, 7, 6) {real, imag} */,
  {32'h42d65881, 32'hc1e549c5} /* (1, 7, 5) {real, imag} */,
  {32'h427019fc, 32'hc045f1e8} /* (1, 7, 4) {real, imag} */,
  {32'hc2020058, 32'h4291487e} /* (1, 7, 3) {real, imag} */,
  {32'hc3330734, 32'h42bf21fe} /* (1, 7, 2) {real, imag} */,
  {32'h4389e06f, 32'hc2b026b4} /* (1, 7, 1) {real, imag} */,
  {32'h434464ac, 32'hc27057d4} /* (1, 7, 0) {real, imag} */,
  {32'hc2960809, 32'h429c3448} /* (1, 6, 31) {real, imag} */,
  {32'hc307a412, 32'hc000b6f8} /* (1, 6, 30) {real, imag} */,
  {32'h42b6e28a, 32'hc1bd9dfc} /* (1, 6, 29) {real, imag} */,
  {32'hc2bd807f, 32'h414ee570} /* (1, 6, 28) {real, imag} */,
  {32'h42a4f2cd, 32'hc2c56e33} /* (1, 6, 27) {real, imag} */,
  {32'h41b60438, 32'hc294a5b1} /* (1, 6, 26) {real, imag} */,
  {32'h4201c5d7, 32'h420a9d40} /* (1, 6, 25) {real, imag} */,
  {32'h4275a856, 32'h42c2d044} /* (1, 6, 24) {real, imag} */,
  {32'hc24381a6, 32'hc2c9d879} /* (1, 6, 23) {real, imag} */,
  {32'hc017d62c, 32'hc1633ee6} /* (1, 6, 22) {real, imag} */,
  {32'hc18f8bba, 32'hc28a7da2} /* (1, 6, 21) {real, imag} */,
  {32'hc0510cb0, 32'h42603589} /* (1, 6, 20) {real, imag} */,
  {32'h422b4863, 32'hc24b79b2} /* (1, 6, 19) {real, imag} */,
  {32'h410e0ce8, 32'h418ad092} /* (1, 6, 18) {real, imag} */,
  {32'hc202a836, 32'h41c9b2e8} /* (1, 6, 17) {real, imag} */,
  {32'h41c35420, 32'h412074de} /* (1, 6, 16) {real, imag} */,
  {32'hc21f8e86, 32'hc14688c4} /* (1, 6, 15) {real, imag} */,
  {32'hc1c8ed14, 32'h4083940e} /* (1, 6, 14) {real, imag} */,
  {32'h3f9495a0, 32'h419b36b3} /* (1, 6, 13) {real, imag} */,
  {32'hc22c3a64, 32'h3f412dc0} /* (1, 6, 12) {real, imag} */,
  {32'h411eb18f, 32'hc289e550} /* (1, 6, 11) {real, imag} */,
  {32'h41a0f210, 32'hc29a249f} /* (1, 6, 10) {real, imag} */,
  {32'h42cefd75, 32'h42d18e23} /* (1, 6, 9) {real, imag} */,
  {32'h3fc764b0, 32'hc17e7220} /* (1, 6, 8) {real, imag} */,
  {32'h42b04220, 32'hc21e5eca} /* (1, 6, 7) {real, imag} */,
  {32'h403041ec, 32'h42bfce51} /* (1, 6, 6) {real, imag} */,
  {32'hc0417d60, 32'h42927f71} /* (1, 6, 5) {real, imag} */,
  {32'h427c825d, 32'hc256fd6c} /* (1, 6, 4) {real, imag} */,
  {32'h4242d701, 32'h42eee06b} /* (1, 6, 3) {real, imag} */,
  {32'hc31d2b10, 32'h42642998} /* (1, 6, 2) {real, imag} */,
  {32'hc29325b3, 32'hc220501c} /* (1, 6, 1) {real, imag} */,
  {32'h431c801d, 32'hc28cc446} /* (1, 6, 0) {real, imag} */,
  {32'hc1db0990, 32'h43cd3627} /* (1, 5, 31) {real, imag} */,
  {32'h42969914, 32'hc3901265} /* (1, 5, 30) {real, imag} */,
  {32'hc22170b8, 32'hc190c4b0} /* (1, 5, 29) {real, imag} */,
  {32'h4291afbc, 32'hc1f57c7a} /* (1, 5, 28) {real, imag} */,
  {32'h42ae1ec9, 32'hc31b092d} /* (1, 5, 27) {real, imag} */,
  {32'h42ae2ef2, 32'hc283e432} /* (1, 5, 26) {real, imag} */,
  {32'h42473b88, 32'h425e5bb1} /* (1, 5, 25) {real, imag} */,
  {32'hc2d12114, 32'h421f2cbf} /* (1, 5, 24) {real, imag} */,
  {32'h3e563080, 32'hc1e1bb00} /* (1, 5, 23) {real, imag} */,
  {32'hc1fa4c93, 32'h3e408b00} /* (1, 5, 22) {real, imag} */,
  {32'hc23ccccc, 32'hc1345c00} /* (1, 5, 21) {real, imag} */,
  {32'h407d94a0, 32'h4216a33a} /* (1, 5, 20) {real, imag} */,
  {32'h41eca6d7, 32'h41cb9320} /* (1, 5, 19) {real, imag} */,
  {32'hc292856e, 32'h4249e69a} /* (1, 5, 18) {real, imag} */,
  {32'hc1ec1130, 32'hc0af7d80} /* (1, 5, 17) {real, imag} */,
  {32'hc12086c0, 32'hc19ef260} /* (1, 5, 16) {real, imag} */,
  {32'hc2248974, 32'hc2016b10} /* (1, 5, 15) {real, imag} */,
  {32'h423c43d4, 32'hc145f258} /* (1, 5, 14) {real, imag} */,
  {32'h41bacf55, 32'hc164d740} /* (1, 5, 13) {real, imag} */,
  {32'hc207e6a6, 32'h41215029} /* (1, 5, 12) {real, imag} */,
  {32'h3f283fc0, 32'hc2435bf4} /* (1, 5, 11) {real, imag} */,
  {32'h42b05481, 32'h410500dc} /* (1, 5, 10) {real, imag} */,
  {32'h425bff98, 32'h42196fa2} /* (1, 5, 9) {real, imag} */,
  {32'hc1b978c0, 32'hc20a04f9} /* (1, 5, 8) {real, imag} */,
  {32'hc2e774a8, 32'h42d82774} /* (1, 5, 7) {real, imag} */,
  {32'h421c768c, 32'h420bf6c1} /* (1, 5, 6) {real, imag} */,
  {32'h4268e23e, 32'hc3252edb} /* (1, 5, 5) {real, imag} */,
  {32'hc3766d3a, 32'h419f2f96} /* (1, 5, 4) {real, imag} */,
  {32'h421c567c, 32'hc121ca1f} /* (1, 5, 3) {real, imag} */,
  {32'h43f16f63, 32'hc28d178c} /* (1, 5, 2) {real, imag} */,
  {32'hc3c41de1, 32'h42fb26d4} /* (1, 5, 1) {real, imag} */,
  {32'hc34884ca, 32'h43144cbc} /* (1, 5, 0) {real, imag} */,
  {32'h43af03ac, 32'h424b0d08} /* (1, 4, 31) {real, imag} */,
  {32'hc3cb132d, 32'h43f8aba3} /* (1, 4, 30) {real, imag} */,
  {32'hc24883e8, 32'h42c7edbc} /* (1, 4, 29) {real, imag} */,
  {32'h433b008e, 32'hc3873a94} /* (1, 4, 28) {real, imag} */,
  {32'hc18b7804, 32'h430ba94b} /* (1, 4, 27) {real, imag} */,
  {32'h42e63a0a, 32'h41cec228} /* (1, 4, 26) {real, imag} */,
  {32'hc21a62c9, 32'hc32f2772} /* (1, 4, 25) {real, imag} */,
  {32'hc37b328c, 32'h42fd723a} /* (1, 4, 24) {real, imag} */,
  {32'hc2908586, 32'hc248c4fc} /* (1, 4, 23) {real, imag} */,
  {32'hc1ef79a6, 32'hc061de20} /* (1, 4, 22) {real, imag} */,
  {32'h41dfbdf8, 32'hc2837e7a} /* (1, 4, 21) {real, imag} */,
  {32'h423856bf, 32'h408cce48} /* (1, 4, 20) {real, imag} */,
  {32'hc128ec28, 32'h42651cc5} /* (1, 4, 19) {real, imag} */,
  {32'hc1f773ea, 32'h4216cc85} /* (1, 4, 18) {real, imag} */,
  {32'h41f4daa8, 32'hc18e50ac} /* (1, 4, 17) {real, imag} */,
  {32'h418e5828, 32'hc2127f1e} /* (1, 4, 16) {real, imag} */,
  {32'hc0d0e3e0, 32'h4183e9ac} /* (1, 4, 15) {real, imag} */,
  {32'hc295448e, 32'h418dd086} /* (1, 4, 14) {real, imag} */,
  {32'h41c9e494, 32'hc1151cac} /* (1, 4, 13) {real, imag} */,
  {32'h42f26024, 32'hc214f70f} /* (1, 4, 12) {real, imag} */,
  {32'hc2d3f798, 32'h42028f55} /* (1, 4, 11) {real, imag} */,
  {32'hc2310815, 32'h412dfee8} /* (1, 4, 10) {real, imag} */,
  {32'h41a356b6, 32'hc20a0e34} /* (1, 4, 9) {real, imag} */,
  {32'hc3143de2, 32'h431a4b6b} /* (1, 4, 8) {real, imag} */,
  {32'hc0943368, 32'h40a8d3c0} /* (1, 4, 7) {real, imag} */,
  {32'h4296bfda, 32'hc31a8b65} /* (1, 4, 6) {real, imag} */,
  {32'hc2b1f275, 32'hc204f2d3} /* (1, 4, 5) {real, imag} */,
  {32'h438ccde8, 32'h42bb54da} /* (1, 4, 4) {real, imag} */,
  {32'h438aaee5, 32'h433f032c} /* (1, 4, 3) {real, imag} */,
  {32'hc3af3ab7, 32'h43c64541} /* (1, 4, 2) {real, imag} */,
  {32'h4252a020, 32'hc3bba6dd} /* (1, 4, 1) {real, imag} */,
  {32'h431b5d25, 32'hc317dda6} /* (1, 4, 0) {real, imag} */,
  {32'h431a3c92, 32'h43cc4450} /* (1, 3, 31) {real, imag} */,
  {32'hc3e80cb8, 32'hc3b69bec} /* (1, 3, 30) {real, imag} */,
  {32'h42a69bc6, 32'hc0ba0920} /* (1, 3, 29) {real, imag} */,
  {32'h430edb2e, 32'hc3427ad2} /* (1, 3, 28) {real, imag} */,
  {32'h42bd5bb6, 32'h42e55d56} /* (1, 3, 27) {real, imag} */,
  {32'h424e7562, 32'h42a529d5} /* (1, 3, 26) {real, imag} */,
  {32'h42b39b60, 32'hc1fb35bb} /* (1, 3, 25) {real, imag} */,
  {32'hc30e3355, 32'h427fac37} /* (1, 3, 24) {real, imag} */,
  {32'h41ed2aec, 32'hc1e426f9} /* (1, 3, 23) {real, imag} */,
  {32'h42bf6f56, 32'h42a86f87} /* (1, 3, 22) {real, imag} */,
  {32'hc25e01ad, 32'hc198a956} /* (1, 3, 21) {real, imag} */,
  {32'h411fe324, 32'h413b623f} /* (1, 3, 20) {real, imag} */,
  {32'h41569752, 32'h41700ae8} /* (1, 3, 19) {real, imag} */,
  {32'hc238809a, 32'h41aee85c} /* (1, 3, 18) {real, imag} */,
  {32'h422fe27c, 32'hc28786c8} /* (1, 3, 17) {real, imag} */,
  {32'hc217f6e5, 32'hc0124100} /* (1, 3, 16) {real, imag} */,
  {32'h41db9841, 32'hc11f6164} /* (1, 3, 15) {real, imag} */,
  {32'hc223f5a6, 32'hc117cc58} /* (1, 3, 14) {real, imag} */,
  {32'hc0abf5ac, 32'hc1dea6e4} /* (1, 3, 13) {real, imag} */,
  {32'h423508b9, 32'hc147e3d1} /* (1, 3, 12) {real, imag} */,
  {32'hc23cfe2f, 32'hc26e8187} /* (1, 3, 11) {real, imag} */,
  {32'hc1e70750, 32'hc2821767} /* (1, 3, 10) {real, imag} */,
  {32'h42e3e133, 32'h423543c8} /* (1, 3, 9) {real, imag} */,
  {32'h41ae92b6, 32'h4097a5f8} /* (1, 3, 8) {real, imag} */,
  {32'hc2735708, 32'h4227e5d6} /* (1, 3, 7) {real, imag} */,
  {32'hc34d37b4, 32'hc328f63e} /* (1, 3, 6) {real, imag} */,
  {32'h420ef24f, 32'hc2995e08} /* (1, 3, 5) {real, imag} */,
  {32'h42a992db, 32'h43775e66} /* (1, 3, 4) {real, imag} */,
  {32'hc2385564, 32'h42c25bec} /* (1, 3, 3) {real, imag} */,
  {32'hc3b8a910, 32'h4210c644} /* (1, 3, 2) {real, imag} */,
  {32'h438588fd, 32'hc34b8050} /* (1, 3, 1) {real, imag} */,
  {32'h417f378c, 32'h42c1a6eb} /* (1, 3, 0) {real, imag} */,
  {32'hc38e423c, 32'h4500541e} /* (1, 2, 31) {real, imag} */,
  {32'hc332d4f8, 32'hc4ad535e} /* (1, 2, 30) {real, imag} */,
  {32'h42962399, 32'h4149e4b4} /* (1, 2, 29) {real, imag} */,
  {32'h435ee2b1, 32'h43462bb4} /* (1, 2, 28) {real, imag} */,
  {32'hc2cc0464, 32'hc339e87d} /* (1, 2, 27) {real, imag} */,
  {32'hc2b34a95, 32'hc218d265} /* (1, 2, 26) {real, imag} */,
  {32'hc2de213c, 32'h4314395d} /* (1, 2, 25) {real, imag} */,
  {32'hc232dd96, 32'hc1b4ccfe} /* (1, 2, 24) {real, imag} */,
  {32'h42b2c984, 32'h428368db} /* (1, 2, 23) {real, imag} */,
  {32'h42774102, 32'hc29a4e1c} /* (1, 2, 22) {real, imag} */,
  {32'hc284c849, 32'hc1f5daea} /* (1, 2, 21) {real, imag} */,
  {32'hc1828b0f, 32'h4224341a} /* (1, 2, 20) {real, imag} */,
  {32'h416ff148, 32'hc298cee6} /* (1, 2, 19) {real, imag} */,
  {32'hc2ab9846, 32'hbe3bec00} /* (1, 2, 18) {real, imag} */,
  {32'h42892af6, 32'h41c209c8} /* (1, 2, 17) {real, imag} */,
  {32'hc175f6b0, 32'hc1f09bf0} /* (1, 2, 16) {real, imag} */,
  {32'hc0990a28, 32'h4153fd70} /* (1, 2, 15) {real, imag} */,
  {32'h4172ce8c, 32'hc2086b14} /* (1, 2, 14) {real, imag} */,
  {32'h40c5b580, 32'hc189ad22} /* (1, 2, 13) {real, imag} */,
  {32'h421e5de8, 32'hc226ef4a} /* (1, 2, 12) {real, imag} */,
  {32'h43318582, 32'h41307034} /* (1, 2, 11) {real, imag} */,
  {32'h41a03630, 32'h420fc229} /* (1, 2, 10) {real, imag} */,
  {32'h42cc6eb0, 32'hc0174080} /* (1, 2, 9) {real, imag} */,
  {32'hc27be38e, 32'h410059bc} /* (1, 2, 8) {real, imag} */,
  {32'hc23677b0, 32'h42f1213e} /* (1, 2, 7) {real, imag} */,
  {32'h41c73c40, 32'hc2c7d336} /* (1, 2, 6) {real, imag} */,
  {32'h43edc3cf, 32'hc3dee1c2} /* (1, 2, 5) {real, imag} */,
  {32'hc34240cb, 32'h4414b23e} /* (1, 2, 4) {real, imag} */,
  {32'hc210f13c, 32'hc1d90f62} /* (1, 2, 3) {real, imag} */,
  {32'h411c0840, 32'hc449d71d} /* (1, 2, 2) {real, imag} */,
  {32'hc1d02f30, 32'h449b2789} /* (1, 2, 1) {real, imag} */,
  {32'hc38e1240, 32'h4457ec80} /* (1, 2, 0) {real, imag} */,
  {32'hc35bce04, 32'hc4c5580c} /* (1, 1, 31) {real, imag} */,
  {32'hc30214a0, 32'h442518a0} /* (1, 1, 30) {real, imag} */,
  {32'h42f61791, 32'hc28da4a9} /* (1, 1, 29) {real, imag} */,
  {32'h436ae8c0, 32'hc3851d1b} /* (1, 1, 28) {real, imag} */,
  {32'hc308860c, 32'h440afaa0} /* (1, 1, 27) {real, imag} */,
  {32'hc2b3a163, 32'hc0039b40} /* (1, 1, 26) {real, imag} */,
  {32'hc26cf686, 32'hc363589e} /* (1, 1, 25) {real, imag} */,
  {32'h4346baa2, 32'h43468e96} /* (1, 1, 24) {real, imag} */,
  {32'h4296f753, 32'h426da69e} /* (1, 1, 23) {real, imag} */,
  {32'hc1fd246c, 32'hc2a463c6} /* (1, 1, 22) {real, imag} */,
  {32'h433427e7, 32'h4304a240} /* (1, 1, 21) {real, imag} */,
  {32'hbfa17720, 32'h41c6a150} /* (1, 1, 20) {real, imag} */,
  {32'hc18890bc, 32'hc12dc4a4} /* (1, 1, 19) {real, imag} */,
  {32'h42262744, 32'h4183d560} /* (1, 1, 18) {real, imag} */,
  {32'h410de2c0, 32'hc1040140} /* (1, 1, 17) {real, imag} */,
  {32'hc175dfc0, 32'hc12871c0} /* (1, 1, 16) {real, imag} */,
  {32'h42725e30, 32'hc0f12d80} /* (1, 1, 15) {real, imag} */,
  {32'hc29746a2, 32'hc22a8e30} /* (1, 1, 14) {real, imag} */,
  {32'h418cbd54, 32'h417487d4} /* (1, 1, 13) {real, imag} */,
  {32'hc2bbb80c, 32'h41e11e30} /* (1, 1, 12) {real, imag} */,
  {32'hc333a85d, 32'hc1bec440} /* (1, 1, 11) {real, imag} */,
  {32'hc30df27a, 32'h42698c9c} /* (1, 1, 10) {real, imag} */,
  {32'hc0dca0d0, 32'h4212975a} /* (1, 1, 9) {real, imag} */,
  {32'hc36d59fe, 32'h408f7240} /* (1, 1, 8) {real, imag} */,
  {32'hc19b0e8c, 32'hc30f2998} /* (1, 1, 7) {real, imag} */,
  {32'hc2e27e31, 32'h43852b92} /* (1, 1, 6) {real, imag} */,
  {32'hc383d7eb, 32'h43a9eb88} /* (1, 1, 5) {real, imag} */,
  {32'h43bf05ba, 32'hc34c6156} /* (1, 1, 4) {real, imag} */,
  {32'hc1ed377c, 32'h42abf697} /* (1, 1, 3) {real, imag} */,
  {32'hc469bb38, 32'h442a540c} /* (1, 1, 2) {real, imag} */,
  {32'h44aee22e, 32'hc5056a4a} /* (1, 1, 1) {real, imag} */,
  {32'h439a3b04, 32'hc4a3775c} /* (1, 1, 0) {real, imag} */,
  {32'hc4206ddd, 32'hc4810077} /* (1, 0, 31) {real, imag} */,
  {32'h43af9926, 32'h43b5e602} /* (1, 0, 30) {real, imag} */,
  {32'h4269853c, 32'hc2319cdf} /* (1, 0, 29) {real, imag} */,
  {32'h42f0c9cc, 32'h426e3936} /* (1, 0, 28) {real, imag} */,
  {32'h42842c5b, 32'h43752670} /* (1, 0, 27) {real, imag} */,
  {32'h4260fc19, 32'h415582d0} /* (1, 0, 26) {real, imag} */,
  {32'hc2ff74e2, 32'h41950bdc} /* (1, 0, 25) {real, imag} */,
  {32'h42e3a46c, 32'hc2595556} /* (1, 0, 24) {real, imag} */,
  {32'h41bca30e, 32'hc11a0180} /* (1, 0, 23) {real, imag} */,
  {32'h42baf7b0, 32'h42845a47} /* (1, 0, 22) {real, imag} */,
  {32'h40d0a398, 32'h43176578} /* (1, 0, 21) {real, imag} */,
  {32'hc1d84c51, 32'hc1a1c50a} /* (1, 0, 20) {real, imag} */,
  {32'hc159cafc, 32'hc21c8662} /* (1, 0, 19) {real, imag} */,
  {32'h42d50241, 32'h411e3c64} /* (1, 0, 18) {real, imag} */,
  {32'hc1351dac, 32'h3e803b00} /* (1, 0, 17) {real, imag} */,
  {32'hc1956bf6, 32'h42a44970} /* (1, 0, 16) {real, imag} */,
  {32'h41d87e6a, 32'h4283157d} /* (1, 0, 15) {real, imag} */,
  {32'hc1ff3ddc, 32'h420bebe7} /* (1, 0, 14) {real, imag} */,
  {32'h41176424, 32'hc1edb32f} /* (1, 0, 13) {real, imag} */,
  {32'hc2120f58, 32'hc1464024} /* (1, 0, 12) {real, imag} */,
  {32'hc1a615fa, 32'h4270ee88} /* (1, 0, 11) {real, imag} */,
  {32'h4154373c, 32'hc1b547cc} /* (1, 0, 10) {real, imag} */,
  {32'hc21f1a11, 32'h3ffde300} /* (1, 0, 9) {real, imag} */,
  {32'hc3899281, 32'h41bc91ec} /* (1, 0, 8) {real, imag} */,
  {32'hc0ac0960, 32'h41b68374} /* (1, 0, 7) {real, imag} */,
  {32'hc08f8df8, 32'hc2c0b8a2} /* (1, 0, 6) {real, imag} */,
  {32'h40be6a30, 32'h43bfd37c} /* (1, 0, 5) {real, imag} */,
  {32'hc2e06a08, 32'h430d5c72} /* (1, 0, 4) {real, imag} */,
  {32'h423a38f4, 32'h4286bc40} /* (1, 0, 3) {real, imag} */,
  {32'hc3d50e90, 32'h42c58df6} /* (1, 0, 2) {real, imag} */,
  {32'h445bc1f9, 32'hc45675ef} /* (1, 0, 1) {real, imag} */,
  {32'h429ac1e8, 32'hc45743c8} /* (1, 0, 0) {real, imag} */,
  {32'hbf89dc18, 32'h4249447b} /* (0, 31, 31) {real, imag} */,
  {32'hc2f83c21, 32'h4287eed2} /* (0, 31, 30) {real, imag} */,
  {32'hc135e7f4, 32'h424941b2} /* (0, 31, 29) {real, imag} */,
  {32'hc1f962b6, 32'h43243ac4} /* (0, 31, 28) {real, imag} */,
  {32'hc2612f44, 32'hc323705a} /* (0, 31, 27) {real, imag} */,
  {32'hc2bed0db, 32'h43130e9d} /* (0, 31, 26) {real, imag} */,
  {32'h40fc13f0, 32'h4165e264} /* (0, 31, 25) {real, imag} */,
  {32'h429a8577, 32'h3e72e900} /* (0, 31, 24) {real, imag} */,
  {32'hc20f9360, 32'hc285def1} /* (0, 31, 23) {real, imag} */,
  {32'hc2eb4f0f, 32'h424bbb5f} /* (0, 31, 22) {real, imag} */,
  {32'hc1cbe943, 32'hc2963721} /* (0, 31, 21) {real, imag} */,
  {32'h42a67dce, 32'h42916894} /* (0, 31, 20) {real, imag} */,
  {32'h426c0e05, 32'h422107a0} /* (0, 31, 19) {real, imag} */,
  {32'hc1c7a8c4, 32'hc0920a54} /* (0, 31, 18) {real, imag} */,
  {32'h40742c50, 32'hc2847f10} /* (0, 31, 17) {real, imag} */,
  {32'hc13e7b18, 32'h4222b66c} /* (0, 31, 16) {real, imag} */,
  {32'h41fb6fa6, 32'hc1b786d2} /* (0, 31, 15) {real, imag} */,
  {32'hc0cf38b0, 32'hc24dc3fe} /* (0, 31, 14) {real, imag} */,
  {32'h420625ff, 32'h425e60de} /* (0, 31, 13) {real, imag} */,
  {32'h4204aac7, 32'hc2ab9f22} /* (0, 31, 12) {real, imag} */,
  {32'hc13730ee, 32'hc284aed5} /* (0, 31, 11) {real, imag} */,
  {32'h42d969bb, 32'hbe868f80} /* (0, 31, 10) {real, imag} */,
  {32'hbeb9f1c0, 32'h42ce36a3} /* (0, 31, 9) {real, imag} */,
  {32'hc22f5f64, 32'h42b11a9a} /* (0, 31, 8) {real, imag} */,
  {32'hc2e736e3, 32'hc05aa32e} /* (0, 31, 7) {real, imag} */,
  {32'h431d356a, 32'h42f769aa} /* (0, 31, 6) {real, imag} */,
  {32'h4354cbc1, 32'hc1c693dc} /* (0, 31, 5) {real, imag} */,
  {32'hc2f63434, 32'h4258ede2} /* (0, 31, 4) {real, imag} */,
  {32'h429d7f74, 32'h42786760} /* (0, 31, 3) {real, imag} */,
  {32'h4160f548, 32'hc2ec5784} /* (0, 31, 2) {real, imag} */,
  {32'h41d10b9a, 32'h41e5df66} /* (0, 31, 1) {real, imag} */,
  {32'h42120475, 32'h419c254c} /* (0, 31, 0) {real, imag} */,
  {32'h4083fa26, 32'hc2ec9816} /* (0, 30, 31) {real, imag} */,
  {32'h420003e0, 32'hc2790026} /* (0, 30, 30) {real, imag} */,
  {32'hc19d89f0, 32'h42874e6a} /* (0, 30, 29) {real, imag} */,
  {32'h42f7a94d, 32'h43501255} /* (0, 30, 28) {real, imag} */,
  {32'hc331f380, 32'h42ea86dc} /* (0, 30, 27) {real, imag} */,
  {32'h42c135e2, 32'hc34af9d2} /* (0, 30, 26) {real, imag} */,
  {32'h42845e4e, 32'h42e01453} /* (0, 30, 25) {real, imag} */,
  {32'hc22b40ad, 32'h428d5710} /* (0, 30, 24) {real, imag} */,
  {32'h429e980a, 32'hc3080882} /* (0, 30, 23) {real, imag} */,
  {32'hbf522380, 32'hc271724b} /* (0, 30, 22) {real, imag} */,
  {32'hc140e48c, 32'hc0b9d1e6} /* (0, 30, 21) {real, imag} */,
  {32'h416d1c3c, 32'hc1be803b} /* (0, 30, 20) {real, imag} */,
  {32'hc22a5c74, 32'h4174d250} /* (0, 30, 19) {real, imag} */,
  {32'h41f39ad6, 32'h41d49f1e} /* (0, 30, 18) {real, imag} */,
  {32'h40f18db6, 32'h412c5a2e} /* (0, 30, 17) {real, imag} */,
  {32'h41124280, 32'h404c7c90} /* (0, 30, 16) {real, imag} */,
  {32'h417977a7, 32'h423b4544} /* (0, 30, 15) {real, imag} */,
  {32'h40a94a70, 32'h4229795d} /* (0, 30, 14) {real, imag} */,
  {32'hc2aebab8, 32'hc20bc80a} /* (0, 30, 13) {real, imag} */,
  {32'h42662f09, 32'h422086a4} /* (0, 30, 12) {real, imag} */,
  {32'h4218c4f9, 32'hc1b0d462} /* (0, 30, 11) {real, imag} */,
  {32'hc22509f0, 32'h41cf0196} /* (0, 30, 10) {real, imag} */,
  {32'hc2c8cbba, 32'hc15f8e88} /* (0, 30, 9) {real, imag} */,
  {32'h426e143b, 32'hc31ea28e} /* (0, 30, 8) {real, imag} */,
  {32'h4293f668, 32'hc08bc050} /* (0, 30, 7) {real, imag} */,
  {32'h423f2e7b, 32'hc2c053e0} /* (0, 30, 6) {real, imag} */,
  {32'h420b8ac6, 32'h429b65cc} /* (0, 30, 5) {real, imag} */,
  {32'h423905ee, 32'hc2a15a3e} /* (0, 30, 4) {real, imag} */,
  {32'h431eb629, 32'hc2e53c96} /* (0, 30, 3) {real, imag} */,
  {32'h42b45046, 32'h42d8886d} /* (0, 30, 2) {real, imag} */,
  {32'hc1b81d1c, 32'h3f4de400} /* (0, 30, 1) {real, imag} */,
  {32'hc25e719e, 32'h41a0901c} /* (0, 30, 0) {real, imag} */,
  {32'h411a31d2, 32'hc2c207b8} /* (0, 29, 31) {real, imag} */,
  {32'h41e33a80, 32'hc3547c98} /* (0, 29, 30) {real, imag} */,
  {32'h410e71b0, 32'h42af889e} /* (0, 29, 29) {real, imag} */,
  {32'h42945764, 32'hc30f5652} /* (0, 29, 28) {real, imag} */,
  {32'hc32ed360, 32'hc3132f7f} /* (0, 29, 27) {real, imag} */,
  {32'hc2e1124f, 32'h4181d03a} /* (0, 29, 26) {real, imag} */,
  {32'hc1925178, 32'h42d0ff18} /* (0, 29, 25) {real, imag} */,
  {32'hc2e24200, 32'hc2801ea5} /* (0, 29, 24) {real, imag} */,
  {32'hc0f0fff8, 32'h42656a95} /* (0, 29, 23) {real, imag} */,
  {32'hc05f6b3c, 32'hc2384564} /* (0, 29, 22) {real, imag} */,
  {32'h40b703c0, 32'h427b4e1e} /* (0, 29, 21) {real, imag} */,
  {32'h42b8efa8, 32'h42cfee72} /* (0, 29, 20) {real, imag} */,
  {32'hc1193c5c, 32'h419078c8} /* (0, 29, 19) {real, imag} */,
  {32'h42362b08, 32'hc24c8475} /* (0, 29, 18) {real, imag} */,
  {32'h4125d43e, 32'h41109c38} /* (0, 29, 17) {real, imag} */,
  {32'h40ff7390, 32'h4213115a} /* (0, 29, 16) {real, imag} */,
  {32'h423b18f4, 32'h408ab520} /* (0, 29, 15) {real, imag} */,
  {32'hc04c9600, 32'h425f8743} /* (0, 29, 14) {real, imag} */,
  {32'h41d577c0, 32'hc1ea65ee} /* (0, 29, 13) {real, imag} */,
  {32'hbf8531e0, 32'hc1f6216a} /* (0, 29, 12) {real, imag} */,
  {32'hc29d864c, 32'h4166c4c8} /* (0, 29, 11) {real, imag} */,
  {32'hc12a4f29, 32'hc1290fd8} /* (0, 29, 10) {real, imag} */,
  {32'hc2596b69, 32'h42d52a4a} /* (0, 29, 9) {real, imag} */,
  {32'h42136c9c, 32'h4236056e} /* (0, 29, 8) {real, imag} */,
  {32'hc343ba7b, 32'hc2fc6ce0} /* (0, 29, 7) {real, imag} */,
  {32'hc2f9699d, 32'hc26c6183} /* (0, 29, 6) {real, imag} */,
  {32'h41fd6164, 32'h4309dca9} /* (0, 29, 5) {real, imag} */,
  {32'h4134f49c, 32'hc2534a88} /* (0, 29, 4) {real, imag} */,
  {32'hc2ab15bc, 32'hc2aaeb3e} /* (0, 29, 3) {real, imag} */,
  {32'h42399068, 32'h41af83d0} /* (0, 29, 2) {real, imag} */,
  {32'h40a07534, 32'h42f26d7c} /* (0, 29, 1) {real, imag} */,
  {32'h4332e222, 32'hc27a93da} /* (0, 29, 0) {real, imag} */,
  {32'h4202d43f, 32'hc29c3656} /* (0, 28, 31) {real, imag} */,
  {32'h4364c487, 32'h40c0be08} /* (0, 28, 30) {real, imag} */,
  {32'hc2b2e114, 32'hc293d46c} /* (0, 28, 29) {real, imag} */,
  {32'h435ff93c, 32'h423e760c} /* (0, 28, 28) {real, imag} */,
  {32'h42636f7c, 32'h4321566c} /* (0, 28, 27) {real, imag} */,
  {32'hc31544fc, 32'hc3469a9e} /* (0, 28, 26) {real, imag} */,
  {32'hc3200156, 32'h41ce27d4} /* (0, 28, 25) {real, imag} */,
  {32'h41fa456e, 32'h41cae9d0} /* (0, 28, 24) {real, imag} */,
  {32'h42beff6b, 32'h424079fb} /* (0, 28, 23) {real, imag} */,
  {32'h4235e490, 32'hc0d53ba8} /* (0, 28, 22) {real, imag} */,
  {32'h42a98e4c, 32'hc2994f57} /* (0, 28, 21) {real, imag} */,
  {32'hc29183c1, 32'h4214a6fe} /* (0, 28, 20) {real, imag} */,
  {32'h427174df, 32'hc2315f4f} /* (0, 28, 19) {real, imag} */,
  {32'hbf5c2760, 32'hc15127fc} /* (0, 28, 18) {real, imag} */,
  {32'hc22d30d6, 32'h41a56855} /* (0, 28, 17) {real, imag} */,
  {32'hc2188e80, 32'hc1cc5be2} /* (0, 28, 16) {real, imag} */,
  {32'h41bc1ed4, 32'hc1d0043b} /* (0, 28, 15) {real, imag} */,
  {32'hc1640326, 32'h4209e4df} /* (0, 28, 14) {real, imag} */,
  {32'hc219bddf, 32'h41c9ee2a} /* (0, 28, 13) {real, imag} */,
  {32'h42a547c9, 32'hc2239546} /* (0, 28, 12) {real, imag} */,
  {32'h41907e14, 32'hc24cc938} /* (0, 28, 11) {real, imag} */,
  {32'hc1b72450, 32'hc13dc914} /* (0, 28, 10) {real, imag} */,
  {32'hc24e8422, 32'h42b8a8e0} /* (0, 28, 9) {real, imag} */,
  {32'h431d3349, 32'h43343331} /* (0, 28, 8) {real, imag} */,
  {32'h422a10ce, 32'hc32b9020} /* (0, 28, 7) {real, imag} */,
  {32'hc3272bdc, 32'h42b00534} /* (0, 28, 6) {real, imag} */,
  {32'h41999cd4, 32'h4327b0e0} /* (0, 28, 5) {real, imag} */,
  {32'hc237be26, 32'h41958871} /* (0, 28, 4) {real, imag} */,
  {32'hc2f34898, 32'h42671ff1} /* (0, 28, 3) {real, imag} */,
  {32'hc34d33e9, 32'hc2f2aebe} /* (0, 28, 2) {real, imag} */,
  {32'hc161885f, 32'h43101885} /* (0, 28, 1) {real, imag} */,
  {32'hc3068865, 32'h427e4191} /* (0, 28, 0) {real, imag} */,
  {32'h415de393, 32'hc33ea688} /* (0, 27, 31) {real, imag} */,
  {32'h42db17fc, 32'h4232db6b} /* (0, 27, 30) {real, imag} */,
  {32'hc24d56ac, 32'h42ae1ab8} /* (0, 27, 29) {real, imag} */,
  {32'hc1bb4ada, 32'hc280016e} /* (0, 27, 28) {real, imag} */,
  {32'h423d3d48, 32'hc284a6f1} /* (0, 27, 27) {real, imag} */,
  {32'hc1a4700e, 32'hc2004834} /* (0, 27, 26) {real, imag} */,
  {32'h42ab0509, 32'hc25474db} /* (0, 27, 25) {real, imag} */,
  {32'h42c53a54, 32'hc299b8a8} /* (0, 27, 24) {real, imag} */,
  {32'h41f6aa0e, 32'h420c4c99} /* (0, 27, 23) {real, imag} */,
  {32'h4084f518, 32'hc2326166} /* (0, 27, 22) {real, imag} */,
  {32'hc1e9c264, 32'h42deb5bd} /* (0, 27, 21) {real, imag} */,
  {32'h41e9d158, 32'h42815bb1} /* (0, 27, 20) {real, imag} */,
  {32'h421d34d5, 32'hc1eb0d34} /* (0, 27, 19) {real, imag} */,
  {32'hc1afd92a, 32'hc21f36f5} /* (0, 27, 18) {real, imag} */,
  {32'hc1d93c3b, 32'hc11a757c} /* (0, 27, 17) {real, imag} */,
  {32'hc1f21e2e, 32'h409147c0} /* (0, 27, 16) {real, imag} */,
  {32'hc1be9f55, 32'h420815e5} /* (0, 27, 15) {real, imag} */,
  {32'hc1c0a70a, 32'hc1c753de} /* (0, 27, 14) {real, imag} */,
  {32'hc0e38038, 32'hc1ea3f24} /* (0, 27, 13) {real, imag} */,
  {32'h417fe458, 32'h429b64bb} /* (0, 27, 12) {real, imag} */,
  {32'h401cd714, 32'h4291fb77} /* (0, 27, 11) {real, imag} */,
  {32'hc2b5c056, 32'h40c54540} /* (0, 27, 10) {real, imag} */,
  {32'hc15b3c90, 32'hc2839f56} /* (0, 27, 9) {real, imag} */,
  {32'hc2bab9ce, 32'h4245e0b3} /* (0, 27, 8) {real, imag} */,
  {32'hc2144bce, 32'hc2ab2b3e} /* (0, 27, 7) {real, imag} */,
  {32'h41b5e852, 32'hc291f5af} /* (0, 27, 6) {real, imag} */,
  {32'hc1a86fe8, 32'hc2e6b42f} /* (0, 27, 5) {real, imag} */,
  {32'hc2d5b18e, 32'hc2bf4066} /* (0, 27, 4) {real, imag} */,
  {32'h426f3f58, 32'hc23b200d} /* (0, 27, 3) {real, imag} */,
  {32'hc342cc6a, 32'h4304d3d2} /* (0, 27, 2) {real, imag} */,
  {32'h413f646f, 32'hc2920b1b} /* (0, 27, 1) {real, imag} */,
  {32'hc2d347a8, 32'hc2ef783e} /* (0, 27, 0) {real, imag} */,
  {32'hc2812561, 32'hc1c48754} /* (0, 26, 31) {real, imag} */,
  {32'h40f5dbbc, 32'h428c06c4} /* (0, 26, 30) {real, imag} */,
  {32'h423ebfaf, 32'h4213d2be} /* (0, 26, 29) {real, imag} */,
  {32'h428949e1, 32'hc0df73a0} /* (0, 26, 28) {real, imag} */,
  {32'hc0ed82a6, 32'hbfc8ce90} /* (0, 26, 27) {real, imag} */,
  {32'hc2835d40, 32'h425e628c} /* (0, 26, 26) {real, imag} */,
  {32'h42d5ffbc, 32'hc318bfc5} /* (0, 26, 25) {real, imag} */,
  {32'hc23e2ce3, 32'h42b80c98} /* (0, 26, 24) {real, imag} */,
  {32'hc18113fa, 32'hc294ba74} /* (0, 26, 23) {real, imag} */,
  {32'hc236859e, 32'hc1b1d28e} /* (0, 26, 22) {real, imag} */,
  {32'hc04da890, 32'hc13fe662} /* (0, 26, 21) {real, imag} */,
  {32'h411fa239, 32'hc120a36e} /* (0, 26, 20) {real, imag} */,
  {32'h423f38d9, 32'h41ef8def} /* (0, 26, 19) {real, imag} */,
  {32'hc0c11024, 32'hc1519af8} /* (0, 26, 18) {real, imag} */,
  {32'h403f26ac, 32'h40649930} /* (0, 26, 17) {real, imag} */,
  {32'hc14dde48, 32'h41abedf3} /* (0, 26, 16) {real, imag} */,
  {32'h3efd5560, 32'h42631f07} /* (0, 26, 15) {real, imag} */,
  {32'h424059f2, 32'hc1affab0} /* (0, 26, 14) {real, imag} */,
  {32'hc0d06248, 32'h4213e77c} /* (0, 26, 13) {real, imag} */,
  {32'hc0a2296a, 32'h414b46ae} /* (0, 26, 12) {real, imag} */,
  {32'hc236d1c9, 32'h41a2a16f} /* (0, 26, 11) {real, imag} */,
  {32'h429cd514, 32'h400df510} /* (0, 26, 10) {real, imag} */,
  {32'h424c3c77, 32'hc2724dd8} /* (0, 26, 9) {real, imag} */,
  {32'hc287ad30, 32'hc0e9bb38} /* (0, 26, 8) {real, imag} */,
  {32'hc207a6bb, 32'hc1324f30} /* (0, 26, 7) {real, imag} */,
  {32'h42449dce, 32'hc2bd39c2} /* (0, 26, 6) {real, imag} */,
  {32'hc1a883de, 32'h4188efd7} /* (0, 26, 5) {real, imag} */,
  {32'h41e194cc, 32'h42e7abca} /* (0, 26, 4) {real, imag} */,
  {32'h4181c17e, 32'h42fda3ab} /* (0, 26, 3) {real, imag} */,
  {32'hc28b6ebd, 32'h41d4e67a} /* (0, 26, 2) {real, imag} */,
  {32'h424dd6c8, 32'hc2e3b94f} /* (0, 26, 1) {real, imag} */,
  {32'h429d7e87, 32'h401d38d0} /* (0, 26, 0) {real, imag} */,
  {32'h42207900, 32'hc2260e94} /* (0, 25, 31) {real, imag} */,
  {32'hc0b5b20e, 32'h41cc8308} /* (0, 25, 30) {real, imag} */,
  {32'hc110cac0, 32'hc3236b70} /* (0, 25, 29) {real, imag} */,
  {32'h42c98ae0, 32'hc1300228} /* (0, 25, 28) {real, imag} */,
  {32'h42bc516f, 32'hc2532e8c} /* (0, 25, 27) {real, imag} */,
  {32'h43060aa0, 32'h4290f07d} /* (0, 25, 26) {real, imag} */,
  {32'hc2891048, 32'h421a2a74} /* (0, 25, 25) {real, imag} */,
  {32'hc050f750, 32'h42add5fb} /* (0, 25, 24) {real, imag} */,
  {32'h428e3b6a, 32'hc2938395} /* (0, 25, 23) {real, imag} */,
  {32'hc1cd4faf, 32'hc2a080a4} /* (0, 25, 22) {real, imag} */,
  {32'hc1668cd4, 32'hc1a58c8e} /* (0, 25, 21) {real, imag} */,
  {32'hc22bc450, 32'h40dda930} /* (0, 25, 20) {real, imag} */,
  {32'hc1d41d5d, 32'hc1cab616} /* (0, 25, 19) {real, imag} */,
  {32'hc228b0ae, 32'hbff8e110} /* (0, 25, 18) {real, imag} */,
  {32'hc19b0db8, 32'hc1bfa57c} /* (0, 25, 17) {real, imag} */,
  {32'h418ce69a, 32'hc114df30} /* (0, 25, 16) {real, imag} */,
  {32'h40e2a432, 32'h40a66c0e} /* (0, 25, 15) {real, imag} */,
  {32'hc0e6a14c, 32'h419ccebd} /* (0, 25, 14) {real, imag} */,
  {32'h3efa92c0, 32'hc25e1527} /* (0, 25, 13) {real, imag} */,
  {32'h41f65a88, 32'h42167622} /* (0, 25, 12) {real, imag} */,
  {32'h4255044f, 32'hc21fd681} /* (0, 25, 11) {real, imag} */,
  {32'hc01050b8, 32'hc2913f02} /* (0, 25, 10) {real, imag} */,
  {32'hc28f8a28, 32'hc3076c44} /* (0, 25, 9) {real, imag} */,
  {32'hc246af30, 32'h42a09c09} /* (0, 25, 8) {real, imag} */,
  {32'hc118599e, 32'hc1d92498} /* (0, 25, 7) {real, imag} */,
  {32'hc287b750, 32'hc197b21c} /* (0, 25, 6) {real, imag} */,
  {32'hc2b1b5e7, 32'hc32140c7} /* (0, 25, 5) {real, imag} */,
  {32'hc3350df4, 32'hc0debcf1} /* (0, 25, 4) {real, imag} */,
  {32'hc2da88d6, 32'hc0a85870} /* (0, 25, 3) {real, imag} */,
  {32'h412aa03d, 32'h430a1c47} /* (0, 25, 2) {real, imag} */,
  {32'hc2bc0cc0, 32'hc1000840} /* (0, 25, 1) {real, imag} */,
  {32'h40cd34ee, 32'h42bc2ce6} /* (0, 25, 0) {real, imag} */,
  {32'hc2b26391, 32'h4151b302} /* (0, 24, 31) {real, imag} */,
  {32'hc16b8a4e, 32'h424148e6} /* (0, 24, 30) {real, imag} */,
  {32'hc27020e9, 32'hc301ad05} /* (0, 24, 29) {real, imag} */,
  {32'hc2c6e4dc, 32'h42096526} /* (0, 24, 28) {real, imag} */,
  {32'hc10663a0, 32'h425ed42d} /* (0, 24, 27) {real, imag} */,
  {32'hc01c6c20, 32'h42a4a017} /* (0, 24, 26) {real, imag} */,
  {32'hc21ec3bb, 32'hc1a488c4} /* (0, 24, 25) {real, imag} */,
  {32'hc29589c9, 32'h427fb001} /* (0, 24, 24) {real, imag} */,
  {32'hc26c0677, 32'hc2ae6d10} /* (0, 24, 23) {real, imag} */,
  {32'h41b43cbd, 32'hc2c45d68} /* (0, 24, 22) {real, imag} */,
  {32'h42f83d82, 32'h41a26c06} /* (0, 24, 21) {real, imag} */,
  {32'h40cb1310, 32'hc1a0e156} /* (0, 24, 20) {real, imag} */,
  {32'hc203a6c3, 32'h42224261} /* (0, 24, 19) {real, imag} */,
  {32'h41472f46, 32'h3f9b6e90} /* (0, 24, 18) {real, imag} */,
  {32'h409abea2, 32'hc225d996} /* (0, 24, 17) {real, imag} */,
  {32'h41666edc, 32'hc1941fef} /* (0, 24, 16) {real, imag} */,
  {32'hc12339e1, 32'hc11d4172} /* (0, 24, 15) {real, imag} */,
  {32'h4205db46, 32'hc1f653db} /* (0, 24, 14) {real, imag} */,
  {32'hc18a05ea, 32'h4175bf54} /* (0, 24, 13) {real, imag} */,
  {32'hc13f0920, 32'hc1d54d6a} /* (0, 24, 12) {real, imag} */,
  {32'h419e05b0, 32'hc28052a2} /* (0, 24, 11) {real, imag} */,
  {32'hc2854029, 32'h4223c59c} /* (0, 24, 10) {real, imag} */,
  {32'h423a60ff, 32'h422e6279} /* (0, 24, 9) {real, imag} */,
  {32'hc24f5afe, 32'h4282ac6b} /* (0, 24, 8) {real, imag} */,
  {32'h4315ef87, 32'h42c6c38e} /* (0, 24, 7) {real, imag} */,
  {32'h42602a2b, 32'hc1e8c361} /* (0, 24, 6) {real, imag} */,
  {32'hc29618d2, 32'h42845eb2} /* (0, 24, 5) {real, imag} */,
  {32'h42a3f06c, 32'hc30a76e0} /* (0, 24, 4) {real, imag} */,
  {32'h4245b5e1, 32'h430af2b7} /* (0, 24, 3) {real, imag} */,
  {32'hc1cfa075, 32'hc2b0558d} /* (0, 24, 2) {real, imag} */,
  {32'hc2afb2c5, 32'h41a8dd53} /* (0, 24, 1) {real, imag} */,
  {32'hc234d54f, 32'hc120a06a} /* (0, 24, 0) {real, imag} */,
  {32'hc267e1cc, 32'h431c3167} /* (0, 23, 31) {real, imag} */,
  {32'hc26ae34e, 32'h43108018} /* (0, 23, 30) {real, imag} */,
  {32'hc1a7aebc, 32'h421357a3} /* (0, 23, 29) {real, imag} */,
  {32'hc23483f2, 32'h419748df} /* (0, 23, 28) {real, imag} */,
  {32'hc2155132, 32'hc2ddc24b} /* (0, 23, 27) {real, imag} */,
  {32'hc1fd3527, 32'h4101a268} /* (0, 23, 26) {real, imag} */,
  {32'h41989fcc, 32'hc28db7ee} /* (0, 23, 25) {real, imag} */,
  {32'hc103e4bd, 32'h4135fd66} /* (0, 23, 24) {real, imag} */,
  {32'h424ebbda, 32'hc2945372} /* (0, 23, 23) {real, imag} */,
  {32'hc1a9f208, 32'h41f22ccc} /* (0, 23, 22) {real, imag} */,
  {32'hc25b9f74, 32'hc1efee26} /* (0, 23, 21) {real, imag} */,
  {32'hc10e07f6, 32'h41e08a6c} /* (0, 23, 20) {real, imag} */,
  {32'hc1a4926a, 32'hc1281056} /* (0, 23, 19) {real, imag} */,
  {32'hc14bccd2, 32'hc14ed8de} /* (0, 23, 18) {real, imag} */,
  {32'hc02cdc40, 32'h41250533} /* (0, 23, 17) {real, imag} */,
  {32'h4212c282, 32'hc1e08dcd} /* (0, 23, 16) {real, imag} */,
  {32'hc1b19550, 32'hc1b87536} /* (0, 23, 15) {real, imag} */,
  {32'h4181bfff, 32'h41501372} /* (0, 23, 14) {real, imag} */,
  {32'h41423097, 32'hc19c434d} /* (0, 23, 13) {real, imag} */,
  {32'h425cab36, 32'h3ee57c60} /* (0, 23, 12) {real, imag} */,
  {32'hc20561c4, 32'h411c3264} /* (0, 23, 11) {real, imag} */,
  {32'hc1f5ae3a, 32'h414f5bd1} /* (0, 23, 10) {real, imag} */,
  {32'hc257cb94, 32'hc26a5d34} /* (0, 23, 9) {real, imag} */,
  {32'hc0a5a76e, 32'h40a218d4} /* (0, 23, 8) {real, imag} */,
  {32'hc13f4ad0, 32'hc146a634} /* (0, 23, 7) {real, imag} */,
  {32'h411327ca, 32'hc16358be} /* (0, 23, 6) {real, imag} */,
  {32'h41838a25, 32'hc191afa4} /* (0, 23, 5) {real, imag} */,
  {32'hc227ddee, 32'hc1222d28} /* (0, 23, 4) {real, imag} */,
  {32'h4253e906, 32'h426a8521} /* (0, 23, 3) {real, imag} */,
  {32'h4321d7bc, 32'hc2bcdea7} /* (0, 23, 2) {real, imag} */,
  {32'hc3062800, 32'hc368271b} /* (0, 23, 1) {real, imag} */,
  {32'hc29957b5, 32'h41b97287} /* (0, 23, 0) {real, imag} */,
  {32'hc2263727, 32'h42cb6011} /* (0, 22, 31) {real, imag} */,
  {32'h420dcfdc, 32'hc18e697c} /* (0, 22, 30) {real, imag} */,
  {32'h41ffd6dc, 32'hc1706b46} /* (0, 22, 29) {real, imag} */,
  {32'h41fc8b07, 32'h4261e242} /* (0, 22, 28) {real, imag} */,
  {32'hc1fd4b14, 32'h41e06bd3} /* (0, 22, 27) {real, imag} */,
  {32'hc1b83a82, 32'hbfa79740} /* (0, 22, 26) {real, imag} */,
  {32'h42ef60db, 32'hc15a4c59} /* (0, 22, 25) {real, imag} */,
  {32'hc13f12c4, 32'hc2300091} /* (0, 22, 24) {real, imag} */,
  {32'h4228747b, 32'h41ce5042} /* (0, 22, 23) {real, imag} */,
  {32'hc20d91b7, 32'hc254bfba} /* (0, 22, 22) {real, imag} */,
  {32'h4224a790, 32'hc0e3fe98} /* (0, 22, 21) {real, imag} */,
  {32'hc2983931, 32'hc0d065fc} /* (0, 22, 20) {real, imag} */,
  {32'h4194d257, 32'h42095596} /* (0, 22, 19) {real, imag} */,
  {32'h414d812c, 32'h415b3501} /* (0, 22, 18) {real, imag} */,
  {32'hc1883e5e, 32'hc138523c} /* (0, 22, 17) {real, imag} */,
  {32'hc181505c, 32'h4022dde4} /* (0, 22, 16) {real, imag} */,
  {32'h417975b5, 32'h4008f0c0} /* (0, 22, 15) {real, imag} */,
  {32'hc13b27f8, 32'hc1168345} /* (0, 22, 14) {real, imag} */,
  {32'h420ff7d0, 32'h408a8e5c} /* (0, 22, 13) {real, imag} */,
  {32'h411ce918, 32'hc0b8cc84} /* (0, 22, 12) {real, imag} */,
  {32'hbf631560, 32'h429678d0} /* (0, 22, 11) {real, imag} */,
  {32'h40d0731e, 32'hbe90e6c0} /* (0, 22, 10) {real, imag} */,
  {32'h419e739a, 32'hc18445a4} /* (0, 22, 9) {real, imag} */,
  {32'hc1e062e2, 32'h41a0dc52} /* (0, 22, 8) {real, imag} */,
  {32'hc26588da, 32'h41c427ba} /* (0, 22, 7) {real, imag} */,
  {32'h41c30f34, 32'h40453c40} /* (0, 22, 6) {real, imag} */,
  {32'h4250ea82, 32'h41b41717} /* (0, 22, 5) {real, imag} */,
  {32'hc2b4a30e, 32'h42dad9a3} /* (0, 22, 4) {real, imag} */,
  {32'hc32e7cac, 32'h4218230c} /* (0, 22, 3) {real, imag} */,
  {32'h4201bd1c, 32'hc1433b13} /* (0, 22, 2) {real, imag} */,
  {32'h41dba34a, 32'hc1189f78} /* (0, 22, 1) {real, imag} */,
  {32'hc1d8c0f8, 32'hc1a493c0} /* (0, 22, 0) {real, imag} */,
  {32'hc1703e0c, 32'h415765aa} /* (0, 21, 31) {real, imag} */,
  {32'hc22de9c8, 32'hc245aecd} /* (0, 21, 30) {real, imag} */,
  {32'h42058806, 32'h41f54182} /* (0, 21, 29) {real, imag} */,
  {32'hc23d9f70, 32'h421611c5} /* (0, 21, 28) {real, imag} */,
  {32'hc255225f, 32'h3fa24548} /* (0, 21, 27) {real, imag} */,
  {32'hc221594c, 32'hc245f477} /* (0, 21, 26) {real, imag} */,
  {32'hc21202b0, 32'hc21f0160} /* (0, 21, 25) {real, imag} */,
  {32'h412824f6, 32'hbfd17230} /* (0, 21, 24) {real, imag} */,
  {32'h41d1d6a2, 32'h41c334ef} /* (0, 21, 23) {real, imag} */,
  {32'hc2257789, 32'hbedf2f58} /* (0, 21, 22) {real, imag} */,
  {32'h4191f004, 32'h410296d6} /* (0, 21, 21) {real, imag} */,
  {32'hc122cb65, 32'h417403f0} /* (0, 21, 20) {real, imag} */,
  {32'hc1d61a1c, 32'hc0435fe8} /* (0, 21, 19) {real, imag} */,
  {32'h411f0ba4, 32'h41f681ef} /* (0, 21, 18) {real, imag} */,
  {32'hbf965940, 32'hc1a4afed} /* (0, 21, 17) {real, imag} */,
  {32'hc1715f56, 32'hc1c16fc6} /* (0, 21, 16) {real, imag} */,
  {32'hbf38dac0, 32'hc150c562} /* (0, 21, 15) {real, imag} */,
  {32'hc0f35d60, 32'h3fd13190} /* (0, 21, 14) {real, imag} */,
  {32'h401cdbb4, 32'h419ab163} /* (0, 21, 13) {real, imag} */,
  {32'h406f8264, 32'hc12fae48} /* (0, 21, 12) {real, imag} */,
  {32'h411fee58, 32'hc24ce3d4} /* (0, 21, 11) {real, imag} */,
  {32'hc1d1d48e, 32'hc03f685b} /* (0, 21, 10) {real, imag} */,
  {32'h41394567, 32'h42806aec} /* (0, 21, 9) {real, imag} */,
  {32'h42125dc4, 32'h418972de} /* (0, 21, 8) {real, imag} */,
  {32'hbf4f4da0, 32'h42367224} /* (0, 21, 7) {real, imag} */,
  {32'h4180c565, 32'h42298559} /* (0, 21, 6) {real, imag} */,
  {32'h42082225, 32'hc02b0f0c} /* (0, 21, 5) {real, imag} */,
  {32'hc1b89c60, 32'hc234f9e7} /* (0, 21, 4) {real, imag} */,
  {32'h40cb56bc, 32'hc1bd2de2} /* (0, 21, 3) {real, imag} */,
  {32'h41be8f2f, 32'h4222955b} /* (0, 21, 2) {real, imag} */,
  {32'h420bb78f, 32'h40b9f904} /* (0, 21, 1) {real, imag} */,
  {32'h40a04798, 32'h4266990d} /* (0, 21, 0) {real, imag} */,
  {32'h429dea4d, 32'hc2655b5d} /* (0, 20, 31) {real, imag} */,
  {32'hc177025a, 32'hc2378cdc} /* (0, 20, 30) {real, imag} */,
  {32'hc29a42f6, 32'h42308486} /* (0, 20, 29) {real, imag} */,
  {32'h41334599, 32'h41eaad07} /* (0, 20, 28) {real, imag} */,
  {32'h4103e0ff, 32'h41be7b77} /* (0, 20, 27) {real, imag} */,
  {32'h404815a0, 32'h4149d800} /* (0, 20, 26) {real, imag} */,
  {32'hbe881540, 32'h419ec235} /* (0, 20, 25) {real, imag} */,
  {32'h41b99174, 32'h3da26100} /* (0, 20, 24) {real, imag} */,
  {32'hc010c938, 32'h41cf7d2c} /* (0, 20, 23) {real, imag} */,
  {32'hc0ab47d0, 32'hc19ebfe4} /* (0, 20, 22) {real, imag} */,
  {32'hc088fdf0, 32'hbfb7c890} /* (0, 20, 21) {real, imag} */,
  {32'h4182f946, 32'hc1338c37} /* (0, 20, 20) {real, imag} */,
  {32'hc1cd3914, 32'h40eedc82} /* (0, 20, 19) {real, imag} */,
  {32'hc0ec7ed6, 32'h4101c036} /* (0, 20, 18) {real, imag} */,
  {32'h4105d3a4, 32'hc15570ea} /* (0, 20, 17) {real, imag} */,
  {32'hc115e8dc, 32'h3e89c380} /* (0, 20, 16) {real, imag} */,
  {32'h41136e20, 32'hc1639402} /* (0, 20, 15) {real, imag} */,
  {32'hc1a67274, 32'hbf940110} /* (0, 20, 14) {real, imag} */,
  {32'h41942d18, 32'hc06e6f44} /* (0, 20, 13) {real, imag} */,
  {32'h4155a995, 32'hc17044f1} /* (0, 20, 12) {real, imag} */,
  {32'hc20043fc, 32'hc206cf2a} /* (0, 20, 11) {real, imag} */,
  {32'h4203c18a, 32'hc0808690} /* (0, 20, 10) {real, imag} */,
  {32'h415f37de, 32'h411fec90} /* (0, 20, 9) {real, imag} */,
  {32'hc232f3a4, 32'hc20d263c} /* (0, 20, 8) {real, imag} */,
  {32'h423ac2cc, 32'h417bd3ee} /* (0, 20, 7) {real, imag} */,
  {32'hc25e277e, 32'h407b9380} /* (0, 20, 6) {real, imag} */,
  {32'h41838c04, 32'h41e0c9c1} /* (0, 20, 5) {real, imag} */,
  {32'hc1b871d8, 32'h42071de3} /* (0, 20, 4) {real, imag} */,
  {32'h412d6588, 32'h425ac7fe} /* (0, 20, 3) {real, imag} */,
  {32'hc1df7ec3, 32'hc1808a87} /* (0, 20, 2) {real, imag} */,
  {32'h416eec18, 32'hc1c07d1e} /* (0, 20, 1) {real, imag} */,
  {32'h42cbe502, 32'h428ff8b4} /* (0, 20, 0) {real, imag} */,
  {32'h41608a66, 32'hc2a69bae} /* (0, 19, 31) {real, imag} */,
  {32'h426c6904, 32'h41f3a8b6} /* (0, 19, 30) {real, imag} */,
  {32'h41e473a4, 32'hc24305cd} /* (0, 19, 29) {real, imag} */,
  {32'hc2830ad2, 32'hc08b9ef8} /* (0, 19, 28) {real, imag} */,
  {32'h40444cd6, 32'h409c940c} /* (0, 19, 27) {real, imag} */,
  {32'h42452db9, 32'h40ef5074} /* (0, 19, 26) {real, imag} */,
  {32'hc206267e, 32'h3ef15080} /* (0, 19, 25) {real, imag} */,
  {32'h421c85fc, 32'hc17168b9} /* (0, 19, 24) {real, imag} */,
  {32'hc2533b94, 32'hc1600899} /* (0, 19, 23) {real, imag} */,
  {32'h40d83714, 32'hc18dc2f0} /* (0, 19, 22) {real, imag} */,
  {32'hc21df1bc, 32'h3f3eedf0} /* (0, 19, 21) {real, imag} */,
  {32'h40fe65fa, 32'hc0dccc9c} /* (0, 19, 20) {real, imag} */,
  {32'h4071aa3a, 32'h40ce1e68} /* (0, 19, 19) {real, imag} */,
  {32'h40d6b49a, 32'h41497bfb} /* (0, 19, 18) {real, imag} */,
  {32'h407cc9cc, 32'h41071837} /* (0, 19, 17) {real, imag} */,
  {32'hc113b298, 32'h408f8faa} /* (0, 19, 16) {real, imag} */,
  {32'hc0b35a16, 32'h40b20c5e} /* (0, 19, 15) {real, imag} */,
  {32'hc16cde33, 32'h4119a38b} /* (0, 19, 14) {real, imag} */,
  {32'h417b183a, 32'hc18b1bcb} /* (0, 19, 13) {real, imag} */,
  {32'hc1bee2f2, 32'h41b3f0b7} /* (0, 19, 12) {real, imag} */,
  {32'h3f9e6860, 32'h40c3308a} /* (0, 19, 11) {real, imag} */,
  {32'h419e7c8d, 32'hc1ce9f00} /* (0, 19, 10) {real, imag} */,
  {32'h4083e99c, 32'hc12d8891} /* (0, 19, 9) {real, imag} */,
  {32'h41af76d9, 32'h41f87d74} /* (0, 19, 8) {real, imag} */,
  {32'h423d2422, 32'hc20466c7} /* (0, 19, 7) {real, imag} */,
  {32'hc2456f9b, 32'h4231a32e} /* (0, 19, 6) {real, imag} */,
  {32'h409dc83b, 32'h4256d35e} /* (0, 19, 5) {real, imag} */,
  {32'hc1b0e07c, 32'hc0f34ca0} /* (0, 19, 4) {real, imag} */,
  {32'hbfac5080, 32'hc17db88c} /* (0, 19, 3) {real, imag} */,
  {32'hc27755d8, 32'hc1c25e7c} /* (0, 19, 2) {real, imag} */,
  {32'hc2115e98, 32'h42aa331a} /* (0, 19, 1) {real, imag} */,
  {32'hc2456a4e, 32'h40bedf62} /* (0, 19, 0) {real, imag} */,
  {32'hc2b9f192, 32'h422327f5} /* (0, 18, 31) {real, imag} */,
  {32'hc1ab0b25, 32'hc0339790} /* (0, 18, 30) {real, imag} */,
  {32'h421fbe52, 32'h41269b76} /* (0, 18, 29) {real, imag} */,
  {32'hc2115a7a, 32'h40d9c366} /* (0, 18, 28) {real, imag} */,
  {32'hc1ce924e, 32'hc1314e89} /* (0, 18, 27) {real, imag} */,
  {32'hc0cfdf50, 32'hc1ab36c1} /* (0, 18, 26) {real, imag} */,
  {32'hc26a8272, 32'h3f2cdf68} /* (0, 18, 25) {real, imag} */,
  {32'h4247e426, 32'h4184be3d} /* (0, 18, 24) {real, imag} */,
  {32'h41b86183, 32'hc16148aa} /* (0, 18, 23) {real, imag} */,
  {32'hc09fc36a, 32'h3e7acda0} /* (0, 18, 22) {real, imag} */,
  {32'hbff4a0c0, 32'hc1059d1c} /* (0, 18, 21) {real, imag} */,
  {32'h4097df3d, 32'h41032aa5} /* (0, 18, 20) {real, imag} */,
  {32'h40a6edf2, 32'h41b245a5} /* (0, 18, 19) {real, imag} */,
  {32'h4047c8be, 32'hc109be8d} /* (0, 18, 18) {real, imag} */,
  {32'h41024b78, 32'h4027159c} /* (0, 18, 17) {real, imag} */,
  {32'hc07351dc, 32'h410f4da0} /* (0, 18, 16) {real, imag} */,
  {32'h3f5b6dc0, 32'hc1078f71} /* (0, 18, 15) {real, imag} */,
  {32'h408fbddd, 32'hc14a631f} /* (0, 18, 14) {real, imag} */,
  {32'hc0f0f59a, 32'hc0dbc21b} /* (0, 18, 13) {real, imag} */,
  {32'h4108a4a6, 32'hc08e8ce6} /* (0, 18, 12) {real, imag} */,
  {32'h4175acdc, 32'h410c57d4} /* (0, 18, 11) {real, imag} */,
  {32'h4097b67e, 32'h4178e9ba} /* (0, 18, 10) {real, imag} */,
  {32'hc10ee8ea, 32'h41c1e12f} /* (0, 18, 9) {real, imag} */,
  {32'h410e218e, 32'h41bfa52b} /* (0, 18, 8) {real, imag} */,
  {32'h40a1076c, 32'h4135541e} /* (0, 18, 7) {real, imag} */,
  {32'h412a7c9a, 32'h3e20fa80} /* (0, 18, 6) {real, imag} */,
  {32'hc11a5700, 32'h40ef56c5} /* (0, 18, 5) {real, imag} */,
  {32'h420d05dc, 32'h41c28fc6} /* (0, 18, 4) {real, imag} */,
  {32'h425aaee6, 32'h41c67e33} /* (0, 18, 3) {real, imag} */,
  {32'hc21caa7e, 32'hc0b4d004} /* (0, 18, 2) {real, imag} */,
  {32'hc0f82000, 32'hc22176a9} /* (0, 18, 1) {real, imag} */,
  {32'h40a4d566, 32'hc26f79b4} /* (0, 18, 0) {real, imag} */,
  {32'h418dad5f, 32'h417469e4} /* (0, 17, 31) {real, imag} */,
  {32'h4237d8b5, 32'h412f1398} /* (0, 17, 30) {real, imag} */,
  {32'h41304344, 32'h4137853e} /* (0, 17, 29) {real, imag} */,
  {32'hc20cdd7e, 32'h40e02cc2} /* (0, 17, 28) {real, imag} */,
  {32'hc2189716, 32'hc151c0d0} /* (0, 17, 27) {real, imag} */,
  {32'h415be322, 32'hc237746e} /* (0, 17, 26) {real, imag} */,
  {32'h41c07d0e, 32'hc18f1502} /* (0, 17, 25) {real, imag} */,
  {32'hbf48a8d8, 32'hc1a18851} /* (0, 17, 24) {real, imag} */,
  {32'hc18322b0, 32'h420c572c} /* (0, 17, 23) {real, imag} */,
  {32'hc1c04688, 32'hc12fb695} /* (0, 17, 22) {real, imag} */,
  {32'h4190d676, 32'h41678b45} /* (0, 17, 21) {real, imag} */,
  {32'h4196be30, 32'h41266248} /* (0, 17, 20) {real, imag} */,
  {32'hbf275450, 32'h4064c50e} /* (0, 17, 19) {real, imag} */,
  {32'h40ba1b3a, 32'h41266bc9} /* (0, 17, 18) {real, imag} */,
  {32'h40327928, 32'hbfe4256c} /* (0, 17, 17) {real, imag} */,
  {32'h401eaa4d, 32'h4108d0f8} /* (0, 17, 16) {real, imag} */,
  {32'hc0bf0c44, 32'hc148747c} /* (0, 17, 15) {real, imag} */,
  {32'h408e19a2, 32'h40f56226} /* (0, 17, 14) {real, imag} */,
  {32'hc06a0984, 32'hc0bc63d9} /* (0, 17, 13) {real, imag} */,
  {32'hc09550ba, 32'hc0d3ea58} /* (0, 17, 12) {real, imag} */,
  {32'hc0131bf0, 32'hc0a568e6} /* (0, 17, 11) {real, imag} */,
  {32'hc1b51f28, 32'hc0b78292} /* (0, 17, 10) {real, imag} */,
  {32'h4104bbe2, 32'h41885add} /* (0, 17, 9) {real, imag} */,
  {32'h4107d1f6, 32'hc1060600} /* (0, 17, 8) {real, imag} */,
  {32'hc0bce246, 32'h408ddd0e} /* (0, 17, 7) {real, imag} */,
  {32'h4196a987, 32'hc1bfdb63} /* (0, 17, 6) {real, imag} */,
  {32'hc2063f74, 32'hc15b4666} /* (0, 17, 5) {real, imag} */,
  {32'h422385d2, 32'h4086f6e4} /* (0, 17, 4) {real, imag} */,
  {32'hc20297e2, 32'hc211a686} /* (0, 17, 3) {real, imag} */,
  {32'hc1de1df6, 32'hc1a7d019} /* (0, 17, 2) {real, imag} */,
  {32'hc243245c, 32'h425dc235} /* (0, 17, 1) {real, imag} */,
  {32'h41151021, 32'h4087c483} /* (0, 17, 0) {real, imag} */,
  {32'h41c2d2ce, 32'h42119f2b} /* (0, 16, 31) {real, imag} */,
  {32'hc1fc9ea4, 32'h41b39b74} /* (0, 16, 30) {real, imag} */,
  {32'hc1d7931d, 32'h41e49801} /* (0, 16, 29) {real, imag} */,
  {32'h41b387cc, 32'h400311be} /* (0, 16, 28) {real, imag} */,
  {32'hc191e924, 32'hc225f412} /* (0, 16, 27) {real, imag} */,
  {32'h410ddfe5, 32'hbfa48abc} /* (0, 16, 26) {real, imag} */,
  {32'hc14cc88f, 32'hc0f8dbb9} /* (0, 16, 25) {real, imag} */,
  {32'hc1a9302c, 32'h41b028c6} /* (0, 16, 24) {real, imag} */,
  {32'hc209de33, 32'hbf6d1008} /* (0, 16, 23) {real, imag} */,
  {32'h3ff279f6, 32'hbefd3610} /* (0, 16, 22) {real, imag} */,
  {32'hbffa4e80, 32'hc0bc51a8} /* (0, 16, 21) {real, imag} */,
  {32'h410bdeaa, 32'hbf951f44} /* (0, 16, 20) {real, imag} */,
  {32'h402272c8, 32'h400dabb8} /* (0, 16, 19) {real, imag} */,
  {32'h41367d30, 32'hc110f4e5} /* (0, 16, 18) {real, imag} */,
  {32'hc06d0ae0, 32'hc0d82242} /* (0, 16, 17) {real, imag} */,
  {32'h3ff4cd40, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hc06d0ae0, 32'h40d82242} /* (0, 16, 15) {real, imag} */,
  {32'h41367d30, 32'h4110f4e5} /* (0, 16, 14) {real, imag} */,
  {32'h402272c8, 32'hc00dabb8} /* (0, 16, 13) {real, imag} */,
  {32'h410bdeaa, 32'h3f951f44} /* (0, 16, 12) {real, imag} */,
  {32'hbffa4e80, 32'h40bc51a8} /* (0, 16, 11) {real, imag} */,
  {32'h3ff279f6, 32'h3efd3610} /* (0, 16, 10) {real, imag} */,
  {32'hc209de33, 32'h3f6d1008} /* (0, 16, 9) {real, imag} */,
  {32'hc1a9302c, 32'hc1b028c6} /* (0, 16, 8) {real, imag} */,
  {32'hc14cc88f, 32'h40f8dbb9} /* (0, 16, 7) {real, imag} */,
  {32'h410ddfe5, 32'h3fa48abc} /* (0, 16, 6) {real, imag} */,
  {32'hc191e924, 32'h4225f412} /* (0, 16, 5) {real, imag} */,
  {32'h41b387cc, 32'hc00311be} /* (0, 16, 4) {real, imag} */,
  {32'hc1d7931d, 32'hc1e49801} /* (0, 16, 3) {real, imag} */,
  {32'hc1fc9ea4, 32'hc1b39b74} /* (0, 16, 2) {real, imag} */,
  {32'h41c2d2ce, 32'hc2119f2b} /* (0, 16, 1) {real, imag} */,
  {32'h426a627e, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'hc243245c, 32'hc25dc235} /* (0, 15, 31) {real, imag} */,
  {32'hc1de1df6, 32'h41a7d019} /* (0, 15, 30) {real, imag} */,
  {32'hc20297e2, 32'h4211a686} /* (0, 15, 29) {real, imag} */,
  {32'h422385d2, 32'hc086f6e4} /* (0, 15, 28) {real, imag} */,
  {32'hc2063f74, 32'h415b4666} /* (0, 15, 27) {real, imag} */,
  {32'h4196a987, 32'h41bfdb63} /* (0, 15, 26) {real, imag} */,
  {32'hc0bce246, 32'hc08ddd0e} /* (0, 15, 25) {real, imag} */,
  {32'h4107d1f6, 32'h41060600} /* (0, 15, 24) {real, imag} */,
  {32'h4104bbe2, 32'hc1885add} /* (0, 15, 23) {real, imag} */,
  {32'hc1b51f28, 32'h40b78292} /* (0, 15, 22) {real, imag} */,
  {32'hc0131bf0, 32'h40a568e6} /* (0, 15, 21) {real, imag} */,
  {32'hc09550ba, 32'h40d3ea58} /* (0, 15, 20) {real, imag} */,
  {32'hc06a0984, 32'h40bc63d9} /* (0, 15, 19) {real, imag} */,
  {32'h408e19a2, 32'hc0f56226} /* (0, 15, 18) {real, imag} */,
  {32'hc0bf0c44, 32'h4148747c} /* (0, 15, 17) {real, imag} */,
  {32'h401eaa4d, 32'hc108d0f8} /* (0, 15, 16) {real, imag} */,
  {32'h40327928, 32'h3fe4256c} /* (0, 15, 15) {real, imag} */,
  {32'h40ba1b3a, 32'hc1266bc9} /* (0, 15, 14) {real, imag} */,
  {32'hbf275450, 32'hc064c50e} /* (0, 15, 13) {real, imag} */,
  {32'h4196be30, 32'hc1266248} /* (0, 15, 12) {real, imag} */,
  {32'h4190d676, 32'hc1678b45} /* (0, 15, 11) {real, imag} */,
  {32'hc1c04688, 32'h412fb695} /* (0, 15, 10) {real, imag} */,
  {32'hc18322b0, 32'hc20c572c} /* (0, 15, 9) {real, imag} */,
  {32'hbf48a8d8, 32'h41a18851} /* (0, 15, 8) {real, imag} */,
  {32'h41c07d0e, 32'h418f1502} /* (0, 15, 7) {real, imag} */,
  {32'h415be322, 32'h4237746e} /* (0, 15, 6) {real, imag} */,
  {32'hc2189716, 32'h4151c0d0} /* (0, 15, 5) {real, imag} */,
  {32'hc20cdd7e, 32'hc0e02cc2} /* (0, 15, 4) {real, imag} */,
  {32'h41304344, 32'hc137853e} /* (0, 15, 3) {real, imag} */,
  {32'h4237d8b5, 32'hc12f1398} /* (0, 15, 2) {real, imag} */,
  {32'h418dad5f, 32'hc17469e4} /* (0, 15, 1) {real, imag} */,
  {32'h41151021, 32'hc087c483} /* (0, 15, 0) {real, imag} */,
  {32'hc0f82000, 32'h422176a9} /* (0, 14, 31) {real, imag} */,
  {32'hc21caa7e, 32'h40b4d004} /* (0, 14, 30) {real, imag} */,
  {32'h425aaee6, 32'hc1c67e33} /* (0, 14, 29) {real, imag} */,
  {32'h420d05dc, 32'hc1c28fc6} /* (0, 14, 28) {real, imag} */,
  {32'hc11a5700, 32'hc0ef56c5} /* (0, 14, 27) {real, imag} */,
  {32'h412a7c9a, 32'hbe20fa80} /* (0, 14, 26) {real, imag} */,
  {32'h40a1076c, 32'hc135541e} /* (0, 14, 25) {real, imag} */,
  {32'h410e218e, 32'hc1bfa52b} /* (0, 14, 24) {real, imag} */,
  {32'hc10ee8ea, 32'hc1c1e12f} /* (0, 14, 23) {real, imag} */,
  {32'h4097b67e, 32'hc178e9ba} /* (0, 14, 22) {real, imag} */,
  {32'h4175acdc, 32'hc10c57d4} /* (0, 14, 21) {real, imag} */,
  {32'h4108a4a6, 32'h408e8ce6} /* (0, 14, 20) {real, imag} */,
  {32'hc0f0f59a, 32'h40dbc21b} /* (0, 14, 19) {real, imag} */,
  {32'h408fbddd, 32'h414a631f} /* (0, 14, 18) {real, imag} */,
  {32'h3f5b6dc0, 32'h41078f71} /* (0, 14, 17) {real, imag} */,
  {32'hc07351dc, 32'hc10f4da0} /* (0, 14, 16) {real, imag} */,
  {32'h41024b78, 32'hc027159c} /* (0, 14, 15) {real, imag} */,
  {32'h4047c8be, 32'h4109be8d} /* (0, 14, 14) {real, imag} */,
  {32'h40a6edf2, 32'hc1b245a5} /* (0, 14, 13) {real, imag} */,
  {32'h4097df3d, 32'hc1032aa5} /* (0, 14, 12) {real, imag} */,
  {32'hbff4a0c0, 32'h41059d1c} /* (0, 14, 11) {real, imag} */,
  {32'hc09fc36a, 32'hbe7acda0} /* (0, 14, 10) {real, imag} */,
  {32'h41b86183, 32'h416148aa} /* (0, 14, 9) {real, imag} */,
  {32'h4247e426, 32'hc184be3d} /* (0, 14, 8) {real, imag} */,
  {32'hc26a8272, 32'hbf2cdf68} /* (0, 14, 7) {real, imag} */,
  {32'hc0cfdf50, 32'h41ab36c1} /* (0, 14, 6) {real, imag} */,
  {32'hc1ce924e, 32'h41314e89} /* (0, 14, 5) {real, imag} */,
  {32'hc2115a7a, 32'hc0d9c366} /* (0, 14, 4) {real, imag} */,
  {32'h421fbe52, 32'hc1269b76} /* (0, 14, 3) {real, imag} */,
  {32'hc1ab0b25, 32'h40339790} /* (0, 14, 2) {real, imag} */,
  {32'hc2b9f192, 32'hc22327f5} /* (0, 14, 1) {real, imag} */,
  {32'h40a4d566, 32'h426f79b4} /* (0, 14, 0) {real, imag} */,
  {32'hc2115e98, 32'hc2aa331a} /* (0, 13, 31) {real, imag} */,
  {32'hc27755d8, 32'h41c25e7c} /* (0, 13, 30) {real, imag} */,
  {32'hbfac5080, 32'h417db88c} /* (0, 13, 29) {real, imag} */,
  {32'hc1b0e07c, 32'h40f34ca0} /* (0, 13, 28) {real, imag} */,
  {32'h409dc83b, 32'hc256d35e} /* (0, 13, 27) {real, imag} */,
  {32'hc2456f9b, 32'hc231a32e} /* (0, 13, 26) {real, imag} */,
  {32'h423d2422, 32'h420466c7} /* (0, 13, 25) {real, imag} */,
  {32'h41af76d9, 32'hc1f87d74} /* (0, 13, 24) {real, imag} */,
  {32'h4083e99c, 32'h412d8891} /* (0, 13, 23) {real, imag} */,
  {32'h419e7c8d, 32'h41ce9f00} /* (0, 13, 22) {real, imag} */,
  {32'h3f9e6860, 32'hc0c3308a} /* (0, 13, 21) {real, imag} */,
  {32'hc1bee2f2, 32'hc1b3f0b7} /* (0, 13, 20) {real, imag} */,
  {32'h417b183a, 32'h418b1bcb} /* (0, 13, 19) {real, imag} */,
  {32'hc16cde33, 32'hc119a38b} /* (0, 13, 18) {real, imag} */,
  {32'hc0b35a16, 32'hc0b20c5e} /* (0, 13, 17) {real, imag} */,
  {32'hc113b298, 32'hc08f8faa} /* (0, 13, 16) {real, imag} */,
  {32'h407cc9cc, 32'hc1071837} /* (0, 13, 15) {real, imag} */,
  {32'h40d6b49a, 32'hc1497bfb} /* (0, 13, 14) {real, imag} */,
  {32'h4071aa3a, 32'hc0ce1e68} /* (0, 13, 13) {real, imag} */,
  {32'h40fe65fa, 32'h40dccc9c} /* (0, 13, 12) {real, imag} */,
  {32'hc21df1bc, 32'hbf3eedf0} /* (0, 13, 11) {real, imag} */,
  {32'h40d83714, 32'h418dc2f0} /* (0, 13, 10) {real, imag} */,
  {32'hc2533b94, 32'h41600899} /* (0, 13, 9) {real, imag} */,
  {32'h421c85fc, 32'h417168b9} /* (0, 13, 8) {real, imag} */,
  {32'hc206267e, 32'hbef15080} /* (0, 13, 7) {real, imag} */,
  {32'h42452db9, 32'hc0ef5074} /* (0, 13, 6) {real, imag} */,
  {32'h40444cd6, 32'hc09c940c} /* (0, 13, 5) {real, imag} */,
  {32'hc2830ad2, 32'h408b9ef8} /* (0, 13, 4) {real, imag} */,
  {32'h41e473a4, 32'h424305cd} /* (0, 13, 3) {real, imag} */,
  {32'h426c6904, 32'hc1f3a8b6} /* (0, 13, 2) {real, imag} */,
  {32'h41608a66, 32'h42a69bae} /* (0, 13, 1) {real, imag} */,
  {32'hc2456a4e, 32'hc0bedf62} /* (0, 13, 0) {real, imag} */,
  {32'h416eec18, 32'h41c07d1e} /* (0, 12, 31) {real, imag} */,
  {32'hc1df7ec3, 32'h41808a87} /* (0, 12, 30) {real, imag} */,
  {32'h412d6588, 32'hc25ac7fe} /* (0, 12, 29) {real, imag} */,
  {32'hc1b871d8, 32'hc2071de3} /* (0, 12, 28) {real, imag} */,
  {32'h41838c04, 32'hc1e0c9c1} /* (0, 12, 27) {real, imag} */,
  {32'hc25e277e, 32'hc07b9380} /* (0, 12, 26) {real, imag} */,
  {32'h423ac2cc, 32'hc17bd3ee} /* (0, 12, 25) {real, imag} */,
  {32'hc232f3a4, 32'h420d263c} /* (0, 12, 24) {real, imag} */,
  {32'h415f37de, 32'hc11fec90} /* (0, 12, 23) {real, imag} */,
  {32'h4203c18a, 32'h40808690} /* (0, 12, 22) {real, imag} */,
  {32'hc20043fc, 32'h4206cf2a} /* (0, 12, 21) {real, imag} */,
  {32'h4155a995, 32'h417044f1} /* (0, 12, 20) {real, imag} */,
  {32'h41942d18, 32'h406e6f44} /* (0, 12, 19) {real, imag} */,
  {32'hc1a67274, 32'h3f940110} /* (0, 12, 18) {real, imag} */,
  {32'h41136e20, 32'h41639402} /* (0, 12, 17) {real, imag} */,
  {32'hc115e8dc, 32'hbe89c380} /* (0, 12, 16) {real, imag} */,
  {32'h4105d3a4, 32'h415570ea} /* (0, 12, 15) {real, imag} */,
  {32'hc0ec7ed6, 32'hc101c036} /* (0, 12, 14) {real, imag} */,
  {32'hc1cd3914, 32'hc0eedc82} /* (0, 12, 13) {real, imag} */,
  {32'h4182f946, 32'h41338c37} /* (0, 12, 12) {real, imag} */,
  {32'hc088fdf0, 32'h3fb7c890} /* (0, 12, 11) {real, imag} */,
  {32'hc0ab47d0, 32'h419ebfe4} /* (0, 12, 10) {real, imag} */,
  {32'hc010c938, 32'hc1cf7d2c} /* (0, 12, 9) {real, imag} */,
  {32'h41b99174, 32'hbda26100} /* (0, 12, 8) {real, imag} */,
  {32'hbe881540, 32'hc19ec235} /* (0, 12, 7) {real, imag} */,
  {32'h404815a0, 32'hc149d800} /* (0, 12, 6) {real, imag} */,
  {32'h4103e0ff, 32'hc1be7b77} /* (0, 12, 5) {real, imag} */,
  {32'h41334599, 32'hc1eaad07} /* (0, 12, 4) {real, imag} */,
  {32'hc29a42f6, 32'hc2308486} /* (0, 12, 3) {real, imag} */,
  {32'hc177025a, 32'h42378cdc} /* (0, 12, 2) {real, imag} */,
  {32'h429dea4d, 32'h42655b5d} /* (0, 12, 1) {real, imag} */,
  {32'h42cbe502, 32'hc28ff8b4} /* (0, 12, 0) {real, imag} */,
  {32'h420bb78f, 32'hc0b9f904} /* (0, 11, 31) {real, imag} */,
  {32'h41be8f2f, 32'hc222955b} /* (0, 11, 30) {real, imag} */,
  {32'h40cb56bc, 32'h41bd2de2} /* (0, 11, 29) {real, imag} */,
  {32'hc1b89c60, 32'h4234f9e7} /* (0, 11, 28) {real, imag} */,
  {32'h42082225, 32'h402b0f0c} /* (0, 11, 27) {real, imag} */,
  {32'h4180c565, 32'hc2298559} /* (0, 11, 26) {real, imag} */,
  {32'hbf4f4da0, 32'hc2367224} /* (0, 11, 25) {real, imag} */,
  {32'h42125dc4, 32'hc18972de} /* (0, 11, 24) {real, imag} */,
  {32'h41394567, 32'hc2806aec} /* (0, 11, 23) {real, imag} */,
  {32'hc1d1d48e, 32'h403f685b} /* (0, 11, 22) {real, imag} */,
  {32'h411fee58, 32'h424ce3d4} /* (0, 11, 21) {real, imag} */,
  {32'h406f8264, 32'h412fae48} /* (0, 11, 20) {real, imag} */,
  {32'h401cdbb4, 32'hc19ab163} /* (0, 11, 19) {real, imag} */,
  {32'hc0f35d60, 32'hbfd13190} /* (0, 11, 18) {real, imag} */,
  {32'hbf38dac0, 32'h4150c562} /* (0, 11, 17) {real, imag} */,
  {32'hc1715f56, 32'h41c16fc6} /* (0, 11, 16) {real, imag} */,
  {32'hbf965940, 32'h41a4afed} /* (0, 11, 15) {real, imag} */,
  {32'h411f0ba4, 32'hc1f681ef} /* (0, 11, 14) {real, imag} */,
  {32'hc1d61a1c, 32'h40435fe8} /* (0, 11, 13) {real, imag} */,
  {32'hc122cb65, 32'hc17403f0} /* (0, 11, 12) {real, imag} */,
  {32'h4191f004, 32'hc10296d6} /* (0, 11, 11) {real, imag} */,
  {32'hc2257789, 32'h3edf2f58} /* (0, 11, 10) {real, imag} */,
  {32'h41d1d6a2, 32'hc1c334ef} /* (0, 11, 9) {real, imag} */,
  {32'h412824f6, 32'h3fd17230} /* (0, 11, 8) {real, imag} */,
  {32'hc21202b0, 32'h421f0160} /* (0, 11, 7) {real, imag} */,
  {32'hc221594c, 32'h4245f477} /* (0, 11, 6) {real, imag} */,
  {32'hc255225f, 32'hbfa24548} /* (0, 11, 5) {real, imag} */,
  {32'hc23d9f70, 32'hc21611c5} /* (0, 11, 4) {real, imag} */,
  {32'h42058806, 32'hc1f54182} /* (0, 11, 3) {real, imag} */,
  {32'hc22de9c8, 32'h4245aecd} /* (0, 11, 2) {real, imag} */,
  {32'hc1703e0c, 32'hc15765aa} /* (0, 11, 1) {real, imag} */,
  {32'h40a04798, 32'hc266990d} /* (0, 11, 0) {real, imag} */,
  {32'h41dba34a, 32'h41189f78} /* (0, 10, 31) {real, imag} */,
  {32'h4201bd1c, 32'h41433b13} /* (0, 10, 30) {real, imag} */,
  {32'hc32e7cac, 32'hc218230c} /* (0, 10, 29) {real, imag} */,
  {32'hc2b4a30e, 32'hc2dad9a3} /* (0, 10, 28) {real, imag} */,
  {32'h4250ea82, 32'hc1b41717} /* (0, 10, 27) {real, imag} */,
  {32'h41c30f34, 32'hc0453c40} /* (0, 10, 26) {real, imag} */,
  {32'hc26588da, 32'hc1c427ba} /* (0, 10, 25) {real, imag} */,
  {32'hc1e062e2, 32'hc1a0dc52} /* (0, 10, 24) {real, imag} */,
  {32'h419e739a, 32'h418445a4} /* (0, 10, 23) {real, imag} */,
  {32'h40d0731e, 32'h3e90e6c0} /* (0, 10, 22) {real, imag} */,
  {32'hbf631560, 32'hc29678d0} /* (0, 10, 21) {real, imag} */,
  {32'h411ce918, 32'h40b8cc84} /* (0, 10, 20) {real, imag} */,
  {32'h420ff7d0, 32'hc08a8e5c} /* (0, 10, 19) {real, imag} */,
  {32'hc13b27f8, 32'h41168345} /* (0, 10, 18) {real, imag} */,
  {32'h417975b5, 32'hc008f0c0} /* (0, 10, 17) {real, imag} */,
  {32'hc181505c, 32'hc022dde4} /* (0, 10, 16) {real, imag} */,
  {32'hc1883e5e, 32'h4138523c} /* (0, 10, 15) {real, imag} */,
  {32'h414d812c, 32'hc15b3501} /* (0, 10, 14) {real, imag} */,
  {32'h4194d257, 32'hc2095596} /* (0, 10, 13) {real, imag} */,
  {32'hc2983931, 32'h40d065fc} /* (0, 10, 12) {real, imag} */,
  {32'h4224a790, 32'h40e3fe98} /* (0, 10, 11) {real, imag} */,
  {32'hc20d91b7, 32'h4254bfba} /* (0, 10, 10) {real, imag} */,
  {32'h4228747b, 32'hc1ce5042} /* (0, 10, 9) {real, imag} */,
  {32'hc13f12c4, 32'h42300091} /* (0, 10, 8) {real, imag} */,
  {32'h42ef60db, 32'h415a4c59} /* (0, 10, 7) {real, imag} */,
  {32'hc1b83a82, 32'h3fa79740} /* (0, 10, 6) {real, imag} */,
  {32'hc1fd4b14, 32'hc1e06bd3} /* (0, 10, 5) {real, imag} */,
  {32'h41fc8b07, 32'hc261e242} /* (0, 10, 4) {real, imag} */,
  {32'h41ffd6dc, 32'h41706b46} /* (0, 10, 3) {real, imag} */,
  {32'h420dcfdc, 32'h418e697c} /* (0, 10, 2) {real, imag} */,
  {32'hc2263727, 32'hc2cb6011} /* (0, 10, 1) {real, imag} */,
  {32'hc1d8c0f8, 32'h41a493c0} /* (0, 10, 0) {real, imag} */,
  {32'hc3062800, 32'h4368271b} /* (0, 9, 31) {real, imag} */,
  {32'h4321d7bc, 32'h42bcdea7} /* (0, 9, 30) {real, imag} */,
  {32'h4253e906, 32'hc26a8521} /* (0, 9, 29) {real, imag} */,
  {32'hc227ddee, 32'h41222d28} /* (0, 9, 28) {real, imag} */,
  {32'h41838a25, 32'h4191afa4} /* (0, 9, 27) {real, imag} */,
  {32'h411327ca, 32'h416358be} /* (0, 9, 26) {real, imag} */,
  {32'hc13f4ad0, 32'h4146a634} /* (0, 9, 25) {real, imag} */,
  {32'hc0a5a76e, 32'hc0a218d4} /* (0, 9, 24) {real, imag} */,
  {32'hc257cb94, 32'h426a5d34} /* (0, 9, 23) {real, imag} */,
  {32'hc1f5ae3a, 32'hc14f5bd1} /* (0, 9, 22) {real, imag} */,
  {32'hc20561c4, 32'hc11c3264} /* (0, 9, 21) {real, imag} */,
  {32'h425cab36, 32'hbee57c60} /* (0, 9, 20) {real, imag} */,
  {32'h41423097, 32'h419c434d} /* (0, 9, 19) {real, imag} */,
  {32'h4181bfff, 32'hc1501372} /* (0, 9, 18) {real, imag} */,
  {32'hc1b19550, 32'h41b87536} /* (0, 9, 17) {real, imag} */,
  {32'h4212c282, 32'h41e08dcd} /* (0, 9, 16) {real, imag} */,
  {32'hc02cdc40, 32'hc1250533} /* (0, 9, 15) {real, imag} */,
  {32'hc14bccd2, 32'h414ed8de} /* (0, 9, 14) {real, imag} */,
  {32'hc1a4926a, 32'h41281056} /* (0, 9, 13) {real, imag} */,
  {32'hc10e07f6, 32'hc1e08a6c} /* (0, 9, 12) {real, imag} */,
  {32'hc25b9f74, 32'h41efee26} /* (0, 9, 11) {real, imag} */,
  {32'hc1a9f208, 32'hc1f22ccc} /* (0, 9, 10) {real, imag} */,
  {32'h424ebbda, 32'h42945372} /* (0, 9, 9) {real, imag} */,
  {32'hc103e4bd, 32'hc135fd66} /* (0, 9, 8) {real, imag} */,
  {32'h41989fcc, 32'h428db7ee} /* (0, 9, 7) {real, imag} */,
  {32'hc1fd3527, 32'hc101a268} /* (0, 9, 6) {real, imag} */,
  {32'hc2155132, 32'h42ddc24b} /* (0, 9, 5) {real, imag} */,
  {32'hc23483f2, 32'hc19748df} /* (0, 9, 4) {real, imag} */,
  {32'hc1a7aebc, 32'hc21357a3} /* (0, 9, 3) {real, imag} */,
  {32'hc26ae34e, 32'hc3108018} /* (0, 9, 2) {real, imag} */,
  {32'hc267e1cc, 32'hc31c3167} /* (0, 9, 1) {real, imag} */,
  {32'hc29957b5, 32'hc1b97287} /* (0, 9, 0) {real, imag} */,
  {32'hc2afb2c5, 32'hc1a8dd53} /* (0, 8, 31) {real, imag} */,
  {32'hc1cfa075, 32'h42b0558d} /* (0, 8, 30) {real, imag} */,
  {32'h4245b5e1, 32'hc30af2b7} /* (0, 8, 29) {real, imag} */,
  {32'h42a3f06c, 32'h430a76e0} /* (0, 8, 28) {real, imag} */,
  {32'hc29618d2, 32'hc2845eb2} /* (0, 8, 27) {real, imag} */,
  {32'h42602a2b, 32'h41e8c361} /* (0, 8, 26) {real, imag} */,
  {32'h4315ef87, 32'hc2c6c38e} /* (0, 8, 25) {real, imag} */,
  {32'hc24f5afe, 32'hc282ac6b} /* (0, 8, 24) {real, imag} */,
  {32'h423a60ff, 32'hc22e6279} /* (0, 8, 23) {real, imag} */,
  {32'hc2854029, 32'hc223c59c} /* (0, 8, 22) {real, imag} */,
  {32'h419e05b0, 32'h428052a2} /* (0, 8, 21) {real, imag} */,
  {32'hc13f0920, 32'h41d54d6a} /* (0, 8, 20) {real, imag} */,
  {32'hc18a05ea, 32'hc175bf54} /* (0, 8, 19) {real, imag} */,
  {32'h4205db46, 32'h41f653db} /* (0, 8, 18) {real, imag} */,
  {32'hc12339e1, 32'h411d4172} /* (0, 8, 17) {real, imag} */,
  {32'h41666edc, 32'h41941fef} /* (0, 8, 16) {real, imag} */,
  {32'h409abea2, 32'h4225d996} /* (0, 8, 15) {real, imag} */,
  {32'h41472f46, 32'hbf9b6e90} /* (0, 8, 14) {real, imag} */,
  {32'hc203a6c3, 32'hc2224261} /* (0, 8, 13) {real, imag} */,
  {32'h40cb1310, 32'h41a0e156} /* (0, 8, 12) {real, imag} */,
  {32'h42f83d82, 32'hc1a26c06} /* (0, 8, 11) {real, imag} */,
  {32'h41b43cbd, 32'h42c45d68} /* (0, 8, 10) {real, imag} */,
  {32'hc26c0677, 32'h42ae6d10} /* (0, 8, 9) {real, imag} */,
  {32'hc29589c9, 32'hc27fb001} /* (0, 8, 8) {real, imag} */,
  {32'hc21ec3bb, 32'h41a488c4} /* (0, 8, 7) {real, imag} */,
  {32'hc01c6c20, 32'hc2a4a017} /* (0, 8, 6) {real, imag} */,
  {32'hc10663a0, 32'hc25ed42d} /* (0, 8, 5) {real, imag} */,
  {32'hc2c6e4dc, 32'hc2096526} /* (0, 8, 4) {real, imag} */,
  {32'hc27020e9, 32'h4301ad05} /* (0, 8, 3) {real, imag} */,
  {32'hc16b8a4e, 32'hc24148e6} /* (0, 8, 2) {real, imag} */,
  {32'hc2b26391, 32'hc151b302} /* (0, 8, 1) {real, imag} */,
  {32'hc234d54f, 32'h4120a06a} /* (0, 8, 0) {real, imag} */,
  {32'hc2bc0cc0, 32'h41000840} /* (0, 7, 31) {real, imag} */,
  {32'h412aa03d, 32'hc30a1c47} /* (0, 7, 30) {real, imag} */,
  {32'hc2da88d6, 32'h40a85870} /* (0, 7, 29) {real, imag} */,
  {32'hc3350df4, 32'h40debcf1} /* (0, 7, 28) {real, imag} */,
  {32'hc2b1b5e7, 32'h432140c7} /* (0, 7, 27) {real, imag} */,
  {32'hc287b750, 32'h4197b21c} /* (0, 7, 26) {real, imag} */,
  {32'hc118599e, 32'h41d92498} /* (0, 7, 25) {real, imag} */,
  {32'hc246af30, 32'hc2a09c09} /* (0, 7, 24) {real, imag} */,
  {32'hc28f8a28, 32'h43076c44} /* (0, 7, 23) {real, imag} */,
  {32'hc01050b8, 32'h42913f02} /* (0, 7, 22) {real, imag} */,
  {32'h4255044f, 32'h421fd681} /* (0, 7, 21) {real, imag} */,
  {32'h41f65a88, 32'hc2167622} /* (0, 7, 20) {real, imag} */,
  {32'h3efa92c0, 32'h425e1527} /* (0, 7, 19) {real, imag} */,
  {32'hc0e6a14c, 32'hc19ccebd} /* (0, 7, 18) {real, imag} */,
  {32'h40e2a432, 32'hc0a66c0e} /* (0, 7, 17) {real, imag} */,
  {32'h418ce69a, 32'h4114df30} /* (0, 7, 16) {real, imag} */,
  {32'hc19b0db8, 32'h41bfa57c} /* (0, 7, 15) {real, imag} */,
  {32'hc228b0ae, 32'h3ff8e110} /* (0, 7, 14) {real, imag} */,
  {32'hc1d41d5d, 32'h41cab616} /* (0, 7, 13) {real, imag} */,
  {32'hc22bc450, 32'hc0dda930} /* (0, 7, 12) {real, imag} */,
  {32'hc1668cd4, 32'h41a58c8e} /* (0, 7, 11) {real, imag} */,
  {32'hc1cd4faf, 32'h42a080a4} /* (0, 7, 10) {real, imag} */,
  {32'h428e3b6a, 32'h42938395} /* (0, 7, 9) {real, imag} */,
  {32'hc050f750, 32'hc2add5fb} /* (0, 7, 8) {real, imag} */,
  {32'hc2891048, 32'hc21a2a74} /* (0, 7, 7) {real, imag} */,
  {32'h43060aa0, 32'hc290f07d} /* (0, 7, 6) {real, imag} */,
  {32'h42bc516f, 32'h42532e8c} /* (0, 7, 5) {real, imag} */,
  {32'h42c98ae0, 32'h41300228} /* (0, 7, 4) {real, imag} */,
  {32'hc110cac0, 32'h43236b70} /* (0, 7, 3) {real, imag} */,
  {32'hc0b5b20e, 32'hc1cc8308} /* (0, 7, 2) {real, imag} */,
  {32'h42207900, 32'h42260e94} /* (0, 7, 1) {real, imag} */,
  {32'h40cd34ee, 32'hc2bc2ce6} /* (0, 7, 0) {real, imag} */,
  {32'h424dd6c8, 32'h42e3b94f} /* (0, 6, 31) {real, imag} */,
  {32'hc28b6ebd, 32'hc1d4e67a} /* (0, 6, 30) {real, imag} */,
  {32'h4181c17e, 32'hc2fda3ab} /* (0, 6, 29) {real, imag} */,
  {32'h41e194cc, 32'hc2e7abca} /* (0, 6, 28) {real, imag} */,
  {32'hc1a883de, 32'hc188efd7} /* (0, 6, 27) {real, imag} */,
  {32'h42449dce, 32'h42bd39c2} /* (0, 6, 26) {real, imag} */,
  {32'hc207a6bb, 32'h41324f30} /* (0, 6, 25) {real, imag} */,
  {32'hc287ad30, 32'h40e9bb38} /* (0, 6, 24) {real, imag} */,
  {32'h424c3c77, 32'h42724dd8} /* (0, 6, 23) {real, imag} */,
  {32'h429cd514, 32'hc00df510} /* (0, 6, 22) {real, imag} */,
  {32'hc236d1c9, 32'hc1a2a16f} /* (0, 6, 21) {real, imag} */,
  {32'hc0a2296a, 32'hc14b46ae} /* (0, 6, 20) {real, imag} */,
  {32'hc0d06248, 32'hc213e77c} /* (0, 6, 19) {real, imag} */,
  {32'h424059f2, 32'h41affab0} /* (0, 6, 18) {real, imag} */,
  {32'h3efd5560, 32'hc2631f07} /* (0, 6, 17) {real, imag} */,
  {32'hc14dde48, 32'hc1abedf3} /* (0, 6, 16) {real, imag} */,
  {32'h403f26ac, 32'hc0649930} /* (0, 6, 15) {real, imag} */,
  {32'hc0c11024, 32'h41519af8} /* (0, 6, 14) {real, imag} */,
  {32'h423f38d9, 32'hc1ef8def} /* (0, 6, 13) {real, imag} */,
  {32'h411fa239, 32'h4120a36e} /* (0, 6, 12) {real, imag} */,
  {32'hc04da890, 32'h413fe662} /* (0, 6, 11) {real, imag} */,
  {32'hc236859e, 32'h41b1d28e} /* (0, 6, 10) {real, imag} */,
  {32'hc18113fa, 32'h4294ba74} /* (0, 6, 9) {real, imag} */,
  {32'hc23e2ce3, 32'hc2b80c98} /* (0, 6, 8) {real, imag} */,
  {32'h42d5ffbc, 32'h4318bfc5} /* (0, 6, 7) {real, imag} */,
  {32'hc2835d40, 32'hc25e628c} /* (0, 6, 6) {real, imag} */,
  {32'hc0ed82a6, 32'h3fc8ce90} /* (0, 6, 5) {real, imag} */,
  {32'h428949e1, 32'h40df73a0} /* (0, 6, 4) {real, imag} */,
  {32'h423ebfaf, 32'hc213d2be} /* (0, 6, 3) {real, imag} */,
  {32'h40f5dbbc, 32'hc28c06c4} /* (0, 6, 2) {real, imag} */,
  {32'hc2812561, 32'h41c48754} /* (0, 6, 1) {real, imag} */,
  {32'h429d7e87, 32'hc01d38d0} /* (0, 6, 0) {real, imag} */,
  {32'h413f646f, 32'h42920b1b} /* (0, 5, 31) {real, imag} */,
  {32'hc342cc6a, 32'hc304d3d2} /* (0, 5, 30) {real, imag} */,
  {32'h426f3f58, 32'h423b200d} /* (0, 5, 29) {real, imag} */,
  {32'hc2d5b18e, 32'h42bf4066} /* (0, 5, 28) {real, imag} */,
  {32'hc1a86fe8, 32'h42e6b42f} /* (0, 5, 27) {real, imag} */,
  {32'h41b5e852, 32'h4291f5af} /* (0, 5, 26) {real, imag} */,
  {32'hc2144bce, 32'h42ab2b3e} /* (0, 5, 25) {real, imag} */,
  {32'hc2bab9ce, 32'hc245e0b3} /* (0, 5, 24) {real, imag} */,
  {32'hc15b3c90, 32'h42839f56} /* (0, 5, 23) {real, imag} */,
  {32'hc2b5c056, 32'hc0c54540} /* (0, 5, 22) {real, imag} */,
  {32'h401cd714, 32'hc291fb77} /* (0, 5, 21) {real, imag} */,
  {32'h417fe458, 32'hc29b64bb} /* (0, 5, 20) {real, imag} */,
  {32'hc0e38038, 32'h41ea3f24} /* (0, 5, 19) {real, imag} */,
  {32'hc1c0a70a, 32'h41c753de} /* (0, 5, 18) {real, imag} */,
  {32'hc1be9f55, 32'hc20815e5} /* (0, 5, 17) {real, imag} */,
  {32'hc1f21e2e, 32'hc09147c0} /* (0, 5, 16) {real, imag} */,
  {32'hc1d93c3b, 32'h411a757c} /* (0, 5, 15) {real, imag} */,
  {32'hc1afd92a, 32'h421f36f5} /* (0, 5, 14) {real, imag} */,
  {32'h421d34d5, 32'h41eb0d34} /* (0, 5, 13) {real, imag} */,
  {32'h41e9d158, 32'hc2815bb1} /* (0, 5, 12) {real, imag} */,
  {32'hc1e9c264, 32'hc2deb5bd} /* (0, 5, 11) {real, imag} */,
  {32'h4084f518, 32'h42326166} /* (0, 5, 10) {real, imag} */,
  {32'h41f6aa0e, 32'hc20c4c99} /* (0, 5, 9) {real, imag} */,
  {32'h42c53a54, 32'h4299b8a8} /* (0, 5, 8) {real, imag} */,
  {32'h42ab0509, 32'h425474db} /* (0, 5, 7) {real, imag} */,
  {32'hc1a4700e, 32'h42004834} /* (0, 5, 6) {real, imag} */,
  {32'h423d3d48, 32'h4284a6f1} /* (0, 5, 5) {real, imag} */,
  {32'hc1bb4ada, 32'h4280016e} /* (0, 5, 4) {real, imag} */,
  {32'hc24d56ac, 32'hc2ae1ab8} /* (0, 5, 3) {real, imag} */,
  {32'h42db17fc, 32'hc232db6b} /* (0, 5, 2) {real, imag} */,
  {32'h415de393, 32'h433ea688} /* (0, 5, 1) {real, imag} */,
  {32'hc2d347a8, 32'h42ef783e} /* (0, 5, 0) {real, imag} */,
  {32'hc161885f, 32'hc3101885} /* (0, 4, 31) {real, imag} */,
  {32'hc34d33e9, 32'h42f2aebe} /* (0, 4, 30) {real, imag} */,
  {32'hc2f34898, 32'hc2671ff1} /* (0, 4, 29) {real, imag} */,
  {32'hc237be26, 32'hc1958871} /* (0, 4, 28) {real, imag} */,
  {32'h41999cd4, 32'hc327b0e0} /* (0, 4, 27) {real, imag} */,
  {32'hc3272bdc, 32'hc2b00534} /* (0, 4, 26) {real, imag} */,
  {32'h422a10ce, 32'h432b9020} /* (0, 4, 25) {real, imag} */,
  {32'h431d3349, 32'hc3343331} /* (0, 4, 24) {real, imag} */,
  {32'hc24e8422, 32'hc2b8a8e0} /* (0, 4, 23) {real, imag} */,
  {32'hc1b72450, 32'h413dc914} /* (0, 4, 22) {real, imag} */,
  {32'h41907e14, 32'h424cc938} /* (0, 4, 21) {real, imag} */,
  {32'h42a547c9, 32'h42239546} /* (0, 4, 20) {real, imag} */,
  {32'hc219bddf, 32'hc1c9ee2a} /* (0, 4, 19) {real, imag} */,
  {32'hc1640326, 32'hc209e4df} /* (0, 4, 18) {real, imag} */,
  {32'h41bc1ed4, 32'h41d0043b} /* (0, 4, 17) {real, imag} */,
  {32'hc2188e80, 32'h41cc5be2} /* (0, 4, 16) {real, imag} */,
  {32'hc22d30d6, 32'hc1a56855} /* (0, 4, 15) {real, imag} */,
  {32'hbf5c2760, 32'h415127fc} /* (0, 4, 14) {real, imag} */,
  {32'h427174df, 32'h42315f4f} /* (0, 4, 13) {real, imag} */,
  {32'hc29183c1, 32'hc214a6fe} /* (0, 4, 12) {real, imag} */,
  {32'h42a98e4c, 32'h42994f57} /* (0, 4, 11) {real, imag} */,
  {32'h4235e490, 32'h40d53ba8} /* (0, 4, 10) {real, imag} */,
  {32'h42beff6b, 32'hc24079fb} /* (0, 4, 9) {real, imag} */,
  {32'h41fa456e, 32'hc1cae9d0} /* (0, 4, 8) {real, imag} */,
  {32'hc3200156, 32'hc1ce27d4} /* (0, 4, 7) {real, imag} */,
  {32'hc31544fc, 32'h43469a9e} /* (0, 4, 6) {real, imag} */,
  {32'h42636f7c, 32'hc321566c} /* (0, 4, 5) {real, imag} */,
  {32'h435ff93c, 32'hc23e760c} /* (0, 4, 4) {real, imag} */,
  {32'hc2b2e114, 32'h4293d46c} /* (0, 4, 3) {real, imag} */,
  {32'h4364c487, 32'hc0c0be08} /* (0, 4, 2) {real, imag} */,
  {32'h4202d43f, 32'h429c3656} /* (0, 4, 1) {real, imag} */,
  {32'hc3068865, 32'hc27e4191} /* (0, 4, 0) {real, imag} */,
  {32'h40a07534, 32'hc2f26d7c} /* (0, 3, 31) {real, imag} */,
  {32'h42399068, 32'hc1af83d0} /* (0, 3, 30) {real, imag} */,
  {32'hc2ab15bc, 32'h42aaeb3e} /* (0, 3, 29) {real, imag} */,
  {32'h4134f49c, 32'h42534a88} /* (0, 3, 28) {real, imag} */,
  {32'h41fd6164, 32'hc309dca9} /* (0, 3, 27) {real, imag} */,
  {32'hc2f9699d, 32'h426c6183} /* (0, 3, 26) {real, imag} */,
  {32'hc343ba7b, 32'h42fc6ce0} /* (0, 3, 25) {real, imag} */,
  {32'h42136c9c, 32'hc236056e} /* (0, 3, 24) {real, imag} */,
  {32'hc2596b69, 32'hc2d52a4a} /* (0, 3, 23) {real, imag} */,
  {32'hc12a4f29, 32'h41290fd8} /* (0, 3, 22) {real, imag} */,
  {32'hc29d864c, 32'hc166c4c8} /* (0, 3, 21) {real, imag} */,
  {32'hbf8531e0, 32'h41f6216a} /* (0, 3, 20) {real, imag} */,
  {32'h41d577c0, 32'h41ea65ee} /* (0, 3, 19) {real, imag} */,
  {32'hc04c9600, 32'hc25f8743} /* (0, 3, 18) {real, imag} */,
  {32'h423b18f4, 32'hc08ab520} /* (0, 3, 17) {real, imag} */,
  {32'h40ff7390, 32'hc213115a} /* (0, 3, 16) {real, imag} */,
  {32'h4125d43e, 32'hc1109c38} /* (0, 3, 15) {real, imag} */,
  {32'h42362b08, 32'h424c8475} /* (0, 3, 14) {real, imag} */,
  {32'hc1193c5c, 32'hc19078c8} /* (0, 3, 13) {real, imag} */,
  {32'h42b8efa8, 32'hc2cfee72} /* (0, 3, 12) {real, imag} */,
  {32'h40b703c0, 32'hc27b4e1e} /* (0, 3, 11) {real, imag} */,
  {32'hc05f6b3c, 32'h42384564} /* (0, 3, 10) {real, imag} */,
  {32'hc0f0fff8, 32'hc2656a95} /* (0, 3, 9) {real, imag} */,
  {32'hc2e24200, 32'h42801ea5} /* (0, 3, 8) {real, imag} */,
  {32'hc1925178, 32'hc2d0ff18} /* (0, 3, 7) {real, imag} */,
  {32'hc2e1124f, 32'hc181d03a} /* (0, 3, 6) {real, imag} */,
  {32'hc32ed360, 32'h43132f7f} /* (0, 3, 5) {real, imag} */,
  {32'h42945764, 32'h430f5652} /* (0, 3, 4) {real, imag} */,
  {32'h410e71b0, 32'hc2af889e} /* (0, 3, 3) {real, imag} */,
  {32'h41e33a80, 32'h43547c98} /* (0, 3, 2) {real, imag} */,
  {32'h411a31d2, 32'h42c207b8} /* (0, 3, 1) {real, imag} */,
  {32'h4332e222, 32'h427a93da} /* (0, 3, 0) {real, imag} */,
  {32'hc1b81d1c, 32'hbf4de400} /* (0, 2, 31) {real, imag} */,
  {32'h42b45046, 32'hc2d8886d} /* (0, 2, 30) {real, imag} */,
  {32'h431eb629, 32'h42e53c96} /* (0, 2, 29) {real, imag} */,
  {32'h423905ee, 32'h42a15a3e} /* (0, 2, 28) {real, imag} */,
  {32'h420b8ac6, 32'hc29b65cc} /* (0, 2, 27) {real, imag} */,
  {32'h423f2e7b, 32'h42c053e0} /* (0, 2, 26) {real, imag} */,
  {32'h4293f668, 32'h408bc050} /* (0, 2, 25) {real, imag} */,
  {32'h426e143b, 32'h431ea28e} /* (0, 2, 24) {real, imag} */,
  {32'hc2c8cbba, 32'h415f8e88} /* (0, 2, 23) {real, imag} */,
  {32'hc22509f0, 32'hc1cf0196} /* (0, 2, 22) {real, imag} */,
  {32'h4218c4f9, 32'h41b0d462} /* (0, 2, 21) {real, imag} */,
  {32'h42662f09, 32'hc22086a4} /* (0, 2, 20) {real, imag} */,
  {32'hc2aebab8, 32'h420bc80a} /* (0, 2, 19) {real, imag} */,
  {32'h40a94a70, 32'hc229795d} /* (0, 2, 18) {real, imag} */,
  {32'h417977a7, 32'hc23b4544} /* (0, 2, 17) {real, imag} */,
  {32'h41124280, 32'hc04c7c90} /* (0, 2, 16) {real, imag} */,
  {32'h40f18db6, 32'hc12c5a2e} /* (0, 2, 15) {real, imag} */,
  {32'h41f39ad6, 32'hc1d49f1e} /* (0, 2, 14) {real, imag} */,
  {32'hc22a5c74, 32'hc174d250} /* (0, 2, 13) {real, imag} */,
  {32'h416d1c3c, 32'h41be803b} /* (0, 2, 12) {real, imag} */,
  {32'hc140e48c, 32'h40b9d1e6} /* (0, 2, 11) {real, imag} */,
  {32'hbf522380, 32'h4271724b} /* (0, 2, 10) {real, imag} */,
  {32'h429e980a, 32'h43080882} /* (0, 2, 9) {real, imag} */,
  {32'hc22b40ad, 32'hc28d5710} /* (0, 2, 8) {real, imag} */,
  {32'h42845e4e, 32'hc2e01453} /* (0, 2, 7) {real, imag} */,
  {32'h42c135e2, 32'h434af9d2} /* (0, 2, 6) {real, imag} */,
  {32'hc331f380, 32'hc2ea86dc} /* (0, 2, 5) {real, imag} */,
  {32'h42f7a94d, 32'hc3501255} /* (0, 2, 4) {real, imag} */,
  {32'hc19d89f0, 32'hc2874e6a} /* (0, 2, 3) {real, imag} */,
  {32'h420003e0, 32'h42790026} /* (0, 2, 2) {real, imag} */,
  {32'h4083fa26, 32'h42ec9816} /* (0, 2, 1) {real, imag} */,
  {32'hc25e719e, 32'hc1a0901c} /* (0, 2, 0) {real, imag} */,
  {32'h41d10b9a, 32'hc1e5df66} /* (0, 1, 31) {real, imag} */,
  {32'h4160f548, 32'h42ec5784} /* (0, 1, 30) {real, imag} */,
  {32'h429d7f74, 32'hc2786760} /* (0, 1, 29) {real, imag} */,
  {32'hc2f63434, 32'hc258ede2} /* (0, 1, 28) {real, imag} */,
  {32'h4354cbc1, 32'h41c693dc} /* (0, 1, 27) {real, imag} */,
  {32'h431d356a, 32'hc2f769aa} /* (0, 1, 26) {real, imag} */,
  {32'hc2e736e3, 32'h405aa32e} /* (0, 1, 25) {real, imag} */,
  {32'hc22f5f64, 32'hc2b11a9a} /* (0, 1, 24) {real, imag} */,
  {32'hbeb9f1c0, 32'hc2ce36a3} /* (0, 1, 23) {real, imag} */,
  {32'h42d969bb, 32'h3e868f80} /* (0, 1, 22) {real, imag} */,
  {32'hc13730ee, 32'h4284aed5} /* (0, 1, 21) {real, imag} */,
  {32'h4204aac7, 32'h42ab9f22} /* (0, 1, 20) {real, imag} */,
  {32'h420625ff, 32'hc25e60de} /* (0, 1, 19) {real, imag} */,
  {32'hc0cf38b0, 32'h424dc3fe} /* (0, 1, 18) {real, imag} */,
  {32'h41fb6fa6, 32'h41b786d2} /* (0, 1, 17) {real, imag} */,
  {32'hc13e7b18, 32'hc222b66c} /* (0, 1, 16) {real, imag} */,
  {32'h40742c50, 32'h42847f10} /* (0, 1, 15) {real, imag} */,
  {32'hc1c7a8c4, 32'h40920a54} /* (0, 1, 14) {real, imag} */,
  {32'h426c0e05, 32'hc22107a0} /* (0, 1, 13) {real, imag} */,
  {32'h42a67dce, 32'hc2916894} /* (0, 1, 12) {real, imag} */,
  {32'hc1cbe943, 32'h42963721} /* (0, 1, 11) {real, imag} */,
  {32'hc2eb4f0f, 32'hc24bbb5f} /* (0, 1, 10) {real, imag} */,
  {32'hc20f9360, 32'h4285def1} /* (0, 1, 9) {real, imag} */,
  {32'h429a8577, 32'hbe72e900} /* (0, 1, 8) {real, imag} */,
  {32'h40fc13f0, 32'hc165e264} /* (0, 1, 7) {real, imag} */,
  {32'hc2bed0db, 32'hc3130e9d} /* (0, 1, 6) {real, imag} */,
  {32'hc2612f44, 32'h4323705a} /* (0, 1, 5) {real, imag} */,
  {32'hc1f962b6, 32'hc3243ac4} /* (0, 1, 4) {real, imag} */,
  {32'hc135e7f4, 32'hc24941b2} /* (0, 1, 3) {real, imag} */,
  {32'hc2f83c21, 32'hc287eed2} /* (0, 1, 2) {real, imag} */,
  {32'hbf89dc18, 32'hc249447b} /* (0, 1, 1) {real, imag} */,
  {32'h42120475, 32'hc19c254c} /* (0, 1, 0) {real, imag} */,
  {32'hc29375ee, 32'h41b5d0e7} /* (0, 0, 31) {real, imag} */,
  {32'hc20c545b, 32'h43070598} /* (0, 0, 30) {real, imag} */,
  {32'h428cbff0, 32'hc2a0f730} /* (0, 0, 29) {real, imag} */,
  {32'h4087e878, 32'hc3834dca} /* (0, 0, 28) {real, imag} */,
  {32'h41c35daa, 32'h42b76ac8} /* (0, 0, 27) {real, imag} */,
  {32'h42e6f1c2, 32'hc273f8f8} /* (0, 0, 26) {real, imag} */,
  {32'h42861ac9, 32'hc30d917d} /* (0, 0, 25) {real, imag} */,
  {32'h4296c380, 32'hc1df69b0} /* (0, 0, 24) {real, imag} */,
  {32'h41dcf09b, 32'h4260eaec} /* (0, 0, 23) {real, imag} */,
  {32'hc2995574, 32'h3ed19c00} /* (0, 0, 22) {real, imag} */,
  {32'hc27766cb, 32'h41e14116} /* (0, 0, 21) {real, imag} */,
  {32'hc1f5df28, 32'hc2751e62} /* (0, 0, 20) {real, imag} */,
  {32'h41d3e0ca, 32'hc265dc6f} /* (0, 0, 19) {real, imag} */,
  {32'h41e3a7ca, 32'h41a076dc} /* (0, 0, 18) {real, imag} */,
  {32'hc14a58ae, 32'h41bf9c5b} /* (0, 0, 17) {real, imag} */,
  {32'h41d0d634, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'hc14a58ae, 32'hc1bf9c5b} /* (0, 0, 15) {real, imag} */,
  {32'h41e3a7ca, 32'hc1a076dc} /* (0, 0, 14) {real, imag} */,
  {32'h41d3e0ca, 32'h4265dc6f} /* (0, 0, 13) {real, imag} */,
  {32'hc1f5df28, 32'h42751e62} /* (0, 0, 12) {real, imag} */,
  {32'hc27766cb, 32'hc1e14116} /* (0, 0, 11) {real, imag} */,
  {32'hc2995574, 32'hbed19c00} /* (0, 0, 10) {real, imag} */,
  {32'h41dcf09b, 32'hc260eaec} /* (0, 0, 9) {real, imag} */,
  {32'h4296c380, 32'h41df69b0} /* (0, 0, 8) {real, imag} */,
  {32'h42861ac9, 32'h430d917d} /* (0, 0, 7) {real, imag} */,
  {32'h42e6f1c2, 32'h4273f8f8} /* (0, 0, 6) {real, imag} */,
  {32'h41c35daa, 32'hc2b76ac8} /* (0, 0, 5) {real, imag} */,
  {32'h4087e878, 32'h43834dca} /* (0, 0, 4) {real, imag} */,
  {32'h428cbff0, 32'h42a0f730} /* (0, 0, 3) {real, imag} */,
  {32'hc20c545b, 32'hc3070598} /* (0, 0, 2) {real, imag} */,
  {32'hc29375ee, 32'hc1b5d0e7} /* (0, 0, 1) {real, imag} */,
  {32'hb7000000, 32'h00000000} /* (0, 0, 0) {real, imag} */};
