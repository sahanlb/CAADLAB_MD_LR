-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Zd36aWReYK0nM7ydOkLmkLjhNB5sS/EmdD5BkDO1CH/RZhl0WDGis+N7lLADG8xwW18/ljS+As1F
yjp29eGdBSEJQYJgSFc86RegajJq+vVWkRugl65ANyzfh1RuK3eXv6ollTNLGSvoW2ve5iFWpKDW
RnzNvZgwQWflc2ql1hr50fGaiWrNq4NiH256yUPIw3eSOSW0zMEmdP1LBu8q40OdpYlirEcvsKMC
zuy0qtrgc+6kZxSe0ik3aUkbcZpSbpk3QVd2passPen2V4KpWJbe2WQ3sjZPEDko7kxVCj9uJMMC
cIZEaRoZF1pQbwypZvQ3nSFFs9LB1ARHW9Q9zA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5712)
`protect data_block
bLedi0hbbbo4AB4tCvwiO+E+FTAleVkrmuUPT1ISPBL1q+AdaEMndtSgROYHmcF5WAq6dQO+bXIY
Ws4tRaARkRRcvYiftATvOyVunaHsoact0+o5yBSz7pdgK+xZw/MzDUj9pkyQr9h9+QlAW5VfW2qw
zJQlY8buLRhOdZ05RdH9ieq0Jki66azPrrpVLD+HYWCVaSWeLD8nqITtCDL9jcvKQsOzOhR9lPQL
T6EOFTFORf3Li7qa5cZrXoccWFW6wahhaxQq7CTN5FWFSX3+fnbAQn27Jwdip4uch+Vu4oVBKI0t
0TiTb4Fh549pL+cvdTcZHJklBap4MaRWFX174lA4ot9fF1FdMO7ORv5za4jeCfW8ie0n2JptkmXe
4ce8bxnfbZxG47dLBPQVkk/QHYAySnFWhG4PZcSQ2D+ve4Qm+6Tkxjz3tPqsgLRr/p4sMYTcEDV6
BEhKlrkZRrqPLxrwASKt+uXeJvHhdwf55NHCWE84Dof3ZA2i7yMosE8mYuPG2EXLeJLLdZZwTjkv
a7QOqqVzjnZsOr69ysKLRSbfNo6icsLPx4Ir7+X+KHBXYawF3Vyk2pWBr45Y50i7wvLHGrtXo6ow
l/PfDtht581rZdsYcmH4GgzQ0sj2hzgIz7y81TyM7VcqRpRGMzQw+MVy4DdjAd0XNFV+BnMb6VAw
Noe9tLa4OMt7XT7tcK7s5pWekGN188kXj5kKIzEZkWEKfphY6VybgRJVsh8Su7+81XmaP/6Gy/TL
5nZMnkA8/n7FTK+gJakZwK9oxDlLx45fAme+oNSZVLzouJgwt3jz167HBZOa7K4UY68HIwTaO5da
WBct73HZZy8A/h5fyujtUl3d98EAHUiAdhhUtG7zCRLgG+kaZSMea6LtMmx+OVYJu/saohSw84lp
ATs45JZkN8Mt5PrOKBcHgFrz18m6nMkuHmJ1SCGH0UI/32DHZPkRjwO1P+vufpZRywW+ebrey1wf
fLYlAsT310Xx9MI85HRsyae27TbUsmG4aXPFwdVCIOmRmOtm8qetSVrEZ8CT+cPO4o12mor6jEDk
x+gZ/rAJN8JrRPL2Gj3tDJlq6wzocIYkXHAOJCIwGWKrsYOQi+PbkWo9x3qSkgztJ99kTO3Ndlzl
9vmtTIL4yLTST56NcTNkwd1LtYBV8Qlfq5WwVwtC42HI2c+52ERfReAZJoY5W/7rdr1LvIr+2FN7
WA6AymdYdMgRnufGfw5ahjvAPKvx0qE4SXRPtE+/9wZ4bsTUgZz/RAKPQh7+SgG8qFG7TTKlpBmD
hr4FcTb2+5olDAQr37W2hzlrZaeVqHqOMR/Ge6ltGkFnzknX8rimCKLd1Rp/aMWt2/qJZgCsj3ab
sp5w59zmuGKGTSHQ3+DSAbsUp4VnF4V+oTdbuuVzvYMEf7ZeApnyfrTswUTYlEoMl8wjDTWSQOOX
KbJdzTOx9+5eyWxzzqicqDQDKcq688Y5+I8xJe8SsQRrQtmh65M/x0aPPfa/V6v1TpezcPoMu53n
TZsfEWS8OOMnE3hLrjdAb9GNGk1OLp3jywTG0P1MW4mZ7i/3G+GXBtsL8IZnnrsWsrs1gSgirrr0
kPTZ/pUlG4lUvcBZLkR4tni5opvvZQBAqY5j1HTGqTa7iECdhpQKgq2p2lMzjpgLdh07TpBbtC5H
Qp2MNEdQmID1WIli4JGk2gHoIOTHysCbVee7QptS9bKXL4CagHbkUGhTTwxskfWmEhbusTU5R9OR
y3xgWYyDdLqEayw41tnD6OrQOaz6V9+OQrUCSv3a9sTZYajpFT8n39RzFlPuA1X11lXoYN2k+hlJ
TGYpstBzITUh6C2U87N+Yj3AKh5EzFaTCM9rqMU0XyBJYaTvoXjT8izFamttR/EYRana7dIFhT5f
7aS1WTN2HM99zXhtrNSBe6dOsWWDhZPeH/dcd2/d0WO0Lv0fark4QrEidFtG4bNz+d+FK0r6t/R+
Ig74x/kdBy4JUxeygj5tDdWEZ7+S2rJIFVmfQ4+woLV2qyeJEg44vXVLVAbIO5IwUkk3BE/ypU/o
IyZ6o2nCQLtiM6VXg2GAPkbWsylgXuaAY7xeftBCYoGKo/Tqa0Xb7bzs2zR5nzgJ6FigpDWVYvDO
JM+pU3rvePlMQNhZSiS63pZJcDZKIhcnTXHHILdcjv/uHAxp1JxwHbAXxCSDUw02DMPpo47tRghX
a26fQO5c4QAlS7pBSDLroVqKsndwpUxRlgbsIzyXfdQbO9+xHGqwC1xtqvdSvTy9iYHb07IV/4H5
Hnrx2kpJEAhDn4PGozidEo7VOaZuUjYXgOiWKTvt6bGDz5G0Y3eCXREMlg5k/CBcoa8h+7zTZKVJ
v0D5WVFnOPD96mPfZDcxskqRm76zDC+3ubfE1ChSp4Daw4/E0/ZJjBygeVXu1f4aTMM0uvTYlamo
+KB3Y/0pIOdCD5cdgPyQKbG7KX2b2TJdZ8rQ7NMR2iGz09ffpMSGeOwzzsAifhhqjD8yFPV5ej8U
XVCAwgW16xmyvBfQNFTtPD8ERakCa4gjcwY+cNQW5GEY8vyuhGKlYjjQlcAu5pOc34mVtCgWRWXN
38oTNH9ICbQh7kTHVnj8i6aiNcSlfjMnhaRALenDBMo8AigU5D5zMxmeSSWEapJvXj0yySzupfHa
2MU/eAON35Ffku2WlLLdckwP6nnU8DBtPrf6z1u6ltonoPNUBBytKM5qrsjghE4uRwEQ28aGIHN9
GrZ3Qs9gUpa1BrhI+T+gsF/+1Vui+rhKSNR+BkcbwflVnalOsnMLgZK2MTF41Yyaws5V9/pYKIls
AHRKf/rYa7pkl1gEYye5ebsrGvzlWBX0DOSHovCXsWX/As5Vq6RJN6uRDhMznGKAq9b3v40RL5F0
g1eUlvGBE3iiRKFgOgtI7jGSMVQOguTXAfClnIE0j5EBLCUhTU00gV0QbRSwmI9VcTgRcH5E019h
98wyK8zPSyoNpkXzfHX70eDoGeVCVTnP66GX2fR/kl8e6QiI7KXr556GDrVcP+mVOdFPAHnLbv3p
SM2p2aHbkbA26vjjewy//iJ7LqpzjnfAJI5mU2ywk+G7rBu7s3dU/XF555+tLHgS0RTnZpYVXkie
mL8p3rAX1YDoDmb1wdypbfPFRQ8CFrkR1dB9lHCp+0FRvUlFQ8+JZYINW49v/YS/zalejEpctQyu
zwsSNerPQBaKodMJR8wUZO0afUjX1pM7WEtoJU6yjCj7duHbwAJ7wncU9IsGup1hLSp0qjHpn6wh
gjw3ewZueopiujDILfK3zS90ScIjEgItLfDijELKA8/HUR/Jj4FauRIlZ4k3aocYkVWYjN2kw6D0
QgvyZKpn9+bVkSikcXxetkdrLL9qi0XwN0Xdq1SxXSAzDqwjtrG0ytGd7zWTaE/OS4hN1sZgp/iS
bWKYYsWSUoDr1rQKYUMqO9pAOd0B06mvncy6fM+49c+C6O908WgfvkGYXNE7Oba4W8+KkiknLScy
ntqr3ECnkkokFDdoz9DfvHtJ7KDDJRmsUqnTW+xfzGD2p5IwFwX9rpOvCKC3G6EMlcyGdEgZsfbk
ak5g/6gMXgkIYFjZu5ac/J2tFVonP+eEd6HEEf4o9wXXPoI8FZmyupnMqSqj1TkbYD5COeVdI5Nm
1uuXq+Cdu4md0slA472XLtbscmIKKE1WRwEaQWJptQe35VguWjIJ2KJKw1WYlXnPxWN8xoM76jGV
VIZodzhh3hGYDnwSFCWUyXd6yPnNehgAHgR5KYoUrT4XiZL7bFNm3PzIiVi2EO8Hw0HTAEIMxC8o
x+Zjfy3gb6oN1kcuhT2zm1ck8l1udwg4D3KAtwtvcXdZKhSwofbzoopHWKXLbNBKbH5rBAZDMefd
7MMbvm2Mi9EdzSlOWcjw5iPYcKFlaVmZEEHjNlPIK91TQa3ixsEvm5ucEGti92JxGIERr7tIy7ju
RoNpEWy3HcNub7/FUb7i72+XRc1OhhB6Vkiz1fuGbDce5iih7RxpHYZ+pinbtoePCHLn6NZYW5l2
i97QKjfl85QkbdVAEpVssdenJdX2gXc0d6RbgHgDkV8W8tSc3MKPynEs0g62d0MMsiqkFUxWnbKk
jXlJUd6nVQ/6Zq0zOTymMVppD02ZF71gknZbaB2eIZkV0/pVSVeJtlQc5X2Z0htfUPDDHKH7hnEK
6INZU1KgeWVTmKLWoxeFMvvBlNZnhh5lnUytkEkavRwuD1CZ1PuAgpRzVBwmubb4w1/R2mrGPPdR
MgED9txGRxubr2LZ+lHJCALHJIP/KORSuTvLl8zjxurLutxHGxeYtdx5cZWd4h3rvk10bbq7FNhr
K9r0y2dSnvoLxAQrJoDKC/NXGDbjW8LJ4YmF6ks4AtZji7yi/uureYRWrvNDf7JzY8BQRGxDJBAr
chPZxlIoLGmiIdLxsC0yysHHnDG+oF2eoc5I3ctHHgegpk/3mt2rIQr4Qhma5HDwV5nftgfkvgEC
smV9s7yQHgNat7yKWRsosi+0y5Kcysmg8K4g1/LtmU8/zy/SWMurtnlBl+pZlH5hVI9UAZuUf8d+
lhM2G9/OToMk8B9L266vekPrgr56HhHbINAY+W8QEAaAs2r7UjOLv9BYV2AlIgAIRTU2I7I3os8v
TTfIGO+05lvTUb7Ma5biabLtN/gJjEjT2OnJfFrjChCtLcZvDI/YOHJzJuto4VEjWIduvpzPUQUz
xqbaQotdTbHRylNeS29FsPW3C6+YCNFJI1u1qMWgxwstxuMRFg8mGixEgNSX4xsE+HUUFzanyhBN
COZZCsyUsHbKFdr85j5KNUqX56lrOd64RzDV4zCIQT/Jf8cpoOOMl8pcZ4lYGwPhCx0XsmkZZcpa
2YDe25hNIjO0cRdJK5CWZ0XgFE12N98bCq4Y0gZ4dnl1W9kSKmP4Zjktc7p7leGnB3yw7zvQOukp
3/VCdolk1AIli9DqyO83QVCKD1wRugueA3BL4DtyWy8x3bsF8QdzWb0vH/aRw4FM1uPNjQHixIhd
W1RQpbtAGxwvHdPcPnXwkUll17sAVVFLm6hVtdQs78vXd98SU8iTkmGq1NdU9WqbJRcRI4gKRueM
+O8hQlvwFd3BNiSTZDn5n3XFwuTMXj/uq1ys81gVjPo6SKgvrAhQq5IAuI1Pw7o2UyBawWEBCH65
2IyVUX24dIL0COlA2lOXyYPqygn2Qvnd1zTKFtLSa8jhAUwE82yKTIkoTYv8Fx0lO2LzmfxKzigB
hWEAYRwERB9ImN776yuCDBqlPqRw8OdOs3fQc4zjIoo1VyQuD7UQWuuIuv69iR0tTBRoGIIglI6D
H0bse6r0zCKPfP/1rePKizXMv4/zTWQRW1Yy0+BspLN6Yh8ZiNWFSezPqf8DHE9t+LeJpxeX5hWC
ebYQX0hg4wKX4TRVVxi6afso2HULYkxFB/KR4xouQPWAVrFiOUO/WBjgFmcsHfmxzyt0ZfQQbk9/
4iv05m8XMxR9g/t8E1h2Bg531pmd9W6dLlK0rMlyL00wfpX02sljAujwoou5xnLrRe0Rqua6Hr9A
4y1JfMbz7oZ9feVw/GORC93Bty8aPTAp7jTZNwIBwmgoVYqdS0/350IBkkSrq2fIgMKfC1TGWARW
OlsbICgBb8Lk1LtK0enyF6921JhN15S/A5jslnAV/nLKzcTn+z4qZzG24X6f+dA0vXIpR2WRvr7W
Ba7NhiARnTkXddEJrM6FYdzo2G27QDqZ9BYtBT91bYmGP/3+psRUzVD3Sqo3skNkOms15+cpIbjv
0sFazz1V9CT/EJL2NkqzlgDxJITtX5hYRRcMV/EsX0VrrmsSFK24X6t/Qgnsm0HjOP78kNEIUHCF
ZK3rVYtkFqjEwGrW7Qqa+FBKNBiWnVZVvRUFSOUXvrzjerGZJeyKQUdU6YDZpXf+vOR0xjHBoBoM
I8N0LJz7OMQI/k4/BV6mAqrzEAZWDhWdt80FOL5Mkd9iCnjpV6nkBiwxT1lZNEvEP0F5ny+OC34D
xFvNro0MueNKLpwzCoHR7Bq+Mes2xfDA+BL/hMfZfRe1w4s+YSroMOndeaf+kbqjq3u0D5HUcf7Q
ydHU+eZz7rXSHPLsDpc6IvedwuTJoB8SAyoVm8h4Z59CjQdfzLVmetIyikXCMzU9vuhEnhRdxY6v
+FlpAo/ty4l3mvFb3rUwKRYzUc5CXo+gyQJ6ymIPfFkPNariHH8qw1fEZTtziOt9MRc0siTJw8uu
JZsZufm63dfAR04uqQGWl3/2zyRzNgSztzduLmou1XNzItSMXcWfPh/7JWn/fPFe8NDkokwcG7zi
dr9FmB2iH9Sf+aGpqhNwDN7qibkiRuQ+KbYZxKGGjeHEr7RnhtjdpEM54o8Oga3g1WBi/A0ZtDvt
9Pl/yCx2Hazi345NzymvBb3qxzIzKLVwvkd1gHQvdhPe3MGj6fYqSg87x936m232ftxxspnuBfsW
fW/Ec1n1JEO1n2UqkcbjfKSNFKPjrsvJhF0u3EdnEL4Nds8R10hMXqULIyb2JkM9x83bZQ7/5CGD
pJ2b08SPwi6lzHlWJOe0hGZk8L/3OnpOIROdc/FZbKG6dlDEkpS8eA+qX+aZGE4G6NZNLPlMtf0H
6GclRVQ++ADN6rHlhUQvPFnSof6YlXa7Dzy+ITGHUKCQr3c/M42bE7xszzlRDNSwyOgXUDq8U9fw
/KZYiVcBUpZsIos0xwfIWKKu4YkPUR4r4SksFbhy629Ffepp3USbqg0m4pAGOrbghT2CQFqFRnOO
0q0a9DelzdaZsVRLtSIQz4Mc3LQsUdCUCgLaq8uVWXwFvRzMcNwY24RUVaXfMJrbxo8oVPtpdKW/
0ZTpVrrimNJpqMNr347OJFO4U2bUgeWplmnBjPzdJnevyb83Pwnqc71o6ahDl0Mw9AFjAIJZPS9x
Ewi7bYmzHNVdwfnV5I+IPqigr7r6wONQqMM85zu8hGM1UrTUFiFxqMUz0dge5tJONGbJdkB7qv53
//PTPtkQf4ls58W+6bEF71NkbXP5EMEDfxa35kErs8VM84ByIOSjg4Io59YWqkF6VZg0EBW0B0ex
8T6QP31Wg941KbKUNQ6YuaTxEPHb+St9D188lvrEBKb0ksF6fFsJ9Mwo9ASw44YtcYr5zfonlzcE
bWYWasBayf4pd8Viw8Dcd6OAn16sJgnCNe066Ayq+Y3XvfLD1x1dclVEaldNaAGDqDwPnKrYw7o4
7np8CkoN+0caGvK+u8logYMqd39DenS6DxbXO17tSG0WVv4lG5ri+elBR1Mv2V6YBFT4rLYxAWDg
LsDHHL94jNfxK8w33OU+Bdke2e1nY3ldS4aasOLBsq7XA0kUHiF0dC7+DLp4cLI+/IJ3sTBbKOXE
6XbmeNK8MiNrvVQNak8JYTo3dEnz/BMewbLMUID48uF3DjoYXuX1ZsMZbk33SKYlcQNr8VHY8i0V
zxZUguGoyBMrQW7uWxgJW3z73Q5TZysruSchoOjYd2jzxgGHihS0Eam8vj+frFPfY9QLdRMJ3Kqn
PQBIzsdEF90cpLilwhdChzj3o+wsDKOo/RVD3KPdqjZIFtUQcFV/RGvP1FqiH1a8lBV2MxmItQTB
SO6qIN3CzJ2zbyvw
`protect end_protected
