-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
lKYvsrdjHf2KKoorersytj1ElmzW3faWszL6cxTFL75jo/iHTLL7r5gmuudblAxH
f/Ix9mwbZ6ag67NlAcImjvBDDQVosJCZuErxkyMgylZZvtdrL8GWnEqOZaqJlH8a
nvhDt5eMyii6DCVV0eVWMpaSb17qFsvHclg4ZWZhSaaLdHujU7GUDA==
--pragma protect end_key_block
--pragma protect digest_block
djmwH5LUwgpWIj8P75+lC7xiyHw=
--pragma protect end_digest_block
--pragma protect data_block
HuyE+1tD2m62XsIfyMAZRldxsO/13Uvy8qsSXUSR5cGRWZPkLhmVLIICp7EBBoI3
8sm+nOY5UKDciDco2Jx07o9r28sOldt4THtLs9lFIMW+qVvg/T1yrbdfaEf0VUZE
OgsB0pjGehcxhTXLFGjdh+z7xmFbkXT7hEozWKu2mj9QUoatYvv+k38ao7MsEZwg
lnjIjShmptxnd/v283ChxeOtZ0aMKUg9XGJ9OiZtEnbrskmtn3WLBILFnruE7qn2
srccXT0GBDBhohMP0rDs6YElXzskb5Ak/Ne/PGLvij8yG3YgkIvbY1dsF+jlvl+q
GB5UTUlXyHlOlIQ3KTwTBome8OONEvYVpPZ6zubw2RVWQlIHGl/qm1sERv7nR1qM
4mzRjBfjLHYwW+tuRLGxJSR2OQa5GBLCvlv75/li93Vw/oIYrO1W8P0ETNM7CQzP
2u7BBFdCo6rEfQLL3+0LiDz4yXH8vW8PP9qACKGKR3jCPNT281VIwJO7e68/nIDa
ybJF2teATUUNg9lf7o67+d2DDgq1hSBX64JN8l1DWJqIcSE96nVPJaSRBwH43JtW
WPTVMynImMJ8zEvl06RjUGSUrzJqMCjwmMG911ziqromJRKlRifOhkfvyApV8Ia4
u/e34NCEG/rXQaQiGWyWzgh3TlNpzkGUP/KTghRjR39vbMhMyB3fS480oU+eZ4pH
iJ929rlfoFgnlw12mhNuSudQHSz1stcWXukZUwZYG1GnrTglf82Oguo3SXtXCUrg
ZDaF9h2Z06zvTTsPRYvLexmvkdot1Wv5UwM2X5xs6EUtS2FaPDJMtQq4vZEwjkB9
fM1L9C81Su+qQBDq7xmXyd8l0MM/9iIh9U+QcKFexbqqjfVc1odBX81lxKR1GgHV
OqRMc/lChWFZ8IhCG+lHJ85FqsnQ53DzueWaCxwoTDRmKM9lM0UyK+c4br+WopAt
fBR455WJe7KEmdP4b75lKcLRAJSCRGVh3K6HX6puqTLLIdJrQkypDk5YcTY3eXER
az3rmH+i0EPEnZxMB5OxVbBbRYWG380fUWAXYSw+f6dgOh5pKEQdotcTkUwkx6hZ
a6ct5rfrpa3lsBbO6y7iML79dUzfuzpb4w/G7EBXlufZ2A0cqRlom74RR2GP5p/Y
1yw99Ni4nPKvp72JxMhdPY9UpPuMjVnHfoFGUCm3Q2LCYA0tvH9Vk+tE+o5XN2aS
rVZs1h1BQhM00taoUJYGjJrCqJlRlP48sPCXVAB95+qLY+RswAKEjpTURZ/CXKAs
Ppq/diZ0El0OsPOr1mdGfNl1M5Id107vIdqpfix+dIw50fsXHMHWFPPFNmLHgs4C
tc6LLwqwg59bJN8BWJ2j2ZrYbHdoPI5FDb3syNLknFwB2h00szJLSGMtoQHVgblo
fRJRoqGEuCY5RA4Mjo0X9QlgqxEB0zrZH2+8uc9Lkxkqm/t5wt/1NbJlvLqMfFmn
0iY1M5AqnkVpsX38g4arDL+3t6/8d0kNvOnaiu6AY9PXM0jTrsP8WGfHstHdUUNa
nbMoSiZ/tnG/1FtUyLjb/udzF1D92aI79blxiqc+nBvXcK48ai57uptvr1tJPb0+
E3/sgftX3Algru5erdGT+yK3GQMBhG6dWZ/JKWUe6l02XqQnewJjtGBMUhSb6wI1
FzdS+XGR0g/wHy943Jxax3HmbEYKONtLs3J3SwVOrJrX/lFHKXtiVPIP4WyY6lXe
F+fq998hr0kjFrvTzoGCqXOKdjosy07rfAaORcpJEjq3DQc1j/ndITDdWBJ4wuH2
Xqjs4RMGLlQ+XzL1VDBUPUcM1tY0b27Nx0mVKnU8aMDTKB1+dvYxMkG3BSkmUcjV
+ArXxzzFDAgt1cDkguCabNbJ8ootOdTwjKGI3JsWKYO3GmezqwHE60jCGMA9rT6D
+uwwczyE9PuQamuQHrn/y8DlwhRZszsF9Bs4AKVb36L7TCSyCxrJYR8+oHdexDxv
LMFEqAoxWHYe1JoYCL770M9InfRZaK4fgnWJIXMu0q9m6JAQNyO/AdjxHhovB7/V
Iyp0+ewOfg18P49KsDUWCCOskTgEKwTnfyrxzIj3hIPA4Tf5KGW4E/UC1eUF01vE
/fYC8SIbZNGEbzzWTYSNSLyUcG8yNP6Fea1g23Gq2qX7e3SesLdykksiolsSnt9E
eucnvibj9Mi7l1bUE+id5Jeh+9MJ74TlIQ5q9mIOpjbZHEI7Km9YKNouSk3x20tw
tOycGGtLpyPYuyhpi0/XwT69pLbz7Z+rPJbQDQh0gK8QzzOMf940Srsh9ntz6gBk
ZLsv2hS2Er8+6vwEf63JRIMYURF/cu33Oj711jAW13MkNXJMuGXw+FMz1I3C9fi1
g/ZtxQw0dJ1rgjOQKMeYeZr1Erkj9J0858ZsO5tcFedZLrv73kEhtq7usU3G7JHn
0G6aejlrC8Ina+Eqnz/2btffqp1+K7OPj9/pWBW11s6JtYlaj3MvG801zHIYlpnk
MYtEE/Ss4fmzQgwHkTWSWBS2bJUWFZ3XqshXg1ePtV3Pe5ObV0xORAObkRkvoUam
8ox7jA6u9t0NK4H4Q5boy6fwxKRcBX9m60e/W9sQfqwmqV4Km6bKoGL7YWwXe8Qn
TctvaYklAfy/niuyZyY6fpMSsIQjp5XySsvfvQbR3EgbOh54NelmlcE8sUNCZA79
XTyA0GksfcMYRcRP18GM8uH9YAWB5giwhDfIxUd/6tSNRRCvUwiWFX+xRELWlds1
9W/X642S2JS2qcfla9Y4ESSYkn2AOqyvz3Wkc4j2nziKLVSxRtPbU7F+SO60ODMN
QI7Tko7SUbF1zoe3FfahfXsVjNECu3FrwmEvHBkjlJer9hHFsZyO+uoYfZLH2Kdj
mY6M372bFuYWLdXId496I/Mgg6LLpfrS3eOfMpUijGJmVYZvjjPrcCcol6DlPuCN
5FBCIL477winrV+o8UnTGy0sI5jxgl3xJuxsBoYLU3GWNv1DabOYfQy8GKNF38b6
2LiJLzWUUZeIEuCz6KvId6LK20Dm9uYoLkn3Zbs2MUefWZOyQDwUoTmr3zlZfWZX
+Q3U53IUxOM1JX8OVMgk2BcJq1gEL4LYBxGQHtSW/EV0+a5pQ4g97dtIQMYv7A7q
wcfHcDNzzAFIhqrdq8LQcW+dmC1FIgIiTb85pgdvzft2iNT36WKXjVehiDpjB0EE
J48my58oPjB3OZf6RTHwtPO+hXn3Mk0Pb0kbl2ggKZ0fjrds2954y1Ub9205PTJb
tlWiPZTzip4+kT4iLWIzArh30vrmrWPw2s32VaIibvN/LaSGcbL7EIIUJMKtdI0d
SxSjxFJxd2K1xJLgByucDIygghSckUD7RrQgzE92SUPXQx3JpmwyF8OvjAJ6Ve1x
nP8uWCnfJeLRvyZ47elcW7BKDuXPB1STJaBH2Nd2ontrve4ZSuGMwQxx3MLRWm4j
dPHaiP/rG0XOFexcxBQinaVXyENE4pgfuBiSG0SZyMBuYj4tt1cz4iRSJp08sFjc
25GVL1Yff6EC4WL5+kpZKTywpfGWmb9ovyPg9M15wNG1IUkn4bhLne8YnSUgJK0v
EJCU2Gal8IbbpnY2hqSfZViN9XNx8sVW1n2Q5nxltSmLdvo/3h+26ZkKc7SFZ8IH
CM3sC7b9xsnKsq7/JT+K2MGWIynEE8WO1ZrCKRhvZVcK4SKhLDwu9NKeWtSwPvID
a5euV/PpG404yzoWeHlda2jyUC1DCAUvMt1UoNtarFVt6KNLaY+9sGJ1G10gZiiB
JocijJd5ULh0bjo/abCuCPetC3U9pPOhh6WsuMgPZWBVF4G2FXJH4GWlMUAppmU0
Y7kKnBRNGiv69L/Ac3wmjILWsf0TlhgMu1n1qncyjTE197P5451gmC0MLZuTC9OZ
CLY+Od+ajEcbRgabvYp2n9Q48a+fVzLBV3JIl0zgNSw2rkhXNmeX/es5AZXnH1Ek
ypKSSJrIRCxO5Kbrt3PFFEMFf9ObVhkdFQZlcj5lK6Rym20lrrvt2C5VaRViRMb6
Q29HB8Kr0hmyovPX7jZvZc4H/SGW0lpV3Dt1bje8bZ2LRwvAlMu5oRl7ucnlv7WG
g1aYX4hg1CwFZxUBNahy1xgPDONRRwXl5PSVcrp0xNTR90W5QIfXJYyQvvrmZoUz
v5LQ+nef9BdOAcyWz5beqqnav5aWiCWam9qOPLgjlOVnlfahGGEDdO3H3+rSoe3d
S4enHWlIxGjeLWWviQs+wbiPdinIoGStiEck6zONccv+IiWXPFLDDi+EL/yp9X8k
6dJjkMf+lUzvnbNapk9xBa3UB4zQSJx27/D+L1EsxWRMfGtavssFkuXTpR3onTOA
3DYks13XMJGr5bUwf/o5EYKofz0O5swbs9N6+TefkVhvfdoJtvtWDUSc+imOJz9S
q3yHVbP79sW1LQ06s5yq39FiKbSkSQClU1nfgS0DKwiH38EQTIaXBcOSj7dQZKEX
k3LEpQZajXnYPNaAVoutRm7lRMJHZyr32ALUlhgllMvk8ca7YpVD84wiuAETXxrp
VbSE2CTTG6cvBJLyq3Wfg5KrauYbo/j/syYBs5NN1I/hc/vJ544xu0IsvlWNwTIp
OwCWBJ3IaWmOMBscQXWfw1ygoGrs9xNpmW6bKzw9xKh4dWS8lT7FyJeZHC4oHqOI
R7SHvVq7xLE9j5mR1gIq+HRZwsZFTmOQjluU504YpCztCFOKCWyyYztu2PhVT1zD
0BA0l4WRytTnpJHjr8i77dWoft40UASKLqp2ibkv7LR78cVqd8Br1+iMKj6r/kli
5bp2Qlgf9Vsg2C0BNuQPKx/gZycSexAc5+dq2kbj2h8Ke97tgDQ/TRmv9QRZL9we
cBNa5ksquUlMl8hZIP+uR+Z5lf8MT1XDEU4BW7wPhKJ2kf0iQyi+NmGZvxXZqCIj
oz+hs7XjKtGRXT6sSrfJLR776+XP8+Ie3bpURjma64dgh29ETp1fLCA4R52H4jzo
TbUoSkkJWZKS/0gNgZTOnWRy5p+Z/1w7IP3R3ytW07f9GbQD1B7IE9LlUlXh8KNf
pvXBgLQErA016s7dm/0Cf/4kFhUzIMAAf+SzI9krsPqvgHe4E1aNpXk5arO1bdZD
3qkUYTxvCFFSptVeZjGc7HTC5b90JwNmBi8IPRed2F15M+PtJSM6oVfdpttA7BKW
DTO7CMcwU/I859764j5oLoheEl8UNnpJ8xmCXPZkstBI5iqlLm+ep7ckZs/pzd4z
+R7vKqsA6QhH9QY3Eb0hBL9B2r4VJ/HJr1hsUftmpAyfzGH/hfq26K37OeYGByYh
gFbX5PsC14lg0Ex+2avKxgexTlumVr1PQOG/b/IkSwpCFVBD3ujrFXhaTyRRLBxw
YNSHkFTiq+sf9fVX+Tbxo15LTE5NEz6JJk97J//kKxl4VIDcv+ITdTjHHN89OC/C
mTKdXgfKyOk6nhjj84U9ef3lvdZK4tUx4gvyqZJdDKFHE7Klz5Dx12YpKiJTOdEj
EJcfhVtUpwUoEMxU8QGnVk425mYk7epoNibkEfe7/wFK59/Y7ik6rTjZhvAJvpjg
qBGTbg/zyGV2DEGrt3Emw/MprThJ6lnGNTDbcuZBFZU4MXXuaFf2xNs40WhXZ5Am
BkEr0527p9dXayaMc/icFcuglJg/ZWzbbBb4ijpb2FjSl+HIoP89NMxNaq6sBadK
rfmuc189HsP8Si3ew8S8sB8yqtIKklOZj6wNZtkPOzuI7Z3p8TDeqT/fnrrNcozk
JhSxtdprn6nW0kcoxISDaU37bymhQxpXb7vCETr0HgqQgCdKiQ7+88QmkUxjjIQF
BwA4RED82OpwtyP5VUzURXaurh85vznz913jZg7kBgVV0C+N9FS8nMiXz6vb6wMJ
BwO5EO72ND2TjfW47H9a4o/mORcq0hJkUijQM/Em17o5jOPR0CN4tVdzwDbeCVoO
gZz2F77eF/6zAqmoA3LgIu8m/bSZ1pYd/n26BZtFxdm8S8RGlF5U4aq9bzuu/m2q
HzeZ+AVA09RyDG4R+gsfbfwVNDz4djF7eCi3TkWR4W8ZVtcllNgS9NB1nz2AIPDZ
gL4D3zjMqRIZQT/hUlO9VRGWWOg946n4N3rhHzwApfccwocPgO7cEi5sHVJRCW9C
myt14lXlsBIgr0F+OeM4UtNIk8LPunlTIvosUHLhIIvFLvJB1RC/l8/Y3SRvHDVJ
bk7JnYwjvdqxtwN+3tkJD3jrPhDa6E16KZTQU/VN6kcRBOrE04FNHvornhDKfzs2
cu09fjrPDxJOs0fGbTDRCuhxx3R9iBLo+tMVMm+eNc76Pa0WMfsNCFS2Xm1nTo4Q
9wBCrDG92oA2gxkIBAcdIhqq4/apPv8Sx2WQF1HKyQwezT3/kgA/wXgJKwYTdRjT
TepA094M+bVH/biIVZd3Rv6okDLnVUbpIzK/G5rC7a6RFaa8FQ0AZCppuOaMuPIq
lhfx8MwQY5E/cTbT9zcDnIq3pYTf222phMV7IBOXwHIGbrkbxFKQQSs97EuV2ZiW
XKyTIKkm/N8seqi/+XR6eyLCZyjlwR8g1uZbYHXHWEOvxjG4xBkroF/a6ZOqfjXQ
MnNVuxJQmr93/RYdn0ZexPBuV+nve9Qivhcjww4MXRAe2IwREGyYa/DCq62Fm8SR
/JY7JvEJjD5KB1vOVGVc35z+IxzQodk0guetGAux58oSA0LtDZ3oP7YUnyl3twSB
ehKXXEnOYLEQBITPQF7OWC3azsgMHQC9roeo2k/QmwVcbpEWhk68Fw+zc9ZvD4fZ
pWIU7Z8EjkRA4QbkSWl3inEseeRhw4a5uZmh+qBvgWrBlQKIPAqXxRd7lpp4/sGD
zropgdY+qU7LvfHCS0xhXJ6CoJxA3QDKaKKeBGi5hf4dtO2rZhujg0trqdHVebBC
la2UgbyJcgU3fGllOp8Qz0Hp4XRDRaNk3b+jRR2ae+NThoT9KbAaOLO2O7f0+jYS
kdiYIyqykcNda6L9Ssn9fm60NOgzgeEOhuFzgVQmGRPKpXxK/ibGHo0AZnv2JpUE
HBbWQVyjqcCYluSXDSG7eiBwYycvlIkfxOmFKYSYheDJ4jdkf3sSkaDo9SRz5VvN
LY/aLLNvRh6sbwHIHomRyGk0Tqo4ulRyexn3IvPukOvaAWDwZwMfdBx3KRjhWFru
N2VfwnjjzCEcv7tm86YDEKQhvFXMsw+VC+LQwddCgcEn8gVxfoEY4CV3QYAvjYNu
E6fSB5BHO3nUaze9rBuM10YCUijY8pxfARZzU7IU6oLmTG1nBtyVx6M51Km+NK++
0EZqdCbb0zr0OHJRnmW9BpbhY9q1Z14lmPleQHJ55hhtHOoQ9LGrosNZpDdC8jCt
tK/QKWDDOudO4zBiT2O0jyClP2ODVaXHm3Z1U9gYmy5+y+ORWKns9hj/M0Y1mKVi
ZxLbpJ6Mr1e/k/uhI7OR0itmSnyO2Wp6bZydzTLZ4/XTFZ7OSRDRXxy5gi2tOV34
EVjgrGc4z7dwi9L9KmyDmMQuP0v9hNMxwUoV5x7P/x4KtjhPhGLBNkBfBsgelbdc
QjIDavwTOEn8jWoKTBei131xDtbf4M6yxpSTBCY5mf+hJmZ41rJqR2dgDSBhr5xD
EbMC/gSAqD1kKbBJdqZvWqMoyjSIQi6m01eiXDcH0ilK4ALhlj90wA6WYdYjWmu3
GkL25EFUJPDW3VdLFwQLaWK8tDM/hdQDwYloX/IEJF7HeqE29hs70QM2CuRODPSy
M1A6v0k+OBD0qWWMtDoX/ROEcKVe2GdllkQgR6OSfT0zEaVlG05MHPwrjrPmBo9N
yXr2iumsPInLdfwWplFVEUldlyNu7w72VhCeilDJRfgNcFcu414/1g5K75GiJeJN
x+Lc8O69N0nxUob+jdoJiWtgdsqoUK9efMFEqHRnkDwwvODmXA5eMV9zco2OWqss
E/3w4wo0BAv5siM/dyOkebdLZFCst14mCn68C+cnB8OMBHcaSxK7PSfwEj4MZwaW
iuXsww6I5qBB5Cb5341kfL+SkIObUdlVDsnf6q6hMTjjg/qvckDoIWN2mIHYgo/U
HNce8S2zLn3Nyo6N1eIt6+JhkaEAg/6n2pxZerdEZApyhq5t7kA1w5oKEqA3SpaP
N0KFa/wLQLh223jvCnmSlcA5bp6n76QA8QdSKxKpo+DlEinbFe3dheqZWnPUtS4U
Jz1QhW87FdhXeVpaenjNbB/HHlVzQE8F6zBXbf2dBKiv8jooaoJdzYuybWdCKdrc
Wwe0Rbi3l0KdVggINNvGONL7GywjuwBUp+236JtaYFkOfdyMzOWtrnu+6UvKM1Hs
bF/WV5VOBdKIp7nyd+zT2kWzyNGYjHfxYkuLpPLwbBz1sAp6YO10lYypi1Hxknnm
uY0xiiJypesNu87LcGuMkrFjoSWPS1VKv3pdRTiS2F/0YIKtY9nCWl8/zvcFqNCc
LdbTmT2v2ERsjrY0wYzwHEYcGQAF7nhHun0DpxpI8XsPXM/+wvaGpXWCq49PpNLX
9ImpD2ruJ5AC8cgFaqrUElBGa7xb8IfG6nngOgU9mw+PCKoPcfvVDn5ezfLLPSQZ
tX67sIZ8L0jg520ON5qI6EqBWf6FM/5df99m7qiicl+HBRau+RvcciuOuLoKi+TR
5ofhIDXgXsoEVDZXp1N/DT/i960yqzE4JZMDmaHlz3Y6txRcVIasS0+zYjU+qjrk
R7cr0iDNTuak1UfV/6FGsvphoPsurSDEmGfsXZG22WLerkbVcdS9XJ/K0wRDWrZJ
vnzcIcbgVPDCtXKQn3vy2aMoI6SyiV62M/9qOh9Sn6d+vgqOf62fONrt2pkWd/ij
U9gM53WXlayQxBcTQ17O+MkuJiErVkAMYS4ibfp8ldw2gFIoQeeAXp8DGV+2IWJE
aWnpW1SszAQerCN2TGTro3LVBCh1rxuOXF6EcJKnqkN6VFr7lZLOA7EiCtt5MAVT
uCOi+9T1YTOKIqqgelPnRdGGIvW+JrFrsdaHAgBg40kspY//gKAWHak33Qm7Co5I
Aat1NzoDBVfONC0ON0dRjxbUrSaxOM0prPm/yD3EzmTpAOJMvvjzhzJgXIzoHuP5
YlBWbTN9LVplOBCJ/q3d3EL1DJvReJNOWXQzuNWLnYQyR5q+Jl2k9hn9VIGts3Bz
gaSNlt35p8b6ozr108DXkYIwZTxj35DmtiwXWOZDaH1pHfZYUcwxBJvVXL6eJ+Sb
klQYgqAUzTwzwGddMmxbbnODHZlwWmKj+i+UJ6eTfSe3/lLrw8gT7gV/0i3ebuH2
XmZd6axmiBYddetw/w5srtGE+wCiHmG+TDz/XTdGPtdONU1HtrZoctr+AUjX2zCx
8cR1SRro1V3KMT8LpL8xnNQZOUxOzk7ak5ss+dhJVV5x0c+eSv79qfNdIhQ2TuZp
0FXAbX4CVWU4uwSHqS/30qB6DH4iUVglFrdX47i6J0C9xDifENpEKmMxT/D4qUkT
JEkfM7dFEhXB4/Xq0/HZ6t3ymmUx6Qc4t8sqjImZOSDk3Mv3l5Ez4/2NVNc+BhUc
EgUba803kXZ/ick6fUeB5+UD0SJeR6diIeq/c/55qO9OEuKqWeBvq7vbwSUy5U2f
ekis/LlqPfeEYPd/pTgSAyPxZUA/+h2BX8UDlUFlMyi9j6N2jV8eh2CYH0L+6poO
cva6nozJxtFJQDFufpEQ2QnxHc4lbeMQcjjkybiIGCSj4kKUWbJT1TFK1yri9DBP
XiXtw2BxepKd/ak0i8g0OFcIi+uUAV5ZpqAiT6r/YCQSBgVynjR8j/zzMrlgEYGz
WdTKoddQD0MGi5NY4jT/WQdPJibP/+iiFT1SthTTWnI3m9WygxapcDpaJkqrKDSF
+xVRS82hY4sOUppPUxmsEPEQepJ785Y1CTY4mEaDoYSTkO56Z5Es8NaKbFnosP/d
NZrr7oEowtTYEl4NSNvw4XZXhHpE7EdYb3HY5Vlgnv1bKiIfXgIS8gM3GTfsqzlO
w2urqOVe9cbdORate46/8j5RJ3x+Sx9cFMGxGVZSSuphqNg3iBizw8suB0c/TeCk
vkDhVYG0GLdlwQSADbGuATrbPo0VzUsBoIRYfuEPjpGRgDzF7XQhn+wYE3Q8MxRC
VG2FV2xdsJDrM+q5N/+zMuk635F4G28SugP8tI1rHCn1TJaXClvuPzjaRNmGsYMk
dMfIFk97bra6EBz3gcO5Da+vZdkvkF3BCq4jXZeDGYK0W2ZWDh+XxH1ODHORkXMj
tlB2nFK+UB+wcleezizB8fqvhILe6HqhZtIafsnsQxD5k+0QuUAtNsruGSvhcm2B
XAVkOHIenbz7euArb6mczWVyQlZqwzxj2vkZ4XqPzoyyk6obUY86gkPExiW1On6e
4F6VpJupKt7EgpEHU3JCSNZixM6XTmLXiM2pHvqcP6P43wtC5q+Bf9r7xCk8Qa9s
qrkDpOeSEi2BH3MhyzggtLjiKXO6ax09u2c+TSQ20+Cbw0ol7cwxAzr9+JBFwyI3
HE2/KUDMchrEPxLORwuq+Vbr/rbm6pXEDIO62qfRZ9fEC9oVu1SN08u4G8bT9XIg
boOhVzex9S/2trAvYSfCAgt3o875BUOZVeUW9qwhkwCGlGfkkSj8j+cXifOKRpIx
LUqDWE+MFmdrSJ2URHu7m+AqLJ2yQjE9Rbu16uA578Wk0rAUW/INAzyRGCrtCCDw
2w+oQ5gHypJW6naWpQdW36C5PwY0B0r2e46SuBja3T0am8fEf4Psl+RJCgdgBeon
jNOJqSLIVkXFQugirzzj8DmHs9T+LX3gKhSmSIoNNu2iWGCJIeH+gJp3fOZK931W
JEckWOaBsWA05/ajiSsL9t8bnwgcolqTopNOqh+HOiVrVKZcojx6u80Q1DJ57ViD
GjZMD1bAXzjR6oGLgSgDLXWrZHQLxet5KLJt7msUuuf/cyrwGjcBC2b3msUFmjJ2
XIRntQnLTo0QjpkygMUwgNwIeMFLvi2ghCaozntwWd8A90g/IZWXgOGw/AECFCtO
y4GnLir8+y73vqgJ0KzR8NgfFqivoDxS6/Zpys8vTdYRet7buYN8OEAaWySl4CrB
EG7DZu1McuPPir1yS8HT4o6HZTblcbsPdlnSJXzqffKtsKmB9+L6zZHHN2dlVCW+
Lpun+ysFjFicl+4jOmos5wgb9dGz2L+y2AiHae/TOGqfyb+V+5doPwI9ZcvG5dL2
pLI90S24uGSIs9mafHiTKuQqpw3TFwVKDYTh7mf1AcfHG+o0H1A06aPWzMSEcufq
zAS27EaaZYG2A4CJyH/R6IUZ1FpT5hI7nayL3593HHpOTO0jE7TYvW5NQeGOjRdm
e9vVoPbU4kT+VZKuT8Z6fPKCHU1dAODRcEUUfk7SnnWpRAMtJBd7O0HBetlwhbhT
u5FUGatR689B+CWkCNY/np2zU32j1BL2o5j5lARKgvpWQA24WXADTqWTphxasP6f
/5IYZp5M/9q3wRPwm8Obf+H5/xWSkxGPyqjbnbDOBq9GEQQLPfpzxb/MtIGOJ27S
jDh/AlcJlVLM1I5PldGU2glg35E2qaVKQP0nPGPXvSFP3q5JlPVlp5vNFwdpmYKO
h+aVhCYazPvvOgqTejmBm3mNaSVwgU4WnSe7tzak3ZMGP93Q+chIUi6FvD7uR9lE
Bi+PLdYYNpX+s1Ija0YSLiWg+hpWj3cKW8T5pPfZ3VKCG/QQHKP0PIsyxFthWvZi
CuxBOChaWPPoASskP6sYESyQIkseroro7BwKWTpNnru4+P6HPoAkRQVED+Otx6Rb
EP+NMPardhz+zkncYeaJH1zoyeHfBZRomazo7DAocnwNCkT6VPHn/9YbY0EexxSE
1OrMHYUa4abxXUIhH7hVZu7dLqxf+7uyNDL9H0AFRzWRf9svPmAZx6v7TKfMa+FX
eHbubVqSnfBA0oQHVefGWqlLTgWYS+MaIaWEn7ODWTyPdOCMnf+a/xexMysRYnOn
ob8ptMws5EddAM9OC3WkrtxG8n9Ja0p0zwARub3aeQEenIeowdIfWtjGF0IpRo9B
+lRzG3nnTqcjW8rnUaXD3ZvSzMx5HqMLQwPD8UL3uCNCDxICJDKfFbnGxJwDSnzC
UXsR8bb4KJuWI6uqHQ9Eh4fVAmiUt8AQhtkP4wwjvY2vkMfijzfa1mFekYml9fKk
UqCkUYtBLZfBH710mitSRTsZm5fuQ23TtwjPp98+wNuKf4JGJFK9y7zrx6Pgrb1Q
bSWYyejRSOd5rVvUi8t0+SG1lUlJsBF0vZOHz9zLAUfbwv/DmdGOo5WlxJunMjSp
VD3eIzO8hvBcAXgNC6mqjyhe9ePjDQuqwZJ2ZMvt7M0QA1OHyHOP0S57HpVD+Urq
S14ozQRxr4Lg33oKsd1A0GKQ6BIANAyV4mbGvYlDy1wO4Qwfzb3Ok/JqzM86VSub
2NmE4Gz/Mnyns+DM+akx89WAw56M+kYw7rrx4oTfJZjAFLtUM+HZalT+zPLtWipL
KklMmFY2PmDbANjjtyAQAh5J3gEWVyZoG4HinQ1+rQfRFfa6tWxQLw/8Yld787L+
9S7CtthCD6mIfdEu1MdmtlpexVd+2Qu5WHMO8DJVYG4kM0HDsTjQPdJfsTPLKPGD
lmM0EGnxTTofhkuz2kPrZPsBgLlWXOBfN3B9IdaVcXvmIqRs2txopcnGnDW+UQML
8sCypoNa/p2i3SON1AwU8cakg1hmTioH75iS3xv+zo+tOCAnO32Zpf6Jo0DuKfd8
/MxQSMyd8ZBdHSWRotY1VaCzI8qcZdKqac3dJjWaBR9ArA2jJhvhHpbyltLjrVwn
o55/rZGkNNYZI4Yy1pKtN4Gzks1QfjojZkKn3PYNmQNdcFMQ4gN9RS2kdIlzdy7H
mqL1Ssi2Tn2QSvyzeiFhVZivECxOli02bhEzGyS3hnMyzUYK3HchplQSvXNm/TJR
+0TGHQokV+UCCLLIK48FacosdH/SqDOxYyguDItFLFH7ZqNkaXrr5NuNupoymcSy
T5+5tdlSMMr3ilhyuERsGyVdGZl6I5kPDglC8VmRSV9i69khYIIEahfAkJuA4L0F
65hZ6dLkj82Ao3KoTtG9qIsHlSXldVlYhe/0hcKqphLqIhsAZuiqCXb0g7bg7Mw9
YnCvhV6SAfUfGEOQRO+FD2iKCF6/CpOVkE9LVI3DJ147KRzkbH7mDf5DgUMF+Cnx
O/ICVvQlLNMrnMo3YKx5JAmk8MFd3NZ7BiTgyhgDsb/qcge6x5ipU9K4E2GfNIqP
wWnZzUy7GGkT5Un5vMCgnZTiJ9ureYxfBphHViov+Q6If0o3/vV8dEoHprf+nGb2
Z8C5V0tzm9cxb4GoMzuM56DHy06fojLblDjFVRVb46Lsd6btKy0E9swy2evsYrZ4
U1i7VcCuLOKOvZ5ia1ToZ2F+CNK60Uxmb/Y/DoCHnSIsPjEPuKNQ0QSSQ8G1ptki
vD/SM6TgVBW/TpmeV+V+LzUggSlnRbGPP4RjtsuyoLr+QtYwov2geTymc0O5lrGD
Wn4ztLm/7iucWk7OUT9yiAYgiDv6XuDSMNLSt65qXaNVywOs234bABEN2TSG2soQ
6gRNH+/oGFQGA1OsrBlkHoeE2ld13PCKA0kYvz6F5FeA/S4RQNZvOJ1zx5BuNY/I
Ok1PFbjsBmuRqslcu8QtC/nP1JC7Bi/IOdBgDM3z7TuQWkso/fKUM+Z9P9iykPHP
GsIXql5rsAWpo0J4OCwEFcXZPfZqdEANsNnGwwkqvIcw3m9+pvMfKZyYt5aqt5Vs
Z07aCFu6gKhy0zz2WuX5ETT9h7Rg6wZHEPUYJNAfIvQDKUN5OzflaeQmBReVXobN
Nt0ZS65Vof0JI+wJzLuXViGdAJN5SRR5+dbIgs18gz8mVTtQu3jaGgnFWB6Gd2Wx
6F514UNbIVofZ099u/pjQC03v81m4XatE61xhCM106xicj9xelK+gHCFQUoAoN91
BsG4cVs2JC9VEJu8jAr9Gip7JknaWzbr5E3vZr37CEz4woQmZAdVIvcbNPP9wwx/
mBayy9f3DqCGlhEaWyTyxLClebWzvaU+wDFTiU1MLF/88sZZs7y8hF5+LXawxlqd
jTwJ7oiRJGYTIMsUjvyBLyySMTWUkniLlgLZpwYa76rALKVK0dpXMe8eQXtqT2ce
kT6Ce8qmtR7OpM6RqU1OwMgcJu3SbNxPwwMNxMjQhAWxmw5anyO/WdU9tkz9/fiM
IY3qb19rQij1EGl/P49GIXtY8bdlkSSi/zdquE5VqCZAOZL1y37sUDxfp8ewCa6c
eFeI3uBSLPfJaYNSgl/+JGG5XmHJpRKMzem6KhKzb07V8I8KoHIz4QsVTg0wzbHX
D8XWDny1wN6UPDKbY3QbBGulihwqe0nthNsldk5VDJFWa8KrsJvpmHiSI2qgKLdm
+Z4rnYMcDNCDN+VLtiJPcfBurZg9MIO1YirMJ5Yzs7OJYu8w3V5NEH2YbrLYTb5h
SIojzZjygutGqZcAKul0OaP1a8aAWoi+rmtQ93TszntcW/yAafNY51XI/Vs8E5lZ
amywfEwxgNLJm6paKsXY5C9Yhk8kAU/glKtgMUQwff8=
--pragma protect end_data_block
--pragma protect digest_block
/e6PCXTo52SNO3wftNshjZLn7Ms=
--pragma protect end_digest_block
--pragma protect end_protected
