-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
xJL34mYwDdJewl/KEOOq2ZwfRQDiKDnY8DVgXNBmV73L9nIZ98n+qXlhkyuXXi9q
/a14A3Md0EgpwYu9/6vJY/iMablJgXH+6qZQVAfby+Ze7rCFLPB9Q9UztIPCdRQt
OD06XCmtYsrnzMpvjAew1CNat8E06MJhw8bJ0n/mMSk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5056)
`protect data_block
2ocq/r3CnG/Ho7AuMh9Mz9pLBQIIDq3DW9b0bqRprWMg6vQ1fmuKZ0kq98M6f722
elf8OI9+1PghvaJBwdTQHryEan4JhGF6B38BhY2Z+1rJozwkrKk6i+/zGOzGtoq2
HeYv6KYMtBbMxpX72zKICDhSRPJevTWfvoBpSeSnFMOiUYvrttqKaRWD6WAoDKID
iDGJH/NFsAs0kcUMEUGiYINNVF37FZ+aI80UKxs90uwW/b3ypXcTq4sQy7Sg47SB
4X48w08N7I7I2DKzGZUJL5zUe1I01yGHKE5UQKp+ra1qpNQp+DQyGP236qrCTVUH
ivoTmQMVyhGnk+KmoCkPtHe3Zph8BYLhXl0Tpr/7so9bAxYUj+nkqKu7mXe6D2rs
X+hWARPoTcU5npMr7kEo7YAi953lzx13g/okfjk9wkdX6Fwe9e/bQnHARQDWmR+L
dw7+tBLMujiCm/amWSqc4g6G7aLE/PAbKluWQ00wNkGIYq/i4QSMCRdmkfrnM7mQ
BtTXSnkFnc1PXy6Igl2V7tJ11RBQlecdY4hWsXsG5WiepIIbxoKauW9ut0vPJjFC
kvY9pPKAKaiO6don8qq6DTaQoJJC8EvAO5xreLsvdg1DjWOJ7LfF4LTefVHgd82U
v9rIBWm5htEnXA79zNM53DGZJ0eLzWwe9pm9eqUejP7YICfEyd0HXCiU34/v2x1m
w9tFPzxt53QWH0ZnVSJ1hpSHXFu+51/0u/BhArFHz0XBIw711xqzQySew/+GCAMq
6Yd94GOIlPOT7OwQpQ2bY/zBiUJ8QLHKYqhdw0hGpD/iosgwWlPykLtOWUWXF+mp
3GhFawHWj3XNAlZS/3eMexplCPTbJskwijz9OzeZ666CJNYva5iSz/GtVCIiWNA9
ABYo4uCrT7fvRfu39iv+OCMlCXxa3UUjtnYMQdB6olNPtWRV+pb9RLsfjdDpOSvV
79CO12FykDMucgbAXAt45oIcfp+ODL7FL6F/C7MoaPB/BkcwGxjtlWQbobFViDSO
A5qkyi+6uL0/BTF5fFMF+w7v25QEfeIgNyKQUeysBIFa8oNo5/6P6HASkD2kbzQU
pM/ullHUfujOMKED+6WLM8e/oq8IwUgWnjN/Uj7kTFLiWk0V5iK4nicAqtFNBPRm
k+/6O7NPKnOXdWuqsaIkoKudLKmI3ADnnYdozZrxsvMrh+yOup/H4pc0od4xkWpM
30P+FcvXoSDrLm3XpLftiR1Qv8ixELmKNcc1W2LOxI4YvPS1qNFqb8x5+a8NB7pd
/Ocb5dwdCPWuvHkWRp8X400vSIspsj38RBLE5Wl8nphGx/CUb52x+zSGmUzyOkdW
1zF/oWf4P8+bacWSL1SDaf+2ITKh7l46W2sNXX5AwjcoJ7rXHkKKFvpGLL/769/N
Za42GDjktevxFtAnsX/lGN7N3xgQnYCjxPwebyOAA0Vd5eJPJrReEy2g1tQ2IaHn
I/LjGpCmqGudFuMdV1ntL0QWXyxoATauu5uC/mG3bdjKp3dzw39poWooBsjhlle4
qHNfNFCrgxspOQY9F6cGqu6qbWjssPtO1brpLKJ3NrvjPtdweF60qA9XK8B+QU4T
LOTJlCBfNAOXoINLu5rF/ZCcfCxLqofJCGnQyq7nXuVfpwdq4VsM4MS2RIlduC6t
qIYCG+n7osiFzo+22/tMI80tgOYYnZdvl/Jgg7Z/dBLB+sZWMPZ5RzMzvG7AUZJc
UHE+zdDVD3Fq5aP0D+HhboGSu7eEjBI3ZY91pIN23q2BOPOfIM46eCDkePbZo8Zs
L9ppx/ojEWkIJvSwOQjt/1PZo33LQ+MspQP3ObVY9hlsUBuiIAOuOy616Q2xUfmE
4/Yz4Ao8r+P5pE2lJjqjT6a+FwY5Q4+JX5uzgQpn9Fd519QLank8Y4lCznGvpk6x
uT/7IEES56tyXRLEUW7DlCDMO4Y3Hd1lj1Mt5uENngs2BOdn8vO5dta0NB0ThrqD
0dzSMZH8zHqH0vI2D0Bg5jL/4K1uPEKCMqJbmMfHna6rMpR7+ZI6lHytAKc1w8S9
be04pxVvpNeoCjB0va08+lte+lJ2GSZ/f71B+FZNCXi0flt2JMY5K+ED+76XAAjc
luQJGypnEG/iRUpJ7mr/g4Gk+3gn0s6xnKw9xa4M9+e8dWcLY0nvgstfeTtqJ9S6
q5fWc5KXOnVub5PZNbbVWL6t8R+keI+mSIOs1+3tKXxsw93VmzIjjEbxG/hqCLJ3
nzDc+SErrCs3eaAOXNs2XepJuwUW0z3YH5IRDLFxewnQbDm94P2LF3LHarfJgpjk
fYlBezqFnLRHw+7VJ6udZIq/Zr3oOnJHIs0hiktiqKJtBo+hsY5QzyG34kppSeO3
2sdEqEhF6IcP3grc+m1xJituQPNLL1fsuYu0OME6MOzp8EVGtxKsBSNcJ9LMlxKy
5nmRz+RmpN/WsC1gYxhOU2uHikqoLte2YbKPvfJ8lNShtqQzYvLw8S18lGJDFv6t
x2AsLx1C9eEMss4S4l8oae99Y544IpDf2HVt8gy53uHhYSFZG6+qBUxq4vkkv9pl
sKblogehidxKSTkIQRdP+FD2X/IztpdFFdSlXaLctWu1uH5fMUBGVez0QUSh/APa
vnOEgtge4qFn7QIhpvFinysXOguhRKy9aB18boK2D6215TM/mDVZZyF1JebwiBfo
fJ+4H/NBNc4VXaM05ADdCjByY0j3g/VyyDu8u8JolExqkTzHnnougVPJ1nHBxZDv
JnLIP0TnYV0cGJN74L75P78egyplodQfyLmyhpJe2y1aoTBaeneNlP1I5Q9WnRXS
xqshm5IxRx210VdmQPYxjWYSV51pQBK9S70uOqNHULRufOfFedwU6xQ2MAslGrlx
EsTnPNNEJO4xuHLpeZtvVvRDz6pqqSr0L2B49NzmgGV6LRbYhGnw/z9k8vPF0LA8
RaYPJ1a49MSSvWW/0QEqJMp4nQV+mpoxmD4yC6Zd74f15TA1RX02pc5ZmGIVUa0L
RrkiEo7lr2FesdLsORo+c1lJJgi+a6QNg0kziBfMUSqO7UxG6mHv54HL9Hlebqfo
DVIjJSMPfk6aYWvrQ4XTT87iwUVvaqbSIROqx3ls1nVepsz2F7236+tCZSXp4okr
07wfFsXTiM8ROclIXn0tlkShdO/C3kkkEnp98eD2pI/H85eC6xwnXnOhS2d2Rmm7
j3g9SabT28gYSnGZHuVTZEz1tt2p6P3tWaIIMo8AZDKr9sx6ylDvAwM6vgLymO6F
0t4My0PGVgxaLk8w0caNsTiqxJqm4LtK9XYe5m+9mAGp4FLoroinwPpgfSJDUfCS
dwip3YIA+22o/vOyf6zI2vDwwzKdK+76cs67l0KqLCmFJ63XJs43P2VeBsiWyfV1
TQ8ZLKARr4QAmV6JupOLs4iZayrOpQ/4OzbAG6hE2R4gl2lg1Me+Bsq8JTCvhxh6
+jj45XxzWN2jDHjg7dziM8ObZYzzVanva469gfyslPxfGfOP8/i59/Um576sh1jR
tOHU8omS/Hz0+G8qo5e35fbX0EOnCti0V10w+44XRsu7AvS4UO7wDPa1pFuFvwrm
uShgGiWOMEwIja5hBO8oYWjTi7vnlDsOzmF8A45ytbZPXeINrIbpLqS8lHKh99sM
JlQOScIoFr/QHkHPvctN1Cip2jDYA2HaOQOd8oHpCyYFg2FjQ94JFbYl9dCUBYv5
MrdNzG4EsYRe4fsAJFJ9IaZFyUykAFEAVBgvZ9uoUOjghgycG6ZU1ZzyHb4a7vQ/
0RTaacz84pbwLTWFL/Z8M7f/eXLnk+DXV5Oq7j76tPQEXgoxD5wlic3DaAcX3pPU
YkxTU5K6BjJTK82BBXlcw7vnpNqAX5bXFSbVgcGtEgl7vrbB9UcHKq2/2t6i3ZUL
rI7QiAB1+B9pJS03CY+Oa8bEbUYmAdCh7WKUZFkeETHH+5QbkRKMcYuwzCyxnl9P
xxK4iymJHC2WUqfs6ElCx7TK2vbR4EwSj29jYi1szsWgJx/7dhzSratck0UiFw9/
5Y8YOAqe7NzgHnah5ha3gwTvcvt1U7grzwcMW9DP8bRRVfBkp1KgE32vBfEgbHVQ
MaSE4K6mME/ImufKGir9tCbfEhwOzCdHdz1+o7QbsVfN/3BvNVfKAV7kHEqkdlcA
mKJwPuMF0a4K8za7QEda3GybnMVZoC/6zCj7uCIknHdZdem+JISc/m1qitMoxchs
nZIo14zt8A/ExAzJOubUNL17LWnqq5qtuuwgDFC4mFkdMebU9VZq0GCVwG2G55Na
JxcbGt4KfxKBck5n/TgHz8XzsqVnZLHVA0mpA/x8JQjVTUrb6Y98v9odNyUGN3mD
rjZGXNhQFfmOe44nuSZfeIKIDPRnHHGQ/iHmAovs0haHv821P2xyHf1Y7CLfd77Q
Yn+QEdALkSLwqu/hv2A+tjSO9GWd/K+ln34IDxg2kowrKSw53Hg3nEyB56MMObvt
X1YekkcUAqPLFGRqqolM6bgCkptRc7Sx7hXv8CRFacZcasHubrYvS1hAd7gDFhIJ
B0kwmSu8rTO87ySxBIKYk82kUBMRG8AniEq6X3pyBKzAM0VZA8lDor+E+qte4v0p
7siHjevs675m6JmZSa4SG9CSJnsdOUxWFUFwT1ufo09F8ZIbC8Zi5h7Ib1eECLfe
b6TzcCjuhUhTlWNjYL2k1XnX9VrLWt8nW6ctztR5KDvZVK/14HHbu3h2xFYu+poA
Y5opEtv1o30Ua5wsT7dqh1gSWWti7t2C8AxtiL/BaVXV4UGH3Yvm0n45m3Yzo4Wu
72/QVmHlqa/t+e8BFlFwyqyktY4C+AfDFJwqWvGzf+VJgEH0UPuGygW32B66O9CU
z6noYN/otZDr3RcMwDdD5ErDpwK5NJncqO+iU40XVIUEZTodPMegt3nD19y+SoIF
oDYYrJvxJJWmnrzFohenAyiDRMDPBYOZOAPkiBSbaoYmQE9rW0JjPXBtN95ByTde
+XoNX0OUkUWpFQniSbuWUS1fKjp8wlkuK9yby26JxOMDp56S2wc/7+QAJFTLMG9h
zrBrkdsMQNarx6jTs7uSwecN/HYyH1XdwjVxa4WGyqtfZSckAZjY70767qc12WT2
IISrf+W/PNM7D9Y8rV94TTI8fJBYUlNYRk8H0zz0Wk2X6vO/H8xqrCJHkZwZByac
3MK0SIlZh40VJWL4x2AOuDhJO53PnfeQZV4ViR7VoQQ7m8waOQcOoVPclqvlwL6t
zbJ0tH4yo+4EtlIoNYqqXfTrGsF8B0L2miwmJDzNXDDYsjG+n7rgVEIHQ5YzT7Sb
uDFMce7+MqBB7sugxcXhHdBAlz68aHX3pTltywqrmkWU3lv86sWm2jWDLa9V/S/e
Lqd7QZVD4YubCRhU3PQqBtC9sTfJchvTqV/CDE28zXiHkypxcYPxzphhpo9QW95K
TkP3j3DX+dTdfnyIMRJvVlRqSlMLJLKLdh8K+Os0lOc0iXLECnLWDq+Fuyymf6rj
OZ9f4nmE/DU2VyhBUTTZSHHHBhvrI+s8VtohimTf9NnyaGX5JeqiDi7HGRFt74Vi
hWBF0WVVx3oXbUiu+vfyIPODGKiQTXaH7aEzeThx6qKe7eDPJSB9gnNlg8ysPdUG
XLLySiz2/bH2/pq738FbfGZMP/9njHaF7ANPetZiuuneT26Qju2xodh1NGzbTl9b
DH1D/1H3ddsZrNcxLLb39VnRlIQJYBTCl8reK0kZ6AP0jr48w5WR5MjNdBVg/8xm
CWR7N4DJLsQWrKsMxJDcPkDscl8Hk1QegH5JGDE6838RcWt9cL/VPskT6k3XdbNB
wxhAtLNnxE0wuNdH9VEBHg0/ZVM8Bxy2+YAiAnlcw/8mrM/x0aMDGLBZMtbBE4rs
BUoat0X+R72MY1wqQUY6lS6gUqLJct5tzXknWF8hvFyzbe9s+2I6wH4e8BcaWei3
ktYR8SHM1uLxyX+/8UCT8byLkE1QQ2yYUfz9FaHuZTsfPXMVEm4nCUj/tgiOMHA1
LemPP8eYzBfOVBKaUxSOhojt3nf8dD29pOOYGGl4+JYff6uCitzLVQoZfR7xRG9e
0F77bij6uafEm81F0Y121z9rGRhX4y4BjqyD6hG+CHKaHq/sgHshjJ5SEtj6fGBt
m3vXsHUjiB2K872kk553nDk1pomGxtAaJcCE5hbpwtIPkpFS1ImXGKwuywm4F030
fiAb3KJNXfpds4871+Ogn7u6MqJvknu+c3iJfXpryD4LX8VAZdOKUb3XzkVpeX10
fK5VYJrkKiT2WT/Na2IrvTHkZobaER552K73SfnzIkIkX6CFqOCQxPPi+kmNUakx
HwjRTvdOjDDKX9jPJEsYy2IGwQ5ww5swxtRiQhz/Jcn5Ui9yPOeHnqY7WQm0RQK7
JzZmiN/3EAhvF/wWaYqSaJnnRuBRtFgMXru0ZUmx1SER++OLwbmB6QxxndSE2rvU
TjwrAD20WgkshAHj4BLT/KMKLrSaPABJTlEXuIyVZJJpl8JOh8k405RtPvSaqPhK
enppnkzQI47Am5Z0Uti6Xn+Ij5PzoPT2RWZIt5dTfmCl/8mfK2rzXQdpHS47j3KQ
mUbfc4F/zQecjErkuQwXgzMPP2Bk7/cP3UDZ/qAmyvLr/sG5mlpyOns9PyZ92vFj
VnZRJxXnO1BbbFlf0I1YMiIBb+j2vRgCJYEEgezvgYv2kvwISHS6+AfYLW2RPA00
ehEKCkMpqka6fWiexmzLfg==
`protect end_protected
