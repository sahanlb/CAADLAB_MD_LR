-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
DuQTJv63ChBuL+KAAzGMUoFoR/gaPQMwwilR4eF/BG8hsP4ao7VcT3oUmAcZrJn9
L+Lx+MZGZDFq5fzgSukGB8nhP2Q8bR7jBiroLbgEh6v4P782oFaKEUIbc6HxPPjp
8Qtpl1XmDK/q/Icfv6J3jGdTwiZbkWCoux+unHSvVSU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13568)
`protect data_block
C3xs00+UHfWhzeHXM8QrgGqTfDvqm4LYWgrJX9qfiZ7DVkVjaf5JO5tThS1xhD6I
AT+wbDu6lUH3sdaSIJwuYqI5x7E1TxgZZbM+wVHN5FxdFAL5CedOSIgJ4jYuvKx4
DAHUwHVqlE2HjwIhvAZUJ0boY+kxVwXpwWhFDA3EJZrAildao2kMpvi7OefSKaV5
00u4I2K2eP8bcXq/+RaJKFmS/0NWhsPQ5I1KUUwTh889GN3DDr7Sez8EWDMwnSMN
8T+bPHWlwRNVqT/2khK1BVPxzqUu0FpTw1M4BuSjDP8zoxo/l0rvEOx3FcCWjkxL
BmH4Yf/HktLbr2hZJyCzsjIb4lweHp+X9krgZEJoaLpwcE5r5rgDyZIoPzU3T0k1
f60rGQFP3Udyh7UERjgWRw9708S6pxpWeeKxxmcVh0Nj3G7wILfIBh/ZMJHoAs+m
iA3KFKCHF090e7PpKJzeAc4pZbCNBe/A7bP/VW/7MHOCCPdsdJwwm9jRQd7v7JPr
oTTGzz7eNQys71keaSMBfn4qsZh7VSWIUuq3NGchoN5xWYCdwX+75eVjEu7AGHXe
Al1WU1PMLo1PogjAPlBAFpFGJ9/WbFhlwq/5/SR6gzbGzQ1HYlq83SumZP2ZKzy6
Oj23OE4EUXrxVIs71eJ9/Q+HZerQ3JBttUTMbmTAhwgVl5xiLsKrnJhjU1hVriks
AoWCVTgZYeJgopyNdQiuIIdj81N6LRTobFfTqkWD48eDiZZGhTEDjJe6A1WljKew
fn3k4w1rCWvOSHyalzdxGqtwSFnFDPmNp3RgPIOzxHgKSdItBNWK7JMFV9+9ahG2
anKLFdgr8RDjJ6BlqO7R4U8FYds66/tcAPYyLZkVLFTJYMdpcNww+KgiI1wgfRcB
U54JlVXgabzIjReXIsG7JrH4sL47tEMta4JjY7vDjw3+VOCFg8+rJG4Z/N8jHu/P
nVCwUoz0bKBkEumGpolUZQ9CCLkLAS4tmVx4vtWxLXjp5LuYyT19eTaUM6fxeMTJ
e/sQbZEn2fTRGTezHGtWvzrK1g5m1lw3NNWl81KPkmR451+U1if7h7qqjnxrX9Lp
5sZUSAaO5FqV1h5RzKF32dq/ps5zaCk2Xj0QUPJ4eHOg9pY6NpnvE3YSLSTDIyfe
FQ0O0TMmofaHfoLPBMXK44fnH2pyZnArPaY7BBr7flCe/h1u4BQLEgMjBHFXk3Aj
phfwflCEpcsqSGps3Rjzh6bv8ETp2+pP9pv7grQmETlxtWsfVdi333U/Y0EBbaFW
91rvYOv6Wmr0dU2ueVv/NESJ8LOMKwUmq3XINP+Dkq+7P+Q1Yn1KvMOQZBeKXegO
rpv/CWSGjis54fzdu5MA0d0xc+YOb4ZaHBQrJxdDlcIgpwYjw50W/Qf5PSTp6ez6
mlmcgkLktGwp8wWJuynN+gZXVJIGZpf7Xo34UB/Idlzi1JzABcxELhJmHms//LrC
qfgaGihjkV5FOS5MMw1lZsvzeI371FMRNJBx9qAwB7IVLfdGjifue+sD0B4Vl1lj
1YYXB/NE8wIQH1cxTEYGF4PPOh6DNH3kWMJ2c/hfGZlZt1N5bMSQ1HSHYhqBrKj7
RpGFzc211142Q3OITYNuBPtshC38lvYhCUUzMYK0GbZk4q5ZP/rc07T2+07yTBAy
CRoGwVZmQ2J47jzzR8ZL6hjvLrBWPvAX7ONFkapTdfwjiK/cROjHixGYz3F191/D
H+kBFqt/7pR6giunVPMhbKaM2/vWHIikEK6+yu8jukPXKRKELZj/0F+qgt5dNjeh
1FmcPUf0qL8RBXj9Cn6iwweOIEvv2e8+e47kYShoWWezKmFRuhUtFwPVpo01hht0
S7kliSNr4o/LLod9205Og+Yh+vJzqqJUvUfMhLTozOREckJCyLZ15Rhp3XZa9VQl
/CcWS1HODHDqrVzydgBwLiRxRJscQFSntHs8upK3zePr1PbF2hECTKsb7RSAYIuT
nBNAYkq7FI5pve/KWcfdt7EMNExuAJLtAP8TP5IHhJT4sA5LjKi/4Ygh/dzOwBXH
r9YbqWKhsLpvbWY8Q186oik3iyfM46uyuX7YHZDG/6DvTrs61IY/XwNZZ1Wn6ZVx
pTYina2kkxKd2k15fJp7SqZY62N5zFQka4x0T85lxiE1CoYHJGusOVC4n3PjbVp7
VR9TUpXZeaGOAao7HevTY3ob8WAzos+q7ZmuoEgC4TNbL256HQEoY7fBRCWdIldK
iURk3oZKrpvcTJopLt8v5ed669Axz+ll9DylSBc+3hWbb3Q//Vx/QRNWK1RxECIP
64RYAQmaf19Os9Y50EAZpMnfhIRp52EN1zkEMSftkT0NcFXlu4QptcRyAgZLVKG4
Dr95TGoJi1FniiYn+mf1IL8TESll5PTGeutIP5MiO64b5Kx8fZifsFvqAWp1MuuE
MWhJKjRuoEcZB1ZQFrgNYoFmGYhNCnW7+S/cNrdJOZK2NqkUyeKsg5RlzFcQxi+X
tmUBpjC68Mzf/gr2tIFh968YxVccWoIg3j1JuiBgwmjVSOLLc+0lGzCPLlAYt6e9
rYRjcdX8uuzq11njsM53OMfTqMKLgiLDBGX41boJagD1cVxS1ikgQ8TkfMbH6bfJ
bGIfFLlTJUZAS4VfVQ6YWISXAOqWGdf2LL7JYrAN9eyL4GWcMCmm04WxkC8uWjSA
TBBxXKgQ3EbzGSiTiQ84Ev6CuLlffKNK+WjYOiSIV3JtN91sQNeOAnFVHUqS/BgM
nWE7X2t8qFf5QRlAfLOyURmhiXHSZ0ousjk5AyzRFTohmzk0G53UhtbT6CHZiXfJ
01VYLUsnOHWQTf+Bz1XRTOMvidE3BEfJngYv1jICqwLWnb4Hb+LOfRtTnozjUf/r
cM/xmi70MnwilFzMZsrdPotpzDF/qSEON0TapS5zReS0A/UjBgm6LvLznK1cak47
e3z7sw0H7yGsWnwVwlNgr0Uc16hnC/PbKLqoxpmFT69VCiiZF5GuJiUpW94Mhga+
aP7Xz2fXPPps6wlQLqw8UbtdAIektX+AAExWUASeh7euWZAImETot2wHpPstiJ6T
gPlf1rfQtCBBXijkvM3QnELAOtm0BI/LtUtTaRpymOTr3gLvBBsfx6kJp4t0DHAl
jaalwO0uEr8e+mBd2lHq/y9M5r0s4Yj73Jt607hF6toRFOkWQETf83NeyP6BT+jZ
iY1x6t8Yo+gxGxrj+deo/qJCrEqP+g9hCvh5941IKYVsau7JD9I3wrx9EDmT3+uT
anMQYULrxuQPBq62qtmFoU50MNo1nNLiXDGKtXIHjeRBlHXYiFATln6Im9FGuonW
m5Yx++7WuR6CJudZIBB//2QDMSxxLHrCMKEpdKOclt25nsLTe+/UM0rlydWEO4wd
KN/HGUvuNnOX2xMxSkST3ZUgJ6Cp75kNQmiCM5ALL7j1BZXtl1SQKZyw0eFa8a72
H1VzuaU+POey6bBvHrmZB6x1y7zUB/VtNe9weUu/GcGHUkukimQUcOW73medpQVp
J9AcQVCWUe9z/ShdxIlb8HVdGflnvTVSjE5DEdRjoG8ydy37ASdQDSV+y/lCZZEt
uGDvt4hYP2PpC/faO4cxceLWzeTKRMiOHSRU4AoQDKFmb8VR+glaA20TklFZKzcK
3K48+KyLep2QNT00H3OE3Qp5tZV6Msmw8jpa/7y2gTxXGwIRJq/isD1aRGarEoXE
WpISqqhuEQcpC4eJBt4gS3bbhN8oZz4kP+4uN3u18UXXyXMtY1r47ZlXxkdtcuN8
kVcKCfoF3r2zU+ysfUsS2xiX7bnTbbJjhYC0ZIzmRw3OnTuRUAtWLDE9ch3zxOAP
M/LKQt5PWASA9ZdaUMSZ4kKsrJ8CF7uojIBPmL3MDelfZJg/YxxpBLlC6jKza7ZX
+cT5P+/rITmZS5KwuvBwD8Lq1c5N+JZRri4IEVZkzulophTq++rRUTj+755D6Cmf
j0JzkJySJixuqhh72YHzHmhd+c+M5EyKVY9srF9qf2YVuh/FqnE6TvQEu4ogjtd7
/jJBsF/LpVGM202JHtARUzULXCEgMEXy1+2jDSrKigl+rCrAIQU4TkIswlwGQkeY
nCJ/XNDC75HaX/WFYxOp9AJkWXygUnIykXErnpxg+vNDaCMjb1gf5gKma5vTyexb
g+gRjC5uzhpe+b411s3r8He4IMp2pnin9lpQflxtNtunZ+TgvDalEYZw5E1UzJs1
TnPgKE9gGmOblBrn0Bu5En/RWfH5LnA7pHEd5PpkZISkhesfd8GncwpGcFV0avkC
IUR5syZWZsG84R4v1Cy3MmO8eneplra1mxlbvyCLOvE7ln2BBz1eZbQSqZRTeA5G
eo0L2xbSeRWXk43LLMlFulvLyUm1UJFThJy/BStj9QiJSnxurF/Lpbt/a7cLwXk/
uT6jsJJoJ3WOwyy0TbxAdjI1iza9ergyY/z7yMhMIf5Nsr8Ov8K/5540LF4/a6fA
HFFMGv9r7d8mCMpA3yJjFuPmRIuQ97wCnF5BW0qIG89cihrnhlm6c8OtL7+rlNy9
7FakW6yIkok8866gRIfDABF1iRVXhg4ysJ86+YLXAdvsp9NrhVweIHXoUteQrvfo
W3iVReAMvXb/ERp9N4aOfHDvDONGCvK+1vpuMIzjzQ4Na2DN9vxl+WSGea/fezI7
hYPPKRpkYhwOl+KfUCEebMDzsi2A2dn09kQYZzFLGnD+SvSp6ZTEnSs2eMyRsINz
vt4tY0J4EVmjWM1J40Jj1/ReQbhevdfZR3qlRjucCgCpp8qTqnGuwV7Fgoq0gpIs
XOGfI6+BCpdJfcybm3WncuvgN9a5f7k9RuNBV4dXX/YifHTJaDRmKGqvuVFzhTqe
owkzkIJDT9dHjtcfLyu4XcLgFqbgJodtclVHcjDuLBIQDuclQGgnI02nDh81kqnV
JzVtR4S7lDfGqbopxXiMx9Qol9obOQYXyJFMlVDLSYtymQfZwhbs5yC6qsT3NR3g
ccjwa6F+dnRBCBw5iNNTUD3G+f6ixUcqaSKxPtQCCNGwMT9K0vjsOybficiUN7R/
byj7u+ViXgLtgiL9fqwWIWAV3VyoW+69oWw+C7x9uRvK6XYleD+EjVjjCEakfpeM
Qs7M0AdDTqUU0/A8xqa7EPG5FPCA7tZP4eQA7+hz1/X1RoO6JcEsuv+ySD0szJLC
+n6GyzmrkejNFFBcUzl6VaT+OKGyMVZ5+FgOEpWJgRJX3eQwFksyp6Dmw1w7rSMp
z9R36XV3KYTXRr08KIYaNz8SWCslKr2nRRMeKuqHYIV9ca7a9ci8LThNV3vgGPLw
iR2tcrx7G8Za/u7N9Lwq8jQao6k8yDxXXZq/jrWhmk/tGwmumylUlYSzcIttz8LZ
uJToGGVuh2rlM8jf0itrunqgMIjOC7NUHJ83TeHNZc39ax29K3x3h/fdlaS//4lR
WeaweXUpY1zAga9sSUYr3g4UMBteYZeVw4MemZUo96WTbYNxt78VbJXwMHxpQZWp
TF3YUPYc1X/P99PcGcHw0iykf2sCmMGEK+HdnixDAY+gcx5QOGzTpez1TAyVAjcb
fMLmrb84Rms8ARpnfW4ycaXbKN0W1xAKrYLM0G6pgc1Bd3hDsvLd8MSUk52ZpVpN
mGEESWg6oGlD4C/N71akF/VBRvue7GKjtJNiZ871nkV4q7YQhhKwzCcYnY3q7HoH
4szqyM2pqXtl73cnnM9q9BMywS1oIE3JRCO0i5EPsTFMyzlS/15ERD830WSUbq6L
YaZoyTX+dCrrlYAefiNo3a5UWZglw1/F6K84qzh2cieSmPbgkoxWemLQAS6mNpXc
qdH1WurXgAS3BgTH9hRUWdW2IpK/BoNsRMicbcE9urZsuWq4/ITvlgNSaE3vV36M
rg5i4HzdxQBqi6aUGDmAlAgEpowtIE+cSSvBjRVYFkgFlOqX2p8RSPBLgBglXSIL
K7ggnND6FHHpVY/PC8XfTwhQgiFT4qJuT71Y9nZkUk+HJobBNNHBlS69H/p+s9iC
WH4kWzc/G0Dxn6QodWhEmSPo3uRFIzNAzwxU+sW2rBwGsT6J7gkQ9477YoOgrJuR
TLuXEWv5A6rATASW95rxxAG9yEGmQ3O4a7sZqqaqJm90p+/5YOAzL9hD18a/5aNU
UG8dlj9OI1sIk7gjXiaH4hoSdcOpje2NvArveL4tApLhyJp0IFb90Anqb80KDeS/
1jXQgIsCmQITAfv7Y8FM2z/3N0/nECH/u4sm4bykQWJRF15AVYqNukmZe45JSNF/
NOFGaYAczKKDQdU2p5dnda/wVFaCDUQ7upiy22k4K64gcZ9o9WeQ2WVCLnFOx6Hr
+09+sMQ0N1m9WYi1s6AnLkUWDHOsHi532X67gq8zE1OlH/4t2/eaWXLjNAEW3d12
a0W7/4UvnPc3s7sOxomDgGd0DE5WeXGxXmggZwLt6kApv8MRkJJK7OZCR+fmT8I7
khs1oFZonXBTT433uYKX/k6IkOsf04Q1Xv2Td+RK2nPds/yqYjDLaCBvAORkDyOV
rnmih7wOxjW3mNbonTHEQ9K+eSrRk8tYB2vKocW1ZODbNTFO1OLDz/yZl0j4/aMY
Ahnj5mBFAier6fVWNLiKFTwDRrtvAA/2WR8UU/uACXFH3S1Peqcomq6ptFvq4+ed
z9qDIpv2s03bjTzbIeSRjCGzkQZRPQWHO014qcy9zyiIJu25e0UcuLXQDDPbi/cl
79ITIv3/ujKC96oTP+Vod7hsHeMZj5G/DHnkj82zDXcskBqhsIZPW6m8akI+iYkZ
gOdl0anR0mK2MIOpKZ96+fHQ+1iyIjoyGdCTaaBytZozClyiBOGiaTBQpn449CbZ
BAqiIgbeq0i8hh4hLpoMGLl8AKMB25CXaBj0Wx2X2PcJqhW397Hrssq0hHlJ3vPV
NTpEkvNw0Al9JDRKbyu5VV3ow2tIGquC6YSt9TslHuMHxm1ZxCCrwXGXd4cGYXcz
fGOUvSrTBQHtScJXmgc+25Zu6n38Onw+ynzr5xFq1zL9hoVEgi8Tf15LdapdQFI9
MtRjSDDSaVneNorTmfi0YidikLc9VR2Bi4epYtHDKOGAM+S1IuUiP0lRBtQoVlxb
w4O9Zpqf+0HjAn91qdF2MVmWoxhhL6FXRvKVmg6d0y6NynOPP5fU+bi+Y9n7VfjG
w3xK7wlKqP6BEoeueZm83ebjfZSUymefNuR1PeJI6UVRsu6jj5UGGw6SYt4SBpZD
MEy8z54UsodQocwA7V49eGIiAhPoSHO68JriODM90TR6TPSSTdaiUXGjFGYg0dzJ
S5zf+qQ6o040WAjBTu9X1EdaCFynJoAmr5gNWaA58ZT+I/GSYdFtg1k5YtXFpZXX
raaZFQ0F5/MMJii2NsQ8+m0+iPEjycXBAgwEIxBoxJppQ/wHeiS1Q4RD6DYcQTlV
GJ+po2Zbr8p2jY2UvEghMRkE6lhsgfL7ybwqztqZCSAAgdUSHe4nCU4CNHklKPFH
zcZIaB+X8MOfrYlYUAKIZN6aKEt7QKTVF6ahRNIqDO6sxAYnyCTAWgP8N9fkL7Q2
UtcEn2ao6z5hjX6rbtwByuiIBl0VB3kipmiBtTk/B1X7f4iG8zH2SfccrMyc63RX
ecWQ5BxdBVtKoKy+WCn2yX6Zf1VoqUekziXiswXQnvpieEpXu7yBSWlZHCuEnrX4
X8FoOBfO6mEG4VSOO1Ce+XpB7ipqRVRBOFhjGGWK3tdAoXPFeqOj2xXnvbGJXmw8
dToPwjve3HYkWQmyK4eQcmJuvKWEgU12Uv1GLpffKYMj069ZELOyvQVzhmqTVfFB
Uic2IQ7LbCOVE6c74QQzzV+9bVvytWyMVRfnKQhqwcHA7njlaT1mScL8ptWlnA7t
OZ7s/l3K2cNwAS/2Qc98L49pEKhCWOrxqOS/f+txRuNH5AtYfDVlYwc2JM46q2iA
o05/XOcH6xmc+5qzE2By9B9DQrK2gAPEPOZJYiHGf/h61c2bJ/Q61bBIaVecc12V
Xgz60LJ1hoqXoWrtH1EGo3mzE/rQ0xd0Pz88gP28L46Q5tsSk7QFm5/g9usWlNLR
+oV/48eeTZLUBQa3JsDniwsyWgbSbjQcUhbQ25ZusyonqA/OfysTSBVrOJGXX1bj
MbTpxappo8qnIG7TIpAMY4/BviOI+07KR7DpVLnD2jAU3fysOJQ4Tkbt4n2E+vFV
rkE1NW5R5tqEsP2RJqbzuLmhn37BXWKvxg4qJJNG/M1X9BCQHj4Id2Ixl/BNLJJ8
PQLse+BaNLegXs4M1V9PLwc4R6wKmgL6NFme6jH+xhqaQGdX7q1O9WVBcDsaRG+0
b/6TU/TtOHe0Y1VvvOK8VRg/R7uAR52UirySqrHOPxxMIITcu1dDOI01hXMA9wvj
ZnAtTuOfDVsYjm2eTiJYXLbpQ1HcLLFgFolqzY3RIngLHhUshcIr2970yRqQGieD
EruQq8/9I3OUvWQWLZgBN6fiY981LX9l7yDHBE5jDiZzj/cxmBNGzKQeNt/Wj1JN
m1IUX0oG8aC1OQgbsoWPi+pnU1XwAuDInNc1BafGJWgI/21D+qzalfjICvoJWxPf
nsfJGrpHGpdjSmPOvkp/CGeP1klT+fj4GhGg4Ys94uSbYyCfb4y3beHCqlRWnWLW
/zlw6EQrXgcS8cMJ8P1jc0O+h200Ui8g6LOsAfebkylIVrpjPhN+lnxJ2Gi8MR9c
e3G3DWTgGmrMJDZSQMC6qC7M2yArdSI4FUplfUKF1UYtjdOBpSii7oOKT8Cl4UwL
M7ObCupUVOlnTUhH9kuiR8cUawiJmt8XC+5U244jaWgKPZEOGNTzuJkd6CLaU6Zc
r2iMGn0j2u6BNFiO2fsOcshdMvSCCLaDwdsICArNC0hFR8/CH49Eku8akYEwqeDr
Ommd3YgR7T+iRfIrHg2s6Zn6DLLevJLY3x0/d3T4GnQM0bswdGqW+/n3S7KZW48c
jCeLGY4Tdlp/SrY+KC3gdvgzizmVVi/YzmDPMc+upcBd6iTbLgEnzmqJ6c3r4w5v
ZLTszr104j6a/6wgYgCiNnLkiR9A+iW+xkLSu0wh8qy8XjJl9ya/GHGNySZXpi16
vBqnOlQoc9VYnvR0w4kdtiVFmmqNN6KRmKof2x6PxOmbG/NeBC960NT1BZ0QrKsT
dz0uhayL9clvVZ34Z0p4aubwBn9B+Vc8kIwFta3zL/KI4SC/TqWuiVrMehPW+BFX
rNLvAwAvckvOg6dgqagcwXiJCn0UDEkmAzh2Ca5O3F7hdzeKNHUerauRYQjbxEF6
cNQmpZHjPAJtjhOs1Vx0/X8CFAMw7YZqM+BLTu/pO2CabwIfcsqZGnyhqGKo5kD0
fDjL9PvXc0G2hBwIilnsWkbI+kwvvfBNRlbVgEIQeuAGb+R7Jwr8HNfpuqzM1B6Q
hGJSFzCi0xs9iFn+5cF4g7qjjrRldwH8Tsz44FdPZVx2fICEm2Uy6TL9Wt0ElWcy
pi8J2L28N+hWD/Bf7CKK3DLNUpnOR6S7YyCEyfQvMsoNvGgSqdr+a84h1pwW6zKx
+WoBhDt3TtUU3lsyFBAevt1k/oRTt5TVEcCoT2Yxp4NdZTyB1qkgiBcX045fv2RH
M+3TdsorGbIkp1rWkGB7kL0KFDOsTojqQBHOcaNUSAJ0dRMBDakKCDlQ+qSwkpGB
/NMsP5qSNBoEbVU0+myM2/cmYtr0HhSDx+qPJErRcQJwWmmy2crdCVVmiyg3W0nx
12qy3n9SOXGRPU+SHYuL07d3w9aOW4b+mepCaLXQ+GMtZvWCjHhvX1va8yi74eVM
IpUMKTNIg4ae2Vnv3wAm2a5gOST5VDGVODhSVm0vbBC3I3B/ao9powoc2v2+qHCO
Xp9i2dB86QmeJJ7/byzeZYwCZJE3BCBIPhhuAHPEHCKkUdP14JvvQhw7aVjpv5I8
z0byowOIZkdb25g73JgHf/6Pajy4nn+ZOF3A3W6odB/o9wQFXt8kl+haqU5Pmm5o
RYgrXdufmAS4w7qPBsmg+Z/npa944789ioluEi5Vj6uF1dT2jR1ZWg+bgdINDhy+
WclOwbsufip9faEQ3c9D71o5MhF1kd9g/vBHkhTxpkh8NqOR7s9HqD3RryU5fYIU
SEuRaMMDT0NfvyjPlR/KWRfFg/A5nH++mBWvLj2waCkKsXlXtYFiGtncs695DmLC
/3Pb244AZnIHvYmyPvakWr7l0eExJtzQOW2Nmya6g7P+8RDXyuZLwax9FdGoK7yg
nD1bzGX9c2BYVt8upGccvSyDBq+DImGZmiewntEyIeT1cS6vgcBXkydzyIo6HghS
v7KoAc2Sl+HAli3+gq07vOBDJw65OMt6wae7As/zbcLwK6F8Px/HJsmuXKnnsWtQ
dYMrNAJujxoBerd+4LqWTt8fbobFMW9V5ZHZUVS11ZPVchWoogOrmHsJjOp9bt9z
5CJqCQhQpXF2AelHuBJXYmFwxrJUh6nwY81HN1jd/syRyv/SWR1zBUPdBB1TO15J
BAkLxCIvGZVC6tqCk+0OJpMZ87z6V/gZbilfhyWnFVfDJoN6XugJNjP7Xi7rT7wd
SSnpp8L49hjnASn4onqP1djm/195qiz5BzQaC6mbjInMj4hPX+UJKXbTqD5q4w3b
IB5loBn4zPN9z3T6xSCtX4vznyQvSDnAJC+KJr6WQ7PiUKLefGFQr67WHhRp2ElG
eAFEAIE0+mgJWNqwlzaU+vK+rfJAicHt7eSzvHazwBy9k+RXAq883sF28QA+Jk5z
iO1u3EsvMidnC1m+59qaQ5d/uYPAtdlSszx1Q0Sa6ECjl5QduKYdEyG+mauYZj9W
LCFKNTZGbWNwXyZsRg0SlUbCacARnRc3kdw3mxX++pypsfQrRxWT9/JMwfero/EP
oKTP0WNe16nxY6LKyabYTalaQAxLAwdmYEp90YBPY91h0lr4iXuOFBRUe8Pol7i1
YuDouYxZc73YiEL2SBm5TZEWKlFQeiA92s1/m1NefArB6d+yF47SQ+YDYRgbs6xi
QuJ6ta5nkFhp2Jkgf3UZOtRTZuNTBadbrk5IxjJH1ITBMVvVV0HXRHHk3Dg4dH7K
/5gL6qWZ4szj6zce5v7itWJ9c97y1P0UaCQAHk1lcaA0UCbG9UqghGXAMSfxkwgs
n2fa1UFzGHO9G6M44MJUDNHAlXUOZAozXL7ZNvMjqLmf4PUirkcG/jgNVqRnTXYq
N5hx7iInuO3zZW32MNT/uGtIe3fyNFWCiLfgLUoQYrLODWO+akgv6ECUyDk/Mxjf
hr2ZHbtBBmTYMTuQgFsdiYrg+H0zoYz0dIpYfzjU24E5KZVou4IcK004kd/3mpQp
uH3wnA1dzj0RoM/ZzBFlKW1FhV1+O+CCbYrZ6pHmrbeQh3VOgeRstCTbvS4oLtER
txWAWXqinHTwfSm62ETlRfMKgqp9fCAAkZbaoaOVY3mm6t+EcrBJ4LjJDe2ZD+j/
R8pUYeq7uHoBU26tcwiBVe6bwhUnSdcBXJJHV1gyChn5+BO6rSFSmooYCxL1rKnv
dmqZt9iDfDmRQn/byy/RUrbni8d5JwxNdw26RWsn6x6jZ6yeKlyXLlZStlrOz8Oz
anZ1+szPYeRSKMQ8LRAu/DzDxjmsoPris/zDs2jQ0W+nsN7KhwN7goIEcJGmhEll
zQnngDqmsqnmDwBnjuHLJte/yc0sBL3dZKO/Rh4OFHRyp9CcMb7UYzxCauFuPAM6
5ZyZyeVoe4uqQgEYFTCpNXMg65x2Z3KsFQTrdBJbxGDw0tqqfTgP4VhrC2M9eNQv
NQie8N2pJA/hAUBNpcY6rYzbVOaft1k2AT1dUa7C1B4yBPUQAQRt1yD/Kzv4HW1O
pyo5ukDVVu67vAHNjoswQ6ka/h2aRwk2+tvxqIva7zsMeAJijhu2iosQbM+jFLO5
szpfYRwdGZE1M3EwHJha9imEKrKKKSqebhFfm9+xowJOjeeZxiXiJb3j7M7QO2va
w5EMLeV/VnizbmpTWN260y83PD57g2NOsoZArvvbYF5GZAWn+iLjg+L0CXJTKI/Z
NZdtUggpLwbSdf6K5SHNwQaGrO1niNsoOPKQ5Dg0UhfhoBKLBthYLH8BExBOE1na
3ylnuvVJDbQRoOa1GnTnom9HwZ03wyIba19I/NlPhXpjY4Pfz6ITnkP0y9muR9LP
LWScCeZN+0JhY2JaO9EU1icqyFU1fyhe7UDlPbDTz/uR68u/qGcgtxbEhLMsH7e7
dz1pncZYY759htz7R2Dsk5CBsNjH1wVKRtHVHiBGuejI8Z8GUSq/pjAMjl1qJbPd
8xaphAG5XDoQvMwdv4RdtyL35cAFiGklFOMqeH9/nHuSBczRESGlqUVI7QxeP/pP
gbF7Dj1vPvHSorciQYas5R0nUuL1uNTbSLXngL/jIl4/MhUenUqq7rBMHSZ5JU8C
qLBgQRPT4sYAXX5PNh3f2QfKfQALueaYYUUvzSrVwPKiOfYs+EBywzR2qPn2NW3p
+2qq4w+l0b7ivxhZS4TIKmdAOKKH1K1igaAwIhCdze4Oawp7M5SCKfG2TArimGv6
flxtH/P4g2HndJ7+msu3vr8w2674WBO/Ga2AvMVSiw++4RfR7a9y9lYXhSUkyWBa
x8FFvPPp59A9QVPiOk2rbcwBXmw3NWIW75PiXaLzyJj+nldcoJEFKAWGJCIP0FTY
xc+orX4qRROfa6VYwbB+MPCpUGvPflUkfMC54tDjN0TG03r6f1th+C389Xxvtiby
M1AIMnRAIHoeFaNeeLtvFHV6uKUCNW+JTA1OwlRIDvFyR7DjrWXMEPdMIQD7+B2u
7iYvEWE3GYKPJSmkz/YUd5+SLM9ZwTHiYI6x++ZQ9UZg6xWOjjymWaNXp2eMNjt3
R8F8cjZjMcWPhvSoPbcIvayA1g4O4If0eAQRP0EwSNZ1mL2jynCloao2qZ2DTMhK
2KGTl77csQ7ya6SrllCa4hvjEeXoggPqVtqCjrtCDNSFTTCOHK4pgpMimN3/70Wf
mzs4eOFjq92cYGiG6riCCl5iJ9vbRDdJj0fcD7gr9rMNjsJBgnDAwnLWsqYVw2tj
Qz1r9E4PJldRNy1btoUy22urqy5kdQMPxm6OWBdcndskzuvQQ1bTWXhw0/9Qmj22
2193l4q8JvvQVhoNvaG1jxcj9YOXDwYOt9JsluPnnM9gZ9tsFr8tR9oIXGKK0lIn
BwEI8fp1K9kKchP/VV5TrApv4KIexB0t4gZl6QbgKtQ8NMeQnxYn7kg/fuMBozH2
DusqbKgaD8vXpwPoegoHo1QHb5janrP4kk8MngQuARuWCnbU9QwBHFv5tpn9CJ0q
JzQLn7mqNqCz/G7zhlVF2EKX7SXf5WSb/znG/R9PWDaqDaosr/eHTJzKU2MZb0ry
NdaAT5Cn96aLgEYbxDF193WPOXVi9GUH8tQATnNUjOrMu14HH8YvUOEGwOCkDi0e
WTS4XWluA8VJcr11G4FO5UG9C536uCzgaLMHW5PEQjX61Yq9TckOrUDYVRcN30IB
n5aEnsvUckIwvEuy0tuyn4baOZkgtXzJfdgscd23IbEAzumboQj1Eh2sJDdHsTwC
tS7Je9PSWKOSOs+DHVDqOZl75BxMgCArCD6LyFvMOkijTYXzViCtu9YhODbKwhE4
1bp6lTffvaTatYfLvOQ54GSH6jTj9uvthBd1hWEt2ha481LiKGJDQoEdgAvJ2BaY
NgeUp0nYplLKykaRAmk5xDj/chTYh6Ew+NOWlb47RbpUHkJvoyGt3TPP6SU/V6jo
HiAy1s/1cDh1ME4vxdfRQkADerGG/wy8N5HggTidVSDtGXYBL1vMYA0QKLdKUuif
wKZAgmM93n0jjUHYGptHX9pg7aDFdbEyNYN3Oc2dwflj7jzua34pryFky3h0eX6/
XtEemf2gcZAOmoJ2J10aM7MIBEkXezNQVfuHEvBd5dIrjXjS5eu8ypBmcOdnb6lj
Dk37Ivi2/HAtCqQvib5VErVcIkyCDC92XcmS4VQjJS/L0QQrz7klSC5BVNsaSbtb
VKPaDrE+8oE5LImX0KP1LJyf1Py5KQeW1CyxaKZAOF6+bO7D0A4f87NIdYseh6/o
ZfZXTxVvigakzcRCxCvdLOIKpjqQ1jj3dj4lfVsXQexdAi67xTqn/kuZlrlMB9nd
wGxxK+mB38Nm42dnMCSsWh3ewVVolEttLOw2zZ5mwJjT6zXnxBJtkyVLpq2bV5Cp
k/j2FYXARHz99TZ/uJxtNI3gpTfSglul32gpTQLbbi6x4nr8MkSycxsKzvdKRyuG
jGAlhkBJ/FZ5JVTcKF9uCO5799pNCJ+rariVOuKfWvbS4c0yulV9kWKODjKKZXwq
LQpZUz33wfiCaa9v5v8DijMO3PmJgxrLguiF7MtI1R4VHVVWWtaU3GsaQ0NLWWCF
MzONTZCnyNBiWjKNJqS2AKxVTznmMSMl58OQ0g7QZ+VVE2W1HObnm0RwXrzWw5tz
FAKQRFvkOWkXLlypSuRR+X34psidjnu8DDu59nk4tDbWoN5G1gpoJU7snLFKSmkY
vGLDtZ6fQl6q+UGQ2tWkG01DYUC0NEwofpvMWvJxqdunfAvlbRXPCp1raBSHhcaI
RlgKtQmTm6UNWPGmbjyl2KXVaMvJdAkLGcugKqEWJY3DsxR0AZzXLqWo04kSWGLQ
S+CbzlGAk9LAAuKpD1EpGkMGh6Za1dX+LBjWFcVJzLtE20j9ZKwqn18fS9kQy6K1
WU9tNO3lnqAJd+JZwS7KQ0mGJzBnZ4PQohi0efv6SOJOfv+5/UOHFEqQdUNh4WK1
IgBzi7p2cMbQFgLgpbzav0LZUdeCXmGALeH6UQbKIyCYAJfjUDHQ7o0sShTGoeRA
LZofGdjvs6epjKkqyyLX0xqILKCNmoM4uzCVHSRIhadyq5pKcF0W6SrzhMGJ7DuE
DkxwBnBGbC6BUkjLW7rSU6UZwyp1GU0xi86Uzi09kp9sbaHyGRJZfC9953JRFLM8
wLwTo0TQm353av1vsHIEbQd/Z62+TRey8FpTcimTnyKBgyl02hkHfcZ8SDkE66pm
oHZGU/QW424skYqVzWIz14lHORx6LG5MKrh79X9iQI8nR4nyZo0vL+QqtZSviwTu
enbDWNnoKIwGyU/+OS1+6sRwN6ds4abu9c2G3QZVyIlWft6AYIEDpVS/uW539z2P
NPcCiYcp4WwT6ttRyhkzPcV5Q0he8pWsiTOHjRvPXxvlsduuOOcmW7SUUwxEMzsN
RnUWJrL7Ycvduholq3GYnudk15l5kknAfaDyCZYW+aU/v6RZSh4xmtXCjwvNUYrt
7od9Dah1zX+2656h3YWEvVujYwjd7E0vV8p85VlR7ONqTAsy4QAF5IBAyt75SySp
UfQDGe7qzPh/F3YUF5JCPpKzvoUQ8s4f1/gRz4VNT48tJJrQVW6bSGCRHD4Gacy6
5OYMhOi6lCBCYDslpfK173hgnKcT08aLBAgBUX2AQpbuH+4bx2nyz2xxFmFRHJJD
sPNG3K3hqgMtz0TAaQsM8qeYrJkYOJo+Ebh9PQlcGz65FFBd6A+V42QzsQIdN8E4
A3yN0t47dleVh3k02hLT/A2yx7KXf9yWJzAyiJWRViW0z8YQjrb82k3H7Ene1KOD
1USmZ0CSeLnncD4y/l7GeAANQ+RQvPS+JC58glMbjSCP/e81zHsA+0fDv86hDj86
6pYG6KxG6DQ0dY0xoX35SK4DW1+hYlBD+WCKi92N+b/1wBFreovN+d/cFXZ68MIK
i/ee+lojB9SVfhzr7qQ1Z1GIppzGtvVq5B20Ndnoy/39jQ5Gpm/gDiWZaI7TxAMc
74APr9aWNXTcIA8RASlm6gNGo9vTWs16R/YJJpPQBwnXUKrFyZG77/UkDqevc4FN
iPZYphU9Rx3eU3a8S8Qa3Re0Rsop08Ody4y389LIHgZX1RIQ9FfM/6fBkOTH7wku
tCE248qx5VqdOeBSxfigQCr+g5ZVYH3g3mNB233AWUWP8upjCnkYa6JI7Gpx9L5d
B0SQmkWdOdymKYlqu6ICoGBD/Bqxeu8lS0NN6sl9yDqy54qzSetGWEekMfbHAtM5
VmEQkqCmLVnR3AUPpBZybFlsAvWiWojiS9PZySxzEsWVaBN43wh9J+yAv8FCOI4R
WTS/rg33KNBh0VhqioCg9cooksyt4IhluJdznFiMGGKx+REnVHSIuRdNHVpLmxhE
PmKSCKUfBcuYJEEUWIk2VQBx4YY44RQNguHRLPgVqH98vOL/hf3mhcc1GVdWRpFH
lW8bhyTHJK2M6+UgwO05kwtKX4jfU+/V3KfW5oJ59CpwgCRDnL+arwfCQN38Dc29
DLDEgzqvm5H4icFLvfDSXMkmfnHpkDrjMAUzWwqXHn4+PWsGc2O8Yr1EUTE8MrQq
gmXIt6R0jpQ4Ys2DwcRPdMSXvT+11MimYtF5FrMFR5s86VT6ZTh5virRgZUFadER
y7o2Pp6ak/D0XkReMq1JJr6dPoxV9yDqF8U6/6KhR9xOCI/iUa3o1NgEY3qdOfoE
kxIK613Hn4qqxMoZyw/LPjsErWUmM+FYXSjx6Iia02zM7w5bI1u/ETbiK2Smx2oo
afQDAuklOsb2+XUPWPWRocWA/N80jqnRxOk3F0AA9rqAudgMB9Ee8p4Cepi0CELL
xnwZtZE0ieuldb+ZWECTfjvES0Thcaegvorui9UPEcN0gmzwYBWgDnHfuTgG+xI6
XtqkkFp5tcswBp2d9oL8xmba3v/0v48fTULZgh2oyd7EvGMOZlMtr/QMaj3s2hWG
HdCIrFsSiAcYPmHZL3lOCGQ8mbfvQ2Gtfzpub+HHw7K4H/6uMNbVy9SoD8n3Q1jJ
TmzmAu0To8Y1rXj/HIltUq37UwnvoQthhKFP7uTj/CSMNROiZ0uSAyQafTEkfqJR
DHY6WZQ3cvCEo/aLKm3M0uZrOTGlb0kSQJlPVGwatN6UELJaXjvHPMYc+YMo6taR
VTzNErxx7vISPZuay3wCSlqh9YpOQhet4tSTRoG+lJT28YLu1/U6azDjqsrqpcoe
H46xuMW0TzOb+SFoPhIWBYLxB3XjUvvNVAk1WJN3ts2cgUwSJims0QT5Dh9OhEwg
LZOfGvWUEQyB7Enu/TE43oC+Fr6M362YZ3VgLAD8X1Z09OoaGmQ28vNtdL+gSBMs
m8fVKvuZ8XTtPJuH63LRa25y0OG0uZfAWWb59XBkXYc7S6Jq+odcVMwIIGVVsMAd
JRzJ34R7d8g6urZKTME7FQPTVrrD2/BH52Ulh6VydVM5ix59vbt2s3jkVYEeVl60
AX4t1Yw/AGAazru76hXE3RF8ay3csM18QRodJ/KLseq55+UxZJjfGHh9BDPdW2Qy
ld292uGesUvOGa1FgqnGU7GdF3JOtt8XQ2aLgDraDN9EzYCEWSQkVpZLtPJyBk9i
oRY3eeFn1tLgkNn/MA3dDWOjTTx9GurYE10YM1g52jViVVe0S1EI+HgjgKEFWbf/
lqxNpBkbJY0QK/0/zIyuUG2YeQSzfJYP92rnwcoiFtxgpYaxMc7RBu3jvVyn9sjw
RHbM2jPLxOUWkDriTBHwg1legwqbUUgrPkaq5pcoWaFlfvrCUWVfJpxf2RaOJtnG
jL5b5WZEey05hYIZ7TLkW7Ccd1ICAfNUeJYSRQimuk7bN6EZ7CV23gnbzg7T/t6P
IraSvzpdCFx9qaC9Xp4vdTPxA1l9dRX0UkvtCUqOdMSWwUWZvNT7iALNaBsGvihB
iTz0fzxeMe38Lj5E1mioD+nc1PB2BfrldyDeOogNMoL0FbHP5pbQhOGlc3qVs0gA
xxNXP8yEp5ULfgyzPkJCXJ9QKQf3aQNmO/d8gAiQSbhNiB9f3dYB0Y6bCx8Chfc8
O6HrV0tC7X1PLikTQcpvSajTjPFuVfYS0KgK/elCe7Ym8QzWzcK1NtX9AU4l4rkO
f983jsKOoDqU9JWjvICf3iYaaC4AkkK4hTTl5011lKZqJsCiFl6+DYlLkPx7c8gb
YDlHvH5ClU1KrZpVmqZGAQ1BqgyZ7+sTVk+f/cND4toTG6cffEdX+SYzMGe8+m2I
p9XvLFXLj5uoNGC7ve8TQrcm34ilYGT6Mu1Bn7q9fJk=
`protect end_protected
