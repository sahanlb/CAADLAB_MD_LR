localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTX_CHK = {
  {32'h41133cb4, 32'hc2bf41e2} /* (15, 15, 15) {real, imag} */,
  {32'hc18072bb, 32'hc0b7fb3c} /* (15, 15, 14) {real, imag} */,
  {32'hc086cd42, 32'hc18904bb} /* (15, 15, 13) {real, imag} */,
  {32'h419c8182, 32'h4187a9ae} /* (15, 15, 12) {real, imag} */,
  {32'h40577c78, 32'h4141cb52} /* (15, 15, 11) {real, imag} */,
  {32'h40e34146, 32'h410fb1b4} /* (15, 15, 10) {real, imag} */,
  {32'hc0f9bfe0, 32'h40a8d559} /* (15, 15, 9) {real, imag} */,
  {32'h4070012c, 32'h411e026f} /* (15, 15, 8) {real, imag} */,
  {32'h405581b0, 32'h40c52940} /* (15, 15, 7) {real, imag} */,
  {32'h40d4e5d3, 32'hc0f388d4} /* (15, 15, 6) {real, imag} */,
  {32'hc12331fc, 32'h417612d7} /* (15, 15, 5) {real, imag} */,
  {32'h4165a016, 32'h40941ed9} /* (15, 15, 4) {real, imag} */,
  {32'hc1d425b4, 32'hc16a4d9f} /* (15, 15, 3) {real, imag} */,
  {32'h4228da55, 32'hc069a060} /* (15, 15, 2) {real, imag} */,
  {32'hc25549ef, 32'h41ea618e} /* (15, 15, 1) {real, imag} */,
  {32'hc2820fcf, 32'hc1194d68} /* (15, 15, 0) {real, imag} */,
  {32'h41d6b02a, 32'h412d5c65} /* (15, 14, 15) {real, imag} */,
  {32'hc1ca6c28, 32'h41558a4c} /* (15, 14, 14) {real, imag} */,
  {32'h403ced98, 32'hc1092452} /* (15, 14, 13) {real, imag} */,
  {32'h40fa846c, 32'hc107dfc0} /* (15, 14, 12) {real, imag} */,
  {32'h41a6afa4, 32'h409efa16} /* (15, 14, 11) {real, imag} */,
  {32'h40aca01e, 32'h40ba2a10} /* (15, 14, 10) {real, imag} */,
  {32'h40809881, 32'hc14353e2} /* (15, 14, 9) {real, imag} */,
  {32'hc1b85b9b, 32'hbfa1ea48} /* (15, 14, 8) {real, imag} */,
  {32'h40620ad8, 32'h40ec7db3} /* (15, 14, 7) {real, imag} */,
  {32'hc15382a8, 32'h415a9c7e} /* (15, 14, 6) {real, imag} */,
  {32'h418590f8, 32'hc0c17918} /* (15, 14, 5) {real, imag} */,
  {32'h403b899c, 32'h409c37fc} /* (15, 14, 4) {real, imag} */,
  {32'h4094d8e0, 32'h3d4dd800} /* (15, 14, 3) {real, imag} */,
  {32'hc100ac50, 32'hc2201f7a} /* (15, 14, 2) {real, imag} */,
  {32'hc233f5a2, 32'h42123894} /* (15, 14, 1) {real, imag} */,
  {32'hc24a8f82, 32'h4181d3b4} /* (15, 14, 0) {real, imag} */,
  {32'hbfbc1620, 32'hc1835195} /* (15, 13, 15) {real, imag} */,
  {32'h41d3a2d1, 32'h409823ca} /* (15, 13, 14) {real, imag} */,
  {32'h412653ce, 32'hc0d4a658} /* (15, 13, 13) {real, imag} */,
  {32'hc1df9f28, 32'h4046c2a0} /* (15, 13, 12) {real, imag} */,
  {32'hc145c183, 32'hc19aea48} /* (15, 13, 11) {real, imag} */,
  {32'hc19f3802, 32'h4108cecb} /* (15, 13, 10) {real, imag} */,
  {32'h40bea4d8, 32'h41153064} /* (15, 13, 9) {real, imag} */,
  {32'h4032c258, 32'hbfa3b8a0} /* (15, 13, 8) {real, imag} */,
  {32'h4191815e, 32'h3fb15e36} /* (15, 13, 7) {real, imag} */,
  {32'hc0d8f6df, 32'h40a11eb9} /* (15, 13, 6) {real, imag} */,
  {32'hc201afe5, 32'hbfcac472} /* (15, 13, 5) {real, imag} */,
  {32'hbdd3be00, 32'h41816688} /* (15, 13, 4) {real, imag} */,
  {32'hc1cbb554, 32'hc0ac1030} /* (15, 13, 3) {real, imag} */,
  {32'hc1b26d4c, 32'h41e2bccb} /* (15, 13, 2) {real, imag} */,
  {32'h3fa254a8, 32'hbe2c3900} /* (15, 13, 1) {real, imag} */,
  {32'h412b9d96, 32'h400d6edc} /* (15, 13, 0) {real, imag} */,
  {32'h416f0d4a, 32'h41fdc881} /* (15, 12, 15) {real, imag} */,
  {32'hc1d17f09, 32'h412722ca} /* (15, 12, 14) {real, imag} */,
  {32'hc16c7136, 32'hc0b1c5ac} /* (15, 12, 13) {real, imag} */,
  {32'hc020a970, 32'h4147cd40} /* (15, 12, 12) {real, imag} */,
  {32'hc1665b5c, 32'hc1acfe76} /* (15, 12, 11) {real, imag} */,
  {32'h40139aa2, 32'h4125322d} /* (15, 12, 10) {real, imag} */,
  {32'h40712cf0, 32'hc0ae1b0e} /* (15, 12, 9) {real, imag} */,
  {32'hc0ad8c03, 32'hc140ae3e} /* (15, 12, 8) {real, imag} */,
  {32'hc12e7e6c, 32'h3f29a420} /* (15, 12, 7) {real, imag} */,
  {32'hc1979367, 32'h402ac290} /* (15, 12, 6) {real, imag} */,
  {32'h3eb5a720, 32'hc1567c44} /* (15, 12, 5) {real, imag} */,
  {32'hc18407a1, 32'h408442b7} /* (15, 12, 4) {real, imag} */,
  {32'h418fb212, 32'h400523f4} /* (15, 12, 3) {real, imag} */,
  {32'h419a9740, 32'h40560908} /* (15, 12, 2) {real, imag} */,
  {32'h41846588, 32'hc14cbe04} /* (15, 12, 1) {real, imag} */,
  {32'hc091eeec, 32'hc0d7def8} /* (15, 12, 0) {real, imag} */,
  {32'hc17c746e, 32'h41e74158} /* (15, 11, 15) {real, imag} */,
  {32'hc0704c38, 32'hc160b642} /* (15, 11, 14) {real, imag} */,
  {32'h41ba6c9b, 32'hc11a8675} /* (15, 11, 13) {real, imag} */,
  {32'h409461f0, 32'hc1a79ac6} /* (15, 11, 12) {real, imag} */,
  {32'h409ac1ec, 32'h412d4d78} /* (15, 11, 11) {real, imag} */,
  {32'h416870cc, 32'hc066edd4} /* (15, 11, 10) {real, imag} */,
  {32'h4049f60a, 32'h4009f95c} /* (15, 11, 9) {real, imag} */,
  {32'h41a0d9f3, 32'h412f68fa} /* (15, 11, 8) {real, imag} */,
  {32'hc162ad37, 32'hc1175a3c} /* (15, 11, 7) {real, imag} */,
  {32'h4180be00, 32'hc1cbba32} /* (15, 11, 6) {real, imag} */,
  {32'hc080b43f, 32'hc2033b46} /* (15, 11, 5) {real, imag} */,
  {32'hc1ac04f7, 32'h402bd37c} /* (15, 11, 4) {real, imag} */,
  {32'h4198ad2a, 32'hc016d5e8} /* (15, 11, 3) {real, imag} */,
  {32'h41141e3b, 32'h4144840a} /* (15, 11, 2) {real, imag} */,
  {32'h40c454dc, 32'hc185db0a} /* (15, 11, 1) {real, imag} */,
  {32'h4170e936, 32'hc077ff90} /* (15, 11, 0) {real, imag} */,
  {32'h40fe99aa, 32'hc167d818} /* (15, 10, 15) {real, imag} */,
  {32'hc1911f0d, 32'hbf8a40b8} /* (15, 10, 14) {real, imag} */,
  {32'h41382562, 32'hc04d3b2e} /* (15, 10, 13) {real, imag} */,
  {32'h409839f8, 32'h412ce053} /* (15, 10, 12) {real, imag} */,
  {32'h4124a951, 32'h3d869240} /* (15, 10, 11) {real, imag} */,
  {32'h40c400cc, 32'h3fd76ce4} /* (15, 10, 10) {real, imag} */,
  {32'h403b030a, 32'hc023fc10} /* (15, 10, 9) {real, imag} */,
  {32'hc08fdbe6, 32'h4138ea00} /* (15, 10, 8) {real, imag} */,
  {32'hc0d97ee8, 32'hc13d87b6} /* (15, 10, 7) {real, imag} */,
  {32'h404a653c, 32'hc1d28fba} /* (15, 10, 6) {real, imag} */,
  {32'hc0bf559c, 32'h419aed23} /* (15, 10, 5) {real, imag} */,
  {32'hc12047b5, 32'hbf10b2d8} /* (15, 10, 4) {real, imag} */,
  {32'h411875dc, 32'hc18a1682} /* (15, 10, 3) {real, imag} */,
  {32'h4197340b, 32'hc06fb5d4} /* (15, 10, 2) {real, imag} */,
  {32'h41270cf0, 32'hc1d3808e} /* (15, 10, 1) {real, imag} */,
  {32'h419989aa, 32'hc1343ef6} /* (15, 10, 0) {real, imag} */,
  {32'h4159dff0, 32'h40fa83f8} /* (15, 9, 15) {real, imag} */,
  {32'hc0e57aa0, 32'hc1668f9a} /* (15, 9, 14) {real, imag} */,
  {32'hc12728df, 32'h4106e2b0} /* (15, 9, 13) {real, imag} */,
  {32'h3fcdc920, 32'hc02b3d66} /* (15, 9, 12) {real, imag} */,
  {32'hc0b17f30, 32'hc149868f} /* (15, 9, 11) {real, imag} */,
  {32'hc0c375e2, 32'hc1819977} /* (15, 9, 10) {real, imag} */,
  {32'h40e397cc, 32'h4069862c} /* (15, 9, 9) {real, imag} */,
  {32'hc0502c9d, 32'h4012385f} /* (15, 9, 8) {real, imag} */,
  {32'hbe597190, 32'h40c7aa82} /* (15, 9, 7) {real, imag} */,
  {32'h40b3b21c, 32'hbfd82fb4} /* (15, 9, 6) {real, imag} */,
  {32'h4093376c, 32'h4043d01c} /* (15, 9, 5) {real, imag} */,
  {32'h41533770, 32'hc15ce22e} /* (15, 9, 4) {real, imag} */,
  {32'hc19b2914, 32'hbfe68fb0} /* (15, 9, 3) {real, imag} */,
  {32'h4123c094, 32'h416bfdc8} /* (15, 9, 2) {real, imag} */,
  {32'h3d9b2a00, 32'hc0882e1c} /* (15, 9, 1) {real, imag} */,
  {32'hc01d33e0, 32'h40f13888} /* (15, 9, 0) {real, imag} */,
  {32'hc16d4490, 32'h410bd150} /* (15, 8, 15) {real, imag} */,
  {32'hc1114462, 32'h3f94677a} /* (15, 8, 14) {real, imag} */,
  {32'h3feff41c, 32'hc1537541} /* (15, 8, 13) {real, imag} */,
  {32'h3ffad6d0, 32'hbf8ba728} /* (15, 8, 12) {real, imag} */,
  {32'hc0f77328, 32'hc102ac58} /* (15, 8, 11) {real, imag} */,
  {32'hc1048d69, 32'h40b6cea8} /* (15, 8, 10) {real, imag} */,
  {32'h413a0402, 32'hc01d7252} /* (15, 8, 9) {real, imag} */,
  {32'hc08dde74, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'h413a0402, 32'h401d7252} /* (15, 8, 7) {real, imag} */,
  {32'hc1048d69, 32'hc0b6cea8} /* (15, 8, 6) {real, imag} */,
  {32'hc0f77328, 32'h4102ac58} /* (15, 8, 5) {real, imag} */,
  {32'h3ffad6d0, 32'h3f8ba728} /* (15, 8, 4) {real, imag} */,
  {32'h3feff41c, 32'h41537541} /* (15, 8, 3) {real, imag} */,
  {32'hc1114462, 32'hbf94677a} /* (15, 8, 2) {real, imag} */,
  {32'hc16d4490, 32'hc10bd150} /* (15, 8, 1) {real, imag} */,
  {32'h3feb5640, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h3d9b2a00, 32'h40882e1c} /* (15, 7, 15) {real, imag} */,
  {32'h4123c094, 32'hc16bfdc8} /* (15, 7, 14) {real, imag} */,
  {32'hc19b2914, 32'h3fe68fb0} /* (15, 7, 13) {real, imag} */,
  {32'h41533770, 32'h415ce22e} /* (15, 7, 12) {real, imag} */,
  {32'h4093376c, 32'hc043d01c} /* (15, 7, 11) {real, imag} */,
  {32'h40b3b21c, 32'h3fd82fb4} /* (15, 7, 10) {real, imag} */,
  {32'hbe597190, 32'hc0c7aa82} /* (15, 7, 9) {real, imag} */,
  {32'hc0502c9d, 32'hc012385f} /* (15, 7, 8) {real, imag} */,
  {32'h40e397cc, 32'hc069862c} /* (15, 7, 7) {real, imag} */,
  {32'hc0c375e2, 32'h41819977} /* (15, 7, 6) {real, imag} */,
  {32'hc0b17f30, 32'h4149868f} /* (15, 7, 5) {real, imag} */,
  {32'h3fcdc920, 32'h402b3d66} /* (15, 7, 4) {real, imag} */,
  {32'hc12728df, 32'hc106e2b0} /* (15, 7, 3) {real, imag} */,
  {32'hc0e57aa0, 32'h41668f9a} /* (15, 7, 2) {real, imag} */,
  {32'h4159dff0, 32'hc0fa83f8} /* (15, 7, 1) {real, imag} */,
  {32'hc01d33e0, 32'hc0f13888} /* (15, 7, 0) {real, imag} */,
  {32'h41270cf0, 32'h41d3808e} /* (15, 6, 15) {real, imag} */,
  {32'h4197340b, 32'h406fb5d4} /* (15, 6, 14) {real, imag} */,
  {32'h411875dc, 32'h418a1682} /* (15, 6, 13) {real, imag} */,
  {32'hc12047b5, 32'h3f10b2d8} /* (15, 6, 12) {real, imag} */,
  {32'hc0bf559c, 32'hc19aed23} /* (15, 6, 11) {real, imag} */,
  {32'h404a653c, 32'h41d28fba} /* (15, 6, 10) {real, imag} */,
  {32'hc0d97ee8, 32'h413d87b6} /* (15, 6, 9) {real, imag} */,
  {32'hc08fdbe6, 32'hc138ea00} /* (15, 6, 8) {real, imag} */,
  {32'h403b030a, 32'h4023fc10} /* (15, 6, 7) {real, imag} */,
  {32'h40c400cc, 32'hbfd76ce4} /* (15, 6, 6) {real, imag} */,
  {32'h4124a951, 32'hbd869240} /* (15, 6, 5) {real, imag} */,
  {32'h409839f8, 32'hc12ce053} /* (15, 6, 4) {real, imag} */,
  {32'h41382562, 32'h404d3b2e} /* (15, 6, 3) {real, imag} */,
  {32'hc1911f0d, 32'h3f8a40b8} /* (15, 6, 2) {real, imag} */,
  {32'h40fe99aa, 32'h4167d818} /* (15, 6, 1) {real, imag} */,
  {32'h419989aa, 32'h41343ef6} /* (15, 6, 0) {real, imag} */,
  {32'h40c454dc, 32'h4185db0a} /* (15, 5, 15) {real, imag} */,
  {32'h41141e3b, 32'hc144840a} /* (15, 5, 14) {real, imag} */,
  {32'h4198ad2a, 32'h4016d5e8} /* (15, 5, 13) {real, imag} */,
  {32'hc1ac04f7, 32'hc02bd37c} /* (15, 5, 12) {real, imag} */,
  {32'hc080b43f, 32'h42033b46} /* (15, 5, 11) {real, imag} */,
  {32'h4180be00, 32'h41cbba32} /* (15, 5, 10) {real, imag} */,
  {32'hc162ad37, 32'h41175a3c} /* (15, 5, 9) {real, imag} */,
  {32'h41a0d9f3, 32'hc12f68fa} /* (15, 5, 8) {real, imag} */,
  {32'h4049f60a, 32'hc009f95c} /* (15, 5, 7) {real, imag} */,
  {32'h416870cc, 32'h4066edd4} /* (15, 5, 6) {real, imag} */,
  {32'h409ac1ec, 32'hc12d4d78} /* (15, 5, 5) {real, imag} */,
  {32'h409461f0, 32'h41a79ac6} /* (15, 5, 4) {real, imag} */,
  {32'h41ba6c9b, 32'h411a8675} /* (15, 5, 3) {real, imag} */,
  {32'hc0704c38, 32'h4160b642} /* (15, 5, 2) {real, imag} */,
  {32'hc17c746e, 32'hc1e74158} /* (15, 5, 1) {real, imag} */,
  {32'h4170e936, 32'h4077ff90} /* (15, 5, 0) {real, imag} */,
  {32'h41846588, 32'h414cbe04} /* (15, 4, 15) {real, imag} */,
  {32'h419a9740, 32'hc0560908} /* (15, 4, 14) {real, imag} */,
  {32'h418fb212, 32'hc00523f4} /* (15, 4, 13) {real, imag} */,
  {32'hc18407a1, 32'hc08442b7} /* (15, 4, 12) {real, imag} */,
  {32'h3eb5a720, 32'h41567c44} /* (15, 4, 11) {real, imag} */,
  {32'hc1979367, 32'hc02ac290} /* (15, 4, 10) {real, imag} */,
  {32'hc12e7e6c, 32'hbf29a420} /* (15, 4, 9) {real, imag} */,
  {32'hc0ad8c03, 32'h4140ae3e} /* (15, 4, 8) {real, imag} */,
  {32'h40712cf0, 32'h40ae1b0e} /* (15, 4, 7) {real, imag} */,
  {32'h40139aa2, 32'hc125322d} /* (15, 4, 6) {real, imag} */,
  {32'hc1665b5c, 32'h41acfe76} /* (15, 4, 5) {real, imag} */,
  {32'hc020a970, 32'hc147cd40} /* (15, 4, 4) {real, imag} */,
  {32'hc16c7136, 32'h40b1c5ac} /* (15, 4, 3) {real, imag} */,
  {32'hc1d17f09, 32'hc12722ca} /* (15, 4, 2) {real, imag} */,
  {32'h416f0d4a, 32'hc1fdc881} /* (15, 4, 1) {real, imag} */,
  {32'hc091eeec, 32'h40d7def8} /* (15, 4, 0) {real, imag} */,
  {32'h3fa254a8, 32'h3e2c3900} /* (15, 3, 15) {real, imag} */,
  {32'hc1b26d4c, 32'hc1e2bccb} /* (15, 3, 14) {real, imag} */,
  {32'hc1cbb554, 32'h40ac1030} /* (15, 3, 13) {real, imag} */,
  {32'hbdd3be00, 32'hc1816688} /* (15, 3, 12) {real, imag} */,
  {32'hc201afe5, 32'h3fcac472} /* (15, 3, 11) {real, imag} */,
  {32'hc0d8f6df, 32'hc0a11eb9} /* (15, 3, 10) {real, imag} */,
  {32'h4191815e, 32'hbfb15e36} /* (15, 3, 9) {real, imag} */,
  {32'h4032c258, 32'h3fa3b8a0} /* (15, 3, 8) {real, imag} */,
  {32'h40bea4d8, 32'hc1153064} /* (15, 3, 7) {real, imag} */,
  {32'hc19f3802, 32'hc108cecb} /* (15, 3, 6) {real, imag} */,
  {32'hc145c183, 32'h419aea48} /* (15, 3, 5) {real, imag} */,
  {32'hc1df9f28, 32'hc046c2a0} /* (15, 3, 4) {real, imag} */,
  {32'h412653ce, 32'h40d4a658} /* (15, 3, 3) {real, imag} */,
  {32'h41d3a2d1, 32'hc09823ca} /* (15, 3, 2) {real, imag} */,
  {32'hbfbc1620, 32'h41835195} /* (15, 3, 1) {real, imag} */,
  {32'h412b9d96, 32'hc00d6edc} /* (15, 3, 0) {real, imag} */,
  {32'hc233f5a2, 32'hc2123894} /* (15, 2, 15) {real, imag} */,
  {32'hc100ac50, 32'h42201f7a} /* (15, 2, 14) {real, imag} */,
  {32'h4094d8e0, 32'hbd4dd800} /* (15, 2, 13) {real, imag} */,
  {32'h403b899c, 32'hc09c37fc} /* (15, 2, 12) {real, imag} */,
  {32'h418590f8, 32'h40c17918} /* (15, 2, 11) {real, imag} */,
  {32'hc15382a8, 32'hc15a9c7e} /* (15, 2, 10) {real, imag} */,
  {32'h40620ad8, 32'hc0ec7db3} /* (15, 2, 9) {real, imag} */,
  {32'hc1b85b9b, 32'h3fa1ea48} /* (15, 2, 8) {real, imag} */,
  {32'h40809881, 32'h414353e2} /* (15, 2, 7) {real, imag} */,
  {32'h40aca01e, 32'hc0ba2a10} /* (15, 2, 6) {real, imag} */,
  {32'h41a6afa4, 32'hc09efa16} /* (15, 2, 5) {real, imag} */,
  {32'h40fa846c, 32'h4107dfc0} /* (15, 2, 4) {real, imag} */,
  {32'h403ced98, 32'h41092452} /* (15, 2, 3) {real, imag} */,
  {32'hc1ca6c28, 32'hc1558a4c} /* (15, 2, 2) {real, imag} */,
  {32'h41d6b02a, 32'hc12d5c65} /* (15, 2, 1) {real, imag} */,
  {32'hc24a8f82, 32'hc181d3b4} /* (15, 2, 0) {real, imag} */,
  {32'hc25549ef, 32'hc1ea618e} /* (15, 1, 15) {real, imag} */,
  {32'h4228da55, 32'h4069a060} /* (15, 1, 14) {real, imag} */,
  {32'hc1d425b4, 32'h416a4d9f} /* (15, 1, 13) {real, imag} */,
  {32'h4165a016, 32'hc0941ed9} /* (15, 1, 12) {real, imag} */,
  {32'hc12331fc, 32'hc17612d7} /* (15, 1, 11) {real, imag} */,
  {32'h40d4e5d3, 32'h40f388d4} /* (15, 1, 10) {real, imag} */,
  {32'h405581b0, 32'hc0c52940} /* (15, 1, 9) {real, imag} */,
  {32'h4070012c, 32'hc11e026f} /* (15, 1, 8) {real, imag} */,
  {32'hc0f9bfe0, 32'hc0a8d559} /* (15, 1, 7) {real, imag} */,
  {32'h40e34146, 32'hc10fb1b4} /* (15, 1, 6) {real, imag} */,
  {32'h40577c78, 32'hc141cb52} /* (15, 1, 5) {real, imag} */,
  {32'h419c8182, 32'hc187a9ae} /* (15, 1, 4) {real, imag} */,
  {32'hc086cd42, 32'h418904bb} /* (15, 1, 3) {real, imag} */,
  {32'hc18072bb, 32'h40b7fb3c} /* (15, 1, 2) {real, imag} */,
  {32'h41133cb4, 32'h42bf41e2} /* (15, 1, 1) {real, imag} */,
  {32'hc2820fcf, 32'h41194d68} /* (15, 1, 0) {real, imag} */,
  {32'h420bdc64, 32'hc3006012} /* (15, 0, 15) {real, imag} */,
  {32'h41fc55ac, 32'h41809a46} /* (15, 0, 14) {real, imag} */,
  {32'h414793bc, 32'h3f8a3e30} /* (15, 0, 13) {real, imag} */,
  {32'hc103065c, 32'hc1945601} /* (15, 0, 12) {real, imag} */,
  {32'h41a62a13, 32'hc03cca30} /* (15, 0, 11) {real, imag} */,
  {32'hc191342a, 32'hc061165a} /* (15, 0, 10) {real, imag} */,
  {32'hc14a8cce, 32'hbfe7f8f0} /* (15, 0, 9) {real, imag} */,
  {32'h41d06860, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'hc14a8cce, 32'h3fe7f8f0} /* (15, 0, 7) {real, imag} */,
  {32'hc191342a, 32'h4061165a} /* (15, 0, 6) {real, imag} */,
  {32'h41a62a13, 32'h403cca30} /* (15, 0, 5) {real, imag} */,
  {32'hc103065c, 32'h41945601} /* (15, 0, 4) {real, imag} */,
  {32'h414793bc, 32'hbf8a3e30} /* (15, 0, 3) {real, imag} */,
  {32'h41fc55ac, 32'hc1809a46} /* (15, 0, 2) {real, imag} */,
  {32'h420bdc64, 32'h43006012} /* (15, 0, 1) {real, imag} */,
  {32'hc2d06031, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h42c8f3d4, 32'hc2b57a14} /* (14, 15, 15) {real, imag} */,
  {32'hc261d021, 32'hc13916f9} /* (14, 15, 14) {real, imag} */,
  {32'hc22d5090, 32'hc1344210} /* (14, 15, 13) {real, imag} */,
  {32'h406f7976, 32'h3cbb3c00} /* (14, 15, 12) {real, imag} */,
  {32'h41d6c25e, 32'hc206fcc7} /* (14, 15, 11) {real, imag} */,
  {32'hc1f7267a, 32'hc18dbfee} /* (14, 15, 10) {real, imag} */,
  {32'hc0d312ac, 32'h40dad2a6} /* (14, 15, 9) {real, imag} */,
  {32'h4195c280, 32'h40e6051e} /* (14, 15, 8) {real, imag} */,
  {32'h40838be9, 32'h4142a5e4} /* (14, 15, 7) {real, imag} */,
  {32'h412f0e14, 32'h410f6024} /* (14, 15, 6) {real, imag} */,
  {32'hbfcc0f74, 32'h42477f2b} /* (14, 15, 5) {real, imag} */,
  {32'hc16a769b, 32'hc1c84a6c} /* (14, 15, 4) {real, imag} */,
  {32'hc1dcb221, 32'hc1b189ee} /* (14, 15, 3) {real, imag} */,
  {32'h42506a3e, 32'h424d2396} /* (14, 15, 2) {real, imag} */,
  {32'hc1fc0dde, 32'h4249202c} /* (14, 15, 1) {real, imag} */,
  {32'hc2abd360, 32'h420042b7} /* (14, 15, 0) {real, imag} */,
  {32'h4224e501, 32'h42238ee0} /* (14, 14, 15) {real, imag} */,
  {32'hc1e9589b, 32'hc099d250} /* (14, 14, 14) {real, imag} */,
  {32'hc0a6fe22, 32'hc224434c} /* (14, 14, 13) {real, imag} */,
  {32'h411d3c78, 32'h4179de30} /* (14, 14, 12) {real, imag} */,
  {32'hc130d24b, 32'hc17bcf46} /* (14, 14, 11) {real, imag} */,
  {32'h41d7cdc0, 32'hc1f4a6a4} /* (14, 14, 10) {real, imag} */,
  {32'hc1a8c688, 32'hc108d2db} /* (14, 14, 9) {real, imag} */,
  {32'hbf7d93d8, 32'h42037aaf} /* (14, 14, 8) {real, imag} */,
  {32'h41cf483b, 32'h4137fdd3} /* (14, 14, 7) {real, imag} */,
  {32'h413b0e47, 32'h42242a26} /* (14, 14, 6) {real, imag} */,
  {32'hc18d42df, 32'h419da7d6} /* (14, 14, 5) {real, imag} */,
  {32'h413b22e6, 32'h41c5b028} /* (14, 14, 4) {real, imag} */,
  {32'h41a888e6, 32'hc1d6d79a} /* (14, 14, 3) {real, imag} */,
  {32'hc2119f62, 32'hc207551e} /* (14, 14, 2) {real, imag} */,
  {32'hc2ba54d5, 32'h4282a730} /* (14, 14, 1) {real, imag} */,
  {32'hc216de42, 32'h4143c002} /* (14, 14, 0) {real, imag} */,
  {32'h41ddfc5a, 32'h409e36f8} /* (14, 13, 15) {real, imag} */,
  {32'hc13bf810, 32'h418eaccb} /* (14, 13, 14) {real, imag} */,
  {32'hc0a06e9a, 32'hc1cfd5b9} /* (14, 13, 13) {real, imag} */,
  {32'hc19e5f2d, 32'hc17e6cb0} /* (14, 13, 12) {real, imag} */,
  {32'hc10927d3, 32'h4173c03a} /* (14, 13, 11) {real, imag} */,
  {32'hc1a6e52e, 32'h417f6163} /* (14, 13, 10) {real, imag} */,
  {32'h4172af60, 32'hc1248a61} /* (14, 13, 9) {real, imag} */,
  {32'hc180871c, 32'hc05c3b64} /* (14, 13, 8) {real, imag} */,
  {32'h40e39179, 32'hc0a2a362} /* (14, 13, 7) {real, imag} */,
  {32'hc1817848, 32'hc25a3668} /* (14, 13, 6) {real, imag} */,
  {32'hc235e460, 32'h41465688} /* (14, 13, 5) {real, imag} */,
  {32'h424167e4, 32'hc19d25c0} /* (14, 13, 4) {real, imag} */,
  {32'hc28a43ca, 32'hc1a21432} /* (14, 13, 3) {real, imag} */,
  {32'h4114e82a, 32'h420f7cf2} /* (14, 13, 2) {real, imag} */,
  {32'hc1ae301e, 32'hc185f902} /* (14, 13, 1) {real, imag} */,
  {32'h41a90ae8, 32'hc190ba7d} /* (14, 13, 0) {real, imag} */,
  {32'h41f23ff0, 32'h42089e32} /* (14, 12, 15) {real, imag} */,
  {32'hc1331ab4, 32'h420ad4d2} /* (14, 12, 14) {real, imag} */,
  {32'h40f13f18, 32'hc09f33cc} /* (14, 12, 13) {real, imag} */,
  {32'h41a50fbe, 32'h41b08493} /* (14, 12, 12) {real, imag} */,
  {32'hc202afc2, 32'h40fae49c} /* (14, 12, 11) {real, imag} */,
  {32'hbfaafb44, 32'hc186c493} /* (14, 12, 10) {real, imag} */,
  {32'hc1f55a5d, 32'hbf3ea128} /* (14, 12, 9) {real, imag} */,
  {32'h4099f8bc, 32'h4187876a} /* (14, 12, 8) {real, imag} */,
  {32'h3f1b7e30, 32'hbf5f270c} /* (14, 12, 7) {real, imag} */,
  {32'h40f50563, 32'hbf858890} /* (14, 12, 6) {real, imag} */,
  {32'hc0e34cf2, 32'h411a3e57} /* (14, 12, 5) {real, imag} */,
  {32'h410725e6, 32'hc1d6b74c} /* (14, 12, 4) {real, imag} */,
  {32'hc1a20f01, 32'hc137f3c6} /* (14, 12, 3) {real, imag} */,
  {32'h418c9ac0, 32'hbef0b4c0} /* (14, 12, 2) {real, imag} */,
  {32'hc027efd2, 32'hc18571d6} /* (14, 12, 1) {real, imag} */,
  {32'hc1afce3c, 32'hc1466486} /* (14, 12, 0) {real, imag} */,
  {32'hc13e77f2, 32'hc1def0b2} /* (14, 11, 15) {real, imag} */,
  {32'h40801816, 32'h41555824} /* (14, 11, 14) {real, imag} */,
  {32'h42224da7, 32'hc0c7ece8} /* (14, 11, 13) {real, imag} */,
  {32'h3fff7200, 32'h412db1fe} /* (14, 11, 12) {real, imag} */,
  {32'hc161a8ba, 32'hc1e94ba2} /* (14, 11, 11) {real, imag} */,
  {32'h413c401f, 32'h4183133e} /* (14, 11, 10) {real, imag} */,
  {32'h4244da24, 32'h40d220b6} /* (14, 11, 9) {real, imag} */,
  {32'hbfde2948, 32'hc0ac7360} /* (14, 11, 8) {real, imag} */,
  {32'hc12ec2d4, 32'hc0a2afc0} /* (14, 11, 7) {real, imag} */,
  {32'h420cc415, 32'hc2320fcd} /* (14, 11, 6) {real, imag} */,
  {32'h414df68c, 32'h4013dac0} /* (14, 11, 5) {real, imag} */,
  {32'h419911e9, 32'hc0642b68} /* (14, 11, 4) {real, imag} */,
  {32'hc11ecd2c, 32'hc1e692cf} /* (14, 11, 3) {real, imag} */,
  {32'h418b686a, 32'h4203445f} /* (14, 11, 2) {real, imag} */,
  {32'h419b1a32, 32'hc2155771} /* (14, 11, 1) {real, imag} */,
  {32'h41aa7f5d, 32'hc0f1f346} /* (14, 11, 0) {real, imag} */,
  {32'h422980aa, 32'h4004a1c5} /* (14, 10, 15) {real, imag} */,
  {32'hc2052362, 32'hc144f745} /* (14, 10, 14) {real, imag} */,
  {32'hc215eeae, 32'hc118f24c} /* (14, 10, 13) {real, imag} */,
  {32'h419a48c3, 32'h4215a4ea} /* (14, 10, 12) {real, imag} */,
  {32'h4145f7da, 32'h41736032} /* (14, 10, 11) {real, imag} */,
  {32'h40f6a4ab, 32'h42293815} /* (14, 10, 10) {real, imag} */,
  {32'h400edd40, 32'h3f2578a2} /* (14, 10, 9) {real, imag} */,
  {32'hc11def9c, 32'hc156ebdf} /* (14, 10, 8) {real, imag} */,
  {32'h40cca121, 32'h4214fe26} /* (14, 10, 7) {real, imag} */,
  {32'h419c79e7, 32'hc12999ab} /* (14, 10, 6) {real, imag} */,
  {32'hc1fe0522, 32'hc1532c7c} /* (14, 10, 5) {real, imag} */,
  {32'hc1066656, 32'h41c760da} /* (14, 10, 4) {real, imag} */,
  {32'h40ba823e, 32'h401d4a58} /* (14, 10, 3) {real, imag} */,
  {32'h40aec5bf, 32'hc1fba17b} /* (14, 10, 2) {real, imag} */,
  {32'hc1292d74, 32'hc1925080} /* (14, 10, 1) {real, imag} */,
  {32'h42529095, 32'h40c9f008} /* (14, 10, 0) {real, imag} */,
  {32'h40677f88, 32'h41247f02} /* (14, 9, 15) {real, imag} */,
  {32'hc12eaa80, 32'h41228f48} /* (14, 9, 14) {real, imag} */,
  {32'h410308cc, 32'h41018196} /* (14, 9, 13) {real, imag} */,
  {32'hc19ec8f0, 32'hc1ea0cfe} /* (14, 9, 12) {real, imag} */,
  {32'hc0ec4b52, 32'h4163f9ac} /* (14, 9, 11) {real, imag} */,
  {32'h411a1556, 32'h3fe8b6b8} /* (14, 9, 10) {real, imag} */,
  {32'hc1c8b037, 32'h41a363c3} /* (14, 9, 9) {real, imag} */,
  {32'h4149837f, 32'hc199daa6} /* (14, 9, 8) {real, imag} */,
  {32'h40225914, 32'h4018ef75} /* (14, 9, 7) {real, imag} */,
  {32'hbee77c00, 32'h41b00e52} /* (14, 9, 6) {real, imag} */,
  {32'hc136b240, 32'hc03aa91e} /* (14, 9, 5) {real, imag} */,
  {32'h413fef34, 32'hc16d023a} /* (14, 9, 4) {real, imag} */,
  {32'h4196c5ac, 32'hc12d9a58} /* (14, 9, 3) {real, imag} */,
  {32'h4090049a, 32'h410f6aa0} /* (14, 9, 2) {real, imag} */,
  {32'h417c3e03, 32'h41a10501} /* (14, 9, 1) {real, imag} */,
  {32'hc0a40a42, 32'hc192ae0d} /* (14, 9, 0) {real, imag} */,
  {32'hc00b2ba4, 32'hc0535c46} /* (14, 8, 15) {real, imag} */,
  {32'h3fea8306, 32'h4052eae0} /* (14, 8, 14) {real, imag} */,
  {32'hc13e2601, 32'h40c96b20} /* (14, 8, 13) {real, imag} */,
  {32'h4181ed07, 32'hc10665ce} /* (14, 8, 12) {real, imag} */,
  {32'h418f57c6, 32'h420ec0e3} /* (14, 8, 11) {real, imag} */,
  {32'hc1b86938, 32'hc132e60c} /* (14, 8, 10) {real, imag} */,
  {32'hc1bd6277, 32'h40a379f0} /* (14, 8, 9) {real, imag} */,
  {32'h414de010, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'hc1bd6277, 32'hc0a379f0} /* (14, 8, 7) {real, imag} */,
  {32'hc1b86938, 32'h4132e60c} /* (14, 8, 6) {real, imag} */,
  {32'h418f57c6, 32'hc20ec0e3} /* (14, 8, 5) {real, imag} */,
  {32'h4181ed07, 32'h410665ce} /* (14, 8, 4) {real, imag} */,
  {32'hc13e2601, 32'hc0c96b20} /* (14, 8, 3) {real, imag} */,
  {32'h3fea8306, 32'hc052eae0} /* (14, 8, 2) {real, imag} */,
  {32'hc00b2ba4, 32'h40535c46} /* (14, 8, 1) {real, imag} */,
  {32'h403dafd0, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h417c3e03, 32'hc1a10501} /* (14, 7, 15) {real, imag} */,
  {32'h4090049a, 32'hc10f6aa0} /* (14, 7, 14) {real, imag} */,
  {32'h4196c5ac, 32'h412d9a58} /* (14, 7, 13) {real, imag} */,
  {32'h413fef34, 32'h416d023a} /* (14, 7, 12) {real, imag} */,
  {32'hc136b240, 32'h403aa91e} /* (14, 7, 11) {real, imag} */,
  {32'hbee77c00, 32'hc1b00e52} /* (14, 7, 10) {real, imag} */,
  {32'h40225914, 32'hc018ef75} /* (14, 7, 9) {real, imag} */,
  {32'h4149837f, 32'h4199daa6} /* (14, 7, 8) {real, imag} */,
  {32'hc1c8b037, 32'hc1a363c3} /* (14, 7, 7) {real, imag} */,
  {32'h411a1556, 32'hbfe8b6b8} /* (14, 7, 6) {real, imag} */,
  {32'hc0ec4b52, 32'hc163f9ac} /* (14, 7, 5) {real, imag} */,
  {32'hc19ec8f0, 32'h41ea0cfe} /* (14, 7, 4) {real, imag} */,
  {32'h410308cc, 32'hc1018196} /* (14, 7, 3) {real, imag} */,
  {32'hc12eaa80, 32'hc1228f48} /* (14, 7, 2) {real, imag} */,
  {32'h40677f88, 32'hc1247f02} /* (14, 7, 1) {real, imag} */,
  {32'hc0a40a42, 32'h4192ae0d} /* (14, 7, 0) {real, imag} */,
  {32'hc1292d74, 32'h41925080} /* (14, 6, 15) {real, imag} */,
  {32'h40aec5bf, 32'h41fba17b} /* (14, 6, 14) {real, imag} */,
  {32'h40ba823e, 32'hc01d4a58} /* (14, 6, 13) {real, imag} */,
  {32'hc1066656, 32'hc1c760da} /* (14, 6, 12) {real, imag} */,
  {32'hc1fe0522, 32'h41532c7c} /* (14, 6, 11) {real, imag} */,
  {32'h419c79e7, 32'h412999ab} /* (14, 6, 10) {real, imag} */,
  {32'h40cca121, 32'hc214fe26} /* (14, 6, 9) {real, imag} */,
  {32'hc11def9c, 32'h4156ebdf} /* (14, 6, 8) {real, imag} */,
  {32'h400edd40, 32'hbf2578a2} /* (14, 6, 7) {real, imag} */,
  {32'h40f6a4ab, 32'hc2293815} /* (14, 6, 6) {real, imag} */,
  {32'h4145f7da, 32'hc1736032} /* (14, 6, 5) {real, imag} */,
  {32'h419a48c3, 32'hc215a4ea} /* (14, 6, 4) {real, imag} */,
  {32'hc215eeae, 32'h4118f24c} /* (14, 6, 3) {real, imag} */,
  {32'hc2052362, 32'h4144f745} /* (14, 6, 2) {real, imag} */,
  {32'h422980aa, 32'hc004a1c5} /* (14, 6, 1) {real, imag} */,
  {32'h42529095, 32'hc0c9f008} /* (14, 6, 0) {real, imag} */,
  {32'h419b1a32, 32'h42155771} /* (14, 5, 15) {real, imag} */,
  {32'h418b686a, 32'hc203445f} /* (14, 5, 14) {real, imag} */,
  {32'hc11ecd2c, 32'h41e692cf} /* (14, 5, 13) {real, imag} */,
  {32'h419911e9, 32'h40642b68} /* (14, 5, 12) {real, imag} */,
  {32'h414df68c, 32'hc013dac0} /* (14, 5, 11) {real, imag} */,
  {32'h420cc415, 32'h42320fcd} /* (14, 5, 10) {real, imag} */,
  {32'hc12ec2d4, 32'h40a2afc0} /* (14, 5, 9) {real, imag} */,
  {32'hbfde2948, 32'h40ac7360} /* (14, 5, 8) {real, imag} */,
  {32'h4244da24, 32'hc0d220b6} /* (14, 5, 7) {real, imag} */,
  {32'h413c401f, 32'hc183133e} /* (14, 5, 6) {real, imag} */,
  {32'hc161a8ba, 32'h41e94ba2} /* (14, 5, 5) {real, imag} */,
  {32'h3fff7200, 32'hc12db1fe} /* (14, 5, 4) {real, imag} */,
  {32'h42224da7, 32'h40c7ece8} /* (14, 5, 3) {real, imag} */,
  {32'h40801816, 32'hc1555824} /* (14, 5, 2) {real, imag} */,
  {32'hc13e77f2, 32'h41def0b2} /* (14, 5, 1) {real, imag} */,
  {32'h41aa7f5d, 32'h40f1f346} /* (14, 5, 0) {real, imag} */,
  {32'hc027efd2, 32'h418571d6} /* (14, 4, 15) {real, imag} */,
  {32'h418c9ac0, 32'h3ef0b4c0} /* (14, 4, 14) {real, imag} */,
  {32'hc1a20f01, 32'h4137f3c6} /* (14, 4, 13) {real, imag} */,
  {32'h410725e6, 32'h41d6b74c} /* (14, 4, 12) {real, imag} */,
  {32'hc0e34cf2, 32'hc11a3e57} /* (14, 4, 11) {real, imag} */,
  {32'h40f50563, 32'h3f858890} /* (14, 4, 10) {real, imag} */,
  {32'h3f1b7e30, 32'h3f5f270c} /* (14, 4, 9) {real, imag} */,
  {32'h4099f8bc, 32'hc187876a} /* (14, 4, 8) {real, imag} */,
  {32'hc1f55a5d, 32'h3f3ea128} /* (14, 4, 7) {real, imag} */,
  {32'hbfaafb44, 32'h4186c493} /* (14, 4, 6) {real, imag} */,
  {32'hc202afc2, 32'hc0fae49c} /* (14, 4, 5) {real, imag} */,
  {32'h41a50fbe, 32'hc1b08493} /* (14, 4, 4) {real, imag} */,
  {32'h40f13f18, 32'h409f33cc} /* (14, 4, 3) {real, imag} */,
  {32'hc1331ab4, 32'hc20ad4d2} /* (14, 4, 2) {real, imag} */,
  {32'h41f23ff0, 32'hc2089e32} /* (14, 4, 1) {real, imag} */,
  {32'hc1afce3c, 32'h41466486} /* (14, 4, 0) {real, imag} */,
  {32'hc1ae301e, 32'h4185f902} /* (14, 3, 15) {real, imag} */,
  {32'h4114e82a, 32'hc20f7cf2} /* (14, 3, 14) {real, imag} */,
  {32'hc28a43ca, 32'h41a21432} /* (14, 3, 13) {real, imag} */,
  {32'h424167e4, 32'h419d25c0} /* (14, 3, 12) {real, imag} */,
  {32'hc235e460, 32'hc1465688} /* (14, 3, 11) {real, imag} */,
  {32'hc1817848, 32'h425a3668} /* (14, 3, 10) {real, imag} */,
  {32'h40e39179, 32'h40a2a362} /* (14, 3, 9) {real, imag} */,
  {32'hc180871c, 32'h405c3b64} /* (14, 3, 8) {real, imag} */,
  {32'h4172af60, 32'h41248a61} /* (14, 3, 7) {real, imag} */,
  {32'hc1a6e52e, 32'hc17f6163} /* (14, 3, 6) {real, imag} */,
  {32'hc10927d3, 32'hc173c03a} /* (14, 3, 5) {real, imag} */,
  {32'hc19e5f2d, 32'h417e6cb0} /* (14, 3, 4) {real, imag} */,
  {32'hc0a06e9a, 32'h41cfd5b9} /* (14, 3, 3) {real, imag} */,
  {32'hc13bf810, 32'hc18eaccb} /* (14, 3, 2) {real, imag} */,
  {32'h41ddfc5a, 32'hc09e36f8} /* (14, 3, 1) {real, imag} */,
  {32'h41a90ae8, 32'h4190ba7d} /* (14, 3, 0) {real, imag} */,
  {32'hc2ba54d5, 32'hc282a730} /* (14, 2, 15) {real, imag} */,
  {32'hc2119f62, 32'h4207551e} /* (14, 2, 14) {real, imag} */,
  {32'h41a888e6, 32'h41d6d79a} /* (14, 2, 13) {real, imag} */,
  {32'h413b22e6, 32'hc1c5b028} /* (14, 2, 12) {real, imag} */,
  {32'hc18d42df, 32'hc19da7d6} /* (14, 2, 11) {real, imag} */,
  {32'h413b0e47, 32'hc2242a26} /* (14, 2, 10) {real, imag} */,
  {32'h41cf483b, 32'hc137fdd3} /* (14, 2, 9) {real, imag} */,
  {32'hbf7d93d8, 32'hc2037aaf} /* (14, 2, 8) {real, imag} */,
  {32'hc1a8c688, 32'h4108d2db} /* (14, 2, 7) {real, imag} */,
  {32'h41d7cdc0, 32'h41f4a6a4} /* (14, 2, 6) {real, imag} */,
  {32'hc130d24b, 32'h417bcf46} /* (14, 2, 5) {real, imag} */,
  {32'h411d3c78, 32'hc179de30} /* (14, 2, 4) {real, imag} */,
  {32'hc0a6fe22, 32'h4224434c} /* (14, 2, 3) {real, imag} */,
  {32'hc1e9589b, 32'h4099d250} /* (14, 2, 2) {real, imag} */,
  {32'h4224e501, 32'hc2238ee0} /* (14, 2, 1) {real, imag} */,
  {32'hc216de42, 32'hc143c002} /* (14, 2, 0) {real, imag} */,
  {32'hc1fc0dde, 32'hc249202c} /* (14, 1, 15) {real, imag} */,
  {32'h42506a3e, 32'hc24d2396} /* (14, 1, 14) {real, imag} */,
  {32'hc1dcb221, 32'h41b189ee} /* (14, 1, 13) {real, imag} */,
  {32'hc16a769b, 32'h41c84a6c} /* (14, 1, 12) {real, imag} */,
  {32'hbfcc0f74, 32'hc2477f2b} /* (14, 1, 11) {real, imag} */,
  {32'h412f0e14, 32'hc10f6024} /* (14, 1, 10) {real, imag} */,
  {32'h40838be9, 32'hc142a5e4} /* (14, 1, 9) {real, imag} */,
  {32'h4195c280, 32'hc0e6051e} /* (14, 1, 8) {real, imag} */,
  {32'hc0d312ac, 32'hc0dad2a6} /* (14, 1, 7) {real, imag} */,
  {32'hc1f7267a, 32'h418dbfee} /* (14, 1, 6) {real, imag} */,
  {32'h41d6c25e, 32'h4206fcc7} /* (14, 1, 5) {real, imag} */,
  {32'h406f7976, 32'hbcbb3c00} /* (14, 1, 4) {real, imag} */,
  {32'hc22d5090, 32'h41344210} /* (14, 1, 3) {real, imag} */,
  {32'hc261d021, 32'h413916f9} /* (14, 1, 2) {real, imag} */,
  {32'h42c8f3d4, 32'h42b57a14} /* (14, 1, 1) {real, imag} */,
  {32'hc2abd360, 32'hc20042b7} /* (14, 1, 0) {real, imag} */,
  {32'h4252ad32, 32'hc3278657} /* (14, 0, 15) {real, imag} */,
  {32'h420d8f4e, 32'h4222ae5b} /* (14, 0, 14) {real, imag} */,
  {32'h40cb6dd4, 32'hc20b68a2} /* (14, 0, 13) {real, imag} */,
  {32'h41d8ba9a, 32'hc1fb3483} /* (14, 0, 12) {real, imag} */,
  {32'h40f5aa16, 32'h415f75ec} /* (14, 0, 11) {real, imag} */,
  {32'h41871d5f, 32'h41ba6848} /* (14, 0, 10) {real, imag} */,
  {32'hc0cf7943, 32'h4115e72e} /* (14, 0, 9) {real, imag} */,
  {32'h419e3201, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hc0cf7943, 32'hc115e72e} /* (14, 0, 7) {real, imag} */,
  {32'h41871d5f, 32'hc1ba6848} /* (14, 0, 6) {real, imag} */,
  {32'h40f5aa16, 32'hc15f75ec} /* (14, 0, 5) {real, imag} */,
  {32'h41d8ba9a, 32'h41fb3483} /* (14, 0, 4) {real, imag} */,
  {32'h40cb6dd4, 32'h420b68a2} /* (14, 0, 3) {real, imag} */,
  {32'h420d8f4e, 32'hc222ae5b} /* (14, 0, 2) {real, imag} */,
  {32'h4252ad32, 32'h43278657} /* (14, 0, 1) {real, imag} */,
  {32'hc29944d1, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h428fafe5, 32'hc1dcad88} /* (13, 15, 15) {real, imag} */,
  {32'hc08ee950, 32'hc23b52f0} /* (13, 15, 14) {real, imag} */,
  {32'hc248ccdd, 32'hc2185719} /* (13, 15, 13) {real, imag} */,
  {32'h4209e3fe, 32'h40c4be50} /* (13, 15, 12) {real, imag} */,
  {32'h416affaa, 32'h415c09f2} /* (13, 15, 11) {real, imag} */,
  {32'h4208cb4c, 32'hc0b09cf4} /* (13, 15, 10) {real, imag} */,
  {32'hc1574d3e, 32'hc11db24d} /* (13, 15, 9) {real, imag} */,
  {32'hc12a4397, 32'h40fe67e1} /* (13, 15, 8) {real, imag} */,
  {32'h419958da, 32'h40f7b2d7} /* (13, 15, 7) {real, imag} */,
  {32'hc09e5cd8, 32'h3ef615c0} /* (13, 15, 6) {real, imag} */,
  {32'h40127980, 32'h4193ac74} /* (13, 15, 5) {real, imag} */,
  {32'h41f3bed6, 32'hc1d02176} /* (13, 15, 4) {real, imag} */,
  {32'h419f0fc0, 32'hc259fe7b} /* (13, 15, 3) {real, imag} */,
  {32'h41d8f004, 32'h42391878} /* (13, 15, 2) {real, imag} */,
  {32'h425a0300, 32'hc0fd560a} /* (13, 15, 1) {real, imag} */,
  {32'hc2670679, 32'h42c0867e} /* (13, 15, 0) {real, imag} */,
  {32'h42d46f71, 32'h41f9d95c} /* (13, 14, 15) {real, imag} */,
  {32'hc1017681, 32'hc1a83714} /* (13, 14, 14) {real, imag} */,
  {32'h3ebf9780, 32'hc1d68292} /* (13, 14, 13) {real, imag} */,
  {32'hc20999ac, 32'h422fd272} /* (13, 14, 12) {real, imag} */,
  {32'hc1a2c0d0, 32'hc0f0e30b} /* (13, 14, 11) {real, imag} */,
  {32'hc053a019, 32'hbfd806b4} /* (13, 14, 10) {real, imag} */,
  {32'h4112761a, 32'hbfa38cf0} /* (13, 14, 9) {real, imag} */,
  {32'h41343e18, 32'hc17b9855} /* (13, 14, 8) {real, imag} */,
  {32'h41871ce0, 32'hc1480cbb} /* (13, 14, 7) {real, imag} */,
  {32'hc0cbbfca, 32'h41aadb56} /* (13, 14, 6) {real, imag} */,
  {32'hc1e43f8a, 32'hc0e08752} /* (13, 14, 5) {real, imag} */,
  {32'hc027559a, 32'h4182de92} /* (13, 14, 4) {real, imag} */,
  {32'h41530160, 32'hc2405430} /* (13, 14, 3) {real, imag} */,
  {32'hc1ce5118, 32'hc15b38f7} /* (13, 14, 2) {real, imag} */,
  {32'hc27561e7, 32'h421ee8b5} /* (13, 14, 1) {real, imag} */,
  {32'hc12d848c, 32'h41e26864} /* (13, 14, 0) {real, imag} */,
  {32'h414803ac, 32'hc1b2a53f} /* (13, 13, 15) {real, imag} */,
  {32'hc13a9680, 32'h3f98719c} /* (13, 13, 14) {real, imag} */,
  {32'h41a63419, 32'hc1fe077c} /* (13, 13, 13) {real, imag} */,
  {32'hc2258271, 32'h4153d4da} /* (13, 13, 12) {real, imag} */,
  {32'h420bac19, 32'h3fc761a0} /* (13, 13, 11) {real, imag} */,
  {32'h40d04d2e, 32'hc1af25c2} /* (13, 13, 10) {real, imag} */,
  {32'h40b4deff, 32'h3f57af80} /* (13, 13, 9) {real, imag} */,
  {32'hc100e106, 32'hc177363a} /* (13, 13, 8) {real, imag} */,
  {32'hc12240db, 32'hc186d662} /* (13, 13, 7) {real, imag} */,
  {32'hc08d490f, 32'hc1d8c734} /* (13, 13, 6) {real, imag} */,
  {32'h40067d3e, 32'hc1958392} /* (13, 13, 5) {real, imag} */,
  {32'h4211cb9e, 32'hc21834e2} /* (13, 13, 4) {real, imag} */,
  {32'hc0d95c5b, 32'h41761f9b} /* (13, 13, 3) {real, imag} */,
  {32'h4200ff2b, 32'hc0c8377c} /* (13, 13, 2) {real, imag} */,
  {32'hc20f6a00, 32'hc271572b} /* (13, 13, 1) {real, imag} */,
  {32'h4216cb18, 32'hc158ea7c} /* (13, 13, 0) {real, imag} */,
  {32'hc16f6608, 32'h409f6f20} /* (13, 12, 15) {real, imag} */,
  {32'h41ff8004, 32'h4188feeb} /* (13, 12, 14) {real, imag} */,
  {32'h4192eaca, 32'hc12a49d4} /* (13, 12, 13) {real, imag} */,
  {32'hc1669d33, 32'hc18cfa53} /* (13, 12, 12) {real, imag} */,
  {32'hc048d010, 32'hbd56e800} /* (13, 12, 11) {real, imag} */,
  {32'h412e1376, 32'hc199a97f} /* (13, 12, 10) {real, imag} */,
  {32'hc1edb448, 32'hc019426f} /* (13, 12, 9) {real, imag} */,
  {32'h4118e6b8, 32'h41b09ddb} /* (13, 12, 8) {real, imag} */,
  {32'hc220825c, 32'h40c263f0} /* (13, 12, 7) {real, imag} */,
  {32'hc0807160, 32'hc167cbdd} /* (13, 12, 6) {real, imag} */,
  {32'hc23e7197, 32'h410c387c} /* (13, 12, 5) {real, imag} */,
  {32'h41c98558, 32'hc2ac317c} /* (13, 12, 4) {real, imag} */,
  {32'hc26e99d0, 32'h4235bb8e} /* (13, 12, 3) {real, imag} */,
  {32'hc216965c, 32'hc17e9604} /* (13, 12, 2) {real, imag} */,
  {32'hc071c05c, 32'h41f0b16f} /* (13, 12, 1) {real, imag} */,
  {32'h409e29f0, 32'hc109d8a7} /* (13, 12, 0) {real, imag} */,
  {32'hc1ac60b9, 32'hc16b0d8a} /* (13, 11, 15) {real, imag} */,
  {32'hc0c909b0, 32'h41ab5b38} /* (13, 11, 14) {real, imag} */,
  {32'hc1a61508, 32'h4180870d} /* (13, 11, 13) {real, imag} */,
  {32'hc0dd6a44, 32'h41558549} /* (13, 11, 12) {real, imag} */,
  {32'h423c8482, 32'hc1d703cf} /* (13, 11, 11) {real, imag} */,
  {32'hc18585fe, 32'hc0929f26} /* (13, 11, 10) {real, imag} */,
  {32'h3e7c0580, 32'hc13c716d} /* (13, 11, 9) {real, imag} */,
  {32'h4051f680, 32'h40b0b7c4} /* (13, 11, 8) {real, imag} */,
  {32'hc157c97a, 32'hc222bf78} /* (13, 11, 7) {real, imag} */,
  {32'h4218779a, 32'h416a8d16} /* (13, 11, 6) {real, imag} */,
  {32'h414962b6, 32'h4212850e} /* (13, 11, 5) {real, imag} */,
  {32'h3f767a84, 32'h41012611} /* (13, 11, 4) {real, imag} */,
  {32'h4181bfda, 32'hc1aa16e3} /* (13, 11, 3) {real, imag} */,
  {32'hc012ed3c, 32'hc0f8f2d4} /* (13, 11, 2) {real, imag} */,
  {32'hc1c00861, 32'hc0ef54ac} /* (13, 11, 1) {real, imag} */,
  {32'h421ecb77, 32'hc1f20859} /* (13, 11, 0) {real, imag} */,
  {32'h40fa9d9f, 32'hc120d8ce} /* (13, 10, 15) {real, imag} */,
  {32'h40997b9f, 32'h41fd4ea2} /* (13, 10, 14) {real, imag} */,
  {32'h40c6e34d, 32'h3fc05ab0} /* (13, 10, 13) {real, imag} */,
  {32'hbf89fd60, 32'hbf5da300} /* (13, 10, 12) {real, imag} */,
  {32'hc0a344d0, 32'h411ae1e8} /* (13, 10, 11) {real, imag} */,
  {32'h42614592, 32'hc14a522c} /* (13, 10, 10) {real, imag} */,
  {32'hc19136c6, 32'hc1a0ea50} /* (13, 10, 9) {real, imag} */,
  {32'hbfd21f12, 32'hbf06dfe8} /* (13, 10, 8) {real, imag} */,
  {32'h421cc475, 32'h420ef559} /* (13, 10, 7) {real, imag} */,
  {32'hc1a19662, 32'h4211aa68} /* (13, 10, 6) {real, imag} */,
  {32'h40fb625a, 32'hc187f808} /* (13, 10, 5) {real, imag} */,
  {32'h4207d670, 32'h416230a4} /* (13, 10, 4) {real, imag} */,
  {32'hc1de6632, 32'hc088c2e3} /* (13, 10, 3) {real, imag} */,
  {32'hc1d7b760, 32'h416d9818} /* (13, 10, 2) {real, imag} */,
  {32'hc25f0e93, 32'hc14cac9a} /* (13, 10, 1) {real, imag} */,
  {32'hc136bfa2, 32'hc1402078} /* (13, 10, 0) {real, imag} */,
  {32'h3f525128, 32'h3f70a13c} /* (13, 9, 15) {real, imag} */,
  {32'hc1b27414, 32'hc20bb4b2} /* (13, 9, 14) {real, imag} */,
  {32'hc13f75ce, 32'hc14a4cb6} /* (13, 9, 13) {real, imag} */,
  {32'hc0e085b1, 32'h414b6412} /* (13, 9, 12) {real, imag} */,
  {32'hbf29ffe0, 32'h41517917} /* (13, 9, 11) {real, imag} */,
  {32'hc05778da, 32'h41e7f086} /* (13, 9, 10) {real, imag} */,
  {32'hc1366f1a, 32'hc073cb13} /* (13, 9, 9) {real, imag} */,
  {32'h411309a7, 32'hc17fcf4f} /* (13, 9, 8) {real, imag} */,
  {32'hc2025fb5, 32'hc15e43e2} /* (13, 9, 7) {real, imag} */,
  {32'hc0451c0c, 32'hc11e33ca} /* (13, 9, 6) {real, imag} */,
  {32'hc1c6076c, 32'hbfbbb070} /* (13, 9, 5) {real, imag} */,
  {32'h4184d39c, 32'h42459f55} /* (13, 9, 4) {real, imag} */,
  {32'h40aaf49d, 32'h417b17dc} /* (13, 9, 3) {real, imag} */,
  {32'hc1787c96, 32'hc185cef9} /* (13, 9, 2) {real, imag} */,
  {32'h411a0b4a, 32'hc1cd993f} /* (13, 9, 1) {real, imag} */,
  {32'h4190e8d7, 32'h415fc01f} /* (13, 9, 0) {real, imag} */,
  {32'hc116e6a0, 32'hc12cac94} /* (13, 8, 15) {real, imag} */,
  {32'h418789d6, 32'hc191de0b} /* (13, 8, 14) {real, imag} */,
  {32'h3ffccd10, 32'h40f0c342} /* (13, 8, 13) {real, imag} */,
  {32'h3f32b318, 32'hbff8c530} /* (13, 8, 12) {real, imag} */,
  {32'h42050920, 32'h404cf250} /* (13, 8, 11) {real, imag} */,
  {32'hc18d0082, 32'h412781c7} /* (13, 8, 10) {real, imag} */,
  {32'h41388fbe, 32'h41ac9cc6} /* (13, 8, 9) {real, imag} */,
  {32'hc1985b0e, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'h41388fbe, 32'hc1ac9cc6} /* (13, 8, 7) {real, imag} */,
  {32'hc18d0082, 32'hc12781c7} /* (13, 8, 6) {real, imag} */,
  {32'h42050920, 32'hc04cf250} /* (13, 8, 5) {real, imag} */,
  {32'h3f32b318, 32'h3ff8c530} /* (13, 8, 4) {real, imag} */,
  {32'h3ffccd10, 32'hc0f0c342} /* (13, 8, 3) {real, imag} */,
  {32'h418789d6, 32'h4191de0b} /* (13, 8, 2) {real, imag} */,
  {32'hc116e6a0, 32'h412cac94} /* (13, 8, 1) {real, imag} */,
  {32'hc1308e2b, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'h411a0b4a, 32'h41cd993f} /* (13, 7, 15) {real, imag} */,
  {32'hc1787c96, 32'h4185cef9} /* (13, 7, 14) {real, imag} */,
  {32'h40aaf49d, 32'hc17b17dc} /* (13, 7, 13) {real, imag} */,
  {32'h4184d39c, 32'hc2459f55} /* (13, 7, 12) {real, imag} */,
  {32'hc1c6076c, 32'h3fbbb070} /* (13, 7, 11) {real, imag} */,
  {32'hc0451c0c, 32'h411e33ca} /* (13, 7, 10) {real, imag} */,
  {32'hc2025fb5, 32'h415e43e2} /* (13, 7, 9) {real, imag} */,
  {32'h411309a7, 32'h417fcf4f} /* (13, 7, 8) {real, imag} */,
  {32'hc1366f1a, 32'h4073cb13} /* (13, 7, 7) {real, imag} */,
  {32'hc05778da, 32'hc1e7f086} /* (13, 7, 6) {real, imag} */,
  {32'hbf29ffe0, 32'hc1517917} /* (13, 7, 5) {real, imag} */,
  {32'hc0e085b1, 32'hc14b6412} /* (13, 7, 4) {real, imag} */,
  {32'hc13f75ce, 32'h414a4cb6} /* (13, 7, 3) {real, imag} */,
  {32'hc1b27414, 32'h420bb4b2} /* (13, 7, 2) {real, imag} */,
  {32'h3f525128, 32'hbf70a13c} /* (13, 7, 1) {real, imag} */,
  {32'h4190e8d7, 32'hc15fc01f} /* (13, 7, 0) {real, imag} */,
  {32'hc25f0e93, 32'h414cac9a} /* (13, 6, 15) {real, imag} */,
  {32'hc1d7b760, 32'hc16d9818} /* (13, 6, 14) {real, imag} */,
  {32'hc1de6632, 32'h4088c2e3} /* (13, 6, 13) {real, imag} */,
  {32'h4207d670, 32'hc16230a4} /* (13, 6, 12) {real, imag} */,
  {32'h40fb625a, 32'h4187f808} /* (13, 6, 11) {real, imag} */,
  {32'hc1a19662, 32'hc211aa68} /* (13, 6, 10) {real, imag} */,
  {32'h421cc475, 32'hc20ef559} /* (13, 6, 9) {real, imag} */,
  {32'hbfd21f12, 32'h3f06dfe8} /* (13, 6, 8) {real, imag} */,
  {32'hc19136c6, 32'h41a0ea50} /* (13, 6, 7) {real, imag} */,
  {32'h42614592, 32'h414a522c} /* (13, 6, 6) {real, imag} */,
  {32'hc0a344d0, 32'hc11ae1e8} /* (13, 6, 5) {real, imag} */,
  {32'hbf89fd60, 32'h3f5da300} /* (13, 6, 4) {real, imag} */,
  {32'h40c6e34d, 32'hbfc05ab0} /* (13, 6, 3) {real, imag} */,
  {32'h40997b9f, 32'hc1fd4ea2} /* (13, 6, 2) {real, imag} */,
  {32'h40fa9d9f, 32'h4120d8ce} /* (13, 6, 1) {real, imag} */,
  {32'hc136bfa2, 32'h41402078} /* (13, 6, 0) {real, imag} */,
  {32'hc1c00861, 32'h40ef54ac} /* (13, 5, 15) {real, imag} */,
  {32'hc012ed3c, 32'h40f8f2d4} /* (13, 5, 14) {real, imag} */,
  {32'h4181bfda, 32'h41aa16e3} /* (13, 5, 13) {real, imag} */,
  {32'h3f767a84, 32'hc1012611} /* (13, 5, 12) {real, imag} */,
  {32'h414962b6, 32'hc212850e} /* (13, 5, 11) {real, imag} */,
  {32'h4218779a, 32'hc16a8d16} /* (13, 5, 10) {real, imag} */,
  {32'hc157c97a, 32'h4222bf78} /* (13, 5, 9) {real, imag} */,
  {32'h4051f680, 32'hc0b0b7c4} /* (13, 5, 8) {real, imag} */,
  {32'h3e7c0580, 32'h413c716d} /* (13, 5, 7) {real, imag} */,
  {32'hc18585fe, 32'h40929f26} /* (13, 5, 6) {real, imag} */,
  {32'h423c8482, 32'h41d703cf} /* (13, 5, 5) {real, imag} */,
  {32'hc0dd6a44, 32'hc1558549} /* (13, 5, 4) {real, imag} */,
  {32'hc1a61508, 32'hc180870d} /* (13, 5, 3) {real, imag} */,
  {32'hc0c909b0, 32'hc1ab5b38} /* (13, 5, 2) {real, imag} */,
  {32'hc1ac60b9, 32'h416b0d8a} /* (13, 5, 1) {real, imag} */,
  {32'h421ecb77, 32'h41f20859} /* (13, 5, 0) {real, imag} */,
  {32'hc071c05c, 32'hc1f0b16f} /* (13, 4, 15) {real, imag} */,
  {32'hc216965c, 32'h417e9604} /* (13, 4, 14) {real, imag} */,
  {32'hc26e99d0, 32'hc235bb8e} /* (13, 4, 13) {real, imag} */,
  {32'h41c98558, 32'h42ac317c} /* (13, 4, 12) {real, imag} */,
  {32'hc23e7197, 32'hc10c387c} /* (13, 4, 11) {real, imag} */,
  {32'hc0807160, 32'h4167cbdd} /* (13, 4, 10) {real, imag} */,
  {32'hc220825c, 32'hc0c263f0} /* (13, 4, 9) {real, imag} */,
  {32'h4118e6b8, 32'hc1b09ddb} /* (13, 4, 8) {real, imag} */,
  {32'hc1edb448, 32'h4019426f} /* (13, 4, 7) {real, imag} */,
  {32'h412e1376, 32'h4199a97f} /* (13, 4, 6) {real, imag} */,
  {32'hc048d010, 32'h3d56e800} /* (13, 4, 5) {real, imag} */,
  {32'hc1669d33, 32'h418cfa53} /* (13, 4, 4) {real, imag} */,
  {32'h4192eaca, 32'h412a49d4} /* (13, 4, 3) {real, imag} */,
  {32'h41ff8004, 32'hc188feeb} /* (13, 4, 2) {real, imag} */,
  {32'hc16f6608, 32'hc09f6f20} /* (13, 4, 1) {real, imag} */,
  {32'h409e29f0, 32'h4109d8a7} /* (13, 4, 0) {real, imag} */,
  {32'hc20f6a00, 32'h4271572b} /* (13, 3, 15) {real, imag} */,
  {32'h4200ff2b, 32'h40c8377c} /* (13, 3, 14) {real, imag} */,
  {32'hc0d95c5b, 32'hc1761f9b} /* (13, 3, 13) {real, imag} */,
  {32'h4211cb9e, 32'h421834e2} /* (13, 3, 12) {real, imag} */,
  {32'h40067d3e, 32'h41958392} /* (13, 3, 11) {real, imag} */,
  {32'hc08d490f, 32'h41d8c734} /* (13, 3, 10) {real, imag} */,
  {32'hc12240db, 32'h4186d662} /* (13, 3, 9) {real, imag} */,
  {32'hc100e106, 32'h4177363a} /* (13, 3, 8) {real, imag} */,
  {32'h40b4deff, 32'hbf57af80} /* (13, 3, 7) {real, imag} */,
  {32'h40d04d2e, 32'h41af25c2} /* (13, 3, 6) {real, imag} */,
  {32'h420bac19, 32'hbfc761a0} /* (13, 3, 5) {real, imag} */,
  {32'hc2258271, 32'hc153d4da} /* (13, 3, 4) {real, imag} */,
  {32'h41a63419, 32'h41fe077c} /* (13, 3, 3) {real, imag} */,
  {32'hc13a9680, 32'hbf98719c} /* (13, 3, 2) {real, imag} */,
  {32'h414803ac, 32'h41b2a53f} /* (13, 3, 1) {real, imag} */,
  {32'h4216cb18, 32'h4158ea7c} /* (13, 3, 0) {real, imag} */,
  {32'hc27561e7, 32'hc21ee8b5} /* (13, 2, 15) {real, imag} */,
  {32'hc1ce5118, 32'h415b38f7} /* (13, 2, 14) {real, imag} */,
  {32'h41530160, 32'h42405430} /* (13, 2, 13) {real, imag} */,
  {32'hc027559a, 32'hc182de92} /* (13, 2, 12) {real, imag} */,
  {32'hc1e43f8a, 32'h40e08752} /* (13, 2, 11) {real, imag} */,
  {32'hc0cbbfca, 32'hc1aadb56} /* (13, 2, 10) {real, imag} */,
  {32'h41871ce0, 32'h41480cbb} /* (13, 2, 9) {real, imag} */,
  {32'h41343e18, 32'h417b9855} /* (13, 2, 8) {real, imag} */,
  {32'h4112761a, 32'h3fa38cf0} /* (13, 2, 7) {real, imag} */,
  {32'hc053a019, 32'h3fd806b4} /* (13, 2, 6) {real, imag} */,
  {32'hc1a2c0d0, 32'h40f0e30b} /* (13, 2, 5) {real, imag} */,
  {32'hc20999ac, 32'hc22fd272} /* (13, 2, 4) {real, imag} */,
  {32'h3ebf9780, 32'h41d68292} /* (13, 2, 3) {real, imag} */,
  {32'hc1017681, 32'h41a83714} /* (13, 2, 2) {real, imag} */,
  {32'h42d46f71, 32'hc1f9d95c} /* (13, 2, 1) {real, imag} */,
  {32'hc12d848c, 32'hc1e26864} /* (13, 2, 0) {real, imag} */,
  {32'h425a0300, 32'h40fd560a} /* (13, 1, 15) {real, imag} */,
  {32'h41d8f004, 32'hc2391878} /* (13, 1, 14) {real, imag} */,
  {32'h419f0fc0, 32'h4259fe7b} /* (13, 1, 13) {real, imag} */,
  {32'h41f3bed6, 32'h41d02176} /* (13, 1, 12) {real, imag} */,
  {32'h40127980, 32'hc193ac74} /* (13, 1, 11) {real, imag} */,
  {32'hc09e5cd8, 32'hbef615c0} /* (13, 1, 10) {real, imag} */,
  {32'h419958da, 32'hc0f7b2d7} /* (13, 1, 9) {real, imag} */,
  {32'hc12a4397, 32'hc0fe67e1} /* (13, 1, 8) {real, imag} */,
  {32'hc1574d3e, 32'h411db24d} /* (13, 1, 7) {real, imag} */,
  {32'h4208cb4c, 32'h40b09cf4} /* (13, 1, 6) {real, imag} */,
  {32'h416affaa, 32'hc15c09f2} /* (13, 1, 5) {real, imag} */,
  {32'h4209e3fe, 32'hc0c4be50} /* (13, 1, 4) {real, imag} */,
  {32'hc248ccdd, 32'h42185719} /* (13, 1, 3) {real, imag} */,
  {32'hc08ee950, 32'h423b52f0} /* (13, 1, 2) {real, imag} */,
  {32'h428fafe5, 32'h41dcad88} /* (13, 1, 1) {real, imag} */,
  {32'hc2670679, 32'hc2c0867e} /* (13, 1, 0) {real, imag} */,
  {32'h41d0bc0d, 32'hc2eb137e} /* (13, 0, 15) {real, imag} */,
  {32'h3fefd9b8, 32'h3fd5b948} /* (13, 0, 14) {real, imag} */,
  {32'hc2304094, 32'h41f23ae6} /* (13, 0, 13) {real, imag} */,
  {32'h42559ef8, 32'hc1410614} /* (13, 0, 12) {real, imag} */,
  {32'h417d250a, 32'hc2310884} /* (13, 0, 11) {real, imag} */,
  {32'hc13be3a1, 32'h40d109eb} /* (13, 0, 10) {real, imag} */,
  {32'h410831b6, 32'h41076509} /* (13, 0, 9) {real, imag} */,
  {32'hc1e5277a, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'h410831b6, 32'hc1076509} /* (13, 0, 7) {real, imag} */,
  {32'hc13be3a1, 32'hc0d109eb} /* (13, 0, 6) {real, imag} */,
  {32'h417d250a, 32'h42310884} /* (13, 0, 5) {real, imag} */,
  {32'h42559ef8, 32'h41410614} /* (13, 0, 4) {real, imag} */,
  {32'hc2304094, 32'hc1f23ae6} /* (13, 0, 3) {real, imag} */,
  {32'h3fefd9b8, 32'hbfd5b948} /* (13, 0, 2) {real, imag} */,
  {32'h41d0bc0d, 32'h42eb137e} /* (13, 0, 1) {real, imag} */,
  {32'h4286bef4, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h41d2b181, 32'hc0e0b230} /* (12, 15, 15) {real, imag} */,
  {32'hc13f1af8, 32'hc2412362} /* (12, 15, 14) {real, imag} */,
  {32'hc1f5d4b3, 32'hc20d3255} /* (12, 15, 13) {real, imag} */,
  {32'h40a8d3a0, 32'hc118987e} /* (12, 15, 12) {real, imag} */,
  {32'hc18e5d9e, 32'h41bb2cee} /* (12, 15, 11) {real, imag} */,
  {32'h4022cbd4, 32'hc06323a0} /* (12, 15, 10) {real, imag} */,
  {32'hc1b35478, 32'h40be31f2} /* (12, 15, 9) {real, imag} */,
  {32'hc0ee72df, 32'h40c60146} /* (12, 15, 8) {real, imag} */,
  {32'hc07aae50, 32'h3fc897bc} /* (12, 15, 7) {real, imag} */,
  {32'hc151f851, 32'hbffecd74} /* (12, 15, 6) {real, imag} */,
  {32'h4091ebde, 32'h41b56bfa} /* (12, 15, 5) {real, imag} */,
  {32'h41926661, 32'h417028c2} /* (12, 15, 4) {real, imag} */,
  {32'h40ed74ea, 32'h3f8ba820} /* (12, 15, 3) {real, imag} */,
  {32'hc21f7192, 32'hbedb3d80} /* (12, 15, 2) {real, imag} */,
  {32'h4293d885, 32'hc28ffed6} /* (12, 15, 1) {real, imag} */,
  {32'hc193e6e7, 32'h418ca2de} /* (12, 15, 0) {real, imag} */,
  {32'h42da37be, 32'hc16ada95} /* (12, 14, 15) {real, imag} */,
  {32'hc1a29234, 32'h4289c010} /* (12, 14, 14) {real, imag} */,
  {32'hc2272724, 32'h41c13a30} /* (12, 14, 13) {real, imag} */,
  {32'hbf882b40, 32'hc0b93779} /* (12, 14, 12) {real, imag} */,
  {32'hc123211e, 32'h41ae4e93} /* (12, 14, 11) {real, imag} */,
  {32'h42019d9e, 32'hc11a3b0f} /* (12, 14, 10) {real, imag} */,
  {32'hc1155497, 32'hc25da01e} /* (12, 14, 9) {real, imag} */,
  {32'h3faeda00, 32'h4089ca01} /* (12, 14, 8) {real, imag} */,
  {32'h409397f0, 32'h3fd907c8} /* (12, 14, 7) {real, imag} */,
  {32'h411dec45, 32'hc1aedc21} /* (12, 14, 6) {real, imag} */,
  {32'h411aceeb, 32'hc027fc5c} /* (12, 14, 5) {real, imag} */,
  {32'hc0b9db42, 32'h40fd7230} /* (12, 14, 4) {real, imag} */,
  {32'h41f83e48, 32'hc1838ed2} /* (12, 14, 3) {real, imag} */,
  {32'h425eb883, 32'hc1b18b9a} /* (12, 14, 2) {real, imag} */,
  {32'hc2a8ca7e, 32'h4240f35e} /* (12, 14, 1) {real, imag} */,
  {32'hc28c7971, 32'h4217478f} /* (12, 14, 0) {real, imag} */,
  {32'hc07dbd10, 32'hc2126a05} /* (12, 13, 15) {real, imag} */,
  {32'hc1ca686c, 32'h418fc59e} /* (12, 13, 14) {real, imag} */,
  {32'h41a09736, 32'h400f2450} /* (12, 13, 13) {real, imag} */,
  {32'hc0f6d28c, 32'h40df04f6} /* (12, 13, 12) {real, imag} */,
  {32'hc1a07e3e, 32'hc17d5419} /* (12, 13, 11) {real, imag} */,
  {32'h41c06f66, 32'h41b357bd} /* (12, 13, 10) {real, imag} */,
  {32'h41db73ec, 32'h413c31d2} /* (12, 13, 9) {real, imag} */,
  {32'h40d6aceb, 32'h3ff683bc} /* (12, 13, 8) {real, imag} */,
  {32'h4207309a, 32'h3fb63b28} /* (12, 13, 7) {real, imag} */,
  {32'hbe7a80c0, 32'h42776474} /* (12, 13, 6) {real, imag} */,
  {32'h41790a75, 32'h416f75f2} /* (12, 13, 5) {real, imag} */,
  {32'h41f8c1c4, 32'h415a0fe4} /* (12, 13, 4) {real, imag} */,
  {32'hc204a8b1, 32'h414d73fa} /* (12, 13, 3) {real, imag} */,
  {32'hc0482df8, 32'hbfb91660} /* (12, 13, 2) {real, imag} */,
  {32'hc23921e4, 32'hc28d0470} /* (12, 13, 1) {real, imag} */,
  {32'h425131c4, 32'hc1a896d0} /* (12, 13, 0) {real, imag} */,
  {32'h41d21b84, 32'hc0b08c19} /* (12, 12, 15) {real, imag} */,
  {32'h412a4df5, 32'hbfd41ec0} /* (12, 12, 14) {real, imag} */,
  {32'h41241712, 32'hc0ffee68} /* (12, 12, 13) {real, imag} */,
  {32'hc0e5068c, 32'h408d829c} /* (12, 12, 12) {real, imag} */,
  {32'hc1db50d8, 32'h40d0ddd6} /* (12, 12, 11) {real, imag} */,
  {32'h41360a4e, 32'hc1104001} /* (12, 12, 10) {real, imag} */,
  {32'h4171df4b, 32'h42193844} /* (12, 12, 9) {real, imag} */,
  {32'h419a3b6f, 32'hc1460072} /* (12, 12, 8) {real, imag} */,
  {32'hc19757c1, 32'hc1976a4e} /* (12, 12, 7) {real, imag} */,
  {32'hc10cb708, 32'hc0ebd462} /* (12, 12, 6) {real, imag} */,
  {32'h3f9ae9f8, 32'h414720d5} /* (12, 12, 5) {real, imag} */,
  {32'h41669b2c, 32'hc2166bda} /* (12, 12, 4) {real, imag} */,
  {32'hc1a3f0f0, 32'h41e6044a} /* (12, 12, 3) {real, imag} */,
  {32'h40939cbe, 32'h400b0f08} /* (12, 12, 2) {real, imag} */,
  {32'h41a710e5, 32'h423743a4} /* (12, 12, 1) {real, imag} */,
  {32'h41169b2d, 32'hc0d80d58} /* (12, 12, 0) {real, imag} */,
  {32'hc20af50a, 32'hc1c21c5e} /* (12, 11, 15) {real, imag} */,
  {32'hc1f46584, 32'h41844c4e} /* (12, 11, 14) {real, imag} */,
  {32'hc0c69650, 32'hc20763dd} /* (12, 11, 13) {real, imag} */,
  {32'h41571980, 32'h41c26343} /* (12, 11, 12) {real, imag} */,
  {32'h40a3dd50, 32'hbf93f6e8} /* (12, 11, 11) {real, imag} */,
  {32'h420246ab, 32'h40953afa} /* (12, 11, 10) {real, imag} */,
  {32'h40ba968c, 32'hc193650d} /* (12, 11, 9) {real, imag} */,
  {32'h4190319a, 32'h40a99d9a} /* (12, 11, 8) {real, imag} */,
  {32'hc2074186, 32'hc181c9b6} /* (12, 11, 7) {real, imag} */,
  {32'hc0561ad6, 32'h41f90b8e} /* (12, 11, 6) {real, imag} */,
  {32'hc08fc9be, 32'hc1d5a3c6} /* (12, 11, 5) {real, imag} */,
  {32'h40b6c748, 32'hbf4b1920} /* (12, 11, 4) {real, imag} */,
  {32'h42511be8, 32'h40819c10} /* (12, 11, 3) {real, imag} */,
  {32'hc10eebf6, 32'h40f4e125} /* (12, 11, 2) {real, imag} */,
  {32'hc173c2e6, 32'hc15e6ec7} /* (12, 11, 1) {real, imag} */,
  {32'h41c283c8, 32'h412904db} /* (12, 11, 0) {real, imag} */,
  {32'hc1478aa1, 32'hc18156d4} /* (12, 10, 15) {real, imag} */,
  {32'h422555d3, 32'hc1a6a93c} /* (12, 10, 14) {real, imag} */,
  {32'hc193f082, 32'h403ec97c} /* (12, 10, 13) {real, imag} */,
  {32'hc13a8e2d, 32'h41c273ba} /* (12, 10, 12) {real, imag} */,
  {32'h4102700f, 32'hc148ca9b} /* (12, 10, 11) {real, imag} */,
  {32'hc1218828, 32'h412463aa} /* (12, 10, 10) {real, imag} */,
  {32'hc0370784, 32'h415166bc} /* (12, 10, 9) {real, imag} */,
  {32'h4085f615, 32'hc1600179} /* (12, 10, 8) {real, imag} */,
  {32'hc19ef7c2, 32'h4211906b} /* (12, 10, 7) {real, imag} */,
  {32'hc11fde58, 32'hc08f6e32} /* (12, 10, 6) {real, imag} */,
  {32'h418bcb95, 32'hc1d8978a} /* (12, 10, 5) {real, imag} */,
  {32'hc15efd5e, 32'h413fb7b5} /* (12, 10, 4) {real, imag} */,
  {32'hc0b47dc2, 32'h4116824e} /* (12, 10, 3) {real, imag} */,
  {32'h41296e44, 32'h404af168} /* (12, 10, 2) {real, imag} */,
  {32'h40d5be92, 32'hc1ad0f3e} /* (12, 10, 1) {real, imag} */,
  {32'h413582f1, 32'h4130f07d} /* (12, 10, 0) {real, imag} */,
  {32'h41b3f531, 32'h41372942} /* (12, 9, 15) {real, imag} */,
  {32'h419fc762, 32'h41cabc25} /* (12, 9, 14) {real, imag} */,
  {32'h40e7e9fc, 32'h41bab51b} /* (12, 9, 13) {real, imag} */,
  {32'hc0413f18, 32'hc1176eb0} /* (12, 9, 12) {real, imag} */,
  {32'h40acf320, 32'h3f9e44a4} /* (12, 9, 11) {real, imag} */,
  {32'hc24939a2, 32'hc12e50db} /* (12, 9, 10) {real, imag} */,
  {32'h411a7a07, 32'hc0cccd82} /* (12, 9, 9) {real, imag} */,
  {32'hc198a2ce, 32'h41724772} /* (12, 9, 8) {real, imag} */,
  {32'h40dbae22, 32'hc18be6da} /* (12, 9, 7) {real, imag} */,
  {32'h416ac664, 32'hc1a40f83} /* (12, 9, 6) {real, imag} */,
  {32'h3f981d8c, 32'h41bb3dcf} /* (12, 9, 5) {real, imag} */,
  {32'hc196042f, 32'hc181ee90} /* (12, 9, 4) {real, imag} */,
  {32'hc162536f, 32'hc1a29f19} /* (12, 9, 3) {real, imag} */,
  {32'hbea9f150, 32'hc0dbf630} /* (12, 9, 2) {real, imag} */,
  {32'h4104a970, 32'hc0bbfe8c} /* (12, 9, 1) {real, imag} */,
  {32'hc0d80d47, 32'hc1548660} /* (12, 9, 0) {real, imag} */,
  {32'h40e01c42, 32'h415dd5e3} /* (12, 8, 15) {real, imag} */,
  {32'h412007bf, 32'hc164fdfb} /* (12, 8, 14) {real, imag} */,
  {32'hc0fc916e, 32'hc1a2feac} /* (12, 8, 13) {real, imag} */,
  {32'h418ab6d6, 32'h401b7458} /* (12, 8, 12) {real, imag} */,
  {32'hc17dfa20, 32'h3e80a840} /* (12, 8, 11) {real, imag} */,
  {32'h404226d4, 32'h411daa67} /* (12, 8, 10) {real, imag} */,
  {32'hc092ca36, 32'h4160b944} /* (12, 8, 9) {real, imag} */,
  {32'h408c93d4, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'hc092ca36, 32'hc160b944} /* (12, 8, 7) {real, imag} */,
  {32'h404226d4, 32'hc11daa67} /* (12, 8, 6) {real, imag} */,
  {32'hc17dfa20, 32'hbe80a840} /* (12, 8, 5) {real, imag} */,
  {32'h418ab6d6, 32'hc01b7458} /* (12, 8, 4) {real, imag} */,
  {32'hc0fc916e, 32'h41a2feac} /* (12, 8, 3) {real, imag} */,
  {32'h412007bf, 32'h4164fdfb} /* (12, 8, 2) {real, imag} */,
  {32'h40e01c42, 32'hc15dd5e3} /* (12, 8, 1) {real, imag} */,
  {32'hc12af5e8, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'h4104a970, 32'h40bbfe8c} /* (12, 7, 15) {real, imag} */,
  {32'hbea9f150, 32'h40dbf630} /* (12, 7, 14) {real, imag} */,
  {32'hc162536f, 32'h41a29f19} /* (12, 7, 13) {real, imag} */,
  {32'hc196042f, 32'h4181ee90} /* (12, 7, 12) {real, imag} */,
  {32'h3f981d8c, 32'hc1bb3dcf} /* (12, 7, 11) {real, imag} */,
  {32'h416ac664, 32'h41a40f83} /* (12, 7, 10) {real, imag} */,
  {32'h40dbae22, 32'h418be6da} /* (12, 7, 9) {real, imag} */,
  {32'hc198a2ce, 32'hc1724772} /* (12, 7, 8) {real, imag} */,
  {32'h411a7a07, 32'h40cccd82} /* (12, 7, 7) {real, imag} */,
  {32'hc24939a2, 32'h412e50db} /* (12, 7, 6) {real, imag} */,
  {32'h40acf320, 32'hbf9e44a4} /* (12, 7, 5) {real, imag} */,
  {32'hc0413f18, 32'h41176eb0} /* (12, 7, 4) {real, imag} */,
  {32'h40e7e9fc, 32'hc1bab51b} /* (12, 7, 3) {real, imag} */,
  {32'h419fc762, 32'hc1cabc25} /* (12, 7, 2) {real, imag} */,
  {32'h41b3f531, 32'hc1372942} /* (12, 7, 1) {real, imag} */,
  {32'hc0d80d47, 32'h41548660} /* (12, 7, 0) {real, imag} */,
  {32'h40d5be92, 32'h41ad0f3e} /* (12, 6, 15) {real, imag} */,
  {32'h41296e44, 32'hc04af168} /* (12, 6, 14) {real, imag} */,
  {32'hc0b47dc2, 32'hc116824e} /* (12, 6, 13) {real, imag} */,
  {32'hc15efd5e, 32'hc13fb7b5} /* (12, 6, 12) {real, imag} */,
  {32'h418bcb95, 32'h41d8978a} /* (12, 6, 11) {real, imag} */,
  {32'hc11fde58, 32'h408f6e32} /* (12, 6, 10) {real, imag} */,
  {32'hc19ef7c2, 32'hc211906b} /* (12, 6, 9) {real, imag} */,
  {32'h4085f615, 32'h41600179} /* (12, 6, 8) {real, imag} */,
  {32'hc0370784, 32'hc15166bc} /* (12, 6, 7) {real, imag} */,
  {32'hc1218828, 32'hc12463aa} /* (12, 6, 6) {real, imag} */,
  {32'h4102700f, 32'h4148ca9b} /* (12, 6, 5) {real, imag} */,
  {32'hc13a8e2d, 32'hc1c273ba} /* (12, 6, 4) {real, imag} */,
  {32'hc193f082, 32'hc03ec97c} /* (12, 6, 3) {real, imag} */,
  {32'h422555d3, 32'h41a6a93c} /* (12, 6, 2) {real, imag} */,
  {32'hc1478aa1, 32'h418156d4} /* (12, 6, 1) {real, imag} */,
  {32'h413582f1, 32'hc130f07d} /* (12, 6, 0) {real, imag} */,
  {32'hc173c2e6, 32'h415e6ec7} /* (12, 5, 15) {real, imag} */,
  {32'hc10eebf6, 32'hc0f4e125} /* (12, 5, 14) {real, imag} */,
  {32'h42511be8, 32'hc0819c10} /* (12, 5, 13) {real, imag} */,
  {32'h40b6c748, 32'h3f4b1920} /* (12, 5, 12) {real, imag} */,
  {32'hc08fc9be, 32'h41d5a3c6} /* (12, 5, 11) {real, imag} */,
  {32'hc0561ad6, 32'hc1f90b8e} /* (12, 5, 10) {real, imag} */,
  {32'hc2074186, 32'h4181c9b6} /* (12, 5, 9) {real, imag} */,
  {32'h4190319a, 32'hc0a99d9a} /* (12, 5, 8) {real, imag} */,
  {32'h40ba968c, 32'h4193650d} /* (12, 5, 7) {real, imag} */,
  {32'h420246ab, 32'hc0953afa} /* (12, 5, 6) {real, imag} */,
  {32'h40a3dd50, 32'h3f93f6e8} /* (12, 5, 5) {real, imag} */,
  {32'h41571980, 32'hc1c26343} /* (12, 5, 4) {real, imag} */,
  {32'hc0c69650, 32'h420763dd} /* (12, 5, 3) {real, imag} */,
  {32'hc1f46584, 32'hc1844c4e} /* (12, 5, 2) {real, imag} */,
  {32'hc20af50a, 32'h41c21c5e} /* (12, 5, 1) {real, imag} */,
  {32'h41c283c8, 32'hc12904db} /* (12, 5, 0) {real, imag} */,
  {32'h41a710e5, 32'hc23743a4} /* (12, 4, 15) {real, imag} */,
  {32'h40939cbe, 32'hc00b0f08} /* (12, 4, 14) {real, imag} */,
  {32'hc1a3f0f0, 32'hc1e6044a} /* (12, 4, 13) {real, imag} */,
  {32'h41669b2c, 32'h42166bda} /* (12, 4, 12) {real, imag} */,
  {32'h3f9ae9f8, 32'hc14720d5} /* (12, 4, 11) {real, imag} */,
  {32'hc10cb708, 32'h40ebd462} /* (12, 4, 10) {real, imag} */,
  {32'hc19757c1, 32'h41976a4e} /* (12, 4, 9) {real, imag} */,
  {32'h419a3b6f, 32'h41460072} /* (12, 4, 8) {real, imag} */,
  {32'h4171df4b, 32'hc2193844} /* (12, 4, 7) {real, imag} */,
  {32'h41360a4e, 32'h41104001} /* (12, 4, 6) {real, imag} */,
  {32'hc1db50d8, 32'hc0d0ddd6} /* (12, 4, 5) {real, imag} */,
  {32'hc0e5068c, 32'hc08d829c} /* (12, 4, 4) {real, imag} */,
  {32'h41241712, 32'h40ffee68} /* (12, 4, 3) {real, imag} */,
  {32'h412a4df5, 32'h3fd41ec0} /* (12, 4, 2) {real, imag} */,
  {32'h41d21b84, 32'h40b08c19} /* (12, 4, 1) {real, imag} */,
  {32'h41169b2d, 32'h40d80d58} /* (12, 4, 0) {real, imag} */,
  {32'hc23921e4, 32'h428d0470} /* (12, 3, 15) {real, imag} */,
  {32'hc0482df8, 32'h3fb91660} /* (12, 3, 14) {real, imag} */,
  {32'hc204a8b1, 32'hc14d73fa} /* (12, 3, 13) {real, imag} */,
  {32'h41f8c1c4, 32'hc15a0fe4} /* (12, 3, 12) {real, imag} */,
  {32'h41790a75, 32'hc16f75f2} /* (12, 3, 11) {real, imag} */,
  {32'hbe7a80c0, 32'hc2776474} /* (12, 3, 10) {real, imag} */,
  {32'h4207309a, 32'hbfb63b28} /* (12, 3, 9) {real, imag} */,
  {32'h40d6aceb, 32'hbff683bc} /* (12, 3, 8) {real, imag} */,
  {32'h41db73ec, 32'hc13c31d2} /* (12, 3, 7) {real, imag} */,
  {32'h41c06f66, 32'hc1b357bd} /* (12, 3, 6) {real, imag} */,
  {32'hc1a07e3e, 32'h417d5419} /* (12, 3, 5) {real, imag} */,
  {32'hc0f6d28c, 32'hc0df04f6} /* (12, 3, 4) {real, imag} */,
  {32'h41a09736, 32'hc00f2450} /* (12, 3, 3) {real, imag} */,
  {32'hc1ca686c, 32'hc18fc59e} /* (12, 3, 2) {real, imag} */,
  {32'hc07dbd10, 32'h42126a05} /* (12, 3, 1) {real, imag} */,
  {32'h425131c4, 32'h41a896d0} /* (12, 3, 0) {real, imag} */,
  {32'hc2a8ca7e, 32'hc240f35e} /* (12, 2, 15) {real, imag} */,
  {32'h425eb883, 32'h41b18b9a} /* (12, 2, 14) {real, imag} */,
  {32'h41f83e48, 32'h41838ed2} /* (12, 2, 13) {real, imag} */,
  {32'hc0b9db42, 32'hc0fd7230} /* (12, 2, 12) {real, imag} */,
  {32'h411aceeb, 32'h4027fc5c} /* (12, 2, 11) {real, imag} */,
  {32'h411dec45, 32'h41aedc21} /* (12, 2, 10) {real, imag} */,
  {32'h409397f0, 32'hbfd907c8} /* (12, 2, 9) {real, imag} */,
  {32'h3faeda00, 32'hc089ca01} /* (12, 2, 8) {real, imag} */,
  {32'hc1155497, 32'h425da01e} /* (12, 2, 7) {real, imag} */,
  {32'h42019d9e, 32'h411a3b0f} /* (12, 2, 6) {real, imag} */,
  {32'hc123211e, 32'hc1ae4e93} /* (12, 2, 5) {real, imag} */,
  {32'hbf882b40, 32'h40b93779} /* (12, 2, 4) {real, imag} */,
  {32'hc2272724, 32'hc1c13a30} /* (12, 2, 3) {real, imag} */,
  {32'hc1a29234, 32'hc289c010} /* (12, 2, 2) {real, imag} */,
  {32'h42da37be, 32'h416ada95} /* (12, 2, 1) {real, imag} */,
  {32'hc28c7971, 32'hc217478f} /* (12, 2, 0) {real, imag} */,
  {32'h4293d885, 32'h428ffed6} /* (12, 1, 15) {real, imag} */,
  {32'hc21f7192, 32'h3edb3d80} /* (12, 1, 14) {real, imag} */,
  {32'h40ed74ea, 32'hbf8ba820} /* (12, 1, 13) {real, imag} */,
  {32'h41926661, 32'hc17028c2} /* (12, 1, 12) {real, imag} */,
  {32'h4091ebde, 32'hc1b56bfa} /* (12, 1, 11) {real, imag} */,
  {32'hc151f851, 32'h3ffecd74} /* (12, 1, 10) {real, imag} */,
  {32'hc07aae50, 32'hbfc897bc} /* (12, 1, 9) {real, imag} */,
  {32'hc0ee72df, 32'hc0c60146} /* (12, 1, 8) {real, imag} */,
  {32'hc1b35478, 32'hc0be31f2} /* (12, 1, 7) {real, imag} */,
  {32'h4022cbd4, 32'h406323a0} /* (12, 1, 6) {real, imag} */,
  {32'hc18e5d9e, 32'hc1bb2cee} /* (12, 1, 5) {real, imag} */,
  {32'h40a8d3a0, 32'h4118987e} /* (12, 1, 4) {real, imag} */,
  {32'hc1f5d4b3, 32'h420d3255} /* (12, 1, 3) {real, imag} */,
  {32'hc13f1af8, 32'h42412362} /* (12, 1, 2) {real, imag} */,
  {32'h41d2b181, 32'h40e0b230} /* (12, 1, 1) {real, imag} */,
  {32'hc193e6e7, 32'hc18ca2de} /* (12, 1, 0) {real, imag} */,
  {32'hc1b25aa2, 32'hc1e82d47} /* (12, 0, 15) {real, imag} */,
  {32'h4051b3e8, 32'hbfc58040} /* (12, 0, 14) {real, imag} */,
  {32'h41094b84, 32'h41df23c3} /* (12, 0, 13) {real, imag} */,
  {32'h41801930, 32'hc2157078} /* (12, 0, 12) {real, imag} */,
  {32'h4199dfe1, 32'hc00c060c} /* (12, 0, 11) {real, imag} */,
  {32'hc1cd4eeb, 32'h41bb4aff} /* (12, 0, 10) {real, imag} */,
  {32'h413965bd, 32'hc1ae9524} /* (12, 0, 9) {real, imag} */,
  {32'hc180b5e0, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'h413965bd, 32'h41ae9524} /* (12, 0, 7) {real, imag} */,
  {32'hc1cd4eeb, 32'hc1bb4aff} /* (12, 0, 6) {real, imag} */,
  {32'h4199dfe1, 32'h400c060c} /* (12, 0, 5) {real, imag} */,
  {32'h41801930, 32'h42157078} /* (12, 0, 4) {real, imag} */,
  {32'h41094b84, 32'hc1df23c3} /* (12, 0, 3) {real, imag} */,
  {32'h4051b3e8, 32'h3fc58040} /* (12, 0, 2) {real, imag} */,
  {32'hc1b25aa2, 32'h41e82d47} /* (12, 0, 1) {real, imag} */,
  {32'h431d99a3, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h3fd074f0, 32'h402abea0} /* (11, 15, 15) {real, imag} */,
  {32'hc23cb9ee, 32'h408a750a} /* (11, 15, 14) {real, imag} */,
  {32'h419f35b6, 32'hc273b61d} /* (11, 15, 13) {real, imag} */,
  {32'h41ce0614, 32'hc08eac00} /* (11, 15, 12) {real, imag} */,
  {32'h42822663, 32'h4127b64a} /* (11, 15, 11) {real, imag} */,
  {32'hc0de508c, 32'h411c9832} /* (11, 15, 10) {real, imag} */,
  {32'hc109069d, 32'hc12ff7b6} /* (11, 15, 9) {real, imag} */,
  {32'h4124ea68, 32'h4073ab56} /* (11, 15, 8) {real, imag} */,
  {32'hc1a67997, 32'h40981aaf} /* (11, 15, 7) {real, imag} */,
  {32'h418a3d00, 32'h42072e82} /* (11, 15, 6) {real, imag} */,
  {32'hc0d4c1a0, 32'h3f9bf378} /* (11, 15, 5) {real, imag} */,
  {32'hc1d177b8, 32'hc11e5ba4} /* (11, 15, 4) {real, imag} */,
  {32'h3fd61680, 32'hc1ec7e0e} /* (11, 15, 3) {real, imag} */,
  {32'hc222e978, 32'h42210b3c} /* (11, 15, 2) {real, imag} */,
  {32'h419bbd30, 32'hc2044f91} /* (11, 15, 1) {real, imag} */,
  {32'hc250e90e, 32'hc2d4e4ce} /* (11, 15, 0) {real, imag} */,
  {32'h41930774, 32'hc2420acf} /* (11, 14, 15) {real, imag} */,
  {32'hc224a756, 32'h415966da} /* (11, 14, 14) {real, imag} */,
  {32'hc153f638, 32'h405a764c} /* (11, 14, 13) {real, imag} */,
  {32'hc1949009, 32'h4187dcbb} /* (11, 14, 12) {real, imag} */,
  {32'hc1cd331d, 32'hc12d7778} /* (11, 14, 11) {real, imag} */,
  {32'h418698f4, 32'h4038bd12} /* (11, 14, 10) {real, imag} */,
  {32'hc137ff8c, 32'hc1dbb188} /* (11, 14, 9) {real, imag} */,
  {32'h3fafc960, 32'h410a7555} /* (11, 14, 8) {real, imag} */,
  {32'h3f7ce0a0, 32'hc1bd2ea6} /* (11, 14, 7) {real, imag} */,
  {32'hc1dfd2be, 32'h413b0ad6} /* (11, 14, 6) {real, imag} */,
  {32'h40a46db8, 32'hc18139d0} /* (11, 14, 5) {real, imag} */,
  {32'hc110b978, 32'h40a8f38c} /* (11, 14, 4) {real, imag} */,
  {32'h423ea443, 32'h422e82d8} /* (11, 14, 3) {real, imag} */,
  {32'h42015d27, 32'hbee38a00} /* (11, 14, 2) {real, imag} */,
  {32'h411d223a, 32'h428fc77b} /* (11, 14, 1) {real, imag} */,
  {32'hc280de48, 32'hc1053b24} /* (11, 14, 0) {real, imag} */,
  {32'h41b4a314, 32'hc0341fe0} /* (11, 13, 15) {real, imag} */,
  {32'hc109a900, 32'h40641dd0} /* (11, 13, 14) {real, imag} */,
  {32'hc1d8268a, 32'h420c580e} /* (11, 13, 13) {real, imag} */,
  {32'h41bb96de, 32'h41e724e2} /* (11, 13, 12) {real, imag} */,
  {32'h418954b2, 32'hbf7b3140} /* (11, 13, 11) {real, imag} */,
  {32'hc162230f, 32'h400f2034} /* (11, 13, 10) {real, imag} */,
  {32'h41a34a45, 32'h3f992188} /* (11, 13, 9) {real, imag} */,
  {32'h41851599, 32'h4180b829} /* (11, 13, 8) {real, imag} */,
  {32'h403cac4b, 32'h40abae0e} /* (11, 13, 7) {real, imag} */,
  {32'hc171372e, 32'h41cc98a1} /* (11, 13, 6) {real, imag} */,
  {32'h41444831, 32'h4197e530} /* (11, 13, 5) {real, imag} */,
  {32'h40d9eeb0, 32'hc1196d6b} /* (11, 13, 4) {real, imag} */,
  {32'hc0e4df63, 32'hc0e2cf42} /* (11, 13, 3) {real, imag} */,
  {32'h4134f660, 32'h4120b304} /* (11, 13, 2) {real, imag} */,
  {32'hc2269ace, 32'hc28637a2} /* (11, 13, 1) {real, imag} */,
  {32'h428cee1a, 32'hc1d6d452} /* (11, 13, 0) {real, imag} */,
  {32'h4238b030, 32'hc1dc48b2} /* (11, 12, 15) {real, imag} */,
  {32'h41de7637, 32'h424f0b14} /* (11, 12, 14) {real, imag} */,
  {32'h4165fd15, 32'hc25100ca} /* (11, 12, 13) {real, imag} */,
  {32'hc1142578, 32'h41d1a3c3} /* (11, 12, 12) {real, imag} */,
  {32'hc2590628, 32'h41e03f26} /* (11, 12, 11) {real, imag} */,
  {32'hbf40db80, 32'hc1f339f4} /* (11, 12, 10) {real, imag} */,
  {32'hbeb46460, 32'h410a383e} /* (11, 12, 9) {real, imag} */,
  {32'h41eab7a4, 32'h3f91ce7c} /* (11, 12, 8) {real, imag} */,
  {32'hc1857508, 32'h414ea6c6} /* (11, 12, 7) {real, imag} */,
  {32'hc1fca4c2, 32'hc1d44bec} /* (11, 12, 6) {real, imag} */,
  {32'h41dd6a86, 32'hc159f28e} /* (11, 12, 5) {real, imag} */,
  {32'h41f0b900, 32'h408d96f8} /* (11, 12, 4) {real, imag} */,
  {32'hc0e5f198, 32'hc15d11f5} /* (11, 12, 3) {real, imag} */,
  {32'h407721a0, 32'h4112782f} /* (11, 12, 2) {real, imag} */,
  {32'h420d4207, 32'hc2267c72} /* (11, 12, 1) {real, imag} */,
  {32'hc19d6a3a, 32'h424ac55c} /* (11, 12, 0) {real, imag} */,
  {32'hc216e064, 32'h41a81c58} /* (11, 11, 15) {real, imag} */,
  {32'h4219a53f, 32'h4195d5ed} /* (11, 11, 14) {real, imag} */,
  {32'hc0c62d72, 32'h40a172ec} /* (11, 11, 13) {real, imag} */,
  {32'hc15977b0, 32'hc237e795} /* (11, 11, 12) {real, imag} */,
  {32'hc19ed70d, 32'hc1095dca} /* (11, 11, 11) {real, imag} */,
  {32'h40d91a74, 32'hc105a3ee} /* (11, 11, 10) {real, imag} */,
  {32'h4168cb94, 32'h423e6b96} /* (11, 11, 9) {real, imag} */,
  {32'h417c5861, 32'h410477ee} /* (11, 11, 8) {real, imag} */,
  {32'h41f9b109, 32'hc105a838} /* (11, 11, 7) {real, imag} */,
  {32'hc0d30734, 32'h3fa51cc8} /* (11, 11, 6) {real, imag} */,
  {32'h40c74ea0, 32'hc1dbfdf3} /* (11, 11, 5) {real, imag} */,
  {32'h415f24a0, 32'hc1071921} /* (11, 11, 4) {real, imag} */,
  {32'hc280e512, 32'hc1b25985} /* (11, 11, 3) {real, imag} */,
  {32'hc10a9b76, 32'h40431348} /* (11, 11, 2) {real, imag} */,
  {32'h41c4ef1e, 32'hc11ed4d4} /* (11, 11, 1) {real, imag} */,
  {32'h41254604, 32'h42118d3c} /* (11, 11, 0) {real, imag} */,
  {32'h41184650, 32'h40cfed42} /* (11, 10, 15) {real, imag} */,
  {32'h419470f5, 32'hc1bef237} /* (11, 10, 14) {real, imag} */,
  {32'hc1e97d57, 32'hc0e8e080} /* (11, 10, 13) {real, imag} */,
  {32'hc13ce15a, 32'h4190c3b8} /* (11, 10, 12) {real, imag} */,
  {32'h41b0b6c3, 32'h416bebc7} /* (11, 10, 11) {real, imag} */,
  {32'h41fdefde, 32'h41656396} /* (11, 10, 10) {real, imag} */,
  {32'h41f11311, 32'hc1dc9bdb} /* (11, 10, 9) {real, imag} */,
  {32'hc17db8c6, 32'hc1d1cade} /* (11, 10, 8) {real, imag} */,
  {32'h4183ff9c, 32'h418acbfe} /* (11, 10, 7) {real, imag} */,
  {32'h40baeb1e, 32'h42453036} /* (11, 10, 6) {real, imag} */,
  {32'hc1f8a3ca, 32'h419ee23e} /* (11, 10, 5) {real, imag} */,
  {32'hc1c2dfdf, 32'hc2244ff6} /* (11, 10, 4) {real, imag} */,
  {32'hc14fbcc4, 32'hbe9f10b0} /* (11, 10, 3) {real, imag} */,
  {32'h418d6158, 32'h4123ad7c} /* (11, 10, 2) {real, imag} */,
  {32'hc14783ac, 32'hc0d4c564} /* (11, 10, 1) {real, imag} */,
  {32'hc12f6b98, 32'h411adf44} /* (11, 10, 0) {real, imag} */,
  {32'hc18e5ace, 32'h414e9516} /* (11, 9, 15) {real, imag} */,
  {32'hc1211449, 32'h419f6621} /* (11, 9, 14) {real, imag} */,
  {32'h41860920, 32'h41923a4e} /* (11, 9, 13) {real, imag} */,
  {32'h4155fbf0, 32'hc19e8e8f} /* (11, 9, 12) {real, imag} */,
  {32'h40c8242c, 32'hc1698dd4} /* (11, 9, 11) {real, imag} */,
  {32'h41c7550f, 32'hc0bf0468} /* (11, 9, 10) {real, imag} */,
  {32'hc18fb764, 32'hc02d881d} /* (11, 9, 9) {real, imag} */,
  {32'h4192de36, 32'h410918fc} /* (11, 9, 8) {real, imag} */,
  {32'h3fcc0560, 32'h413d7cbb} /* (11, 9, 7) {real, imag} */,
  {32'hc19db550, 32'hc04ce5f6} /* (11, 9, 6) {real, imag} */,
  {32'hc172d946, 32'h40958a24} /* (11, 9, 5) {real, imag} */,
  {32'hc10237e0, 32'h41f8f275} /* (11, 9, 4) {real, imag} */,
  {32'h3ffff2da, 32'hc13d9ced} /* (11, 9, 3) {real, imag} */,
  {32'h41a0105d, 32'hc2419430} /* (11, 9, 2) {real, imag} */,
  {32'h41a23e16, 32'h4093252a} /* (11, 9, 1) {real, imag} */,
  {32'hc165d144, 32'h4144c850} /* (11, 9, 0) {real, imag} */,
  {32'hc0e4a370, 32'hc13f6f2c} /* (11, 8, 15) {real, imag} */,
  {32'h3f06b6a0, 32'hc0772680} /* (11, 8, 14) {real, imag} */,
  {32'h409b17e1, 32'h3f03bbc0} /* (11, 8, 13) {real, imag} */,
  {32'h405c2898, 32'h3ff34efc} /* (11, 8, 12) {real, imag} */,
  {32'h415a2b28, 32'hc1276e22} /* (11, 8, 11) {real, imag} */,
  {32'h417835e5, 32'hc15ef31f} /* (11, 8, 10) {real, imag} */,
  {32'h40877360, 32'hc16b2aba} /* (11, 8, 9) {real, imag} */,
  {32'hc16de6aa, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'h40877360, 32'h416b2aba} /* (11, 8, 7) {real, imag} */,
  {32'h417835e5, 32'h415ef31f} /* (11, 8, 6) {real, imag} */,
  {32'h415a2b28, 32'h41276e22} /* (11, 8, 5) {real, imag} */,
  {32'h405c2898, 32'hbff34efc} /* (11, 8, 4) {real, imag} */,
  {32'h409b17e1, 32'hbf03bbc0} /* (11, 8, 3) {real, imag} */,
  {32'h3f06b6a0, 32'h40772680} /* (11, 8, 2) {real, imag} */,
  {32'hc0e4a370, 32'h413f6f2c} /* (11, 8, 1) {real, imag} */,
  {32'hc0f797d7, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h41a23e16, 32'hc093252a} /* (11, 7, 15) {real, imag} */,
  {32'h41a0105d, 32'h42419430} /* (11, 7, 14) {real, imag} */,
  {32'h3ffff2da, 32'h413d9ced} /* (11, 7, 13) {real, imag} */,
  {32'hc10237e0, 32'hc1f8f275} /* (11, 7, 12) {real, imag} */,
  {32'hc172d946, 32'hc0958a24} /* (11, 7, 11) {real, imag} */,
  {32'hc19db550, 32'h404ce5f6} /* (11, 7, 10) {real, imag} */,
  {32'h3fcc0560, 32'hc13d7cbb} /* (11, 7, 9) {real, imag} */,
  {32'h4192de36, 32'hc10918fc} /* (11, 7, 8) {real, imag} */,
  {32'hc18fb764, 32'h402d881d} /* (11, 7, 7) {real, imag} */,
  {32'h41c7550f, 32'h40bf0468} /* (11, 7, 6) {real, imag} */,
  {32'h40c8242c, 32'h41698dd4} /* (11, 7, 5) {real, imag} */,
  {32'h4155fbf0, 32'h419e8e8f} /* (11, 7, 4) {real, imag} */,
  {32'h41860920, 32'hc1923a4e} /* (11, 7, 3) {real, imag} */,
  {32'hc1211449, 32'hc19f6621} /* (11, 7, 2) {real, imag} */,
  {32'hc18e5ace, 32'hc14e9516} /* (11, 7, 1) {real, imag} */,
  {32'hc165d144, 32'hc144c850} /* (11, 7, 0) {real, imag} */,
  {32'hc14783ac, 32'h40d4c564} /* (11, 6, 15) {real, imag} */,
  {32'h418d6158, 32'hc123ad7c} /* (11, 6, 14) {real, imag} */,
  {32'hc14fbcc4, 32'h3e9f10b0} /* (11, 6, 13) {real, imag} */,
  {32'hc1c2dfdf, 32'h42244ff6} /* (11, 6, 12) {real, imag} */,
  {32'hc1f8a3ca, 32'hc19ee23e} /* (11, 6, 11) {real, imag} */,
  {32'h40baeb1e, 32'hc2453036} /* (11, 6, 10) {real, imag} */,
  {32'h4183ff9c, 32'hc18acbfe} /* (11, 6, 9) {real, imag} */,
  {32'hc17db8c6, 32'h41d1cade} /* (11, 6, 8) {real, imag} */,
  {32'h41f11311, 32'h41dc9bdb} /* (11, 6, 7) {real, imag} */,
  {32'h41fdefde, 32'hc1656396} /* (11, 6, 6) {real, imag} */,
  {32'h41b0b6c3, 32'hc16bebc7} /* (11, 6, 5) {real, imag} */,
  {32'hc13ce15a, 32'hc190c3b8} /* (11, 6, 4) {real, imag} */,
  {32'hc1e97d57, 32'h40e8e080} /* (11, 6, 3) {real, imag} */,
  {32'h419470f5, 32'h41bef237} /* (11, 6, 2) {real, imag} */,
  {32'h41184650, 32'hc0cfed42} /* (11, 6, 1) {real, imag} */,
  {32'hc12f6b98, 32'hc11adf44} /* (11, 6, 0) {real, imag} */,
  {32'h41c4ef1e, 32'h411ed4d4} /* (11, 5, 15) {real, imag} */,
  {32'hc10a9b76, 32'hc0431348} /* (11, 5, 14) {real, imag} */,
  {32'hc280e512, 32'h41b25985} /* (11, 5, 13) {real, imag} */,
  {32'h415f24a0, 32'h41071921} /* (11, 5, 12) {real, imag} */,
  {32'h40c74ea0, 32'h41dbfdf3} /* (11, 5, 11) {real, imag} */,
  {32'hc0d30734, 32'hbfa51cc8} /* (11, 5, 10) {real, imag} */,
  {32'h41f9b109, 32'h4105a838} /* (11, 5, 9) {real, imag} */,
  {32'h417c5861, 32'hc10477ee} /* (11, 5, 8) {real, imag} */,
  {32'h4168cb94, 32'hc23e6b96} /* (11, 5, 7) {real, imag} */,
  {32'h40d91a74, 32'h4105a3ee} /* (11, 5, 6) {real, imag} */,
  {32'hc19ed70d, 32'h41095dca} /* (11, 5, 5) {real, imag} */,
  {32'hc15977b0, 32'h4237e795} /* (11, 5, 4) {real, imag} */,
  {32'hc0c62d72, 32'hc0a172ec} /* (11, 5, 3) {real, imag} */,
  {32'h4219a53f, 32'hc195d5ed} /* (11, 5, 2) {real, imag} */,
  {32'hc216e064, 32'hc1a81c58} /* (11, 5, 1) {real, imag} */,
  {32'h41254604, 32'hc2118d3c} /* (11, 5, 0) {real, imag} */,
  {32'h420d4207, 32'h42267c72} /* (11, 4, 15) {real, imag} */,
  {32'h407721a0, 32'hc112782f} /* (11, 4, 14) {real, imag} */,
  {32'hc0e5f198, 32'h415d11f5} /* (11, 4, 13) {real, imag} */,
  {32'h41f0b900, 32'hc08d96f8} /* (11, 4, 12) {real, imag} */,
  {32'h41dd6a86, 32'h4159f28e} /* (11, 4, 11) {real, imag} */,
  {32'hc1fca4c2, 32'h41d44bec} /* (11, 4, 10) {real, imag} */,
  {32'hc1857508, 32'hc14ea6c6} /* (11, 4, 9) {real, imag} */,
  {32'h41eab7a4, 32'hbf91ce7c} /* (11, 4, 8) {real, imag} */,
  {32'hbeb46460, 32'hc10a383e} /* (11, 4, 7) {real, imag} */,
  {32'hbf40db80, 32'h41f339f4} /* (11, 4, 6) {real, imag} */,
  {32'hc2590628, 32'hc1e03f26} /* (11, 4, 5) {real, imag} */,
  {32'hc1142578, 32'hc1d1a3c3} /* (11, 4, 4) {real, imag} */,
  {32'h4165fd15, 32'h425100ca} /* (11, 4, 3) {real, imag} */,
  {32'h41de7637, 32'hc24f0b14} /* (11, 4, 2) {real, imag} */,
  {32'h4238b030, 32'h41dc48b2} /* (11, 4, 1) {real, imag} */,
  {32'hc19d6a3a, 32'hc24ac55c} /* (11, 4, 0) {real, imag} */,
  {32'hc2269ace, 32'h428637a2} /* (11, 3, 15) {real, imag} */,
  {32'h4134f660, 32'hc120b304} /* (11, 3, 14) {real, imag} */,
  {32'hc0e4df63, 32'h40e2cf42} /* (11, 3, 13) {real, imag} */,
  {32'h40d9eeb0, 32'h41196d6b} /* (11, 3, 12) {real, imag} */,
  {32'h41444831, 32'hc197e530} /* (11, 3, 11) {real, imag} */,
  {32'hc171372e, 32'hc1cc98a1} /* (11, 3, 10) {real, imag} */,
  {32'h403cac4b, 32'hc0abae0e} /* (11, 3, 9) {real, imag} */,
  {32'h41851599, 32'hc180b829} /* (11, 3, 8) {real, imag} */,
  {32'h41a34a45, 32'hbf992188} /* (11, 3, 7) {real, imag} */,
  {32'hc162230f, 32'hc00f2034} /* (11, 3, 6) {real, imag} */,
  {32'h418954b2, 32'h3f7b3140} /* (11, 3, 5) {real, imag} */,
  {32'h41bb96de, 32'hc1e724e2} /* (11, 3, 4) {real, imag} */,
  {32'hc1d8268a, 32'hc20c580e} /* (11, 3, 3) {real, imag} */,
  {32'hc109a900, 32'hc0641dd0} /* (11, 3, 2) {real, imag} */,
  {32'h41b4a314, 32'h40341fe0} /* (11, 3, 1) {real, imag} */,
  {32'h428cee1a, 32'h41d6d452} /* (11, 3, 0) {real, imag} */,
  {32'h411d223a, 32'hc28fc77b} /* (11, 2, 15) {real, imag} */,
  {32'h42015d27, 32'h3ee38a00} /* (11, 2, 14) {real, imag} */,
  {32'h423ea443, 32'hc22e82d8} /* (11, 2, 13) {real, imag} */,
  {32'hc110b978, 32'hc0a8f38c} /* (11, 2, 12) {real, imag} */,
  {32'h40a46db8, 32'h418139d0} /* (11, 2, 11) {real, imag} */,
  {32'hc1dfd2be, 32'hc13b0ad6} /* (11, 2, 10) {real, imag} */,
  {32'h3f7ce0a0, 32'h41bd2ea6} /* (11, 2, 9) {real, imag} */,
  {32'h3fafc960, 32'hc10a7555} /* (11, 2, 8) {real, imag} */,
  {32'hc137ff8c, 32'h41dbb188} /* (11, 2, 7) {real, imag} */,
  {32'h418698f4, 32'hc038bd12} /* (11, 2, 6) {real, imag} */,
  {32'hc1cd331d, 32'h412d7778} /* (11, 2, 5) {real, imag} */,
  {32'hc1949009, 32'hc187dcbb} /* (11, 2, 4) {real, imag} */,
  {32'hc153f638, 32'hc05a764c} /* (11, 2, 3) {real, imag} */,
  {32'hc224a756, 32'hc15966da} /* (11, 2, 2) {real, imag} */,
  {32'h41930774, 32'h42420acf} /* (11, 2, 1) {real, imag} */,
  {32'hc280de48, 32'h41053b24} /* (11, 2, 0) {real, imag} */,
  {32'h419bbd30, 32'h42044f91} /* (11, 1, 15) {real, imag} */,
  {32'hc222e978, 32'hc2210b3c} /* (11, 1, 14) {real, imag} */,
  {32'h3fd61680, 32'h41ec7e0e} /* (11, 1, 13) {real, imag} */,
  {32'hc1d177b8, 32'h411e5ba4} /* (11, 1, 12) {real, imag} */,
  {32'hc0d4c1a0, 32'hbf9bf378} /* (11, 1, 11) {real, imag} */,
  {32'h418a3d00, 32'hc2072e82} /* (11, 1, 10) {real, imag} */,
  {32'hc1a67997, 32'hc0981aaf} /* (11, 1, 9) {real, imag} */,
  {32'h4124ea68, 32'hc073ab56} /* (11, 1, 8) {real, imag} */,
  {32'hc109069d, 32'h412ff7b6} /* (11, 1, 7) {real, imag} */,
  {32'hc0de508c, 32'hc11c9832} /* (11, 1, 6) {real, imag} */,
  {32'h42822663, 32'hc127b64a} /* (11, 1, 5) {real, imag} */,
  {32'h41ce0614, 32'h408eac00} /* (11, 1, 4) {real, imag} */,
  {32'h419f35b6, 32'h4273b61d} /* (11, 1, 3) {real, imag} */,
  {32'hc23cb9ee, 32'hc08a750a} /* (11, 1, 2) {real, imag} */,
  {32'h3fd074f0, 32'hc02abea0} /* (11, 1, 1) {real, imag} */,
  {32'hc250e90e, 32'h42d4e4ce} /* (11, 1, 0) {real, imag} */,
  {32'hc0ca1a00, 32'h42868a2a} /* (11, 0, 15) {real, imag} */,
  {32'h42254019, 32'hc17256ac} /* (11, 0, 14) {real, imag} */,
  {32'h412970a8, 32'hc0009420} /* (11, 0, 13) {real, imag} */,
  {32'h40ffd994, 32'hc29fb157} /* (11, 0, 12) {real, imag} */,
  {32'h41a1f135, 32'h4272a7b7} /* (11, 0, 11) {real, imag} */,
  {32'hc227078d, 32'h41e16db4} /* (11, 0, 10) {real, imag} */,
  {32'h42071d1f, 32'hc0ed3016} /* (11, 0, 9) {real, imag} */,
  {32'hc244283d, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'h42071d1f, 32'h40ed3016} /* (11, 0, 7) {real, imag} */,
  {32'hc227078d, 32'hc1e16db4} /* (11, 0, 6) {real, imag} */,
  {32'h41a1f135, 32'hc272a7b7} /* (11, 0, 5) {real, imag} */,
  {32'h40ffd994, 32'h429fb157} /* (11, 0, 4) {real, imag} */,
  {32'h412970a8, 32'h40009420} /* (11, 0, 3) {real, imag} */,
  {32'h42254019, 32'h417256ac} /* (11, 0, 2) {real, imag} */,
  {32'hc0ca1a00, 32'hc2868a2a} /* (11, 0, 1) {real, imag} */,
  {32'h43a442d4, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'hc21aa9de, 32'h41616fc4} /* (10, 15, 15) {real, imag} */,
  {32'hc21dcc5b, 32'hc1d34251} /* (10, 15, 14) {real, imag} */,
  {32'h42b003dc, 32'h41ebd09a} /* (10, 15, 13) {real, imag} */,
  {32'h41368ed4, 32'h413de04e} /* (10, 15, 12) {real, imag} */,
  {32'h41c1adda, 32'h41d609f6} /* (10, 15, 11) {real, imag} */,
  {32'h4201a4db, 32'h4216b578} /* (10, 15, 10) {real, imag} */,
  {32'hc13616ba, 32'hc0c7fa4c} /* (10, 15, 9) {real, imag} */,
  {32'h4013cf7e, 32'h40d04ad1} /* (10, 15, 8) {real, imag} */,
  {32'hc2042963, 32'hc091c1b8} /* (10, 15, 7) {real, imag} */,
  {32'hc0963523, 32'h41cf6ae4} /* (10, 15, 6) {real, imag} */,
  {32'h41ab8eef, 32'hc145e945} /* (10, 15, 5) {real, imag} */,
  {32'hc15fc80c, 32'h41b112cc} /* (10, 15, 4) {real, imag} */,
  {32'h423c7210, 32'hc202eca7} /* (10, 15, 3) {real, imag} */,
  {32'hc1d13b00, 32'hc1c5d15a} /* (10, 15, 2) {real, imag} */,
  {32'h40848258, 32'h4020acf0} /* (10, 15, 1) {real, imag} */,
  {32'hc26afe61, 32'hc30a1600} /* (10, 15, 0) {real, imag} */,
  {32'hc15b148c, 32'hc2f9bb7c} /* (10, 14, 15) {real, imag} */,
  {32'hc29e55f4, 32'h42869f7c} /* (10, 14, 14) {real, imag} */,
  {32'hc1dbe5b5, 32'hc1dc524d} /* (10, 14, 13) {real, imag} */,
  {32'hc01f0cb8, 32'hc142dbfe} /* (10, 14, 12) {real, imag} */,
  {32'hc01cf218, 32'h4220f315} /* (10, 14, 11) {real, imag} */,
  {32'hc199fa4e, 32'hc1a77fef} /* (10, 14, 10) {real, imag} */,
  {32'h4107b165, 32'h40fe5c9e} /* (10, 14, 9) {real, imag} */,
  {32'hc10715b6, 32'h413f2115} /* (10, 14, 8) {real, imag} */,
  {32'hc01a6702, 32'h3fb1d258} /* (10, 14, 7) {real, imag} */,
  {32'hc1c793d8, 32'h421ddd2c} /* (10, 14, 6) {real, imag} */,
  {32'h40ebc958, 32'hc19c0ad7} /* (10, 14, 5) {real, imag} */,
  {32'h403a64c4, 32'h42260ece} /* (10, 14, 4) {real, imag} */,
  {32'hc13419a0, 32'hc13c423c} /* (10, 14, 3) {real, imag} */,
  {32'h428a0c78, 32'h41e9133f} /* (10, 14, 2) {real, imag} */,
  {32'h42cce91e, 32'h425a699f} /* (10, 14, 1) {real, imag} */,
  {32'hc0df8168, 32'h41c6e46f} /* (10, 14, 0) {real, imag} */,
  {32'hc15b8bf4, 32'hc113f31c} /* (10, 13, 15) {real, imag} */,
  {32'hc1b23504, 32'hc0acd458} /* (10, 13, 14) {real, imag} */,
  {32'h421b44e8, 32'hc1a5cb64} /* (10, 13, 13) {real, imag} */,
  {32'h422d2814, 32'h42087a99} /* (10, 13, 12) {real, imag} */,
  {32'h4080181a, 32'hc0c9a35c} /* (10, 13, 11) {real, imag} */,
  {32'hc1eba97f, 32'h40fa3af2} /* (10, 13, 10) {real, imag} */,
  {32'h41c8efd2, 32'h3ef13e40} /* (10, 13, 9) {real, imag} */,
  {32'h4137a9fa, 32'hbde01110} /* (10, 13, 8) {real, imag} */,
  {32'h4122e7d6, 32'hbff16298} /* (10, 13, 7) {real, imag} */,
  {32'hc0bdd894, 32'hc19c2f1f} /* (10, 13, 6) {real, imag} */,
  {32'h3fb1ad58, 32'h422d6e7c} /* (10, 13, 5) {real, imag} */,
  {32'h3f940640, 32'h400d4e70} /* (10, 13, 4) {real, imag} */,
  {32'h40db5cd6, 32'h41a6dffc} /* (10, 13, 3) {real, imag} */,
  {32'hc16c2cc3, 32'hc0d089ef} /* (10, 13, 2) {real, imag} */,
  {32'hc12735ac, 32'hc29c2018} /* (10, 13, 1) {real, imag} */,
  {32'h41b994fc, 32'h40d1464c} /* (10, 13, 0) {real, imag} */,
  {32'h41e681d6, 32'h416fc218} /* (10, 12, 15) {real, imag} */,
  {32'h420e17b3, 32'h422be2a4} /* (10, 12, 14) {real, imag} */,
  {32'hc1910cd8, 32'h41894cfe} /* (10, 12, 13) {real, imag} */,
  {32'hbf8c14c6, 32'h4051c310} /* (10, 12, 12) {real, imag} */,
  {32'hc119ab68, 32'h4029f36f} /* (10, 12, 11) {real, imag} */,
  {32'hc14f7f06, 32'h419b9273} /* (10, 12, 10) {real, imag} */,
  {32'hc178bb33, 32'hc1cf46db} /* (10, 12, 9) {real, imag} */,
  {32'hc1f1c3c3, 32'hc11b4578} /* (10, 12, 8) {real, imag} */,
  {32'h40703cb4, 32'h415c732c} /* (10, 12, 7) {real, imag} */,
  {32'h4209cdda, 32'hc1c15390} /* (10, 12, 6) {real, imag} */,
  {32'h40d9d4b4, 32'hc0d1cef6} /* (10, 12, 5) {real, imag} */,
  {32'hc1d36c30, 32'h41120eef} /* (10, 12, 4) {real, imag} */,
  {32'h40a7164c, 32'h41b79f6d} /* (10, 12, 3) {real, imag} */,
  {32'h41e3b156, 32'hc1a1feac} /* (10, 12, 2) {real, imag} */,
  {32'hc0af66bb, 32'h41c6cddc} /* (10, 12, 1) {real, imag} */,
  {32'hc13a519e, 32'h4149bf3c} /* (10, 12, 0) {real, imag} */,
  {32'h422acdc4, 32'h42080ede} /* (10, 11, 15) {real, imag} */,
  {32'h413b4254, 32'hc08be040} /* (10, 11, 14) {real, imag} */,
  {32'h40ae093c, 32'h40000acc} /* (10, 11, 13) {real, imag} */,
  {32'hbfd17e60, 32'hc1caba20} /* (10, 11, 12) {real, imag} */,
  {32'h3f0538f0, 32'hc150388a} /* (10, 11, 11) {real, imag} */,
  {32'hc0b49a12, 32'h418a6780} /* (10, 11, 10) {real, imag} */,
  {32'hc1b1b08b, 32'h415f3860} /* (10, 11, 9) {real, imag} */,
  {32'h41bd2d90, 32'hbf7ccca8} /* (10, 11, 8) {real, imag} */,
  {32'hc1789c8b, 32'hc1bbedf6} /* (10, 11, 7) {real, imag} */,
  {32'h419837ed, 32'hc0f82ab4} /* (10, 11, 6) {real, imag} */,
  {32'h421aeb40, 32'hc13901fa} /* (10, 11, 5) {real, imag} */,
  {32'hc1d49793, 32'h40fec690} /* (10, 11, 4) {real, imag} */,
  {32'hc193ab52, 32'hc184478b} /* (10, 11, 3) {real, imag} */,
  {32'hc16a2e1f, 32'hc243d25f} /* (10, 11, 2) {real, imag} */,
  {32'h4228c309, 32'h41a62177} /* (10, 11, 1) {real, imag} */,
  {32'h41e5bf71, 32'h4216aec2} /* (10, 11, 0) {real, imag} */,
  {32'hc18af2f1, 32'hc1b9590c} /* (10, 10, 15) {real, imag} */,
  {32'hc20bc61c, 32'hc07ed398} /* (10, 10, 14) {real, imag} */,
  {32'h41700354, 32'hc0ab23cb} /* (10, 10, 13) {real, imag} */,
  {32'hc06e9d88, 32'h41a2494f} /* (10, 10, 12) {real, imag} */,
  {32'h3fad6ff0, 32'h420a8fc1} /* (10, 10, 11) {real, imag} */,
  {32'hc1a59ff2, 32'h41174db0} /* (10, 10, 10) {real, imag} */,
  {32'hc0a05502, 32'hc061cfb2} /* (10, 10, 9) {real, imag} */,
  {32'hc144bd79, 32'h4182477e} /* (10, 10, 8) {real, imag} */,
  {32'hc11af240, 32'hc1ca601e} /* (10, 10, 7) {real, imag} */,
  {32'h414e94d8, 32'hc0bbbb82} /* (10, 10, 6) {real, imag} */,
  {32'h3ed1b750, 32'h41dcb272} /* (10, 10, 5) {real, imag} */,
  {32'h4213866a, 32'h40d960c2} /* (10, 10, 4) {real, imag} */,
  {32'hc182894c, 32'h41b12876} /* (10, 10, 3) {real, imag} */,
  {32'hc0e64405, 32'h40d894f2} /* (10, 10, 2) {real, imag} */,
  {32'hc227d602, 32'h4201f27c} /* (10, 10, 1) {real, imag} */,
  {32'h40af6c3c, 32'h408482ac} /* (10, 10, 0) {real, imag} */,
  {32'hc0cee951, 32'hc0ee9fc7} /* (10, 9, 15) {real, imag} */,
  {32'h418c2dec, 32'hbece6800} /* (10, 9, 14) {real, imag} */,
  {32'hc10aeaee, 32'hc027dda2} /* (10, 9, 13) {real, imag} */,
  {32'hc0f0017f, 32'hc12005a0} /* (10, 9, 12) {real, imag} */,
  {32'hc139f0da, 32'hc05e3fdd} /* (10, 9, 11) {real, imag} */,
  {32'h41b08b10, 32'hc1bef6a4} /* (10, 9, 10) {real, imag} */,
  {32'h41ea80cf, 32'hc0494ba8} /* (10, 9, 9) {real, imag} */,
  {32'hc155e262, 32'hc0bb2cfa} /* (10, 9, 8) {real, imag} */,
  {32'h41840594, 32'hc1a82b72} /* (10, 9, 7) {real, imag} */,
  {32'h41209493, 32'h3fdbd3f8} /* (10, 9, 6) {real, imag} */,
  {32'h4187c8a8, 32'hc1e1cac2} /* (10, 9, 5) {real, imag} */,
  {32'h40da3e19, 32'h4197e23e} /* (10, 9, 4) {real, imag} */,
  {32'hc10f3412, 32'h40ee75e4} /* (10, 9, 3) {real, imag} */,
  {32'hc1e1e3e4, 32'h41a345eb} /* (10, 9, 2) {real, imag} */,
  {32'h41cff254, 32'h410d9d8c} /* (10, 9, 1) {real, imag} */,
  {32'hc1597065, 32'hc111105c} /* (10, 9, 0) {real, imag} */,
  {32'hc004e562, 32'hc09c0a50} /* (10, 8, 15) {real, imag} */,
  {32'h3fe37e0c, 32'hc1968525} /* (10, 8, 14) {real, imag} */,
  {32'h3f0307f0, 32'h40e93ae1} /* (10, 8, 13) {real, imag} */,
  {32'h4188c3f2, 32'h406e62b0} /* (10, 8, 12) {real, imag} */,
  {32'hc10185f8, 32'hc1791d98} /* (10, 8, 11) {real, imag} */,
  {32'hc144a9bb, 32'hc15c4872} /* (10, 8, 10) {real, imag} */,
  {32'hc13877fa, 32'hc0b48e16} /* (10, 8, 9) {real, imag} */,
  {32'hc016f250, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'hc13877fa, 32'h40b48e16} /* (10, 8, 7) {real, imag} */,
  {32'hc144a9bb, 32'h415c4872} /* (10, 8, 6) {real, imag} */,
  {32'hc10185f8, 32'h41791d98} /* (10, 8, 5) {real, imag} */,
  {32'h4188c3f2, 32'hc06e62b0} /* (10, 8, 4) {real, imag} */,
  {32'h3f0307f0, 32'hc0e93ae1} /* (10, 8, 3) {real, imag} */,
  {32'h3fe37e0c, 32'h41968525} /* (10, 8, 2) {real, imag} */,
  {32'hc004e562, 32'h409c0a50} /* (10, 8, 1) {real, imag} */,
  {32'hc0cf279c, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h41cff254, 32'hc10d9d8c} /* (10, 7, 15) {real, imag} */,
  {32'hc1e1e3e4, 32'hc1a345eb} /* (10, 7, 14) {real, imag} */,
  {32'hc10f3412, 32'hc0ee75e4} /* (10, 7, 13) {real, imag} */,
  {32'h40da3e19, 32'hc197e23e} /* (10, 7, 12) {real, imag} */,
  {32'h4187c8a8, 32'h41e1cac2} /* (10, 7, 11) {real, imag} */,
  {32'h41209493, 32'hbfdbd3f8} /* (10, 7, 10) {real, imag} */,
  {32'h41840594, 32'h41a82b72} /* (10, 7, 9) {real, imag} */,
  {32'hc155e262, 32'h40bb2cfa} /* (10, 7, 8) {real, imag} */,
  {32'h41ea80cf, 32'h40494ba8} /* (10, 7, 7) {real, imag} */,
  {32'h41b08b10, 32'h41bef6a4} /* (10, 7, 6) {real, imag} */,
  {32'hc139f0da, 32'h405e3fdd} /* (10, 7, 5) {real, imag} */,
  {32'hc0f0017f, 32'h412005a0} /* (10, 7, 4) {real, imag} */,
  {32'hc10aeaee, 32'h4027dda2} /* (10, 7, 3) {real, imag} */,
  {32'h418c2dec, 32'h3ece6800} /* (10, 7, 2) {real, imag} */,
  {32'hc0cee951, 32'h40ee9fc7} /* (10, 7, 1) {real, imag} */,
  {32'hc1597065, 32'h4111105c} /* (10, 7, 0) {real, imag} */,
  {32'hc227d602, 32'hc201f27c} /* (10, 6, 15) {real, imag} */,
  {32'hc0e64405, 32'hc0d894f2} /* (10, 6, 14) {real, imag} */,
  {32'hc182894c, 32'hc1b12876} /* (10, 6, 13) {real, imag} */,
  {32'h4213866a, 32'hc0d960c2} /* (10, 6, 12) {real, imag} */,
  {32'h3ed1b750, 32'hc1dcb272} /* (10, 6, 11) {real, imag} */,
  {32'h414e94d8, 32'h40bbbb82} /* (10, 6, 10) {real, imag} */,
  {32'hc11af240, 32'h41ca601e} /* (10, 6, 9) {real, imag} */,
  {32'hc144bd79, 32'hc182477e} /* (10, 6, 8) {real, imag} */,
  {32'hc0a05502, 32'h4061cfb2} /* (10, 6, 7) {real, imag} */,
  {32'hc1a59ff2, 32'hc1174db0} /* (10, 6, 6) {real, imag} */,
  {32'h3fad6ff0, 32'hc20a8fc1} /* (10, 6, 5) {real, imag} */,
  {32'hc06e9d88, 32'hc1a2494f} /* (10, 6, 4) {real, imag} */,
  {32'h41700354, 32'h40ab23cb} /* (10, 6, 3) {real, imag} */,
  {32'hc20bc61c, 32'h407ed398} /* (10, 6, 2) {real, imag} */,
  {32'hc18af2f1, 32'h41b9590c} /* (10, 6, 1) {real, imag} */,
  {32'h40af6c3c, 32'hc08482ac} /* (10, 6, 0) {real, imag} */,
  {32'h4228c309, 32'hc1a62177} /* (10, 5, 15) {real, imag} */,
  {32'hc16a2e1f, 32'h4243d25f} /* (10, 5, 14) {real, imag} */,
  {32'hc193ab52, 32'h4184478b} /* (10, 5, 13) {real, imag} */,
  {32'hc1d49793, 32'hc0fec690} /* (10, 5, 12) {real, imag} */,
  {32'h421aeb40, 32'h413901fa} /* (10, 5, 11) {real, imag} */,
  {32'h419837ed, 32'h40f82ab4} /* (10, 5, 10) {real, imag} */,
  {32'hc1789c8b, 32'h41bbedf6} /* (10, 5, 9) {real, imag} */,
  {32'h41bd2d90, 32'h3f7ccca8} /* (10, 5, 8) {real, imag} */,
  {32'hc1b1b08b, 32'hc15f3860} /* (10, 5, 7) {real, imag} */,
  {32'hc0b49a12, 32'hc18a6780} /* (10, 5, 6) {real, imag} */,
  {32'h3f0538f0, 32'h4150388a} /* (10, 5, 5) {real, imag} */,
  {32'hbfd17e60, 32'h41caba20} /* (10, 5, 4) {real, imag} */,
  {32'h40ae093c, 32'hc0000acc} /* (10, 5, 3) {real, imag} */,
  {32'h413b4254, 32'h408be040} /* (10, 5, 2) {real, imag} */,
  {32'h422acdc4, 32'hc2080ede} /* (10, 5, 1) {real, imag} */,
  {32'h41e5bf71, 32'hc216aec2} /* (10, 5, 0) {real, imag} */,
  {32'hc0af66bb, 32'hc1c6cddc} /* (10, 4, 15) {real, imag} */,
  {32'h41e3b156, 32'h41a1feac} /* (10, 4, 14) {real, imag} */,
  {32'h40a7164c, 32'hc1b79f6d} /* (10, 4, 13) {real, imag} */,
  {32'hc1d36c30, 32'hc1120eef} /* (10, 4, 12) {real, imag} */,
  {32'h40d9d4b4, 32'h40d1cef6} /* (10, 4, 11) {real, imag} */,
  {32'h4209cdda, 32'h41c15390} /* (10, 4, 10) {real, imag} */,
  {32'h40703cb4, 32'hc15c732c} /* (10, 4, 9) {real, imag} */,
  {32'hc1f1c3c3, 32'h411b4578} /* (10, 4, 8) {real, imag} */,
  {32'hc178bb33, 32'h41cf46db} /* (10, 4, 7) {real, imag} */,
  {32'hc14f7f06, 32'hc19b9273} /* (10, 4, 6) {real, imag} */,
  {32'hc119ab68, 32'hc029f36f} /* (10, 4, 5) {real, imag} */,
  {32'hbf8c14c6, 32'hc051c310} /* (10, 4, 4) {real, imag} */,
  {32'hc1910cd8, 32'hc1894cfe} /* (10, 4, 3) {real, imag} */,
  {32'h420e17b3, 32'hc22be2a4} /* (10, 4, 2) {real, imag} */,
  {32'h41e681d6, 32'hc16fc218} /* (10, 4, 1) {real, imag} */,
  {32'hc13a519e, 32'hc149bf3c} /* (10, 4, 0) {real, imag} */,
  {32'hc12735ac, 32'h429c2018} /* (10, 3, 15) {real, imag} */,
  {32'hc16c2cc3, 32'h40d089ef} /* (10, 3, 14) {real, imag} */,
  {32'h40db5cd6, 32'hc1a6dffc} /* (10, 3, 13) {real, imag} */,
  {32'h3f940640, 32'hc00d4e70} /* (10, 3, 12) {real, imag} */,
  {32'h3fb1ad58, 32'hc22d6e7c} /* (10, 3, 11) {real, imag} */,
  {32'hc0bdd894, 32'h419c2f1f} /* (10, 3, 10) {real, imag} */,
  {32'h4122e7d6, 32'h3ff16298} /* (10, 3, 9) {real, imag} */,
  {32'h4137a9fa, 32'h3de01110} /* (10, 3, 8) {real, imag} */,
  {32'h41c8efd2, 32'hbef13e40} /* (10, 3, 7) {real, imag} */,
  {32'hc1eba97f, 32'hc0fa3af2} /* (10, 3, 6) {real, imag} */,
  {32'h4080181a, 32'h40c9a35c} /* (10, 3, 5) {real, imag} */,
  {32'h422d2814, 32'hc2087a99} /* (10, 3, 4) {real, imag} */,
  {32'h421b44e8, 32'h41a5cb64} /* (10, 3, 3) {real, imag} */,
  {32'hc1b23504, 32'h40acd458} /* (10, 3, 2) {real, imag} */,
  {32'hc15b8bf4, 32'h4113f31c} /* (10, 3, 1) {real, imag} */,
  {32'h41b994fc, 32'hc0d1464c} /* (10, 3, 0) {real, imag} */,
  {32'h42cce91e, 32'hc25a699f} /* (10, 2, 15) {real, imag} */,
  {32'h428a0c78, 32'hc1e9133f} /* (10, 2, 14) {real, imag} */,
  {32'hc13419a0, 32'h413c423c} /* (10, 2, 13) {real, imag} */,
  {32'h403a64c4, 32'hc2260ece} /* (10, 2, 12) {real, imag} */,
  {32'h40ebc958, 32'h419c0ad7} /* (10, 2, 11) {real, imag} */,
  {32'hc1c793d8, 32'hc21ddd2c} /* (10, 2, 10) {real, imag} */,
  {32'hc01a6702, 32'hbfb1d258} /* (10, 2, 9) {real, imag} */,
  {32'hc10715b6, 32'hc13f2115} /* (10, 2, 8) {real, imag} */,
  {32'h4107b165, 32'hc0fe5c9e} /* (10, 2, 7) {real, imag} */,
  {32'hc199fa4e, 32'h41a77fef} /* (10, 2, 6) {real, imag} */,
  {32'hc01cf218, 32'hc220f315} /* (10, 2, 5) {real, imag} */,
  {32'hc01f0cb8, 32'h4142dbfe} /* (10, 2, 4) {real, imag} */,
  {32'hc1dbe5b5, 32'h41dc524d} /* (10, 2, 3) {real, imag} */,
  {32'hc29e55f4, 32'hc2869f7c} /* (10, 2, 2) {real, imag} */,
  {32'hc15b148c, 32'h42f9bb7c} /* (10, 2, 1) {real, imag} */,
  {32'hc0df8168, 32'hc1c6e46f} /* (10, 2, 0) {real, imag} */,
  {32'h40848258, 32'hc020acf0} /* (10, 1, 15) {real, imag} */,
  {32'hc1d13b00, 32'h41c5d15a} /* (10, 1, 14) {real, imag} */,
  {32'h423c7210, 32'h4202eca7} /* (10, 1, 13) {real, imag} */,
  {32'hc15fc80c, 32'hc1b112cc} /* (10, 1, 12) {real, imag} */,
  {32'h41ab8eef, 32'h4145e945} /* (10, 1, 11) {real, imag} */,
  {32'hc0963523, 32'hc1cf6ae4} /* (10, 1, 10) {real, imag} */,
  {32'hc2042963, 32'h4091c1b8} /* (10, 1, 9) {real, imag} */,
  {32'h4013cf7e, 32'hc0d04ad1} /* (10, 1, 8) {real, imag} */,
  {32'hc13616ba, 32'h40c7fa4c} /* (10, 1, 7) {real, imag} */,
  {32'h4201a4db, 32'hc216b578} /* (10, 1, 6) {real, imag} */,
  {32'h41c1adda, 32'hc1d609f6} /* (10, 1, 5) {real, imag} */,
  {32'h41368ed4, 32'hc13de04e} /* (10, 1, 4) {real, imag} */,
  {32'h42b003dc, 32'hc1ebd09a} /* (10, 1, 3) {real, imag} */,
  {32'hc21dcc5b, 32'h41d34251} /* (10, 1, 2) {real, imag} */,
  {32'hc21aa9de, 32'hc1616fc4} /* (10, 1, 1) {real, imag} */,
  {32'hc26afe61, 32'h430a1600} /* (10, 1, 0) {real, imag} */,
  {32'hc178ea98, 32'h42a25b98} /* (10, 0, 15) {real, imag} */,
  {32'h41b14680, 32'hc2aaf258} /* (10, 0, 14) {real, imag} */,
  {32'h40edab5d, 32'hc1483ef1} /* (10, 0, 13) {real, imag} */,
  {32'h41774d6d, 32'hc17e3b66} /* (10, 0, 12) {real, imag} */,
  {32'h3f856f50, 32'h422f9ec4} /* (10, 0, 11) {real, imag} */,
  {32'hc00b3875, 32'h413302c2} /* (10, 0, 10) {real, imag} */,
  {32'h41a8e612, 32'hc17cc0d1} /* (10, 0, 9) {real, imag} */,
  {32'hc0461e1e, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'h41a8e612, 32'h417cc0d1} /* (10, 0, 7) {real, imag} */,
  {32'hc00b3875, 32'hc13302c2} /* (10, 0, 6) {real, imag} */,
  {32'h3f856f50, 32'hc22f9ec4} /* (10, 0, 5) {real, imag} */,
  {32'h41774d6d, 32'h417e3b66} /* (10, 0, 4) {real, imag} */,
  {32'h40edab5d, 32'h41483ef1} /* (10, 0, 3) {real, imag} */,
  {32'h41b14680, 32'h42aaf258} /* (10, 0, 2) {real, imag} */,
  {32'hc178ea98, 32'hc2a25b98} /* (10, 0, 1) {real, imag} */,
  {32'h43b998eb, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'hc2369551, 32'hc0e8f370} /* (9, 15, 15) {real, imag} */,
  {32'h411285f8, 32'hc19b7e90} /* (9, 15, 14) {real, imag} */,
  {32'h40f9e0c6, 32'h41317aad} /* (9, 15, 13) {real, imag} */,
  {32'h4229c686, 32'hc0bc97fe} /* (9, 15, 12) {real, imag} */,
  {32'h41820989, 32'h41f5cc7f} /* (9, 15, 11) {real, imag} */,
  {32'hc1752223, 32'hc1b4e9df} /* (9, 15, 10) {real, imag} */,
  {32'hc0f29e54, 32'hbf34b138} /* (9, 15, 9) {real, imag} */,
  {32'h4171f126, 32'h3e780840} /* (9, 15, 8) {real, imag} */,
  {32'hc18b9149, 32'hc18110ea} /* (9, 15, 7) {real, imag} */,
  {32'h413b6dc0, 32'h4113252a} /* (9, 15, 6) {real, imag} */,
  {32'hc19e9a20, 32'hc14083ab} /* (9, 15, 5) {real, imag} */,
  {32'hc17b72f2, 32'h419e374f} /* (9, 15, 4) {real, imag} */,
  {32'h4220bfaf, 32'h414c5c33} /* (9, 15, 3) {real, imag} */,
  {32'hc25c1d96, 32'hc274b1a6} /* (9, 15, 2) {real, imag} */,
  {32'hc1d9c586, 32'h420c9720} /* (9, 15, 1) {real, imag} */,
  {32'hc27ba610, 32'hc2f2de73} /* (9, 15, 0) {real, imag} */,
  {32'hc2638e86, 32'hc1c00c18} /* (9, 14, 15) {real, imag} */,
  {32'hc28addee, 32'h4296581d} /* (9, 14, 14) {real, imag} */,
  {32'hc090f6c4, 32'h3f1935d8} /* (9, 14, 13) {real, imag} */,
  {32'h421fce7e, 32'hc1fce845} /* (9, 14, 12) {real, imag} */,
  {32'hc2416022, 32'hc08bc242} /* (9, 14, 11) {real, imag} */,
  {32'hc1914fc0, 32'h406626d8} /* (9, 14, 10) {real, imag} */,
  {32'h418873c7, 32'hc00f1108} /* (9, 14, 9) {real, imag} */,
  {32'hc0b49dbe, 32'hc053c701} /* (9, 14, 8) {real, imag} */,
  {32'hc1a912d2, 32'hc1a0ccc0} /* (9, 14, 7) {real, imag} */,
  {32'h42090cf0, 32'h40827a50} /* (9, 14, 6) {real, imag} */,
  {32'h42596f3c, 32'hc1a914ae} /* (9, 14, 5) {real, imag} */,
  {32'hc2208411, 32'h4234dd3a} /* (9, 14, 4) {real, imag} */,
  {32'hc228442d, 32'hc255251d} /* (9, 14, 3) {real, imag} */,
  {32'h42a6e6c2, 32'h42584bd9} /* (9, 14, 2) {real, imag} */,
  {32'h42c26353, 32'h41fedf96} /* (9, 14, 1) {real, imag} */,
  {32'hc034d3bc, 32'hc0b7f8e0} /* (9, 14, 0) {real, imag} */,
  {32'h4148637f, 32'hc182d85a} /* (9, 13, 15) {real, imag} */,
  {32'hc1ecf0df, 32'h41cf15ae} /* (9, 13, 14) {real, imag} */,
  {32'h417d34ee, 32'hc1ccfd60} /* (9, 13, 13) {real, imag} */,
  {32'hc161ff1d, 32'h3e372400} /* (9, 13, 12) {real, imag} */,
  {32'hc1159250, 32'hc0632600} /* (9, 13, 11) {real, imag} */,
  {32'hc1b02644, 32'hc13d0e9f} /* (9, 13, 10) {real, imag} */,
  {32'hc1d8971e, 32'hc2324ea4} /* (9, 13, 9) {real, imag} */,
  {32'h41043719, 32'h4082b0ac} /* (9, 13, 8) {real, imag} */,
  {32'hc11ae98a, 32'hc0339a02} /* (9, 13, 7) {real, imag} */,
  {32'hc1bfc40a, 32'hc0ad3aef} /* (9, 13, 6) {real, imag} */,
  {32'h421b24ea, 32'h41810e5e} /* (9, 13, 5) {real, imag} */,
  {32'hc10e4ac8, 32'h420bcc4a} /* (9, 13, 4) {real, imag} */,
  {32'hc15d0f70, 32'h424475b8} /* (9, 13, 3) {real, imag} */,
  {32'hc0b3e4bb, 32'h3f73a820} /* (9, 13, 2) {real, imag} */,
  {32'hc1bc1492, 32'hc204f95c} /* (9, 13, 1) {real, imag} */,
  {32'h422722e0, 32'hc0c6dbc4} /* (9, 13, 0) {real, imag} */,
  {32'hc15fe5ba, 32'hc19f1a52} /* (9, 12, 15) {real, imag} */,
  {32'h3f46e508, 32'h40786fde} /* (9, 12, 14) {real, imag} */,
  {32'h41059202, 32'h413a0d1e} /* (9, 12, 13) {real, imag} */,
  {32'h41a2776e, 32'hc1ced134} /* (9, 12, 12) {real, imag} */,
  {32'hc1ba835a, 32'h410747ea} /* (9, 12, 11) {real, imag} */,
  {32'h4103a372, 32'h41317767} /* (9, 12, 10) {real, imag} */,
  {32'h40db6694, 32'hc0a53044} /* (9, 12, 9) {real, imag} */,
  {32'h412edfb4, 32'h41374761} /* (9, 12, 8) {real, imag} */,
  {32'hc13e8ef8, 32'hbf5c4960} /* (9, 12, 7) {real, imag} */,
  {32'h41e87ede, 32'h41ea0c85} /* (9, 12, 6) {real, imag} */,
  {32'h41e7e9f8, 32'h411a40a4} /* (9, 12, 5) {real, imag} */,
  {32'h3f9dfe28, 32'h423f1fd4} /* (9, 12, 4) {real, imag} */,
  {32'hc0308872, 32'h4093b0be} /* (9, 12, 3) {real, imag} */,
  {32'hc1b8ae33, 32'hc01b1ab2} /* (9, 12, 2) {real, imag} */,
  {32'hc022bc54, 32'hc2071116} /* (9, 12, 1) {real, imag} */,
  {32'hc176fc38, 32'h4176b746} /* (9, 12, 0) {real, imag} */,
  {32'h41478dae, 32'hc130a024} /* (9, 11, 15) {real, imag} */,
  {32'h423a66c2, 32'hc1efa8b3} /* (9, 11, 14) {real, imag} */,
  {32'hc212feee, 32'hc17c356e} /* (9, 11, 13) {real, imag} */,
  {32'h4187e490, 32'h415a4e7a} /* (9, 11, 12) {real, imag} */,
  {32'h41708fa1, 32'h41726023} /* (9, 11, 11) {real, imag} */,
  {32'hc109042c, 32'h419ebf15} /* (9, 11, 10) {real, imag} */,
  {32'h42041db1, 32'hc1bc7616} /* (9, 11, 9) {real, imag} */,
  {32'hc17af6ad, 32'h410ee299} /* (9, 11, 8) {real, imag} */,
  {32'h4083823e, 32'h41edf3c2} /* (9, 11, 7) {real, imag} */,
  {32'hc0cd0f6b, 32'hc1ac135e} /* (9, 11, 6) {real, imag} */,
  {32'hc1a79a89, 32'h41d5a0af} /* (9, 11, 5) {real, imag} */,
  {32'h4221706a, 32'hc002f1fc} /* (9, 11, 4) {real, imag} */,
  {32'hc1e0bf63, 32'hc2122572} /* (9, 11, 3) {real, imag} */,
  {32'hc1591d79, 32'hc23c8d10} /* (9, 11, 2) {real, imag} */,
  {32'hc1150432, 32'h40a9af9d} /* (9, 11, 1) {real, imag} */,
  {32'hc21dfd49, 32'h413042ba} /* (9, 11, 0) {real, imag} */,
  {32'h40deae24, 32'hc08570c4} /* (9, 10, 15) {real, imag} */,
  {32'h4208c9fe, 32'hc12b97b5} /* (9, 10, 14) {real, imag} */,
  {32'h4217479a, 32'h414a3ba7} /* (9, 10, 13) {real, imag} */,
  {32'hc26cbed2, 32'h4255f01b} /* (9, 10, 12) {real, imag} */,
  {32'hc156eaaa, 32'hc0d98992} /* (9, 10, 11) {real, imag} */,
  {32'hc20f0de8, 32'hc1ab5341} /* (9, 10, 10) {real, imag} */,
  {32'h4159441e, 32'h4182d972} /* (9, 10, 9) {real, imag} */,
  {32'hc134adb2, 32'hc2326c74} /* (9, 10, 8) {real, imag} */,
  {32'hc0347b61, 32'hc11ed01c} /* (9, 10, 7) {real, imag} */,
  {32'h40765628, 32'h41a010ca} /* (9, 10, 6) {real, imag} */,
  {32'h402f0e8a, 32'h415d9761} /* (9, 10, 5) {real, imag} */,
  {32'hc1a70a0e, 32'hc185c185} /* (9, 10, 4) {real, imag} */,
  {32'h409b76a0, 32'h41a2d28a} /* (9, 10, 3) {real, imag} */,
  {32'h4163865e, 32'hc14a572f} /* (9, 10, 2) {real, imag} */,
  {32'hc08f9152, 32'h3fa2fc38} /* (9, 10, 1) {real, imag} */,
  {32'hc09c3670, 32'h41786972} /* (9, 10, 0) {real, imag} */,
  {32'h41b882a7, 32'hc1c0f74a} /* (9, 9, 15) {real, imag} */,
  {32'hc104dcbb, 32'h40ad8374} /* (9, 9, 14) {real, imag} */,
  {32'h4186f0a8, 32'hc1199416} /* (9, 9, 13) {real, imag} */,
  {32'h3f1bd050, 32'h41d06174} /* (9, 9, 12) {real, imag} */,
  {32'h4109b540, 32'hc1e3beca} /* (9, 9, 11) {real, imag} */,
  {32'hc0e6ad30, 32'hc21c17c0} /* (9, 9, 10) {real, imag} */,
  {32'hc1b82299, 32'h421c2fcf} /* (9, 9, 9) {real, imag} */,
  {32'h40ef50aa, 32'hc13bb24a} /* (9, 9, 8) {real, imag} */,
  {32'h3f4663dc, 32'h40e6f39a} /* (9, 9, 7) {real, imag} */,
  {32'h41e6b2c1, 32'h410c83b8} /* (9, 9, 6) {real, imag} */,
  {32'hc1d43e55, 32'hbfdd58d0} /* (9, 9, 5) {real, imag} */,
  {32'hc1900ffa, 32'h41751462} /* (9, 9, 4) {real, imag} */,
  {32'h3f903308, 32'hc09c59c8} /* (9, 9, 3) {real, imag} */,
  {32'h40b0385c, 32'h41c8dad2} /* (9, 9, 2) {real, imag} */,
  {32'hc1ca7578, 32'hc21fc830} /* (9, 9, 1) {real, imag} */,
  {32'h41359ff8, 32'h40fe8104} /* (9, 9, 0) {real, imag} */,
  {32'hc030ff56, 32'hc1a42da5} /* (9, 8, 15) {real, imag} */,
  {32'hbfe97828, 32'hc10c59a2} /* (9, 8, 14) {real, imag} */,
  {32'h419019ef, 32'hbf04fac0} /* (9, 8, 13) {real, imag} */,
  {32'hc0bb9f7e, 32'hc0931b8a} /* (9, 8, 12) {real, imag} */,
  {32'h4111613e, 32'hc07b923e} /* (9, 8, 11) {real, imag} */,
  {32'hc1ca06d2, 32'hc0d2901e} /* (9, 8, 10) {real, imag} */,
  {32'hc15bd916, 32'h414aa452} /* (9, 8, 9) {real, imag} */,
  {32'hc0a8e092, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'hc15bd916, 32'hc14aa452} /* (9, 8, 7) {real, imag} */,
  {32'hc1ca06d2, 32'h40d2901e} /* (9, 8, 6) {real, imag} */,
  {32'h4111613e, 32'h407b923e} /* (9, 8, 5) {real, imag} */,
  {32'hc0bb9f7e, 32'h40931b8a} /* (9, 8, 4) {real, imag} */,
  {32'h419019ef, 32'h3f04fac0} /* (9, 8, 3) {real, imag} */,
  {32'hbfe97828, 32'h410c59a2} /* (9, 8, 2) {real, imag} */,
  {32'hc030ff56, 32'h41a42da5} /* (9, 8, 1) {real, imag} */,
  {32'hc1805e18, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'hc1ca7578, 32'h421fc830} /* (9, 7, 15) {real, imag} */,
  {32'h40b0385c, 32'hc1c8dad2} /* (9, 7, 14) {real, imag} */,
  {32'h3f903308, 32'h409c59c8} /* (9, 7, 13) {real, imag} */,
  {32'hc1900ffa, 32'hc1751462} /* (9, 7, 12) {real, imag} */,
  {32'hc1d43e55, 32'h3fdd58d0} /* (9, 7, 11) {real, imag} */,
  {32'h41e6b2c1, 32'hc10c83b8} /* (9, 7, 10) {real, imag} */,
  {32'h3f4663dc, 32'hc0e6f39a} /* (9, 7, 9) {real, imag} */,
  {32'h40ef50aa, 32'h413bb24a} /* (9, 7, 8) {real, imag} */,
  {32'hc1b82299, 32'hc21c2fcf} /* (9, 7, 7) {real, imag} */,
  {32'hc0e6ad30, 32'h421c17c0} /* (9, 7, 6) {real, imag} */,
  {32'h4109b540, 32'h41e3beca} /* (9, 7, 5) {real, imag} */,
  {32'h3f1bd050, 32'hc1d06174} /* (9, 7, 4) {real, imag} */,
  {32'h4186f0a8, 32'h41199416} /* (9, 7, 3) {real, imag} */,
  {32'hc104dcbb, 32'hc0ad8374} /* (9, 7, 2) {real, imag} */,
  {32'h41b882a7, 32'h41c0f74a} /* (9, 7, 1) {real, imag} */,
  {32'h41359ff8, 32'hc0fe8104} /* (9, 7, 0) {real, imag} */,
  {32'hc08f9152, 32'hbfa2fc38} /* (9, 6, 15) {real, imag} */,
  {32'h4163865e, 32'h414a572f} /* (9, 6, 14) {real, imag} */,
  {32'h409b76a0, 32'hc1a2d28a} /* (9, 6, 13) {real, imag} */,
  {32'hc1a70a0e, 32'h4185c185} /* (9, 6, 12) {real, imag} */,
  {32'h402f0e8a, 32'hc15d9761} /* (9, 6, 11) {real, imag} */,
  {32'h40765628, 32'hc1a010ca} /* (9, 6, 10) {real, imag} */,
  {32'hc0347b61, 32'h411ed01c} /* (9, 6, 9) {real, imag} */,
  {32'hc134adb2, 32'h42326c74} /* (9, 6, 8) {real, imag} */,
  {32'h4159441e, 32'hc182d972} /* (9, 6, 7) {real, imag} */,
  {32'hc20f0de8, 32'h41ab5341} /* (9, 6, 6) {real, imag} */,
  {32'hc156eaaa, 32'h40d98992} /* (9, 6, 5) {real, imag} */,
  {32'hc26cbed2, 32'hc255f01b} /* (9, 6, 4) {real, imag} */,
  {32'h4217479a, 32'hc14a3ba7} /* (9, 6, 3) {real, imag} */,
  {32'h4208c9fe, 32'h412b97b5} /* (9, 6, 2) {real, imag} */,
  {32'h40deae24, 32'h408570c4} /* (9, 6, 1) {real, imag} */,
  {32'hc09c3670, 32'hc1786972} /* (9, 6, 0) {real, imag} */,
  {32'hc1150432, 32'hc0a9af9d} /* (9, 5, 15) {real, imag} */,
  {32'hc1591d79, 32'h423c8d10} /* (9, 5, 14) {real, imag} */,
  {32'hc1e0bf63, 32'h42122572} /* (9, 5, 13) {real, imag} */,
  {32'h4221706a, 32'h4002f1fc} /* (9, 5, 12) {real, imag} */,
  {32'hc1a79a89, 32'hc1d5a0af} /* (9, 5, 11) {real, imag} */,
  {32'hc0cd0f6b, 32'h41ac135e} /* (9, 5, 10) {real, imag} */,
  {32'h4083823e, 32'hc1edf3c2} /* (9, 5, 9) {real, imag} */,
  {32'hc17af6ad, 32'hc10ee299} /* (9, 5, 8) {real, imag} */,
  {32'h42041db1, 32'h41bc7616} /* (9, 5, 7) {real, imag} */,
  {32'hc109042c, 32'hc19ebf15} /* (9, 5, 6) {real, imag} */,
  {32'h41708fa1, 32'hc1726023} /* (9, 5, 5) {real, imag} */,
  {32'h4187e490, 32'hc15a4e7a} /* (9, 5, 4) {real, imag} */,
  {32'hc212feee, 32'h417c356e} /* (9, 5, 3) {real, imag} */,
  {32'h423a66c2, 32'h41efa8b3} /* (9, 5, 2) {real, imag} */,
  {32'h41478dae, 32'h4130a024} /* (9, 5, 1) {real, imag} */,
  {32'hc21dfd49, 32'hc13042ba} /* (9, 5, 0) {real, imag} */,
  {32'hc022bc54, 32'h42071116} /* (9, 4, 15) {real, imag} */,
  {32'hc1b8ae33, 32'h401b1ab2} /* (9, 4, 14) {real, imag} */,
  {32'hc0308872, 32'hc093b0be} /* (9, 4, 13) {real, imag} */,
  {32'h3f9dfe28, 32'hc23f1fd4} /* (9, 4, 12) {real, imag} */,
  {32'h41e7e9f8, 32'hc11a40a4} /* (9, 4, 11) {real, imag} */,
  {32'h41e87ede, 32'hc1ea0c85} /* (9, 4, 10) {real, imag} */,
  {32'hc13e8ef8, 32'h3f5c4960} /* (9, 4, 9) {real, imag} */,
  {32'h412edfb4, 32'hc1374761} /* (9, 4, 8) {real, imag} */,
  {32'h40db6694, 32'h40a53044} /* (9, 4, 7) {real, imag} */,
  {32'h4103a372, 32'hc1317767} /* (9, 4, 6) {real, imag} */,
  {32'hc1ba835a, 32'hc10747ea} /* (9, 4, 5) {real, imag} */,
  {32'h41a2776e, 32'h41ced134} /* (9, 4, 4) {real, imag} */,
  {32'h41059202, 32'hc13a0d1e} /* (9, 4, 3) {real, imag} */,
  {32'h3f46e508, 32'hc0786fde} /* (9, 4, 2) {real, imag} */,
  {32'hc15fe5ba, 32'h419f1a52} /* (9, 4, 1) {real, imag} */,
  {32'hc176fc38, 32'hc176b746} /* (9, 4, 0) {real, imag} */,
  {32'hc1bc1492, 32'h4204f95c} /* (9, 3, 15) {real, imag} */,
  {32'hc0b3e4bb, 32'hbf73a820} /* (9, 3, 14) {real, imag} */,
  {32'hc15d0f70, 32'hc24475b8} /* (9, 3, 13) {real, imag} */,
  {32'hc10e4ac8, 32'hc20bcc4a} /* (9, 3, 12) {real, imag} */,
  {32'h421b24ea, 32'hc1810e5e} /* (9, 3, 11) {real, imag} */,
  {32'hc1bfc40a, 32'h40ad3aef} /* (9, 3, 10) {real, imag} */,
  {32'hc11ae98a, 32'h40339a02} /* (9, 3, 9) {real, imag} */,
  {32'h41043719, 32'hc082b0ac} /* (9, 3, 8) {real, imag} */,
  {32'hc1d8971e, 32'h42324ea4} /* (9, 3, 7) {real, imag} */,
  {32'hc1b02644, 32'h413d0e9f} /* (9, 3, 6) {real, imag} */,
  {32'hc1159250, 32'h40632600} /* (9, 3, 5) {real, imag} */,
  {32'hc161ff1d, 32'hbe372400} /* (9, 3, 4) {real, imag} */,
  {32'h417d34ee, 32'h41ccfd60} /* (9, 3, 3) {real, imag} */,
  {32'hc1ecf0df, 32'hc1cf15ae} /* (9, 3, 2) {real, imag} */,
  {32'h4148637f, 32'h4182d85a} /* (9, 3, 1) {real, imag} */,
  {32'h422722e0, 32'h40c6dbc4} /* (9, 3, 0) {real, imag} */,
  {32'h42c26353, 32'hc1fedf96} /* (9, 2, 15) {real, imag} */,
  {32'h42a6e6c2, 32'hc2584bd9} /* (9, 2, 14) {real, imag} */,
  {32'hc228442d, 32'h4255251d} /* (9, 2, 13) {real, imag} */,
  {32'hc2208411, 32'hc234dd3a} /* (9, 2, 12) {real, imag} */,
  {32'h42596f3c, 32'h41a914ae} /* (9, 2, 11) {real, imag} */,
  {32'h42090cf0, 32'hc0827a50} /* (9, 2, 10) {real, imag} */,
  {32'hc1a912d2, 32'h41a0ccc0} /* (9, 2, 9) {real, imag} */,
  {32'hc0b49dbe, 32'h4053c701} /* (9, 2, 8) {real, imag} */,
  {32'h418873c7, 32'h400f1108} /* (9, 2, 7) {real, imag} */,
  {32'hc1914fc0, 32'hc06626d8} /* (9, 2, 6) {real, imag} */,
  {32'hc2416022, 32'h408bc242} /* (9, 2, 5) {real, imag} */,
  {32'h421fce7e, 32'h41fce845} /* (9, 2, 4) {real, imag} */,
  {32'hc090f6c4, 32'hbf1935d8} /* (9, 2, 3) {real, imag} */,
  {32'hc28addee, 32'hc296581d} /* (9, 2, 2) {real, imag} */,
  {32'hc2638e86, 32'h41c00c18} /* (9, 2, 1) {real, imag} */,
  {32'hc034d3bc, 32'h40b7f8e0} /* (9, 2, 0) {real, imag} */,
  {32'hc1d9c586, 32'hc20c9720} /* (9, 1, 15) {real, imag} */,
  {32'hc25c1d96, 32'h4274b1a6} /* (9, 1, 14) {real, imag} */,
  {32'h4220bfaf, 32'hc14c5c33} /* (9, 1, 13) {real, imag} */,
  {32'hc17b72f2, 32'hc19e374f} /* (9, 1, 12) {real, imag} */,
  {32'hc19e9a20, 32'h414083ab} /* (9, 1, 11) {real, imag} */,
  {32'h413b6dc0, 32'hc113252a} /* (9, 1, 10) {real, imag} */,
  {32'hc18b9149, 32'h418110ea} /* (9, 1, 9) {real, imag} */,
  {32'h4171f126, 32'hbe780840} /* (9, 1, 8) {real, imag} */,
  {32'hc0f29e54, 32'h3f34b138} /* (9, 1, 7) {real, imag} */,
  {32'hc1752223, 32'h41b4e9df} /* (9, 1, 6) {real, imag} */,
  {32'h41820989, 32'hc1f5cc7f} /* (9, 1, 5) {real, imag} */,
  {32'h4229c686, 32'h40bc97fe} /* (9, 1, 4) {real, imag} */,
  {32'h40f9e0c6, 32'hc1317aad} /* (9, 1, 3) {real, imag} */,
  {32'h411285f8, 32'h419b7e90} /* (9, 1, 2) {real, imag} */,
  {32'hc2369551, 32'h40e8f370} /* (9, 1, 1) {real, imag} */,
  {32'hc27ba610, 32'h42f2de73} /* (9, 1, 0) {real, imag} */,
  {32'hc100d040, 32'h42d0c5b4} /* (9, 0, 15) {real, imag} */,
  {32'hc01b7338, 32'hc2da62a5} /* (9, 0, 14) {real, imag} */,
  {32'h41e68cc8, 32'h41364aca} /* (9, 0, 13) {real, imag} */,
  {32'h411f3da0, 32'h4218a23e} /* (9, 0, 12) {real, imag} */,
  {32'hc18d28c4, 32'hbd189c00} /* (9, 0, 11) {real, imag} */,
  {32'hc1ed16d8, 32'h425ed050} /* (9, 0, 10) {real, imag} */,
  {32'h41cd78b0, 32'hc0d20eb7} /* (9, 0, 9) {real, imag} */,
  {32'hc159adfe, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'h41cd78b0, 32'h40d20eb7} /* (9, 0, 7) {real, imag} */,
  {32'hc1ed16d8, 32'hc25ed050} /* (9, 0, 6) {real, imag} */,
  {32'hc18d28c4, 32'h3d189c00} /* (9, 0, 5) {real, imag} */,
  {32'h411f3da0, 32'hc218a23e} /* (9, 0, 4) {real, imag} */,
  {32'h41e68cc8, 32'hc1364aca} /* (9, 0, 3) {real, imag} */,
  {32'hc01b7338, 32'h42da62a5} /* (9, 0, 2) {real, imag} */,
  {32'hc100d040, 32'hc2d0c5b4} /* (9, 0, 1) {real, imag} */,
  {32'h4373f914, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'hc27650ea, 32'hc19b964b} /* (8, 15, 15) {real, imag} */,
  {32'h426d3b23, 32'hc22359ac} /* (8, 15, 14) {real, imag} */,
  {32'hc127cac3, 32'hc0a96f1c} /* (8, 15, 13) {real, imag} */,
  {32'h41138378, 32'hbfc0a3ec} /* (8, 15, 12) {real, imag} */,
  {32'hc05f21b0, 32'hc234f0ba} /* (8, 15, 11) {real, imag} */,
  {32'hc1bbca2e, 32'hc0dd78b2} /* (8, 15, 10) {real, imag} */,
  {32'h40d216b2, 32'h412f59ce} /* (8, 15, 9) {real, imag} */,
  {32'hbfd7dd60, 32'h41946720} /* (8, 15, 8) {real, imag} */,
  {32'h42083cfc, 32'h4144fcc7} /* (8, 15, 7) {real, imag} */,
  {32'h409ff782, 32'hc1824636} /* (8, 15, 6) {real, imag} */,
  {32'h406d9b98, 32'h41ba1be4} /* (8, 15, 5) {real, imag} */,
  {32'hc195bed8, 32'h41140b4a} /* (8, 15, 4) {real, imag} */,
  {32'h41ca3ad2, 32'h41f0d250} /* (8, 15, 3) {real, imag} */,
  {32'hc288aabe, 32'hc25df78e} /* (8, 15, 2) {real, imag} */,
  {32'hc1a9e8e1, 32'hc202d607} /* (8, 15, 1) {real, imag} */,
  {32'hc28197b0, 32'hc236a9c0} /* (8, 15, 0) {real, imag} */,
  {32'hc2abebe0, 32'hc235ffbd} /* (8, 14, 15) {real, imag} */,
  {32'hc2019256, 32'h41b57f52} /* (8, 14, 14) {real, imag} */,
  {32'h420618bb, 32'h40c60a20} /* (8, 14, 13) {real, imag} */,
  {32'h41370c46, 32'hc0bc9a7b} /* (8, 14, 12) {real, imag} */,
  {32'hc128e2aa, 32'h41839f9e} /* (8, 14, 11) {real, imag} */,
  {32'h40beee0f, 32'hc1aaf372} /* (8, 14, 10) {real, imag} */,
  {32'hc1181c5b, 32'hc0b7746a} /* (8, 14, 9) {real, imag} */,
  {32'hbf8f1ce8, 32'hc06b2cca} /* (8, 14, 8) {real, imag} */,
  {32'hc1a41a3d, 32'hc1260640} /* (8, 14, 7) {real, imag} */,
  {32'h40fcfa2c, 32'h4050cfca} /* (8, 14, 6) {real, imag} */,
  {32'hc19054ca, 32'h41a37754} /* (8, 14, 5) {real, imag} */,
  {32'h4109ee07, 32'hc18aab09} /* (8, 14, 4) {real, imag} */,
  {32'h40893155, 32'hc26b70fd} /* (8, 14, 3) {real, imag} */,
  {32'h41ded4f2, 32'h41feaafb} /* (8, 14, 2) {real, imag} */,
  {32'h4293e829, 32'h416e3ba8} /* (8, 14, 1) {real, imag} */,
  {32'hc131873b, 32'h414c183e} /* (8, 14, 0) {real, imag} */,
  {32'h40b35b50, 32'hc161dc62} /* (8, 13, 15) {real, imag} */,
  {32'hc0b494fb, 32'h41cba1ca} /* (8, 13, 14) {real, imag} */,
  {32'hc1e8bb72, 32'hc1b76fc2} /* (8, 13, 13) {real, imag} */,
  {32'hc0f50c08, 32'h41d40f6e} /* (8, 13, 12) {real, imag} */,
  {32'h42165b4e, 32'h3ef5fed0} /* (8, 13, 11) {real, imag} */,
  {32'h40dca578, 32'hc19b69d3} /* (8, 13, 10) {real, imag} */,
  {32'h3f1ff690, 32'hbf8c8498} /* (8, 13, 9) {real, imag} */,
  {32'hc199d948, 32'h4131d8c7} /* (8, 13, 8) {real, imag} */,
  {32'h3ffbdf04, 32'h417df9a8} /* (8, 13, 7) {real, imag} */,
  {32'hc0abb572, 32'hc1b52fee} /* (8, 13, 6) {real, imag} */,
  {32'hc1565c94, 32'hc17c8826} /* (8, 13, 5) {real, imag} */,
  {32'hc10a7a6a, 32'hc0e42dcd} /* (8, 13, 4) {real, imag} */,
  {32'hc2120010, 32'h422653fc} /* (8, 13, 3) {real, imag} */,
  {32'h4139a909, 32'hbf3ddc98} /* (8, 13, 2) {real, imag} */,
  {32'hc0aeaed6, 32'hc20512d7} /* (8, 13, 1) {real, imag} */,
  {32'h419d9a68, 32'hc1ea49d2} /* (8, 13, 0) {real, imag} */,
  {32'hc20a81f9, 32'hc21b3e68} /* (8, 12, 15) {real, imag} */,
  {32'h40cdcf1e, 32'hc2057f1e} /* (8, 12, 14) {real, imag} */,
  {32'hc1fa425f, 32'h41ec27dd} /* (8, 12, 13) {real, imag} */,
  {32'hc1a8917a, 32'h419f2320} /* (8, 12, 12) {real, imag} */,
  {32'h4264042e, 32'h41f21644} /* (8, 12, 11) {real, imag} */,
  {32'hc13581ab, 32'hc1f1a7ee} /* (8, 12, 10) {real, imag} */,
  {32'h41ac2a14, 32'h419804b9} /* (8, 12, 9) {real, imag} */,
  {32'hbfe9009c, 32'h40ee1506} /* (8, 12, 8) {real, imag} */,
  {32'h409d46e7, 32'hc13dc01f} /* (8, 12, 7) {real, imag} */,
  {32'hc17b1a4c, 32'h4163d795} /* (8, 12, 6) {real, imag} */,
  {32'h41ad5c0c, 32'hc2242f31} /* (8, 12, 5) {real, imag} */,
  {32'h42303566, 32'hc03d2164} /* (8, 12, 4) {real, imag} */,
  {32'hc20df5f7, 32'hc061ed28} /* (8, 12, 3) {real, imag} */,
  {32'hc125992f, 32'hc104fffc} /* (8, 12, 2) {real, imag} */,
  {32'h41f121b0, 32'h4175f346} /* (8, 12, 1) {real, imag} */,
  {32'h41512d55, 32'h40fe191e} /* (8, 12, 0) {real, imag} */,
  {32'hc1382adc, 32'hbeb8a680} /* (8, 11, 15) {real, imag} */,
  {32'h419f921a, 32'h418d2b80} /* (8, 11, 14) {real, imag} */,
  {32'hc0d11b09, 32'hc1522d15} /* (8, 11, 13) {real, imag} */,
  {32'h415627bb, 32'h41767ace} /* (8, 11, 12) {real, imag} */,
  {32'h41127db6, 32'hbff34b14} /* (8, 11, 11) {real, imag} */,
  {32'hc0efa462, 32'hc015763e} /* (8, 11, 10) {real, imag} */,
  {32'hc18037ae, 32'h41099786} /* (8, 11, 9) {real, imag} */,
  {32'h418b2b2e, 32'h3ff78dd9} /* (8, 11, 8) {real, imag} */,
  {32'h40ae1608, 32'h418f5b9a} /* (8, 11, 7) {real, imag} */,
  {32'h3fb65ad4, 32'h40411528} /* (8, 11, 6) {real, imag} */,
  {32'hc20962cc, 32'h420caaef} /* (8, 11, 5) {real, imag} */,
  {32'h41a56004, 32'hc094e3a6} /* (8, 11, 4) {real, imag} */,
  {32'h3fd94bf8, 32'hc2419fd0} /* (8, 11, 3) {real, imag} */,
  {32'hc16f7f78, 32'h416aad80} /* (8, 11, 2) {real, imag} */,
  {32'hc22d1036, 32'hc1eea46c} /* (8, 11, 1) {real, imag} */,
  {32'h420c75bd, 32'h4135722c} /* (8, 11, 0) {real, imag} */,
  {32'h411821b4, 32'h418affba} /* (8, 10, 15) {real, imag} */,
  {32'h4145298a, 32'hc184be90} /* (8, 10, 14) {real, imag} */,
  {32'h4130a777, 32'h4049b5e0} /* (8, 10, 13) {real, imag} */,
  {32'h419f91ea, 32'h3fcb06c8} /* (8, 10, 12) {real, imag} */,
  {32'hc201d378, 32'hc1c8cf24} /* (8, 10, 11) {real, imag} */,
  {32'h41591f33, 32'hc18e0d57} /* (8, 10, 10) {real, imag} */,
  {32'hc146d382, 32'h40a7b8e8} /* (8, 10, 9) {real, imag} */,
  {32'hc090a4e8, 32'hc1b1518e} /* (8, 10, 8) {real, imag} */,
  {32'h413e36ae, 32'h40fb80ae} /* (8, 10, 7) {real, imag} */,
  {32'h41921687, 32'h419d6806} /* (8, 10, 6) {real, imag} */,
  {32'hc1c42b1a, 32'hc11e9779} /* (8, 10, 5) {real, imag} */,
  {32'h3ec92cd0, 32'hc1037680} /* (8, 10, 4) {real, imag} */,
  {32'h4198958a, 32'hc1fcc70c} /* (8, 10, 3) {real, imag} */,
  {32'hc0b5e188, 32'h418b8c1c} /* (8, 10, 2) {real, imag} */,
  {32'hc0612f02, 32'hc1414079} /* (8, 10, 1) {real, imag} */,
  {32'hc18728e8, 32'hc16a12cc} /* (8, 10, 0) {real, imag} */,
  {32'h3fbbcb38, 32'h40bb45b1} /* (8, 9, 15) {real, imag} */,
  {32'hc11cf704, 32'hc08ff7e9} /* (8, 9, 14) {real, imag} */,
  {32'hc24c425c, 32'hc1c8ecbb} /* (8, 9, 13) {real, imag} */,
  {32'hbef79400, 32'hc20fdaee} /* (8, 9, 12) {real, imag} */,
  {32'h42309964, 32'h41164c08} /* (8, 9, 11) {real, imag} */,
  {32'h410e31da, 32'h4102219b} /* (8, 9, 10) {real, imag} */,
  {32'hc0f983ca, 32'h40e6fdcc} /* (8, 9, 9) {real, imag} */,
  {32'h418a04e6, 32'h41352be8} /* (8, 9, 8) {real, imag} */,
  {32'h41c779a6, 32'hc13bc8e9} /* (8, 9, 7) {real, imag} */,
  {32'hc0b04be8, 32'hbf920b74} /* (8, 9, 6) {real, imag} */,
  {32'hc0ec217c, 32'hc12beb6f} /* (8, 9, 5) {real, imag} */,
  {32'hc1c361ef, 32'h41dfe2af} /* (8, 9, 4) {real, imag} */,
  {32'h41720298, 32'h40f00082} /* (8, 9, 3) {real, imag} */,
  {32'hc0b20223, 32'h40215c7c} /* (8, 9, 2) {real, imag} */,
  {32'hc1978649, 32'h409b117a} /* (8, 9, 1) {real, imag} */,
  {32'h4175875a, 32'h4140e708} /* (8, 9, 0) {real, imag} */,
  {32'h417bf736, 32'h41176adc} /* (8, 8, 15) {real, imag} */,
  {32'hc065ad14, 32'hc100914f} /* (8, 8, 14) {real, imag} */,
  {32'hc1cb7a5e, 32'h4115b68a} /* (8, 8, 13) {real, imag} */,
  {32'hc16997f8, 32'hbf6a4ff0} /* (8, 8, 12) {real, imag} */,
  {32'hc1545ecf, 32'h416ea371} /* (8, 8, 11) {real, imag} */,
  {32'h425687e0, 32'hbf75a4a8} /* (8, 8, 10) {real, imag} */,
  {32'hc17d3d92, 32'hc1134fa4} /* (8, 8, 9) {real, imag} */,
  {32'hc065df32, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'hc17d3d92, 32'h41134fa4} /* (8, 8, 7) {real, imag} */,
  {32'h425687e0, 32'h3f75a4a8} /* (8, 8, 6) {real, imag} */,
  {32'hc1545ecf, 32'hc16ea371} /* (8, 8, 5) {real, imag} */,
  {32'hc16997f8, 32'h3f6a4ff0} /* (8, 8, 4) {real, imag} */,
  {32'hc1cb7a5e, 32'hc115b68a} /* (8, 8, 3) {real, imag} */,
  {32'hc065ad14, 32'h4100914f} /* (8, 8, 2) {real, imag} */,
  {32'h417bf736, 32'hc1176adc} /* (8, 8, 1) {real, imag} */,
  {32'hc10053d8, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'hc1978649, 32'hc09b117a} /* (8, 7, 15) {real, imag} */,
  {32'hc0b20223, 32'hc0215c7c} /* (8, 7, 14) {real, imag} */,
  {32'h41720298, 32'hc0f00082} /* (8, 7, 13) {real, imag} */,
  {32'hc1c361ef, 32'hc1dfe2af} /* (8, 7, 12) {real, imag} */,
  {32'hc0ec217c, 32'h412beb6f} /* (8, 7, 11) {real, imag} */,
  {32'hc0b04be8, 32'h3f920b74} /* (8, 7, 10) {real, imag} */,
  {32'h41c779a6, 32'h413bc8e9} /* (8, 7, 9) {real, imag} */,
  {32'h418a04e6, 32'hc1352be8} /* (8, 7, 8) {real, imag} */,
  {32'hc0f983ca, 32'hc0e6fdcc} /* (8, 7, 7) {real, imag} */,
  {32'h410e31da, 32'hc102219b} /* (8, 7, 6) {real, imag} */,
  {32'h42309964, 32'hc1164c08} /* (8, 7, 5) {real, imag} */,
  {32'hbef79400, 32'h420fdaee} /* (8, 7, 4) {real, imag} */,
  {32'hc24c425c, 32'h41c8ecbb} /* (8, 7, 3) {real, imag} */,
  {32'hc11cf704, 32'h408ff7e9} /* (8, 7, 2) {real, imag} */,
  {32'h3fbbcb38, 32'hc0bb45b1} /* (8, 7, 1) {real, imag} */,
  {32'h4175875a, 32'hc140e708} /* (8, 7, 0) {real, imag} */,
  {32'hc0612f02, 32'h41414079} /* (8, 6, 15) {real, imag} */,
  {32'hc0b5e188, 32'hc18b8c1c} /* (8, 6, 14) {real, imag} */,
  {32'h4198958a, 32'h41fcc70c} /* (8, 6, 13) {real, imag} */,
  {32'h3ec92cd0, 32'h41037680} /* (8, 6, 12) {real, imag} */,
  {32'hc1c42b1a, 32'h411e9779} /* (8, 6, 11) {real, imag} */,
  {32'h41921687, 32'hc19d6806} /* (8, 6, 10) {real, imag} */,
  {32'h413e36ae, 32'hc0fb80ae} /* (8, 6, 9) {real, imag} */,
  {32'hc090a4e8, 32'h41b1518e} /* (8, 6, 8) {real, imag} */,
  {32'hc146d382, 32'hc0a7b8e8} /* (8, 6, 7) {real, imag} */,
  {32'h41591f33, 32'h418e0d57} /* (8, 6, 6) {real, imag} */,
  {32'hc201d378, 32'h41c8cf24} /* (8, 6, 5) {real, imag} */,
  {32'h419f91ea, 32'hbfcb06c8} /* (8, 6, 4) {real, imag} */,
  {32'h4130a777, 32'hc049b5e0} /* (8, 6, 3) {real, imag} */,
  {32'h4145298a, 32'h4184be90} /* (8, 6, 2) {real, imag} */,
  {32'h411821b4, 32'hc18affba} /* (8, 6, 1) {real, imag} */,
  {32'hc18728e8, 32'h416a12cc} /* (8, 6, 0) {real, imag} */,
  {32'hc22d1036, 32'h41eea46c} /* (8, 5, 15) {real, imag} */,
  {32'hc16f7f78, 32'hc16aad80} /* (8, 5, 14) {real, imag} */,
  {32'h3fd94bf8, 32'h42419fd0} /* (8, 5, 13) {real, imag} */,
  {32'h41a56004, 32'h4094e3a6} /* (8, 5, 12) {real, imag} */,
  {32'hc20962cc, 32'hc20caaef} /* (8, 5, 11) {real, imag} */,
  {32'h3fb65ad4, 32'hc0411528} /* (8, 5, 10) {real, imag} */,
  {32'h40ae1608, 32'hc18f5b9a} /* (8, 5, 9) {real, imag} */,
  {32'h418b2b2e, 32'hbff78dd9} /* (8, 5, 8) {real, imag} */,
  {32'hc18037ae, 32'hc1099786} /* (8, 5, 7) {real, imag} */,
  {32'hc0efa462, 32'h4015763e} /* (8, 5, 6) {real, imag} */,
  {32'h41127db6, 32'h3ff34b14} /* (8, 5, 5) {real, imag} */,
  {32'h415627bb, 32'hc1767ace} /* (8, 5, 4) {real, imag} */,
  {32'hc0d11b09, 32'h41522d15} /* (8, 5, 3) {real, imag} */,
  {32'h419f921a, 32'hc18d2b80} /* (8, 5, 2) {real, imag} */,
  {32'hc1382adc, 32'h3eb8a680} /* (8, 5, 1) {real, imag} */,
  {32'h420c75bd, 32'hc135722c} /* (8, 5, 0) {real, imag} */,
  {32'h41f121b0, 32'hc175f346} /* (8, 4, 15) {real, imag} */,
  {32'hc125992f, 32'h4104fffc} /* (8, 4, 14) {real, imag} */,
  {32'hc20df5f7, 32'h4061ed28} /* (8, 4, 13) {real, imag} */,
  {32'h42303566, 32'h403d2164} /* (8, 4, 12) {real, imag} */,
  {32'h41ad5c0c, 32'h42242f31} /* (8, 4, 11) {real, imag} */,
  {32'hc17b1a4c, 32'hc163d795} /* (8, 4, 10) {real, imag} */,
  {32'h409d46e7, 32'h413dc01f} /* (8, 4, 9) {real, imag} */,
  {32'hbfe9009c, 32'hc0ee1506} /* (8, 4, 8) {real, imag} */,
  {32'h41ac2a14, 32'hc19804b9} /* (8, 4, 7) {real, imag} */,
  {32'hc13581ab, 32'h41f1a7ee} /* (8, 4, 6) {real, imag} */,
  {32'h4264042e, 32'hc1f21644} /* (8, 4, 5) {real, imag} */,
  {32'hc1a8917a, 32'hc19f2320} /* (8, 4, 4) {real, imag} */,
  {32'hc1fa425f, 32'hc1ec27dd} /* (8, 4, 3) {real, imag} */,
  {32'h40cdcf1e, 32'h42057f1e} /* (8, 4, 2) {real, imag} */,
  {32'hc20a81f9, 32'h421b3e68} /* (8, 4, 1) {real, imag} */,
  {32'h41512d55, 32'hc0fe191e} /* (8, 4, 0) {real, imag} */,
  {32'hc0aeaed6, 32'h420512d7} /* (8, 3, 15) {real, imag} */,
  {32'h4139a909, 32'h3f3ddc98} /* (8, 3, 14) {real, imag} */,
  {32'hc2120010, 32'hc22653fc} /* (8, 3, 13) {real, imag} */,
  {32'hc10a7a6a, 32'h40e42dcd} /* (8, 3, 12) {real, imag} */,
  {32'hc1565c94, 32'h417c8826} /* (8, 3, 11) {real, imag} */,
  {32'hc0abb572, 32'h41b52fee} /* (8, 3, 10) {real, imag} */,
  {32'h3ffbdf04, 32'hc17df9a8} /* (8, 3, 9) {real, imag} */,
  {32'hc199d948, 32'hc131d8c7} /* (8, 3, 8) {real, imag} */,
  {32'h3f1ff690, 32'h3f8c8498} /* (8, 3, 7) {real, imag} */,
  {32'h40dca578, 32'h419b69d3} /* (8, 3, 6) {real, imag} */,
  {32'h42165b4e, 32'hbef5fed0} /* (8, 3, 5) {real, imag} */,
  {32'hc0f50c08, 32'hc1d40f6e} /* (8, 3, 4) {real, imag} */,
  {32'hc1e8bb72, 32'h41b76fc2} /* (8, 3, 3) {real, imag} */,
  {32'hc0b494fb, 32'hc1cba1ca} /* (8, 3, 2) {real, imag} */,
  {32'h40b35b50, 32'h4161dc62} /* (8, 3, 1) {real, imag} */,
  {32'h419d9a68, 32'h41ea49d2} /* (8, 3, 0) {real, imag} */,
  {32'h4293e829, 32'hc16e3ba8} /* (8, 2, 15) {real, imag} */,
  {32'h41ded4f2, 32'hc1feaafb} /* (8, 2, 14) {real, imag} */,
  {32'h40893155, 32'h426b70fd} /* (8, 2, 13) {real, imag} */,
  {32'h4109ee07, 32'h418aab09} /* (8, 2, 12) {real, imag} */,
  {32'hc19054ca, 32'hc1a37754} /* (8, 2, 11) {real, imag} */,
  {32'h40fcfa2c, 32'hc050cfca} /* (8, 2, 10) {real, imag} */,
  {32'hc1a41a3d, 32'h41260640} /* (8, 2, 9) {real, imag} */,
  {32'hbf8f1ce8, 32'h406b2cca} /* (8, 2, 8) {real, imag} */,
  {32'hc1181c5b, 32'h40b7746a} /* (8, 2, 7) {real, imag} */,
  {32'h40beee0f, 32'h41aaf372} /* (8, 2, 6) {real, imag} */,
  {32'hc128e2aa, 32'hc1839f9e} /* (8, 2, 5) {real, imag} */,
  {32'h41370c46, 32'h40bc9a7b} /* (8, 2, 4) {real, imag} */,
  {32'h420618bb, 32'hc0c60a20} /* (8, 2, 3) {real, imag} */,
  {32'hc2019256, 32'hc1b57f52} /* (8, 2, 2) {real, imag} */,
  {32'hc2abebe0, 32'h4235ffbd} /* (8, 2, 1) {real, imag} */,
  {32'hc131873b, 32'hc14c183e} /* (8, 2, 0) {real, imag} */,
  {32'hc1a9e8e1, 32'h4202d607} /* (8, 1, 15) {real, imag} */,
  {32'hc288aabe, 32'h425df78e} /* (8, 1, 14) {real, imag} */,
  {32'h41ca3ad2, 32'hc1f0d250} /* (8, 1, 13) {real, imag} */,
  {32'hc195bed8, 32'hc1140b4a} /* (8, 1, 12) {real, imag} */,
  {32'h406d9b98, 32'hc1ba1be4} /* (8, 1, 11) {real, imag} */,
  {32'h409ff782, 32'h41824636} /* (8, 1, 10) {real, imag} */,
  {32'h42083cfc, 32'hc144fcc7} /* (8, 1, 9) {real, imag} */,
  {32'hbfd7dd60, 32'hc1946720} /* (8, 1, 8) {real, imag} */,
  {32'h40d216b2, 32'hc12f59ce} /* (8, 1, 7) {real, imag} */,
  {32'hc1bbca2e, 32'h40dd78b2} /* (8, 1, 6) {real, imag} */,
  {32'hc05f21b0, 32'h4234f0ba} /* (8, 1, 5) {real, imag} */,
  {32'h41138378, 32'h3fc0a3ec} /* (8, 1, 4) {real, imag} */,
  {32'hc127cac3, 32'h40a96f1c} /* (8, 1, 3) {real, imag} */,
  {32'h426d3b23, 32'h422359ac} /* (8, 1, 2) {real, imag} */,
  {32'hc27650ea, 32'h419b964b} /* (8, 1, 1) {real, imag} */,
  {32'hc28197b0, 32'h4236a9c0} /* (8, 1, 0) {real, imag} */,
  {32'hc287cf04, 32'h42bb89fc} /* (8, 0, 15) {real, imag} */,
  {32'hc1d4a362, 32'hc2b751b2} /* (8, 0, 14) {real, imag} */,
  {32'h4202fbf6, 32'h40b85572} /* (8, 0, 13) {real, imag} */,
  {32'hc084a4ae, 32'h42015a03} /* (8, 0, 12) {real, imag} */,
  {32'hc07457f8, 32'hc225f70c} /* (8, 0, 11) {real, imag} */,
  {32'hc16f553c, 32'h41ff001a} /* (8, 0, 10) {real, imag} */,
  {32'hbf9c9fa8, 32'hc10c366c} /* (8, 0, 9) {real, imag} */,
  {32'h4135e4da, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hbf9c9fa8, 32'h410c366c} /* (8, 0, 7) {real, imag} */,
  {32'hc16f553c, 32'hc1ff001a} /* (8, 0, 6) {real, imag} */,
  {32'hc07457f8, 32'h4225f70c} /* (8, 0, 5) {real, imag} */,
  {32'hc084a4ae, 32'hc2015a03} /* (8, 0, 4) {real, imag} */,
  {32'h4202fbf6, 32'hc0b85572} /* (8, 0, 3) {real, imag} */,
  {32'hc1d4a362, 32'h42b751b2} /* (8, 0, 2) {real, imag} */,
  {32'hc287cf04, 32'hc2bb89fc} /* (8, 0, 1) {real, imag} */,
  {32'h42cc4e64, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h41906432, 32'hc299cc79} /* (7, 15, 15) {real, imag} */,
  {32'h421b3c95, 32'hc2c5be56} /* (7, 15, 14) {real, imag} */,
  {32'h419d75b2, 32'h42247f63} /* (7, 15, 13) {real, imag} */,
  {32'hc145c1d6, 32'h3fe83218} /* (7, 15, 12) {real, imag} */,
  {32'hc112cafe, 32'hc09289dc} /* (7, 15, 11) {real, imag} */,
  {32'hc1405733, 32'h40cee7a4} /* (7, 15, 10) {real, imag} */,
  {32'h418e89c5, 32'h4121c4b2} /* (7, 15, 9) {real, imag} */,
  {32'h41266fb0, 32'hc0935ed0} /* (7, 15, 8) {real, imag} */,
  {32'hc0d8c3c0, 32'hc081dd5e} /* (7, 15, 7) {real, imag} */,
  {32'h40aec653, 32'hc105e7fa} /* (7, 15, 6) {real, imag} */,
  {32'h4110c703, 32'h418b1730} /* (7, 15, 5) {real, imag} */,
  {32'hbf8b9e70, 32'h4205dd74} /* (7, 15, 4) {real, imag} */,
  {32'h40b8ef78, 32'h413c88dd} /* (7, 15, 3) {real, imag} */,
  {32'hc241e1f0, 32'h414a50e0} /* (7, 15, 2) {real, imag} */,
  {32'hc208817f, 32'hc233fb2a} /* (7, 15, 1) {real, imag} */,
  {32'hc28f7b5e, 32'hc281abef} /* (7, 15, 0) {real, imag} */,
  {32'hbffba540, 32'h412deb3d} /* (7, 14, 15) {real, imag} */,
  {32'h418742e0, 32'hc213c13e} /* (7, 14, 14) {real, imag} */,
  {32'h422ac872, 32'hc106871a} /* (7, 14, 13) {real, imag} */,
  {32'hc0f28100, 32'hc1ad197b} /* (7, 14, 12) {real, imag} */,
  {32'hc0c2e5b0, 32'h413967bd} /* (7, 14, 11) {real, imag} */,
  {32'h41f1e772, 32'hc1d73d7a} /* (7, 14, 10) {real, imag} */,
  {32'hc20274cc, 32'h41f9b61f} /* (7, 14, 9) {real, imag} */,
  {32'hbea41828, 32'h4008216f} /* (7, 14, 8) {real, imag} */,
  {32'h4028a0e8, 32'hc0d50ff8} /* (7, 14, 7) {real, imag} */,
  {32'hc2117c90, 32'h418abbb0} /* (7, 14, 6) {real, imag} */,
  {32'h411f43ea, 32'h41a575ba} /* (7, 14, 5) {real, imag} */,
  {32'hc1541545, 32'h4202d0b6} /* (7, 14, 4) {real, imag} */,
  {32'hc0c40848, 32'hc229fff9} /* (7, 14, 3) {real, imag} */,
  {32'hc0ee47e0, 32'hc2a657a7} /* (7, 14, 2) {real, imag} */,
  {32'h41cf5ca4, 32'h413f80a0} /* (7, 14, 1) {real, imag} */,
  {32'hc17a118d, 32'h426e8682} /* (7, 14, 0) {real, imag} */,
  {32'h3f670820, 32'h41d45fa6} /* (7, 13, 15) {real, imag} */,
  {32'h40a04c4c, 32'h419e4c0a} /* (7, 13, 14) {real, imag} */,
  {32'h3fbc295c, 32'hc23a1e4c} /* (7, 13, 13) {real, imag} */,
  {32'h4229bc89, 32'h410e8e8c} /* (7, 13, 12) {real, imag} */,
  {32'h42057dbc, 32'h425c98e4} /* (7, 13, 11) {real, imag} */,
  {32'h3fb59fe8, 32'hc1ee5bf6} /* (7, 13, 10) {real, imag} */,
  {32'h41186f8b, 32'hc12ffba8} /* (7, 13, 9) {real, imag} */,
  {32'h4064e930, 32'h41e43023} /* (7, 13, 8) {real, imag} */,
  {32'h415d9bba, 32'h41350eca} /* (7, 13, 7) {real, imag} */,
  {32'hc21e6324, 32'hc0efeeb5} /* (7, 13, 6) {real, imag} */,
  {32'hc0ce5da0, 32'h40263f00} /* (7, 13, 5) {real, imag} */,
  {32'hc02e7934, 32'h40979cba} /* (7, 13, 4) {real, imag} */,
  {32'hc13fa45c, 32'h414cd528} /* (7, 13, 3) {real, imag} */,
  {32'h41a05a77, 32'hc1a88a61} /* (7, 13, 2) {real, imag} */,
  {32'hc13e37ec, 32'hc1d46250} /* (7, 13, 1) {real, imag} */,
  {32'hc08b10b4, 32'hc25001da} /* (7, 13, 0) {real, imag} */,
  {32'hc1eacd9f, 32'hc1457f34} /* (7, 12, 15) {real, imag} */,
  {32'hc117207c, 32'h414e6868} /* (7, 12, 14) {real, imag} */,
  {32'hbfea400c, 32'h4167a882} /* (7, 12, 13) {real, imag} */,
  {32'hc0ab4b91, 32'h4228bb92} /* (7, 12, 12) {real, imag} */,
  {32'h420e777e, 32'hc14fcb60} /* (7, 12, 11) {real, imag} */,
  {32'hc219681e, 32'hbfb137a8} /* (7, 12, 10) {real, imag} */,
  {32'h41a4b397, 32'hc161a242} /* (7, 12, 9) {real, imag} */,
  {32'hc0e91be8, 32'h412285df} /* (7, 12, 8) {real, imag} */,
  {32'h414617e8, 32'hc0aa752c} /* (7, 12, 7) {real, imag} */,
  {32'h41c9b936, 32'hc270cf46} /* (7, 12, 6) {real, imag} */,
  {32'hc0a5f93a, 32'h40a1d485} /* (7, 12, 5) {real, imag} */,
  {32'h41d207e4, 32'h418fb043} /* (7, 12, 4) {real, imag} */,
  {32'hc098d3a7, 32'h41881d9e} /* (7, 12, 3) {real, imag} */,
  {32'h41565b6e, 32'hc12f2c96} /* (7, 12, 2) {real, imag} */,
  {32'h41da9a78, 32'h4055a098} /* (7, 12, 1) {real, imag} */,
  {32'h4202520e, 32'h41b94757} /* (7, 12, 0) {real, imag} */,
  {32'hc20fd062, 32'hc1f1a546} /* (7, 11, 15) {real, imag} */,
  {32'hc0dccd74, 32'h41496b5a} /* (7, 11, 14) {real, imag} */,
  {32'h41741a56, 32'hbf9385b0} /* (7, 11, 13) {real, imag} */,
  {32'h41b35f56, 32'h41ac8b0f} /* (7, 11, 12) {real, imag} */,
  {32'h407b121c, 32'h41692851} /* (7, 11, 11) {real, imag} */,
  {32'h41c4141a, 32'h40df6cc8} /* (7, 11, 10) {real, imag} */,
  {32'hc088dfbe, 32'hc148b893} /* (7, 11, 9) {real, imag} */,
  {32'h41c079ae, 32'h411140eb} /* (7, 11, 8) {real, imag} */,
  {32'hc080a052, 32'h41adb6e6} /* (7, 11, 7) {real, imag} */,
  {32'h4150272a, 32'hc1afc5b2} /* (7, 11, 6) {real, imag} */,
  {32'hc1110816, 32'h41973e4f} /* (7, 11, 5) {real, imag} */,
  {32'hc1e1cd84, 32'hc1d320b6} /* (7, 11, 4) {real, imag} */,
  {32'hc1204fae, 32'hc08f81bc} /* (7, 11, 3) {real, imag} */,
  {32'hc0e819c6, 32'hc2498480} /* (7, 11, 2) {real, imag} */,
  {32'hc05fa037, 32'h3e76a6a0} /* (7, 11, 1) {real, imag} */,
  {32'h421a2cd3, 32'h41c4fabb} /* (7, 11, 0) {real, imag} */,
  {32'hc12f5a3a, 32'h4208acf4} /* (7, 10, 15) {real, imag} */,
  {32'h4120fe2a, 32'h41ab4fe8} /* (7, 10, 14) {real, imag} */,
  {32'hc0af02a0, 32'h41845c1a} /* (7, 10, 13) {real, imag} */,
  {32'h40de0d30, 32'h418eac06} /* (7, 10, 12) {real, imag} */,
  {32'hc2022692, 32'hbefb5f80} /* (7, 10, 11) {real, imag} */,
  {32'hc0909384, 32'h41f9f1e3} /* (7, 10, 10) {real, imag} */,
  {32'hc19e639b, 32'h4125f574} /* (7, 10, 9) {real, imag} */,
  {32'h416eb03a, 32'hc047ed58} /* (7, 10, 8) {real, imag} */,
  {32'h4083b028, 32'hc09546c9} /* (7, 10, 7) {real, imag} */,
  {32'h41f14227, 32'h418f63be} /* (7, 10, 6) {real, imag} */,
  {32'h415650d6, 32'hc2148b15} /* (7, 10, 5) {real, imag} */,
  {32'h3fc51188, 32'h3fdc5364} /* (7, 10, 4) {real, imag} */,
  {32'hc13e3a44, 32'h40bd822e} /* (7, 10, 3) {real, imag} */,
  {32'h4102bb6e, 32'h41592b0b} /* (7, 10, 2) {real, imag} */,
  {32'hc023d280, 32'h412303ad} /* (7, 10, 1) {real, imag} */,
  {32'h420b2996, 32'hc1b059a3} /* (7, 10, 0) {real, imag} */,
  {32'h40f5d304, 32'h40e64430} /* (7, 9, 15) {real, imag} */,
  {32'hc0354bb9, 32'h4120f1e4} /* (7, 9, 14) {real, imag} */,
  {32'h41813f68, 32'hc16f32a6} /* (7, 9, 13) {real, imag} */,
  {32'h41901788, 32'hc1a2411e} /* (7, 9, 12) {real, imag} */,
  {32'hc2251d9c, 32'hc1523205} /* (7, 9, 11) {real, imag} */,
  {32'h425a0962, 32'hc03fa8c0} /* (7, 9, 10) {real, imag} */,
  {32'h401e5970, 32'h4176fcc3} /* (7, 9, 9) {real, imag} */,
  {32'hc0c0bf82, 32'hc13dd962} /* (7, 9, 8) {real, imag} */,
  {32'h40746cbf, 32'h41c8dafe} /* (7, 9, 7) {real, imag} */,
  {32'hc201e8b7, 32'h4188aeff} /* (7, 9, 6) {real, imag} */,
  {32'hc0cb96e4, 32'h41b94df2} /* (7, 9, 5) {real, imag} */,
  {32'hc16935c0, 32'hc199a6ef} /* (7, 9, 4) {real, imag} */,
  {32'h40bef68a, 32'hc181c914} /* (7, 9, 3) {real, imag} */,
  {32'hc1220631, 32'hc044fdd4} /* (7, 9, 2) {real, imag} */,
  {32'h41845e08, 32'h414dedd8} /* (7, 9, 1) {real, imag} */,
  {32'hc1e86500, 32'hbe947d88} /* (7, 9, 0) {real, imag} */,
  {32'h401ff23a, 32'h40f09e9d} /* (7, 8, 15) {real, imag} */,
  {32'h41803b96, 32'h41908103} /* (7, 8, 14) {real, imag} */,
  {32'hc166193e, 32'hc122eeaa} /* (7, 8, 13) {real, imag} */,
  {32'h420047f3, 32'h41d1c456} /* (7, 8, 12) {real, imag} */,
  {32'h40d6d200, 32'hc111fcfc} /* (7, 8, 11) {real, imag} */,
  {32'h40d161aa, 32'h40f59a66} /* (7, 8, 10) {real, imag} */,
  {32'h40e13935, 32'hbfb377cc} /* (7, 8, 9) {real, imag} */,
  {32'hc0ba0286, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'h40e13935, 32'h3fb377cc} /* (7, 8, 7) {real, imag} */,
  {32'h40d161aa, 32'hc0f59a66} /* (7, 8, 6) {real, imag} */,
  {32'h40d6d200, 32'h4111fcfc} /* (7, 8, 5) {real, imag} */,
  {32'h420047f3, 32'hc1d1c456} /* (7, 8, 4) {real, imag} */,
  {32'hc166193e, 32'h4122eeaa} /* (7, 8, 3) {real, imag} */,
  {32'h41803b96, 32'hc1908103} /* (7, 8, 2) {real, imag} */,
  {32'h401ff23a, 32'hc0f09e9d} /* (7, 8, 1) {real, imag} */,
  {32'h408dd290, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h41845e08, 32'hc14dedd8} /* (7, 7, 15) {real, imag} */,
  {32'hc1220631, 32'h4044fdd4} /* (7, 7, 14) {real, imag} */,
  {32'h40bef68a, 32'h4181c914} /* (7, 7, 13) {real, imag} */,
  {32'hc16935c0, 32'h4199a6ef} /* (7, 7, 12) {real, imag} */,
  {32'hc0cb96e4, 32'hc1b94df2} /* (7, 7, 11) {real, imag} */,
  {32'hc201e8b7, 32'hc188aeff} /* (7, 7, 10) {real, imag} */,
  {32'h40746cbf, 32'hc1c8dafe} /* (7, 7, 9) {real, imag} */,
  {32'hc0c0bf82, 32'h413dd962} /* (7, 7, 8) {real, imag} */,
  {32'h401e5970, 32'hc176fcc3} /* (7, 7, 7) {real, imag} */,
  {32'h425a0962, 32'h403fa8c0} /* (7, 7, 6) {real, imag} */,
  {32'hc2251d9c, 32'h41523205} /* (7, 7, 5) {real, imag} */,
  {32'h41901788, 32'h41a2411e} /* (7, 7, 4) {real, imag} */,
  {32'h41813f68, 32'h416f32a6} /* (7, 7, 3) {real, imag} */,
  {32'hc0354bb9, 32'hc120f1e4} /* (7, 7, 2) {real, imag} */,
  {32'h40f5d304, 32'hc0e64430} /* (7, 7, 1) {real, imag} */,
  {32'hc1e86500, 32'h3e947d88} /* (7, 7, 0) {real, imag} */,
  {32'hc023d280, 32'hc12303ad} /* (7, 6, 15) {real, imag} */,
  {32'h4102bb6e, 32'hc1592b0b} /* (7, 6, 14) {real, imag} */,
  {32'hc13e3a44, 32'hc0bd822e} /* (7, 6, 13) {real, imag} */,
  {32'h3fc51188, 32'hbfdc5364} /* (7, 6, 12) {real, imag} */,
  {32'h415650d6, 32'h42148b15} /* (7, 6, 11) {real, imag} */,
  {32'h41f14227, 32'hc18f63be} /* (7, 6, 10) {real, imag} */,
  {32'h4083b028, 32'h409546c9} /* (7, 6, 9) {real, imag} */,
  {32'h416eb03a, 32'h4047ed58} /* (7, 6, 8) {real, imag} */,
  {32'hc19e639b, 32'hc125f574} /* (7, 6, 7) {real, imag} */,
  {32'hc0909384, 32'hc1f9f1e3} /* (7, 6, 6) {real, imag} */,
  {32'hc2022692, 32'h3efb5f80} /* (7, 6, 5) {real, imag} */,
  {32'h40de0d30, 32'hc18eac06} /* (7, 6, 4) {real, imag} */,
  {32'hc0af02a0, 32'hc1845c1a} /* (7, 6, 3) {real, imag} */,
  {32'h4120fe2a, 32'hc1ab4fe8} /* (7, 6, 2) {real, imag} */,
  {32'hc12f5a3a, 32'hc208acf4} /* (7, 6, 1) {real, imag} */,
  {32'h420b2996, 32'h41b059a3} /* (7, 6, 0) {real, imag} */,
  {32'hc05fa037, 32'hbe76a6a0} /* (7, 5, 15) {real, imag} */,
  {32'hc0e819c6, 32'h42498480} /* (7, 5, 14) {real, imag} */,
  {32'hc1204fae, 32'h408f81bc} /* (7, 5, 13) {real, imag} */,
  {32'hc1e1cd84, 32'h41d320b6} /* (7, 5, 12) {real, imag} */,
  {32'hc1110816, 32'hc1973e4f} /* (7, 5, 11) {real, imag} */,
  {32'h4150272a, 32'h41afc5b2} /* (7, 5, 10) {real, imag} */,
  {32'hc080a052, 32'hc1adb6e6} /* (7, 5, 9) {real, imag} */,
  {32'h41c079ae, 32'hc11140eb} /* (7, 5, 8) {real, imag} */,
  {32'hc088dfbe, 32'h4148b893} /* (7, 5, 7) {real, imag} */,
  {32'h41c4141a, 32'hc0df6cc8} /* (7, 5, 6) {real, imag} */,
  {32'h407b121c, 32'hc1692851} /* (7, 5, 5) {real, imag} */,
  {32'h41b35f56, 32'hc1ac8b0f} /* (7, 5, 4) {real, imag} */,
  {32'h41741a56, 32'h3f9385b0} /* (7, 5, 3) {real, imag} */,
  {32'hc0dccd74, 32'hc1496b5a} /* (7, 5, 2) {real, imag} */,
  {32'hc20fd062, 32'h41f1a546} /* (7, 5, 1) {real, imag} */,
  {32'h421a2cd3, 32'hc1c4fabb} /* (7, 5, 0) {real, imag} */,
  {32'h41da9a78, 32'hc055a098} /* (7, 4, 15) {real, imag} */,
  {32'h41565b6e, 32'h412f2c96} /* (7, 4, 14) {real, imag} */,
  {32'hc098d3a7, 32'hc1881d9e} /* (7, 4, 13) {real, imag} */,
  {32'h41d207e4, 32'hc18fb043} /* (7, 4, 12) {real, imag} */,
  {32'hc0a5f93a, 32'hc0a1d485} /* (7, 4, 11) {real, imag} */,
  {32'h41c9b936, 32'h4270cf46} /* (7, 4, 10) {real, imag} */,
  {32'h414617e8, 32'h40aa752c} /* (7, 4, 9) {real, imag} */,
  {32'hc0e91be8, 32'hc12285df} /* (7, 4, 8) {real, imag} */,
  {32'h41a4b397, 32'h4161a242} /* (7, 4, 7) {real, imag} */,
  {32'hc219681e, 32'h3fb137a8} /* (7, 4, 6) {real, imag} */,
  {32'h420e777e, 32'h414fcb60} /* (7, 4, 5) {real, imag} */,
  {32'hc0ab4b91, 32'hc228bb92} /* (7, 4, 4) {real, imag} */,
  {32'hbfea400c, 32'hc167a882} /* (7, 4, 3) {real, imag} */,
  {32'hc117207c, 32'hc14e6868} /* (7, 4, 2) {real, imag} */,
  {32'hc1eacd9f, 32'h41457f34} /* (7, 4, 1) {real, imag} */,
  {32'h4202520e, 32'hc1b94757} /* (7, 4, 0) {real, imag} */,
  {32'hc13e37ec, 32'h41d46250} /* (7, 3, 15) {real, imag} */,
  {32'h41a05a77, 32'h41a88a61} /* (7, 3, 14) {real, imag} */,
  {32'hc13fa45c, 32'hc14cd528} /* (7, 3, 13) {real, imag} */,
  {32'hc02e7934, 32'hc0979cba} /* (7, 3, 12) {real, imag} */,
  {32'hc0ce5da0, 32'hc0263f00} /* (7, 3, 11) {real, imag} */,
  {32'hc21e6324, 32'h40efeeb5} /* (7, 3, 10) {real, imag} */,
  {32'h415d9bba, 32'hc1350eca} /* (7, 3, 9) {real, imag} */,
  {32'h4064e930, 32'hc1e43023} /* (7, 3, 8) {real, imag} */,
  {32'h41186f8b, 32'h412ffba8} /* (7, 3, 7) {real, imag} */,
  {32'h3fb59fe8, 32'h41ee5bf6} /* (7, 3, 6) {real, imag} */,
  {32'h42057dbc, 32'hc25c98e4} /* (7, 3, 5) {real, imag} */,
  {32'h4229bc89, 32'hc10e8e8c} /* (7, 3, 4) {real, imag} */,
  {32'h3fbc295c, 32'h423a1e4c} /* (7, 3, 3) {real, imag} */,
  {32'h40a04c4c, 32'hc19e4c0a} /* (7, 3, 2) {real, imag} */,
  {32'h3f670820, 32'hc1d45fa6} /* (7, 3, 1) {real, imag} */,
  {32'hc08b10b4, 32'h425001da} /* (7, 3, 0) {real, imag} */,
  {32'h41cf5ca4, 32'hc13f80a0} /* (7, 2, 15) {real, imag} */,
  {32'hc0ee47e0, 32'h42a657a7} /* (7, 2, 14) {real, imag} */,
  {32'hc0c40848, 32'h4229fff9} /* (7, 2, 13) {real, imag} */,
  {32'hc1541545, 32'hc202d0b6} /* (7, 2, 12) {real, imag} */,
  {32'h411f43ea, 32'hc1a575ba} /* (7, 2, 11) {real, imag} */,
  {32'hc2117c90, 32'hc18abbb0} /* (7, 2, 10) {real, imag} */,
  {32'h4028a0e8, 32'h40d50ff8} /* (7, 2, 9) {real, imag} */,
  {32'hbea41828, 32'hc008216f} /* (7, 2, 8) {real, imag} */,
  {32'hc20274cc, 32'hc1f9b61f} /* (7, 2, 7) {real, imag} */,
  {32'h41f1e772, 32'h41d73d7a} /* (7, 2, 6) {real, imag} */,
  {32'hc0c2e5b0, 32'hc13967bd} /* (7, 2, 5) {real, imag} */,
  {32'hc0f28100, 32'h41ad197b} /* (7, 2, 4) {real, imag} */,
  {32'h422ac872, 32'h4106871a} /* (7, 2, 3) {real, imag} */,
  {32'h418742e0, 32'h4213c13e} /* (7, 2, 2) {real, imag} */,
  {32'hbffba540, 32'hc12deb3d} /* (7, 2, 1) {real, imag} */,
  {32'hc17a118d, 32'hc26e8682} /* (7, 2, 0) {real, imag} */,
  {32'hc208817f, 32'h4233fb2a} /* (7, 1, 15) {real, imag} */,
  {32'hc241e1f0, 32'hc14a50e0} /* (7, 1, 14) {real, imag} */,
  {32'h40b8ef78, 32'hc13c88dd} /* (7, 1, 13) {real, imag} */,
  {32'hbf8b9e70, 32'hc205dd74} /* (7, 1, 12) {real, imag} */,
  {32'h4110c703, 32'hc18b1730} /* (7, 1, 11) {real, imag} */,
  {32'h40aec653, 32'h4105e7fa} /* (7, 1, 10) {real, imag} */,
  {32'hc0d8c3c0, 32'h4081dd5e} /* (7, 1, 9) {real, imag} */,
  {32'h41266fb0, 32'h40935ed0} /* (7, 1, 8) {real, imag} */,
  {32'h418e89c5, 32'hc121c4b2} /* (7, 1, 7) {real, imag} */,
  {32'hc1405733, 32'hc0cee7a4} /* (7, 1, 6) {real, imag} */,
  {32'hc112cafe, 32'h409289dc} /* (7, 1, 5) {real, imag} */,
  {32'hc145c1d6, 32'hbfe83218} /* (7, 1, 4) {real, imag} */,
  {32'h419d75b2, 32'hc2247f63} /* (7, 1, 3) {real, imag} */,
  {32'h421b3c95, 32'h42c5be56} /* (7, 1, 2) {real, imag} */,
  {32'h41906432, 32'h4299cc79} /* (7, 1, 1) {real, imag} */,
  {32'hc28f7b5e, 32'h4281abef} /* (7, 1, 0) {real, imag} */,
  {32'hc2e65d14, 32'h42fc7ac6} /* (7, 0, 15) {real, imag} */,
  {32'hc217eaae, 32'hc2b88883} /* (7, 0, 14) {real, imag} */,
  {32'h4212ea30, 32'hc1e8d7c1} /* (7, 0, 13) {real, imag} */,
  {32'h40ce38f0, 32'h4211a6d6} /* (7, 0, 12) {real, imag} */,
  {32'h40a54a66, 32'hc204ff77} /* (7, 0, 11) {real, imag} */,
  {32'h416edd1f, 32'h41dc52a9} /* (7, 0, 10) {real, imag} */,
  {32'h419eceb6, 32'hc18b4234} /* (7, 0, 9) {real, imag} */,
  {32'hc1c7bb33, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'h419eceb6, 32'h418b4234} /* (7, 0, 7) {real, imag} */,
  {32'h416edd1f, 32'hc1dc52a9} /* (7, 0, 6) {real, imag} */,
  {32'h40a54a66, 32'h4204ff77} /* (7, 0, 5) {real, imag} */,
  {32'h40ce38f0, 32'hc211a6d6} /* (7, 0, 4) {real, imag} */,
  {32'h4212ea30, 32'h41e8d7c1} /* (7, 0, 3) {real, imag} */,
  {32'hc217eaae, 32'h42b88883} /* (7, 0, 2) {real, imag} */,
  {32'hc2e65d14, 32'hc2fc7ac6} /* (7, 0, 1) {real, imag} */,
  {32'h40ea2910, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h41d831e9, 32'hc2cd9354} /* (6, 15, 15) {real, imag} */,
  {32'hc11b2543, 32'hc232a726} /* (6, 15, 14) {real, imag} */,
  {32'hc2116003, 32'h41584797} /* (6, 15, 13) {real, imag} */,
  {32'hc19fefe6, 32'h41db24ab} /* (6, 15, 12) {real, imag} */,
  {32'hc01f54a4, 32'h41a9361e} /* (6, 15, 11) {real, imag} */,
  {32'h41d55d32, 32'h4082f7f8} /* (6, 15, 10) {real, imag} */,
  {32'h4211ae90, 32'h4193beb1} /* (6, 15, 9) {real, imag} */,
  {32'h414afe60, 32'h40abdadf} /* (6, 15, 8) {real, imag} */,
  {32'hc1938b02, 32'h41f26daa} /* (6, 15, 7) {real, imag} */,
  {32'h40690396, 32'h41842d58} /* (6, 15, 6) {real, imag} */,
  {32'h41bc9c4d, 32'hbfe2e7f8} /* (6, 15, 5) {real, imag} */,
  {32'h423d61db, 32'hc25084e0} /* (6, 15, 4) {real, imag} */,
  {32'hc10de4cc, 32'h4013ce70} /* (6, 15, 3) {real, imag} */,
  {32'hc2985cae, 32'h410fcb04} /* (6, 15, 2) {real, imag} */,
  {32'hc28fb836, 32'h40eb5358} /* (6, 15, 1) {real, imag} */,
  {32'hc2c037e4, 32'hc2b35a79} /* (6, 15, 0) {real, imag} */,
  {32'hc19835f2, 32'h4269b690} /* (6, 14, 15) {real, imag} */,
  {32'h41b5f22e, 32'hc205336c} /* (6, 14, 14) {real, imag} */,
  {32'h41a6a6bb, 32'hc24a709e} /* (6, 14, 13) {real, imag} */,
  {32'h40d4568c, 32'h405becd8} /* (6, 14, 12) {real, imag} */,
  {32'h410b4f0c, 32'hc210819d} /* (6, 14, 11) {real, imag} */,
  {32'hc1e63dbe, 32'hc17da9d2} /* (6, 14, 10) {real, imag} */,
  {32'h40c3dfe2, 32'h414b04f5} /* (6, 14, 9) {real, imag} */,
  {32'hc1453c8a, 32'hc102005b} /* (6, 14, 8) {real, imag} */,
  {32'h40cd739d, 32'hc1877002} /* (6, 14, 7) {real, imag} */,
  {32'h3fc01a20, 32'hc153ac3c} /* (6, 14, 6) {real, imag} */,
  {32'hc0d067a6, 32'hbfb119e0} /* (6, 14, 5) {real, imag} */,
  {32'h418122c4, 32'h421dcef0} /* (6, 14, 4) {real, imag} */,
  {32'hc20530c2, 32'hc19977b5} /* (6, 14, 3) {real, imag} */,
  {32'h3f9507a0, 32'hc2a250a7} /* (6, 14, 2) {real, imag} */,
  {32'h41c13c28, 32'hc1707f04} /* (6, 14, 1) {real, imag} */,
  {32'h41d9f946, 32'h42a06e65} /* (6, 14, 0) {real, imag} */,
  {32'hc0efc2a0, 32'h4253f02b} /* (6, 13, 15) {real, imag} */,
  {32'hc16343e1, 32'hc20dc9ff} /* (6, 13, 14) {real, imag} */,
  {32'hc11e6700, 32'hc237b4aa} /* (6, 13, 13) {real, imag} */,
  {32'h420c84a0, 32'hc0da37d8} /* (6, 13, 12) {real, imag} */,
  {32'hc172c207, 32'h4224cd6c} /* (6, 13, 11) {real, imag} */,
  {32'hbf4f84e0, 32'h41da3c18} /* (6, 13, 10) {real, imag} */,
  {32'h401a8a60, 32'h410dcd4c} /* (6, 13, 9) {real, imag} */,
  {32'h414aa02e, 32'h3e019928} /* (6, 13, 8) {real, imag} */,
  {32'hc157b8de, 32'hc17c5bd5} /* (6, 13, 7) {real, imag} */,
  {32'h3eb23580, 32'h40645bf0} /* (6, 13, 6) {real, imag} */,
  {32'h410a70e5, 32'h41f3c709} /* (6, 13, 5) {real, imag} */,
  {32'h41304ac4, 32'hc1f544fa} /* (6, 13, 4) {real, imag} */,
  {32'hc16382c1, 32'h410d8133} /* (6, 13, 3) {real, imag} */,
  {32'hc124f9ed, 32'hc0b9daa7} /* (6, 13, 2) {real, imag} */,
  {32'h42328b61, 32'hc10eaf8c} /* (6, 13, 1) {real, imag} */,
  {32'h4193c0b8, 32'hc25ed294} /* (6, 13, 0) {real, imag} */,
  {32'hc20a6066, 32'hc28fd876} /* (6, 12, 15) {real, imag} */,
  {32'hbfb48900, 32'hc2042ab8} /* (6, 12, 14) {real, imag} */,
  {32'h41a244b2, 32'hc1a27e1c} /* (6, 12, 13) {real, imag} */,
  {32'h3fb4e50e, 32'h422fa231} /* (6, 12, 12) {real, imag} */,
  {32'hc1b111d5, 32'hc0328633} /* (6, 12, 11) {real, imag} */,
  {32'h4123e22a, 32'hc23f0130} /* (6, 12, 10) {real, imag} */,
  {32'h419e62c8, 32'h41882775} /* (6, 12, 9) {real, imag} */,
  {32'h409fa01c, 32'h40a2d0e2} /* (6, 12, 8) {real, imag} */,
  {32'hc15a410f, 32'hc025bfd8} /* (6, 12, 7) {real, imag} */,
  {32'hc18c533e, 32'hc0858170} /* (6, 12, 6) {real, imag} */,
  {32'hc1bc0a29, 32'h412765af} /* (6, 12, 5) {real, imag} */,
  {32'h41620020, 32'hc15991db} /* (6, 12, 4) {real, imag} */,
  {32'hc123e878, 32'h41512a0a} /* (6, 12, 3) {real, imag} */,
  {32'hc079e5cc, 32'h4176f178} /* (6, 12, 2) {real, imag} */,
  {32'hc0dd883f, 32'hc1e5a53a} /* (6, 12, 1) {real, imag} */,
  {32'h4147b4ec, 32'h410c9ff8} /* (6, 12, 0) {real, imag} */,
  {32'hc1103ba6, 32'h41b60794} /* (6, 11, 15) {real, imag} */,
  {32'h4094c544, 32'h41d57b78} /* (6, 11, 14) {real, imag} */,
  {32'h423e264a, 32'hc0a6d540} /* (6, 11, 13) {real, imag} */,
  {32'hc2484ac7, 32'h41d62024} /* (6, 11, 12) {real, imag} */,
  {32'hc179e549, 32'h4207cb72} /* (6, 11, 11) {real, imag} */,
  {32'hbfb6fcb2, 32'hc2453104} /* (6, 11, 10) {real, imag} */,
  {32'hc1c56c7d, 32'hbf0bd410} /* (6, 11, 9) {real, imag} */,
  {32'hc0f7d576, 32'h415a3bba} /* (6, 11, 8) {real, imag} */,
  {32'h41f3c7ce, 32'h411543af} /* (6, 11, 7) {real, imag} */,
  {32'h41937cf7, 32'hc125204e} /* (6, 11, 6) {real, imag} */,
  {32'hc195d698, 32'hc0b52485} /* (6, 11, 5) {real, imag} */,
  {32'h41138e96, 32'hc020026f} /* (6, 11, 4) {real, imag} */,
  {32'hc121b3f4, 32'hc15c3a18} /* (6, 11, 3) {real, imag} */,
  {32'hc10b9dcb, 32'hc24c4c97} /* (6, 11, 2) {real, imag} */,
  {32'h420392b7, 32'h420f369c} /* (6, 11, 1) {real, imag} */,
  {32'h41a18bb7, 32'hc0f9748c} /* (6, 11, 0) {real, imag} */,
  {32'h4196961d, 32'hc1370a1b} /* (6, 10, 15) {real, imag} */,
  {32'hbf61fa80, 32'hc1b0abe3} /* (6, 10, 14) {real, imag} */,
  {32'h41c8fb86, 32'h4109a6f8} /* (6, 10, 13) {real, imag} */,
  {32'hc213ada4, 32'h41593762} /* (6, 10, 12) {real, imag} */,
  {32'hc0731c40, 32'hc2301683} /* (6, 10, 11) {real, imag} */,
  {32'h413eb37f, 32'hc196caf7} /* (6, 10, 10) {real, imag} */,
  {32'h41b6eb02, 32'hbec1a434} /* (6, 10, 9) {real, imag} */,
  {32'hc1898254, 32'h411adda6} /* (6, 10, 8) {real, imag} */,
  {32'h40d639df, 32'hc1ffe7ae} /* (6, 10, 7) {real, imag} */,
  {32'hc095947b, 32'h41cd434a} /* (6, 10, 6) {real, imag} */,
  {32'hc1731478, 32'hc2222381} /* (6, 10, 5) {real, imag} */,
  {32'hbefdd1c0, 32'h41208e05} /* (6, 10, 4) {real, imag} */,
  {32'hbf66b4f0, 32'hbf772c60} /* (6, 10, 3) {real, imag} */,
  {32'hc0cfb63f, 32'h41119d03} /* (6, 10, 2) {real, imag} */,
  {32'hc1088390, 32'h4179f7f8} /* (6, 10, 1) {real, imag} */,
  {32'hc105ad60, 32'h42067d6c} /* (6, 10, 0) {real, imag} */,
  {32'hc15ee1c8, 32'h3fe253bc} /* (6, 9, 15) {real, imag} */,
  {32'hbf7b4cf0, 32'hc10db853} /* (6, 9, 14) {real, imag} */,
  {32'h417b962c, 32'h41476b5a} /* (6, 9, 13) {real, imag} */,
  {32'h40df2247, 32'h41ac65d3} /* (6, 9, 12) {real, imag} */,
  {32'h408db9fc, 32'h40f9b78e} /* (6, 9, 11) {real, imag} */,
  {32'hc0d4255f, 32'h420dde2c} /* (6, 9, 10) {real, imag} */,
  {32'h41931bb9, 32'hc17a93d2} /* (6, 9, 9) {real, imag} */,
  {32'hc10ee1b0, 32'hc137630b} /* (6, 9, 8) {real, imag} */,
  {32'hc1bfc2de, 32'h411a13cb} /* (6, 9, 7) {real, imag} */,
  {32'hc112836b, 32'h41d7b70a} /* (6, 9, 6) {real, imag} */,
  {32'h40526bc4, 32'h4058dea4} /* (6, 9, 5) {real, imag} */,
  {32'h414f84a4, 32'h41d20280} /* (6, 9, 4) {real, imag} */,
  {32'h408de450, 32'hc1d2c16d} /* (6, 9, 3) {real, imag} */,
  {32'h41a16876, 32'hc142f4d6} /* (6, 9, 2) {real, imag} */,
  {32'h411d7fe7, 32'hc1068c92} /* (6, 9, 1) {real, imag} */,
  {32'hbe1dfac0, 32'hc0766b31} /* (6, 9, 0) {real, imag} */,
  {32'hc0d412cf, 32'h3f17398c} /* (6, 8, 15) {real, imag} */,
  {32'hc1458974, 32'h3fec3260} /* (6, 8, 14) {real, imag} */,
  {32'h418e09ea, 32'h408fd527} /* (6, 8, 13) {real, imag} */,
  {32'h412156fb, 32'hc1951e3e} /* (6, 8, 12) {real, imag} */,
  {32'h4178a418, 32'hc124e5c8} /* (6, 8, 11) {real, imag} */,
  {32'hc097d062, 32'h405887e0} /* (6, 8, 10) {real, imag} */,
  {32'hbf644cf0, 32'hc0a1049e} /* (6, 8, 9) {real, imag} */,
  {32'h40a01c64, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'hbf644cf0, 32'h40a1049e} /* (6, 8, 7) {real, imag} */,
  {32'hc097d062, 32'hc05887e0} /* (6, 8, 6) {real, imag} */,
  {32'h4178a418, 32'h4124e5c8} /* (6, 8, 5) {real, imag} */,
  {32'h412156fb, 32'h41951e3e} /* (6, 8, 4) {real, imag} */,
  {32'h418e09ea, 32'hc08fd527} /* (6, 8, 3) {real, imag} */,
  {32'hc1458974, 32'hbfec3260} /* (6, 8, 2) {real, imag} */,
  {32'hc0d412cf, 32'hbf17398c} /* (6, 8, 1) {real, imag} */,
  {32'h410f0836, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h411d7fe7, 32'h41068c92} /* (6, 7, 15) {real, imag} */,
  {32'h41a16876, 32'h4142f4d6} /* (6, 7, 14) {real, imag} */,
  {32'h408de450, 32'h41d2c16d} /* (6, 7, 13) {real, imag} */,
  {32'h414f84a4, 32'hc1d20280} /* (6, 7, 12) {real, imag} */,
  {32'h40526bc4, 32'hc058dea4} /* (6, 7, 11) {real, imag} */,
  {32'hc112836b, 32'hc1d7b70a} /* (6, 7, 10) {real, imag} */,
  {32'hc1bfc2de, 32'hc11a13cb} /* (6, 7, 9) {real, imag} */,
  {32'hc10ee1b0, 32'h4137630b} /* (6, 7, 8) {real, imag} */,
  {32'h41931bb9, 32'h417a93d2} /* (6, 7, 7) {real, imag} */,
  {32'hc0d4255f, 32'hc20dde2c} /* (6, 7, 6) {real, imag} */,
  {32'h408db9fc, 32'hc0f9b78e} /* (6, 7, 5) {real, imag} */,
  {32'h40df2247, 32'hc1ac65d3} /* (6, 7, 4) {real, imag} */,
  {32'h417b962c, 32'hc1476b5a} /* (6, 7, 3) {real, imag} */,
  {32'hbf7b4cf0, 32'h410db853} /* (6, 7, 2) {real, imag} */,
  {32'hc15ee1c8, 32'hbfe253bc} /* (6, 7, 1) {real, imag} */,
  {32'hbe1dfac0, 32'h40766b31} /* (6, 7, 0) {real, imag} */,
  {32'hc1088390, 32'hc179f7f8} /* (6, 6, 15) {real, imag} */,
  {32'hc0cfb63f, 32'hc1119d03} /* (6, 6, 14) {real, imag} */,
  {32'hbf66b4f0, 32'h3f772c60} /* (6, 6, 13) {real, imag} */,
  {32'hbefdd1c0, 32'hc1208e05} /* (6, 6, 12) {real, imag} */,
  {32'hc1731478, 32'h42222381} /* (6, 6, 11) {real, imag} */,
  {32'hc095947b, 32'hc1cd434a} /* (6, 6, 10) {real, imag} */,
  {32'h40d639df, 32'h41ffe7ae} /* (6, 6, 9) {real, imag} */,
  {32'hc1898254, 32'hc11adda6} /* (6, 6, 8) {real, imag} */,
  {32'h41b6eb02, 32'h3ec1a434} /* (6, 6, 7) {real, imag} */,
  {32'h413eb37f, 32'h4196caf7} /* (6, 6, 6) {real, imag} */,
  {32'hc0731c40, 32'h42301683} /* (6, 6, 5) {real, imag} */,
  {32'hc213ada4, 32'hc1593762} /* (6, 6, 4) {real, imag} */,
  {32'h41c8fb86, 32'hc109a6f8} /* (6, 6, 3) {real, imag} */,
  {32'hbf61fa80, 32'h41b0abe3} /* (6, 6, 2) {real, imag} */,
  {32'h4196961d, 32'h41370a1b} /* (6, 6, 1) {real, imag} */,
  {32'hc105ad60, 32'hc2067d6c} /* (6, 6, 0) {real, imag} */,
  {32'h420392b7, 32'hc20f369c} /* (6, 5, 15) {real, imag} */,
  {32'hc10b9dcb, 32'h424c4c97} /* (6, 5, 14) {real, imag} */,
  {32'hc121b3f4, 32'h415c3a18} /* (6, 5, 13) {real, imag} */,
  {32'h41138e96, 32'h4020026f} /* (6, 5, 12) {real, imag} */,
  {32'hc195d698, 32'h40b52485} /* (6, 5, 11) {real, imag} */,
  {32'h41937cf7, 32'h4125204e} /* (6, 5, 10) {real, imag} */,
  {32'h41f3c7ce, 32'hc11543af} /* (6, 5, 9) {real, imag} */,
  {32'hc0f7d576, 32'hc15a3bba} /* (6, 5, 8) {real, imag} */,
  {32'hc1c56c7d, 32'h3f0bd410} /* (6, 5, 7) {real, imag} */,
  {32'hbfb6fcb2, 32'h42453104} /* (6, 5, 6) {real, imag} */,
  {32'hc179e549, 32'hc207cb72} /* (6, 5, 5) {real, imag} */,
  {32'hc2484ac7, 32'hc1d62024} /* (6, 5, 4) {real, imag} */,
  {32'h423e264a, 32'h40a6d540} /* (6, 5, 3) {real, imag} */,
  {32'h4094c544, 32'hc1d57b78} /* (6, 5, 2) {real, imag} */,
  {32'hc1103ba6, 32'hc1b60794} /* (6, 5, 1) {real, imag} */,
  {32'h41a18bb7, 32'h40f9748c} /* (6, 5, 0) {real, imag} */,
  {32'hc0dd883f, 32'h41e5a53a} /* (6, 4, 15) {real, imag} */,
  {32'hc079e5cc, 32'hc176f178} /* (6, 4, 14) {real, imag} */,
  {32'hc123e878, 32'hc1512a0a} /* (6, 4, 13) {real, imag} */,
  {32'h41620020, 32'h415991db} /* (6, 4, 12) {real, imag} */,
  {32'hc1bc0a29, 32'hc12765af} /* (6, 4, 11) {real, imag} */,
  {32'hc18c533e, 32'h40858170} /* (6, 4, 10) {real, imag} */,
  {32'hc15a410f, 32'h4025bfd8} /* (6, 4, 9) {real, imag} */,
  {32'h409fa01c, 32'hc0a2d0e2} /* (6, 4, 8) {real, imag} */,
  {32'h419e62c8, 32'hc1882775} /* (6, 4, 7) {real, imag} */,
  {32'h4123e22a, 32'h423f0130} /* (6, 4, 6) {real, imag} */,
  {32'hc1b111d5, 32'h40328633} /* (6, 4, 5) {real, imag} */,
  {32'h3fb4e50e, 32'hc22fa231} /* (6, 4, 4) {real, imag} */,
  {32'h41a244b2, 32'h41a27e1c} /* (6, 4, 3) {real, imag} */,
  {32'hbfb48900, 32'h42042ab8} /* (6, 4, 2) {real, imag} */,
  {32'hc20a6066, 32'h428fd876} /* (6, 4, 1) {real, imag} */,
  {32'h4147b4ec, 32'hc10c9ff8} /* (6, 4, 0) {real, imag} */,
  {32'h42328b61, 32'h410eaf8c} /* (6, 3, 15) {real, imag} */,
  {32'hc124f9ed, 32'h40b9daa7} /* (6, 3, 14) {real, imag} */,
  {32'hc16382c1, 32'hc10d8133} /* (6, 3, 13) {real, imag} */,
  {32'h41304ac4, 32'h41f544fa} /* (6, 3, 12) {real, imag} */,
  {32'h410a70e5, 32'hc1f3c709} /* (6, 3, 11) {real, imag} */,
  {32'h3eb23580, 32'hc0645bf0} /* (6, 3, 10) {real, imag} */,
  {32'hc157b8de, 32'h417c5bd5} /* (6, 3, 9) {real, imag} */,
  {32'h414aa02e, 32'hbe019928} /* (6, 3, 8) {real, imag} */,
  {32'h401a8a60, 32'hc10dcd4c} /* (6, 3, 7) {real, imag} */,
  {32'hbf4f84e0, 32'hc1da3c18} /* (6, 3, 6) {real, imag} */,
  {32'hc172c207, 32'hc224cd6c} /* (6, 3, 5) {real, imag} */,
  {32'h420c84a0, 32'h40da37d8} /* (6, 3, 4) {real, imag} */,
  {32'hc11e6700, 32'h4237b4aa} /* (6, 3, 3) {real, imag} */,
  {32'hc16343e1, 32'h420dc9ff} /* (6, 3, 2) {real, imag} */,
  {32'hc0efc2a0, 32'hc253f02b} /* (6, 3, 1) {real, imag} */,
  {32'h4193c0b8, 32'h425ed294} /* (6, 3, 0) {real, imag} */,
  {32'h41c13c28, 32'h41707f04} /* (6, 2, 15) {real, imag} */,
  {32'h3f9507a0, 32'h42a250a7} /* (6, 2, 14) {real, imag} */,
  {32'hc20530c2, 32'h419977b5} /* (6, 2, 13) {real, imag} */,
  {32'h418122c4, 32'hc21dcef0} /* (6, 2, 12) {real, imag} */,
  {32'hc0d067a6, 32'h3fb119e0} /* (6, 2, 11) {real, imag} */,
  {32'h3fc01a20, 32'h4153ac3c} /* (6, 2, 10) {real, imag} */,
  {32'h40cd739d, 32'h41877002} /* (6, 2, 9) {real, imag} */,
  {32'hc1453c8a, 32'h4102005b} /* (6, 2, 8) {real, imag} */,
  {32'h40c3dfe2, 32'hc14b04f5} /* (6, 2, 7) {real, imag} */,
  {32'hc1e63dbe, 32'h417da9d2} /* (6, 2, 6) {real, imag} */,
  {32'h410b4f0c, 32'h4210819d} /* (6, 2, 5) {real, imag} */,
  {32'h40d4568c, 32'hc05becd8} /* (6, 2, 4) {real, imag} */,
  {32'h41a6a6bb, 32'h424a709e} /* (6, 2, 3) {real, imag} */,
  {32'h41b5f22e, 32'h4205336c} /* (6, 2, 2) {real, imag} */,
  {32'hc19835f2, 32'hc269b690} /* (6, 2, 1) {real, imag} */,
  {32'h41d9f946, 32'hc2a06e65} /* (6, 2, 0) {real, imag} */,
  {32'hc28fb836, 32'hc0eb5358} /* (6, 1, 15) {real, imag} */,
  {32'hc2985cae, 32'hc10fcb04} /* (6, 1, 14) {real, imag} */,
  {32'hc10de4cc, 32'hc013ce70} /* (6, 1, 13) {real, imag} */,
  {32'h423d61db, 32'h425084e0} /* (6, 1, 12) {real, imag} */,
  {32'h41bc9c4d, 32'h3fe2e7f8} /* (6, 1, 11) {real, imag} */,
  {32'h40690396, 32'hc1842d58} /* (6, 1, 10) {real, imag} */,
  {32'hc1938b02, 32'hc1f26daa} /* (6, 1, 9) {real, imag} */,
  {32'h414afe60, 32'hc0abdadf} /* (6, 1, 8) {real, imag} */,
  {32'h4211ae90, 32'hc193beb1} /* (6, 1, 7) {real, imag} */,
  {32'h41d55d32, 32'hc082f7f8} /* (6, 1, 6) {real, imag} */,
  {32'hc01f54a4, 32'hc1a9361e} /* (6, 1, 5) {real, imag} */,
  {32'hc19fefe6, 32'hc1db24ab} /* (6, 1, 4) {real, imag} */,
  {32'hc2116003, 32'hc1584797} /* (6, 1, 3) {real, imag} */,
  {32'hc11b2543, 32'h4232a726} /* (6, 1, 2) {real, imag} */,
  {32'h41d831e9, 32'h42cd9354} /* (6, 1, 1) {real, imag} */,
  {32'hc2c037e4, 32'h42b35a79} /* (6, 1, 0) {real, imag} */,
  {32'hc28dc9c0, 32'h43147d8c} /* (6, 0, 15) {real, imag} */,
  {32'h41a76f04, 32'hc2541ce5} /* (6, 0, 14) {real, imag} */,
  {32'h4185145b, 32'hc2288d37} /* (6, 0, 13) {real, imag} */,
  {32'hc134a2b5, 32'hc1017d52} /* (6, 0, 12) {real, imag} */,
  {32'hc09bdd98, 32'hc0f18a20} /* (6, 0, 11) {real, imag} */,
  {32'h3ff7e70a, 32'h41c7e50f} /* (6, 0, 10) {real, imag} */,
  {32'hc117af14, 32'hc1896c80} /* (6, 0, 9) {real, imag} */,
  {32'hc0f335c3, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'hc117af14, 32'h41896c80} /* (6, 0, 7) {real, imag} */,
  {32'h3ff7e70a, 32'hc1c7e50f} /* (6, 0, 6) {real, imag} */,
  {32'hc09bdd98, 32'h40f18a20} /* (6, 0, 5) {real, imag} */,
  {32'hc134a2b5, 32'h41017d52} /* (6, 0, 4) {real, imag} */,
  {32'h4185145b, 32'h42288d37} /* (6, 0, 3) {real, imag} */,
  {32'h41a76f04, 32'h42541ce5} /* (6, 0, 2) {real, imag} */,
  {32'hc28dc9c0, 32'hc3147d8c} /* (6, 0, 1) {real, imag} */,
  {32'hc326eafe, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h42448106, 32'hc2df6874} /* (5, 15, 15) {real, imag} */,
  {32'hc1e0fec4, 32'h406b98a4} /* (5, 15, 14) {real, imag} */,
  {32'h40b45ec9, 32'h4225adf1} /* (5, 15, 13) {real, imag} */,
  {32'hc02edfbc, 32'h41684d0c} /* (5, 15, 12) {real, imag} */,
  {32'h4172dd3a, 32'hc1c23111} /* (5, 15, 11) {real, imag} */,
  {32'h41ba21df, 32'h41d3d481} /* (5, 15, 10) {real, imag} */,
  {32'hc09e2a70, 32'hc0c333e8} /* (5, 15, 9) {real, imag} */,
  {32'hc00b0d5a, 32'hc05593da} /* (5, 15, 8) {real, imag} */,
  {32'h41cb79d9, 32'h40a04773} /* (5, 15, 7) {real, imag} */,
  {32'h4141c261, 32'hc1667592} /* (5, 15, 6) {real, imag} */,
  {32'h40ae2c54, 32'hc119181f} /* (5, 15, 5) {real, imag} */,
  {32'h4263f9b4, 32'hc1bc92de} /* (5, 15, 4) {real, imag} */,
  {32'hc21c6d87, 32'hc1c26bfe} /* (5, 15, 3) {real, imag} */,
  {32'hc295ba32, 32'hbf807370} /* (5, 15, 2) {real, imag} */,
  {32'hc2d7a90c, 32'hc1982198} /* (5, 15, 1) {real, imag} */,
  {32'hc28b142b, 32'hc1a307c0} /* (5, 15, 0) {real, imag} */,
  {32'hc02f0420, 32'h422cb651} /* (5, 14, 15) {real, imag} */,
  {32'hc0b5d1f4, 32'hc1aa1f9d} /* (5, 14, 14) {real, imag} */,
  {32'hc1e6f256, 32'hc1c76cde} /* (5, 14, 13) {real, imag} */,
  {32'h419fec4f, 32'h41dd6637} /* (5, 14, 12) {real, imag} */,
  {32'h41cbf47b, 32'hc0fd86e9} /* (5, 14, 11) {real, imag} */,
  {32'hc0e335b6, 32'hc1148e68} /* (5, 14, 10) {real, imag} */,
  {32'h414a5014, 32'hc0d6f3c0} /* (5, 14, 9) {real, imag} */,
  {32'h4121f3c4, 32'hc1f4332a} /* (5, 14, 8) {real, imag} */,
  {32'hc216dee2, 32'hbeb6bae0} /* (5, 14, 7) {real, imag} */,
  {32'hc17fa545, 32'h3fb1cec0} /* (5, 14, 6) {real, imag} */,
  {32'hc083e36c, 32'hc212e32b} /* (5, 14, 5) {real, imag} */,
  {32'h41ec94ba, 32'hc21a598e} /* (5, 14, 4) {real, imag} */,
  {32'h4130e2cc, 32'h417b8d66} /* (5, 14, 3) {real, imag} */,
  {32'h421f82fb, 32'hc2863a22} /* (5, 14, 2) {real, imag} */,
  {32'hc143d1b6, 32'hc1b3bc65} /* (5, 14, 1) {real, imag} */,
  {32'h428bf210, 32'h4256b62d} /* (5, 14, 0) {real, imag} */,
  {32'hc1a6be2a, 32'h41aafe58} /* (5, 13, 15) {real, imag} */,
  {32'hc101cc98, 32'hc18487a2} /* (5, 13, 14) {real, imag} */,
  {32'hbf1c3e80, 32'hc1f79235} /* (5, 13, 13) {real, imag} */,
  {32'h41b6cede, 32'hc1359874} /* (5, 13, 12) {real, imag} */,
  {32'hc0cafa8a, 32'hc211c061} /* (5, 13, 11) {real, imag} */,
  {32'hbf3d6a70, 32'h416c9fb7} /* (5, 13, 10) {real, imag} */,
  {32'hc13260f4, 32'hc165c5c8} /* (5, 13, 9) {real, imag} */,
  {32'h41f520d3, 32'hc01aef48} /* (5, 13, 8) {real, imag} */,
  {32'h4021a6d9, 32'hc187ddb4} /* (5, 13, 7) {real, imag} */,
  {32'hc10ed68a, 32'hc08f1bdc} /* (5, 13, 6) {real, imag} */,
  {32'hc1308d3f, 32'h419f6728} /* (5, 13, 5) {real, imag} */,
  {32'h40e62800, 32'h40e86096} /* (5, 13, 4) {real, imag} */,
  {32'h4066dd42, 32'hc1e80358} /* (5, 13, 3) {real, imag} */,
  {32'hc2625672, 32'h401c6622} /* (5, 13, 2) {real, imag} */,
  {32'h40fbe70c, 32'hc1882a8a} /* (5, 13, 1) {real, imag} */,
  {32'hc16732c6, 32'hc206b5d6} /* (5, 13, 0) {real, imag} */,
  {32'h4222cc74, 32'hc20b4bff} /* (5, 12, 15) {real, imag} */,
  {32'h4147802a, 32'hc102ccc6} /* (5, 12, 14) {real, imag} */,
  {32'hc1307823, 32'hc20d0fca} /* (5, 12, 13) {real, imag} */,
  {32'hc21609e4, 32'hc1ba89bf} /* (5, 12, 12) {real, imag} */,
  {32'hc19b2de9, 32'h4178cfe5} /* (5, 12, 11) {real, imag} */,
  {32'h4148232d, 32'hc1902f34} /* (5, 12, 10) {real, imag} */,
  {32'h41659c19, 32'h413f34c6} /* (5, 12, 9) {real, imag} */,
  {32'h40c98fe0, 32'h410ec442} /* (5, 12, 8) {real, imag} */,
  {32'hc19c5b44, 32'h418f3e90} /* (5, 12, 7) {real, imag} */,
  {32'hc1d20b5a, 32'h4220478a} /* (5, 12, 6) {real, imag} */,
  {32'hc10f20d5, 32'h3ff34f70} /* (5, 12, 5) {real, imag} */,
  {32'hc202aa36, 32'h40a7c6e0} /* (5, 12, 4) {real, imag} */,
  {32'hc21647c2, 32'hc158224b} /* (5, 12, 3) {real, imag} */,
  {32'h413cfaa0, 32'h3fbe4008} /* (5, 12, 2) {real, imag} */,
  {32'hc16b2ee1, 32'hc0d4d1fc} /* (5, 12, 1) {real, imag} */,
  {32'h419e0982, 32'hc0f88e34} /* (5, 12, 0) {real, imag} */,
  {32'hc1075eda, 32'hc1e24dd6} /* (5, 11, 15) {real, imag} */,
  {32'h410abe63, 32'h41d7a2f3} /* (5, 11, 14) {real, imag} */,
  {32'h406eed34, 32'h421d5a64} /* (5, 11, 13) {real, imag} */,
  {32'hc24f64e8, 32'hc13f3cf4} /* (5, 11, 12) {real, imag} */,
  {32'h41e870f3, 32'hc13877a4} /* (5, 11, 11) {real, imag} */,
  {32'h40b55850, 32'hc23fe2d4} /* (5, 11, 10) {real, imag} */,
  {32'hc21fdea9, 32'hc09cf960} /* (5, 11, 9) {real, imag} */,
  {32'hc1846dd5, 32'h41813c4f} /* (5, 11, 8) {real, imag} */,
  {32'hc1934f3f, 32'hc225d922} /* (5, 11, 7) {real, imag} */,
  {32'h42227004, 32'hc168c7a7} /* (5, 11, 6) {real, imag} */,
  {32'hc2051c2c, 32'hc18acb53} /* (5, 11, 5) {real, imag} */,
  {32'hc1bc71b4, 32'hc1e98aae} /* (5, 11, 4) {real, imag} */,
  {32'hc17c474e, 32'h420827f5} /* (5, 11, 3) {real, imag} */,
  {32'h41a7450e, 32'h4183131d} /* (5, 11, 2) {real, imag} */,
  {32'h41c005c4, 32'h414a3772} /* (5, 11, 1) {real, imag} */,
  {32'hc032da70, 32'h418d3426} /* (5, 11, 0) {real, imag} */,
  {32'h42506117, 32'h40768d5c} /* (5, 10, 15) {real, imag} */,
  {32'h41875aef, 32'h41b379d5} /* (5, 10, 14) {real, imag} */,
  {32'h41916435, 32'h424c5d7e} /* (5, 10, 13) {real, imag} */,
  {32'hbff2f9a0, 32'hc28f24ee} /* (5, 10, 12) {real, imag} */,
  {32'hc1b22147, 32'hc146a9e1} /* (5, 10, 11) {real, imag} */,
  {32'h41b98ba2, 32'h41152b82} /* (5, 10, 10) {real, imag} */,
  {32'hc19db32f, 32'h41020222} /* (5, 10, 9) {real, imag} */,
  {32'hc09bf14c, 32'hc12e3c2c} /* (5, 10, 8) {real, imag} */,
  {32'h41f9cce8, 32'h3fa06e38} /* (5, 10, 7) {real, imag} */,
  {32'h4212351d, 32'hc1b29f07} /* (5, 10, 6) {real, imag} */,
  {32'h417ef340, 32'h41a59ede} /* (5, 10, 5) {real, imag} */,
  {32'h40931f84, 32'h422eb868} /* (5, 10, 4) {real, imag} */,
  {32'h40d4c387, 32'h41087bcc} /* (5, 10, 3) {real, imag} */,
  {32'h4122b868, 32'hbf3ed320} /* (5, 10, 2) {real, imag} */,
  {32'hc2377409, 32'h41237f02} /* (5, 10, 1) {real, imag} */,
  {32'hc132fb44, 32'hbfc0623c} /* (5, 10, 0) {real, imag} */,
  {32'h41ab1d12, 32'h41d49edf} /* (5, 9, 15) {real, imag} */,
  {32'h403d54b4, 32'hc1020956} /* (5, 9, 14) {real, imag} */,
  {32'hc213c41a, 32'h3e3efc40} /* (5, 9, 13) {real, imag} */,
  {32'hc154ce20, 32'hc18c1ff7} /* (5, 9, 12) {real, imag} */,
  {32'hc1c98e46, 32'h40ed6ea4} /* (5, 9, 11) {real, imag} */,
  {32'h410176b2, 32'h41c08130} /* (5, 9, 10) {real, imag} */,
  {32'hc0b0008e, 32'h403c0ba9} /* (5, 9, 9) {real, imag} */,
  {32'hc1c15a0e, 32'h419d1bef} /* (5, 9, 8) {real, imag} */,
  {32'h3f8a05b0, 32'h4180c3e8} /* (5, 9, 7) {real, imag} */,
  {32'h41c55ce0, 32'h4118349a} /* (5, 9, 6) {real, imag} */,
  {32'h415bf400, 32'h41a5ace8} /* (5, 9, 5) {real, imag} */,
  {32'h418084c6, 32'h3f2a8e60} /* (5, 9, 4) {real, imag} */,
  {32'hc0e22aa6, 32'hc11aac09} /* (5, 9, 3) {real, imag} */,
  {32'h41092afe, 32'h41a759a1} /* (5, 9, 2) {real, imag} */,
  {32'hc1689590, 32'hbfad28e8} /* (5, 9, 1) {real, imag} */,
  {32'h40931c70, 32'h401c2910} /* (5, 9, 0) {real, imag} */,
  {32'hbdde8ea0, 32'h421747d0} /* (5, 8, 15) {real, imag} */,
  {32'h411c05ce, 32'hc18c77c8} /* (5, 8, 14) {real, imag} */,
  {32'hbf659c38, 32'hc1630e33} /* (5, 8, 13) {real, imag} */,
  {32'h41e7b6a5, 32'hc0c68373} /* (5, 8, 12) {real, imag} */,
  {32'hc1dc2442, 32'h417d650c} /* (5, 8, 11) {real, imag} */,
  {32'hc06c696c, 32'hbfea0d38} /* (5, 8, 10) {real, imag} */,
  {32'h41b5e940, 32'hc18cf4cf} /* (5, 8, 9) {real, imag} */,
  {32'hc11addba, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h41b5e940, 32'h418cf4cf} /* (5, 8, 7) {real, imag} */,
  {32'hc06c696c, 32'h3fea0d38} /* (5, 8, 6) {real, imag} */,
  {32'hc1dc2442, 32'hc17d650c} /* (5, 8, 5) {real, imag} */,
  {32'h41e7b6a5, 32'h40c68373} /* (5, 8, 4) {real, imag} */,
  {32'hbf659c38, 32'h41630e33} /* (5, 8, 3) {real, imag} */,
  {32'h411c05ce, 32'h418c77c8} /* (5, 8, 2) {real, imag} */,
  {32'hbdde8ea0, 32'hc21747d0} /* (5, 8, 1) {real, imag} */,
  {32'h41a76bb3, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'hc1689590, 32'h3fad28e8} /* (5, 7, 15) {real, imag} */,
  {32'h41092afe, 32'hc1a759a1} /* (5, 7, 14) {real, imag} */,
  {32'hc0e22aa6, 32'h411aac09} /* (5, 7, 13) {real, imag} */,
  {32'h418084c6, 32'hbf2a8e60} /* (5, 7, 12) {real, imag} */,
  {32'h415bf400, 32'hc1a5ace8} /* (5, 7, 11) {real, imag} */,
  {32'h41c55ce0, 32'hc118349a} /* (5, 7, 10) {real, imag} */,
  {32'h3f8a05b0, 32'hc180c3e8} /* (5, 7, 9) {real, imag} */,
  {32'hc1c15a0e, 32'hc19d1bef} /* (5, 7, 8) {real, imag} */,
  {32'hc0b0008e, 32'hc03c0ba9} /* (5, 7, 7) {real, imag} */,
  {32'h410176b2, 32'hc1c08130} /* (5, 7, 6) {real, imag} */,
  {32'hc1c98e46, 32'hc0ed6ea4} /* (5, 7, 5) {real, imag} */,
  {32'hc154ce20, 32'h418c1ff7} /* (5, 7, 4) {real, imag} */,
  {32'hc213c41a, 32'hbe3efc40} /* (5, 7, 3) {real, imag} */,
  {32'h403d54b4, 32'h41020956} /* (5, 7, 2) {real, imag} */,
  {32'h41ab1d12, 32'hc1d49edf} /* (5, 7, 1) {real, imag} */,
  {32'h40931c70, 32'hc01c2910} /* (5, 7, 0) {real, imag} */,
  {32'hc2377409, 32'hc1237f02} /* (5, 6, 15) {real, imag} */,
  {32'h4122b868, 32'h3f3ed320} /* (5, 6, 14) {real, imag} */,
  {32'h40d4c387, 32'hc1087bcc} /* (5, 6, 13) {real, imag} */,
  {32'h40931f84, 32'hc22eb868} /* (5, 6, 12) {real, imag} */,
  {32'h417ef340, 32'hc1a59ede} /* (5, 6, 11) {real, imag} */,
  {32'h4212351d, 32'h41b29f07} /* (5, 6, 10) {real, imag} */,
  {32'h41f9cce8, 32'hbfa06e38} /* (5, 6, 9) {real, imag} */,
  {32'hc09bf14c, 32'h412e3c2c} /* (5, 6, 8) {real, imag} */,
  {32'hc19db32f, 32'hc1020222} /* (5, 6, 7) {real, imag} */,
  {32'h41b98ba2, 32'hc1152b82} /* (5, 6, 6) {real, imag} */,
  {32'hc1b22147, 32'h4146a9e1} /* (5, 6, 5) {real, imag} */,
  {32'hbff2f9a0, 32'h428f24ee} /* (5, 6, 4) {real, imag} */,
  {32'h41916435, 32'hc24c5d7e} /* (5, 6, 3) {real, imag} */,
  {32'h41875aef, 32'hc1b379d5} /* (5, 6, 2) {real, imag} */,
  {32'h42506117, 32'hc0768d5c} /* (5, 6, 1) {real, imag} */,
  {32'hc132fb44, 32'h3fc0623c} /* (5, 6, 0) {real, imag} */,
  {32'h41c005c4, 32'hc14a3772} /* (5, 5, 15) {real, imag} */,
  {32'h41a7450e, 32'hc183131d} /* (5, 5, 14) {real, imag} */,
  {32'hc17c474e, 32'hc20827f5} /* (5, 5, 13) {real, imag} */,
  {32'hc1bc71b4, 32'h41e98aae} /* (5, 5, 12) {real, imag} */,
  {32'hc2051c2c, 32'h418acb53} /* (5, 5, 11) {real, imag} */,
  {32'h42227004, 32'h4168c7a7} /* (5, 5, 10) {real, imag} */,
  {32'hc1934f3f, 32'h4225d922} /* (5, 5, 9) {real, imag} */,
  {32'hc1846dd5, 32'hc1813c4f} /* (5, 5, 8) {real, imag} */,
  {32'hc21fdea9, 32'h409cf960} /* (5, 5, 7) {real, imag} */,
  {32'h40b55850, 32'h423fe2d4} /* (5, 5, 6) {real, imag} */,
  {32'h41e870f3, 32'h413877a4} /* (5, 5, 5) {real, imag} */,
  {32'hc24f64e8, 32'h413f3cf4} /* (5, 5, 4) {real, imag} */,
  {32'h406eed34, 32'hc21d5a64} /* (5, 5, 3) {real, imag} */,
  {32'h410abe63, 32'hc1d7a2f3} /* (5, 5, 2) {real, imag} */,
  {32'hc1075eda, 32'h41e24dd6} /* (5, 5, 1) {real, imag} */,
  {32'hc032da70, 32'hc18d3426} /* (5, 5, 0) {real, imag} */,
  {32'hc16b2ee1, 32'h40d4d1fc} /* (5, 4, 15) {real, imag} */,
  {32'h413cfaa0, 32'hbfbe4008} /* (5, 4, 14) {real, imag} */,
  {32'hc21647c2, 32'h4158224b} /* (5, 4, 13) {real, imag} */,
  {32'hc202aa36, 32'hc0a7c6e0} /* (5, 4, 12) {real, imag} */,
  {32'hc10f20d5, 32'hbff34f70} /* (5, 4, 11) {real, imag} */,
  {32'hc1d20b5a, 32'hc220478a} /* (5, 4, 10) {real, imag} */,
  {32'hc19c5b44, 32'hc18f3e90} /* (5, 4, 9) {real, imag} */,
  {32'h40c98fe0, 32'hc10ec442} /* (5, 4, 8) {real, imag} */,
  {32'h41659c19, 32'hc13f34c6} /* (5, 4, 7) {real, imag} */,
  {32'h4148232d, 32'h41902f34} /* (5, 4, 6) {real, imag} */,
  {32'hc19b2de9, 32'hc178cfe5} /* (5, 4, 5) {real, imag} */,
  {32'hc21609e4, 32'h41ba89bf} /* (5, 4, 4) {real, imag} */,
  {32'hc1307823, 32'h420d0fca} /* (5, 4, 3) {real, imag} */,
  {32'h4147802a, 32'h4102ccc6} /* (5, 4, 2) {real, imag} */,
  {32'h4222cc74, 32'h420b4bff} /* (5, 4, 1) {real, imag} */,
  {32'h419e0982, 32'h40f88e34} /* (5, 4, 0) {real, imag} */,
  {32'h40fbe70c, 32'h41882a8a} /* (5, 3, 15) {real, imag} */,
  {32'hc2625672, 32'hc01c6622} /* (5, 3, 14) {real, imag} */,
  {32'h4066dd42, 32'h41e80358} /* (5, 3, 13) {real, imag} */,
  {32'h40e62800, 32'hc0e86096} /* (5, 3, 12) {real, imag} */,
  {32'hc1308d3f, 32'hc19f6728} /* (5, 3, 11) {real, imag} */,
  {32'hc10ed68a, 32'h408f1bdc} /* (5, 3, 10) {real, imag} */,
  {32'h4021a6d9, 32'h4187ddb4} /* (5, 3, 9) {real, imag} */,
  {32'h41f520d3, 32'h401aef48} /* (5, 3, 8) {real, imag} */,
  {32'hc13260f4, 32'h4165c5c8} /* (5, 3, 7) {real, imag} */,
  {32'hbf3d6a70, 32'hc16c9fb7} /* (5, 3, 6) {real, imag} */,
  {32'hc0cafa8a, 32'h4211c061} /* (5, 3, 5) {real, imag} */,
  {32'h41b6cede, 32'h41359874} /* (5, 3, 4) {real, imag} */,
  {32'hbf1c3e80, 32'h41f79235} /* (5, 3, 3) {real, imag} */,
  {32'hc101cc98, 32'h418487a2} /* (5, 3, 2) {real, imag} */,
  {32'hc1a6be2a, 32'hc1aafe58} /* (5, 3, 1) {real, imag} */,
  {32'hc16732c6, 32'h4206b5d6} /* (5, 3, 0) {real, imag} */,
  {32'hc143d1b6, 32'h41b3bc65} /* (5, 2, 15) {real, imag} */,
  {32'h421f82fb, 32'h42863a22} /* (5, 2, 14) {real, imag} */,
  {32'h4130e2cc, 32'hc17b8d66} /* (5, 2, 13) {real, imag} */,
  {32'h41ec94ba, 32'h421a598e} /* (5, 2, 12) {real, imag} */,
  {32'hc083e36c, 32'h4212e32b} /* (5, 2, 11) {real, imag} */,
  {32'hc17fa545, 32'hbfb1cec0} /* (5, 2, 10) {real, imag} */,
  {32'hc216dee2, 32'h3eb6bae0} /* (5, 2, 9) {real, imag} */,
  {32'h4121f3c4, 32'h41f4332a} /* (5, 2, 8) {real, imag} */,
  {32'h414a5014, 32'h40d6f3c0} /* (5, 2, 7) {real, imag} */,
  {32'hc0e335b6, 32'h41148e68} /* (5, 2, 6) {real, imag} */,
  {32'h41cbf47b, 32'h40fd86e9} /* (5, 2, 5) {real, imag} */,
  {32'h419fec4f, 32'hc1dd6637} /* (5, 2, 4) {real, imag} */,
  {32'hc1e6f256, 32'h41c76cde} /* (5, 2, 3) {real, imag} */,
  {32'hc0b5d1f4, 32'h41aa1f9d} /* (5, 2, 2) {real, imag} */,
  {32'hc02f0420, 32'hc22cb651} /* (5, 2, 1) {real, imag} */,
  {32'h428bf210, 32'hc256b62d} /* (5, 2, 0) {real, imag} */,
  {32'hc2d7a90c, 32'h41982198} /* (5, 1, 15) {real, imag} */,
  {32'hc295ba32, 32'h3f807370} /* (5, 1, 14) {real, imag} */,
  {32'hc21c6d87, 32'h41c26bfe} /* (5, 1, 13) {real, imag} */,
  {32'h4263f9b4, 32'h41bc92de} /* (5, 1, 12) {real, imag} */,
  {32'h40ae2c54, 32'h4119181f} /* (5, 1, 11) {real, imag} */,
  {32'h4141c261, 32'h41667592} /* (5, 1, 10) {real, imag} */,
  {32'h41cb79d9, 32'hc0a04773} /* (5, 1, 9) {real, imag} */,
  {32'hc00b0d5a, 32'h405593da} /* (5, 1, 8) {real, imag} */,
  {32'hc09e2a70, 32'h40c333e8} /* (5, 1, 7) {real, imag} */,
  {32'h41ba21df, 32'hc1d3d481} /* (5, 1, 6) {real, imag} */,
  {32'h4172dd3a, 32'h41c23111} /* (5, 1, 5) {real, imag} */,
  {32'hc02edfbc, 32'hc1684d0c} /* (5, 1, 4) {real, imag} */,
  {32'h40b45ec9, 32'hc225adf1} /* (5, 1, 3) {real, imag} */,
  {32'hc1e0fec4, 32'hc06b98a4} /* (5, 1, 2) {real, imag} */,
  {32'h42448106, 32'h42df6874} /* (5, 1, 1) {real, imag} */,
  {32'hc28b142b, 32'h41a307c0} /* (5, 1, 0) {real, imag} */,
  {32'hc2b83918, 32'h42b8b23c} /* (5, 0, 15) {real, imag} */,
  {32'h42067767, 32'hc2b9e0fc} /* (5, 0, 14) {real, imag} */,
  {32'h423235a9, 32'hc250e8c4} /* (5, 0, 13) {real, imag} */,
  {32'hc1cca129, 32'h4191d05c} /* (5, 0, 12) {real, imag} */,
  {32'hc11481fe, 32'h422a7a8b} /* (5, 0, 11) {real, imag} */,
  {32'h41d3bd4e, 32'hc08b4d76} /* (5, 0, 10) {real, imag} */,
  {32'h41899c3c, 32'h41135301} /* (5, 0, 9) {real, imag} */,
  {32'hc18c49c6, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'h41899c3c, 32'hc1135301} /* (5, 0, 7) {real, imag} */,
  {32'h41d3bd4e, 32'h408b4d76} /* (5, 0, 6) {real, imag} */,
  {32'hc11481fe, 32'hc22a7a8b} /* (5, 0, 5) {real, imag} */,
  {32'hc1cca129, 32'hc191d05c} /* (5, 0, 4) {real, imag} */,
  {32'h423235a9, 32'h4250e8c4} /* (5, 0, 3) {real, imag} */,
  {32'h42067767, 32'h42b9e0fc} /* (5, 0, 2) {real, imag} */,
  {32'hc2b83918, 32'hc2b8b23c} /* (5, 0, 1) {real, imag} */,
  {32'hc3a59416, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'h42974444, 32'hc2c6b285} /* (4, 15, 15) {real, imag} */,
  {32'hc2a39a71, 32'h42432b46} /* (4, 15, 14) {real, imag} */,
  {32'h41ac8845, 32'h42091ab1} /* (4, 15, 13) {real, imag} */,
  {32'h420dac70, 32'hc184c959} /* (4, 15, 12) {real, imag} */,
  {32'h41aa6f56, 32'hc114b6ec} /* (4, 15, 11) {real, imag} */,
  {32'hc18ac7b8, 32'hc0cbaea8} /* (4, 15, 10) {real, imag} */,
  {32'h40dfef5e, 32'h419db238} /* (4, 15, 9) {real, imag} */,
  {32'h410665f2, 32'h411c2665} /* (4, 15, 8) {real, imag} */,
  {32'hc1d17b11, 32'h415a6afc} /* (4, 15, 7) {real, imag} */,
  {32'h42288867, 32'hc14731f4} /* (4, 15, 6) {real, imag} */,
  {32'hc1ada05c, 32'hc11a3680} /* (4, 15, 5) {real, imag} */,
  {32'h40db553c, 32'hc1146f42} /* (4, 15, 4) {real, imag} */,
  {32'hc20d3c95, 32'hc1bd5ec0} /* (4, 15, 3) {real, imag} */,
  {32'hc1c91913, 32'h413c507c} /* (4, 15, 2) {real, imag} */,
  {32'hc2f26e6f, 32'hc2163df8} /* (4, 15, 1) {real, imag} */,
  {32'hc2304d46, 32'hc2bfdbd0} /* (4, 15, 0) {real, imag} */,
  {32'h4293959a, 32'hc09c30aa} /* (4, 14, 15) {real, imag} */,
  {32'h41fceb00, 32'hc20dfe74} /* (4, 14, 14) {real, imag} */,
  {32'hc1e25d75, 32'hc20375b0} /* (4, 14, 13) {real, imag} */,
  {32'hc21374bc, 32'h4132f536} /* (4, 14, 12) {real, imag} */,
  {32'hc142b586, 32'h41a52a6d} /* (4, 14, 11) {real, imag} */,
  {32'h41f6e2af, 32'hc0a13120} /* (4, 14, 10) {real, imag} */,
  {32'hc18380ba, 32'h413c6938} /* (4, 14, 9) {real, imag} */,
  {32'hc10b288a, 32'h405b6b72} /* (4, 14, 8) {real, imag} */,
  {32'h418b9ac3, 32'h418bf73c} /* (4, 14, 7) {real, imag} */,
  {32'hc1cb04cc, 32'h41fc35f5} /* (4, 14, 6) {real, imag} */,
  {32'h41237077, 32'hc182e734} /* (4, 14, 5) {real, imag} */,
  {32'h4080f9b4, 32'h4084fea2} /* (4, 14, 4) {real, imag} */,
  {32'hc10a28f8, 32'h420d7e8c} /* (4, 14, 3) {real, imag} */,
  {32'h41db1096, 32'hc0bc5812} /* (4, 14, 2) {real, imag} */,
  {32'hc1fa97f6, 32'h414d6028} /* (4, 14, 1) {real, imag} */,
  {32'h41205c4a, 32'h418503de} /* (4, 14, 0) {real, imag} */,
  {32'hc2088f47, 32'h41ca2f92} /* (4, 13, 15) {real, imag} */,
  {32'h417e4738, 32'hc112a660} /* (4, 13, 14) {real, imag} */,
  {32'hc0eafec6, 32'hc25b1cc9} /* (4, 13, 13) {real, imag} */,
  {32'hc20a21bc, 32'h412ab7f5} /* (4, 13, 12) {real, imag} */,
  {32'h416f3e63, 32'h40c6dc9e} /* (4, 13, 11) {real, imag} */,
  {32'h4166b97b, 32'hc1057168} /* (4, 13, 10) {real, imag} */,
  {32'hc1d009a8, 32'h3fc79380} /* (4, 13, 9) {real, imag} */,
  {32'h401d5ffe, 32'hc118d834} /* (4, 13, 8) {real, imag} */,
  {32'hc1030832, 32'h416b0d87} /* (4, 13, 7) {real, imag} */,
  {32'h40fec88a, 32'hc143e5c0} /* (4, 13, 6) {real, imag} */,
  {32'hc186a0a1, 32'hc1121b96} /* (4, 13, 5) {real, imag} */,
  {32'h40328f90, 32'hc1da33be} /* (4, 13, 4) {real, imag} */,
  {32'hc1b1cbb4, 32'h40680f9a} /* (4, 13, 3) {real, imag} */,
  {32'hc23b785e, 32'h41cd4c22} /* (4, 13, 2) {real, imag} */,
  {32'hc1a6eb18, 32'hc235601a} /* (4, 13, 1) {real, imag} */,
  {32'h420e6b0c, 32'hc15fbac7} /* (4, 13, 0) {real, imag} */,
  {32'hc1331f0b, 32'hc1057d5a} /* (4, 12, 15) {real, imag} */,
  {32'hc09e4e82, 32'h40adf31c} /* (4, 12, 14) {real, imag} */,
  {32'h3fafdf90, 32'hc20bc505} /* (4, 12, 13) {real, imag} */,
  {32'hc08b44a8, 32'h422e5d34} /* (4, 12, 12) {real, imag} */,
  {32'hc1d2d1f8, 32'hc13a3d21} /* (4, 12, 11) {real, imag} */,
  {32'h41062954, 32'h4100544b} /* (4, 12, 10) {real, imag} */,
  {32'hc15bb71d, 32'hc1ca16ba} /* (4, 12, 9) {real, imag} */,
  {32'hc14b53b0, 32'h40aa3f99} /* (4, 12, 8) {real, imag} */,
  {32'h4176fe7e, 32'hc25252cd} /* (4, 12, 7) {real, imag} */,
  {32'hc02bf52a, 32'h417aa447} /* (4, 12, 6) {real, imag} */,
  {32'h415a846d, 32'h412f3b37} /* (4, 12, 5) {real, imag} */,
  {32'hc2220fc5, 32'hc1ab4359} /* (4, 12, 4) {real, imag} */,
  {32'h41c81aac, 32'h412c818c} /* (4, 12, 3) {real, imag} */,
  {32'h3ff4d37a, 32'h412df00e} /* (4, 12, 2) {real, imag} */,
  {32'h41958b8f, 32'hc0104c18} /* (4, 12, 1) {real, imag} */,
  {32'h42000b33, 32'hbd97f1e0} /* (4, 12, 0) {real, imag} */,
  {32'hc1d7ee7c, 32'h3f7fde00} /* (4, 11, 15) {real, imag} */,
  {32'h41745960, 32'hc078422c} /* (4, 11, 14) {real, imag} */,
  {32'hc1afd56d, 32'hc17871cc} /* (4, 11, 13) {real, imag} */,
  {32'h41bf4bbc, 32'hc1df0f79} /* (4, 11, 12) {real, imag} */,
  {32'h410358c8, 32'hc0746970} /* (4, 11, 11) {real, imag} */,
  {32'h4189dc57, 32'hbe6c94d0} /* (4, 11, 10) {real, imag} */,
  {32'h4159f5ae, 32'h416572bd} /* (4, 11, 9) {real, imag} */,
  {32'h41b9cd9c, 32'h40fc8ce6} /* (4, 11, 8) {real, imag} */,
  {32'h415205ef, 32'h4144c81a} /* (4, 11, 7) {real, imag} */,
  {32'h40e1ad07, 32'hc0298d30} /* (4, 11, 6) {real, imag} */,
  {32'h3ecf74e0, 32'h40d96688} /* (4, 11, 5) {real, imag} */,
  {32'h4161320c, 32'h41991fbe} /* (4, 11, 4) {real, imag} */,
  {32'hc23b4550, 32'h42144ae6} /* (4, 11, 3) {real, imag} */,
  {32'h4183a851, 32'hc1921b13} /* (4, 11, 2) {real, imag} */,
  {32'hc172147e, 32'h41acfd99} /* (4, 11, 1) {real, imag} */,
  {32'hc1edaebc, 32'h417f5f3d} /* (4, 11, 0) {real, imag} */,
  {32'hc1a9cfb6, 32'h421975f1} /* (4, 10, 15) {real, imag} */,
  {32'h41a40886, 32'hc0b1a4c2} /* (4, 10, 14) {real, imag} */,
  {32'h419eb212, 32'h413c6e48} /* (4, 10, 13) {real, imag} */,
  {32'hc1279eb5, 32'hc227e85d} /* (4, 10, 12) {real, imag} */,
  {32'h4033100c, 32'h41830702} /* (4, 10, 11) {real, imag} */,
  {32'hc1e99ae6, 32'h4192d519} /* (4, 10, 10) {real, imag} */,
  {32'h41a8b4ec, 32'h4110ee9e} /* (4, 10, 9) {real, imag} */,
  {32'h417c71b8, 32'hc181dc55} /* (4, 10, 8) {real, imag} */,
  {32'hc1d679aa, 32'h419f9338} /* (4, 10, 7) {real, imag} */,
  {32'hc1d8a9f8, 32'h40522bbc} /* (4, 10, 6) {real, imag} */,
  {32'h41a49841, 32'h4161f79c} /* (4, 10, 5) {real, imag} */,
  {32'hbfb7d92c, 32'h419e9084} /* (4, 10, 4) {real, imag} */,
  {32'h4016b42c, 32'h3ee9e310} /* (4, 10, 3) {real, imag} */,
  {32'h41822f3a, 32'h423fc55a} /* (4, 10, 2) {real, imag} */,
  {32'h410064ad, 32'hc2037405} /* (4, 10, 1) {real, imag} */,
  {32'hbf09d0b0, 32'hc21e57f7} /* (4, 10, 0) {real, imag} */,
  {32'h4134d79e, 32'h410e1d7e} /* (4, 9, 15) {real, imag} */,
  {32'h417ca86c, 32'h40d0046c} /* (4, 9, 14) {real, imag} */,
  {32'hc139c772, 32'h4199e6c7} /* (4, 9, 13) {real, imag} */,
  {32'hbfbb5ae8, 32'h40e90790} /* (4, 9, 12) {real, imag} */,
  {32'hc02f0bd0, 32'h3f9556e4} /* (4, 9, 11) {real, imag} */,
  {32'hbfed26a0, 32'h418e702c} /* (4, 9, 10) {real, imag} */,
  {32'h41153333, 32'hbfc4743a} /* (4, 9, 9) {real, imag} */,
  {32'hc0a1b0ef, 32'hc0ea54f1} /* (4, 9, 8) {real, imag} */,
  {32'h410e7c85, 32'hc1705ef4} /* (4, 9, 7) {real, imag} */,
  {32'h41b054c2, 32'h41602a7a} /* (4, 9, 6) {real, imag} */,
  {32'hc0302be0, 32'hc188bb15} /* (4, 9, 5) {real, imag} */,
  {32'h414d926e, 32'hc081e45a} /* (4, 9, 4) {real, imag} */,
  {32'hc19de767, 32'hc1914f81} /* (4, 9, 3) {real, imag} */,
  {32'h415b382a, 32'hc14e3fee} /* (4, 9, 2) {real, imag} */,
  {32'hc1223d64, 32'hc160597a} /* (4, 9, 1) {real, imag} */,
  {32'hc15f83a0, 32'h4148392c} /* (4, 9, 0) {real, imag} */,
  {32'h4196effa, 32'hc0920642} /* (4, 8, 15) {real, imag} */,
  {32'h3fd6c548, 32'h404a0be4} /* (4, 8, 14) {real, imag} */,
  {32'h41f6f5fc, 32'hc10fc590} /* (4, 8, 13) {real, imag} */,
  {32'h3f946b00, 32'h41d38c48} /* (4, 8, 12) {real, imag} */,
  {32'hc149ad82, 32'h4132b8bc} /* (4, 8, 11) {real, imag} */,
  {32'h40f66cc6, 32'h416518dd} /* (4, 8, 10) {real, imag} */,
  {32'hc1fe7cee, 32'hc18ce0df} /* (4, 8, 9) {real, imag} */,
  {32'hc0946a30, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'hc1fe7cee, 32'h418ce0df} /* (4, 8, 7) {real, imag} */,
  {32'h40f66cc6, 32'hc16518dd} /* (4, 8, 6) {real, imag} */,
  {32'hc149ad82, 32'hc132b8bc} /* (4, 8, 5) {real, imag} */,
  {32'h3f946b00, 32'hc1d38c48} /* (4, 8, 4) {real, imag} */,
  {32'h41f6f5fc, 32'h410fc590} /* (4, 8, 3) {real, imag} */,
  {32'h3fd6c548, 32'hc04a0be4} /* (4, 8, 2) {real, imag} */,
  {32'h4196effa, 32'h40920642} /* (4, 8, 1) {real, imag} */,
  {32'hc213ade2, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hc1223d64, 32'h4160597a} /* (4, 7, 15) {real, imag} */,
  {32'h415b382a, 32'h414e3fee} /* (4, 7, 14) {real, imag} */,
  {32'hc19de767, 32'h41914f81} /* (4, 7, 13) {real, imag} */,
  {32'h414d926e, 32'h4081e45a} /* (4, 7, 12) {real, imag} */,
  {32'hc0302be0, 32'h4188bb15} /* (4, 7, 11) {real, imag} */,
  {32'h41b054c2, 32'hc1602a7a} /* (4, 7, 10) {real, imag} */,
  {32'h410e7c85, 32'h41705ef4} /* (4, 7, 9) {real, imag} */,
  {32'hc0a1b0ef, 32'h40ea54f1} /* (4, 7, 8) {real, imag} */,
  {32'h41153333, 32'h3fc4743a} /* (4, 7, 7) {real, imag} */,
  {32'hbfed26a0, 32'hc18e702c} /* (4, 7, 6) {real, imag} */,
  {32'hc02f0bd0, 32'hbf9556e4} /* (4, 7, 5) {real, imag} */,
  {32'hbfbb5ae8, 32'hc0e90790} /* (4, 7, 4) {real, imag} */,
  {32'hc139c772, 32'hc199e6c7} /* (4, 7, 3) {real, imag} */,
  {32'h417ca86c, 32'hc0d0046c} /* (4, 7, 2) {real, imag} */,
  {32'h4134d79e, 32'hc10e1d7e} /* (4, 7, 1) {real, imag} */,
  {32'hc15f83a0, 32'hc148392c} /* (4, 7, 0) {real, imag} */,
  {32'h410064ad, 32'h42037405} /* (4, 6, 15) {real, imag} */,
  {32'h41822f3a, 32'hc23fc55a} /* (4, 6, 14) {real, imag} */,
  {32'h4016b42c, 32'hbee9e310} /* (4, 6, 13) {real, imag} */,
  {32'hbfb7d92c, 32'hc19e9084} /* (4, 6, 12) {real, imag} */,
  {32'h41a49841, 32'hc161f79c} /* (4, 6, 11) {real, imag} */,
  {32'hc1d8a9f8, 32'hc0522bbc} /* (4, 6, 10) {real, imag} */,
  {32'hc1d679aa, 32'hc19f9338} /* (4, 6, 9) {real, imag} */,
  {32'h417c71b8, 32'h4181dc55} /* (4, 6, 8) {real, imag} */,
  {32'h41a8b4ec, 32'hc110ee9e} /* (4, 6, 7) {real, imag} */,
  {32'hc1e99ae6, 32'hc192d519} /* (4, 6, 6) {real, imag} */,
  {32'h4033100c, 32'hc1830702} /* (4, 6, 5) {real, imag} */,
  {32'hc1279eb5, 32'h4227e85d} /* (4, 6, 4) {real, imag} */,
  {32'h419eb212, 32'hc13c6e48} /* (4, 6, 3) {real, imag} */,
  {32'h41a40886, 32'h40b1a4c2} /* (4, 6, 2) {real, imag} */,
  {32'hc1a9cfb6, 32'hc21975f1} /* (4, 6, 1) {real, imag} */,
  {32'hbf09d0b0, 32'h421e57f7} /* (4, 6, 0) {real, imag} */,
  {32'hc172147e, 32'hc1acfd99} /* (4, 5, 15) {real, imag} */,
  {32'h4183a851, 32'h41921b13} /* (4, 5, 14) {real, imag} */,
  {32'hc23b4550, 32'hc2144ae6} /* (4, 5, 13) {real, imag} */,
  {32'h4161320c, 32'hc1991fbe} /* (4, 5, 12) {real, imag} */,
  {32'h3ecf74e0, 32'hc0d96688} /* (4, 5, 11) {real, imag} */,
  {32'h40e1ad07, 32'h40298d30} /* (4, 5, 10) {real, imag} */,
  {32'h415205ef, 32'hc144c81a} /* (4, 5, 9) {real, imag} */,
  {32'h41b9cd9c, 32'hc0fc8ce6} /* (4, 5, 8) {real, imag} */,
  {32'h4159f5ae, 32'hc16572bd} /* (4, 5, 7) {real, imag} */,
  {32'h4189dc57, 32'h3e6c94d0} /* (4, 5, 6) {real, imag} */,
  {32'h410358c8, 32'h40746970} /* (4, 5, 5) {real, imag} */,
  {32'h41bf4bbc, 32'h41df0f79} /* (4, 5, 4) {real, imag} */,
  {32'hc1afd56d, 32'h417871cc} /* (4, 5, 3) {real, imag} */,
  {32'h41745960, 32'h4078422c} /* (4, 5, 2) {real, imag} */,
  {32'hc1d7ee7c, 32'hbf7fde00} /* (4, 5, 1) {real, imag} */,
  {32'hc1edaebc, 32'hc17f5f3d} /* (4, 5, 0) {real, imag} */,
  {32'h41958b8f, 32'h40104c18} /* (4, 4, 15) {real, imag} */,
  {32'h3ff4d37a, 32'hc12df00e} /* (4, 4, 14) {real, imag} */,
  {32'h41c81aac, 32'hc12c818c} /* (4, 4, 13) {real, imag} */,
  {32'hc2220fc5, 32'h41ab4359} /* (4, 4, 12) {real, imag} */,
  {32'h415a846d, 32'hc12f3b37} /* (4, 4, 11) {real, imag} */,
  {32'hc02bf52a, 32'hc17aa447} /* (4, 4, 10) {real, imag} */,
  {32'h4176fe7e, 32'h425252cd} /* (4, 4, 9) {real, imag} */,
  {32'hc14b53b0, 32'hc0aa3f99} /* (4, 4, 8) {real, imag} */,
  {32'hc15bb71d, 32'h41ca16ba} /* (4, 4, 7) {real, imag} */,
  {32'h41062954, 32'hc100544b} /* (4, 4, 6) {real, imag} */,
  {32'hc1d2d1f8, 32'h413a3d21} /* (4, 4, 5) {real, imag} */,
  {32'hc08b44a8, 32'hc22e5d34} /* (4, 4, 4) {real, imag} */,
  {32'h3fafdf90, 32'h420bc505} /* (4, 4, 3) {real, imag} */,
  {32'hc09e4e82, 32'hc0adf31c} /* (4, 4, 2) {real, imag} */,
  {32'hc1331f0b, 32'h41057d5a} /* (4, 4, 1) {real, imag} */,
  {32'h42000b33, 32'h3d97f1e0} /* (4, 4, 0) {real, imag} */,
  {32'hc1a6eb18, 32'h4235601a} /* (4, 3, 15) {real, imag} */,
  {32'hc23b785e, 32'hc1cd4c22} /* (4, 3, 14) {real, imag} */,
  {32'hc1b1cbb4, 32'hc0680f9a} /* (4, 3, 13) {real, imag} */,
  {32'h40328f90, 32'h41da33be} /* (4, 3, 12) {real, imag} */,
  {32'hc186a0a1, 32'h41121b96} /* (4, 3, 11) {real, imag} */,
  {32'h40fec88a, 32'h4143e5c0} /* (4, 3, 10) {real, imag} */,
  {32'hc1030832, 32'hc16b0d87} /* (4, 3, 9) {real, imag} */,
  {32'h401d5ffe, 32'h4118d834} /* (4, 3, 8) {real, imag} */,
  {32'hc1d009a8, 32'hbfc79380} /* (4, 3, 7) {real, imag} */,
  {32'h4166b97b, 32'h41057168} /* (4, 3, 6) {real, imag} */,
  {32'h416f3e63, 32'hc0c6dc9e} /* (4, 3, 5) {real, imag} */,
  {32'hc20a21bc, 32'hc12ab7f5} /* (4, 3, 4) {real, imag} */,
  {32'hc0eafec6, 32'h425b1cc9} /* (4, 3, 3) {real, imag} */,
  {32'h417e4738, 32'h4112a660} /* (4, 3, 2) {real, imag} */,
  {32'hc2088f47, 32'hc1ca2f92} /* (4, 3, 1) {real, imag} */,
  {32'h420e6b0c, 32'h415fbac7} /* (4, 3, 0) {real, imag} */,
  {32'hc1fa97f6, 32'hc14d6028} /* (4, 2, 15) {real, imag} */,
  {32'h41db1096, 32'h40bc5812} /* (4, 2, 14) {real, imag} */,
  {32'hc10a28f8, 32'hc20d7e8c} /* (4, 2, 13) {real, imag} */,
  {32'h4080f9b4, 32'hc084fea2} /* (4, 2, 12) {real, imag} */,
  {32'h41237077, 32'h4182e734} /* (4, 2, 11) {real, imag} */,
  {32'hc1cb04cc, 32'hc1fc35f5} /* (4, 2, 10) {real, imag} */,
  {32'h418b9ac3, 32'hc18bf73c} /* (4, 2, 9) {real, imag} */,
  {32'hc10b288a, 32'hc05b6b72} /* (4, 2, 8) {real, imag} */,
  {32'hc18380ba, 32'hc13c6938} /* (4, 2, 7) {real, imag} */,
  {32'h41f6e2af, 32'h40a13120} /* (4, 2, 6) {real, imag} */,
  {32'hc142b586, 32'hc1a52a6d} /* (4, 2, 5) {real, imag} */,
  {32'hc21374bc, 32'hc132f536} /* (4, 2, 4) {real, imag} */,
  {32'hc1e25d75, 32'h420375b0} /* (4, 2, 3) {real, imag} */,
  {32'h41fceb00, 32'h420dfe74} /* (4, 2, 2) {real, imag} */,
  {32'h4293959a, 32'h409c30aa} /* (4, 2, 1) {real, imag} */,
  {32'h41205c4a, 32'hc18503de} /* (4, 2, 0) {real, imag} */,
  {32'hc2f26e6f, 32'h42163df8} /* (4, 1, 15) {real, imag} */,
  {32'hc1c91913, 32'hc13c507c} /* (4, 1, 14) {real, imag} */,
  {32'hc20d3c95, 32'h41bd5ec0} /* (4, 1, 13) {real, imag} */,
  {32'h40db553c, 32'h41146f42} /* (4, 1, 12) {real, imag} */,
  {32'hc1ada05c, 32'h411a3680} /* (4, 1, 11) {real, imag} */,
  {32'h42288867, 32'h414731f4} /* (4, 1, 10) {real, imag} */,
  {32'hc1d17b11, 32'hc15a6afc} /* (4, 1, 9) {real, imag} */,
  {32'h410665f2, 32'hc11c2665} /* (4, 1, 8) {real, imag} */,
  {32'h40dfef5e, 32'hc19db238} /* (4, 1, 7) {real, imag} */,
  {32'hc18ac7b8, 32'h40cbaea8} /* (4, 1, 6) {real, imag} */,
  {32'h41aa6f56, 32'h4114b6ec} /* (4, 1, 5) {real, imag} */,
  {32'h420dac70, 32'h4184c959} /* (4, 1, 4) {real, imag} */,
  {32'h41ac8845, 32'hc2091ab1} /* (4, 1, 3) {real, imag} */,
  {32'hc2a39a71, 32'hc2432b46} /* (4, 1, 2) {real, imag} */,
  {32'h42974444, 32'h42c6b285} /* (4, 1, 1) {real, imag} */,
  {32'hc2304d46, 32'h42bfdbd0} /* (4, 1, 0) {real, imag} */,
  {32'hc2ce49d4, 32'h42325a82} /* (4, 0, 15) {real, imag} */,
  {32'h410718be, 32'hc2c081d7} /* (4, 0, 14) {real, imag} */,
  {32'h4270dddf, 32'h41b80ef7} /* (4, 0, 13) {real, imag} */,
  {32'h41f48cc0, 32'h421a1448} /* (4, 0, 12) {real, imag} */,
  {32'h4216de66, 32'hc1dfd626} /* (4, 0, 11) {real, imag} */,
  {32'h4158d042, 32'hc108e516} /* (4, 0, 10) {real, imag} */,
  {32'h411c336d, 32'h41b1c1ec} /* (4, 0, 9) {real, imag} */,
  {32'hc10e5c08, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'h411c336d, 32'hc1b1c1ec} /* (4, 0, 7) {real, imag} */,
  {32'h4158d042, 32'h4108e516} /* (4, 0, 6) {real, imag} */,
  {32'h4216de66, 32'h41dfd626} /* (4, 0, 5) {real, imag} */,
  {32'h41f48cc0, 32'hc21a1448} /* (4, 0, 4) {real, imag} */,
  {32'h4270dddf, 32'hc1b80ef7} /* (4, 0, 3) {real, imag} */,
  {32'h410718be, 32'h42c081d7} /* (4, 0, 2) {real, imag} */,
  {32'hc2ce49d4, 32'hc2325a82} /* (4, 0, 1) {real, imag} */,
  {32'hc395039e, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'h425b8548, 32'hc26db8da} /* (3, 15, 15) {real, imag} */,
  {32'hc2831813, 32'h428a4ac6} /* (3, 15, 14) {real, imag} */,
  {32'hc1aae2b6, 32'h424f03a1} /* (3, 15, 13) {real, imag} */,
  {32'h400ddc20, 32'hc1c06a8c} /* (3, 15, 12) {real, imag} */,
  {32'hc22ac254, 32'h402cddba} /* (3, 15, 11) {real, imag} */,
  {32'h41db05c4, 32'hc1f3dfb1} /* (3, 15, 10) {real, imag} */,
  {32'h408b9357, 32'hc0dc558a} /* (3, 15, 9) {real, imag} */,
  {32'h41537aaf, 32'hc0475ad6} /* (3, 15, 8) {real, imag} */,
  {32'h419869d6, 32'h408c9073} /* (3, 15, 7) {real, imag} */,
  {32'h420c5dd3, 32'h41b45dfd} /* (3, 15, 6) {real, imag} */,
  {32'hc1903797, 32'h419782a6} /* (3, 15, 5) {real, imag} */,
  {32'h4019dbf0, 32'hc1d5772a} /* (3, 15, 4) {real, imag} */,
  {32'hc11d21cc, 32'hc27fdabf} /* (3, 15, 3) {real, imag} */,
  {32'hc1b136bc, 32'h417fa7aa} /* (3, 15, 2) {real, imag} */,
  {32'hc2919c40, 32'hc1e35ee4} /* (3, 15, 1) {real, imag} */,
  {32'hc211292f, 32'hc31910ac} /* (3, 15, 0) {real, imag} */,
  {32'h41a4b9cc, 32'h40fd3fa0} /* (3, 14, 15) {real, imag} */,
  {32'hc05d30ac, 32'hc242df0e} /* (3, 14, 14) {real, imag} */,
  {32'hc169f51f, 32'hc1836876} /* (3, 14, 13) {real, imag} */,
  {32'hc1f9ab28, 32'h41585ef4} /* (3, 14, 12) {real, imag} */,
  {32'hc040d100, 32'hc0762ad2} /* (3, 14, 11) {real, imag} */,
  {32'h406d66e3, 32'h4106a138} /* (3, 14, 10) {real, imag} */,
  {32'h413b2652, 32'h3f889b00} /* (3, 14, 9) {real, imag} */,
  {32'h4109ba58, 32'h4103bf6b} /* (3, 14, 8) {real, imag} */,
  {32'hc18662aa, 32'h41d31888} /* (3, 14, 7) {real, imag} */,
  {32'hc0a35fa2, 32'hc18a2d76} /* (3, 14, 6) {real, imag} */,
  {32'h415bfddd, 32'hbf72d130} /* (3, 14, 5) {real, imag} */,
  {32'hc18cbb3b, 32'hc135df69} /* (3, 14, 4) {real, imag} */,
  {32'hc107ea3a, 32'h41a52c53} /* (3, 14, 3) {real, imag} */,
  {32'h41797b27, 32'hbf98aac8} /* (3, 14, 2) {real, imag} */,
  {32'hc104bb54, 32'h421624bf} /* (3, 14, 1) {real, imag} */,
  {32'h41f336ec, 32'h418654ec} /* (3, 14, 0) {real, imag} */,
  {32'h41bf1400, 32'h4105e9ce} /* (3, 13, 15) {real, imag} */,
  {32'h40c90180, 32'h40d20a32} /* (3, 13, 14) {real, imag} */,
  {32'hc1bf969d, 32'hc125183c} /* (3, 13, 13) {real, imag} */,
  {32'hc1d4d092, 32'hc0f78e23} /* (3, 13, 12) {real, imag} */,
  {32'h42773205, 32'h42076eb3} /* (3, 13, 11) {real, imag} */,
  {32'hc1318531, 32'hc024dc2c} /* (3, 13, 10) {real, imag} */,
  {32'h408441a3, 32'hc16fa7f3} /* (3, 13, 9) {real, imag} */,
  {32'hc05970a2, 32'h3ff38750} /* (3, 13, 8) {real, imag} */,
  {32'hc0bde42a, 32'hbf1bc870} /* (3, 13, 7) {real, imag} */,
  {32'hc07606ee, 32'h41f5be6c} /* (3, 13, 6) {real, imag} */,
  {32'hc11c0294, 32'h416f545b} /* (3, 13, 5) {real, imag} */,
  {32'h41a22d7f, 32'hc2211802} /* (3, 13, 4) {real, imag} */,
  {32'h411246c4, 32'hc186d606} /* (3, 13, 3) {real, imag} */,
  {32'hc2309def, 32'hc20aae46} /* (3, 13, 2) {real, imag} */,
  {32'h3ea87240, 32'h406e50f0} /* (3, 13, 1) {real, imag} */,
  {32'h41282d0b, 32'hbfb747fc} /* (3, 13, 0) {real, imag} */,
  {32'hc03c72a0, 32'h41ab2758} /* (3, 12, 15) {real, imag} */,
  {32'hc0b1b3ea, 32'hc20f5f92} /* (3, 12, 14) {real, imag} */,
  {32'hc237388f, 32'h4034d1be} /* (3, 12, 13) {real, imag} */,
  {32'hc11d131b, 32'h42140e0e} /* (3, 12, 12) {real, imag} */,
  {32'hbe92eb00, 32'h422aee0a} /* (3, 12, 11) {real, imag} */,
  {32'h40e999d3, 32'hc120c322} /* (3, 12, 10) {real, imag} */,
  {32'hc17a4d68, 32'hc080a67e} /* (3, 12, 9) {real, imag} */,
  {32'h418e86c0, 32'h41a2ebad} /* (3, 12, 8) {real, imag} */,
  {32'hbf03e880, 32'hc0d1363c} /* (3, 12, 7) {real, imag} */,
  {32'h41eabfb0, 32'hc19c394a} /* (3, 12, 6) {real, imag} */,
  {32'hbfb47460, 32'h414496ac} /* (3, 12, 5) {real, imag} */,
  {32'hc1619769, 32'hc2017cc0} /* (3, 12, 4) {real, imag} */,
  {32'h412b8482, 32'h40973000} /* (3, 12, 3) {real, imag} */,
  {32'hc1fa45cb, 32'h4224245f} /* (3, 12, 2) {real, imag} */,
  {32'h41a833b6, 32'h41a0f8e1} /* (3, 12, 1) {real, imag} */,
  {32'h4215bf94, 32'h418e5986} /* (3, 12, 0) {real, imag} */,
  {32'h42264f9e, 32'h411e819a} /* (3, 11, 15) {real, imag} */,
  {32'hc227fc66, 32'h4099f906} /* (3, 11, 14) {real, imag} */,
  {32'h41b4fdf4, 32'hc0d2671c} /* (3, 11, 13) {real, imag} */,
  {32'h41bbeb43, 32'h41ebd640} /* (3, 11, 12) {real, imag} */,
  {32'hc0e09454, 32'hc10f4a96} /* (3, 11, 11) {real, imag} */,
  {32'hc17586bd, 32'h41585499} /* (3, 11, 10) {real, imag} */,
  {32'hbf287640, 32'h41717f45} /* (3, 11, 9) {real, imag} */,
  {32'hc18fae62, 32'h41abcde7} /* (3, 11, 8) {real, imag} */,
  {32'hc194955d, 32'hc157c7fe} /* (3, 11, 7) {real, imag} */,
  {32'hc23510a8, 32'h4233bc6e} /* (3, 11, 6) {real, imag} */,
  {32'hc0769612, 32'hc1b78a71} /* (3, 11, 5) {real, imag} */,
  {32'hc07fd5b7, 32'h41863a5e} /* (3, 11, 4) {real, imag} */,
  {32'hc1ba15f4, 32'hc18f5ea7} /* (3, 11, 3) {real, imag} */,
  {32'h4164a473, 32'hc251f1e6} /* (3, 11, 2) {real, imag} */,
  {32'h419c5217, 32'hc102bb44} /* (3, 11, 1) {real, imag} */,
  {32'hc117b79c, 32'h405af0d8} /* (3, 11, 0) {real, imag} */,
  {32'hc0bdb337, 32'h42034e44} /* (3, 10, 15) {real, imag} */,
  {32'h40cd4461, 32'hc189a982} /* (3, 10, 14) {real, imag} */,
  {32'h4112d43c, 32'hc11a5f50} /* (3, 10, 13) {real, imag} */,
  {32'h423127e1, 32'h421c5bcc} /* (3, 10, 12) {real, imag} */,
  {32'hc106db3c, 32'hc18b6dca} /* (3, 10, 11) {real, imag} */,
  {32'hc04ab020, 32'h42604461} /* (3, 10, 10) {real, imag} */,
  {32'hc093c072, 32'hc1a74f6c} /* (3, 10, 9) {real, imag} */,
  {32'hbff8ecae, 32'h403f5242} /* (3, 10, 8) {real, imag} */,
  {32'hc0e219c8, 32'h4134426c} /* (3, 10, 7) {real, imag} */,
  {32'hc11cef49, 32'hc14d6982} /* (3, 10, 6) {real, imag} */,
  {32'hc1136d37, 32'hc245a5c6} /* (3, 10, 5) {real, imag} */,
  {32'h4090e194, 32'hc0ab7388} /* (3, 10, 4) {real, imag} */,
  {32'h412f11b0, 32'h41708e38} /* (3, 10, 3) {real, imag} */,
  {32'hc10d57af, 32'hc19b2ce8} /* (3, 10, 2) {real, imag} */,
  {32'h419d313e, 32'hc09fde69} /* (3, 10, 1) {real, imag} */,
  {32'h41fc7e73, 32'h401fbb72} /* (3, 10, 0) {real, imag} */,
  {32'h40b80f59, 32'hc0b16e48} /* (3, 9, 15) {real, imag} */,
  {32'h4118cf7f, 32'h407ad7c8} /* (3, 9, 14) {real, imag} */,
  {32'hc1aed185, 32'hc1af9ab1} /* (3, 9, 13) {real, imag} */,
  {32'h3fce9c1c, 32'h41cc0131} /* (3, 9, 12) {real, imag} */,
  {32'h40fcee48, 32'h41e375e8} /* (3, 9, 11) {real, imag} */,
  {32'hc0b817c3, 32'hc1f01550} /* (3, 9, 10) {real, imag} */,
  {32'h417f14d4, 32'hc0bbebc8} /* (3, 9, 9) {real, imag} */,
  {32'h41afd654, 32'hc0be97be} /* (3, 9, 8) {real, imag} */,
  {32'h3fc3d968, 32'h41e78a2b} /* (3, 9, 7) {real, imag} */,
  {32'hc14b48e9, 32'hc1f63ba1} /* (3, 9, 6) {real, imag} */,
  {32'hc0766968, 32'hc212f496} /* (3, 9, 5) {real, imag} */,
  {32'h4150e7a8, 32'hc1f1d596} /* (3, 9, 4) {real, imag} */,
  {32'hc01fa348, 32'h41a3271e} /* (3, 9, 3) {real, imag} */,
  {32'hbf5189e0, 32'h416f27aa} /* (3, 9, 2) {real, imag} */,
  {32'h4170e9aa, 32'h416c22ba} /* (3, 9, 1) {real, imag} */,
  {32'h4002e2d8, 32'h40c657fa} /* (3, 9, 0) {real, imag} */,
  {32'hc0bb549a, 32'hc1ae3b7e} /* (3, 8, 15) {real, imag} */,
  {32'hc1a85148, 32'hc1839f35} /* (3, 8, 14) {real, imag} */,
  {32'h41d8f985, 32'hc00c63a0} /* (3, 8, 13) {real, imag} */,
  {32'h415088b6, 32'h40e46e8a} /* (3, 8, 12) {real, imag} */,
  {32'hbfc58a90, 32'h417d1d8e} /* (3, 8, 11) {real, imag} */,
  {32'h4022dcd0, 32'hc168c659} /* (3, 8, 10) {real, imag} */,
  {32'hc116b232, 32'h40e39a7e} /* (3, 8, 9) {real, imag} */,
  {32'h41e8a4e2, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'hc116b232, 32'hc0e39a7e} /* (3, 8, 7) {real, imag} */,
  {32'h4022dcd0, 32'h4168c659} /* (3, 8, 6) {real, imag} */,
  {32'hbfc58a90, 32'hc17d1d8e} /* (3, 8, 5) {real, imag} */,
  {32'h415088b6, 32'hc0e46e8a} /* (3, 8, 4) {real, imag} */,
  {32'h41d8f985, 32'h400c63a0} /* (3, 8, 3) {real, imag} */,
  {32'hc1a85148, 32'h41839f35} /* (3, 8, 2) {real, imag} */,
  {32'hc0bb549a, 32'h41ae3b7e} /* (3, 8, 1) {real, imag} */,
  {32'hc17e5f69, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'h4170e9aa, 32'hc16c22ba} /* (3, 7, 15) {real, imag} */,
  {32'hbf5189e0, 32'hc16f27aa} /* (3, 7, 14) {real, imag} */,
  {32'hc01fa348, 32'hc1a3271e} /* (3, 7, 13) {real, imag} */,
  {32'h4150e7a8, 32'h41f1d596} /* (3, 7, 12) {real, imag} */,
  {32'hc0766968, 32'h4212f496} /* (3, 7, 11) {real, imag} */,
  {32'hc14b48e9, 32'h41f63ba1} /* (3, 7, 10) {real, imag} */,
  {32'h3fc3d968, 32'hc1e78a2b} /* (3, 7, 9) {real, imag} */,
  {32'h41afd654, 32'h40be97be} /* (3, 7, 8) {real, imag} */,
  {32'h417f14d4, 32'h40bbebc8} /* (3, 7, 7) {real, imag} */,
  {32'hc0b817c3, 32'h41f01550} /* (3, 7, 6) {real, imag} */,
  {32'h40fcee48, 32'hc1e375e8} /* (3, 7, 5) {real, imag} */,
  {32'h3fce9c1c, 32'hc1cc0131} /* (3, 7, 4) {real, imag} */,
  {32'hc1aed185, 32'h41af9ab1} /* (3, 7, 3) {real, imag} */,
  {32'h4118cf7f, 32'hc07ad7c8} /* (3, 7, 2) {real, imag} */,
  {32'h40b80f59, 32'h40b16e48} /* (3, 7, 1) {real, imag} */,
  {32'h4002e2d8, 32'hc0c657fa} /* (3, 7, 0) {real, imag} */,
  {32'h419d313e, 32'h409fde69} /* (3, 6, 15) {real, imag} */,
  {32'hc10d57af, 32'h419b2ce8} /* (3, 6, 14) {real, imag} */,
  {32'h412f11b0, 32'hc1708e38} /* (3, 6, 13) {real, imag} */,
  {32'h4090e194, 32'h40ab7388} /* (3, 6, 12) {real, imag} */,
  {32'hc1136d37, 32'h4245a5c6} /* (3, 6, 11) {real, imag} */,
  {32'hc11cef49, 32'h414d6982} /* (3, 6, 10) {real, imag} */,
  {32'hc0e219c8, 32'hc134426c} /* (3, 6, 9) {real, imag} */,
  {32'hbff8ecae, 32'hc03f5242} /* (3, 6, 8) {real, imag} */,
  {32'hc093c072, 32'h41a74f6c} /* (3, 6, 7) {real, imag} */,
  {32'hc04ab020, 32'hc2604461} /* (3, 6, 6) {real, imag} */,
  {32'hc106db3c, 32'h418b6dca} /* (3, 6, 5) {real, imag} */,
  {32'h423127e1, 32'hc21c5bcc} /* (3, 6, 4) {real, imag} */,
  {32'h4112d43c, 32'h411a5f50} /* (3, 6, 3) {real, imag} */,
  {32'h40cd4461, 32'h4189a982} /* (3, 6, 2) {real, imag} */,
  {32'hc0bdb337, 32'hc2034e44} /* (3, 6, 1) {real, imag} */,
  {32'h41fc7e73, 32'hc01fbb72} /* (3, 6, 0) {real, imag} */,
  {32'h419c5217, 32'h4102bb44} /* (3, 5, 15) {real, imag} */,
  {32'h4164a473, 32'h4251f1e6} /* (3, 5, 14) {real, imag} */,
  {32'hc1ba15f4, 32'h418f5ea7} /* (3, 5, 13) {real, imag} */,
  {32'hc07fd5b7, 32'hc1863a5e} /* (3, 5, 12) {real, imag} */,
  {32'hc0769612, 32'h41b78a71} /* (3, 5, 11) {real, imag} */,
  {32'hc23510a8, 32'hc233bc6e} /* (3, 5, 10) {real, imag} */,
  {32'hc194955d, 32'h4157c7fe} /* (3, 5, 9) {real, imag} */,
  {32'hc18fae62, 32'hc1abcde7} /* (3, 5, 8) {real, imag} */,
  {32'hbf287640, 32'hc1717f45} /* (3, 5, 7) {real, imag} */,
  {32'hc17586bd, 32'hc1585499} /* (3, 5, 6) {real, imag} */,
  {32'hc0e09454, 32'h410f4a96} /* (3, 5, 5) {real, imag} */,
  {32'h41bbeb43, 32'hc1ebd640} /* (3, 5, 4) {real, imag} */,
  {32'h41b4fdf4, 32'h40d2671c} /* (3, 5, 3) {real, imag} */,
  {32'hc227fc66, 32'hc099f906} /* (3, 5, 2) {real, imag} */,
  {32'h42264f9e, 32'hc11e819a} /* (3, 5, 1) {real, imag} */,
  {32'hc117b79c, 32'hc05af0d8} /* (3, 5, 0) {real, imag} */,
  {32'h41a833b6, 32'hc1a0f8e1} /* (3, 4, 15) {real, imag} */,
  {32'hc1fa45cb, 32'hc224245f} /* (3, 4, 14) {real, imag} */,
  {32'h412b8482, 32'hc0973000} /* (3, 4, 13) {real, imag} */,
  {32'hc1619769, 32'h42017cc0} /* (3, 4, 12) {real, imag} */,
  {32'hbfb47460, 32'hc14496ac} /* (3, 4, 11) {real, imag} */,
  {32'h41eabfb0, 32'h419c394a} /* (3, 4, 10) {real, imag} */,
  {32'hbf03e880, 32'h40d1363c} /* (3, 4, 9) {real, imag} */,
  {32'h418e86c0, 32'hc1a2ebad} /* (3, 4, 8) {real, imag} */,
  {32'hc17a4d68, 32'h4080a67e} /* (3, 4, 7) {real, imag} */,
  {32'h40e999d3, 32'h4120c322} /* (3, 4, 6) {real, imag} */,
  {32'hbe92eb00, 32'hc22aee0a} /* (3, 4, 5) {real, imag} */,
  {32'hc11d131b, 32'hc2140e0e} /* (3, 4, 4) {real, imag} */,
  {32'hc237388f, 32'hc034d1be} /* (3, 4, 3) {real, imag} */,
  {32'hc0b1b3ea, 32'h420f5f92} /* (3, 4, 2) {real, imag} */,
  {32'hc03c72a0, 32'hc1ab2758} /* (3, 4, 1) {real, imag} */,
  {32'h4215bf94, 32'hc18e5986} /* (3, 4, 0) {real, imag} */,
  {32'h3ea87240, 32'hc06e50f0} /* (3, 3, 15) {real, imag} */,
  {32'hc2309def, 32'h420aae46} /* (3, 3, 14) {real, imag} */,
  {32'h411246c4, 32'h4186d606} /* (3, 3, 13) {real, imag} */,
  {32'h41a22d7f, 32'h42211802} /* (3, 3, 12) {real, imag} */,
  {32'hc11c0294, 32'hc16f545b} /* (3, 3, 11) {real, imag} */,
  {32'hc07606ee, 32'hc1f5be6c} /* (3, 3, 10) {real, imag} */,
  {32'hc0bde42a, 32'h3f1bc870} /* (3, 3, 9) {real, imag} */,
  {32'hc05970a2, 32'hbff38750} /* (3, 3, 8) {real, imag} */,
  {32'h408441a3, 32'h416fa7f3} /* (3, 3, 7) {real, imag} */,
  {32'hc1318531, 32'h4024dc2c} /* (3, 3, 6) {real, imag} */,
  {32'h42773205, 32'hc2076eb3} /* (3, 3, 5) {real, imag} */,
  {32'hc1d4d092, 32'h40f78e23} /* (3, 3, 4) {real, imag} */,
  {32'hc1bf969d, 32'h4125183c} /* (3, 3, 3) {real, imag} */,
  {32'h40c90180, 32'hc0d20a32} /* (3, 3, 2) {real, imag} */,
  {32'h41bf1400, 32'hc105e9ce} /* (3, 3, 1) {real, imag} */,
  {32'h41282d0b, 32'h3fb747fc} /* (3, 3, 0) {real, imag} */,
  {32'hc104bb54, 32'hc21624bf} /* (3, 2, 15) {real, imag} */,
  {32'h41797b27, 32'h3f98aac8} /* (3, 2, 14) {real, imag} */,
  {32'hc107ea3a, 32'hc1a52c53} /* (3, 2, 13) {real, imag} */,
  {32'hc18cbb3b, 32'h4135df69} /* (3, 2, 12) {real, imag} */,
  {32'h415bfddd, 32'h3f72d130} /* (3, 2, 11) {real, imag} */,
  {32'hc0a35fa2, 32'h418a2d76} /* (3, 2, 10) {real, imag} */,
  {32'hc18662aa, 32'hc1d31888} /* (3, 2, 9) {real, imag} */,
  {32'h4109ba58, 32'hc103bf6b} /* (3, 2, 8) {real, imag} */,
  {32'h413b2652, 32'hbf889b00} /* (3, 2, 7) {real, imag} */,
  {32'h406d66e3, 32'hc106a138} /* (3, 2, 6) {real, imag} */,
  {32'hc040d100, 32'h40762ad2} /* (3, 2, 5) {real, imag} */,
  {32'hc1f9ab28, 32'hc1585ef4} /* (3, 2, 4) {real, imag} */,
  {32'hc169f51f, 32'h41836876} /* (3, 2, 3) {real, imag} */,
  {32'hc05d30ac, 32'h4242df0e} /* (3, 2, 2) {real, imag} */,
  {32'h41a4b9cc, 32'hc0fd3fa0} /* (3, 2, 1) {real, imag} */,
  {32'h41f336ec, 32'hc18654ec} /* (3, 2, 0) {real, imag} */,
  {32'hc2919c40, 32'h41e35ee4} /* (3, 1, 15) {real, imag} */,
  {32'hc1b136bc, 32'hc17fa7aa} /* (3, 1, 14) {real, imag} */,
  {32'hc11d21cc, 32'h427fdabf} /* (3, 1, 13) {real, imag} */,
  {32'h4019dbf0, 32'h41d5772a} /* (3, 1, 12) {real, imag} */,
  {32'hc1903797, 32'hc19782a6} /* (3, 1, 11) {real, imag} */,
  {32'h420c5dd3, 32'hc1b45dfd} /* (3, 1, 10) {real, imag} */,
  {32'h419869d6, 32'hc08c9073} /* (3, 1, 9) {real, imag} */,
  {32'h41537aaf, 32'h40475ad6} /* (3, 1, 8) {real, imag} */,
  {32'h408b9357, 32'h40dc558a} /* (3, 1, 7) {real, imag} */,
  {32'h41db05c4, 32'h41f3dfb1} /* (3, 1, 6) {real, imag} */,
  {32'hc22ac254, 32'hc02cddba} /* (3, 1, 5) {real, imag} */,
  {32'h400ddc20, 32'h41c06a8c} /* (3, 1, 4) {real, imag} */,
  {32'hc1aae2b6, 32'hc24f03a1} /* (3, 1, 3) {real, imag} */,
  {32'hc2831813, 32'hc28a4ac6} /* (3, 1, 2) {real, imag} */,
  {32'h425b8548, 32'h426db8da} /* (3, 1, 1) {real, imag} */,
  {32'hc211292f, 32'h431910ac} /* (3, 1, 0) {real, imag} */,
  {32'hc2b196b3, 32'hc26b01d8} /* (3, 0, 15) {real, imag} */,
  {32'hc1763149, 32'hc19bbea8} /* (3, 0, 14) {real, imag} */,
  {32'h42443d78, 32'h41b6cb6e} /* (3, 0, 13) {real, imag} */,
  {32'h424f49c2, 32'h40fb9218} /* (3, 0, 12) {real, imag} */,
  {32'h40b467dd, 32'hc1e9f4ac} /* (3, 0, 11) {real, imag} */,
  {32'h41bdb71a, 32'hc0d70667} /* (3, 0, 10) {real, imag} */,
  {32'hc1c8a79d, 32'hbe1ad340} /* (3, 0, 9) {real, imag} */,
  {32'hc05a95dc, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'hc1c8a79d, 32'h3e1ad340} /* (3, 0, 7) {real, imag} */,
  {32'h41bdb71a, 32'h40d70667} /* (3, 0, 6) {real, imag} */,
  {32'h40b467dd, 32'h41e9f4ac} /* (3, 0, 5) {real, imag} */,
  {32'h424f49c2, 32'hc0fb9218} /* (3, 0, 4) {real, imag} */,
  {32'h42443d78, 32'hc1b6cb6e} /* (3, 0, 3) {real, imag} */,
  {32'hc1763149, 32'h419bbea8} /* (3, 0, 2) {real, imag} */,
  {32'hc2b196b3, 32'h426b01d8} /* (3, 0, 1) {real, imag} */,
  {32'hc3663dc2, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc10a34dc, 32'hc129ce5c} /* (2, 15, 15) {real, imag} */,
  {32'hc28b34d2, 32'h421f0a7b} /* (2, 15, 14) {real, imag} */,
  {32'hc0e0e0dc, 32'h41d69af8} /* (2, 15, 13) {real, imag} */,
  {32'hc1681882, 32'hc041a1d8} /* (2, 15, 12) {real, imag} */,
  {32'h3fcdac18, 32'h4121c573} /* (2, 15, 11) {real, imag} */,
  {32'hc1a0b94a, 32'hc0ab075f} /* (2, 15, 10) {real, imag} */,
  {32'h40333a18, 32'hc0ef1108} /* (2, 15, 9) {real, imag} */,
  {32'h40a53031, 32'hc06838a4} /* (2, 15, 8) {real, imag} */,
  {32'hc0b60a3d, 32'hc1660a96} /* (2, 15, 7) {real, imag} */,
  {32'h4082ef7f, 32'h4085f648} /* (2, 15, 6) {real, imag} */,
  {32'h41857457, 32'h41fa935a} /* (2, 15, 5) {real, imag} */,
  {32'hc103e1d9, 32'h4107ba31} /* (2, 15, 4) {real, imag} */,
  {32'h4223cda7, 32'hc2635e55} /* (2, 15, 3) {real, imag} */,
  {32'h4277586a, 32'hc14c0328} /* (2, 15, 2) {real, imag} */,
  {32'hc2f30a72, 32'hc1fdd204} /* (2, 15, 1) {real, imag} */,
  {32'hc2deb010, 32'hc2b19c74} /* (2, 15, 0) {real, imag} */,
  {32'hc11e94a9, 32'hc00dd368} /* (2, 14, 15) {real, imag} */,
  {32'hc1e4a961, 32'hc2813e8b} /* (2, 14, 14) {real, imag} */,
  {32'hc112dc17, 32'hc00f0038} /* (2, 14, 13) {real, imag} */,
  {32'hc21d2655, 32'hc287ee98} /* (2, 14, 12) {real, imag} */,
  {32'h41722523, 32'h40302a52} /* (2, 14, 11) {real, imag} */,
  {32'hc1ae27c4, 32'h4202a039} /* (2, 14, 10) {real, imag} */,
  {32'h42198c38, 32'h3f99b6d6} /* (2, 14, 9) {real, imag} */,
  {32'hc0d0dc84, 32'h3fdbd320} /* (2, 14, 8) {real, imag} */,
  {32'h41dbb729, 32'h41a3104a} /* (2, 14, 7) {real, imag} */,
  {32'hc0fc080a, 32'hc15dfe3e} /* (2, 14, 6) {real, imag} */,
  {32'h414b3fc2, 32'h40c3aedc} /* (2, 14, 5) {real, imag} */,
  {32'hc1a1d2ae, 32'hc080f16e} /* (2, 14, 4) {real, imag} */,
  {32'hc16b0fd1, 32'h41d29616} /* (2, 14, 3) {real, imag} */,
  {32'hc091dac4, 32'hc1a5c427} /* (2, 14, 2) {real, imag} */,
  {32'hc1978b14, 32'h41d04a74} /* (2, 14, 1) {real, imag} */,
  {32'h428841cf, 32'h42431cd6} /* (2, 14, 0) {real, imag} */,
  {32'h40b4c232, 32'hc108fd54} /* (2, 13, 15) {real, imag} */,
  {32'h41e6077c, 32'h4103c6ea} /* (2, 13, 14) {real, imag} */,
  {32'hbf855498, 32'h41f58ca3} /* (2, 13, 13) {real, imag} */,
  {32'h41072a7a, 32'h42857162} /* (2, 13, 12) {real, imag} */,
  {32'h4135b10d, 32'hc1304f18} /* (2, 13, 11) {real, imag} */,
  {32'hc2103256, 32'h40541c54} /* (2, 13, 10) {real, imag} */,
  {32'h40df93a9, 32'hbfa55fd8} /* (2, 13, 9) {real, imag} */,
  {32'h40890039, 32'hc0aa6652} /* (2, 13, 8) {real, imag} */,
  {32'hc1441048, 32'h41ce46e4} /* (2, 13, 7) {real, imag} */,
  {32'hc1add1d4, 32'hc030e340} /* (2, 13, 6) {real, imag} */,
  {32'hc1a43208, 32'h420a7c25} /* (2, 13, 5) {real, imag} */,
  {32'hc08da028, 32'h40a4621d} /* (2, 13, 4) {real, imag} */,
  {32'h41e23e02, 32'hc1c2aee0} /* (2, 13, 3) {real, imag} */,
  {32'hc22b3226, 32'hc20f4ade} /* (2, 13, 2) {real, imag} */,
  {32'hbfa1a7d8, 32'h4185abd6} /* (2, 13, 1) {real, imag} */,
  {32'hc20200f0, 32'hc1038cea} /* (2, 13, 0) {real, imag} */,
  {32'hc237feb6, 32'h41104fc8} /* (2, 12, 15) {real, imag} */,
  {32'h40590c62, 32'h41b4b3eb} /* (2, 12, 14) {real, imag} */,
  {32'hc2029338, 32'h41c737c7} /* (2, 12, 13) {real, imag} */,
  {32'h40537cb0, 32'h408d1864} /* (2, 12, 12) {real, imag} */,
  {32'h40b80982, 32'h41a68757} /* (2, 12, 11) {real, imag} */,
  {32'hc1370a14, 32'hc20ffcd8} /* (2, 12, 10) {real, imag} */,
  {32'hc140c7ce, 32'hc119df88} /* (2, 12, 9) {real, imag} */,
  {32'hc1e18cff, 32'hc12f7eb1} /* (2, 12, 8) {real, imag} */,
  {32'h41c4b940, 32'h400360fb} /* (2, 12, 7) {real, imag} */,
  {32'h40dbbfab, 32'hc1c1b5af} /* (2, 12, 6) {real, imag} */,
  {32'h40af1ec0, 32'h3fcb4698} /* (2, 12, 5) {real, imag} */,
  {32'hc1786948, 32'hc1a8808c} /* (2, 12, 4) {real, imag} */,
  {32'hc18210d7, 32'h42350b94} /* (2, 12, 3) {real, imag} */,
  {32'hc0a3906e, 32'hc11a3dcc} /* (2, 12, 2) {real, imag} */,
  {32'h40ca55bb, 32'hc1a00976} /* (2, 12, 1) {real, imag} */,
  {32'h422fe5c6, 32'hbf8a7e54} /* (2, 12, 0) {real, imag} */,
  {32'h41dbc67f, 32'h4206fc35} /* (2, 11, 15) {real, imag} */,
  {32'hc19604b0, 32'h41d63ac8} /* (2, 11, 14) {real, imag} */,
  {32'h4208a5ab, 32'h41e7e298} /* (2, 11, 13) {real, imag} */,
  {32'h41e35790, 32'hc09ae253} /* (2, 11, 12) {real, imag} */,
  {32'h4192cb0b, 32'hc1f0972c} /* (2, 11, 11) {real, imag} */,
  {32'hc0ee530e, 32'h418e98ea} /* (2, 11, 10) {real, imag} */,
  {32'h40ce873c, 32'hbe532c80} /* (2, 11, 9) {real, imag} */,
  {32'h413bc0c1, 32'h407234ec} /* (2, 11, 8) {real, imag} */,
  {32'hc2149203, 32'h4150bfda} /* (2, 11, 7) {real, imag} */,
  {32'h41565374, 32'h421e4b1f} /* (2, 11, 6) {real, imag} */,
  {32'h41344436, 32'h41abd908} /* (2, 11, 5) {real, imag} */,
  {32'hc119bff2, 32'hc0f1eaec} /* (2, 11, 4) {real, imag} */,
  {32'h41e8e76a, 32'hc10f31d2} /* (2, 11, 3) {real, imag} */,
  {32'hc11a6bfd, 32'hc09c24d8} /* (2, 11, 2) {real, imag} */,
  {32'h3f791900, 32'h3f1f39c0} /* (2, 11, 1) {real, imag} */,
  {32'hc00a0b10, 32'hc2020b28} /* (2, 11, 0) {real, imag} */,
  {32'h41a78ca3, 32'hc0957222} /* (2, 10, 15) {real, imag} */,
  {32'hc1b3e9bf, 32'hc09be4b6} /* (2, 10, 14) {real, imag} */,
  {32'hbf68f780, 32'hc1948880} /* (2, 10, 13) {real, imag} */,
  {32'hc12b7c66, 32'hc1a00c92} /* (2, 10, 12) {real, imag} */,
  {32'h419264e0, 32'h40b6b70c} /* (2, 10, 11) {real, imag} */,
  {32'h40cb8365, 32'hbf46f0c0} /* (2, 10, 10) {real, imag} */,
  {32'hc1156d3c, 32'h407c0f84} /* (2, 10, 9) {real, imag} */,
  {32'h41e79d5e, 32'hc14bd3af} /* (2, 10, 8) {real, imag} */,
  {32'h4189bd9a, 32'h409b1710} /* (2, 10, 7) {real, imag} */,
  {32'hc11bfa10, 32'h415e7b01} /* (2, 10, 6) {real, imag} */,
  {32'hc1bd91ea, 32'h41f1e386} /* (2, 10, 5) {real, imag} */,
  {32'h41e4445b, 32'h4100a214} /* (2, 10, 4) {real, imag} */,
  {32'hc1bbad5e, 32'hc19bc4c8} /* (2, 10, 3) {real, imag} */,
  {32'hbf539b18, 32'hc1fc85bb} /* (2, 10, 2) {real, imag} */,
  {32'h42030981, 32'hbf5f14f0} /* (2, 10, 1) {real, imag} */,
  {32'h3f6720c0, 32'h41e8c41c} /* (2, 10, 0) {real, imag} */,
  {32'h405ade22, 32'h3f95570c} /* (2, 9, 15) {real, imag} */,
  {32'hc11da962, 32'h41500098} /* (2, 9, 14) {real, imag} */,
  {32'hc1a6f211, 32'h41c0a9d9} /* (2, 9, 13) {real, imag} */,
  {32'h40839c12, 32'hc162fd53} /* (2, 9, 12) {real, imag} */,
  {32'hc165ac59, 32'h4014ed68} /* (2, 9, 11) {real, imag} */,
  {32'h41f202b5, 32'hc18a569e} /* (2, 9, 10) {real, imag} */,
  {32'h412ab316, 32'h41ab539f} /* (2, 9, 9) {real, imag} */,
  {32'hc154a76d, 32'h41be564a} /* (2, 9, 8) {real, imag} */,
  {32'hc1c61424, 32'hc0b53882} /* (2, 9, 7) {real, imag} */,
  {32'h41907cf1, 32'hc1454987} /* (2, 9, 6) {real, imag} */,
  {32'hc0216db0, 32'h4050092a} /* (2, 9, 5) {real, imag} */,
  {32'h4212737b, 32'hc18339f1} /* (2, 9, 4) {real, imag} */,
  {32'hc1df3238, 32'h41127bf4} /* (2, 9, 3) {real, imag} */,
  {32'h413f7165, 32'hc11ffcf6} /* (2, 9, 2) {real, imag} */,
  {32'h419a78fe, 32'hc0f15370} /* (2, 9, 1) {real, imag} */,
  {32'h41c70c52, 32'hc1233362} /* (2, 9, 0) {real, imag} */,
  {32'hc007fd9e, 32'h40d8bd4d} /* (2, 8, 15) {real, imag} */,
  {32'h4077a901, 32'hc1ccee31} /* (2, 8, 14) {real, imag} */,
  {32'h41174b53, 32'hc0af0bc2} /* (2, 8, 13) {real, imag} */,
  {32'hc1e3fcbd, 32'hc1ab559f} /* (2, 8, 12) {real, imag} */,
  {32'hc11c3914, 32'hc22b7b75} /* (2, 8, 11) {real, imag} */,
  {32'hc1b0c94a, 32'h41be2c06} /* (2, 8, 10) {real, imag} */,
  {32'hc0aebd0c, 32'h4207cfb6} /* (2, 8, 9) {real, imag} */,
  {32'h41afe364, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'hc0aebd0c, 32'hc207cfb6} /* (2, 8, 7) {real, imag} */,
  {32'hc1b0c94a, 32'hc1be2c06} /* (2, 8, 6) {real, imag} */,
  {32'hc11c3914, 32'h422b7b75} /* (2, 8, 5) {real, imag} */,
  {32'hc1e3fcbd, 32'h41ab559f} /* (2, 8, 4) {real, imag} */,
  {32'h41174b53, 32'h40af0bc2} /* (2, 8, 3) {real, imag} */,
  {32'h4077a901, 32'h41ccee31} /* (2, 8, 2) {real, imag} */,
  {32'hc007fd9e, 32'hc0d8bd4d} /* (2, 8, 1) {real, imag} */,
  {32'h414454d0, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'h419a78fe, 32'h40f15370} /* (2, 7, 15) {real, imag} */,
  {32'h413f7165, 32'h411ffcf6} /* (2, 7, 14) {real, imag} */,
  {32'hc1df3238, 32'hc1127bf4} /* (2, 7, 13) {real, imag} */,
  {32'h4212737b, 32'h418339f1} /* (2, 7, 12) {real, imag} */,
  {32'hc0216db0, 32'hc050092a} /* (2, 7, 11) {real, imag} */,
  {32'h41907cf1, 32'h41454987} /* (2, 7, 10) {real, imag} */,
  {32'hc1c61424, 32'h40b53882} /* (2, 7, 9) {real, imag} */,
  {32'hc154a76d, 32'hc1be564a} /* (2, 7, 8) {real, imag} */,
  {32'h412ab316, 32'hc1ab539f} /* (2, 7, 7) {real, imag} */,
  {32'h41f202b5, 32'h418a569e} /* (2, 7, 6) {real, imag} */,
  {32'hc165ac59, 32'hc014ed68} /* (2, 7, 5) {real, imag} */,
  {32'h40839c12, 32'h4162fd53} /* (2, 7, 4) {real, imag} */,
  {32'hc1a6f211, 32'hc1c0a9d9} /* (2, 7, 3) {real, imag} */,
  {32'hc11da962, 32'hc1500098} /* (2, 7, 2) {real, imag} */,
  {32'h405ade22, 32'hbf95570c} /* (2, 7, 1) {real, imag} */,
  {32'h41c70c52, 32'h41233362} /* (2, 7, 0) {real, imag} */,
  {32'h42030981, 32'h3f5f14f0} /* (2, 6, 15) {real, imag} */,
  {32'hbf539b18, 32'h41fc85bb} /* (2, 6, 14) {real, imag} */,
  {32'hc1bbad5e, 32'h419bc4c8} /* (2, 6, 13) {real, imag} */,
  {32'h41e4445b, 32'hc100a214} /* (2, 6, 12) {real, imag} */,
  {32'hc1bd91ea, 32'hc1f1e386} /* (2, 6, 11) {real, imag} */,
  {32'hc11bfa10, 32'hc15e7b01} /* (2, 6, 10) {real, imag} */,
  {32'h4189bd9a, 32'hc09b1710} /* (2, 6, 9) {real, imag} */,
  {32'h41e79d5e, 32'h414bd3af} /* (2, 6, 8) {real, imag} */,
  {32'hc1156d3c, 32'hc07c0f84} /* (2, 6, 7) {real, imag} */,
  {32'h40cb8365, 32'h3f46f0c0} /* (2, 6, 6) {real, imag} */,
  {32'h419264e0, 32'hc0b6b70c} /* (2, 6, 5) {real, imag} */,
  {32'hc12b7c66, 32'h41a00c92} /* (2, 6, 4) {real, imag} */,
  {32'hbf68f780, 32'h41948880} /* (2, 6, 3) {real, imag} */,
  {32'hc1b3e9bf, 32'h409be4b6} /* (2, 6, 2) {real, imag} */,
  {32'h41a78ca3, 32'h40957222} /* (2, 6, 1) {real, imag} */,
  {32'h3f6720c0, 32'hc1e8c41c} /* (2, 6, 0) {real, imag} */,
  {32'h3f791900, 32'hbf1f39c0} /* (2, 5, 15) {real, imag} */,
  {32'hc11a6bfd, 32'h409c24d8} /* (2, 5, 14) {real, imag} */,
  {32'h41e8e76a, 32'h410f31d2} /* (2, 5, 13) {real, imag} */,
  {32'hc119bff2, 32'h40f1eaec} /* (2, 5, 12) {real, imag} */,
  {32'h41344436, 32'hc1abd908} /* (2, 5, 11) {real, imag} */,
  {32'h41565374, 32'hc21e4b1f} /* (2, 5, 10) {real, imag} */,
  {32'hc2149203, 32'hc150bfda} /* (2, 5, 9) {real, imag} */,
  {32'h413bc0c1, 32'hc07234ec} /* (2, 5, 8) {real, imag} */,
  {32'h40ce873c, 32'h3e532c80} /* (2, 5, 7) {real, imag} */,
  {32'hc0ee530e, 32'hc18e98ea} /* (2, 5, 6) {real, imag} */,
  {32'h4192cb0b, 32'h41f0972c} /* (2, 5, 5) {real, imag} */,
  {32'h41e35790, 32'h409ae253} /* (2, 5, 4) {real, imag} */,
  {32'h4208a5ab, 32'hc1e7e298} /* (2, 5, 3) {real, imag} */,
  {32'hc19604b0, 32'hc1d63ac8} /* (2, 5, 2) {real, imag} */,
  {32'h41dbc67f, 32'hc206fc35} /* (2, 5, 1) {real, imag} */,
  {32'hc00a0b10, 32'h42020b28} /* (2, 5, 0) {real, imag} */,
  {32'h40ca55bb, 32'h41a00976} /* (2, 4, 15) {real, imag} */,
  {32'hc0a3906e, 32'h411a3dcc} /* (2, 4, 14) {real, imag} */,
  {32'hc18210d7, 32'hc2350b94} /* (2, 4, 13) {real, imag} */,
  {32'hc1786948, 32'h41a8808c} /* (2, 4, 12) {real, imag} */,
  {32'h40af1ec0, 32'hbfcb4698} /* (2, 4, 11) {real, imag} */,
  {32'h40dbbfab, 32'h41c1b5af} /* (2, 4, 10) {real, imag} */,
  {32'h41c4b940, 32'hc00360fb} /* (2, 4, 9) {real, imag} */,
  {32'hc1e18cff, 32'h412f7eb1} /* (2, 4, 8) {real, imag} */,
  {32'hc140c7ce, 32'h4119df88} /* (2, 4, 7) {real, imag} */,
  {32'hc1370a14, 32'h420ffcd8} /* (2, 4, 6) {real, imag} */,
  {32'h40b80982, 32'hc1a68757} /* (2, 4, 5) {real, imag} */,
  {32'h40537cb0, 32'hc08d1864} /* (2, 4, 4) {real, imag} */,
  {32'hc2029338, 32'hc1c737c7} /* (2, 4, 3) {real, imag} */,
  {32'h40590c62, 32'hc1b4b3eb} /* (2, 4, 2) {real, imag} */,
  {32'hc237feb6, 32'hc1104fc8} /* (2, 4, 1) {real, imag} */,
  {32'h422fe5c6, 32'h3f8a7e54} /* (2, 4, 0) {real, imag} */,
  {32'hbfa1a7d8, 32'hc185abd6} /* (2, 3, 15) {real, imag} */,
  {32'hc22b3226, 32'h420f4ade} /* (2, 3, 14) {real, imag} */,
  {32'h41e23e02, 32'h41c2aee0} /* (2, 3, 13) {real, imag} */,
  {32'hc08da028, 32'hc0a4621d} /* (2, 3, 12) {real, imag} */,
  {32'hc1a43208, 32'hc20a7c25} /* (2, 3, 11) {real, imag} */,
  {32'hc1add1d4, 32'h4030e340} /* (2, 3, 10) {real, imag} */,
  {32'hc1441048, 32'hc1ce46e4} /* (2, 3, 9) {real, imag} */,
  {32'h40890039, 32'h40aa6652} /* (2, 3, 8) {real, imag} */,
  {32'h40df93a9, 32'h3fa55fd8} /* (2, 3, 7) {real, imag} */,
  {32'hc2103256, 32'hc0541c54} /* (2, 3, 6) {real, imag} */,
  {32'h4135b10d, 32'h41304f18} /* (2, 3, 5) {real, imag} */,
  {32'h41072a7a, 32'hc2857162} /* (2, 3, 4) {real, imag} */,
  {32'hbf855498, 32'hc1f58ca3} /* (2, 3, 3) {real, imag} */,
  {32'h41e6077c, 32'hc103c6ea} /* (2, 3, 2) {real, imag} */,
  {32'h40b4c232, 32'h4108fd54} /* (2, 3, 1) {real, imag} */,
  {32'hc20200f0, 32'h41038cea} /* (2, 3, 0) {real, imag} */,
  {32'hc1978b14, 32'hc1d04a74} /* (2, 2, 15) {real, imag} */,
  {32'hc091dac4, 32'h41a5c427} /* (2, 2, 14) {real, imag} */,
  {32'hc16b0fd1, 32'hc1d29616} /* (2, 2, 13) {real, imag} */,
  {32'hc1a1d2ae, 32'h4080f16e} /* (2, 2, 12) {real, imag} */,
  {32'h414b3fc2, 32'hc0c3aedc} /* (2, 2, 11) {real, imag} */,
  {32'hc0fc080a, 32'h415dfe3e} /* (2, 2, 10) {real, imag} */,
  {32'h41dbb729, 32'hc1a3104a} /* (2, 2, 9) {real, imag} */,
  {32'hc0d0dc84, 32'hbfdbd320} /* (2, 2, 8) {real, imag} */,
  {32'h42198c38, 32'hbf99b6d6} /* (2, 2, 7) {real, imag} */,
  {32'hc1ae27c4, 32'hc202a039} /* (2, 2, 6) {real, imag} */,
  {32'h41722523, 32'hc0302a52} /* (2, 2, 5) {real, imag} */,
  {32'hc21d2655, 32'h4287ee98} /* (2, 2, 4) {real, imag} */,
  {32'hc112dc17, 32'h400f0038} /* (2, 2, 3) {real, imag} */,
  {32'hc1e4a961, 32'h42813e8b} /* (2, 2, 2) {real, imag} */,
  {32'hc11e94a9, 32'h400dd368} /* (2, 2, 1) {real, imag} */,
  {32'h428841cf, 32'hc2431cd6} /* (2, 2, 0) {real, imag} */,
  {32'hc2f30a72, 32'h41fdd204} /* (2, 1, 15) {real, imag} */,
  {32'h4277586a, 32'h414c0328} /* (2, 1, 14) {real, imag} */,
  {32'h4223cda7, 32'h42635e55} /* (2, 1, 13) {real, imag} */,
  {32'hc103e1d9, 32'hc107ba31} /* (2, 1, 12) {real, imag} */,
  {32'h41857457, 32'hc1fa935a} /* (2, 1, 11) {real, imag} */,
  {32'h4082ef7f, 32'hc085f648} /* (2, 1, 10) {real, imag} */,
  {32'hc0b60a3d, 32'h41660a96} /* (2, 1, 9) {real, imag} */,
  {32'h40a53031, 32'h406838a4} /* (2, 1, 8) {real, imag} */,
  {32'h40333a18, 32'h40ef1108} /* (2, 1, 7) {real, imag} */,
  {32'hc1a0b94a, 32'h40ab075f} /* (2, 1, 6) {real, imag} */,
  {32'h3fcdac18, 32'hc121c573} /* (2, 1, 5) {real, imag} */,
  {32'hc1681882, 32'h4041a1d8} /* (2, 1, 4) {real, imag} */,
  {32'hc0e0e0dc, 32'hc1d69af8} /* (2, 1, 3) {real, imag} */,
  {32'hc28b34d2, 32'hc21f0a7b} /* (2, 1, 2) {real, imag} */,
  {32'hc10a34dc, 32'h4129ce5c} /* (2, 1, 1) {real, imag} */,
  {32'hc2deb010, 32'h42b19c74} /* (2, 1, 0) {real, imag} */,
  {32'hc1b7f2d0, 32'hc311faa5} /* (2, 0, 15) {real, imag} */,
  {32'h40f65024, 32'hc217157f} /* (2, 0, 14) {real, imag} */,
  {32'h41fdd9bf, 32'h4208115c} /* (2, 0, 13) {real, imag} */,
  {32'h42374ed9, 32'hc13c851a} /* (2, 0, 12) {real, imag} */,
  {32'h418ade70, 32'h420506b7} /* (2, 0, 11) {real, imag} */,
  {32'h3f4b9300, 32'h4035b784} /* (2, 0, 10) {real, imag} */,
  {32'hc0eb1267, 32'hbfe20e20} /* (2, 0, 9) {real, imag} */,
  {32'hc1bfa82f, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'hc0eb1267, 32'h3fe20e20} /* (2, 0, 7) {real, imag} */,
  {32'h3f4b9300, 32'hc035b784} /* (2, 0, 6) {real, imag} */,
  {32'h418ade70, 32'hc20506b7} /* (2, 0, 5) {real, imag} */,
  {32'h42374ed9, 32'h413c851a} /* (2, 0, 4) {real, imag} */,
  {32'h41fdd9bf, 32'hc208115c} /* (2, 0, 3) {real, imag} */,
  {32'h40f65024, 32'h4217157f} /* (2, 0, 2) {real, imag} */,
  {32'hc1b7f2d0, 32'h4311faa5} /* (2, 0, 1) {real, imag} */,
  {32'hc29cdeb1, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc2729f75, 32'hc193a1c0} /* (1, 15, 15) {real, imag} */,
  {32'hc253d6e2, 32'h3fb7d670} /* (1, 15, 14) {real, imag} */,
  {32'hc1b89010, 32'h419a0c5f} /* (1, 15, 13) {real, imag} */,
  {32'h40d03162, 32'h413775d3} /* (1, 15, 12) {real, imag} */,
  {32'hc25f40ae, 32'h40e572ab} /* (1, 15, 11) {real, imag} */,
  {32'h41c666ec, 32'h41cb2d66} /* (1, 15, 10) {real, imag} */,
  {32'hc0378640, 32'h4100a2be} /* (1, 15, 9) {real, imag} */,
  {32'hc0bfd506, 32'h40a3c9a8} /* (1, 15, 8) {real, imag} */,
  {32'hc1c87e6b, 32'h4246da04} /* (1, 15, 7) {real, imag} */,
  {32'hc0246506, 32'hc0b34f52} /* (1, 15, 6) {real, imag} */,
  {32'h41ac2fd3, 32'h41e0c1b4} /* (1, 15, 5) {real, imag} */,
  {32'hc2274fce, 32'h419d2324} /* (1, 15, 4) {real, imag} */,
  {32'h4244732c, 32'hc20cfabe} /* (1, 15, 3) {real, imag} */,
  {32'h41f526aa, 32'h4227c624} /* (1, 15, 2) {real, imag} */,
  {32'hc2d34768, 32'hc0e5f238} /* (1, 15, 1) {real, imag} */,
  {32'hc2fa6a7f, 32'hc29c4211} /* (1, 15, 0) {real, imag} */,
  {32'h414c6744, 32'hc1189737} /* (1, 14, 15) {real, imag} */,
  {32'h413514ef, 32'hc25b046d} /* (1, 14, 14) {real, imag} */,
  {32'h421054f2, 32'hc23225da} /* (1, 14, 13) {real, imag} */,
  {32'hc113ea48, 32'hc1c3b7c0} /* (1, 14, 12) {real, imag} */,
  {32'h41119717, 32'hc14d7d1f} /* (1, 14, 11) {real, imag} */,
  {32'hc181e3b6, 32'hc175d83a} /* (1, 14, 10) {real, imag} */,
  {32'hc0b7a7ff, 32'h41a2dfe7} /* (1, 14, 9) {real, imag} */,
  {32'hc0f2c1c4, 32'hc10b3f4d} /* (1, 14, 8) {real, imag} */,
  {32'h4126ae00, 32'hc183199d} /* (1, 14, 7) {real, imag} */,
  {32'hc18f8462, 32'h4148173e} /* (1, 14, 6) {real, imag} */,
  {32'hc235065b, 32'hc0a5deac} /* (1, 14, 5) {real, imag} */,
  {32'h4110e681, 32'hc0ae6d6c} /* (1, 14, 4) {real, imag} */,
  {32'h40a682a4, 32'hc0c153d0} /* (1, 14, 3) {real, imag} */,
  {32'hc0075950, 32'h40831320} /* (1, 14, 2) {real, imag} */,
  {32'hc26170ee, 32'hc251a3b8} /* (1, 14, 1) {real, imag} */,
  {32'h41cace17, 32'h423c4bd4} /* (1, 14, 0) {real, imag} */,
  {32'hc14cfc17, 32'h412712c6} /* (1, 13, 15) {real, imag} */,
  {32'hc0ead5a4, 32'hc1fcd2b6} /* (1, 13, 14) {real, imag} */,
  {32'hc09ff6d9, 32'h4207321e} /* (1, 13, 13) {real, imag} */,
  {32'hbfc6cd38, 32'h428d51bd} /* (1, 13, 12) {real, imag} */,
  {32'hc083bfaa, 32'hbfd630c0} /* (1, 13, 11) {real, imag} */,
  {32'h40f52b4a, 32'h4198a854} /* (1, 13, 10) {real, imag} */,
  {32'hc24bb973, 32'h415d4ac4} /* (1, 13, 9) {real, imag} */,
  {32'hc012a874, 32'hc0ad201e} /* (1, 13, 8) {real, imag} */,
  {32'hc183431c, 32'h40f561d0} /* (1, 13, 7) {real, imag} */,
  {32'hbfaf9c64, 32'h410c3fde} /* (1, 13, 6) {real, imag} */,
  {32'hc1147b9c, 32'h40fc0314} /* (1, 13, 5) {real, imag} */,
  {32'h41c68ae8, 32'h418e8aae} /* (1, 13, 4) {real, imag} */,
  {32'h40b87788, 32'hc1810501} /* (1, 13, 3) {real, imag} */,
  {32'hc127c630, 32'h405ea578} /* (1, 13, 2) {real, imag} */,
  {32'h41587dda, 32'h42155c11} /* (1, 13, 1) {real, imag} */,
  {32'h3f80697c, 32'hc1f82c2a} /* (1, 13, 0) {real, imag} */,
  {32'h40fa1bf7, 32'h41cfcaeb} /* (1, 12, 15) {real, imag} */,
  {32'hc1cb4b7f, 32'h41bfbdbb} /* (1, 12, 14) {real, imag} */,
  {32'hc1cb445b, 32'h425370e0} /* (1, 12, 13) {real, imag} */,
  {32'hbfafe2c8, 32'h41f108d8} /* (1, 12, 12) {real, imag} */,
  {32'h418cc7ac, 32'hc197b78a} /* (1, 12, 11) {real, imag} */,
  {32'hc0470b7e, 32'hc1d1583c} /* (1, 12, 10) {real, imag} */,
  {32'hc1495788, 32'hc0bd6260} /* (1, 12, 9) {real, imag} */,
  {32'hc0972b39, 32'hc0c88e9d} /* (1, 12, 8) {real, imag} */,
  {32'h418697c0, 32'hc1d10eaf} /* (1, 12, 7) {real, imag} */,
  {32'hbf3cc8a0, 32'h422b2a60} /* (1, 12, 6) {real, imag} */,
  {32'hc1a7666e, 32'hc0c53f0d} /* (1, 12, 5) {real, imag} */,
  {32'hc192f67b, 32'hbfe46aec} /* (1, 12, 4) {real, imag} */,
  {32'h3fca6000, 32'h41ae6dc0} /* (1, 12, 3) {real, imag} */,
  {32'hc1ad66b6, 32'hc214735c} /* (1, 12, 2) {real, imag} */,
  {32'h42c92624, 32'hc261aa6f} /* (1, 12, 1) {real, imag} */,
  {32'hc16dca2a, 32'h4205c508} /* (1, 12, 0) {real, imag} */,
  {32'hc08e368c, 32'hc2124cfa} /* (1, 11, 15) {real, imag} */,
  {32'h4223ef08, 32'h3e8e33f0} /* (1, 11, 14) {real, imag} */,
  {32'hc20ccd02, 32'hc0df0a4e} /* (1, 11, 13) {real, imag} */,
  {32'hc1e58a12, 32'hc13947ac} /* (1, 11, 12) {real, imag} */,
  {32'hc11ff478, 32'hc1822f6e} /* (1, 11, 11) {real, imag} */,
  {32'h404e539e, 32'h41e322ae} /* (1, 11, 10) {real, imag} */,
  {32'h410fa710, 32'hc0dc9782} /* (1, 11, 9) {real, imag} */,
  {32'h40c49fc8, 32'h3ebba490} /* (1, 11, 8) {real, imag} */,
  {32'h41e0e9c0, 32'hc1497742} /* (1, 11, 7) {real, imag} */,
  {32'hc0bdf697, 32'hc1654c3d} /* (1, 11, 6) {real, imag} */,
  {32'hc002b5c2, 32'hc0fae564} /* (1, 11, 5) {real, imag} */,
  {32'h419274f7, 32'h41aab85c} /* (1, 11, 4) {real, imag} */,
  {32'h40f7c851, 32'h40b17a84} /* (1, 11, 3) {real, imag} */,
  {32'h414a5559, 32'hc08dd52c} /* (1, 11, 2) {real, imag} */,
  {32'h41c40eb9, 32'h4181e45c} /* (1, 11, 1) {real, imag} */,
  {32'hc1b16d8b, 32'h41577b44} /* (1, 11, 0) {real, imag} */,
  {32'hbf92e5ee, 32'hc1c98dca} /* (1, 10, 15) {real, imag} */,
  {32'h41129206, 32'hc1e2c9e8} /* (1, 10, 14) {real, imag} */,
  {32'hc0558c90, 32'hc0895de3} /* (1, 10, 13) {real, imag} */,
  {32'hc21587db, 32'h403ce22c} /* (1, 10, 12) {real, imag} */,
  {32'hc1fe877a, 32'h409a5b5d} /* (1, 10, 11) {real, imag} */,
  {32'hc17fd956, 32'hbf47eed8} /* (1, 10, 10) {real, imag} */,
  {32'h418c9b2b, 32'hc1c03324} /* (1, 10, 9) {real, imag} */,
  {32'h411987e0, 32'hc1857ff9} /* (1, 10, 8) {real, imag} */,
  {32'hc0985640, 32'h40062b62} /* (1, 10, 7) {real, imag} */,
  {32'hc10cf926, 32'hc2846cbe} /* (1, 10, 6) {real, imag} */,
  {32'h40e2bb9e, 32'h41e6f015} /* (1, 10, 5) {real, imag} */,
  {32'h41cc7108, 32'h41756044} /* (1, 10, 4) {real, imag} */,
  {32'hbfb19a4c, 32'h4221373c} /* (1, 10, 3) {real, imag} */,
  {32'hc13cd022, 32'h41c49840} /* (1, 10, 2) {real, imag} */,
  {32'hc1b391fc, 32'h419752c6} /* (1, 10, 1) {real, imag} */,
  {32'h4193160e, 32'h40a4d301} /* (1, 10, 0) {real, imag} */,
  {32'h41b229dc, 32'h41fdd1d8} /* (1, 9, 15) {real, imag} */,
  {32'hc1bdf7ee, 32'hc008af30} /* (1, 9, 14) {real, imag} */,
  {32'h40fa32fe, 32'hc1006d90} /* (1, 9, 13) {real, imag} */,
  {32'h40a7cb65, 32'hc0dfd3cb} /* (1, 9, 12) {real, imag} */,
  {32'h41cb9893, 32'hc13c9979} /* (1, 9, 11) {real, imag} */,
  {32'hc1a97bb4, 32'hbf3ff140} /* (1, 9, 10) {real, imag} */,
  {32'h417ee88c, 32'hc19f2b42} /* (1, 9, 9) {real, imag} */,
  {32'h3fe08b66, 32'hc06801af} /* (1, 9, 8) {real, imag} */,
  {32'h4087330c, 32'hc0ea2e96} /* (1, 9, 7) {real, imag} */,
  {32'h4151bb6e, 32'h3ead6b10} /* (1, 9, 6) {real, imag} */,
  {32'hc186fe2d, 32'hc1ebbc64} /* (1, 9, 5) {real, imag} */,
  {32'hc1175890, 32'hc128e3c6} /* (1, 9, 4) {real, imag} */,
  {32'h416294a4, 32'hc217e74c} /* (1, 9, 3) {real, imag} */,
  {32'h417f4804, 32'h414a7a6e} /* (1, 9, 2) {real, imag} */,
  {32'h4042ff58, 32'h4122a9b2} /* (1, 9, 1) {real, imag} */,
  {32'h3fab8250, 32'hc1457686} /* (1, 9, 0) {real, imag} */,
  {32'hc116e038, 32'h3fc1f118} /* (1, 8, 15) {real, imag} */,
  {32'hc1549f48, 32'hc0312757} /* (1, 8, 14) {real, imag} */,
  {32'hc1462ff0, 32'hc1880548} /* (1, 8, 13) {real, imag} */,
  {32'hc1ae419e, 32'hc0a953ea} /* (1, 8, 12) {real, imag} */,
  {32'h41277e4a, 32'h40c8b5a2} /* (1, 8, 11) {real, imag} */,
  {32'hc15ee1c1, 32'h40df4f48} /* (1, 8, 10) {real, imag} */,
  {32'h414e2232, 32'hc189d4bb} /* (1, 8, 9) {real, imag} */,
  {32'h3f9141c6, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'h414e2232, 32'h4189d4bb} /* (1, 8, 7) {real, imag} */,
  {32'hc15ee1c1, 32'hc0df4f48} /* (1, 8, 6) {real, imag} */,
  {32'h41277e4a, 32'hc0c8b5a2} /* (1, 8, 5) {real, imag} */,
  {32'hc1ae419e, 32'h40a953ea} /* (1, 8, 4) {real, imag} */,
  {32'hc1462ff0, 32'h41880548} /* (1, 8, 3) {real, imag} */,
  {32'hc1549f48, 32'h40312757} /* (1, 8, 2) {real, imag} */,
  {32'hc116e038, 32'hbfc1f118} /* (1, 8, 1) {real, imag} */,
  {32'hc1dc1fcc, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'h4042ff58, 32'hc122a9b2} /* (1, 7, 15) {real, imag} */,
  {32'h417f4804, 32'hc14a7a6e} /* (1, 7, 14) {real, imag} */,
  {32'h416294a4, 32'h4217e74c} /* (1, 7, 13) {real, imag} */,
  {32'hc1175890, 32'h4128e3c6} /* (1, 7, 12) {real, imag} */,
  {32'hc186fe2d, 32'h41ebbc64} /* (1, 7, 11) {real, imag} */,
  {32'h4151bb6e, 32'hbead6b10} /* (1, 7, 10) {real, imag} */,
  {32'h4087330c, 32'h40ea2e96} /* (1, 7, 9) {real, imag} */,
  {32'h3fe08b66, 32'h406801af} /* (1, 7, 8) {real, imag} */,
  {32'h417ee88c, 32'h419f2b42} /* (1, 7, 7) {real, imag} */,
  {32'hc1a97bb4, 32'h3f3ff140} /* (1, 7, 6) {real, imag} */,
  {32'h41cb9893, 32'h413c9979} /* (1, 7, 5) {real, imag} */,
  {32'h40a7cb65, 32'h40dfd3cb} /* (1, 7, 4) {real, imag} */,
  {32'h40fa32fe, 32'h41006d90} /* (1, 7, 3) {real, imag} */,
  {32'hc1bdf7ee, 32'h4008af30} /* (1, 7, 2) {real, imag} */,
  {32'h41b229dc, 32'hc1fdd1d8} /* (1, 7, 1) {real, imag} */,
  {32'h3fab8250, 32'h41457686} /* (1, 7, 0) {real, imag} */,
  {32'hc1b391fc, 32'hc19752c6} /* (1, 6, 15) {real, imag} */,
  {32'hc13cd022, 32'hc1c49840} /* (1, 6, 14) {real, imag} */,
  {32'hbfb19a4c, 32'hc221373c} /* (1, 6, 13) {real, imag} */,
  {32'h41cc7108, 32'hc1756044} /* (1, 6, 12) {real, imag} */,
  {32'h40e2bb9e, 32'hc1e6f015} /* (1, 6, 11) {real, imag} */,
  {32'hc10cf926, 32'h42846cbe} /* (1, 6, 10) {real, imag} */,
  {32'hc0985640, 32'hc0062b62} /* (1, 6, 9) {real, imag} */,
  {32'h411987e0, 32'h41857ff9} /* (1, 6, 8) {real, imag} */,
  {32'h418c9b2b, 32'h41c03324} /* (1, 6, 7) {real, imag} */,
  {32'hc17fd956, 32'h3f47eed8} /* (1, 6, 6) {real, imag} */,
  {32'hc1fe877a, 32'hc09a5b5d} /* (1, 6, 5) {real, imag} */,
  {32'hc21587db, 32'hc03ce22c} /* (1, 6, 4) {real, imag} */,
  {32'hc0558c90, 32'h40895de3} /* (1, 6, 3) {real, imag} */,
  {32'h41129206, 32'h41e2c9e8} /* (1, 6, 2) {real, imag} */,
  {32'hbf92e5ee, 32'h41c98dca} /* (1, 6, 1) {real, imag} */,
  {32'h4193160e, 32'hc0a4d301} /* (1, 6, 0) {real, imag} */,
  {32'h41c40eb9, 32'hc181e45c} /* (1, 5, 15) {real, imag} */,
  {32'h414a5559, 32'h408dd52c} /* (1, 5, 14) {real, imag} */,
  {32'h40f7c851, 32'hc0b17a84} /* (1, 5, 13) {real, imag} */,
  {32'h419274f7, 32'hc1aab85c} /* (1, 5, 12) {real, imag} */,
  {32'hc002b5c2, 32'h40fae564} /* (1, 5, 11) {real, imag} */,
  {32'hc0bdf697, 32'h41654c3d} /* (1, 5, 10) {real, imag} */,
  {32'h41e0e9c0, 32'h41497742} /* (1, 5, 9) {real, imag} */,
  {32'h40c49fc8, 32'hbebba490} /* (1, 5, 8) {real, imag} */,
  {32'h410fa710, 32'h40dc9782} /* (1, 5, 7) {real, imag} */,
  {32'h404e539e, 32'hc1e322ae} /* (1, 5, 6) {real, imag} */,
  {32'hc11ff478, 32'h41822f6e} /* (1, 5, 5) {real, imag} */,
  {32'hc1e58a12, 32'h413947ac} /* (1, 5, 4) {real, imag} */,
  {32'hc20ccd02, 32'h40df0a4e} /* (1, 5, 3) {real, imag} */,
  {32'h4223ef08, 32'hbe8e33f0} /* (1, 5, 2) {real, imag} */,
  {32'hc08e368c, 32'h42124cfa} /* (1, 5, 1) {real, imag} */,
  {32'hc1b16d8b, 32'hc1577b44} /* (1, 5, 0) {real, imag} */,
  {32'h42c92624, 32'h4261aa6f} /* (1, 4, 15) {real, imag} */,
  {32'hc1ad66b6, 32'h4214735c} /* (1, 4, 14) {real, imag} */,
  {32'h3fca6000, 32'hc1ae6dc0} /* (1, 4, 13) {real, imag} */,
  {32'hc192f67b, 32'h3fe46aec} /* (1, 4, 12) {real, imag} */,
  {32'hc1a7666e, 32'h40c53f0d} /* (1, 4, 11) {real, imag} */,
  {32'hbf3cc8a0, 32'hc22b2a60} /* (1, 4, 10) {real, imag} */,
  {32'h418697c0, 32'h41d10eaf} /* (1, 4, 9) {real, imag} */,
  {32'hc0972b39, 32'h40c88e9d} /* (1, 4, 8) {real, imag} */,
  {32'hc1495788, 32'h40bd6260} /* (1, 4, 7) {real, imag} */,
  {32'hc0470b7e, 32'h41d1583c} /* (1, 4, 6) {real, imag} */,
  {32'h418cc7ac, 32'h4197b78a} /* (1, 4, 5) {real, imag} */,
  {32'hbfafe2c8, 32'hc1f108d8} /* (1, 4, 4) {real, imag} */,
  {32'hc1cb445b, 32'hc25370e0} /* (1, 4, 3) {real, imag} */,
  {32'hc1cb4b7f, 32'hc1bfbdbb} /* (1, 4, 2) {real, imag} */,
  {32'h40fa1bf7, 32'hc1cfcaeb} /* (1, 4, 1) {real, imag} */,
  {32'hc16dca2a, 32'hc205c508} /* (1, 4, 0) {real, imag} */,
  {32'h41587dda, 32'hc2155c11} /* (1, 3, 15) {real, imag} */,
  {32'hc127c630, 32'hc05ea578} /* (1, 3, 14) {real, imag} */,
  {32'h40b87788, 32'h41810501} /* (1, 3, 13) {real, imag} */,
  {32'h41c68ae8, 32'hc18e8aae} /* (1, 3, 12) {real, imag} */,
  {32'hc1147b9c, 32'hc0fc0314} /* (1, 3, 11) {real, imag} */,
  {32'hbfaf9c64, 32'hc10c3fde} /* (1, 3, 10) {real, imag} */,
  {32'hc183431c, 32'hc0f561d0} /* (1, 3, 9) {real, imag} */,
  {32'hc012a874, 32'h40ad201e} /* (1, 3, 8) {real, imag} */,
  {32'hc24bb973, 32'hc15d4ac4} /* (1, 3, 7) {real, imag} */,
  {32'h40f52b4a, 32'hc198a854} /* (1, 3, 6) {real, imag} */,
  {32'hc083bfaa, 32'h3fd630c0} /* (1, 3, 5) {real, imag} */,
  {32'hbfc6cd38, 32'hc28d51bd} /* (1, 3, 4) {real, imag} */,
  {32'hc09ff6d9, 32'hc207321e} /* (1, 3, 3) {real, imag} */,
  {32'hc0ead5a4, 32'h41fcd2b6} /* (1, 3, 2) {real, imag} */,
  {32'hc14cfc17, 32'hc12712c6} /* (1, 3, 1) {real, imag} */,
  {32'h3f80697c, 32'h41f82c2a} /* (1, 3, 0) {real, imag} */,
  {32'hc26170ee, 32'h4251a3b8} /* (1, 2, 15) {real, imag} */,
  {32'hc0075950, 32'hc0831320} /* (1, 2, 14) {real, imag} */,
  {32'h40a682a4, 32'h40c153d0} /* (1, 2, 13) {real, imag} */,
  {32'h4110e681, 32'h40ae6d6c} /* (1, 2, 12) {real, imag} */,
  {32'hc235065b, 32'h40a5deac} /* (1, 2, 11) {real, imag} */,
  {32'hc18f8462, 32'hc148173e} /* (1, 2, 10) {real, imag} */,
  {32'h4126ae00, 32'h4183199d} /* (1, 2, 9) {real, imag} */,
  {32'hc0f2c1c4, 32'h410b3f4d} /* (1, 2, 8) {real, imag} */,
  {32'hc0b7a7ff, 32'hc1a2dfe7} /* (1, 2, 7) {real, imag} */,
  {32'hc181e3b6, 32'h4175d83a} /* (1, 2, 6) {real, imag} */,
  {32'h41119717, 32'h414d7d1f} /* (1, 2, 5) {real, imag} */,
  {32'hc113ea48, 32'h41c3b7c0} /* (1, 2, 4) {real, imag} */,
  {32'h421054f2, 32'h423225da} /* (1, 2, 3) {real, imag} */,
  {32'h413514ef, 32'h425b046d} /* (1, 2, 2) {real, imag} */,
  {32'h414c6744, 32'h41189737} /* (1, 2, 1) {real, imag} */,
  {32'h41cace17, 32'hc23c4bd4} /* (1, 2, 0) {real, imag} */,
  {32'hc2d34768, 32'h40e5f238} /* (1, 1, 15) {real, imag} */,
  {32'h41f526aa, 32'hc227c624} /* (1, 1, 14) {real, imag} */,
  {32'h4244732c, 32'h420cfabe} /* (1, 1, 13) {real, imag} */,
  {32'hc2274fce, 32'hc19d2324} /* (1, 1, 12) {real, imag} */,
  {32'h41ac2fd3, 32'hc1e0c1b4} /* (1, 1, 11) {real, imag} */,
  {32'hc0246506, 32'h40b34f52} /* (1, 1, 10) {real, imag} */,
  {32'hc1c87e6b, 32'hc246da04} /* (1, 1, 9) {real, imag} */,
  {32'hc0bfd506, 32'hc0a3c9a8} /* (1, 1, 8) {real, imag} */,
  {32'hc0378640, 32'hc100a2be} /* (1, 1, 7) {real, imag} */,
  {32'h41c666ec, 32'hc1cb2d66} /* (1, 1, 6) {real, imag} */,
  {32'hc25f40ae, 32'hc0e572ab} /* (1, 1, 5) {real, imag} */,
  {32'h40d03162, 32'hc13775d3} /* (1, 1, 4) {real, imag} */,
  {32'hc1b89010, 32'hc19a0c5f} /* (1, 1, 3) {real, imag} */,
  {32'hc253d6e2, 32'hbfb7d670} /* (1, 1, 2) {real, imag} */,
  {32'hc2729f75, 32'h4193a1c0} /* (1, 1, 1) {real, imag} */,
  {32'hc2fa6a7f, 32'h429c4211} /* (1, 1, 0) {real, imag} */,
  {32'h411b616c, 32'hc3336f08} /* (1, 0, 15) {real, imag} */,
  {32'h41124ffd, 32'h41f30546} /* (1, 0, 14) {real, imag} */,
  {32'h420c0a2f, 32'h425f3afc} /* (1, 0, 13) {real, imag} */,
  {32'h4280fd98, 32'hc1533dfa} /* (1, 0, 12) {real, imag} */,
  {32'h4222404e, 32'h423ae381} /* (1, 0, 11) {real, imag} */,
  {32'h402fa4b4, 32'hbf9171ec} /* (1, 0, 10) {real, imag} */,
  {32'h4121c26a, 32'h41752166} /* (1, 0, 9) {real, imag} */,
  {32'h41874c2e, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'h4121c26a, 32'hc1752166} /* (1, 0, 7) {real, imag} */,
  {32'h402fa4b4, 32'h3f9171ec} /* (1, 0, 6) {real, imag} */,
  {32'h4222404e, 32'hc23ae381} /* (1, 0, 5) {real, imag} */,
  {32'h4280fd98, 32'h41533dfa} /* (1, 0, 4) {real, imag} */,
  {32'h420c0a2f, 32'hc25f3afc} /* (1, 0, 3) {real, imag} */,
  {32'h41124ffd, 32'hc1f30546} /* (1, 0, 2) {real, imag} */,
  {32'h411b616c, 32'h43336f08} /* (1, 0, 1) {real, imag} */,
  {32'h410b1848, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hc148663a, 32'hc2a08bab} /* (0, 15, 15) {real, imag} */,
  {32'hc1d7e852, 32'hc1a12a76} /* (0, 15, 14) {real, imag} */,
  {32'hc040d86c, 32'hc0469b90} /* (0, 15, 13) {real, imag} */,
  {32'h4168c156, 32'h410edf9e} /* (0, 15, 12) {real, imag} */,
  {32'hc1bbb0de, 32'h4142cba8} /* (0, 15, 11) {real, imag} */,
  {32'h41eb3b2e, 32'hc14f95e3} /* (0, 15, 10) {real, imag} */,
  {32'h41067df5, 32'hc0c0631c} /* (0, 15, 9) {real, imag} */,
  {32'hc17f3528, 32'hbf8e9db8} /* (0, 15, 8) {real, imag} */,
  {32'h403969c8, 32'hbfd58478} /* (0, 15, 7) {real, imag} */,
  {32'hc117a7c7, 32'h3fa1353c} /* (0, 15, 6) {real, imag} */,
  {32'hc178744e, 32'hbf7756b0} /* (0, 15, 5) {real, imag} */,
  {32'h41ab869e, 32'h414aa3b2} /* (0, 15, 4) {real, imag} */,
  {32'hc1da57e4, 32'hc2164e64} /* (0, 15, 3) {real, imag} */,
  {32'hc162391c, 32'h4248eb2a} /* (0, 15, 2) {real, imag} */,
  {32'hc28f887c, 32'hc2192641} /* (0, 15, 1) {real, imag} */,
  {32'hc2938ef8, 32'hc20e29b0} /* (0, 15, 0) {real, imag} */,
  {32'h40b35588, 32'hc12de8ac} /* (0, 14, 15) {real, imag} */,
  {32'hbf09ece0, 32'hc18b10fa} /* (0, 14, 14) {real, imag} */,
  {32'h421849af, 32'hc1d7a008} /* (0, 14, 13) {real, imag} */,
  {32'h3fa556c0, 32'h408a3769} /* (0, 14, 12) {real, imag} */,
  {32'hc11fa8ca, 32'h41089cc3} /* (0, 14, 11) {real, imag} */,
  {32'hbedbbd70, 32'h3f072a80} /* (0, 14, 10) {real, imag} */,
  {32'h412c9331, 32'h41d03f7a} /* (0, 14, 9) {real, imag} */,
  {32'h41912a30, 32'hc1223bfc} /* (0, 14, 8) {real, imag} */,
  {32'hc13468b0, 32'h4109cdb0} /* (0, 14, 7) {real, imag} */,
  {32'hc0a1c68c, 32'hc0ccb583} /* (0, 14, 6) {real, imag} */,
  {32'h416a2dd5, 32'h41dbd34c} /* (0, 14, 5) {real, imag} */,
  {32'h4164d91d, 32'h4116d3be} /* (0, 14, 4) {real, imag} */,
  {32'h400a09ba, 32'hc1aae2c6} /* (0, 14, 3) {real, imag} */,
  {32'hc173acfc, 32'hc1b18dcd} /* (0, 14, 2) {real, imag} */,
  {32'hc1b751d5, 32'hc25def86} /* (0, 14, 1) {real, imag} */,
  {32'hc12b5071, 32'h41ce7c89} /* (0, 14, 0) {real, imag} */,
  {32'hc14763a0, 32'h414721c6} /* (0, 13, 15) {real, imag} */,
  {32'hc0d9473d, 32'hc15cbd1c} /* (0, 13, 14) {real, imag} */,
  {32'h411ffeb4, 32'h41259684} /* (0, 13, 13) {real, imag} */,
  {32'hc12e08e2, 32'h41de11be} /* (0, 13, 12) {real, imag} */,
  {32'h40528378, 32'h41343c80} /* (0, 13, 11) {real, imag} */,
  {32'h40a90114, 32'h40ed5047} /* (0, 13, 10) {real, imag} */,
  {32'hc18eae6c, 32'h4191062a} /* (0, 13, 9) {real, imag} */,
  {32'h40de5b79, 32'hc1458d91} /* (0, 13, 8) {real, imag} */,
  {32'hc101291e, 32'h417e065c} /* (0, 13, 7) {real, imag} */,
  {32'hc0c046ca, 32'hc0f20bcc} /* (0, 13, 6) {real, imag} */,
  {32'h41da327a, 32'h418a297d} /* (0, 13, 5) {real, imag} */,
  {32'h4204cb62, 32'h40ccd6db} /* (0, 13, 4) {real, imag} */,
  {32'h3f76eec0, 32'hc1662bc0} /* (0, 13, 3) {real, imag} */,
  {32'h419717b4, 32'hbf5cc798} /* (0, 13, 2) {real, imag} */,
  {32'hc11e91f7, 32'h412ab6a4} /* (0, 13, 1) {real, imag} */,
  {32'hc1a9a434, 32'hc14b6f83} /* (0, 13, 0) {real, imag} */,
  {32'h41daad56, 32'h412eb4ea} /* (0, 12, 15) {real, imag} */,
  {32'hc1bf81de, 32'hbeca2d00} /* (0, 12, 14) {real, imag} */,
  {32'hc1e533d3, 32'h42533cf4} /* (0, 12, 13) {real, imag} */,
  {32'hc212ea4d, 32'h4001e814} /* (0, 12, 12) {real, imag} */,
  {32'h41a527f3, 32'hc10f9637} /* (0, 12, 11) {real, imag} */,
  {32'hc0e51646, 32'hc11fc4d4} /* (0, 12, 10) {real, imag} */,
  {32'h409f0ad6, 32'h4182a235} /* (0, 12, 9) {real, imag} */,
  {32'h4173c34a, 32'h4159b36d} /* (0, 12, 8) {real, imag} */,
  {32'h40da61c3, 32'hc1bad7e6} /* (0, 12, 7) {real, imag} */,
  {32'h4183150e, 32'h40c4195a} /* (0, 12, 6) {real, imag} */,
  {32'hc16b4847, 32'h41c072be} /* (0, 12, 5) {real, imag} */,
  {32'hbf652420, 32'hc07bfa5c} /* (0, 12, 4) {real, imag} */,
  {32'hc08dae78, 32'h401536b0} /* (0, 12, 3) {real, imag} */,
  {32'hc0338013, 32'hc1898d7e} /* (0, 12, 2) {real, imag} */,
  {32'h424994ae, 32'hc1a21cb5} /* (0, 12, 1) {real, imag} */,
  {32'hc0ef97f6, 32'h41cff6e2} /* (0, 12, 0) {real, imag} */,
  {32'h40e9fee8, 32'hc1e264b0} /* (0, 11, 15) {real, imag} */,
  {32'hc10383cd, 32'h41593999} /* (0, 11, 14) {real, imag} */,
  {32'hc121d186, 32'hc0a51d06} /* (0, 11, 13) {real, imag} */,
  {32'hc0de35da, 32'h410f5f3e} /* (0, 11, 12) {real, imag} */,
  {32'h41d5d57d, 32'hc13c9566} /* (0, 11, 11) {real, imag} */,
  {32'hc18e7828, 32'h40f55f7b} /* (0, 11, 10) {real, imag} */,
  {32'hc0472e0c, 32'hc02d0627} /* (0, 11, 9) {real, imag} */,
  {32'hbe190540, 32'h408f785a} /* (0, 11, 8) {real, imag} */,
  {32'h41534a2e, 32'hbfe70e68} /* (0, 11, 7) {real, imag} */,
  {32'hc0075632, 32'hc04b4b54} /* (0, 11, 6) {real, imag} */,
  {32'h41183a3e, 32'h3febac20} /* (0, 11, 5) {real, imag} */,
  {32'h4154a3d0, 32'h406222d4} /* (0, 11, 4) {real, imag} */,
  {32'hc1e1d1d2, 32'hc16a73c2} /* (0, 11, 3) {real, imag} */,
  {32'h3f015cb8, 32'h41701a78} /* (0, 11, 2) {real, imag} */,
  {32'hc11bc63e, 32'h41250887} /* (0, 11, 1) {real, imag} */,
  {32'hc13545ac, 32'h401e2caa} /* (0, 11, 0) {real, imag} */,
  {32'hc19139b4, 32'h3ff51570} /* (0, 10, 15) {real, imag} */,
  {32'h418aca8f, 32'h40d3af97} /* (0, 10, 14) {real, imag} */,
  {32'hc1902350, 32'h41d98768} /* (0, 10, 13) {real, imag} */,
  {32'h401b016c, 32'hc12d24b7} /* (0, 10, 12) {real, imag} */,
  {32'hc0f5941c, 32'h419fb8f8} /* (0, 10, 11) {real, imag} */,
  {32'hc10a60ff, 32'hc184600b} /* (0, 10, 10) {real, imag} */,
  {32'h3fc7876c, 32'hc12b4b2a} /* (0, 10, 9) {real, imag} */,
  {32'h4139b89e, 32'hc0c2c9a8} /* (0, 10, 8) {real, imag} */,
  {32'h410c8048, 32'hc035614c} /* (0, 10, 7) {real, imag} */,
  {32'h4194a831, 32'h415e6a74} /* (0, 10, 6) {real, imag} */,
  {32'hc1b25178, 32'hc1368a87} /* (0, 10, 5) {real, imag} */,
  {32'h410e5752, 32'h40886821} /* (0, 10, 4) {real, imag} */,
  {32'h4029185c, 32'h41ddd5d2} /* (0, 10, 3) {real, imag} */,
  {32'hc16aab08, 32'h411bf8c6} /* (0, 10, 2) {real, imag} */,
  {32'hc1443ffc, 32'h41510833} /* (0, 10, 1) {real, imag} */,
  {32'hc09764a4, 32'hc1260e8e} /* (0, 10, 0) {real, imag} */,
  {32'hc100e875, 32'h419009b4} /* (0, 9, 15) {real, imag} */,
  {32'hc058223a, 32'h40541016} /* (0, 9, 14) {real, imag} */,
  {32'hbf9a9db0, 32'hc11c45ee} /* (0, 9, 13) {real, imag} */,
  {32'h40cca518, 32'hc128a738} /* (0, 9, 12) {real, imag} */,
  {32'h40f83304, 32'h4196dd2c} /* (0, 9, 11) {real, imag} */,
  {32'hbf43dae0, 32'h41135607} /* (0, 9, 10) {real, imag} */,
  {32'h40e7a27e, 32'hc10a1218} /* (0, 9, 9) {real, imag} */,
  {32'h410fe7c4, 32'hc0bf0fd9} /* (0, 9, 8) {real, imag} */,
  {32'hc1d282a2, 32'h415c97cb} /* (0, 9, 7) {real, imag} */,
  {32'h41bca1b6, 32'h41726b42} /* (0, 9, 6) {real, imag} */,
  {32'hc0e5ca50, 32'hc0437bb7} /* (0, 9, 5) {real, imag} */,
  {32'hc1c0d0b3, 32'h40e5a51c} /* (0, 9, 4) {real, imag} */,
  {32'h41da5b12, 32'hc0448294} /* (0, 9, 3) {real, imag} */,
  {32'hc104bbc0, 32'hc1d0fc74} /* (0, 9, 2) {real, imag} */,
  {32'h3ef7aac0, 32'h3faca5c0} /* (0, 9, 1) {real, imag} */,
  {32'h41cb79a5, 32'h3fe5925c} /* (0, 9, 0) {real, imag} */,
  {32'h41d719b5, 32'hc156d468} /* (0, 8, 15) {real, imag} */,
  {32'hc10776a1, 32'h4109a9bf} /* (0, 8, 14) {real, imag} */,
  {32'h4082ee36, 32'hbfbfec8c} /* (0, 8, 13) {real, imag} */,
  {32'h40602296, 32'hc10395db} /* (0, 8, 12) {real, imag} */,
  {32'hc05f225c, 32'h412a9755} /* (0, 8, 11) {real, imag} */,
  {32'h417949e8, 32'hc16cca12} /* (0, 8, 10) {real, imag} */,
  {32'h411678d0, 32'h41825999} /* (0, 8, 9) {real, imag} */,
  {32'hc1143e24, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'h411678d0, 32'hc1825999} /* (0, 8, 7) {real, imag} */,
  {32'h417949e8, 32'h416cca12} /* (0, 8, 6) {real, imag} */,
  {32'hc05f225c, 32'hc12a9755} /* (0, 8, 5) {real, imag} */,
  {32'h40602296, 32'h410395db} /* (0, 8, 4) {real, imag} */,
  {32'h4082ee36, 32'h3fbfec8c} /* (0, 8, 3) {real, imag} */,
  {32'hc10776a1, 32'hc109a9bf} /* (0, 8, 2) {real, imag} */,
  {32'h41d719b5, 32'h4156d468} /* (0, 8, 1) {real, imag} */,
  {32'hc1a24fac, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h3ef7aac0, 32'hbfaca5c0} /* (0, 7, 15) {real, imag} */,
  {32'hc104bbc0, 32'h41d0fc74} /* (0, 7, 14) {real, imag} */,
  {32'h41da5b12, 32'h40448294} /* (0, 7, 13) {real, imag} */,
  {32'hc1c0d0b3, 32'hc0e5a51c} /* (0, 7, 12) {real, imag} */,
  {32'hc0e5ca50, 32'h40437bb7} /* (0, 7, 11) {real, imag} */,
  {32'h41bca1b6, 32'hc1726b42} /* (0, 7, 10) {real, imag} */,
  {32'hc1d282a2, 32'hc15c97cb} /* (0, 7, 9) {real, imag} */,
  {32'h410fe7c4, 32'h40bf0fd9} /* (0, 7, 8) {real, imag} */,
  {32'h40e7a27e, 32'h410a1218} /* (0, 7, 7) {real, imag} */,
  {32'hbf43dae0, 32'hc1135607} /* (0, 7, 6) {real, imag} */,
  {32'h40f83304, 32'hc196dd2c} /* (0, 7, 5) {real, imag} */,
  {32'h40cca518, 32'h4128a738} /* (0, 7, 4) {real, imag} */,
  {32'hbf9a9db0, 32'h411c45ee} /* (0, 7, 3) {real, imag} */,
  {32'hc058223a, 32'hc0541016} /* (0, 7, 2) {real, imag} */,
  {32'hc100e875, 32'hc19009b4} /* (0, 7, 1) {real, imag} */,
  {32'h41cb79a5, 32'hbfe5925c} /* (0, 7, 0) {real, imag} */,
  {32'hc1443ffc, 32'hc1510833} /* (0, 6, 15) {real, imag} */,
  {32'hc16aab08, 32'hc11bf8c6} /* (0, 6, 14) {real, imag} */,
  {32'h4029185c, 32'hc1ddd5d2} /* (0, 6, 13) {real, imag} */,
  {32'h410e5752, 32'hc0886821} /* (0, 6, 12) {real, imag} */,
  {32'hc1b25178, 32'h41368a87} /* (0, 6, 11) {real, imag} */,
  {32'h4194a831, 32'hc15e6a74} /* (0, 6, 10) {real, imag} */,
  {32'h410c8048, 32'h4035614c} /* (0, 6, 9) {real, imag} */,
  {32'h4139b89e, 32'h40c2c9a8} /* (0, 6, 8) {real, imag} */,
  {32'h3fc7876c, 32'h412b4b2a} /* (0, 6, 7) {real, imag} */,
  {32'hc10a60ff, 32'h4184600b} /* (0, 6, 6) {real, imag} */,
  {32'hc0f5941c, 32'hc19fb8f8} /* (0, 6, 5) {real, imag} */,
  {32'h401b016c, 32'h412d24b7} /* (0, 6, 4) {real, imag} */,
  {32'hc1902350, 32'hc1d98768} /* (0, 6, 3) {real, imag} */,
  {32'h418aca8f, 32'hc0d3af97} /* (0, 6, 2) {real, imag} */,
  {32'hc19139b4, 32'hbff51570} /* (0, 6, 1) {real, imag} */,
  {32'hc09764a4, 32'h41260e8e} /* (0, 6, 0) {real, imag} */,
  {32'hc11bc63e, 32'hc1250887} /* (0, 5, 15) {real, imag} */,
  {32'h3f015cb8, 32'hc1701a78} /* (0, 5, 14) {real, imag} */,
  {32'hc1e1d1d2, 32'h416a73c2} /* (0, 5, 13) {real, imag} */,
  {32'h4154a3d0, 32'hc06222d4} /* (0, 5, 12) {real, imag} */,
  {32'h41183a3e, 32'hbfebac20} /* (0, 5, 11) {real, imag} */,
  {32'hc0075632, 32'h404b4b54} /* (0, 5, 10) {real, imag} */,
  {32'h41534a2e, 32'h3fe70e68} /* (0, 5, 9) {real, imag} */,
  {32'hbe190540, 32'hc08f785a} /* (0, 5, 8) {real, imag} */,
  {32'hc0472e0c, 32'h402d0627} /* (0, 5, 7) {real, imag} */,
  {32'hc18e7828, 32'hc0f55f7b} /* (0, 5, 6) {real, imag} */,
  {32'h41d5d57d, 32'h413c9566} /* (0, 5, 5) {real, imag} */,
  {32'hc0de35da, 32'hc10f5f3e} /* (0, 5, 4) {real, imag} */,
  {32'hc121d186, 32'h40a51d06} /* (0, 5, 3) {real, imag} */,
  {32'hc10383cd, 32'hc1593999} /* (0, 5, 2) {real, imag} */,
  {32'h40e9fee8, 32'h41e264b0} /* (0, 5, 1) {real, imag} */,
  {32'hc13545ac, 32'hc01e2caa} /* (0, 5, 0) {real, imag} */,
  {32'h424994ae, 32'h41a21cb5} /* (0, 4, 15) {real, imag} */,
  {32'hc0338013, 32'h41898d7e} /* (0, 4, 14) {real, imag} */,
  {32'hc08dae78, 32'hc01536b0} /* (0, 4, 13) {real, imag} */,
  {32'hbf652420, 32'h407bfa5c} /* (0, 4, 12) {real, imag} */,
  {32'hc16b4847, 32'hc1c072be} /* (0, 4, 11) {real, imag} */,
  {32'h4183150e, 32'hc0c4195a} /* (0, 4, 10) {real, imag} */,
  {32'h40da61c3, 32'h41bad7e6} /* (0, 4, 9) {real, imag} */,
  {32'h4173c34a, 32'hc159b36d} /* (0, 4, 8) {real, imag} */,
  {32'h409f0ad6, 32'hc182a235} /* (0, 4, 7) {real, imag} */,
  {32'hc0e51646, 32'h411fc4d4} /* (0, 4, 6) {real, imag} */,
  {32'h41a527f3, 32'h410f9637} /* (0, 4, 5) {real, imag} */,
  {32'hc212ea4d, 32'hc001e814} /* (0, 4, 4) {real, imag} */,
  {32'hc1e533d3, 32'hc2533cf4} /* (0, 4, 3) {real, imag} */,
  {32'hc1bf81de, 32'h3eca2d00} /* (0, 4, 2) {real, imag} */,
  {32'h41daad56, 32'hc12eb4ea} /* (0, 4, 1) {real, imag} */,
  {32'hc0ef97f6, 32'hc1cff6e2} /* (0, 4, 0) {real, imag} */,
  {32'hc11e91f7, 32'hc12ab6a4} /* (0, 3, 15) {real, imag} */,
  {32'h419717b4, 32'h3f5cc798} /* (0, 3, 14) {real, imag} */,
  {32'h3f76eec0, 32'h41662bc0} /* (0, 3, 13) {real, imag} */,
  {32'h4204cb62, 32'hc0ccd6db} /* (0, 3, 12) {real, imag} */,
  {32'h41da327a, 32'hc18a297d} /* (0, 3, 11) {real, imag} */,
  {32'hc0c046ca, 32'h40f20bcc} /* (0, 3, 10) {real, imag} */,
  {32'hc101291e, 32'hc17e065c} /* (0, 3, 9) {real, imag} */,
  {32'h40de5b79, 32'h41458d91} /* (0, 3, 8) {real, imag} */,
  {32'hc18eae6c, 32'hc191062a} /* (0, 3, 7) {real, imag} */,
  {32'h40a90114, 32'hc0ed5047} /* (0, 3, 6) {real, imag} */,
  {32'h40528378, 32'hc1343c80} /* (0, 3, 5) {real, imag} */,
  {32'hc12e08e2, 32'hc1de11be} /* (0, 3, 4) {real, imag} */,
  {32'h411ffeb4, 32'hc1259684} /* (0, 3, 3) {real, imag} */,
  {32'hc0d9473d, 32'h415cbd1c} /* (0, 3, 2) {real, imag} */,
  {32'hc14763a0, 32'hc14721c6} /* (0, 3, 1) {real, imag} */,
  {32'hc1a9a434, 32'h414b6f83} /* (0, 3, 0) {real, imag} */,
  {32'hc1b751d5, 32'h425def86} /* (0, 2, 15) {real, imag} */,
  {32'hc173acfc, 32'h41b18dcd} /* (0, 2, 14) {real, imag} */,
  {32'h400a09ba, 32'h41aae2c6} /* (0, 2, 13) {real, imag} */,
  {32'h4164d91d, 32'hc116d3be} /* (0, 2, 12) {real, imag} */,
  {32'h416a2dd5, 32'hc1dbd34c} /* (0, 2, 11) {real, imag} */,
  {32'hc0a1c68c, 32'h40ccb583} /* (0, 2, 10) {real, imag} */,
  {32'hc13468b0, 32'hc109cdb0} /* (0, 2, 9) {real, imag} */,
  {32'h41912a30, 32'h41223bfc} /* (0, 2, 8) {real, imag} */,
  {32'h412c9331, 32'hc1d03f7a} /* (0, 2, 7) {real, imag} */,
  {32'hbedbbd70, 32'hbf072a80} /* (0, 2, 6) {real, imag} */,
  {32'hc11fa8ca, 32'hc1089cc3} /* (0, 2, 5) {real, imag} */,
  {32'h3fa556c0, 32'hc08a3769} /* (0, 2, 4) {real, imag} */,
  {32'h421849af, 32'h41d7a008} /* (0, 2, 3) {real, imag} */,
  {32'hbf09ece0, 32'h418b10fa} /* (0, 2, 2) {real, imag} */,
  {32'h40b35588, 32'h412de8ac} /* (0, 2, 1) {real, imag} */,
  {32'hc12b5071, 32'hc1ce7c89} /* (0, 2, 0) {real, imag} */,
  {32'hc28f887c, 32'h42192641} /* (0, 1, 15) {real, imag} */,
  {32'hc162391c, 32'hc248eb2a} /* (0, 1, 14) {real, imag} */,
  {32'hc1da57e4, 32'h42164e64} /* (0, 1, 13) {real, imag} */,
  {32'h41ab869e, 32'hc14aa3b2} /* (0, 1, 12) {real, imag} */,
  {32'hc178744e, 32'h3f7756b0} /* (0, 1, 11) {real, imag} */,
  {32'hc117a7c7, 32'hbfa1353c} /* (0, 1, 10) {real, imag} */,
  {32'h403969c8, 32'h3fd58478} /* (0, 1, 9) {real, imag} */,
  {32'hc17f3528, 32'h3f8e9db8} /* (0, 1, 8) {real, imag} */,
  {32'h41067df5, 32'h40c0631c} /* (0, 1, 7) {real, imag} */,
  {32'h41eb3b2e, 32'h414f95e3} /* (0, 1, 6) {real, imag} */,
  {32'hc1bbb0de, 32'hc142cba8} /* (0, 1, 5) {real, imag} */,
  {32'h4168c156, 32'hc10edf9e} /* (0, 1, 4) {real, imag} */,
  {32'hc040d86c, 32'h40469b90} /* (0, 1, 3) {real, imag} */,
  {32'hc1d7e852, 32'h41a12a76} /* (0, 1, 2) {real, imag} */,
  {32'hc148663a, 32'h42a08bab} /* (0, 1, 1) {real, imag} */,
  {32'hc2938ef8, 32'h420e29b0} /* (0, 1, 0) {real, imag} */,
  {32'h42037162, 32'hc3091250} /* (0, 0, 15) {real, imag} */,
  {32'h40767560, 32'h4216b3e4} /* (0, 0, 14) {real, imag} */,
  {32'h41f51d6b, 32'h41c242fa} /* (0, 0, 13) {real, imag} */,
  {32'h41425cad, 32'hc11562b4} /* (0, 0, 12) {real, imag} */,
  {32'h3f0e6ea0, 32'h414f6ff7} /* (0, 0, 11) {real, imag} */,
  {32'hc0969d7b, 32'h415a50fb} /* (0, 0, 10) {real, imag} */,
  {32'h41175ad1, 32'hc04442ca} /* (0, 0, 9) {real, imag} */,
  {32'hc1129416, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h41175ad1, 32'h404442ca} /* (0, 0, 7) {real, imag} */,
  {32'hc0969d7b, 32'hc15a50fb} /* (0, 0, 6) {real, imag} */,
  {32'h3f0e6ea0, 32'hc14f6ff7} /* (0, 0, 5) {real, imag} */,
  {32'h41425cad, 32'h411562b4} /* (0, 0, 4) {real, imag} */,
  {32'h41f51d6b, 32'hc1c242fa} /* (0, 0, 3) {real, imag} */,
  {32'h40767560, 32'hc216b3e4} /* (0, 0, 2) {real, imag} */,
  {32'h42037162, 32'h43091250} /* (0, 0, 1) {real, imag} */,
  {32'hc061ade0, 32'h00000000} /* (0, 0, 0) {real, imag} */};
