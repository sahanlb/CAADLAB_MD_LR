-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kRVDptRRA60+3RYOeyOPK2VCO+XsQ9N+7O8no+eaxPSuxkLkS8mvAM6XZQwNVJOCyHhVi+iw/Wdl
Hxn8wz9IUkwAgS92aLKZLmi0i5bjRXpuMRqS82BOJkJ9IpEVkxA64iH9yA60YjGASS+xunURUY13
zrocAVQvRPXUOoxTpvsROY8DqX9thlbO4bfq7xx3UEnGyvw/+XB8whLxbRyuJzXM/9mECyTIDKET
7jzKvkrYFc4bGXLSn4bFw5nQdUhoz44tFv3sFbO2vlQf86nAy/BYhJOhhuWmLfHj5/IYIZgTGZJU
KwK/KU6AwJCtKYQqJXaJ/ipW0XIGnjGAYO82lQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4304)
`protect data_block
rK+9i/SqwqvbkMlog/8xv2Dt8+wG7lo0id1dzIckEgI/GWOrHmfLLAnMwxsWqAJ/W6+pAl+07t2q
e4sGKiXz3Jxd8YsDjAxsAG1+ODPB0B6V0VEoTEYZNBcxNi+ZgOkRtz4qoTULfd7pP1jolnhf2Iru
D6t+weMcxsbdS8nfDbsEWAbU8+DrdHVxaapLRbleZyddo42/moqEboBS7W48MnRoq9efHu4Skqzt
XmSp9GmhL+pUiL7yAa/bJyzPf6n60joRVRpoAhkPh70MuxqH65zIyi51nZckoTqzEcRcGZkkWVRx
cBuLm2VRyKkWwbcRaX/qG7FAj4GkIRYyrd3LXXoDKKeScOjAzM3uBh97krVxLWj4q6/VvAtlSVtg
J/UwZhr5wu0TR8TG1/o/qYvrSTVR5SVk6jsQ6Sqy4L1GeEgaXNPsvVFMOosOyigeZ087BOKqQ4Qq
usyKJzvMohPANbXn473i1QHARR8OLUcbU7VQWBNrRn/OMLzHkv1ztjmHSEH/AvaxbL/TqDbhL6FV
7C+ePqZmkSic+6OAfsojxeJebsmr9YkASMPlJqU2S5e6kfjHW7ZjBxw+tLWD1BlVMGnwFu87+pFd
7djxdMtYA698xGmeAHh4QAI6OLQfhcGA+6mvqADIlfeDWs/eZs49UW3W2zyht7lSYIBYNWQoXhYO
JpITY5XWsnonAAmiZgTJqPFwEwA+L1/93rbkjX+KIP6Hj40GWzm6jFh3oJhyucltY/MsC8AmfDQ5
5P38ffMCeTK5CfaNOlmSNS6v2iIk1jcAVrYtIPGledXzfXDbDYGbd5e8Nc8gwt9dMHUtmaLyjYjS
WvSAFAUj6DX9tNEA3WKy2ZfMBttudAvK+4y8yeA0+GjPvZYNgytYZqZd/VIZ9akuJT77S74xhhIE
nK1A2z/q3w3V4Sue8IXZQcQhUyrZakwQ1VO06sM5okxXlIG5DoMkhS569Od/lSNWozSihYCVLTlN
svdxzuLFqeg+KrlCTE8WFJ7c1jNSvBqMiy1dqhpbNWuJJYKh/XeOlNEuvVstf18GRZ22VqNPQAOd
GvcqmX/wLOaByyLpAPX02PpYnZCniPT4Nogc2MPGJu4SCclX2V+YPhM/1L1UxoPuPLIKbv9YDLjH
cnQKsGFKT1okFSg831kyDZddbZJJ3vSoOBnOnfHMQYsidBxYM8BHpnEAeq3RB5L7m6e5zn6BALPy
m91jGrr43GV/gfxC4uL2icr4uMDiBXZizVeo6a2sbuKMx1Rd/S1RjqbYlXqIxBApqCk9axyqHwji
7VHpNZGV6BF6z38TKIa3o7Su2WZ6/Rup1geboUX6HWYZFiKG8bWdELcUfVAOMJDmHPyKulydVKt/
BH4BVAcaRLrDyu0ahEJd6DCFIkCfIKyozAI0sCGrt+dPyXzbs1gCxiaEZykZ0gH4ll1kVcvVsiBd
hHd0G+ZI3Gj5YjZaY197eJFnpotJJJWezyE/H3T9yyUExmKJeBg5tOUwV38vgaI7CWuc4HI9gyAz
QF7Ud2+hEswJP+OaFLAFC1TyKqNete/jDPWtNOLonanCogYxs0HkQfaNgGv0lMeQNjubjHRMZeJv
TP2PSlIyyUvBeVJjBKvFTKH2TCTefYsnQ78x1yyBBPlxwK1AkvkO4fcuJjrFavviRSsbTSZZZ/0r
baUQ7Gn5nViDY4pzraT/TgXHRZIAaP8z4CnivDSTjFAP0TffkVnytwVg4pUYLW4H+Rm/3umQ1Rpn
iiQx50zRY4ign1sOmLlG/Bh3TdJugsixcVkpmbkrzsxY4sAwjJ4JKPpg31DhHUCp43QTRfqPZiha
zn1M9LYIJSbaTP08ipGT8+lQDkgK6ZFttPLXrjW5QsRhcIDTD3Esgx1ptIlTk0bvhSv/HSNS1mtn
p8BCE1GqyD6EmqUFdmaE7v7PznGYiXdC6W+eZgCskjw+k5mRInVjqPnRTEi+NO5oyZfB5naYZR7X
+dySjp9gsJoprwpQbOJsWUXMPNA0OKiYBY+PgdX0dbmMxqXg/dE9Hs9xVfJPjDtuRoqVjL+/PmYs
7LONTDdH9A1QNMZ0ylzMRXJ6s7V20KvY1I2fyQypEhVLH1dgpYGRicQTwZpriwd3ib6hFLfgPRgA
eTG1Cso9slud9AFMV3mZnS5heI+XHR/Vxd9gQabrferuotS7s9IaA3iTsqqI9OyXR0P+lGyDTb+7
W46+NwWTTQeyzJvJ4lNAq2xFjec4NJg5z6YPhMPHSYp7oGtfmHRVxG7NH0WUBQALgMa4MDbypLWF
jABoaABtoup3PfQwOwVzDlHFWeLkYDfTq55YohIeiY615pRQ7U6KYCmk0SeiRmFuVf7LFatLwOVS
OIp1H6o2UDxG5+BFIOxIXi7ovDVRmQhXP1EnoJyeiG0Yf5Lq/Yigfo3m4TcWRIH75kq6txuocmr4
w1cTH/ofLME878vFIXTdJDXAjPWFeTvuNMziGwPL5B9F2FXL4koQrgfk56r44E+ATvCnUAtaybKr
JndsbKMFiT9kXELZkcK7e9tCQY6LQNW7PK6t8JxW55r4Y0q7y7810hZtPljdFCM1e838ceTLpr+Z
SpHulUiKb9X8kAD8bP4dtbDqFX//cFfNQU1kruPNPuteEZcnVnMs1+5rkr1fWKeJqr3J7IoJ+OZC
hVnquvVSg1eqvTkBXxpLmD6lvNUDTagl+pxd76C8+tGAFgfxpLOGzp5qoc2l4RJH96vnUqSbQOC5
Jx4StYZDKhEJDcAQQUmghDVwwkdXCDuaPWlZt2D0zD7wi73mBE2FkzKm6Cq4mJwDyimmLPH7eWfP
BRU1TEAt54s0b4+s2IV7f+oUVeSe4hkNjgdhfK/Qh5KnMvWEZdJLQTjwkZWlyqU33C6qo/yep21J
OWG485FMh3aeh7rS8eN/L90YedOSHhUjorB6fxfkw/TKJXT45yU/Xgkqnxf2kUxzNzXFzLXvqPTG
Cv+vbGOnOZEtzqZHpHLydFz5RIm7Mv2Iga+pDS5rtZRlEeBivHxnVhndijpZoRnALrhSap5/PnJK
yH5juIi4ARbqKf/skDhM2eytJ/DlGjy+cuyVcqCJG4o3LmAZAk8jWm/Ovek0WMFB+D29DC7Nij2W
ExJQdRe0WX4aeYrj1R82duKFk/oAO5vUDYiRgkO0N6it9c8iAtDiki3Q7vwusRbNH/KS0VoV9nFV
goGeQrhPuH6aTH8co78f07iySCYZsSfFtOP4fW95WTjHtCBeQBoMIDcLcQOcuoIAlfEYvDH/jAQr
+Bkp7qsU2E9BdDm4pGM79rJAZ+LWJO8Xoy+7lOludSW77WjS0BxKVNd2Mb8F7R7YyfpaNjRJpPpc
UH0zMd/7yB/RBT6bMXUPq/1RCreX+IIZyOnEsj5J+nXVnf4dvpyt25lp/mn5t3OwCXI/OAiuItju
PPISMPHvkFTZek8rliO3NifPKqTxM/2uLEa2KjlHvvnBUELCstfTYxBwRHaYvm7CS3F+nBUBLvxZ
xrwWkZr9BuJTqPR8Gpj78zXR1cw3anOlarq1gIyElTbhrbEP51udBTJ9IUs+QmWFCo5o8h6v1S2g
l3sXxc+WYLt4VeRLK414ajPps+XY+pnvkserNHgpQoZW1CIhalGoiysnGlXAePR8HdGTKwzcSPEA
3w+Juh4vpSutbObJYsvsqIGxBCGCak2Lfvxp+xX8AqeTUusDIRIrpN9tbwTa6o9o2tPswYHc7lF5
YBIqAe2kl89+eiO9aijw82iA3xAllX9o5Y5zpGfWub1cuc1XJGBBL4LJQ25ZfVqm0YLpJN+dyg5t
v9+UHAeu62Err1Gtgso0xmlb+sRUTCgAgrviFJbzJrKn/bHXapK0Dw54b6V3RX175by7BuwZ2VYU
D4E+SKTxhw3CLmrhh4aU3+ElZwcJFxSOaGMxUs+Po52y7XMEw3NeLX5pDI5PJuXb+clGqEAvM+Zz
NQ4hJnHT41N/SHpXkcr4vrwuRusho3GgBVPNdGuKY8mbIT6/Am1Jg7Kq73307r2SfgqJr1nsb2XA
wKJ62sS6IEKHwW1z9GzDY+PUI9g02Kd1dcIxRCj6a0PmLZhfYwcdo5+LLjBaPqUTKJp9XQXZWmMs
DDpeAGD5SxL7D2jXZqLZAzPUhALHSdYCiHhPlUVVrl3X79bEQQWrVobDUSkQhDdW7CLYLXHL+rHK
BI8cxKFdarpCdr1yjeAuCp+ltO22XAu4qaM27RhQKPycxCPoGxqewjWCORBodOAoE9AucF1TdWwC
OJX5wuvBK1UsJ/0EWGa+SIdYrEPxSWfNLWaLQQocIbA4Tvp7rR0mAX0gE5lBQVG9c/cxZvEuN+CC
Qe9rGYkZnMJoS662Pez7Ah/V4Gf83bF2RZOIECwkP2OfuZf/pL+xnDarKqa7nvxq1D8ZO9dxBbiB
/TF4PbEkWoyIWH3fqg0duf9Q82wTpPL4K0zXV50uf8ba8hlyZm3lviAkG3wXHlk/8YVK58HIaGH8
93cOMg6tJAD5t5QtbNgYlDtUzs+18xSunsrypglQnlhDuGI873+MYsRG7DDZa+5bhTEotVQiDiBH
QwnBlbMq1BtxvD0hX6axRqjO8vndpZU4JTarSG9qGik9b/5LHaifMzz+a6mhadNfZOt8I2qUuiLH
qjpyAT9Wg++RnP5v68RELUGN7TQF/F0DGfZY4CExaA/j4X4HTCLi0cJiG9J9ajwzZtjXkv2rQ36t
ZnnqmuhMCJ1+b9r7PiasJ7zOb42xlOK51njrzasu9gaIkZaN0EcbYrS17/rlTrQ8zjOK1BrZ3WK/
/vmcSFN+L/AlTZ+IGjDZ7MVAnWIoiHjXXtfWXzUBICbyn5W3C+dsYP0EA+oTl1MoRuY+cwyzneWT
erSGBVXBV4KAg3c7vJvQA3TN84dkpevqmoQcUvFrjr4lz0+ydVhxPc2WsOVVi8/CyvFrt90fO5rf
XkPZ03Yy7p0aPz+qR7RZt40CTEH9sRq1zy3bGouUctzLhabFnsBNrCtI16spA6+vVXnvlZDshQIc
u2Kzru/rVtN5wK0VjSiEsYZy6S/x3Z94GrmSptkHNPFWPW1wmmn0RMM6sWNdEHWZlaLoTK+R8OGk
hkXVsu3hR92fy2+LS1BbIaoRI0K58dqIT3C07Ls4SrhrVPERInTqiBzHXsDoXmWWvMOeBA+R1aQd
jU7iSulHNefy9L6H/jQIuyXgeFEuag5WzbCu7TkRKT4S7dJDP971N4nUAQQdhtx4CRZSvD+xyVzy
NZHiLV4modI0EBQTWqz2KuGLEMAmnLDHgnCbzrplGMr/2OTLLmsPsR7Vl2pJWtSdDR48iMh94UbV
N5V67RGNM3XXWu8zgBgWUPv9pbVG9aLnszPJlISnyfg8ALzWA5Y9sTK3BZslgyELUsofaEP9J2KS
Du2vDDJR7Z0EviOPFf73ymLSjlhI0DJPo7Jyi2z0ll2Q9nMOhSz3bJwJFtRLzqxhFLPbREcAQZjr
48Tb0TpT3+O8qKcNpkHjfxms2oVp4WqqCEEdvKjvYzTXxTwp2F5Od56oeTZfFQUVS+cm1LVpKoz9
g2iR4tRaRzKEizEyDpy7hqmXWhLOTYYrA9Fihf1TTFYmKfuyLQRW0wdZ5Lr3zRF428OWJu0du0oG
FcBd+kSVuaywb9nr8A92l+d4AY1Y8vKQZA+vigQh8GvidBSxSNrDrN6ibJ8uZCXYaoV7Za3dVsF6
peDqEkZuVD8iuRBMQVCQ+8HSWO89mMfI9vJjfZ8=
`protect end_protected
