-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vQ/oeuqh/8QPrIJeptEDnMuLHWfcikmGV3o8k+Uu1ekH+aDMk/ewzxhkmisAfHES
NcIss+MmWXwXlXTkYSOS1QuD5RoKD9GcDwcMW7QxrIKDIRkcyETsKAjidzwdFt+q
War6IN32Wy1SRAumDXQudTdBPKoGVRjXhOOvSUfPLTvLOj47kJKzxQ==
--pragma protect end_key_block
--pragma protect digest_block
5QyCZE4iibkSxh4CxeIWk+1QJMQ=
--pragma protect end_digest_block
--pragma protect data_block
bgSvNojQcvwvJOg27PL30I0vpfIcS19crBg6tj167/XvO2fzdo0tWoo1pApA5tyT
pa7CUuMkVO+Fz2Kch4k+h2TxoyzlfbCOBO4GHeTj2+R1jN33OAbqp9PP/FY8baee
SGQdxZaQ6Wjsiu7LOYepXxSeosha5MymfICiK1IuyXKi3sy8IK72feaqD6sVpMls
oT80dbgdpR+uWp+PG7HQjem1MUW/Kkcf486x2oSwMXPe4yeBsi1uwprwWa9AK41z
YfO70fRA5XY82H0PtDvkvlfKECzJdJXAp1yQG8q5NPvqBGh6Nje07x4x531OiUbW
2WQYuFSgTIzjJEAZMBeU6LLPsHzLkYor7R+s8y9s9gMfeCx7GPA7pAImOBm+0aSQ
vVGhHTTHQj7BwoKXR2QIaF/8/7+oKjQ+SqgM9I29Nbu9RtYEGX24SzkST5MQAXEA
x7oC8dpRVUn0N4VN5WJiOHzykOeCJe93RXU45+EK5KGNoTEXw8Gybsh3MHFf72uE
D/f9XJQVArzXv+g/RsjIK7F7+GKLGRb6J6hUzNScbC9dADKEHFJqr8ZiP4rC417R
xHs3kvvb1kmbQyICZjwRSL/fpFwEcJIjlH9D3B36gN9vrvyUvokslkhNoYn/RBia
5wLBTAqY4uVJsNQ9x2MZEfS/Kr3kaaGL87VAVWq3mdyTWO3nZdByD0pXmOTi81u0
GIypXYepLf7AZ+stuURiOmc0IUX9akMdNdIPtkiU6ymotqfc6zRGOWK6UoGQjGls
UhqgsE4/22QwdKUqc210IYJHGEbIWIjhsxoOjG+3zIi9BpdXlMVYMbRc75fAeUIO
pPiy2FXfKbc6dP3pA/dhT1LxCJbVm5ebQ/cklSPxvC7PYA4BFQTtIjr4Vr2Hw5g7
lxuVTZ4VQxIXuV4LzidorpmmGVuWM0QAPTBo7Yx6U6UuAc/vVaWQ0r6ETDQfCDkC
DjYn/gEMDQzmFEPT52Wg8Kh8hI8IS8cwcyeUs2x/xcBOsGZW5O4tCtZFp/KsCWkQ
R8FiKI2Ftk0uJOsbqVDTlSbqH6vLjSB+T0CKL8V46cC1y+F+OlkpHSrrPm8LJht1
AvoPE8sys/l1sRGnrhWq5+Q/JDHcBAg6wCJTEbDdEL23nwGEJDldnyRS26w+Gsqv
6WZn2iH6sXlFTym21WYefijN2ACB2cDh3VFfA6Ik7mNpXpDsceeA96wRBOEToxAw
9BiHUSz8TUSgTusIKVRO7RjtLZ71zOa1nk+ZTcJ/7PNwMhN1MthrOuTgwFtoXctd
hvjnBP9JHhzG0VG3X0X2eZ2TECmKM/E3vJzR6TbX3VbA7cN7hR9S2J/Ud5WQspDr
SgVI0wHg1UaD9fKm3i7pL/v9zUWDSrUbNrHZKjkBKtIszXWhZvsmemVBw6nCopMr
jAsUq4yqXtPn+3WOKYowyK1irIFokg5Q5xXP27nKxnSZvVeLYg6HOt3h2zAz/FD8
frjgChClfmY5yVgbBh7KYf5qwYj+K9lhx+zwzGbij2AV6vzHfgwRkgZ2FD1ExagY
y7ix+aDv97fWSRtDSPMUl4T8brANPFk3xRi7Hq+HqCdgTAlCEjoBkjEaNWjcbYxF
YlMepTBwjm7ejPujfWtd096A5GvO0wB42wR6Tcx3VmdgfVQwwdV96zWKdAfxB5HQ
PEb5rMhL+C1keKuPFxe1mFmhv+W7sqmdyomdPfKbU1/nqJyu4CjiyCETwzU02D50
1dbkS+m3e9sgdjC98SmAikrSSjlwL1onLMS888GhtCq3kXUETwlUF7vQJPuGIeGw
EoSPgw7kYcGz823rUnQ/L5/lt2gXLrLyS+BED+wQaksL2UDgtjZLYyW6XII7ZuST
0fsyby1dbgtk+C+IegVpiz4OWSHaRi401gN5d1tRcgMoRLqbRCuG4XwvaoY1f+o4
DNblPbuf3uV1MRh8hxWpRS8Rtl2qvvzv242N79HQvM0YYbvUNlyAYG7P/rCndOmY
65p0bpfJJY4xZgoBDNF60x9i/AgmagHwedMF5ioBcFQA9H+WGAlaH8C2+GxN+3Wc
cfpScK+l44oJjDcs2FM51EF9Lntx4N3xqH+CKSlpGTASnxLijjTro6nmeLk+oe5D
kwJ5hlJjRtEj6sAF9hc4LaqkuMAchlJKapnUjzzknLmNczNxzgqHS8nqgdCZu2Ff
9AdAujLx8dEobAPznW/ylV53QzP36rkkX9piXkyWlpq9yq/r+unNP1Zepk+RDinM
SPPLVzUKTC3jVvOjDvfWm1Vtr1TO+knCNp3sILqOkL11PyWqisxFMmHZJ55dE9up
b5FkXaKyube2iS6fkRkl1zdNHjo7D8Rc7mpZCsDRdiBu0suzutc0yy0h+F4kVzzN
1QFM43QCPw07EoudbGzl7JKVxSugusaclJNLbJfWifhvRHpAKJZqEV6k9DhRQpOD
5CE4r3T3pasRZGq2qtGkjwA7lnCtFteDZ9zgYiHTiIqrHOw8oIdCDIngg+x27kK4
gEhTZIr0EX7wLntTDhb+Et/ncltPYzn6qYHg1uXMHRzLdBRzu9U56DWh1CyMJGBo
rNPxVgSL4sNicUvxIPAy9YQbuqdouoh9D/Zi70hqsf1LS79kEJZxQIBYLFaFejg3
loHwc4KqqRg7NfKlg2qIrWQMOGMKg87aOCTuWweFCwmzLFWOJonCyFk+DcpMrGPi
rChAep6s+H/VWeWfDiLuyNRXfx1NMczvS5mdTb/cACeJs4aE5QnvBO34Qc3bsM5y
uHNzv7lKvUa4UwUW1g8CoYSJaLkxhuOYn1S4gKdEKaVb06YvH3ipFy3jDz3180MG
1Xv1AA8QD4on3mJDTW0EkqWGcOoMJu90QodT+ClnmKHPJrW4oYd47MrKbz73cdoM
4iiif4RHiiGxLE6jU9FdMrWBCXT2gWmGz8W/8FeDPyE5kIxiPscof2S2P75lJ2lk
ExbMq83SI2zZ0ut9tR7Fr2adqoJULyCXwEec8bFkfxQ8iO+y7LS46YkXNv3+o/eX
6C+QUymb4Zw1FhPQCw+NOxA4TeTSnZQI71l9xOR8q+XQnBNnUHqzGq9AIjK8dMa7
usQtAhmqTL5/gXei6WtX+G96Ldk8wGnk6S2FKZvZoeldC60FnfUzU+FfN97gNGtp
2rU5A47bq3XC7LEA9HKNwyGG6sI0Sn1a/s3xpy2o5NWWCAgwEFElGmOBhqRRjx4Z
8w1E0w+96uagNuB/VB7+WX5VxTYUpgdUN8zAoJv9m3+Z5kEa4BKxHg3wX+zGkd0w
juZMXVfJP3KydN8M3o2sN0FejcyHiPA303oGvSdWxSbEC97gloz8T1I6PqsdGkjA
j/1RBW1thjUaIT0UgpG7LMvBQLqDJW5feal05rW2/EeNSay4VjJygL+GQqyTh7jz
U9F2GI0WSLUv57cEcDo3BGJQxWB2WyvXAJsUOgDEpnMhFUMT+fop/cQ/FOgHTf8j
AYb0Dsf/Y4WWZERIOyc5wu8Gqpw+f39rnLXjCSftSOTYj1afXu9EUGtGdx19oQDS
nDDf6TpvlpB4YmAmW340vnj0SvNv4xWrhSH9w1KWsFDKsEu2qP8RCNrz9PqqWcbn
w1QLdykmvJZaBhqoO5UnMP98Q8qq6099zC28N5UpPq+XW+Wb547YuldMKoKBJUo1
J9touSMWAhJNS3pws4Cr7oSxfRj/6PTfaFyAim20IxqDI9gFPPmvfbGmZiF5JFWU
E/ubiyNOF8x6h/ZIDLAd5GeBerz5A1CLYsyKALAxcgrB0gEgn1UjZkTS7cNOaH4H
KNFHl373s3uOdaGdU+/Lu0mr7qOzxlYGq1EyOvzQFpOxtK2kQZSozTy0WLMdNEkL
jv08j876sjIW/QdSmAR8+cpZF2/uivl2ivv2WTPOf4a1308Muqdu0GDDFzmoCgv1
6w3tO7aAGaR3XDjoSZPvrtmTkBdofDgiqQttty3RPeY1M4ICPjR4ZY1iN4Abztgi
TRgaatxps6hvlsdV0j8oWj0cEG5ufhou9fXgyfUWFMO3ejJ9kdV9gO9yv8BD5YAb
qQLe4NpQkZHHeE14J0zZa4qtIv5fy0b9y0+fqrkzU31nBJJ8On7VfHqVwM/oGyxv
KIkU67LW7bVd+W9EQ16qwrZDC57EU/FTsgxtp8OiYOEBB/HiWGGER76nh2sZFfSI
QWY+vNHsRqZzXOinEwam/u26ujwCZnbE8FtIXvN+khTHOC2ej9R5Ol60TGs6UYCM
I8wRXrf3uRsPUrM+JkSLKNWotqSHgI2vtdPZkbZDqzABoNMS9tuD76ACi3nZEltN
MZ61aWVR9RFJeVVZhyfm29SKg27TrqFCWZF4N5Uha5AP7Gx8V2jcwxDkbuHicD+g
manu51Idd8/7DBtwdfKp4x4rCtSnk7ZZskWuiPRs3J2BgBI5yw08H0dksXFXqcLy
89GBHHPWSuiolAlaLfLjYy3uHykNHnj3e8Jc4B/JcYgiQJ9RjLQQi2/fH8HEbGKX
3wU/SXJw6pfwOUdOKpLn/xoqj45fQa83TC1lMbLvGP2NVJxqIAz+1ajIYe+CnuO/
yaCYIq61Eb3vdMHY1hFfthvz1Cqb3fBqlZBnHVXuclPb4pUY1uJRxZex+aLJXBhM
ppcjtU5Y+PrrlNG5PPhpj5foGKfTS8KoLNHRk+RgSrpOlU7wJtf2/mwhHnCKcl6f
B8L4OHtLY6NTTBebLSWuX3sUQJLsmxO0LzsFssvPZhToGHLCUomQOsdJYQYzVIHR
HlOCcxlavcna4eya2pt99YlvyJY9Wc6LuBbzJnsqZ+1qda49HkI0me4aMXK8PSr5
yw+tUOvtTCrz3/0FiF7oBiAXe3eFyXOh+2Ki7su5llko6n13INl1idFDOGw+KAGA
OdNjzTGXpJf/s/g+0cSyxQiPTdmUQgip+i5i9o50Eng8lMakL33xdTXxWSevuSJ+
zXU7XViMwHG75evNrRb57EhAkMWNyklm23ZCVyO9PlWjj02aP6yGYr+UDTfeAC1P
YFs+jWINFuGSZ0xs5sF46p0ascdQrjT4YU2jQziutvv1bLNidjK98JCtfL05UDjW
bG9TLtnFL0t/VOuw9y57hOMjmn8C0LG/y6Grx0wxW24FQPLWWa4GQkMwAHnKSdzI
CR1Mx8VyyV0B84QMX47qqj19zBSU2tbduEESbzRtF3fr1oMavS70VFyx6UvPvWvU
SEpb+7PcZz0bVnCngmjikockAX2NL6pzK4xSiW9bdDwxuWGLgr2UoK6+hkaq1EeZ
b9VyAhdFWkI4Raw6RsXkMTD9kHK7cfX7PTGk7/9vMXMn2vR8NFisW+ljogTx0IK6
7fK9RKteRjviSGZU0niHiClZ4oXBZsxsQpC6ztDL0AhvMs4/0rxXDwqDAqOux7SH
Ug2+kNCG4VZ9IUWYQ4VgOuUT8jW2tWuITizo0iFfOS4KKhrCgW9eYVyYuiweCuc1
itrVves2GC9X3IcOtyYnp776pS3mwHght9/QhgmVAjJ677VxaOAnQ1u6CcsSanrI
YsZHI6WUk+i0sBxsHWhkvYkk6HP+0uk3RvRKowBXDw6dupGwDz67fuyuk1W/DATA
U3yvKKn2hgQjDyEKqohoKYRS1W8IVUL64V3jce7NLT/uWCnfva0dcnToD0TvmD3e
lxSM+Lojj1UTHgKHHGxNr9Vrg9AH+8MIZRFW5AgFzVimf41i9aOjGIzgpk3IZgK8
7nz6N4HycszWyAa0VxjNIERqACTJpHU4D7342vXlmtCwMaLB/SnzaLFp6t/3rrVe
xdmsF+xLItjO8lpjtrvaUmYSYeF3QSXuladz9IFjDFWmD3vyEqi/mCrWgaf00zVa
3F2BMbJ5Mzn6g9KG1YZlD68YQ/gvNsXTSOm/Kmq/HtfRWDN7vnCGGPQh09d19bFa
Ojr4O0QGovrQlugyqkU94Um1osmoRV28pBTjVSnND1ZwSIDx8ahdmt1P1uu3wzvT
x0qdxV6eFdVFUSUM2MspSiSN76qHZYSJfr5fCaoKbBaDqMrDU8/+5/c2eUhZAEHP
DhpKt10qC5SV5Ac4gJpqbmTu0vymSbGP9egR8C25z8eDEYDhns3fsmyQd/Wndoj0
lWjj+0zRwqCPfIAF6nawtA6Nn0hDaBVFVFNG8Bp9EFol7t99aoacQefIRr2xOJtw
3VPGOo3K8x1BD8LY4Y7DrSB+Za2srDKfWVjuu1g5ggCniUZDzpEMMkDDTFhzgG93
beI3Syj+NRf42bfkocn6sb/gPd2DY32cexCqzcZSw7nokN6IDVUDyGjPuYq+f6Sc
eVKfSk0wpdljQlROq4o5yluw7ITbhiO70MKIDSdv4HxVaIdFMQPpIaSD51sUoP79
esWxeYkSuythIExANOLMkecenWjY5STMygZ4xU0I5COsP2bMFtZUqf3OjjwjyD6g
XZlYxK6HvNeiv1niTlD96Ef+SHOIVv/1JPEYyEhIkyE5GEf89YIuVMKoT/npjCPm
tXDbefORgAYDfBVQsQd1k29p6AIV7PMy33wicvBAGCqmXJk5HbwSZ3iaONK6+Vbc
NNnVgXhhzW4Yo24pS1Jkj608mXz0Mrd6TybDBlKSLFc4l36IZ7vCqx0sAhP7hCqp
dkNqGRoelRhybgz4POKXlHfiKJ+Clnqg2co+c1CkKqU60TzPxU6fmfl+2t31zxu2
dYYlnmGwZuGt8S2WOMeShO10A8pfxkrPm6cg1HBb8x1LgosYCcd3zcbQlAp2E61X
dorlmF14h7g9vBC07k+oHph27gYFQPUpw53S0xd3AFZ2EX6QSC6RumRXXrXmroYS
v0PphwKZ/eh6P4YeLvgVEeEr9C86zPIC94NlL/2L88T+Tk8y4g2LD3MxtIp3QYvc
n1BX9Uhz0iXKkO2W8YwEi50hxomYyX2mUYAKwzMdEf28MKYJ6i8a/mdDmbD1neYE
BZ62fOae6DQpPptPPMywS5+1kG1DlQO8irPRaZFJTdrunDFwrB6M7NwkpCskYhHo
PARtrieu5EXtBsrmXL0an8PzaoUu+Kd4Jh+GnRl2rovBNhUqhND6vlR+i6fk5BgJ
yHJb0V0r2XZEISnCsyCtdes4yhpjavaJpWlcsbUleHFa29t5k7nCPCEC3BHMZ3/F
Fc586DntI5AxWnk1z4cQx5tT4pwU5LwW6EEZqsQBVcC65JzyIcONPo0e/FFwa2eV
GNU6C1UUNeUDLWHkYBRMo0thF1BzbJpbZsa/TbgE3m/OA58dTrJ+Y6q1JYD8Qtwb
AmjjrcaG6DbvbH1XJuxJHJZz6gkMYOPx9KJ/nUjayyrUZHPehXpqBzEIOBOCf6oQ
dQDNAol95pRx2QMIcxe5PmYmzql7mzcy7JpH7//mnDLJWO9Q1Gu6fAviCjpZas8d
K8dMZineXcHOArf0ouezy97WDiUQSNGCpWTOWsWh7CWlb3axH79O8VAVcGlqJuok
zpgHAvUSMQRGjk3kCe6jKag3XGM9/KxNnTjKwpnPH+4G1MzuIGjA3Lomyud7PuyH
5FERSwkbLKGuq8PwKoA4WalPOT+051l77uNrFIPLeP0+z0F1qTFpMOkK7+GAshqH
4OPRHYEWyiUrYU/nYjWQBzNFWvX/phxf8WtgtarsnmyN7DhZo1W5exx8449jh7eh
LUpCWS7HNRRAVxeMgq2Vk1BytKPW9sf1/WWDRk7tnU9Vyb94XxZngo3/K21EzMiC
ZWzkbWUOhYOuufpSQL9TqvAOsSN9xoQqtd+IAY7jXabf5NCmOqjj3lIrYWtFCvJP
ke/kKZYrkbgVYyrT3p4cO2smjyPz6DMszfwQCfTf2HfmGYj8aihbp4gpeHKwHZuA
fpaiFW8pu5kh3X+zEuKi5gvumgXY9LStaPIicGeDq+8dxmH7NbbFWYynw3VGXevV
gfNOmy4lnYVz19bm1Fq7fUu+z0NSXZiDv2TGGyvxbm3pZtq6sq8hPJcb0QNO5oMd
8YBFWPUWnjAUgUZjmRhQEKXhP+D8cMKQ7mWZPWTkN/5wbgnPR3HB9kuif9L9T8I2
FEUObDaCJQzM5tJ40cUvRavpKyob0/RhyAD2SPjvuF5Lz9LQrv0AId4lRb5Vywu6
+emV7CPltSBW0DLcEqBCRs5OgISp+UUGd2BL/RRHfLaCwaRD6eg3iU3WL3fLBkvE
1gpVymA+17gpIcAYBrIMDnpGnnwfPbk/d2hahD4aKOAWLvd1kDZ3q1zVLu+hlnv7
s/wCzWAyKZLMDGnSYBru3KksfJ/P/V15IRqdU4jFl90tv04OMi9aRt0sKybx2qOH
ZCAMHno5X+734pKC6y3Wnd6EM3fm3ojUjpDhw20A6gXM89q+2/t6ElbQ36Wm/Wf2
qZBjA9bjQwa8Y/3f5DjFbYBr9zvWGlHBlOjnrDeKTOO2CGlymlj91W0UWInNef2c
TDMln4UZbDKmuGzD2zJkx6c0QI60j7Olsr2Vr0syZ67AkMmra9GgeLy7ImHUVhkK
+wIDoi1Pyv5qQTjFDdeYAfd5Va+cKexdyb0fR4Zed8z+FfBKbOmUbZNtheRs40o2
YdPcOJVaWZC1Z+/SPdHQ+HlRfUAOFcdgjopF8UInWFjRTqFic50QplLft45qvj/P
Ssm/xpYOnjbDZnVDf5S/XSPwP0jheGa3/2reHLR2e4PrmmocrpXNXNp5pRWuWveg
wvxrROjQtq6W9QyccO+spB/qge0KKLVAacOfp2hiXo1jFJy5xG7tFVkwOzi02S6u
jszYwXsMgA6v3KgVA4M1xgRXh61MSSSmWfcOVfXBEPaZX+Z3vs2ciSez02l5AhFP
YqSgOTAdpaz4sJLqMhXotmlU7vPPN33dcsXoLaLZ0ZP5/Q+z5kqEaJlcT382ZFER
aEDO4i9QeRnU5kbhOBr4OogQnpK1XEAiNLTKlLGX2N/vgD4rCMbEkk3MD6KfgyE3
+Zselbv3RDXTaaTzIy9IPviXao9GlZAc5+u1loGfIIv5YHYf5xoLEGagWlIkow4Q
EzRqAP1Y8szskQK98daMrH4XqX/od/Pjq7Xz2OaDIR6++hxuBZdIOwxKVMejAwAi
KfMLOx5Cea9FvaK0o7IdpR6TV0NZHM2ZalksyA3Ssld5Sbr5Iziw0j2YWcpsMVuC
9VdI/K5gud6JGEqmEUQ9fl9Sgt7I92Rb5OZQVchuC/ucyr37NxFOUZrN4N6pnJdb
JmBkN3SCVgmNbOYhTxX3VUwkA9JbIfIfbzI8DmWZ1qJWcWA7/4WntJ1tE7BRSRys
ZTUrRpG1rRS0RNjWCLanjZ27TLt71LjvEekJPre7ThMksfDOi1PveFvkBpoOD8qM
fgHYPsegnfud/RmzZyrOm3mOvIuxgS1x4UG3bfxNNRKRnw0ax3eCCkqyGBwWnWev
Wiu2D3M/rKHHKdvQdWbedKmwP7ZLRXYrYuPUAOZF1FiULRq2DVXzDd/EffMcBYBA
uacWllBb3Z+ktS0itpOXeycmUWC2YneMJqOtFdkQgkjbS0Ihx2G4dk05kR+5KSXl
eweGfhBMjvLdcnBoIq7PyQ==
--pragma protect end_data_block
--pragma protect digest_block
9LESHjBxx9sSLr7i3JyyNkkFUu0=
--pragma protect end_digest_block
--pragma protect end_protected
