-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
DilCODeyDkT3wmRU+VEgmbizyT3Lo3gS+wGqZOAyxEuwY2x7Sqy19uXVztVyf7Wi
0HlGZUeLP/wMMRWHqvDF5Mkt9P0e540kH17kUYl+wWYQcTqsEUjkG1LujaE8X0zP
CwRDocew6WVFmqXsh5iSERWXMEHzCaz7QHHb9wM3XkpNTDPZeFljuw==
--pragma protect end_key_block
--pragma protect digest_block
TH5W56vaRtfESOp9imO6kHyg4cM=
--pragma protect end_digest_block
--pragma protect data_block
5M4lro0CqisKH3rBI4BXXNxZHd6FKzMWElEooOaxRt14VJs822skTC5pm+XRJqS4
UlydL3JlghB9GPURJdZwVLkGNX1K2eFmVgRy3FI6eAGqhuQNwki/lG9avaR9FNS5
WXi0Qx63SkfLmq1oH6g0BEvAeLuxNnOeaHMDEafzu6QN3EbhmIcg2lkvmYpJzVMg
1JF8/d77ehLQWj+eKYnPCRKz69aU0kYlG70s7mlb3Uwdw8yeal70T+RCzEIt2oJa
9IzP2+EeKLLJISIwEeM7a4PqSe8W3skGEsYrDa5VfX4/gCmOGqtkGqWywH1NLzim
pp5wnRI/dGMvjwGFPMr+PCDnAIBnhAV4/yX2vukbqn8Z2Bx+c1fPi+D+ComvRZVR
44Bj2nzclvM4JzVpYqH1RSj/e7F5tewb7DY2VP/uKf2v4R/NQ0kMPCKdhb5W3pBt
16E8juR8fP6F+3gV0JqrdwhaBXemjJsTNLJi0k72muPOSGwjxPH1PH694uQRWMm8
ESE5b0OkKhhiHA3ocmvhoI622JVyJMudLhpUGCZ1op/Mm/VczJYb/b4QpxEjmG2R
a3iTJQdRkFcwdw1Z1JCEJwJj4cDRCUXhAiDBDnHjQC07wbGvy1BlufJ+JPUzkHdb
Kyf7NyAg3eFsHzf1Jmo3bCxsPtfdfe0M915kTxR+ju4unigoibKj94tZCN6znJuE
f9eLDIoCpp6M5CkgKVr1l9njhUmqfhTb+iBjTuzjAQ7DGbctwZLwyXKvR7XgBEoD
WOHaQH/qSLKHkOLibK3WbQZFcAsPNepDT4lm+JMxMciZ0J2GX5dFbrKrQCWuKN5r
uQoSM4aoEIGfu5rZLWsP+412475OmdgTjbbn7Ntgagw35SpN8XO2SsjAyfyVncG1
5cXML3Xu4Pw31Zv48VPvB+y3bs+FkukMDdGAs3O0ldREpcpDJJvteotUqyt6t2H2
BljzTEWxOT7zjlxn/D0RNP8htUsLSUSlwHR8PJT83lVbQoAbOvgVipTeSf18ULJ8
y9aQHCBuAhNaMNL1jTaZxL6XFqYtfW5xysKo4vSrvxNpRXaePw45inv73aFNjSaS
Ie5uGSeP5iI3d7lfW2+A58qXd7oJ9DC+17gxYLjpDDTLyiD6siBF04+MEVHNJR8w
AAO8mKv/YP2oCNNIuXJyvArI/MQoTzlMY77zbd3I5ycSEWW0y37B8iWhIR7ClwSJ
LorTUwZa4wDPST/HGMtog++J40aRDrS6wx3D1fZLf2xhEHvy1BYlyzgN83vDyfom
OhWK7H1rgC4QlsyeYks3HtvcFSwpotijWvFonQhH6BrQnhI8he8CV8ZHLY2iaiaS
BJgHMOTgp+zvOMXsoR2/bIBbw0pcSjIxR72qa4lWRUDbNXQcfdHExgd/7OqoPcbk
8kqbSSLDKgoL50AqWqppRRE9+07JyBX1Z1UFij2b6o6d/qQdMj2V2rprSjSjb37r
U23oxHBYC+jaoLg1dWSuCVKcQ4ZqBBeFDgQduZcks8GCK0hWDaNSU6dax7r1E9ez
ZaRnqiTOKYwqntV+Tdw9sHrkOr9d5b0C7iim6QR0BOHA59awtsqLCrK6PteQt/Pv
9kU7ytiTU1IeJcgLE9Vk2gTkSL2Jtvj4UHBFHfC8JsF/1ovz2/rfCNd6xlwrZEct
rvWU+zVdEFo4WqAtbnR3kfw3Y62YXMTFFX/G7RXoEM/4qaBjJpFwRNOcYK+Ul+2b
/JUIo2SqXQNW1LUiyzXx6ZMuJBDELZpII6J39Bt6OXXEzGI5XuJ8IGwNCpYRw5ep
lu+DFNaGglPTU0/OvDupH4HWsQZqCaeh+qiY4JiiTTt/HNpohmidh0/BR/KIM7za
v0FvGuMF1J6bWZQW7ExftBKk3yA98dXfecqxT8M55WifWNH5o20WXUQ1hdR2JQUr
KVBwSE4+k1eYCF+B8rcNIjxREqc7/l/SkxNTBOGbQHG7Lb36eXu/0M+mdANJmUtH
TteFH9VBTb9q8TH1QUCsC8SkMySDxJ7VWNjJbZXJaVq+64KjNAvyjwn6RXmTar/v
DqWN6b+QKFp+jCF16S4SnnImWyF7cEDpXaINTAphPldi2pQfo26pE4LHwTcNa1jG
VOqfHddWHEr7H5RBAwjdM5ynG0Pm9Zl+nhMDontMV9Oo028ve1tENE4feIq24tES
az+H+niEHaE/e9slVJLFw2q1HX+DwvCJ7V10AfiVilDApV2PI917lEaqJoH0r1iG
jkTIoVplnqjafQG+n4xyP5WkaPvYwK8HBxB/hG4bRLnXmgVVAh42hcImwqWfgJnl
akDvXi5WjvPbG77phaCa3s2z/OpJg0zGTWerPPihKCsPbGOIxhkAuUVMCp5TD8ug
JVR/SrP6+cIWx1S3FyB1Ap5w3wqPeA7MTs5K+npZyoL0Rsr9ekzQoFBEYlCjSPZG
7StpDuC2Qcn9OSSADr6t+xZeoCVNmeyVBQqZ1JiplU5YMrKqpYEwQmmOReXsl7xV
kW8ur1RTUQ3nAqgmsx5XG1Cw7PTSMzG5AYwxSydBMtM+tF4cY+zh5s0qjusCbY9r
YCD37lQUkLtgBu6CEQneRcyXA2t8/Jy1s8uBRSZrPyD4fuP0bRX7MO8mySykDggQ
iTXD4r1IB3LgkIEpNoAu8Y4eH+g3Uq8q2hCHHpa3vd8N4hwuD9/VbsKHHf2vx27H
rUJEo99PLWgU6BRFERh1044q/Cld6Zn4Btl+lQ96wmQrGAAl72V1ZWK7k+Nvwxza
/bfyLN4xpB/iBt7hVp/8w10CAmag0DdGgc+pZc+Hfz9J7Mjgc/ftI5i3dbDj6rW0
UdmeEIqKet0Nlz2yD/orx5iIqGhtqcI+sv2+u7QXeFcTnWWt9D6OZecICQe5BpKV
0WNXGfkgp7Ghkgdpb1hT5Numfd93whUDRX+Zqg1QX13+2ud+PG0NJTlExpxZAvcG
X8YSkrZqkQwi3wEb6/pmMB3IJ7IbXTSZiFZBkeXYgrqtYZIyFk7mGUDhFrv0BUpG
td2JhfanLo7tVzxmgzyhDvHjbGoPEvEnN+Gbgk0ykNFzG7Cb3mJOtRUvEcGvhEDk
Oh3PJYmrH+lXC9h6Ln0rTI0aE2afbH2rh8sq71jWqXz4l7RXfGXr4h6xUPVmkB5x
QZQPasGxJioWV4yuRJU3g5Q1ZlZQ/XPlhtS6VuLX4aRWiO/kUGUmoTh2RmdlJsYZ
000Wd7hfJ5JvrCWCSme3+pd4TjVKVx4akCqf+zwJQCaEJAEMqlxHEBGHrVeGN2QD
llEHB9nEEBWCF1kxujqMBjgrNp55n0w+L67jwdnBQFcoIVfqOv20wBiejZREC5Pr
Ppyloq0VoJxEWdsFfsypSeHpNsytqEUrj65WcKRQO8OUx1XvWjpRKqkmUv0HcDgR
P4/YXBd4glTcS+jTePoPEGaSULHxxZM993NbhuXts7SFHbjU1LEYEJVcWsvfAtfD
BFpIiF+kgvqifJ5s0tryqj9UAOsC/JuqpN44ZRPMvAPypLw2wYwcK60EqfQeUBs9
T92HDxT5/HkQIucDEN/Z7+gtDZq9HA7EbAjr7zpuf1MaqWLpxon77dePJoBBfDHe
zqSOAR0JSGHCTXpRR7lZDOz8qxs7KzDtnVzN+EppH116+aEPsqTWW7QKMRN5rsSV
VYLBnzS8yjIK3nfwEPJsR5QWIdbp7PeIfkt+m80fcZGbMRuk3yr14Nqw4EwGBzmc
2UzcO9KCPmM5/0h7hEYwd3jyEHBEaXSQf2+Ia02gqBsGkOUk4I7RwNH8yKrghXua
ltW10gCKGkoD2FxaSzjApRFqPx4SxXfDofTj2s6jAwKF0EQS/0AhX8ldHt2f36JB
QBO7gLTC/04yWga3MeW+AhtxTV+xEOHIIWUzbrAdyPoFaV4nZpqr23tqzsqoZBs3
14alw3wHlvS037bD7H+Oz5ETEeJegYORJQYKG1mScFR84AB6IMZVeD2f+sgSxIv6
nl/GnMMg1mWOcr+Wd9itUZZ2XqGhIFjV8PwjAP3DWezVHbUXbDki/BR/mWjPzKVx
pBR6HNJBZSihmYOS0yS2/P1EZTOzvimGWrhd/7FUu5QSm2/5UOxpHeiyziYaHHG+
dyBtVYhYYy26qlXRUdNwQvUfYWbzsIIqNW5jxVS4qeOkKVRTd2Qwmh7/YpvY3PH3
cTtKBQUzx/bW9DZ0yC3VV88VjyFAE1wgyxSmDqvbbWx/q7vALZkMdbQs2tjd3npL
fOIT/nAw+zIL2qWSLU0BYvzyGoVw76WQOp/PJ3+8qI13DPkXyOejV0kOJeB8q47R
jlaT89lRU53xNjaBQey/u44c99PCSz9vi9DKlmpIxBblsNzDNklOHqAPWwvzNXPT
Q+jKDFKkGJrNDyqafuKJrt5aodTv/B46CD8y40g4Ndbxr/70I3PHXk70oVAT6c6F
KP0HKTrB872fTB4bVviZzHwoR8r1CS+pBJ7Z9zpZmmLn57ciGJNOy/95+a2BTy6V
GDDziwFv7Pbv4FdPr+RgnasuPT0Qq7nVU3HJRHZhSm6jqOP9yZV93/tJZoLoqWII
hl01AC6ZDGhOEpn96hvGZ/OAJ1XUwSiSBpzWH0SIie9tM9ZEffnev1NE7OTF37rz
b56qJmIY0DEIZ5NFvdpcm+ZvD/m0kv+qszTEO7Mh3d47JPwiB6DIoAR4Ifb00K0l
djfyhdAGOh+Sc9oHWBoiXGjtIB5jLF2Z8LkaxaxSCx0H5PFFOTlGmEo3LcUaD9tw
GdNC8YCmOsD5BpI/OkVLKfEXHnmnC8vWE9aYMmwkNIvU4xm3bqADRExpz+i8Y6hN
iN0Pz8Xp6qEID1TSEsPDdDPYWmochrtgIe5fRQz8yF+gohpgoANhN+EBTpGcw+fF
aOhdcrrpFOMC/fuFFfSDMPZLVa+/rdT27qZunlN7cj1qdb7AGePPlB40uND3P0Z9
os6X+SXaReu3PLcaovCiFffOZktiDMLo6iDQu6t9FDKa2+9Be43jlInxZYaLO7ez
2zoSftacC541+jUuYqs6PwZjVm0jtqO+3zRDw+l81QrDk6hfXQojFaFGRkdh6Gzp
ZAd6bqMp8FTnG4JqZn2rx6o3KyOLc4aPYjjiTCQNJkT7k3X5Je6xjpeATQwF5n4l
d/D7658ql8xLC5uW3GOjXxmbfT7jhosdSyjclHg6YbwbA8SLY3gw4hjOXlm8MZRB
1kS3PvLw0HJ8jlKU6DiKoav5AN7hveeoKafDRVRZzxsNN+/CZlFiVvkz001+vFJU
9taRtyKt/1Nbr8Q+Bs52OaGkLbXjh/BbVtSF49abuU3CafVaE6cIFqxr/xaXDNSf
fHh5GWJ1GpP2NOp1cs/7t8JSV8aIjhsja2UtuL4ILQI1Q32wn8/62FX9y3m8L9cD
CSZuo4sHfYuZ9immjKtnPypi+SsiF5SkTTNDqBA66gVCzjeDo7nYxglXXjtjCtf/
RrkZPWpPHIZyzCyulkkZhCf/XpHqb3Iwf0WHK7MZM/wgoNDajWEakhG9mZ9npmZu
YOf8HSSustiazIGnCiT5yhKt6m7F89MaDFhayZoyvNMh18Jw5v6R9vwXoHleMnrL
npvwS1MDSO7aHanudyWVPdI7PtOJQGf+kNGkXSzaWdSXtk6wtZYeShSjY8o6Adok
ZRpwFomVriP1EXkdwnAPt9IgJsk9BDul2LHwXZa4Xk8M6tG0EAquSUp422wc2XSV
DOayjt6DnRbjObCBiN36baxuLDouDLROedzf4HwWnJie1rFVvSc7DQ7s/779Q3A9
w6BPDGy/JUnPekAIP8PrRTNBma87wvMMFPPNSaFRGaKKn4J+JbWOtM7cMa3l9PgY
Ey49jaSogb6pSa7Dq83juMQSxg1FJja43n2H4x0DOVcPVYwuAapEGy4FKBWJZkfQ
QhFd/KNIyiHOh+7HzDEsBDjxJ+Js5i9/74PeOhHE2/0JOrnaoounv1LuvAbqix51
J1rCK2I5Hgn3m9vcWO01o2HmMk9y/GHJJjyOCe7OSf05emCOELRsLlGdalxiMZZ1
bCpTdwohlbzYzuPwUdxc/TEMZZv0L4fMFtzYq6eqBN6m+duHdQrujLq6ViBwgVgw
krWi5d7oOkA2oMRGgsG8vLY+4iaUImDOCf7+kX3IvQgb+xLxl4gNoTDGe0SFuFnC
2xNxQI2Y7yws/x505TRi4BqhZdqyI0UJaXuvTaALi+nfJ8po+NQdYzkljV/od4UR
pgV0sOQznKCxuh8JeA/h8bZgndYJ/Ve51RBdRKf87YP5IrVaM4hKrSjWkGFi2BHk
gNaOwhzHqhjzXmsF9tpHHpKjEhr9INcazhL6VJ0tzjBMbqks4BcB3SiY+Vf8vYfb
SjKSgbkvBccqBGczxdzhiQzIeb0KBr61bg73ey2fDEyUbCBR+wjUNCToDzXfkoUK
Wr1d22j0MqTn3LZ+Mjnl/h1xJRzpqkxsJecKMw3ziWPSbtfm2QoydZSa+7v0+cUr
zdY7bl6uKvedjmLZuCH/OKOGlyl1Faxt4qikiWYef6mR/ksrQKszzM8MFfh3dCDK
msBNG1AYz7ZmjPRz40BxwG/+hA6yfDhdZ1kcrf8mlAfMR3Igk8joPq2+gSmFZ/nw
dPPP/1FuCusf5YsH/1pGfP+8B5YmbVIPyk+toeW6o4s7x0kxu8morglgo1/2WciH
KhnN/wn1ZoYxudN0saUh8/7kcAcGCvAovcA6rXOKq3k0ar4WYr0Qan2fcU8emMVp
d06nOjbd+e/h0EVn5raH7AoI40igmWVH+vnMXstje4JIxTZXDHvZJHvaoiVjWU/Q
mW0c3m2yNQLmnUZompAjvVeBcQeru0VXTyHNJ1PdkRv4atxLwjrkc3Mpx3ahx+nJ
quLw6XfmNyJmm/RYnUBjZrwOo8lqf0RNkOlT5bde8St7CcgUoyJqfv1Fe5cna+gm
e5nYJZhEdhLW9wPim/cumFP9XikCghBTMvFs/lvavYAmimzXKz1pTfM77r/lgYVe
ngpahFLbkiDBWvMyFbJ7gfrowr/fS9TXLYmFOH2fbRYeX8r+KYQI7dOA23pkejN/
LMmynBhoKcB3wf2AuOMf/1fFFRGawrMSFH4OY7uuyMudAA9EV6mRyPwZvbLzXTmr
aa6+tmgzN18a+GWYqOUcctXbsazf67XmFdNz2giNFBrfNV8s1LJbwkbo7wf7AtU4
+2GyEvn88U6egfF9rpD3mg==
--pragma protect end_data_block
--pragma protect digest_block
/IRlrveZgxaUnjllojwJganF/kA=
--pragma protect end_digest_block
--pragma protect end_protected
