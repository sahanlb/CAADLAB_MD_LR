-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
FGMI03RYGM4+aXQgu2rD6puQg9xZrDDI3iIBwDbfNg5WLAUF3Y3DNygnRKzytXPZ
8U25pMGa7mvuSwYKg65TEdClFX2qshaIwpGoOKQysks3yguV3A49T/p5xwZtriQP
m40OLc2rdJ4yuWCkSFEbpW64aVJAi9s9IWQGhgFtzqg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5175)

`protect DATA_BLOCK
1dr8CpyV75w0Ov+mjOqy+P4U3HAWpt4drGwLSwIWaL+1fZfA5aMNU/aBysOSFRzF
zdTOEwdP32VHD00d7SoGUMzifHUdxqRcAbSb2ygBlUjkek5mA2JOYmqBcsx8WTyG
V+E008wiPKiMis0PUo0WDbhHTYmrSJs83tosjNT5hYw6RTdg8v6CDOv3VpfOO9Fb
rWjxr5Wm512Bu2FYYo8C0gmdzi9nonZeX3ZEwEKrlNBI0L9N6Vk5Eq3myaYWiZBL
cpghdH/rbRmrqcdKTdMmrDZL/V6dx+DCQA7M/CiJNheZ76/x6XrcI/5h8Dr2X63y
+Q0cjKl7OikIZkJOc3XPjYxl++fbaXDTvcCUQbC4zW56KB0zrTI8r44tX+1nmai2
IjvbCET5Qkqrqg7bLT9Ag6vUo8ZcxwmbahuA2IvWJ5WFfygwbCnNoSuuL0SFU21i
2QdDop2+x1t36A3Tx32yYavrngskRj7leyrwIr7/mdbG11qVBuh/TCFz6yFq0yWc
2AYBLWMQTQ7Rr3vcTse1hVX8ud54eh0MfqOy+Zu+6OGyO/upylewC5KmKvdvyI5w
z9skEgMpv30TxHCcXB8teXckVrQrNcxnjK1QHfg4b0yPLY733U8WfBbMjexjfpNW
hWFC7ND51BdukGjwQZujQpoir8eSwj16tAeZGZVeqFYYaGcYYXd8Bt3K+iXFHkx4
i3ib9qt0JQXMxmAN6jacMaPerQhxrmidolqlOp0gOndz6RBOo+e1cJLxc8L2rtoI
jcxoZUkS3p//5c0uVmTYqEIrztvBmm86bSphI8h0yuGGKTZss4Lmgxt8zKG0hX0Y
HhaQJUstTY/u2LIdMCsA9O75wWMNp0B5moS9Xeitl8aEzELqmYnt+Sjk/5+vtzt2
gnJTCoqPs3DkRVh9hT3ww09wNQYBVHg20htgudpGFhUR2LSI719H3PQTtjOMIpxp
6m4fokfk2A/SQdF7qmL/CoxSpXnaiK0caGQe+xwg44M2enUXDJQ/Wl/+Vpon2zvV
CGw+zwXTM0YmN+P4UoZh7rHS5Mrsa+PPWBaVbzXSaxQwPUNeRFX0Exph7u0aZpqA
iaT6s0Ggf7wOYUHhSrgSgsy51J/emAql7QQ0A1xYf0IEwjxOFAb4atUJxEQYN//u
v6hTaZ6y3NGn6DWLRnZwHCPPj1sUKW5oZAGMRRVOvBO0KBEU2jm82TUyR28An6kB
8ECHDqpV3sDhAuEuH70xeeaJtxndy7hEaxwElaBhIosb34PeZVTrddmS3451sEpN
KxgUalZN7sJfFXn5vx/4IiPALN3rVZQvumpV1qS1gbk6wUZFft4zdqpNo+IC2Yuo
o8LHvxwI9wHJ+6t7gH3pFmPJZne+5+QabfALJu4g4y801VOoFBnyhDEYg019oHEo
yysqpss1y6T/ZamGvtKdJjdFqDJVLcMi8ZEfl0H+iwHnz8QyYHcPt3/TjBbbBYh9
Caan0m4y24r5zdhHMmJgiqsLXFlh9+KTqk11a3Z565O6CPU6ej/IuWE/WJDop3mg
She87m8OVZEB2Jx406gqKAV1mDMGK9kuLh0jDaQhg7R7Xd6Yz9GJv11iLZIo0Kh5
V0chwW+98fJ7XLnCiOzmLFnyuBLEeAWaI4ECsfl7NSAOT06o+BNXsmhw6Vl8Symf
/LswTx6HJfsI3sWRzhooKQc+duNYzm41Potn69o26cz8C5MmNMmSequcikL2JEv7
8ipi/qE+VLMz1j3r0mz3Njqxd5wxb+EFkZsv/2TDWgPCZAuiWeofEhIcHOXuv+mO
msdU626iDQSXYVEyK5rankjFugVOI3I0HUYHusHBMsnUZjys2Yta3xjG9rMMPd/O
NDz6Xa992sqos4p4451JhnclGDcWCVA2VOQNgc4UwMv+7GAa6U/Gz0cRPAzeSD7/
MIG41+eDRwofKjcrE6EwM8lMy5uePFImn/man1zhonLyRENzSiOKTnPsucZqQpw2
Z+vvEYj5rUFv1pVkLnzCijjKNZQ/9h10yzhpW4haJyICzEjOdyh+H9WEZkjJqLjP
WykjCnMt1iIIDRHJuhMWbpxyLB4E+5ZBDbMl1x2HbH+ZgwPxP6FqaHXBjCN3oL9q
TRKgTRSYZzmC2F9aPXxMbGsS41hckw0ibyE3ZPJluq2PIyHxlYoPMybxV8xyUZUT
YMI24/hxJLlTJDBmtM9r+40pzX3/60BS6GOPP+qOfQl7+ulG3Uu0H5wvDNpIHDXS
AH1nPN+u9uHNZqIvt/0WY5FbCJi9JYz9rvpFKJeTy9AnyJTk3A1AIEsD0RDXW0HU
A1LVSdlRg6KbOh9LBRl66eIB2MeVcg64h1AJ4EYeJk+OsQzclJtv/77syHzcjzVY
WMDYvkokTjPLOKp5waaCpPsrDxe19+M1xVh3wt+9HaX4O5fEs3F9YYkvE7r4LmIG
g1UGNaEabXpv5pV++X0I/44wpQ7S3hKHXcU2TJzPvJ0zTiuG8yaFoMFdmWQJQoFf
OVZt8oxNeERHPjIbED5HNf6j30dcxnMaHY81h/NCFkUNVa53z1Muh3Tj8DzyEGI4
yp9lpcHBC86eF3OBOp0qyF5ZHH6crJLBH5BxYaf4yQpIALv2fmMrt0FZuC3nyDjl
E0e0PEKua+jfhR5+QffA7MEuxOBe0Xe6WBuW6kvYUEqxdvrw7iSsyAVSPnk/vH1s
jz19nNU+mkPPZe589Q5uHMPEfkAm12qZDPk8QCJ5FUN6cXjTu7o0nqSygVk4R7vH
fofgYT7Toxdg67V7dm4IRe+D6sZUs1tYB2uwJBJDx0nvAY/5JcuiMCZ94Cc7qNtd
9aoKunMXhfirA32v0QLZCWoCCby1LOWIreKIB3t5bP78tk5X46ry7VfWxZ9frKwi
qLnB4dc5C3DdTNnGE2q0p+coKLGmUTBKX1MBbnePOnBX8i0tRCJmztyE1IKfPWIC
ZzZW+g/2l0DG8Vdogi0pcOUhoe6PoM8BJAA/VWielotJB1DmL3Drr44Oprpntl0P
KhEF1Zr/UZVcc8pLFmwr8SxmyzuhiMWjjnGPGZ62Su7v6pcFtAZzY+Sz5ZquNJDT
gn3tEDLMJU3/pXDCeIdTN4WwZCdm+C6agBiJxkGhQxjHNKJC9d5iCoqjZOURJoiB
nqdp2CQLseRJm3xCscgZMLubM5fs6I2Gc0CR7ZNbW0qz0Yc05jvntB4MMeEHY/sF
YeFb6QYYpxIEtqD6z/WU4kLtF2N8HJLE4LskXht/fN+T23R1SxUfCFIU4zxWPkc8
gkaiha4mECyVV6+Zpk5yEIvUeh11zgEbQoutTHKEJp+tvpb1lIFg8/98I4gomoWB
hIEbCIHH15hTMai8L1ujhYJdpxI2QqWAmKzvI+ZW+Ax+8Gd2BwWgr7FQF0Y+5iMf
YA0zvm3LrX/pw8eU3UQOabpt2Rn8mbNIx5Wd7xtYTa8CMJL5gbW5bhhL3bTBMRCS
2JzYa2RqWZ3LjCN9wUM4xe5oVakif/UHZFrr7NlL6lELDELxdOKf9/2ATuiEc3nV
7DRqtVQm04qenV33lHBaGgxKr+6sMwdeJnD++eImJqQWbH0D0QMt+23qRBEQqrck
hqJAZuwbWtNC4g77wnNtCygiFmEOED0chuGw4nUrXu0+XOXDc57qRghh3DW4vj/+
1WujHeu4t5A2mbNOpuuEOdpv4dHt/0GWO273EZNh47NySYg7gXJG8WRbmNBVnAlN
S/AJsrIFRfJ1WkSD+bKeqhTszlaXL8cO5gwcmHf0qS7zhFKZygbKBw1zmd/TXHtc
bZgDO3BmXNXxA3us9t3b4lxGBrUP9fpPuI3VW8ak6Qwr/2iGF4Yl5uVaFYg3cMc1
dDZFu0rgS/CHwHIsTl0+HaLRCkNnkNFY8Tb5ims6JYkcZLp+jZ2K2iO7+I5/fT3n
IzMP1QhRdPtkEtH/umMUJQX++/0fYF+bW7crEue8liioOSP/WBVs2i8tIEy9M/jb
cEnBFi0+lHjkRDVsowceeyWZFWibuVo3a0EUjt8KgnDz+aAa+qbL9IesKezqicpM
Mg/vyGVqmh8PbAmK1vM0Y67fKjjcXnpY7Cqao1i9cx8AXOAeVDUDLGHT1NOkqpsS
rqSSWQvNLyf4lfebJL9aP/h3o6xWniqdo7xp9Cjwk/nC2XlsoBMsWMzuoQL5L9fl
3HQQK1XE3qdpgf0rdYXelByRHJ/mm/hW5enXWEJyOl8NarWhFcZFYp0/MT6cfD7A
3qpc+DseJIeVv3TfdFo1PgaXiGuqOe9GgleKYzHMBBAH2DKJKHdIt8ZS7JwsKuus
dc2qm4VKyU9fYUOwmS9lFd3ExM2qUDyHW1r01ZBTQBGxg57L4HC3HphnlR2WMrHL
GuhRABnbd0OLqgvraqOElAWmVYTXXj4hGxRVxxF8ElpnsHF85gZcxWId1aYzxVHk
HxpeDVab3fsKggzDgE3IKpom+uIWTh0w0UlNgmPSfIE8xtIrpc2/NWWAep42S2SI
3qg0tkMeKQbQc7/XTLdYBwhVhGzol1XKjXcuWyUm9CopFi8Q8RRG/QenHHseXTWc
AiD/CCQnWSvqwCIhCS0dDZa1TTWEHYmeUpBeWsb+xNYTois29GRkHXdDXtg/cNFr
msjAYZZywpk9UEDOylbcHnZ3ZczNFPaIqdsYcp/4jLbaweHoi1i87UHuxWuo0C+N
w9q87uB7T5yAJ56kQhGcG6FtqmOoNCWGy4j0WjQ0i8M/pZtNKqeHdZdQUqjAdi9V
uzv9SfQm2XQZrChsKFembg6+f2wxaUlzo3q2Q97P1Z6TXbwfMPMSKGnv79u5hUNK
f9n5V59W9LJel/uEmRpVkYej/h+p3e2d+Xk88LgjshSqsoCDLUpd86ICiOwZn2t7
ABamKWs1V5tH8r1TQ1b00sHIQYiD3zJZOe3FIRAnzdn7UQdOJAh8HRREEw4WRKz4
xYIBmtsnvsLrlm7NNK67sGCyULn6kWP5Ck9wKpmiqz28ICNNOrkg/nOppxAV7AcC
B647NYhd+SN5I1Jo9hwi5gKXlIWoTeLB2QZmlApDSxx0oOgMZylVOSkyNdEE57ga
pRDS7NuP16Oh6HhRMrGrToP5AIdnOhSXRlahAUu2SEglDHwAwRnAvxdp5o1zWZgS
416NgSdsKOx73InvwqvqjoITYyRfVm65qX0gn6jTZ4khvRbvXStuNZOheI6QuF3X
hmBskGGqNmrnsEKAnUbeZjdL0BB5/xBzfunuMTMCntsVXGFbfUPoeffO11rRp92B
lp2f+sjB09KEDXVq9PE3KjwuYHM4ywk40uiheGABAJiZNZ+1pMkzYKDdloA3vIGy
eWHFhrA33ElyITlmRPcwCd58Ka/us9E63+a4PH9sK11X90qFuEMZ4JM+f9whrxR/
iPyidN8exquCnA7pxh8y4bYu1C9UzxjTSrYJU3SxXFYLom6/bK9bJvAs77Jd0UPl
9P6Z/EagybxeNK3haTcgYsPFhAqO0r1evlM14KREpN91nkHnkYHv96iJN3m0ETV5
J+VX+n0jOKgV05Okvrf3WtMQhJ5h/twduq1X5mo16147LOGPY+tfALYx6l7kd6SS
W4Bj/vW0AbCm7gzB9XE8aculyMB/uff2TzI+/7VA4km3iKPVetUcCrLHO0pbR7y4
NiEF9FJ1V6C3Dwd3TqVnfe3ePte0ibIfKgAZ1myMuNMTmRFh20Exl3wEEtZoPDeR
JgRYUctrVMzW8oqcxCOp7agd2UYJC4LVKH5dhNYGzO6gAckyUYEpj0zZoxtbmB6h
vqZRyT1N1TQhxF2KNdobTiGhD1iBFKlICXFAqGCcBNnVU7Sfdy045RxnGtznFEl2
S4+3VvugQS5Xhte/P0SjzQs/6dISmE6pNrEowVozKHp0vK26I7hpskCpITbZn0+y
QEZh6HfFalCgmcGONQXq9d7pSeVGaL/IeQLUb444PMmmU4MLVPy7B8DyzB0slCbh
f8sH3LkOQewG1WxfPOVOIkvbv9duo6+ebCPnlhpGrZYHyZsSIbgefElnTQABRsym
9dx1EBZPpgT/rO3KjsMJzS7SfEy733Lt9ri5tu58fR17wXd0d2RJSzPwtW4Odstp
H8WxR1nT+k9lL+w0WzrwPAyc6okW7ibSvAS/cL8P1M/XRgwfZdn7fuphoTNdoRdh
XSevoz6iIX1s6OXLofrhC1CGGtE0H443Ei/suVN7Wf59lmvvyMrBlPcaIYNNNZjA
wK3rMasRlGruGhfZfYiDNEg1pmSkzYPuyc+zvgV4O2g6hqT8GMkftR+ayW1/hHoR
irME2F5WZAo9VvDZLg6s6Gh77fhUSgwpd3RQmOWtXH6KD3rt6h7ZXdvudXBQcHnr
0oVTjQowDGjfxMfR+rMARcK0lsUvumUZXiiTGlaq2k2+KIPHK80qGONQZUJ3o2pR
JUsspl98HbwC28mEbSqc2s1rL3lJRq8z+zmh0S6SG7gzO/vTxrF/AEVTRZo+vkxg
CSec3ykuS1BibHds3nJ/NeC6J43ihZBE15SAQ1egbze1WPlRlJ2YDidDZyMBx9ap
rBzExSZrMawyarvCKhCRWVw81lwYZHl8w5wYRNzW3+Am9LI7xY9YwNtLGYIAhXQi
szTjDTYn2mFw24qbPu79joR+WlVZm7zR1NFEk+BW1mDSGCkBHvephWjL1ty7qOxb
qhHUjzVHwn77pHn9qEF7QNRnDWiZU29tc0/P4fFGG9oUU6S27e/tBSbhyw8CZcLG
k+OHnIK4+m8OXUK+6a3sj/Tl4mjpRIWJuAYJiJdTaqVylQl00v8fQctdoaP6B8Uc
6yxB5BsPYGL9UNL/OnsOmQoUEh0V4btytFn4HQGDlq+BvSkiTtSf6ubVLmILrP1t
wzpU0xlH4tLEYzVYJPS1qI4h3QSTwOADjGudJn4jx0HETSgPscoJyMJGCwDPnpeF
ZqElBsUgJLZLh084b+9+MQ==
`protect END_PROTECTED