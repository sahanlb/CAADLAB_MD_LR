-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
w4uGDTufmWHMAB+Fq6aH5eP7LrpubQfsrtOGpNb3sVOxm1JG/yWIDD5mSprQdkl+
r4mZJv1NtTMowCxPJqxY6tDibYAgZafQEmi0JsEl5csW0n3uX/bUn05k5tg1ovYQ
VOsaYVhye0OEzDI89OcXiBeDYid3rmvyYcNUtkZr/WE4IGUT/F3lWw==
--pragma protect end_key_block
--pragma protect digest_block
y4xneJUmktGTv24/1lSr06jfqXw=
--pragma protect end_digest_block
--pragma protect data_block
BxPo6MW2rSgokWtinOjO757hpW59qRKMd3Nt4ikINAfQUK8t5GGSjsR5LODry9ze
hhHbuKsMvPwd5qGfX6cAQvHasBw+FAvG6FT3Giib+qGwGjgVGIhYerjC5HeCC+Zk
I+ahRUTTxhvshf2j6XfZ+yuFaebrg0e/dlNrkIkl5BFA1F6JNC42GjApdGTnmlvi
M/ZxK7BhlcMzET4sr5UD0Bc3Lwe3Zdbih8IDJUo/8jOOpVjswEF9rBMKodi6d6WC
SOOkPcxLe91RrvtDfkkH73r8IYa7E7tjFFCRUHZOtgnZ+FV16g9Mp8krjOP5YF9/
s4LMts0f6F89vx41QqMbSKbaQy17FXuLwBDk2hWXrUQXYZPr9pLu+ojzXfuFBk/a
DdwkenD8+fTgFtbGsh04GP41/xGQZDpK6oNdGeq+PJYePXxyz75BATzf1VrarWPn
nf0yQYq9WEoOjVdDIwskHSaxZGLepLdfZRAlkVH55G3JHUJn7796mgpdaFlJHAsV
LJ5WW75vm8BMhMaeeR1yq4fA4jIPLc0lFD8x8S4nSjPoB0INTDoeyYHFatP95Ar0
+x1WzL7JOG+M9OIm3Jg+IQGXZLTXfFzDwDubgHrZUtPqU87t/N/pq9lvKVgpLvlY
FH9UfsLp298RXDXuKGrHllV+OUMLfEGznGnxts3nA8AwyUR22+3igUXRw3L6pVBv
soBwdbJ4QOig9j49Q82CUHJ8iDJPRi4BrzEd/7cYyVFp93aOVZalaGwyA2kaHLCN
eESYbxUVker5mqhlAvOdsJEeY7CDdN1kjq9WqrmKxtCa+wXU4GEuTTfB//qnmO3u
y3PXe8epkD8schkw7x3y9V052WKn9lhJD2pQ+0l6XQfK4I9/iiOgPFls66I5sGH8
FVgwcJcDFhke79FLm3Cf6TIjs2GZGAsWGLQz7sT40Gv5ajg9AdubBH3EY98ZnQNe
sfIsal7/+pohVVvtF470gAuJnvqPrTFJLxXJPQbkvPKVhqG8j0FddUaNSCkTCDsQ
4N2M+1lZ3tRy1w2Bv9PZfZB3LOWRyCg/isbFKkwydNNNXZUvhKIp9gxxUCy1oCgW
fhFc7SbMEPqKJ+FCTWtAABrAYfF8RyYqBWDgXCN3DGVYg2JfAynj+d1D1abEiu4t
G6WZ+JFTEWzAP3kFoRjb1+bf1KbpeV5O/XFEQd+9JO6psyHFPthnVmAwm2duHyOZ
G9ZjmYSUxLqKMINdZPwl98oDzRRjNktjUKecXNTdkXTYAIyvvj60lEkIrXzx4wO1
VDznSNzw+FzP3US/1kygjBDEpHSRFpTNZVw8YqGvSGXU2FlvVJZy56b3hP5qljeb
cOObxWveqOdi8ItYk91eHQz8gz1yqZtVcU+xkbEBzLMIk+TcYPN++rSEjOGA7egC
AKQjy7gxW6QqoUfeGOQXIzlhEYjNZDUnlpusf036VG/O3jCxqXyUrp5UoXseoBkk
UQbU8HjjOFkLEBFNUOwPkjsS93h2bJJxXf8w1wrdgppYlGLaWVwW2hJsvUeKyBwG
zUfWZZO3dTrkAbKyXQccL4gYsBeJkL0nn4bF2w5kJ8/9PK4R1cepGg6a2qzWh/V5
dEWe2+WmB3BpSPhDE/EEpE3HTQUrFCIixO1nKABI7hDsv+Lw/WAq2RF5kqrKvBOW
bYDoJfa7s9D5At5sgLMB+gJ6kWbCtjKQuQuSZj4NFdjsW2Za415rplKgLWxcr3zu
AQdTzahhHqDcvEpjZwIYkestVwvjhG+rZi68+UQlU6HHSe0ozkLZFq1XTlidU4PW
orLcxmTdCKIoSV0dXmAHjig96VDif3LFzjFlsgIx+ta1FNA+NMz+k8uPUUEn9ro6
S7GcnAIG8HS9rvZbAaK3P703N4Ae/O5KeZceCaM61NokdvPA4vti9tTmsRi1pr1M
3g+Ttmjb2Biizykpmln9nBpYWrpIGpoK/K15OIk3Yn+W8xOCAsMV+1R1WtoF1A63
cib9msrF5thsP6B7e5NCZKOt476C0h4YZ385pQsvFKiHDEl3J7jBbRsPWEZVtJXF
agNzGEhYBx6oOiQ3F97CtpPBjMjt89+w46UyBMZmaXYSqZ+dYkN9af3QlafItk1I
UZIM5zXoZXVYKWz1w/rZPOvDMnKmW9ywI03kAdrm4nqRRKtwb8uT3Y0U2O33D+aR
/sWLv5ClGfGIdTXHv2Edv1cOpH+Oitu+Qt3Ks+3YJYbTkkxdBOyF547HYkk3xhkG
pvrBYhh9e+kPVZ92cnAK2OjrpZlf1Zy1JgWuEXl7MjC/h2wletQc6lGmTpl0dThS
chz1cg2AzfHtLn1PaARnxlLqDH+4wxUr317dED9tw4dUchI6llMuCV4IipfINlmC
OQjFAxzFpAKmw5rN8VpBie53dgFeBMejWQf5Aosl4TPU3VmtLYG8jzk9bsfiYl1k
/f315cN6MOqFsRuJsbr3PfrFlhSTB+cRzccNvkCGCWzFVmRiIDEjv+UBY1mJI2OQ
7Xxy8Tln6MM1ZeoevK/SAETzYunX7QB9NToMIAePxwau95Ucq3jbPzIFnr4gpkNO
axCee9SLbjhLsp3ScA2gbrRwEwnV9HSGJmayxgxIAj8UnA5JzmQX3GfZrgYaAEJ1
e9J1eZ+nrkfq0MtQ61oLv0JVweBYD4Sb9fDeExwtHErkApxdupuyGYSeMZ9Mp+rH
M1E9/8fEKXDjosddndvcajA7x50YYUruyZ8/qTT6AfQvRC3ryJggpCV9j4UMvVUb
EOLHLSUl0JAEFZfBzH8V/OimCqkpsn2GA6uESB2dyjL2eSnHZYEmB/ZPQ9/d4xgT
dgv0r3fEpQZX+b62WQPbDqHE6805CjOe5GsPDQYLvNwY37xZtJOWQB+3KeMkSpJ5
asHNgmMHvTJwVXqfZHPL5RvDputnTVIBYiGtAiIGv1SrrQlPfPAVfJ8Q9aL3L8nz
vfBnodWoDgYgp8kSOyW617UiGqrYfl2J8o8Src5nmU9qXAhKmvYyP6wy9U81jin4
zyrlh172ptbNRKGpLBj6rL/97NJqUudslkkgl5wic/Y7HhAZ9paYe8Gmwqkf7wQd
/UmjVtJtI+YVKW3+hYAUwHaV/1x/CLujWrpLPpva3ghzbUmA08crHeXIQo6O+vXJ
Be4YpGAAHQTqXlW43Nzmye9/54zLkUX/9wmBiehlYRwbWeSjBZZOVLs+6xJar1uo
kT/ly+UYb3FTN+BKuQXIvhvSMvYvK7JQCRCXCgCFka7yIP7MqzXyv+K75zPX3hvM
INBx9Vr2laKjsUuN1TM6PXCSJoc6AhIdgG+EJb95bAixJ1lxzdR6SLNzzgtSKLiv
PAbvTdIgPpEiqVnTZ2Rk3gnZknm21dyRuhimgUE/MawPhYkysggoj4dp0dNpVcbh
VgeKzu0FxAEy5MBEE8pZdwW4zQtZPZ/zwbsGhNhzBXsY8VtKmPPdwP2ZcZAtUG/+
c2dlpttke1Q2ybEfeaeGxCrcycevXAPhd2Ijm4mJW/ITADF7RXyLhnoECKICid9C
TZVYiYHfsSf/0eWr92viZwnqdnWNvny7Rzvxy3HBbkr/krftnFlipMmgZt8l0W8X
4DGMPTpPgYBjV1juQup9l555FaVcPXraZcEc38vPTuRAqa3hQO2y+UnPs0dFb8eA
p0l111G2rlbCFbgami6/e6v9uCfAqBRcFJzB1uRP+0KO63p7yOcpcwF/Z0XmRZ1f
zuuChivORlZz6sMkYrTfdJrZ9BoJ/yDu7bz0E3PVhX41jV4JjXU4JpHNhp26FYQy
6HR1n2yCN+QTKe+18Hl95HgBOHcQtgaRC0DXueYP2hZZVU7n1pehewlrYKM7u1Cj
89WktBsb5eueGtbjqSIS8Ql88fSVex2eAT1gPS8Iw6lPJA1onZwzu7swWPiBw5LB
lmLku3rIv3TwZgboUoTUUF83jY4zjnOKdP9aBQVvlrWj9ITmOr0P87JGoRU9nDSS
mEnKWxI72PSPE9LpYWN99fPBtt7K/3GGcfYvwRZDoubg9hN0CfUBDVLpAWgiC1vo
f8kp5QspkgO4fb8mV7aIhQy9/jIc7P/DOGJmbnxJaK+bUnW9RfVjIA4o/RUjIbQV
6cZQEzV2MzKKJH421n3BqMPxiXryDKa9AemxXwh0IPZ/+EpTj/lrtgFubE1LNzwn
eK1uRl692AMeOuKnlvNeRiuTamwPTt82o9DJBJZwc9/pEAvyJCoBo94kbMMT29r2
duNHI8NMPlsuybiZS5+rVzPiv4CIEt1KZSUs2BtL51OWUN375OVk4/nyjqWa/C57
JtvfHEDaQmmmH+3uHHRiLn/V3e08X7adVliO8rWazFjH2uRoihB71vW+RETYKZHy
dfSjvIVnEfMWpxSthtsdWdSdYC4zqeYphJreZewmm6yN9mPYRKezQsTHegbBEzqv
CnJgI2k+pblZ9hZyT1EZxsI1EImQajBCvImudfxPaPJOtMp1pXUMWKm7k0kuYMYB
zlg7yFQ2nnKvJkKEngAx1KF/ynHeLJGkklZeDY8MGJqMdov0u9FeJhechYanR/9z
KQO9yag8YHlE3Zs7L3ewbprsQulhXfNwIBiZMhdk0wRjlTbaiDcuuBK6tRNxPD2B
D1CV/Tqk2hd6gUVEtMR/76OpcExw90Y7GS0Qdj9xyFy4xJxyALEQHK+HnjEPYECJ
zVRwjGDua/cFdcxgyHnTwmNbxiogRiM6RkazwjaBWWMGo2zZgW3cgmZ78Rxi9zE3
bLbRANElIy7g/Dtb54BBD+W4WKqT8n0q79xwX6dIeg1Dtgei+IDiLIs7UBy8KLgl
vXgf6ng45rtqXF/T9FHD5vbKGuEVF6vGs8PmZOreieW/X+/MzaIeXKbYFlH9z6Z8
lEw7fUA76zOI7KJ+0qvtdsNgyvUJCo0cLbA72xMz/hmQufDUdDhefrcj9yRmg8Iw
5SIQ/R1uA41M6GOSSICf//hUZFTZG2IBaWGsUjH9Vu5VvAMGHVuC4cJo96HQtRjn
R/mQIK3GbyE5BObHA6eq92uib0KO3XosfOYkj2UkRsvkoSzCtXSd7BoEx2TN4ptm
XJWpe5Dl+uU8Bqa9A3I3+zaMCAkwmxvFcmir0+afWaXk2sHSrhRslxkobV5Xv/nt
D6d4QL/fysDGhqYrfYDUi24VQocrIqV3QwCY/ewMWp0udfAcQom0O6yZmJilUEan
xmS3vOwIrHeNGFiS3AupiAG965wLV6INjbwPNMAvPA34OryeaHcssJCiUHI1tEkp
EkUMhXE7woSf1U1gTjJUoX0KkCqHC1F3ZxUVlD+j6uf/RVeSpoT7SpAU+lP3I3zY
lB+ByyXSfsMmz7R6lcdWs4xopWa09mo1O3YAXFx5Ud5mEXoHZKOtqyo4R0KLIlvp
h18AxZMgjUEL4BCtcNbewvJ2v6r0yIgPUvCK8eXyZosF54NXLQhtS1/fM8XoCwVJ
4xEI/OCM998Nzl/fkfV0QQBHTVvl3/DrMWRyW17yyFifn6EZr1jpBMiw0KmTxLgv
pWAD9fP1jMELo6RRi3ZOFDGfsEcqSfawKe2sANgL1uMty067ulBgHEjIuSht+Afl
ALYfF6yrMPlhfIqsA6u/n50fgE6aL0GdNjEkobqmTDRlq1L4GCbb6fRo13JsEWMW
TtKmfUjJdyFztElC/UYRa39ahPfkM/vcBdbK09jSpaq/+UBQcvitjSwXdhIqUQOr
6fL8GmqxH8IRXZ6rQ8jpIO1D9Uf5B/urzkLMhBzgbvnNaJxwFrrWKBvMF7U02OUs
W4PLw0cI87TtZxPAV7hzvcSb9qE7h/3y5/jMzidTGekiVsqpkBsCCaZjzxBtYW3E
+UbkOQm6LkkQCr0yMQe4cmJssuUUuQhH+t5TeY6cYKcUwqYcC9+Ht7+0BDJ4MjFj
nDGbXP4Q8j8ehl+C5YiAA2eMYGrhlymVs47kRDdUMbMTHn7/HksOT2xGZAcSeef3
4WR4kEk3vDGQ+vM7pMEu/x75rBKKKKak/zsN8HUSNP2dAL78ZsNhr3pjMx9cToan

--pragma protect end_data_block
--pragma protect digest_block
VUmMlrwn1LEotoUtanhbt7Tz37Q=
--pragma protect end_digest_block
--pragma protect end_protected
