-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
SaJLFQM1yPQp2g1ylqX8WCDbQIHkVRW9v3gAyXOYhP7n9+6M7HT/C4WqIAcGS05/
zrInrfoudy/lPEvWRgbO+R5j6QI1WEMmzdfN0nmywBGMuQK1xClLve8qrE7zVBL7
6mjkLMTEuJ5mWoA3N9ElglDmSBn56uBOW0FwBaaHsmw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 81696)
`protect data_block
AbrDt2VFHspCEAwZnukO9GiraVrdBuRf+vGK+TGYuVa8BaThoDRvb7LP23/D5v3O
o9mt9jJXUF8Vxak900loyGC4FbU/kxuYGLI0VfQQzmZ3/cABCZM4YHsDqRF8mr5X
0yj+Utencd0dkS30nC4pBjmtNls6jSVaPfYadenK/TwQprndqQOTIOTcE0TwnBML
lY/afBCaV2X2yVVG0uTVZyizAwIeBPdkqONG/ooo+OSDajJid70bDHXucGy2fWa3
EYQQIsofpvPHjRdWXBbdFhWt7vsJMbWJqd+MvPi6UrdBYsxXJYiPdF3x4ZhrNC0c
bA6Fbc/OAuQ5ZsFnsxwwJSX3mndZpHNbfDUc8gHQmo03cnS7A7T4zeZRjmqlxtqB
ysKCklD/ZASR+1UHwQS3rTn/38fIxdRuCBKVuXqgfZZCYXodJzcMyHC3JfTr+2Y8
agCpZjGuFGHhpKGyeShraW1lpLj434tvu4mBf8VO9i0WrGGSxBSYS7X5RaYuecIG
xCai2zlt+rSdRZ0gex+VcSzx7dWlxd8dZ1250ZfMWSRG4pMCoaSgdCthcltZAmRo
o6YEMyDDlYSpHQV0POFg/4frqa3zn4e+FuBvRt5gIra8s5YocQdsSELT9PLIZnjX
zQFeJgG5Cy7JOtkQ9Y/9299ouDc2scKcDEqMyjQlFOduEW0ezcEf7z1Hrt306kqT
I8SOl3Zv2X28aGKMDpUUnCt9Pi+tp9Zz4aLbI8coIiThzyEzLDokZTvBQIdkS5Jy
eIafonQkcPbBCax73QeOrPMLtyEf/Ayl4Wz9Zztwe0MKcVBbfQO6PW/Vt2rb74kY
sB1OICINe5Gheh/wi4gAVK8vNDmQxQuiGNIGH4nOrgSuAAETpbyGcYRCix8MGX2N
K8IrOx7hoWGksbDFTp6gOXGaOaNuipDfZ+wIEKqR4bRJp1NlY1FjJe3r1/50GdRV
Wsi6CJwt5bFHEbX2FRYnz3Pw0bImYPCo8w0FCcu20j91LlUA1wVP31pwz6r/7e6L
qqgvAXLU16dJeJWfTq/Qqb8DSLtmu+cWYIq9RkfcjnFPfIX2dbEdu23h5ILwpDpw
65IpmloLjJWuPQ/I/UU+aQ2rbRKxe3ugxOUmJUou7xct81G79B3voiBIduFlksll
n4jNwU2Bj8cfvVz6nZQWbkd6vOXrymYe/CA4zpM7O9L88DyKvfHflr/02l+cZ3Eg
D9TCGEbR6291sD1VAHqQ6FHyYo+PRiq4iDCsio1SexARJTaphB+SMrYKh1Li01lr
SKbCqNY8Z4hEHeNwkqlX0FmnlzB1DoQNmr86qLxGnrZ3Lm42FGkwQ/D+WBth9z8z
3q9YeppGMQs2DSnZxrVFWKdaPAwMKz3wiRSA1XerX9eb6SZE8QKSfI0NmslAiYdX
R5YaKpKZtNYOQRHgU5F/3xm8zuAgpwK49lLvWwZdSV1p0IFRsJk5qC1hTGu6dONO
4fDY8WzQGsywHEWPwsdgYcTW+UTDH1+u2IXYXSIK7IL9YXkmR5OgFkwpw2OkOrY0
HhT9xwvzSiVif1ToYhVhzFjgQo3rBPtxO18FtnC0u9NM5d6ll4lRPBbdlbMc5Snz
4ORuwDdHf9FHBbrsJxOgK3zJ7YiG0wUMKPP+6MqTCAkmk7F03aspoBQ7V6WorkQ0
wM0EaSyRy594GGoqi/hRn6i/QkzQajGedwxpgiwPxKnEWlI3fN2FTYM/57u9oFHb
WLKuadtjXyVOKFkV6cTGl/KJd5kipn0st3Ik63bt3peqNFkNVEGQLzk+upZg0gK9
RPNYzoazjPqyQZVvwZWlX4oFfPQUPy7fO0PX+aMAUg0YHUCk76ANqoOAyFURPWJh
2coiNq5zI43p+asyTB3KmElKK7P+WoafNZPBeCRBRDtVTe6A/JkYt4D32LfAFQnw
iCZCqPC4yqJiUAF+ZH3S80yTsdycKl01aBKVhNGS3BFh/N/Z7uK9rXYS1rx/5L4k
h1pEIWOR71gzx5x7SGslJBXDki3UcgzUMPLw3K418CVhmg5mFZ04thzHQVz8YmxP
As1yJM9E53/NraLQ5SgBMZcsRSQ5pY9jWFPu5pd/fVZ4TcpE8QvtJq8F4W/3iloq
5Ez09Sk5SqtesCCYHpSMrCXchdc//bxH+Usrr63e+LY4DK/I5xY/9kMNs/idD3jK
YJwSY9EfXe253kOHS/dfIIn83WPKKWPiiWZ4fyZQ3XnjWaggOpocEx/HsQfHGDx4
/WpnKqf9zUnSPSi65UahlL7Onn9WdmCOYZaoJAEGT+4ScvMGpqM/U9dqGuqdETpn
1lBLEb4wpQt5sna2WI0WGJTWEXxk/XDc5qiWQeg3Twxv4rP3f3MQoPHnC2cfsiv2
dwmiZM8kU6QXAEWheILz30rW11CHkqHBbnEjeXelR3YSLu36DyZeca5d3vPyweoY
TAdqtqWqjsUNe8Vl0VxJMNECxuMI6HAMUw/0+FNNYOBayFSYH91sLTFRj6ObFMxm
rr3usKnPQSfe9Va1VkSNbRx5e87BUVh2E8ZTEWZZDsg+OI/bQC63yTeiFPQiw4OA
/ygeCd73uv9wxAHHkaXCb9zFZyhfgoxt61TtXFgRBk6cBvlVtpVAFhrTnRqpl+ub
+mB68KTdq/cu6aFo4CvXwAJSOpTl+otw62EyxbCAogFUQ4oq9XuhIk/fNCXKnxrR
Sh6ZWHgckP7OuUzLDyVu8ZPNaEWZIovKlCaVwi+KOgQtsIM2KZE/6jsJ1obKyLwK
FPpRv10R5R+dK0FEpN1EeaEJyX6A/YZ1LuvdhVMnA59OeGeVUQwnrE70ied5uqKq
YDDgEf6TowsABC9arpKzfORSqauRzfIh//zZOw82h2rRU3zJwZAklgaXqd3yIFef
R4bl4OWmKdUIjn8cNyIqYtTGOxVcmcENnfHiiqwW89CF58swcvyWFdag9H8GwLWR
oN+9aSVZTm9jkfblqSURSjCyUTY+M4gSNAqX4jccU/S9/GTW/eeoi6asKud00/iG
OY8RQzHYxMTqu4/n33XheRwSyG5Q3OX/6fwFXYNesmTwPUda3O+l7TatdE8mpG3M
o2HbfdLuR2Rzl0Dm0Hu5V+3Al8yRAzkeR4XlP1JU7zrifCSC1mDP9qVDIp89KkII
gKPGAuVeUh1ibb8IATmUqR/WoysXWUxS3PwI0glnazTH3bvMegaic2GcWndkd+Q4
ZCHWrTctK9S//EsHJ5qSYb0sIOrlgkW1WGubMWxN/sT0M7THKqmyqls0ID42BRVU
gM3WCb6WKUAsBWs1m2QbT0LwggBi32F4fRT0RHi171KsGVhQATklmphQTcSBD4J/
pqA9drdkAI3m73rkpYZXbVzH/ZuOkqIFPRP2CvxaBab8el1qrCvYKrRetaUwDo5v
r3xH6hmLFZhvmEhSX9/p8LwxuOW9F7o8bjqS0iN39MQ0w4+IoUgzaHRoSVJTMiCy
+rLGsymi8uKNuop9X38triZY/mAUOUVkVMLc+z0URD9mKDbp8boYY4f65QYg4+fq
qx53DQFqacDAyeV8w+ytVJaABeSIi+eVdRRrfHUJBe0+X1u1HGCbfC5qySVYlHLU
IVJLdx+KcV0tTuPeMFf2Cm2uu83o68M4MKdC1rPL0Sijl/G5hlL9P1DAErkALc/4
3ueTQqlbFw2rWAvovQCWeSXQJvBWTLwY+C8QfQ8Xcc4LatL5ZCEV9rzpDUYieOnS
d07qU4HbEtswpm5BmGl5/y4gYQxgqJkkJVhcici+2z04wlhbhNefQOo4hhK9I59n
Yo1yX7o3wSHYX/oZixY57eHbC7xiMFOQ73aH6j177rt0eub51isGguQ290iL7DKy
+Nc08mgwrBtSIo+oXI66TPsAe2Y5k4jfr0li4Yd8zxzJ2iYCglkB5/+W1N7yRzT+
8AfEMlwf/Eiq0y9Q+8ESwh9i9ssMKG0ALjiFuzK4Mt8YiABHdeE3A46B1uYDS0PC
SpTOEzCPcy2TuoYQh9OJAXluLzsDafrslitHe86FOjhz/Kamfns74gkz+dAICfUY
pVnNGCYz5Sp1T5ZkUuBEjwJGwPmGlnsbxS3ysepSX3aP2+5a3HacvrCcEtnsJ8ph
x1EUcLtd2lNmkPpNBNgcILt1nzLJOPHRN1WiWemWgwl5ZUWC9MJPVL+VzBKj0yRe
2braEt46OSxX33l3Cml/qHW+jwibKB9GHae336TmazotzBJyjnfgSDuX1T8i2Ysj
hJ3iwkEFuWIBNyQCPPkFA+9YZkS4+HACISus4nR3KtiaI+TOarS+W4tLbAbUVvSJ
UpKWosdLE81qv0EwudhyhDbikgtcw6x1eiwGyGdSOUkqhGNQExG51LvCHY4MIsJU
O6Qv6/T0JBYAgL8k94mvcgV2TJDwjlVBEI794smKegSrQ8q78N6DoyU/fxImEYYv
rempgOmD2xWQPxNecKbhInI8TDd4rwaacvU7D0LT8MW7WvTSX97xTuT1ZX0vXtid
x71MTxZQ53AHAk4oVWKvve87+BbHzwKXOpUxZjacEx53FEtg9lMY0GeC4P3DJur7
lTO908aGUxnsuSLyAmS+2qjvbtnEvBnycqzTGL0ZlTJ9QcNTurjjWM8/LjnVhg+m
dm4Dp2wA2YGziKamcQOmcWQF7MjXppG9FgDXoUMB2TAAkm3AKvTY0BtqZT9lgisG
b1qhaludj+OtObYcSNE9GoTTPaJHMc7JwwyHT5yonAvqSC4MBibAXu+DCXFmY2ek
h339s2BzXsGBygRntqb9K3EzBCwCFu1H6HvDSwxJQu89t6havICL0DT+tCCLJmq9
/Oc8mY4KD9yHWgl/xVyBwkjdRx3+1BKW5drVOQ/H2yaMecerwLb/yvagdLqT5pn5
xSCjEdbRiJ3WcWQMMKb99B2L9RW4/qSbMCEm74HAMUD4rrGPzO57jV2GBVBo/Ux1
pu6Bb0CVnpwvXJoQBrsQnGCFsBc4yKb3Ge9gPK686HlJ69CdpqabR7GyRcp0OO4Y
om280Puc0zvgkcqDgXCIkTF/M+P5bo/zZCHy8dy/qt/vebVDB3n8ogluW6Ta/apF
04MDhfzc95Ae39dafQzUNRZpuxkWkGHcAV5/Y+qOa5tlP5ubqvKseaJsqmIVXw0Q
4UzHYV8oExX9o2NIJXw79aGbA3/yVl3sVYnN8hmqzXNIxqS+EmL2i77CA5PLmpW/
Veajav76XWv35S+4xzIh+Q8fUOf6XGyulKnQwwmCcQ4wXvxAial526HRFPUw0V20
CcMWnjiS2j5kZvQqEWD6kIzwFZRSNaOqTBA1QgtTr6JVAGUYfuhZ//lkWeY3Zz4W
uvoGDppglWeof0ddC8QZsuTbuXmIvQ37eCggFFuEFoupAgnqAFzIJsjvgpBWBna7
JG9xkM/hbMUJcwzNdjQcBRbS27BO8zv6TuUJyHFu1TDjFspmuDE4LmGMMWdZYjZC
nCoyOYwa0AoFtph2Ycxop7/goh4l7z2p3UhXIHBsvqjNqUj9dja+szZ+LLwalO0m
+FK9nquq5swBum0z0br1nhK7YHrLryl6X8HgLGvYParRH+Jl8G66z/1zo5rJfyjF
WI4W/23UoAdG+8/mpYZd4VJm5NOrCUJTq1DuLF1FOwd7Y5bjcE1ymMXoqqqLg1SU
P6Z59rcYExlxtKvnCax/gB6DDJpbX9q8fYLXrmbMFoHaMSMffnwjxILqUjXuN4ms
QnDB8BcT1p5pzJmHphC6AvUdiH+S6hHmJQqfTF2UXyeZELhUMvozoCApW+W6Rd/l
p1fOKDZHMkrucJC/XN57lrXXghOY0rZ5s65SwqeDLHPhHcxOzdwVpofzU+BpEwdD
8zN5FCCg2tu+6ghQGwmILu09QyKR64By7RRnJMy3H7cQ4o74qk8ZaZCDwGBYh7lb
TPrSWyXcKa95XrfrdgSAeFBQGMWM17XP4dnctjViG4V97rOcNjxlMk7KJny1Xq87
LPMzgYJ0sSHSdIUwykHRXqu4UkndyvJZKyMP6q9iuhRK4ydMklPj+NGMKYN+7/ly
A60kWSINKHXj3ElCXGKkUUhzDbfbv9nZCaw2Jkaob3Pfoaf2gibl0Uo0ImS9Nnhf
TIcif+DnudgQn8D1DhzFLTM7A0FF510iIVdQQ16JfJ8m/7vFFqZ6OAZStb29zGjq
Iw5n3QolXycIJUvH1lP1jLOGUdpLjY1b7PSCJn8oSl3Q6Bd8hKJ2FdfqHcSqQzCh
5VjD6XWV2QqHcn9mgmuXh3CzJFTcgupcsQYkFD2jlWv9YjFHYcGg/U3OeOrySmVW
i8M3yQpLd8M57pNm9ZqfoCZ8eGz6f6yfJvDrew2iz5YmYnBjOwAWv/Pe38sgMaGQ
1JLLdpMjppMl+OwV2owos6dFOTt0OFK4qNiPtyAtpKJsQ5yc7DpSE5pDb2WReQMJ
fE/i3xXgbd2lb/Blcwbbp/KELVv7mEbXkyoJrtnWW5YX4x8QX71BoBjX+D6SO+QQ
l4GtCfKi3UudJZTBrV4bVNRoZuPdiAjXf6jtRPPTuoErKs8MEMBSGaY8rc1BWBjp
7ET8IXBeuofgkorMNnNY+L9CHtp+gA8vHXI+ePZXUr4/X2c9P2jXYfNut4VoiOZ1
VBVjO5JYs2vFr4sazuCS236hFuTARGFGUmblAGtC9wlQPLVVnZJW9MU0DLOJFTxq
rCacRymaqeScLsKP0zh/skaiSeI+fpSyDYJqTJsgfSVFic+eZY1PfiLig1Gl6zft
cmke4knTQS+NtLlvY86YUYFjLAsVqsPg2FoCOqlpK+Sn5QWzeI1jfjc0Bj9vx47q
0bDm/0LF0XCZcghTE6RgWqDZ8pp/IvWVXHTFXuK01JcmRWyzPqaJ/Tk4wFtut/z+
Tjxk2+ezi95SQRx4OhLUm7cOKOUWwmFRJdt0UMpn+fd40RkV5dmPZlFmhCMMUU1/
hR7fvO/YwVqATWjsC/HHEmRIAgedg2jhI5gOYbElyH08Xf4DgeLEqlf8LfLpwpyK
4MuljXe1/xSr8+Wgl+6zt0sWTw0iLbGMDCnX1RFOS/k+V/Zg1GXFrBincrAC46Qh
JzoC5iRpokWmhtAI+Un5SB3QPffZVHubXd3YzQiGLqZiUE/mLusLuwdchwA9MLRE
I+ZjYM6u2N3ppyK6grHHaHvxp+qSaRQ3WNfz56Rf67Uy3bF1wnjNOFQmIbgfSCjq
1FrG3d7B1hXSMhH5Q1ybG2VkBgiDJyld77npGXxwgLklBxctXnJqxCZC3I4b36BG
ft9JIeWuD2IL+RGxsntZzY0qJwZu3/il4hQ3geoyekxJGmXJBm3Q6AvKfT6BrrIU
JQ35IxwKMgyaTsJFU/FbOZEEpAGqsKwTgn57akGgETzJgxClohio771WkuhZNLbx
Sl1MyUrmXjwH5UMvwJY3U3qYqZxk0d+JKreJ1yjMB63hf3RQ0SXp6rqk2aWRSi53
71ZXwCdQ6wMPApUYfbjFKO6UNm0CM56hbzal2u2eIXXVRwBliFA2vrJ8wHqujgGr
KSqz23Rn2DWwHaF7c0MFTAP0Yg9vDpvuUlzPKCf70p9ovpP8iI6bZbYU6vyzhpNb
2AxsPidcwKkDqR/eNFylxC225I3XP7+tRFwHGVQFisAZFXr3UOnS63giX5oQYbY/
fmU/WxPb11p66XVUPakpKFRS0Wzld8fqhTmGYwNJ34YQmzVBNcYA1yiarvNMS+aN
ximur9M0pf/t0Ozx4tfdyj2mIFRkT/fQ8By32V0pNdcXv/0zTCwqjFmkIq/hkyBy
E+GvEUUYK2tfDWYi0gty4kSwR0c46ULIhrVNNDblifzcSUvn+l5ARTBHSGVkJFtQ
DYPV/zf0vXu55aWEFwBAqxhV6EsT7qMoVqsfg4Rd+jq9JL207hxpx7u9r3gE8oG/
e8dNoUbh+ABQJrRzJleuYvY/N8colDTSFDFs3tIcAlTg9WeYpMAugmqAxkbXZTb7
ja2JGYw2nYFO0zyxUrnNEYYm+zGyq1bjcBJISeYwagbYd6fTdyFdAoWgKWd+WOuY
0ZEfsGZjj+30sn1iCtoG+0cFCLUOniY+NppCZnzVtZjucTKP6L8EmxW76GNq2NMu
3GG+c6UYX9XKrNJy9vhs6kjrj3Ut2P8J91HTbcIFis2eVfcrGRjb7TpKBBEGTyMF
y3wr+N9AIIbGXNpKWapinLc2fLE8APCNW3JeCe4tNxdNKbsE3htPWSShoB7XeW11
eV7TPA0cMk5rHfyCtAM31gPIdFZhx35VY7t9Ysy9G2EVe01Ndxx6gXq+CVNMu35Q
Djv4M+WO/TAwxCWQlBf/Kb3g/Ij4o2GZL0Xr+aNIxBJU2xaTSS1jdOVWi5B/IcKW
6//8oQNkpLusBXcwLmqVMaVgQx7iP5NvR2oKkT3xvtGvNSKNDrfkZSRist7Y0F6J
bmL/f+lb6hJ0+5RbQbHWTXTwm8cazh2tvZkjsIdaef7axNPxjngQNGgYOW3BDTB8
mUXqsx2LWNA60mw2ZJ70WD8nA8xQYYh1e8lyriCB4MwC9XCZQNY23quyfSQ72hYH
G7spTtdrBCqRX660baF6OWlr2a6/iFfWyh1RqTi2J7oDpNMdXMaSyOigUHyvxe68
IqcHeF/3/S76ijbgKvD3TM69GsI5AOayYk1pQCKv7WeoFzHG320EZ7dqLLeSZQaQ
07f632SkUWcDiwD4Go/AKtrj8C5UogzSTycWdzUbYyWLygiD/WUlsfq/ejcUdgNx
zt97kyVGvOZ8qp28xPiPSpp8hqy4mCJk+Pb9IYmFHVrgRzd5mXo0Tm0q3LIg1thb
0jnfD1IIYcMC+I8fYj9sv066iG/7jvYN1tqkAA+J3wJ9I3uZNYdyuUaZy2XKiIo6
1A1kuB3Dm7NHSOW8hMiI0WioTp+gWxSUxcussN0YYpu8pU0L7DE794ODXTpqwSFs
8fwpg/P0xLzmiIvYWHhPcUg6vln9a/LoY1gPgWOSuWpiSGQOS5dcaBHzVZ7CMiiJ
dyTZmnHF36fXGN74tGMcUb2wgs3JUaXLlEjxpdnZFEdC72mpi1T8aOv6Ek6dzDw3
ec0bDTWYvwg1QuXo9G8tFBSkYTyeuzy7BuJsSxDKTC8cUN5xRNbeswgHWULdnoFk
Tfl4ta+eY6exE9C8Ovg3rwnNLF0VS9K/Mtrdpo8haWfhe5BD5TaPDslb/tebKyvc
u/LLjO8dIdO0wFSAIqurqYPg9DjspiQ36JoLQwURTKJRy87UYiz7pEzzmjGtGSHD
W+r9eef//FcPRgSfQqr29yghafoCnj5Y+FQldvduSj1F0Rh80xz9zcfU9b5/XBji
81x9TCNHJH6Eacan7OpSosjPQ8gPQJBEE9h6ZO0thqIy8Jwf+kiKNYSfA8pNqQmp
tUDAW6zxCpxDxKlRVnoPm/rUPKUzDo/Q2YJtN9pxy3mni8o+VlL6WRsNoltrjLAu
ESTmdnLRbiO5kUZIcXv7XkCODTW3egU/swRWKsAQTV65Le0uMDC1ylm/B4F5+zqb
5Glah1wANut/mw4zDspZe/g6sKkZrQTFaA1TeUUODtTsr+18tQvz6f/mVX2yM7Mc
xonQ2DYjYUsnBVsEFphv+/iPd92ndXRHmiST746xFDWfkqBtAFAKuQQYX8LdWiqg
HKxDVLlx2nqYGWPAqvAnKh66qDGd+UY5SUbwNmLmQpXHsM5WXjlsSAW4nSDguwnX
hBEup0NVL/VyuvBHP17g8pXJDvicF3QlyyfSAXT8nUktBfENhm8gZd+uw/aSSH1E
58eR+OHKCuH/bAuFBZUcN7z+SMINaBpcpuXXTPo7Up0FY6dX83zHcwxDdR91mdKt
jtn2gOkelHbVaq9aFcUlXAmPhx3ra4pjUyozeRkrIbjI2tnI8D9G/vkCsnBHPaQQ
2qC3r2AmOmzCG0eTxgb4Q3GiVdZUWD/FxLTDKxN2IyAHXL0WqaT5lyQFpK1m7J8P
CXqdrfZyozQU1mLMf8HCxomf5Fsnxh3m55ShK4Wt3VW3+enaCGDgd+x4SZNVYHf8
tLbnVoml5Z4LCXzhy7jDYtCIeCBiSvpMKbXmlz1nbIpuqAYtAydltQNBqVwPqdWB
nuBBzi3X2YLj7F80DlYVhkDJYpzbb0FyMKMsSA4mp0bJqwdG28sXNu3D4QsWROJ+
Or+0t27lPdS3+P9/XvuoqZ8d56LSfnsQQI3z34LArbTJToVKMaHBxZiU+nAzwbiE
FhNBCJJ30gbzMU3GZMonnHB/xJXDMQWWN06HzJFyZdZr9bTtPeP1aRFdtY2utJdM
w3qGq3nM13jrY/9Alk5nepYzUXUGfOF4oOUrwAorRzuYVNdZ+uLjsQejkznTnFzV
3jBuVZMdkw4+QcDjOcyZtVM266nOJ1/PCRI3DmSL8VNVjFmMICqU1b3LgrhT4/Kq
dYTwCanANeTrnourMW5TTvZHXAktI27NYQfYC0WZy+0BGqgBdgoArVp7iScArs6v
zcVBSXPnaop9GdgrtxV2QXNK5eUZWe5V7GlU03KZFvYifmxjHyg7KbsgzBqo9ojO
+td49+6iagQUnwXSFp7GDnwAWXUyIXrCdQPPbaKxMwcEdB/YkfniC6/Ka30hjaAZ
UCYqyEdktVY6CCnVxfRqLNZzxUVTQ4Cuq9Vx8QrQNf//wzjK0FPal3nnMNt9TN0f
1HND99GmiLoXCgPEfhHpwSqsK6kr6XrDNM1o3n7i4GSJLCC2hbHqlbbASgjqTKFc
rZ0A/6yIylhpLiBO8l0lugeFOluhntqR9/m95hw8XUsa9jw80uQrHXmKWLxkF/op
sduI8bRJy2D+VdSEoS81XWN2Wtc0f4VrKnww/8wYLyyMdc8E6lPRbP8LR8Cg5p6i
9fVa1oBRmOZY8TcNrezLdWPVgo0H9wtAzUlQZNRTHUb9OJwo9I3bbEOrr+RXPked
aWQThN43riJzDHOlmfNUHNbanuUbwQQs0k0uWXpDlY9iV0ctSol8rBoO9sp6TP7I
1aGa6Q9fp585GJvC/mb1kZPif6kJUc2ou9pfqMbOnMZa0gyb7h2xG8fmlAwxto55
QlJMBaHml2HqUgjsxQkgreTZYVSdcG2pjt93RInCf0Mpsa+BTFO4n8oDbunh8GUK
yBLFNfZKO5uupHMpInbCVanOxKb3Zo9h0QCLS072MD1KcRFKXFvx348h9U6wX2Su
rOQmFL9ACvIKMWFKW8OSwfensipedcqgjvvmBXRFoFwWBIGLBCCCHrSZ45QkKu0a
Nn4VbhQBiLmhcdHpkIc+sYkl3HI9oomByGAfHGxYNJ+Y7YDn+GHPdJX5vzIemgGF
gVK8a3lg4UAaIl2BW0KC/auLykPQowduZV+HzYDpyEnB2+8m6ZgZn330YIcaxQiR
JYIiAUXZnpEyJi02CSowYEVQglQJk6NwaIWJ7a0vbxvSM509fclvxVrphj1tR4Hu
dZmLA3zFg/PTtgXSEJBXaQFQxaZ6e/0s43a4XF9ZtTyjQumTqUxysdEgflvDi4/2
kBXJ7gkNFC+yGe90jCBehUgVMhrsQ+LpFELOSfFYtpmRc6gLN6OBFlodahyOwnSS
AQLcQgn2WY9mTaHsRoxy80B5BCHhnIRcluXwamKwGwXxIDWgRL7odL2UcndrsJA1
7R1SwLy1YjbZALNI4iLb69cXnjj+22psCLhv26pch83EnxEwgr16BhXYU0kFYxuM
GF1pdXIwecvr4sq75x48A2owXOXc7BCZm5muL8DGW+rfeyGAtBx003kNzF/u0fPi
fldDdCjM6hedyNsAwMYefkR0n+yIOzyyhjvAhbbbmFZ8WentheXz/7l1xldjnpKi
1eOTJvjT2/k/kHwLLT7ISHCsPNWOHpvIjMekcjpBqKFn5ayK/rfuqJNdLct072Im
gCCCmTc+cFFK0dNiMHuejl/z9qt8Rg97Pr92mZiwpxbtY4wdIblLFsC5ZPkPrTpH
malg2IaLt3bJ0eVWFCyCQImgSBxqXQ65yGe1C6tMIfLNBBADkj8yLIP9qTtoIgdn
6l97m6J5fJ/RX0/zDE67id/GqE4KbhugrwmX0l14rH7ziLgXmwmEfE7tZZcFd0DP
9G3ZJ57J4pVaCgEKjbMqemw09oYxfOFIiztP3V9BQt2xklTWBKyg/NasCa9ZeWjZ
WwrQrznjDUo+beYPVWqEbPzsvctvUzEfA5QdKdjkqHGNmZMUbaEGsrVhq97X5A8u
41zPwdxRtQ1uBMOzw00rXw41KZH234MLvc47fvdLINRCazP9YQpg+wHD/lU9XKLf
EGCGbTm/lKqQTmOPHOYYoAq2ZvU3e9U+CSWLb2tRHW62FM/B+yqNExkNJgXnf61N
Ufyul2IlB6H+3Uw9iXNkllcGDx2BEuAITEA6/q7rIx2Bhzg/biTRHzDCQxdufJCW
L6umEK8QZXuidj/pfJRNMH+Sv0guhoBot1fSkZV0UHr9mb98qWJw0HpK/q5HkyHx
qXY0zzCNJOZu9S37L7HAVdWr3qVGYQSNtl9V9MyehaWQlNkTiV/sRu5f53VnDJYZ
GTpgGITJpg6eicyfqwrjX6hAlqejbcjnaU4JlrR7aI9G36rEU4lUqrDecgG3VwIK
0ihsbsAPdppMdtFSFzqazj5ne8FEQ0NlL27lyQN8SHTjLeA3vAMYuX0BPd3jXRiD
q4/vAg5gdrEwHN7ABZk2Zjjc6z/7h0xxVmjijvD2MsJgJBE7bVEFndtAUqk9aM66
bZdFOtOONlfdted2E4K0k1FthxuElNWY0n6zkRCVhBAl/TL3W4wiIPvSSeTngxrR
p5vQ7BzOILKdhY9DU1nwIoFHm3HCVZR8d327opMEakPtqWWzY3KisG0MpbfVNrp/
61cJSmT6u2xu2tIPZHU9muAJWkX2NVsIu0/keBnFltFTvJPe4iLpjZ/N4CEEzPJV
46KS6LLfFO+u0LEgNFis5TkqzPL4yqjgR2/4Xvxn5xgHj3XOPpm+Ty95T0gSyzrr
khm2e3CQdPKA8ad4KKW1qL95i5X4n0IOnoZ3pujvW3ruKzQwBBzCwDCTYghApJ/A
T46mWfxDhtzS6EvCL59OCSmst1guEgpeXJ4Kw0Em6wNyKiTTOCeVhLhoRLMwFU9h
3HyCdoKTwiwe4cGI9WXwA6zjF1c2ek3Y9D2MKno/hdMzTsLDM9mIbdr6mS7sNylA
pRNdWmyVspbUS6yvcTChv/4c7AAgOGFQR0ymaRh9ohr46BULLIycxqY/4yiZdkQg
bToFhwPF1MsYSIh39zQQDW8UEtu+h/A6y1Ka/S7/Bz/iYCP7AZKNu7Nx+Ce1gh3j
ov+BsbbUo7nlPVDEtpKXR6+ERXvbyVa8TnTYRoje7x1h2T5owW3+cpubvixT2eFY
rtMedufpfuo5kooCRXdQ+M1p0LvhDukP4YCiXP37V9QeriLgOSz7k7r72/A7kVgK
HCq1fNQ+Lny82doCxnyjV/NZGyEJ9r8x/qgHYbzAusa/mufwyXUD2ye0yEvIVVh2
JFppSBYPGUlbrn7RSvyNtAjUQkQQggMEHiR/S61QnRldRNAFQxyNfVMqinLRqPaS
EQ5TW6Ilx8WZMQjC19ld+CH762fyxlH/wFu+mlNB9di8H0yEGKuSy/9Pen4THa2I
SyYIGR6mmxUE2ZUMxRipsrrbhizdzIjayEpAckV0K6T33MO9dy4lchghMgILFyfi
4YfPNJ7TLEwzjKTGYVV4pddKyh+kn5ozbm6p+kqQ1FCJCWDTf0NUhSj4r3v2bHaD
DM92jLXzlWlaP5YhWFO5bKkdG1tmeGC698zJU1E4YFO1/99mZLgkpS+szaBxxNlz
ehrZPP9q5IJawiS8AXIr1T1ei4Y2qVxTb7YzrmMiDRHIhWcE+RcvtYUSQCqsFcLm
YFCU1UIVIxQ/mPXgUj0tK70hkGvtoBJkr5az4NK/Qp7cPLU112p9hG+tW9/vUWz8
vLyF0eUlV/BtRDKWCxSWiLJpg7g2qZFaK9nI42uMWIsZoxamBGV9XIfrTHOgp5md
cqlbS+p3gyKrsz/fVpR4cAiEfYBOxyAaAas6GHQeVbo6WGRfnZSQCQTFxbRAglBM
eiSOK520yx5Zrwmrd1eZCKndbDSruEXr6e6f3yGCIDqzQc+bgHYSMjBBJiAaI0lK
6S3Bp728AXeT7BVJ/jNjm+fq5A8VqYXHaj7AUj3o4OFyUV5xbnKNuRD1Ur1wq6Mu
ZZhEqg33NBVwjM2JCyNA1ayuEZTwV0QkR+9Qu+ePgoAzWzGYg5vO200dnKbCCC5m
Gzo5jquLPErD9ExEDjtlQsKfaDRlIst5tpf4PkSduWvbpc3VjNNcDndIFW1lpM9n
gNo60LAPao3liGfCHUVHn+ApxqBsGnp4o82zJ7rYdscNTXXU8YKuS1WypOFQW3ql
sDiVGlldr2BV9KspAPi0Sch/MTOZXXHTkeoC5gsGLjsOOjF2wOVlMvK03T+gf0zw
/ccJa6n2qlDeB/VFyK2IN6goMNJp8aaqd6KVya6sImnPn2zIDZ5Lp7ZqXkfAIYKZ
fHIqdV+dc8Udyv0sK356jMnbe/SFGrA0AyjnNf47eM/0APByIf68lW0MdG6x3/+k
e47jFxbpsps+KHcSWtg/ku/inTMivE0uRRCeWHG41NoYcaaoo9xgq9JZb/+H7/sB
qH/A/qgPmbTTROZw950Vu4/svbM1PjqHY+BcVhlQZ8moH5sfhMqAqj5S8CPwau9W
6ijc0o/rRrIv4VNZWmbqYH2PD1VrVCMPXhGQMUElC07OtsGN4x7OmPy46DYy3yP1
ErpBv9EgHh51Bkq4cPJtWMnr1pzXHU5vizWYL1L8L0Ovsgzzr2rGZN4gaimfhgM+
BM6OpARQowT+HjCFehIWk80D6IubBoVpvAqN3K8smpuoyfKVV89TlYz656OKw22p
pJCaUPBQAF9Rx4XXV8tSj2T3ngt4YoDdTs7Ajko9BDc24voo1LOpzEkL88QdSK8/
/ppZPx3ENU6GlNVPWCbvjejcffKI8P8ZeuAiZwFMmF80pP65UY9XdpGYcb11oMfT
I52hnS/h4yf/2IawYKX3b+v588zATEZRrcL5YzGC1fyPEgf1kxaeil+OaNO4sAVe
VoxgegRXbi06f0IVjhDY0sq5bKXOFtPTX0InIlkQnHJ8Ox9vSnq6p5puoDiqqafU
rcyPLejkjAXE4egWsMV1on3xWCisrxh1Txk111tx3/G+2BbAGbRffrSZ3A1Nqqc/
RWIdm53tiN81jLxlIfIc/tXtBwfio+aGgE7bRm257QnHkc+Oi7P8au/ZIbSyz4zm
HkNFZC6jfamnxy3O4xbTfsYRkB09cB+eiMuEsZ6bnOTd8iPYndX2rVNW8+NNu1iq
oh56moR2F8ZHJPPLfM13M6Q5obDYDrkTrWQlS674uii/QV47zDDDhFLPCtUB74vM
EH8Y4Nmc4lQJ0JkS+oYlgab0nKngmhtY7S2CiuW7RlEfJoE+IonjkuX3P6i8Nt/H
w5U2ZOh1NQ/QInUw6TWq662BGiDuzlE0Zrvww0rfaOWw3zrP2jfY2ennvUMEK9oC
r911rj3O+mrri3r84FoY86O8Z4YcHstnkKXJHikcvC+LunGSWgucvwYggrDyydCL
VHzu2cLb32cNp5IhLuxYeFj37U67Dno8mpe31LRiQteAaskWMR7aVc6iCOqLS6oK
1ADqwf9y+yBvPwPvIaFGaTIIe42rO+aP/kZQU9cyix2kPBgjtvgj0135gwKrYjo/
8URjRRxek4ETXZTtM7/hKBglkgId46cwY09tZys2FqCmhQG97M/QBB3EJhohWa3Z
Y37NhjMVd9lVkVoSv7722at0cu79BBeTa+ZZAQ5ci96czPbHbDVA3bfPoo451BCG
ZPMZzmabcsV5JnUzu/9fzFfFjySVyTe/fcNppl0xhDpsub8KgfrMoRX0Ly8FxU7j
KNw+qfm1zutOlefY0zLC6of2UeCfsNhMnCZGdr3dd7lllek83p/v55R1zCosyFSJ
R+kWB3yIfV4KsaCFXzHffM/OAOQD/gpRb1xSVln3AeN6hob5zsOEYuAcrtDgoq+7
wVZMwU5fzITQlYyxawvhe085PMwWZwd1pBrwZDxrqE+XWqNfl/Sch+Yogf3qIar2
gtgbMfN5vahNUIZ6BX14KrTDjj+rW2uXbNLiFFWWj5w5D2hGCT5qzGRBkzgvpaU2
CKspPSrg9ALV+g+u2Xc4195YL1Ykxy0QR0126D2gdT8g6QLBv3VCbeDt0V9mWxYX
ggkpaYrold1kv8hSS/yDDEDx8K1eFvCbOqC6Dm71o+V8j3uEIAWpw54Y1Vqk9OUD
AOnVzEr0hi7DEqRMhpX/S9CM500ueU1hnhi4FPQyzAb3oMR2E72QvBogDjYzZJLC
dQYg5zRHLJxcrR+XDUduJVT3MBqvcYZGi9hPg/szGfCwTBMzS+DSPtgSIqlIyKmS
m1g218pBynOQ7owssBc1ND7dap4YTtreYgupWURfNPY78CYRXFwB2Pkr80YuBGB1
3js4SSFmTqQq2sB5hWZFmyVVziTmEl0JGO40xmZwb4C56MVEntH896MazvhrchwG
qbTza08nQSxT+JqzRbpIeZz3wxgs8a9PANBzv3hOO0nEp/Eymfudv6ifwSvc4hM1
H44DNGlPEMc97dVsp4YJyYgVBiS+NEWGLpdE2Em1O/bpSt8fHmmBu82goxK/bZyd
FCs+rnXybQRzWzFxCtmkktnq5dCBB5T/V0yTvYOA2Y/JRZ20iIX3l15b9cchksTa
qpoJtbM7cG8eGgCuxAyzbUZ2plHm45Z4ou/Vz3/+FPBEDqObWCHYQsmgvh+Ad7Sq
tSIlfP9grzcCclFAEZi9PDgt1JKEAO4C34vFVRql+S+kZON2gM94MQRCLAbte6Y1
GAqVjux8PsIsRXj46lFBuvuS3T8svGrpWJj98+MgZC0Bb+0UeIUqE7vnT0skPBoo
f32g2JAO29St/mRQf0/A/9y6UtgGkcZSodiKmhmTImwgMLPNDLk3kw6YaNZ7sOya
IGgonB4PBAAR9wtsqcdqlLKcL1C3LELSYF3rwiNp7/CPYMjF33spg6NAuemHCh/H
2UZS4J2/nFlAW9yR4VvxQ+mVYFriVUVn4Y1rdZIwk41EhIdhkHE64EoqUFYTz+cl
V/rE9OWD9QW7AmKf0MuCtQQ2cf6Tog60jjZCg0vN44/BPpExnwZyS5UDO3XJfs5r
by95OUzLMc/1UqRfwKcWCtRaMpjeBqJe9iwNRKxuki4iXWIe4Bqlv6HY5rkchdo/
zeOVroW5i+aGLtZVx1ih6dJyRh3o3TA38va3SB5shjY53Im7k9dQghUvNWa93g2O
OZYzmMexUKyHGhZsKIQy4MrDU0JS4TVvGUSgMNJBI2J4wGrYKDdFANTIRnVP0r7u
kroRSKSa2WHziWBpf2kARhqXx+G0/CH8N04xhiLbYrv2vZVMwszcxu/1E/r9LbKR
RTt/ufZYsDny3zt07NT8MjOioYpHcXvekHVmR28c/z760ix/obbMMySeK0pPRv+1
+4r1+cP/MgCN1KLbWbwXUSADixYC8ianDhZoS8CKQXtcRUY9GM6T8B6ctZsC3X+I
BP58v/B8EmLUzob8SOZWDIDyFhKpBQcjv/mGeKUO5AhvFe9xto077oVpG2YxlHY7
DsuA20Fk+zx+rCdeCXH/UbZz1mSTAHyyYRGsOb93WR2Gi6Ww9s2mpaGc7ibPshy/
bRTRgYHim5thq3H7MVoT2f6liTrFSHVeYxM+IXL39PDV84vIw4jq7UGbZ6+fq1wU
3z2BvliHwYu0f+puLSVVXUNhvk1u2csT2PCzoVdp0xd4x9FktO6cwscQibeuzbSp
7QG6KPSuIJeJ1pi+V4XaqJzxc1DzJ80k+uaPiCk882gK/UAOmsARc2cMyLkp0oei
kJNw89ea/gfqMx18HiLIuF0ogZZuGtJ3UoW1FtnkQOrJBqbOscTo0xpsJZypBt5H
/KsXRDMy4BEg/d5YvtPrQGi9vLBzy2CDUoqqBR8tgbm483qJO1wHYS0iwOYpnpSr
L887r38fu/FbKBi4JQXRjvgxKlfkwrtqYwUOci50CFHgU9mFmG4lghhH5Xtc5cit
56AkPLIpF3TgMB4vrcFDLmNnShUaPUBVkfhfal/KsjN6T5YVFNYrN90UYOnw3dkK
jSlAOkJGD0dUhUage2gtzkdEeK1CzCMf/4NqXnKVN0RY11lkUDRXl+5PVnBng7n4
Ar2aLCwxcARDJ8Gces3CUDrJYifj69oJlkpzZFvEvk2QTreIUm382v4sgfKFZiwc
ISsvowUkENcjHCJWExiL7OuVSvk+WgNm5ZGoEJwDIpg5NoXpE/GKdo3/eIKdXgwS
i6CsBJ2nO3p6YoEF7s/pnf+U6xK7x71TG2QQsD4FytwRqrzd/TZ6IoI/WgRNN/t6
szXDkHzM5suBFpe+FCuQUthVwc21Q7kjeSQCnjjl3BxgWxLZev2P2iDANFRdoYFl
vdmOO6ArLQIRD+dp+GcyzVMrt9nSoMePKQKocn1II+8YHdMnBxPDcrzdVfbuHrv1
vked0YXM7xPKgJqFDPnN70hZxyulhvWgi1HsPBSXH8pb49afElAuVBYNVPym/buX
pCyzCJQFgm1KoB7xvw8HtlNd2KVumE3fMoouijL43lRLWQ9L/ru6FQdR0s5+LIov
Uz7IkWa/NentiIPYVC2mFBX3eKydxYWYptkZFkkfLnLNriiCRBJAgn3JeuynL+Ue
FSCPeu0+pLLiK4Hl3iAjxBEoPd1KCXfx9Rbivfzr7Egh4bnUnqSyqivrXLJKQnIO
cpMpqVkzAgrDY4jgNJb7PKIQGCwmBTGDdelVkiTpqHpu9JuMiNEQVMPAhE+i7Qsa
2yQ1XOZLrQWUeVCnDYfT2HclOLcw8v3QRjvCrYzoCMlYPaWCvs42ZjOmhgOIY/c8
DOpQ42MuZMttfSUxM4w0Hw41YTKH8i3rAV6lWELo6N+z4AYmsw0/EUqggWWcL00c
xwojRS7+2tn+/IDeCWfwEPZWPZAXXR5iAh6J+GBtVOV6T2Odw8MxWBsoeW1fBD0g
ibVaFUdz1K7uxG/cXmW/1kYqTQ738SXvFilC7fcA+kqvp5KLvjJzOleZ4QtxhTi8
MXBeWPgusaYS8bTW0KCKKQwjaW/jYFK+S+i13waY0Tpg8lQJbNOTnafd7q3PXWz/
i1LVS/uqHKZAhDHUos4a+0it+2Ar3mEavm1jR+8w5KKNbD5hCDO4raXfkc3XbsMh
6k4XcHVGzZRO3wHmJoewe0YRjp8Zf0sFMCRbcHfa221nNJi87GP292HJa3P8p083
HZRQZYs89FAKgaz47RSP2yjxi/lrXZvVCtjpW8lZVPfIRy5AW5xBtNjJSmrY6ftK
G/dPEr0EUIp6uPuOfjpBzuNMh1DO6bPtPHj+EIGAuhauqkxmD+uq/0UxXuKtkL8d
xolDgnEFJdQFLylpVxrdrs0htnHIWBtaxJ5ac8TAX7IY/D88QT8T38HLatksR03s
ZQxrqeqzu++PmuAYL+9X/QucOYJoD3jRj7KoahT276TQuoboOmaLYTCPKECHreAi
LWYs1JKoBlp3iGwlcq5PJSfM0hyq4/JK97yNck0yMvlOmGMP/5EJEBerGS5/cGY7
3+8hgVD9RzCnFFMtQz+RHH9d0Tr1WyHFIF6GhioOV6OZm5GLjHk9kOAl/mavaFDz
R35HMC8MoC8fQkvTNDgy7LzBpLchK+OGPA+pQ1a3rj1bLYS1nwxgqY/16itjM139
t3HB8TkBZap8qK8bgJ/OkX4Plf84pXm7AudXxHRvq+u5NgD0BChnk7EUirXQClFo
vxMvGLTAh/ZWEDBwqygF3ifmWVKsvoVyGXI5hVMuSx0imA/iCzF9xbfbiLKy4hN9
v7dtmvHncAXp8op+LhPunYpUK9QqdbKLrVE8GAVr52gJT2eMVTwo2Qer7Fe+aCXc
br9xBcFLYnf73s07FVoFn8jV5Suai8aVVgQTQOtKBCLEeCZF8xwqlkU99kftilN5
0rompSAOfVNGi8FJZ94eyaz/y+GwRT1UIfwGyPvn1jVjVHiR8FE/Vv/YGTwYwjct
mojwAs8pVwf7NFXx9+A5gcanvAICgXlvLLnZw5+3e2V83QaBoY8rv9CSp1JLQyxg
w0Mr2AsTkXmJ5Z/u4w89KPsTwLo2kohIPBfxR+jJ5Ieh5QcTpkU0E8AatPJtevle
QujbYVwcy6oFdIz0e46kys37vdfoKQHD6CYStSAifIcuFTi2R03Cb3hCcpmkdPTe
xEpq3cF9ghA0cO5eqprbTj2LipvjtOwODvtfSCD+clvRp5v2Kzb1hA9mHuIjBCJP
zf255RL2eiD67yUuH2kYCTQ+UbN8zJee39Yz/0viNIEkzcekXc8ubYZTYxPjuMyv
uFpX+4tMH9WbC6IiwDYSlNppuLMhoUSgPZ5+ffjhBINCB6U83r+luzDpYkf+2Srm
TXoVshg5uOPfrooPyDcJZay2Tn1rPPEeo5V3DQ6ZH+wLlUNbsTVT+d+IexLaP6o9
K7cHMsTC3RfSt+eAASE3+DI0QIspLkjBSkOoH8w1JwVyLXxpuz6UQ9f7vEFmeOcP
jFVwW9GgxEV79kZZhjJ8wOPLresMFDvMO0pPteSojyja/quvLLKI8bUkB3HMszsx
EecLjA/Rs/C81V++WuVnhIGEPwqaOPybkGOD/6rJcsyloazgWpMnDEPU50xe6UTH
0INjJZ0G7CXm4xKKwOCnv3KRvB/nYnBPC1p9EGcSZcfahU6tSUS/VtKuTSnBqZqp
PJL2wOgfKl3LDTETcMRdgSRh+MMxHGpJFj9Bx3Rde3mMp4puCpsp9NugR78KwUg8
A7cDTaxq4NKz16VRzrkRpKtJVWq31DBLLHfRgF3pqoGE7tMveYpOobCBoGCL8mt/
1G78mSoWwvUGNNN+esj+QfzqxbXVbdS8/FN9UkzusG66LE9tM4hrNR7+jmVemBo0
HxZ+A+PHPzjDGMjlV+cYsu0JDADMeW9SL8Y8qaLCK3eBXpYqMbDz5iYZ3B/sDV56
YeuBrw20nGgpsm+iRXneiA52e0uH7vBioBfv7/oIg9ZXr+W6mJRve9g+npUeZ2gY
9VJnt9Kf3olvxN+FnprqBOKGJxyd5Y/5Uiax7moAN6jdSr17rKZfeWEZS7czTDs6
pN7RAdOPBHoR86dbs2loZMuYD7oK3+1L9bEyUQcOyO9pQT6R/iGC7BbVLKS1OcrJ
heEyIe7qZo422lx/l1F5jf1lon55AcySmT3o5jDKvyvZv/mC1eY2eiSEjTy3DAys
9sEDvmHZJCnM4aZeU/CA2wOf/a+M2yCenBKeDYrPQIejaB9jt8ONcqqAwu8rq/VS
XO73mjqN3Orri7Htbs28rGP/WJuUqJS1OqfDsChURHr/Me2gGxASoJsag/r1rFrD
y+KEvZrDEUyFH16iy2O7r9o+K+V3SkItD+S1a4TVXuUl2OBndoM47msYLheWeFXN
PdcD7xqz6ZHeIN3q06gzXCm1ALOWd2jnGKQjnz8cZ2V8471Plpg+4Tl84/eJe0DD
t1+qsoJBdLpCaZdvcEtMeOsrjlXeA+ZXr4SGBRX0gCLGKJGcYSYyNOZiLLXYlvmJ
irXWyGbJmwID7TgzhdTNg9jUXYk8RtXLXTwEJxIJTQ69+i+DTJF05xqw2YqdRO0i
UPv9ce02veiiKotHDTB36gIjUFby5wVGwT8qG502pJ6KxQ01AatMApBWuPsqyjVN
TccCdStV+/q2lkouQ+gcfOYSBCcLcfAOOVbkmswFm4OVVaUlAsssWr+15zi4NZk6
oGOUzq9T9WxykWimM64wGrukrrEDBetTC5wT49tl1QyqeWnyGatTd2CXeFQj34Mf
ic6dINodSKj9VMno7sx5cUlG0DpVAQD1mnPz9plFYHIhVkN7B/jns20whr4W7jPa
4Jt9DR1bIJSrNZR7L5vI3yyBIhckV4xy90yjMf5GdbsYZlm5eKqRqKYCOykHXpa5
DJ53IilgxUhd8gSuOvKPJT67fKmm8ki05T9DWoeyLUhWoG8NpnwKXsdOWaZEHMaG
1S7kjHDrnLAcF/Km0Ts3Zx3ld3KkJXO/3at4HHlLTS41xw4VcuXiSUNzs4xqcEGr
JuB9RJF63BETojXxP0OiBLZWTMj8IL2F7Ik0EtU9pjrnzW+9EfIOqnuka/kD+V5L
Ckd0AGAKrRjnSFBG5lg43EgY++bicrDoeCHeJUSJVsQ+uVCfyl8mQLwXeLh7rp43
F1jjueUPkocMP14UlEjfSGZoYaZ1Twk+6QO0EgCUEbTh9pxxscPCZLTrZyCvOM3m
oTQzCIilkwU6mE9Fac8Kj0LNCjE91wGSvfv+CY8vBiPFRoornVQBiZFRG/dMzJyf
3eMHfU3iCNHKwMoJIyjyEYt/kXnlADXalKdlvvJZ5WhAaLocf2VV9niqNx5f6lk4
VIXgDbotY1ANWRDfCc6lG7C4aGGL4P0/c4kxBAK7qi/sBS+IWnFVx7k0RDBfkeiI
VWJ/OlEjIwyeUzdnx1Jr8f0psRSnVhmgN/2LG1Ej/QRxElsVn6p8G2S/gQ4FsfgB
0byVnPUI3TagunTDXpXrP+MuTxRfPfBYe2FbIzAAySiKm/5uhOi9pmUf+kud4CiS
lI0O7aiifesXHQv8wNRDnwBUr0FiH19LJAud33FFPF7jdxzOUE9jyG24z6p3eIiP
f4lkE1KMqJin+XWVWVWxVrI+WKzAp+YaRX6UCB23GZiD44akeLBwAEUQceia+Cc+
0geVe6eqR1SG9RGA6rTPJF+yuV+ZonitdYotakdCcgiAvcolwPMP92lEcc97SJbN
ogS89Wx2G8dILtK+QUNlKUopLp/y+7roJ50Wf2k9UKiO5b7zUSaewqzY8kSvPQOK
M55iuYH3xQsfCZ+kAumYGdga07NJOBAH/AAjItqd3kSle2fbP/1rzM90i9amyRAq
K82AvZRzIJkLwobPu/T5lRtgUkL29mwXp9K03f7HYodkzv4VrxV1OXX7sq0SXY28
xPTiYlzbmUSCPkSs7/RbpbtgKbXZuG454JwescdTpK10YMRarcNyki442OZiJcnJ
uO75INv+8CntAMdWCNvco2pFWnsu1JF7TAA5DwlWOih+ati1DIytO2He65CXCZ1K
bfWyIHgXJSbNZmp1C4uyFz5V0Mgz+RWhLNKoG6Z5nss7/6I8ShWPw5mwexzD8oax
LzDxrII2tizs7qkb1L/dePwOB5NOtF9CNKsB5alQpRPMv6HnBhd5NRucvJZ7NGpp
DUknruE+XQYI2PystxYWqv8cf5tpNrQDCD/RfTX2kL8QpVC040/khRZPBh+5+q0P
v92HZ4yB2l2lBTwu7lyKbtKSuDvUI/S/PLSbPqi3yf6ZrLddk+6KT548KUSqhlkj
pLN/5HTOxWXAbVnY4EpNeTrazh6ulxP3PfeD+5rljZH34X7DxZOSZXS1C42QKOE8
kKCN4x1mOPwNJT742iPa+8g2J49Z4M+bgmUvPgJ55gjh3KfghDsrU5xSMrrQ/nQ+
chW1Z0ejUjV43K/pUdV4Av5pwRB5wHv3em3cqdrTqa3pWLC7oOS6sKgtdLTI1Uvz
QuhaYHKd3Hj4eW8uHOfju+ktXcKOVIH/NHUHWma1WhafqzgvuCKM/CV/vJEwx/f9
GeZ+xp1gxf8S6cmE6yfK/SpvIHWbp5uozE3+4xRve7ZJa/gyfwp9JzuMQ72D55/R
CymhAwcDHxn1S1ZGozEIyLjHjz4ceuOnZw9g/jDGIMAbxXtNIlX8FnQJQFitJdWD
rUoCrleaTZP+GZsCKzdATeJMmKF4fCaAyygeC/1dr68x1/fZAllvVyx5kOr4AcoP
ZkbhsN8n6SpzatTS1livtD1/R3oCVhZseVQnvstIw0B6d5xujN6sfnOYOfBTc/s4
ShoNzmdtmZLK89rOG1FGEAR49BAZmaEBkaFO/RnFdgNexNrNP9SsCCKuiKjLXtXa
8FK7FcCqPGe/q3tuRkX61kcHSfuftAMSu0YZ1Dw6QWAoj7/HcRoiGNHg3shVcskR
LaacGEKKeKnj7MgTa71BR+eSgOf795WPNovtrU7AYq+/z0eEpJHpwRC70/aI/GEq
sn0XOyXtGS2ZTRIMo/dhRwTJh+2tJX5Qlu/rA+56PNqCB+4E2+MKprMTdQLb5x3B
P6zZQdArtrIBPxQ87fJWyAGfPQZRPkEr5DgVqmCXYVIFCn1PYUQFEqs7AnFxsnRG
LT9KcRuFKVviHA5UFqWNiuicINkVAe6KhCrcgRFPq73oal+Du0vXdumVA3yRqCY7
VzeyJr/F1VENvxW0szc3OrFoMD6r/5dKjCTX4gpPjxsseQnpMZe4GD8Yr2eePz7e
ew80rW/dQQns0UIBNnLdVJWhimpVyOYqzIXtISCT8PDtBGETX4qRMEVNGjd4ruBD
JCeWDgsVyWFEjCWvQsb1PdEe0620xKfsLmBgagximw3thAJcc2JyNVrt0jIOCKyg
78geG+M+bzSaDtkaIVkb5Ums4eXAxzYgcsQ7/JutlAwVJ2uBDxQRIK/4O5PNzRph
sbhVB88N8DMkN0VwNKaTmCU/btPzDWLorCMm2Xm1MWeRIvEkugAIfeygAdHHaTxw
TnHLcYMfVNnOyLZ1bMVDkC8HcOyF4oDUjOzhv2pvRjcqmR9PHVe6qxtF+W6J3SG1
IOHRMGaefYhFLdvvnv4vjqeC4+aW9DX6qkf26vZ5+OeeyrX8GUk5raAMEp0H36Ps
Hr/uvYu7rZmUMzQFNR3uUL8/RNUzcUBPaKBD8wkLqq6cmnSH6LIPe1NG6QYEQwKu
wwYErjL3AvuGwBsC3dHtLFwzX18pPmdXWUlDroxWKzhngI+eaZgge4qch0Kh+p35
EXum6q8huElQ4b/IFVWNCk2FGb9WdafHYBG1DXFos0flMMo3rsxxmpOCoDQSR73Y
d+v38GKUewDc5HNSjewtrArLwFj/hKPm3PzgYL52vg2Hm1kl8lnaGAJw3zU1v53e
7upemEBY5gs3JTlibvrmqhFq9jNiVsJYhWNCPCPfYNY64Jlu46rVb4QNp6LUtkoO
yBacSyTHXdy8B1IGng+cSWGQP3vqwNS7Tmu80ILKOewP0JTkaSdWBTG8aTDfaUMf
3xcK3gs4fw0PTsV/I1EJOVJQ2MXzpTF+8z9gGmM9xh9lqQnscDJ6i7UpKVwP15IP
2P5r/YBwGVUJ5gkMNXb3j7hmHvf7c+pIKn/ervXIgTO45s2xTaD6/s+yXkwNSvCN
U1Sm8klDEjG32byqh2dLDwoVzg5/nNC1u9StMJncMhVIcccCCQqBXDJe+W/g3AKY
w2Fo4TuRkzNFYI5bk0m/0HHMn/hepnEYOTOOyT596HAKpFKwUNiHH3txzsCjpnyq
r/bz6cEDgO6FG1PsFK++1bezRcVbEqz82FwRRfM/fOx60Cp4+cZFiIKoApFxdnno
mPPChW5Mact8sKryoQvY6ZLdg43Dp76s0H4Edcwz1wRZyUUjAkB0QjXkC14+GqyF
cYQB/yRZEhnX2Nar15s6q2EJcX3yBR7POp7UnGBkxDusQyaNk9iqYRk+G0AN7BkT
ChccAfmXeV6J0uZPgIh8RGO4OYC40wiUEKPcDVNxt8HTX/I0nemAWs6H+IqzrW6k
Rhy36lB5W0d44yByrtVH10pIV8D0PeFjrVzlOcEg4YYY66qf1D1DryCfrYywWmz2
txv8QZovlbUe39OL+jqw+nvuEfpnj8UkKU9uGE0r78asRJ88BysMSQBL8VkLLlhz
1CFcHq2uoo2w6gIq2tVwfK8vX390TlNtS4L/Wock2n0FlbF1rjhrEUQdoCHlaLtf
6oGGe87MOwKwKSK2NLt31hnlAK9G/alDq1Es+ElK0o9GjCf3FiXUM1nsn+B2UprA
s9/yEjAUeBE1bEgyod/Yqx9wgfne/j9UfmzA0Z91BnyrVUMcGpIkKnvrExmjT0UU
BTiHjNQVna3sraRUx2fFLFy2LpCUSzSuhqpGHlZscJEbMCQT9/71p9HEY9XSwQlt
TvvWg7IEaD4mvjy2V11CZ/B4nEZaL84U4it4yrzfHWOD/Rr9kB/LJz+bkKcId8xO
cQoI2U57zhRoqp//GU0GAyTHmvrsfa7p/NOcCL7LBq5CQvWHUjsm07s2LAIXKQfX
iODlCt+gFDPVJhKYT0n5wWcMaEuFkme2ioesyD2V12v1c56XizhfLv21veKW/TDy
gQ7d2B7P/0XMKr/ekOAmEVkB3bw3kgme4oOY0qVVtLdXkssrGatfwwcQuHAHBPxo
VK46ffjHaTfyCMj6+NcG098N4ixBIx4dpXh1QnRSWHvSsBh0JFCnvRXC3jSLi8fE
Dq2KT3egGJrcOxaPtOtILxcujJ0M0eG9zDQhi4DDXWPfrHIIqX/aCR1vZz09KIQ8
oEKIZV5pYjhTdA/Yss2Lp7E5eBAzgycUT4Gf5SJTw3sgf2igyAbGaXy1yqKgHxV0
hhUZrwBRakSEkF4dMmrUkzojkBZl9FktQGM4Y4ZMgOvmWsx1TxtVjT1TUrybi31z
UaG6GyIB+DIp/U8kCoxcFIlZi4bxx2/xrjfjemLGtiVPPDK5gK0uRHDlA4T8AM7r
iSVD0Vwe+7yNYpEeO3YJUS1FqaxMDcAgB7fh7WdVZEDWH0ZZ5rKjybJtWm+vS6oe
RpkJSddds7gBPgWqTN0e72xP6twfhZFzCoWSUnhkpuCgqKg+AWxqfCyTqSdFbkzC
uS5tyOV2CWcNCjOYQw1JWjvGN+3AULxJe+PruFshMC/pAW0tCowPZ43chg7T+xis
Q3bJNnkGQEop9OcpbAP1FUnj+Btyl+1BKMMfAn+ff0nr25EOKxbiWmy1o+ycx4J7
IffCz4mOf/l5/oN3Mi/goRTXFtF5VIN37goKWoeQTp0mxQtZDBk2exPxyPNKTN1W
xHxVsyyB1ahFfhCEKCumqN6P7Eh9wow9h/GcPRasQsMbD1BobI5fDbXTu+GhA5+M
F/fWm37fn32XfPn6+varOkU8e0Xajpnf9DeGfufSwPI7RPcO2pfIKUCCeo98+rWi
sJlXH65s6R6H8dFLHrSDmHuvX2pypjxy10ekyeXSg1WPpTWxjTGXy9haKQ0k5Wc/
WjO6q97e9gVJcYjKRWx1CaMAe2dZbZ+yGJIAaArQsi2mWhyiVW/U4bixDBWWNvQ+
GmjK985otIjh/AUtaHAOIwvpuFC83ZSLOCwWbYxQM+ZNMzJQVsYmuQJ+9M1x23VC
3ix5PBg4fo1w8mF/u3uX+BGX5EcSIiVCSfCRMdV8Hm3UQQBC4obHh4nCvSkUhJ0w
vFFWDNNR/zppdCjiLxIpUcajjVRycRxgrTyvBWmVdvu/1X9I+mMGGvgyZedN0zqc
8T33BxRTuMNJibls9X5BYzdnZpah3wJiyNH91NTKHWcK1hSBnoLlw1MweA3EFbH8
X9XTaYWy2gEat0YwbF510DA6gKpiCddqeXpJreuurWJl5iF+2M7EQM/2HRoMB8U9
1/2B8Uz96pgVy+BXb1HCeelFABMGTqCf35W1srg8dzJkvS9B9Vghl6R3kv8Np4JC
KAZ5Fq2JKQS/PK8lduI77hEmQQ1TiBViKTlCulSZZekpqKStDrFvlzc8ccCqL6u0
CYxfCFsyFrvp2/9AiMXPtMbTG6RUDWcxw3YLflaqPqbc0fZ00UPC4Bhx3u7QCw0Q
krH0gPuu6voIrIzQIdXHg7djLI6GOHQfZQWe2JywUoqRW4EVdLDd5mY5TFK9YEsz
XlJRSqY3bP/EA30ptfLFJgAz7VZ3NFVYZs9TaOFdUlimXzs1zd8r01kdGFYPI/R1
H9Qbgd1Eor2cVZUMELO7/HOjUKvuOMfrb2eVIcB6ppSJf3W4i7Pq4yTrrxuyWYBs
wtWG/xWEH7KZS464QaFG2DRtUoM6bB7fwbQM7Z34iotwHFArseQmtCFmADSTMoG2
yQpB/Z9rvb7k3lAb7oSad9PJfe0bIJw9+EKoeNehv5dKTGXF+0VWy8E3N625wrxN
Po2vFG2e2E3oVFXFS2u8U+n4SW8/E1tCUmnxNcfeI2u6Je+Gbci0GNWliy0WpKUg
xxK6WlTRJq6baWNQLxIk03ciknUXnbrEdixLWtUt0RfDaCmBRLwWPU53E//mIHFw
9N9x8ImOxxslxJL6BDE9DddcitjRFMMWflw/1u0nQR+9tTPWXdQ18QiUH9zMM8cy
VkDHObD0KPaP3jGAh4fZxLjcjKNpPcJBk6Pmv2NB8QspP8MwnD/QmK/9ZgMGqeyd
trw8Xub05g2u83vm/SZ5q+tRYlqhj+uCS1xVywqeA1shSFUh7Wb3zDNAX03NyrR9
tUW6iGoex94ZhXjhmVWKetSBfplPqD4IbGgVRTMjSImZdMzow334AJq/kxtU8SIn
U8XRANJ0RqdjGHVY5zQVFZSXU73kZf8CDnWzxr0VXLkEQ7NKLQgZ0ujytmFzdgYo
gsicw/jMw65V9YWITs2OMPcWcsGHYMK+mBgcGWe/Kp6Hl/TsE7u3pYrw3EcfvJGZ
eAWMVxhHbJ+sVymfk/dmHiSdLh6TFguzg9glCKi6BDPDpifitrreE0Y1CQmL1vBf
dnsJRNB3Od213xFCzbzcRWnDRUFKCywwv94Lc6iucsNHg5mEUcqvd7QIDzr/9ldx
D1EZZroX/kMsCBqh0ZAfxGxmE925p+SFZot2AEmok6fhNjxz5MJeYS8ZUi1NL68L
QxZGWTdwZLsVsH8uN2X2Vikny3bKdGNeMVgt193Lb0anSMHzQUgIxb0OwpXOd9wm
MwrX13z9a9Drpjj9nFkdvSqQMrvrjZhfwCHyPFV8/HAJPFERt+IMiNayP8MQp3y7
CBacMp7A7wGU6KjIROHtFnp1yt7LPZmTxhTtdp2iuqBnRj3IE2y+PpkMYKDYMsZE
DS11Hhg0tWPOexUU2UrM02wIK/yEyudI+dCklxjg6jBIq4riwdk556hGrcwFM4kJ
qm0lNoWl515zjFU2I0Ez+FCivYpx9J6zTh7Mi+bLYQVnXR/ZpqDI7mlayM8sZw3n
zDXgA/B5C2qQBzJwQj3rKFMuGcJM1X+FeN7fm1smqr5oObUJLQFIt0Hnb4APwh1y
N41hQ50BH9uooksXcCM+311oFbZyqnApLTizj8Nkq3BzRp1YL67qnq+HjaxGUJam
oySZTMHmDrVwnYd6tPJRwDpR5oQPnShKe4WMpsGTxYbkVM2bPKMAv22uHkIfZqTg
NMwMj55BUApbibjRqVx1t0UfXDjc+UOLJ5Mk15GghW45/ZClsBXGiIEzxaohaifl
8R/f77UfSQ2PAv5kWiZSN9KOuearamAVRQiamDaIEZpYC5jR/hJ0/jVXfPb6eSGI
fwcKmTnteEVA9S9wSfo+fJy3DJQ+vFnIV/I1z/kbMiwYGTNQT+DWcX93WCskFssq
OT1B7DFxLCdhronzQqU4NLL4Qwr5rcXWPaiQVy5gBFyOKKMfwqSsNGI7Qoe/2JHL
kNeUEhj1AV9XSLcS1guTljynQyfekrRbhufzQ3nfRP/2GpPw0L5Me4zbaCKuQLU3
Xq76/UdCp8ZzdHlXxPZnqiITMstTkxEPAN6IY2y4Jx/g+IT+kTIDSoJbXyS2tgrg
y8slVVZ8XVL2niBSEY5yplYTuUF+kVo2qip7sq318VPtO6vp1jX4aNDhhvqYoJ72
bvga6dhA1QRyS4s8c7qxS3iGqkDQilGwMRIFlQISLoHGZsw+qY/3SLvq9OXhczCi
R+pAFJFDM22XZZTO2/1ftkS/jLZ78n8wz3bdJo63klzllrlGmvkUn3YgPuqinewq
C6hZVjz+up6duUYQxz1j1eNfi3wW4miblfXERsrOs7PrJDDbGpavATaFr03KU3qR
UJd2v7ZKddureBB7ah1zwE8FADfBKE9X7m8Ig++uW+lOuRD5PFkUSIyiMgJVjgep
0Mzitr2dgs1i8sQwU01XUL42+l6opWy58FLMJgGZgw/XKlWZWV6vRtk5XGyMdldE
WncT9PnM49SLlRYZA4CNHDPvb/YV3PgOkkFtNOdQhE6VuaJtY8gclwgFtmScCk+3
BIZbvxEOZPZoIKiANxFOuuYSVG6z2jgtBoq2Dm3aXrvbLgupsyOMdmzgrbD5q2I9
0lDBOUpEzbcjfbEwo7pqbIucuD/q/bG4XpEAgFeBCGniozM3vG/rizkNT0B7RaD5
sbBgfW4om17Y0Swu9jRLOo6UW15TFtq+kCErLZX2hn/LMd6TupUHXavCpbr+Yyew
JYXyPgw0CKu8sgIXCOD8AQKMOv5CpXEDQXrZIJIPH8TCJEMwG8RQWlm1RyPa9FUA
gkOhv3oGyp7hCRF2eaK5vTPwmdV5yqTUl5nLab4mMUg0/n3jvIBDNb5HfIKZYhAW
9g8MRD1UEFatJ3nvFLPDhzSCSSbaRgoT6GpM7hb/hFHrE/bFsK0KtLVYhltiwn0l
simb5lihZx5+jCIDBop+j+SisOOuVIdgmVeNPXGgkjCcG4mAuKpELz2P1w5ZNlra
O+3cI58CwplumqhAXU7bMGgFmfNhu8hT74H1iIU1aGS0yHZ6BUcVfSX0GY1P+QHN
P8ehRUEQFrdhCHRD4A9p73Q2qWVlXyBh2lIvDgV++JH8CiBiNQAgImO4oOXS9FbN
5Bae6oznQDTck8+oVA0gYeBEi9DgCqqbPZydD1xfavl0s0ePEW64BbJExpuLUjEI
hKLX7CKIwa3IALsb7FLrHTZRCAuEFGpRVsqvwWd4wj0MNCT4hJGFG7nqbTmoBHjD
5Ady+r4N+yg2QSdAB2t9+sfWJhNqgQ+M777i+RSoKxD9+Yhl0Wt4hnxWoFl5K/Ax
nNFwJZ9aH5HgSv9616AW8UDqHM43xT+cybQDK2FQXEdCTUBD4O1eBQG10uVSCd76
5XFQjVFOlu1WLzbIxVcoP1gqBSfcbuDf60kyxRRT4htFtS+uKvVQCMxDSGYo1wYA
d3z+tj+cicEGl4fiV+BTstaQF40fe5ANX66t5TR+CFxUQ81cHBZiW14JtGXq2ZQj
8WShlThUDbSGByK1gDX3jmqtpk6MbNxBboTVhXrN73M9NzXXBCCAJCXt7Dggl3+8
eUwWKx43VU/BowPkKMWvDKrm5Ua2nk4ILS7CTPTrgWy8YvOpoYTN9LgNj8Y4kP/Z
2N6hyJL6lR8K/2PREFMIZiXwNSbJzWIL1Rpcm0FU1JePVrC4nC3NiPWyVUsCGTZI
kwRyHB7ScydPGmpA7Oqlj8DoyGSKgXOUsDVs6nKLAp2ax4ZPbeWfIATxFgT1p57w
mv0mL0VZksAVBYU4i+HPDV4zEzPEM0jfqeyX2ySwztBnTAoqLe+4pYE7QB1z5nTS
geCnJ0YIPrcErj6JWkReH8HTiVcJu7kcVEscILfD8o3R1uoSFhN6M9G7fMQOX7Z4
LTIM0ncvF6gkXShl9f3An4rNFC2JQi2hjKCMlmau4hujwSlJ9KzLdH9EHBFzIOEt
suFKRY38jDjZx4/jr14jcqB5ystpigBclX+nwCydR4cfF1YI/9LuEFV7CjWI7iYm
EoV86K4yaCPp6Tq2/S685iTwioab8sttr1fwSpPwxkS8bVDUQ8xK/Oel09wIXDQ6
TQTdOvV1qKOpCKoU2MfypM5wpy+jMB/vX7yPqr+p8VUbdb8W7/qW7QsD9AHNiJq4
k1Hz9unPhQPH7j3e8eip4jQD35Q2jDSnW23l0BsiBhAceJJnF1ieM493Z47aN9Ej
8InLGibKGEu6ulwgkO9yEE6ON1Ekp26yy6rU5TNdsR4nqjNvYnRSBvIg8Mbi/eS/
kSRG0VWx/MI7Vv7kInvkH/Y9nwedc/hQb3YQK6htWg9D9TjisF2P7wUiq7DrmI0g
YehRPwm/0qc+blVmNoY1UdRRfIpSonhsSeryuIk7hNplpE8C/hREJmQ+vWAj3NU5
r4BzJBx2SPvieUt7ubP+Rxef0xdJxQJyRc0mJGVJDXmKJqSPp7pZHEDFb7g9oE/V
kzWPMUa0vAA4gVHQpxgRfF/N0Ny4OY7/rrL0mnE2y0BS3Rem9DnlVjfek9t9gPtI
8oJ0K2qEXMl3YcYQa6iLnzzp3OqMksHMo9b+HldrBubpT2fcbxKzHwsHLB47M2BC
gO/l1TEEAmul2f6LpO2Do/vu78zIPOm8zORjNThEOIudGPxK+xDzp3AHLPnIHTEm
RrUycZ1dbIIwKNhLmTSSWInQH3GONpWpEWuT+fxRzXpsWxF64wSQFnaeVTHkNpY+
11Ez4w4xBl9rGgtUOXfXS5QYTtKD3oYqF/s8hpD9jMmAuj2yI04cUuzZqH5cj9S3
FljFceWjkk+/Fdy2faaHIDUbnlQ2C1xBQJqoifQE/ffSJO+kTyWmmZwICwcnS9fq
eK1IIDsug2776qZkMgYObfdekvBrPnC7hapgrVVslIa2EbTxrJwS/X81u1DrjUtY
sxr/UjpG3IdUEA3f386tRVsKWtWzRTjcerGdNdDfld8RJshhktHiuUUGnXZFa8ry
hETNVoleQo0dl4O1xCAEmIpsiyM5nCCwRmyKGd1WgHBBEJM6kg1bpg54ehrWQ48m
OQGh5MOJJ/A8MIrCTkQibdhM2fd2DLiQbejhdVUYb517iB/4NCtTkDibSA50YpW1
WrPKgcaxsJauDCjfL0tZvqXSMIe3xwD+KEVe3T29XtFZ5ZHdpG61J1bHhrXaUKgs
SV9z2ZjcRSkYe2fhKdHejdzooxPUwOaagQZ1ECGzS4VvFAK1JTtZ3MYKIinXGjpO
k8V9YcdXPeDax6majnCZK23tewJEILcbTvqFW92L4a1MXEDTs6UQX/Jq2/bsD8WD
+tJMoBa1byKlQC/uohdasbCa5hpDz5t/tl1N4iqFALQTGF26qwfsMFaCy9EZt7Tu
/k0JT93a0blao5NW7roq1h5cet7M88IvTbSEdKeAtdTPrkpZezkbyoH2IPCIbi5T
Qxo5R/y+0KVofFQE7Dn48jBtFRVZgufLY8PVmPUa7w6Fa00XyryhpRyKrIQyiHyB
jaOwSMvatZPMLM+s/5s/UPWaYh+Bg8R+xbsYOjG5581qWNI3CZwfwZnWzxRIcD1Z
UpBInLq7SWUBI6HCLB8uF+fc1w69PGIxLhpp7+qBD1yJ3XS8oWco109qRztOHOSO
vZH6mhiD3O1kVljZHmTZBLMH4hvDAN/wZmHF8OjDxfVGiEwIRMjY66JAo8ZOBf8j
dvDZFOQ1cZRVg09iDo8wjr3z0NCjjD6g2RnyxzNPYJtjTMfDo2QC1PDhL8iZUiD9
woLwgdN6gFavgKMNhNhG33NSVjs+PbVIObOrVDC44ujzmou3GlouwoWpBE1OhxXr
1sOWWex4PtXVXXy8esaLS9t5igUYxXbvRP+QXnV++bwayifV3+nLOpjnaCQiyYZU
vssTZrgUrKnOs3PCTjGycfj7yc0kCj+qyzAitlmhploNnjD3hEoudsowwceTtn52
Bi/qFyZVgwRTuvRsMOFYHYObyR6TRUzqhxZS2WUVYt2M9QPP7SGYd+bvhQfmtE4t
tP/u/opsYGUWebVjtPEmzU2JAfMzi1UTiWe/P4twCNO2Sxr2xQ9bdiJc9uJNCpff
LJ5iH8c54pZcxtEiqM3N7eeAYhhlkNrhp8iG8TmA6uEMxCkDLWyNh+787lEyGhZ6
9Y+N1GwMplIvbWYMG3/aQDPSU1YAHYILyo5qLURFdCPseZjChmHKErR3zA3cjhdn
70Bh+Zj3y95tm3HPAtDkBzyXOFfjaouzd8mgTtxyOjF3tsN/UfiJrSxt1NStv1Mz
widK23XrU4vu4FRCwRfCv7bgt66vAtfj3NNdo5YrXhs9LVeQVvIxsvt/ToxwwnbR
pkmdpvuzJ4A6Bmw4HIIvmOHl6bgkbOb6ePA8um2bSXADZb6ZE9Cb2+bQ5dtkKoFU
VdrO8cCFTWUMa18jdAvfl11NwpShemR+olxN8YglMMZjKP04ormMTx3jBsmykTGM
H4FhN7WY4YFUs5fa/KW8k+HcgVFXs+rXP6f0rY2jvWaZoJKNVPcqqrEhaogMWwV2
wNzM5tm2LNfDpGNRSOgjTBwW2WWg16gU/h69ieJCuJI7GhhxXtooG0wGXUAOmnLx
5t2zwZC7Ki3poT3LT10H0ZKYsiU2Xv68z5+qm0LexMltolVsbF4Xk4dzGz+l2DE+
k6to6R1zS5G2nhs4CvvzpPCfHaq7NkN87+c4SnOnxqHR21yRElJKtq9mujMZPobo
u0mHCTg5aYLaeBzzyvlcJKCPyzUkb/HvnMLXL5C/r0n6FUjB2RZ4VRPWywIxIdTn
PoVtNutbGUoIEmI7bbgUhgX1fj1d8t9lGlBFIkdvSIJI02TArEnI69ME+6QzZ3oL
2fxEq3IbX2xxATo2M83HGxgPBenUfsxu14kq6+0vW47Z/FIs/tDKBPJ2DVQTJfHk
iQg72Nigr7auDFyhEyjycnPtQuwH2Ev2qG9nzWqpsD8kppm3u+bpvwVP24swSN5b
LI7dK/Sf34K7pGMNTzPRaOsw5d6SepwGhFUmarotFNo5va6THXdJy/p9o7X51tjT
WsSDVX7QsoqtzQp6FJKR5hfirxntWZ1UkQYjP5ZlamjmlyfI6M+t3ZU/xvDlc0n7
13AeIRh+Wayxw3NuLRGYIrcIsZP7m01ZqU7JcpUbFzNJGL9Y07m3Acp7RA+op/2G
yxNgEzXOxjLRFyGrgzAdSICUHA54W9Ji83qSY0h4mu8yX5BuOSs7UnfX+yrvcu38
kok1z9xRDKEth6w4rbnvHRPgzHWxy+VxFP0seCNTcKOG6+yOENchBZO3o4DeN900
F6ckymJBS+A0LojMdG5ETvPM8ncy+4RtmEWBnm9ge7kYF7tjrqa3eXO4aHpB9JLd
mk9EyPvZbH0Byq4ARpp+2JLwmcaFP7OaGvgC3GUIgy8STjrfMwNds6DPkedsWGSi
9lJlNo3c5HYVos1RRGw5GMpN84DAoo/EOu1PXXsXjH0Gz9g4acTlAxatF6ifQvcX
mp/9lB1T0bwThRmsFf0BWYotzKL6htdBZ0cSLP9PfgrW5T1F/vFE4fBztWqJa49H
vucJWDTQo7iOc/+W8NKbi06XhFJPLt0lI5kQwUoVxm+7xLSMkFkRxy7G1Xg1UaE4
KpZ0kgZ4mqs7hUMooL1gK77B122gQzJVkqc/yduVROAZ4yzxUaOGrRO3sgPGWylF
RBSqOCK7JBBQscdu5SVksyg+RV1h73Pkt0/Pt9cRd/Dca8/bmYTaICfoCxMJgJkG
SOQyg80xV8Clvti8AzJDjnPTZEJHwEoN6YidkpHhifSFO+9Dx3E2Q4MqdtAhRe6o
gOM3xMd3pparhUGDsCnCApmS8bYCZ2ZPSsENHcwyqqa7WrIZc7o+Vdw+0RWilSZ3
RfByvnkO6vWFkXby1XpKouU0tqInSTdhNh3jXgKVw31Y9d5dqT7t+4ubtWJk3squ
xM9geTcVkHq/5VrMITo4Mvqv++h89ovsDWduntEwVhHc5I79dp71PBbFaG3VZShc
Z2rOH7veXmIxfTI3eKs3vMRXAdsakQYhtafRtlL7yB9WZdGUjINCG58k/Fw8L3F3
a/nl9uAsuvvXgoveL09xt6oDYxGxtLzCMT3PIsp4tlKMpLyPNPOWTm/oDxp8TTCd
1ghktemW2F3kZzn2AOPXlsy8+j+bvPX0nne8jspWByzebptu0zdVk5OwStHZUKRx
Dsp9zSZ1qK+e75uTjkk5l0sxIySKX0JKoM9iSXqd8MnAJxS8/m/mV56CrI+ZuFIt
MFwSpdb8Qg/Hlp1nU0gkACYMACNSplCS+sbKGXnbs9SGhd2TIGQtuMg7R/hafSsA
tJ5MHkTZ6C0LUKPERyqFhi4+KB78poAryJjaKaGAqHoxsP1Q7zUtY7Dc6OVF882u
0Yw+tgZOrEOu6x6l+QfnriAcczN0KKLRprfWFjRuSxfVFKp8qsc62dYM6Z8uenkM
G88BoZnIt6EgDDK3zvyuAO56hh3hKEzHDg/p6JjwNLArrIDQV1VePeZavAEXfyhH
kaXSO/o0Plw0GZx99uf+yMCJAOh9p7kiBkL9BBHmPqn9ttW613m9tIUFNkcTpSKj
gYyFIN1pj7HIYhMgJSh+MZM258rEjgExzoxmjt8xb3gaKCKxMLmMe+W6WGpXs08T
QXu9bNjI07yE73jog66fX4jnKZfEO1ZIjef3zZ0cN49G/srs5m4PqIxv4kJDfzC7
0v4waQ2M63slGR1LhS4kN0COjOFf1C/AGzAIvvKnYVZUJkE7Q1oZxV5Lw2Jfokan
VhWmGtTL5eIW9HVvPzKApSWKJS3Q1Ze1QDA5bxiQuqFr0l9DTzWT2UwRpp8D0Kvr
Ii7lHEk5m26djUe310hYEC7WKtN1JPrbhoC3u8lNDGjJxg08U+YmfPyAHEQ5mRZ9
DEaCO68jogBQg1QJhsnQCNySO89lYU2k/M9ZSs5u+n+JGEcDmJ4PIutRBoI3qVCq
SzVdWoRvsjCzQ9VhYCmFkIVq6Qbe/dI6ppQ8D/qftan+MuG50Z9jskGGEZUfiEuc
TLTZSlRKe/TXdPUSfPioNrTP8Ltn8GEilZRazErCg3GIJ/UtZYUwHZAsPRifLpMO
dZoYHm/PRfnsjAxK9hBcFwLNS0bHqE8+F6vJaMpbOq1xJNUYyYA4PSGAZtKhG76Q
iCKBbhzXyrS1jzJozQhZiCarZBu0ihWGblRNOskB4WjqfFy4WbxZJnf2OPNc/ruS
ZnmjEsnwOZHv53uZLnmBpHkRmi493XONuljumGxFh7TlUzPYT2sAimajbPzl0IMy
TP9ScHAtP/T8dPgy+k1/Xmwq2HHAcri8+tATD5EnwBuak/Zn8xygnHDq6L0ZieQ0
ItUM7kX+JmNg5mZzkqcWZpOxfuxH8ejuPP5vdSxUgwVcIBf04fknIAEyzVvV1bzE
zcB5R60wQOnIc93PIVIJy0eLiHc/QZxCaaHMeqMTI/BiN01NbsD3wT7uGmiPpVH4
0puFQ4OpLrrTvBI7O9Ox5ngMH2R4gFlDTuXvooGqOcjBkU7sF4pPciH9uLzRos2y
lji4jfEYTksE2AmEC4oXGp86e0YiuwTSMsUjU9vlh7SqJMRuoFbIbpTNitf66SkH
tybEORo2YhKIVfKNI25e4rclTbSljQwowAnubTxHzs0QNflXuBjbViLnc+yHrYXu
b8On+PobAq8I8ppzUi5FN0VzuJta3YTBSRmdasutdg5xh/miFy9rtfD1AKena6YQ
gban6yeEjtL5tY3Vw9qcFHYnQLEguh4amD4+GC60xmxYDmAoHbwcoS6NI89dvj/z
PVQinCNNqvKdERb+CVB6t+e6PEw7c1Ml3YGt7uqBkV1OqHHAR3TUxwIymjeo2Hzn
n4PNaH2nGUSlP8jgNPzGLg8kQrTECTFRbmwubiu4oWH4DYqw2lbdESJe1YPB5whn
nmdpIOL1hGeohDZpOXoBIfNhscLTXWSmPwUdJ8/zKacKSxj7TFKc4Ouzx6i0wfbc
m7BY2a8jmSfIUCmUj5rdbRjAUaS/oOZw8EgvLlk9yZIqRWii7cVfDD212zTSBeLp
aZyC0wIZhHxHLi4ho4IPAk7tBP2rmSNjSlvdmE5DxU5Q4sxhvSIOC4qkEN6Ao5V5
IfqiB5qCTAa1VA3w9KnH7vnOQGy84rbVe1Xn1sYZuEyNTPb5UXjENgNdi6PcUHUv
Liy02AD3qWGVYbbs3/KC7fjyQwMw1TrCGwBnStpnUJRsVHfH7x8wjm3yy5/ol65I
vjDT16SU/MbtF7GgPsHvmiCYhwUSoVodYNqO/B4ipzraZAYnUbuV1W2BiQIHFZZ6
eYE56khlztFgnUj3oOAvXc4159w0ZL5kPC0yWcIHKfXGsDwsZz16yR8kBnqu6lEa
4SZ159ORbBmAsqzK0auUUhFAd6FBmRsfNANkgjKS8mMTiVIX1CegT5gw8MCzDYAI
+91/tV45opu7P6gOLAmzt7R5LXiHn0z6m7pVoR9bLIppBUyZ9VAkdR1gPRye0fyE
LPNMaPDkgO4JCDDl5cMkGISckhzPxbf0H2A2t6t1tVlyu/diEjLtQlRhZ9MQZqg7
NjPfXwnnqbIWxPoUIalJCaJi4Kel/tmMBpENcIuYAue+tttCONhzihyor9vZpM2R
pOaC70zJXyjSaco7KiRJoN0jR5sGYPtUV0vexK2iWRTP+xyvlKceuewxjXLRgOjC
KLDkO/QDiz2rgxRUMeZwNQ+ZWjZMEUjC+Njr1nie5xxO1e11F66w2Ex4CEkCZ7V2
EHdWa6KKmF+TlMeyy7Iu7JM2LM1HJo2eXpgIGvGMPAUQ9GkFGS9gdXMRyAsbOkWy
tloogILWuDGsegeEOlom/arY3GP6gyWO80lCNsHHtaX10s/Fzy/ilvMWELsOX39p
+S33KmPyLczKn3MRDpXkXsI1v+QbZZMGTu7N7OGXw/4kKJUeu41iZgeC1fVoDJUH
kSMXg2WUeKqLCcqCw8vf5Gouigu8IYe/ss+TbscC1jI9D/kf+K6DltByHBjNNhj1
LOq04pVZzTqTnXYonwuvXCMrXID8c+VG3LWJ3DaLkksxalmhpPbGUiVmphmwyepD
1h9UXymCbgsnaFLmrexujY/yqOQsDabplr8Iw2iLNMrj2XY6VN0BJh6oup540nQ5
PZVSGni6/H805Rl/4mvOOCBsmVIGlvZY8aTQjKeDNJNG8PM9SzLB8dW93XkNviBz
/ZaIdvxb8/fHf7j5FadtheSfAOVD+/rbilv++qAxW2XnKCTSUpHRujKJhSBCIJpo
X+XZ3JL+MWS25QzpjccejGs5VQjkXFTkOrUbw0p9A3AGR8fMCPhPGO4karp2Z/2z
JJGZeUcc9JMpR/MZzraIvdpiF3/JH4MBnZbTritiahBa9HcWfsE7/yXPFQnikCYN
9Rag7IZGa4EnNEJcL68FVARgoGtKuJnorIJn6p4tuXEzMuIFDQM7aG4hkEXN/Zsj
aJDIXw1dbHXfpLPt+rQfSPDlvPGq7EZKcjXnRQd22YoMXCpeclLbDXQLJiwB/eNl
OLlwqazOOKtc4fSNeqKL1+J2p1/UDYrWQ+0QKuJ0t8iHxxTZ0N1E1oxGuGOkk410
iJNcLgTcxdmNCZzZ8BohuO4m11WK10enkwYo3GynxMWJBXVSliy6UnvqgsAOTTXu
SkrjoHLg5nt07xd1982wAxhfFOhiIuR9aanwC4lrVfkYpSpd8rV2o3mBHcTk+IPF
GO+3b2MGyX7VMf4Ftii8F3wD/NAvNTU5jTFyr5H5QeVRnzNiMO1gHak4MoYMtdp/
wpq+SyKsvEwgJEwOUl4J9FSubSVhrb5mvLrb3pjzJFz3G+lccr6N62L+YQLt5Tov
+y6Fct30+ZQIy58JIv1XPtv/MJ65oPFxQFlQVLThfmgWR8g6bYi1QI+fZ1LQMMQ7
iG49nNoppkf5NTzPC2Ha2r7vGDyaObsgWVifVzk1SMR1U7Q2XWyf0W+J5Hahbfsv
I3FNKEPRpYsUVE4rlJZFpRiHccg8iJtHts0GZrf4eepRdvnugP1j2hsGMxU8hUcT
e9qqWRrhuAPyTu44msUz4WlbR73lIAwEl1FpACPn/jRyMjY+w8bg+d5/zCX+ZuvQ
ur2PKnyrvTaRa15akdXnZQZFxZpwO9RRc3bnlYJtKZyJSBc+ZmARPS8p3YdSGfGh
M5HvWj9SvmZGsGG62/RfcujFwKuZxX4JgmppJkLgofaMb4cs9+/v4f0w5PVp3VYh
cfQ6O0bFnM9U/GOlPHJE6QXP6u3Wp47MSCv62jsHdLjKTNnw5Dy3uX/wCuJMi5FR
S1TASj2H9ValHjsH/MUS+yNsMF94gjp08LVIqL4W8+JhCzwJZMM4byX8K/wbtkHr
Zg1ACNFrRIHjITe5D8UOawDXJYBr2JaBgQj09JnH1EMMLaErYr99YRl4UsPLbr4T
dRjT5OHyXcibmerdJiQ4+ESzKI18vZzerYzpoSfsPz5BVei8S6EDg8vhXxOO6gkV
lF3KTAhQAR7Eu/3w32LBtQ6D0Mt7HqUsAHFUdd2HqMJ/gwnxQyoqnajBEiI3t7Iu
Lvto+0Mbb/9ze3DBCV/JmTI/2xGY9Yc62qTOOKKOaei0BR0VEplWFOtNQ+zfnlq/
SKwMELCNDNS/IyIKTDehDbT03WHo1W5fE3pQbGcOXSlW+6D/kYuo+RW9p2ppFtkN
dwun/og0+MqnrVO2FsR4gEqPDZ29wSogalFSh5cIQTwO/vUxWfpUmdFe2hkEG9pP
WFM5U7olzsNZGnvm0PxN5pDJYj8WcVQJGwHpevZpz81lflSV1bTpZPPIRXp0b8wh
3fV27U5gkBBt1fD5VAF/fQnBisbr28WVZYqreAIoxhASBz7vSR/aKS41o0qu8hJj
sO91aPvKmeq7HDOw5IkCi+sZ8AaQm3gVl9QNKFvb1HdqNuM8WJKYpAp9FfJk3CmJ
XXzEjcZ07z6SQBhmne9RausPty0NbakIX0ckd8xH6thuaZygPsZyp9SUXfDpW5ls
usZ7fNG8L/Lu6Ixh7hGFC/QQ9/8/YsMNB1c7h8tlb/D7zslezUMajScLZsJ4b/gH
uqzwN9QZqnPPnLZfPZJWr9MYhMgPwTqsItf+Tfa+cjQjwOZRIqaoKAM2VJBpHtP2
TBeyOMZ1HLgVx9XLXWoc8aSyq44K4jvjchBW1jb+Hf9NIovnlK9fH2UZC3L4W9Of
r9s0s6snmshi7ViEOwZLLhRK/yqNriRvFiqScjydHLXg6Za8bEBWmC35QZjZw071
W0z03S9RtdZXwBjF9OlG3K4XctV9yX9iW4CUCixB0zv4IcrCOOVFDF6jUIIi2jyn
hVPL28CQq3mrVIWvGCDvBP5kNMSpNIMIhDeZHgm/U6yZR7W+nculNdMpnNo3hFgz
gmTjQyzDlvEmZAATS35L6Hklncc7YHM6rA5wOGI5jVxMpCVZeGyFUhLcvGbkdgZo
o6n+1MCla5ltaWhP/LppYADNlPPwE/7hhqsWpP0lQDGuFRXy/T2fIJskdqIB2V74
tMRPgSrGGzOl3RG3WgXq5Ne+44hYIGLvOWbTWDdxzh5X2GPCcok6LEyBBTA/GWsL
dtjESlrkZR8TmfHyRcyWLq1tVVANyWgqkaZWS+R+dauJ5nL9Ao2yV26n1JkzeFo3
oBXQlN76D5oyLCV2PFnYS/n+owWi5s+7NY1dbKRgOJHQmMcEckrAZjHBb0f1fudD
2TnajP8/tRbwypz0Ct2ga6NHkOSSgLl+kPWB23UtE01Jb7O+FCa1AxJRIQclve7r
k1Oxaky1Otx9440kbU2yKppr8V6n/+BzCPMfj6Mr4S0ffvnjQtrcbZiFwQpmPOtK
FoiETwxox9zSL4kEDIb9hbJUntdw/m/Luf9pi0Wxp2HWhkHj89zgrekTl5JEgJvY
hNdWS3b6LIo0qK0s07mhuy/HRCIhNLfYuRPbHnOvNuhseC7mcKnVzm4/A7dUP9Bw
ZI72vCCvpW83DJM0zmOL1HVqoXmQ2M56zNVMdABct46aIq7Wm+zdH0gj/BKOiMC+
02zxbBWOcLt+NHNy8rYJjnbkZfQKhrBxjDbCnAaRnH5AB96oJYeQ9TYCtYvI5KUW
dBactoARXBNzVGMMavWhtCiBYtnKTum5KhiAI+VsPo5Gd98LMSGFFLkcFNRVIxPA
03hNLd8F8xW7chOjZeZDaGm2RoUiZoBefqJsYZWbE/jxS2ceiLyDYysCXSaaBmz0
33ujayYYEJptaK1RDK34+ozUL5Npqm8XImK8oqIt7YruAvLG1GKMIVheqjjG8MBp
idN2yheiLxBgPVd+s0SeoQf7A2zjdc/FvTSTh0oJnRMCvP0yA25OpFGPEVLNo7JW
0KSbKHC+ThDk2qNEf2sLi4vE4yskbKPQ+cYvcVfrnd4VFc/5b31Ejr46CaTndWKX
ade5oSYzOwQD0hj6a9rPDM2lvdVAxKCI2SLfPMWiV8UGS5h/K0x/UoeNhlrUKYNJ
0hiYdLBTcOD89McePw7sQpzv448Sd3vNT8cDB43wEtIX7r828bAHSZeJW030TSC7
oEssMeTsJAqjI36+6gI+DvSum5qykR7ZepHKiq7QBMZ3ZBBztCuJCw1XXT6wxiqi
W5myyxlp76ZDAWVenPVJJJ6kTJhjPvV4Yj7nJVtE7pFSdaEhYLQGiOP7Mh+eHlJP
2/xPNceaTq2x6wPecvGriqzrRE9wj18egM7xVgC95tYSmbAPEsqEJmO0LnXNEmDI
cmrLRJn/a4kOEZc+KjGanWxd13yzCteP1GgaZ+JXtCBMt++Z5iihjJQ3FjOXXK7W
02aj8xgcRYYe691hXC0THKCulxrZLoZoh5DOlpPSaqbW4HX5cjLuhPIYM5NpxGVA
ehIMnAYRP4drxh+2TPS2fDVkT5phVFA8xj/X25d8V7c8Lw2wfw/u5CDt0Z4Z2jFR
NoWHg7LGTJ1ucGdkdJemicLoJoph6IzjLHyA+sWYXISTzk40fkweTIHRT0YmclE5
8TNAK2/1W75/p2lpjOv+LnXjKoNA2BX8r5djdu+EPXdY+LS+GFAIp/DQDVCKFtyy
3EkLcjYcIokgYoN8A2Z+gOFJF8JgwgnVRFXUZot/nG0wlPPMylUXlSSYZeXXEoHL
Z+/hlTi1/vstmBiX0bWo9WK8NGLlqq7OtbJI/Cs3E8NFobNoS+3WPlU1UWK+VRvX
QNYZeq4DeifK+tUo91E02lKXmM2MlDQUrT7SfhFyyLJxhJ1YmRe1IJgHSRZGwKn+
a7RxiucRrbLZ0gbWSOv0huTd6eq4p9D2wswUIL3NTok7hr2WaS2ALzqq1KkJ8sMe
eCoybrKNLKGEPAjHc946dzf8Sv23FwLefKUGAex+6Hs/llrnjOELm3QLN5Woi9Wh
8s4XzSlHGDxQVj9s70CXioAuqGPzqL2awc3aRZ120fFm4bHOPk03M5msU+TDUxH8
DHsopWNfXbnfaFG/PagL0pWztxz7g4ULsZ1ya0MEN1a3iEJ4IWf1IoFlCipwH7Kc
NvX+6DQ6pv5AJ3L0ysppKOLnWZt259FgeAsy87M+mlISo/onPI4VwKqaKkEeh3Yo
HKtgtptvAYY9JEGQhk11eIiluxnrATV5S3sSVUXWbcU2f31HhXSZIFOKICN5aJfS
G48vLF5qAxp4ZucUHTqD9qDchahIEcKKc79z5okibtF8M8wFDJJrquAGWN664GNK
sEOczNJ9ThJ8mhpS/x283W1l6ne81pYbAp3hnYF89uC7Wnr/2SDpeE+LXjf2XHNY
qq/6crXCNA4hP9ULO0i/dcqE0dQnNiOIdJ1ybI7YrDG48bFp+ycPZwD0y5DRtNA3
G3R2mAqHeRk7ArE5kyyThWnHk6toozndn3mWxRiIpUI+ZGRxnoWnHH9jzu2x5puQ
GndJK6/nsLFV/BAeXCTpUfLtpX9bt8s5t1NJIGTZZ5s6fhs4UxUFSs+Ixbxi7umQ
ScZRHQ3V5U/WlYX5kC0jf/RF6PuI9J0rXbuzLsv7BhrWaebdIVbyI3IuVI/Kw3av
UO5jUGuMeK8qVDw1KyJRrqnfPwmvYz+G7EUkilo7KsITxDkX03iFE7ff0BH9QCgs
xdxzXcaj8ho9L4/UbkpwudZH2/vfWxsP0/XHXFdFQJiisbro6LR2njlW3q6Lr+bC
nL6CR0wRzyUilms7o7SlTKt0mFKsUI69gPX3XpFjc5EfIfS9vjlmnLPaBEAb6hl7
3LOTtnv1OQiLlKgUIq2Lq/zHAfWQURiICPE5aWVkfhqh2iChy0WB3QJOVZ0oNoZX
i0fKzXQjvU6I20f26+f/f81lkiwY06qHKjA87VUlvzPWd2wsLLZOWdKwHoKYZm9J
Ys7jXwgKxNotkLL8xrluoMomr9GNVV9Cx5VXnKPw40Weij/0KbSlwB3bsHYyFY3b
iSQ9Qngwc1Yn7ifkErCzPUgyLBcLWKPufbtc9SA9RQKS1CmJTH5D7+AoTVgHaMKq
tQTiDhFnf6A/0UjHHKsIfxSmoSC9tMeoDzPJpa/Yh4/JSwGMdW9fVJ+3B86I1aLV
F4QcB6x7JHTeMmFh8XwwTO2s87ONi+1EbakLotUQSzj5yw+5Gn8VDDifh7FL2u/w
Qx+2HkKI+GSj7BZeKeHgnuFU1LZ4a4gO1DQ4Cgq/IdiIxXSxbxO4u3RbarstXoNS
bwRg34VV2q7b6haWh6qgBzaW3zV1JKiQReb3DYuoCtdMlwI0wMZr1NwiwWXkxuVf
Zx4uQwnDAoZ9VCRRZth6+cCDB+sFZRmUNFeCorhCjWrMZrmHD0o9ecpchgQsu9Tw
fxP9P16+IYUQiY93K7hJKDQobx+ic4qjgW8oC6VUpNaLuBqTDTiiWdnbZ+CVNNJ7
pQWxISsungX9Jc6acMGe/EBJtg7FmLtLRWLxjt8YH2RMxXkIrvbFaO7HD3LcUQR9
7iphEJcpWUE1ECGhP7+grPH9ihsc1icCFnhN6NKoftj/MyRU5fZuTt5Wk3Y0jHmR
shQymK+v/7Qg6xS6bmGyiRgPQ7iLhSzcCZzARJ3iHiq3cewpaDe1wJaMua6sgbXl
EPJcvDYIHABBFYQcE3aMBd9Vf4nC1p2zjyswB+i608eSi46o3eGfy2S78l5RA4bs
8SAJMKBmpfAFkj39Zrlv+LNvX4z3qRXQ9SErgs1UWkZhC56llP7ktqIzHtAYz0YD
EjMD0O/1QPPMWOVous2DF9eyt49J47qcdn3J7v8rJC5fPNIQVWBOal1RsMMU9fff
uuXcoeJulOH4QRoVq9FLzMyWckEpwRcFDnx3VDhzIWVWD9yqau+T+12nmBC05WpN
vUO7ZQiR839FQIdjRlhpWeeqIniE3kUZqMqInM3polAXJikwZXloYtGQzimDH49t
JGNKNL1RiTvVXR1wrTJOv7JnThE7EE/PU1aLX0iwlUKIV3lq+LD+Pph/TY72Sl8C
NMyVBSUK2Xi8+lj+5TFTDppS4RysAhX8JxkrXVK/OqjzbyXtKnAj9a621la6DEUG
j7quTjLCQtlXZeRhaqR1bhE2kffQkTlc3fwoWVFG3Ylvv7EwiHjQ58i+I2XPPVyP
K61/bTmguL9bWuluDiByjo57EeMFAZtBfiXtOxnXpl71G8qgD5Ecq0GX+Ai9vGzw
lMiajQb2gqBKQVfTvHS0K70X3DgBDoB5+tGKvyOm0H/yfqrsi2oFFEui4BIvGyED
fDcfCxAdA8Nt7tiRPJfgoQK2c9g1w2jBQc34mxSvQxs7jEphet76to5ZktUye6GY
xhOitf2N2qY2P5M8pMQkgYgNy0d8cr5hCW5ArI/OaSMiTayhWerX/g6p0dY/Wf1I
bzMn2mh/Hi0LepCrIho14k5RR8GZWMb9jQTgieuuDSNdL7yqU9DuVjZPmIGYgfKW
RXJIDFi3FXZwRlaNixAQEkT2QVOR3rC0B7Lphv9EzinvD8GdkVrVc2l1aQaS0zoQ
1fiAqu48mJMud1cWlI1vYIW2heQsIanObr5RIeU7bnarNKuiCCz67sVqJIKzQ7jN
PgHtiSqjSi8vRtvfbUMiVNaFFAypHih/7dB668F6U+p1FfmFIkVPTvfMsM1OvJUm
7QrjbTPjsaxuwi7xhLPTjewPc2BeNXhtKvx/oeGe7zW5RJCMmpBo0z3FkL1luLT8
F0jIILWkmuKGSvacpeEMrpC16A4NYBuUMtkweSQ6YoQH+johYMMf0pbh9zsUqkB8
1+Jfx/AcklzJKjrlhvMiavuDw89PxITAGBLiyYZ7/ESnWiUDlqiWZVssrmBMpBI3
5ar9H8a6EniV4dztCOyUKbDUDCRbx6gjuUOdxtm6Lr3pxQAOF8ZukqJIswbWK72W
EaHyFp+qGcEeDaNMakL39Kt3iFk5jdzbgjbR54ekRh+mL0sBR9unENM6YVFUPeze
E997+sY9bYdsvporD1XjHLe7B814rP+F0fUmQ2rMniXEcdMooZSr5isJKtX0imO0
JOirJrSFDQNUP5KfX1yobQlRI2MPNIhY4BlmoUfgZozofgXs2dzqq/tTCIR9UeZe
wRAG9jb3me1/0ORi3EJH6fMd+YoAXP8TnZ4pbqxhjpgUmqAxvTqv5RT1EHy8gIOV
EBowLo/HBfPL2nLlI21JpX0d4v/WavqqFq8/pLSLZDvOwpvgaibTYPqvafp0qfJf
TPfUpilnXfdDRqlnu3FmsPdG19qjuD0f4KUhh2NvMkv3f8gkv6CRbL6nB9oDC7yY
WddAHIYRQQcul4PFh+ppgMPTCwqZmIqtrp1B4GL5HNTo+T0eqn7UEKUxqPsfi5oD
92i/wojy9vN4pMGNFlqy0g9aUXersp5D4Nq1FP77C0zxa8hSiPLI8cLa4y+a7u4l
HiJvIME0Xww94zwbQZcBwvnC7lJEkyLo2g7KUGJkqRcn/8a7jL9mb5qIFayYdh2S
L7T2e0ifCP0qxkWO0hwKA5vLpVgzNdA9/SWOcTIfKS/2zFJW1sKNZjrXmtdYf4dd
RTcGASPs7xApRSh3lk1Ng4JvpPT315syadQu+xogkFS2r2jI3As1KFi638+28M7Z
8s4+w+Rdu44g5ugCCH3G9PsiYTBKActgBn5k7Kx/wwtneUYQAj0zLjwVUvexKWkm
5GqSKMPseZgvmt1LKQo2MpEbkChxGS+1Y1S0kceX+AAVmgKg3ibe6MpO9BW6zEiH
MKkfqrueZKItNbk89/JhhE6CcSs1nmAFJBPvjKMi9i1IUcTtGV9S7oDBJ1FWGYaO
uOA7wwWQvKBzFpeGd6Y2ekX6Tpb1KL2FclZFJXvnGzVaNBaLklumP+/co6BsEdcv
NimXhGmL6iEU8OBukXAlNh5EMpGYKWF6nanQBxhJvDUvVIcqS5rXhPydvyQmb175
HMkOOhtYb6dHSpqSBu7Q1OYbZabQ4SoEwYl4W5QJRiIC34Eb3HIvdqLwC3dO7qXO
MNTpw7jRjr8gbFwkAz8YCz2al0nnDpFuVxDGBlshodIoIUjwj6ft4k1kIT/kO46c
Ma0jQao5bc8FByBjwEEqMqoyGSNYJjUnZocY6fI3K7OsmqHWuHMm0cPU+L2S+xgn
ZisHRlW2ZUvDWAOr7rLbhl7wyc+mhmtR4g/bvMJUYOijcZQ96YMaE9SPgf02o2xW
hldXk7bgvFOyOHb+1SfgOUc5ThIZPjPM4dtNoNrLNMnPfNsjG2TITGzdlIQZLQc3
gRLPjsoPkQNKsSixLXOUeC3Ao3D0Ll49F0MDW+ctHuAmNucMtftvjVS8AWuOv6FP
zfA+S/4XH5f8r5XqhQN1Nd4Wv3grkwQYpM93LwuFmsl0ugsjvW9JtwqUZrBdVp5h
YEhOP9xv1kiLohggcA+yAlp/JYE6wyiqI4VU0MaAauU4VFZZI7vqovRDNH38QAus
AJS4j79RCKTu78v2Mxh3gmjcymTDYqvXQom6GjdCPojjQPGYA1q4vfJn3r5k4qpu
ioRYS9YHIfcDkEDK5wIGuzFwRKf+/7dyjPbhmaa+Y767w26VzOXLeImm/d3/Zc04
XHd34Qy7NauRpm+hLBfYXLCAUiw8sjOlwjTGWI6Kmbgfw6Ig0REUX7U52fq+XLos
Y+XuC5iQvpsu0ss+Iz8yE//4LpPFkSPgJKgGS4xIuV6cEH3qhllrtrure7weCduO
jL/lf3sC6A27SRVrfGe8bJx57VtNt6WIJeoNHiEZZX3w/0gWtOaqGy1OG5EZXodq
FttEMtGxEXmyM0MOTFX8n/vmwaRmSPn7rZ5PjmD7aMYGjSu90p8KHUERwuE0/qZ8
B3IplCyCsB9XOSk+aBytevZNInX4cRuq5CIlUp7gpC/Wu0pEp0Zn2bEJwaWKUrMv
lD+dNMt//BPRbYUDy3IDAmJXBhH9J9weYYcz4sRyI9rWVYRQF7ZEAuyI/3fvP3Bz
e2+OenwLJc1XMP2BgDzJGY/ONn5lFr2Qs2ZuVgvJpWRoaC/TBB+duM3hdgUMWI98
enVeti2rGFwuJ5WN/87HMNn769DpVNIR44y0yRG7BBx4j5AtWzN8ncOCjf9O0VHk
xuTqmdEFOcKUT+Vz8ZTA9ONYEf3EePCWHltJIMji6UmZy/5Ah2aviH9UChuJQVDl
fbs1O29mH0Ey9jXQRLmJyndzZKwWAoTg+gr74ReAQT2xVlT6iRR0E0zHRpe9ddmm
CuOorek6OpV23maekJ5mRMf8NHoAxXKMw7zUXEiv/DRzX7/UHWRNR7UUX9wicVpU
8PF5XcW0NONnBE/O7hx7WiNUNAKaCs7TzPH6vWuGqiWAxafduglyznBlyCS51VA2
LvIGBn31W4Ei1NMA8NIL/FEPEwgTRDHxJS8kl+sxXIJMzBi6GEK/qUtLp5Mnyb0i
3L5C8IhDG8wfaxmvPLR1IHRNVtsKAEbMzq6qM9zftjDjikvVCe1dUMxL4vscRD7I
bHlNy5EeSeKz+HSrquDxhm2ZuY+jM5rZU2zHhs1P7iMQid8rOZagCAIIcOymQN8s
e9n1iJRTdWOLbgKJ3MG/sdzuj6gm30j59TWqJiC/lFuXq3vAMEulgViCITe3NpAc
GFn7SwEZuJ5TasM8415EHpxSrRcYOfq8WbSN82k1VDDOcDRt2u6SwbuCDN9adUzG
VOdgIhhBaOfzK8dnu/CGWmX2S1vy9F1U3wwwvkFwDmHOcfhxmQ9crVjyjudLpKiM
wKSZxS5JKa/iwmWpXGowegzPxduGGWNvcEAD2prP2u8PfhYIAG8dJKnkHfVy0k9N
Jb7jX0lC6XzvBOseb4LIqxmZnFIOcYgWLxo7ilkn/2ulEV8O6xIKnTlc+KrYuFA/
6yhp8ZaZ28AJ9fNqU8QAK9/Fgpms9+F994WNVOmxCzukGkYOX25cpAdurLE/pSVn
KBKjFZCSY/XXEdYJPTtauYpLkkkLQrhrf9EDWwgsV/OsLqi9rwiYPK6yfOyQQXy1
5XIEbsiqNlYn95/Xrhf4TisWjpC4Lu+mkNHjxcoB6JxshkcTSGXDXyr1Ik8/rMa0
wUmvaIhqYTSN7udmuF/pbe337Z3IceM3+VfPCYNcvY6iIHJ38/PPmHFm5xBsUR2F
DD5Bh0p9dL/f1L+mENUl2Ebyedc3ssePdLeMtGBn1mJsq5Eew8PCx0otGZVn0yy2
q/Yv7h81glUp5RWOV0K7g1kfKobesxXcy4R96xtQCrVdRBOp7GTB2ZqWMtlm7FEo
wGvYnHEpmUfgL5THqGXvpJNMHYrsRU62BMLMWMkHgIfWJ/ebdCRSnDqOx8c5bu0e
WFNf47wWTbQ1sK70muMsfvy+YVCom804TdU0J0QEGIEzAcPQvIAId6Vd+GEo8+Pc
Q7TEh/KrJsUusjk4I62gC5kndmzdROy2I4ZxPgzm7ChRxu+YxozbeFzu6kvmO4Dz
9u8J8dbYzUyvsxONX37GpNh/fdRgV4yMOfPEMzUcnUGXQweDC6FELUi9dJ28doUT
g881GxYF5wlj0k615djRG4KvumKerXqxispyyFTOU8ydO798+0EPMA/WBDeRGYc0
JH1upzsynwYj5klzvSwaO08IRqgPEaUH7+CXnmptVUhWjG3Cv5Gc9TK8R+YGWAnw
ODmXZJYyUvaitZEQRUQTaxV0LlJpUBUeny6TsZ0sGD7rbyQmmCNqvMjDRnJXs9rY
8IhGg0jOo248+GjslRR4aWnxSvzKThG+h2G8Bj28LWZIx9YN50hdys/SKl++OtFT
11kWbPTOTCVU+y4vW6AAWvNIV0G8LltHSrryuZ3JVfzyKNgqwkVgEN1BFhcoPAnK
blOyZA/pUp8xrk3I+OOscPqWbBE02itT3TwNcGmcpoPwdT4ObBCUhUtKiS8VFv5S
h5WuG3eNtpdMKftPyiTbneFQ1FTlD23zOU7y67fMRTgz/FCTLGdaaiF2MSqHQL6l
pAAN581deq7ziM7p+HtgPb2Hq4mQXFg+A5T+U9fkHMJ562RsmP3MzmonGzAtFbCe
QzPSMoIOCHaGdF0ss8Snn59xex3cEAhbXXJFU0xpWVrUa57rFMn5W92Y/nC9HNLu
IwvY+vYV287RtuFSpecHu9f3EH5Ks3opjrpI3gvEPRSSvohpXPmDki5vrqI8osEi
CQ0jn2s2FLVGOS76d4kcJJD+/ATHIy2qYahx7NeLh4Z4Dk+xUbJRNY4fGk+hCGwo
AwPcgsq4JY/4poW/YBBy699EMuX5eN0xwVJL7TcoOQOrCHHNNVHqNLVzcltWgZVA
2BlUk9C36IU/LFc8+VUfb7G+KPyH8jo3GsFauUbpWLHmlUG9xiL3HRoGCckpidoO
f007uVgqWzR9Mvh1tVtJjGrrst8juKCXBt+UeDVWQr/FLFkROZ51CjUxznJfWQ4I
ZdlwRfiGSPj2Jv1OXDXMpP4KKmgURcyZk2vZ0cp76bcZiGXBhN2XKWxulY0N3yEH
4h5ZSVM233EdehBPZktEjkD8EFC1Cos8+drDRcelBYctSxUZ+S5DWJgeep5o2MY+
JG8m+xfVS36di/EWovSFKGUgdEh+7UDTcX/Xnq0OYZQrB2EmVGPFPopDBlULf+eo
tBJTof5urJ/itfawBw3jzyVRlcNH/BJwQavYPIkhSAGBBM/ARNCWRrRGnsP0eYlw
tRbSAhAyxWmuuh/Ys2k6U5k+NaB69rlXsAOhNBvOdxPKuRcs23AhXyvvAfZIU+qw
B2AzKaJEC658GpuUmcYM0W6wcon+H25d5IebOdJrjfkHBTVdQ+PWTgWg/nRpj0ZI
7+ndUkGQFT38nZi5zOf/d2uaxhWxYz+C0b0btAYKY+ztVrTjptrAWRtfYXb+yPij
uxA1xFYqbkhHhUUhSTQ9eyKMvtCVQuAFqtTj9xoOvc0SUBYbRr9lw+TRDhz+o+GQ
k/BrmJ2OxuqDYzsV1C14vYLlks0PCsG3bxUx3nYnQGM0GCmelrRuvMBiiMZ5j9og
THIDRy00IpJUkeYWd15+oFZceCOk3XVbPSptocil65Mp0hOkTPnuTZHK7j49baGU
5cNx4udo2prHg7Mi5egjW+XyBmd8ZPT6t39cVLoHc+Nd21avhUkeZ0Zb/Ol+eJJF
gUhK+wJIJgwg781/ki58fM03v00XJOQducaCRMgkuJukBCOL5MzJaHLQL7GJVJTY
hiq7uj1IF3AGcYXaj3ZB4Ux9USBigV89QemSLqlBYfzDy/ceofkRD4wH9Y/PPcKg
n/QqQCmAHSHp0lZZkhW3TgrVjOBuL3q5fNk0FiEvU50vS5CfhKZ+jUG+JF8pU/nj
HYQIxgyHjMncV96VAbBWUD5tpymEuW+bBht6ZI2HQRXKB33uh3p22GL02CG9tuDC
Rk+B0YhrwiKA8pn0GctZtQfRWwkFxlHEqbiycAZl889BgtJT5X/U6FERCq5pdaPs
zBtMtcgPaC08v8/wYE29jOO/fch9rS9Wjhl/Ag+njvKRcsha7UaxAXzYYlSEFOte
+VHGVJzrJtNwJHk9GI5p78S1aoZfHnCckGffc2hamTsdwnNuUT/VL6kv9w80bBOc
aWhsqfEYXxnnoIf8jTcz5K3sK8aBqkqqbfcLNj5lNoSXCzdgTwuKqxuqgn6VpRyt
0ajuQmDWqp45oUnrgBNB0jHRjQuSG/lIv68e70Lk5Q0EAI41nACIosmHBp4Bb0Sl
Q9CQuhBDq8J8b0n2kw3OVC7fG0K7n8MvWSDpAfhjRF+S6uaDgN/BAwsJP3tt9trx
wAh6zoMqLxVa9jv/TIUJMdpEiotG+iflty8/G0tfoQXPyZEJXLlVAkTus7E3wozj
EgoUEi3BwY3dLPtAYNjwQGN+7dVHF6k6vbZz2uZE7FFVQbONibV35O0ZA53xMOBE
hSU9Z1e7J5o7mhVt9+lADkTL4SCEls3wg03rUeW+h8O1AZbA2g9JXCthrpV5csRb
R/1I4NoyPGBCb4ijw9wFRVjxkpbW8Ure7cRbwOtZ2uEQEiun/CP5/dOhJNhhDAzc
B5UIXSl8OOEB7IreHYYOtiWfviY4wH7PRvcNF2J2pcGNbwH/A932hilCXEkjMu96
TN1KjneqvbRGsvwdybyf8UcWfKAFVSyaMiVCwV+zkTDHCZzboVOsIOFGRoZYAOSF
Pd3Mk62RMrHap7xJDMiCR7JwPPCC9U2pqkrkyAF2XQbkWDTfxkfI0aYlbTO+Iqu8
wD/gRy6mwV1MGoQyAeXYaE5ICIG8wZfqsEfkrkAPQHxjkPlEuGRGsdfi0O5Skjuk
3g0jhaBK+9VJMbhSyMd70CIFimH/XmpLH+tQwcTMDvWLdFHZn19bpFvWP2KAmV62
nmQpC4PAeMZUrpNkE+0O0lfoWGcsLEHyov2V3dKioPfBchUCTYC8Nfi0QugKPkwr
jAX6D+NXQ+cSZ92QjEFctQiE/YbG8PBizTT9uH2XZQ6vnEASsW/t2ECbesGDZ1s5
waH3yAxvLHmkX/sGeeqQZFs1nVuRtm0N+ZEt2w1m2hjmMcIjN5GOZKyaT2UmbB/2
7wAlyaG+j1ebomDhRm3aDqEXuyf1ZkB54ovmjuaRAdvb/tmcFdooxXYacsFHDkLA
6r5+k8dajI5Kj+ohoTmgR9psbSD9umd/pfoFgc+PTqdd+lHA7WgDryJZUGAnBNJH
x16SXhDQbve0pwCMbeeuWKCI6SnHrYwz2tdqJAzH7rRvTyXe7vTxAijsphvb9h41
jyCS/YdKW9sb2JijE9AT+6bAq0273IQJEIaclTtJUjTx08ynmfqxQiiVRNvjJz3L
xhcAryKVJae466SBR/o19R6R/8RMCOmU092unioJX5BLCfT9A2vz+qwNo+9fGw68
8RU+jNDUIk/TS3UVRT/rCh8SvUFjlM1eaHfGwVemWeNmtaNEI0xGsd7CTwge7CtN
cdvTKWZ+W7DLSeyACEGX/aPHPertEiDWWildAVMo0zyFvf4YolMvI6exOveEv/mi
Y7Dj1+4HsEvfYFIXeEkRA5/aQ4Mh0RA0gGVhsMEo/65X2JTIsj0PVQuNfw19CCLm
baZW3LEc5VsXUJHREEQJYqOBEzbYqJ7w1amfZ3nrYlCZmzEv76TzYL2JJ1veQ3x0
ds1EyVLWX0MWNyUTOoMY2O4jNp4ZoWEC3/6tyb35ZRPunE1deFXzupSWDLV/USvc
AKdAxUw1F3NAXqwoc1x9QNZuz8Rl73QCgCmlsSwVS0Cu8JOgnwJQx2rIQB0mjn6g
1Rtw+bDQID/Fadtc/7pAy9IYUMzK7KFYhjyTPS2Zfem0inyVujO9K42ti5AVlPdl
/8OTmpxUTq+wh2n1K+x+PDrBn+Tlrxh2l1CXyU8VoQOQ0O1je2JUMpkUYFQRP07i
c34NOcy7g1fNvcfE+sCcWy+Kfv5jMFRgHyqlafK/TDSEjKzz9j229OgyaCjXAqX0
k3kM16n5VmDROBVYriqRegHzx6jM+MLQEJOadzTMwG31DZC9jW/Px1mBYCta38s9
gXswLPtnHbe5vvZHMKFXdboyGeBjB2MPHcrA2fG6TpNWWYzAZHhL1NvRAZdiAu0S
/rHPfaFZyFabv6CMBj7QoT3EDir7XG75MIMvLuD3itMNgnfa/x8CsDZNp4O0QLeR
9ODt79rwi5Xm4TagQrj43pvdffC6HGEMKN4g6B1QXyPmoHJe1LBd10hsYjXh2pXX
CW92K1KuJVt7AaD0WKl4zdMxQYxOlgRKJ6Yag5uizdVEF/VgI1bYzggWZ6lhzntP
Dr/zQHBsMtzkpUfP9ktuxuBzkPDRGho1Pb+e3oMVuE4QiI9KRpqhu30h03w/pqWE
ocWFdoZjIqiP2x8lRwFk7lChzvoqHuSDrYtrTqqMUlIoaaitzRGtZ7ekv1AS9kx/
SxPDfn4z0jxrM5J5PPL9bAyXKAym5FlvLwwpsEttZjkLUYktnUd4j18UYnBqmUyU
85uoxszhWKlO6V7W3jsrdSIB0vEOlWdc29jRaXP7fq0fdGF135Jzoqna0v3xfsN9
h0li2IvAu7xUUk58CGbmcAfaiWBMpslPziTQq/yxZhubhnjn+EXHHdD3Tpgrgo54
YWjomccRVLcR5LnYsWr0BN0zZJyCU1CvfUDdcs6rUGeWECS54Wvg2j44fUlqQUip
G4isdei4yL/BUCdGPkRCG7SmwLCYJ0B5nJZ7Q90uW+Gpw+ue3dJGZMs8rjtYPugh
25588C7zTMGgDEyZO2DB45nQldSyPGyfhvhCnoPInAF14tDId5QwiDDb7MUXOt6u
fbEz5SYdRq/gBd6UpAPlBADKpf38bOCl+B/37r3dRmI+87UeBgdviYvIHOF/WFN+
Hs5J3dyl2h4OrdOceiJ8ZIV5bjV+IniZUDQPoHzlsY9qLDzNTHc0f4Y6N0JFLwxM
fy0aK8ASoK6EIkJwz6+Os/ox8ksoksk1ZgZ5lArc0ozrBf9bgPWWhTw21sJGHqNx
DKl+Kwo/i0htlEjnEIfKGHvfF+b20qvewZHTZN7vtDywXfgd4rMivTEQX4plD+bQ
Dts1sh0Yg++b/Psg+XWjwzxbEI7Y0YbctwD70pFaWUVDmnnurWeY9iCdy7R4BvVb
dOvSy9KxDTqM9HiFdXkedEmW6IVWx+QiOesnQcI0Cw15Xqr6FW0gwGqv9MA4W0Zr
ABqVqQvRWjHeozwAYrd/1m8DfTbsep7RdTFu2RmaHkYuzkjWW7QG6DaQOhZXP1JR
zIZ31hQPQEewh4PGOp8DgrJKo1Ug1/JDxktcAHma7/nDbCdNlZ+Ixl7GfxeHZmJu
Q9Bp3W2z90jAbfFgQPXK8FoTswYRAvIU7/IEn0nsbtLEY3WDdXK+aDbTTxthQE/M
7eQoydfoajIUN9PUUy7L6RxMOYpbqY/8TMOMRItDKLcAtNRjMKZbJp9aVmrzlpG1
rlO+JUDdsTrVHkvAFkigNPpjzZDQ/F8TmBnGOrZdPlpxli+dN0aW0Yb6JfdoiL+q
jDbzREKBTXcG3TpAW04EjosH3JIdw4AJO3DUarE76hyrN9ctPCVEPKGf3LJw89vA
M4YadIwb6Shb0KZZmzw2rnOTTHSday2CEl7ow/y7FnC/AQG9W5KPVJYM37q0QQ1L
BEFryVIEZd8O71sK0LjAH7inEOkb3Dd91N87FqAl89pQ+crjlq4ERKN+jxOgtqKa
lP23HBkNoyIM6qSjBKd4ktq3cMIB+5hviAkslRQJEzRGvOl42gSlwqBCcjPaR3km
Rp93pdtNr6RjGHC043xE2sHbhI1i3x8eVSQpnnF2zyTNmCXijCfICeLYsNxWGj0b
zTAXjt+cOdhYmM17laZVqLXz2X38a/NOSGfc4x6SEwI8yBuvQ4KjdoedLt0PAoGy
rXMzjWpO+dow7QW+eQJKNl1OTR2R6hH3LouU8xjrkQ8yJ7KH0tkhw3LxeD314o9o
npc4qcxXCNwYJh7A2s1lRYEC8sJVrmT2K3D2zrBmMlAbki9lPI1+BXO0rcKqjw/4
2hGqrPU6YyuOMgaZTmxuOqX1r0Fo6Ert//tMo7gu2kJOc5Yjvf7y+Coa2sqyMDy1
QQ1EjF/1hI4DMRz9vOzNIjftwHnyj61wgpP8+Qoj7lHBYvmcbeUO8kJ0s59y/gnJ
W/P/Ct9phGeKKm2ScCXQIjwOu+NxEhWaJLkfM7NLUXnkMfm/CnJTG+edwQkhZ0g6
K8tg2TmIe1CB5BOxKvzvwK3xECQPiL1eY6f91YwaJFzhV1QSjVlI1V0F6NXiuUi7
tHUchHoYco61Z6rKEqJG5YaNWLPtYmfaCoXjaamVO58CPl2BovnZtIFoV+VabvG+
Ofr5OmJB36wvNEdksQpVCSKIo8+Y2NU1CraAbLMLjLY0Pfsy7zZdPUwK83JWUrjv
3diEFQ42XhuunfVFPuRUGjFnVCciTzDH6qrnZ5bAoJQuleyzxkK8rbL64HNfqDOM
699pIEL5V8ZjfT5FsLYsZueS5xXCbBy73IQUAcwZJrExdQp0xmjhY7vdw9VBRjpQ
us7cZ6y4Qg+w8IOTHSOWHiASzxSbQZd2r8ynsrZrLhswgx/ij9SyZrmqol/kcXkX
sUK44fAuK9w2K/M50ecMF4gSvhELZVWBdL4hpWHIJq+AVsKnywJiw1RqpQ44xCzC
VtHezmQAr6id5PICpDq7vzjriCDpyNktqVV2LWmz0Iy1tTAL9VlL/XLC68Mlm0tV
sN6Ngv16iBjFJaRVLjkQ/TW/u7F7ADNOWtyVb1ytdFEnF++hU0AuNtkkIBm1TFkv
+wcV+cn2ztSZZUPmljHF7F9+3r6Bmg6xY6qvom6TWPiktW5ZQufjJvSozeLepyEK
gRqtrtx3iNq4uTojpjZ5VsKoFcWWkB/s1N2E/jNEM3hr9zPkEcVeBLtAWY5ufbQD
WEQ4C8Mn/0EqQtrt5wKnHhgGpr0ZLVl0uEX7PbJfPWHszQzIMRCtbUHmUoe/oXyL
RRcgbZFGl8tcU202H0tUwOCxYKxhRYLSVxqqEWKQjZxBXQNxAVQv2XuamB/lP9Wl
q0iiLA5yepMoU1tD7/xv4SPpONvx477EWjROzAqS4ldId4vPoFA1IvaborXiwQcY
8y2usnp/JALbX4vKz5kKB4mbXUdIXOMaF11doe1ugVae1rx89hjV2d74eD/CaH2w
LFluojZ1H25YfXTWZwsyJbowar9mWxtftGqnKcNYYtZFebIPdYrLW7pqLSmeVJB7
C/FKONyJjwdUH3FCZXXJOhOhuzzezTWvKhXPZGBseoS8j2PKrk4gIZvmqXX2VvUE
XozZSAl3qLj4oQAZhg2twJDEMGx/mfxqZUB0aVHtj0w5cwnRopA+04MCBKlBAKfG
p+0dj9848dlsavA+n/5iynzXh63bbY43Zb7HlU1olbcO1R1lHpKVcW0wRp/gWyI2
yJkyqNLB0+yR0LdkSpREovdn+4gSWoxBkwZ3OyzXzQsHS+E3fPo56l/+5R88SV7c
sl5uwP/YnXBI3DV2SGQX8IKTo5rv6mDXdxXhkfIkemDeaws9D3M/oPGuvw9V5xqM
VLCPU6VJj7jO+Wa8NWy5QkCwtpFxx6yrd+3RiNhMCbp9ccuyhM6HkR0wrnB4Y26V
Yr3RRQnDvkCzguZteKyBMbbMRaL7Fd7veYlDaUsib7wcEsj/yf8Tk1dd8SOheaKa
Lr8esiaS3cOoeNny8X0pU1uwHXZfF7+/ktrnT6x3UmMqvKktdy3imWx3oLKc/3oa
FFX1Cp+zLWGPBuob9ix8SE88d1w6E6YSN9yZdhKElJxqlr5XEFrBenHQUzVQ6W8v
K37KzXLxalWHK3kKy2l1CpFeS0dovp8N6DTin1K4Nu/WnEPj2UCwsKI4oTEckXVd
6K12+Tq8spTEiS33l//XFwqxLd6qsuT9vZ5v1iLXWG64GpWbaiff1f5G8kpk/3Hu
WdHyufKbP39AXzJ0mSe9i/VQ++Ce25fHYGuMQY6tJE1KNsFSsjSkg278NSF/+uMF
QEqP8MrPnQHiClELwGK7EDsOEJWFQaowS/ahXQMxq65CTtwl2PLzTMyv0D0MR5iE
knlKNSThn30Gmgw6OvLfVT9qF0OisfkbZr2GQWxZyAGVIaLZBfLCWYEPnsNn0jwi
+zBN7lHbVdpVsJ7T2ZO0T+JsQU510iTuxkqsYCsXR1DeX1751wjm/CGfngxD6ycW
zoYJrAMlXbGFwqQcI3JagHqm0mnky15gEyX3mO6TkdciqxP9qCe7rdtwr4n5/kcj
hT0/7k8mfIefHsbzUMUVwH/Y1pUxBQlVosHhhhNsDAZXVCj03RtvoEctYHh50zjd
6Wa2H+bVUjBRp8QWJhzGN/HtUM/aACPC+0hdVETCsgD/R5hgN8TejUk6TVzR+J0c
QFXkPgCx2jhFjZWaL1yJq6MkrCUCeNcvBY4hRygrvfLl+67UVgs3DVnkdyXk/DBB
veKUPUt52XsFfILZ6e3Ca2G9oTrtJtzuTBjsVNyt4dAPvC2y2SFUyFP3xeFs3WlI
yoZQrAYwh5DoSZAV8Hk+yTuwxI7JE5aMFMZmQcnwH1+06p0IKQIAKqsXUTN3tEQy
to9aYJ9FwAw/tQb0p2njZDSyZpWaOKqaCsiV2eVaL9MJLf4v/JnzH5pFI2wOmAjH
1ChCNZSNi6Y9P/63/nbNHGlazwLKci9nJSifYRq8u03gWA619FhXYYqBVeWm1mcF
yqkyy/WDxkR0Q7Jv+6Vjedw421xxK0Zlsta6OODZR+G6/OCZkVAk5qA0pgVWqFTr
zrCa+6bj07zO00mHCuqNiJxRBq1J9gS3NgBuIakc3aq4GTmfwzw03wOp0cLZKfZK
q41px3La8GUalF3Zq0g5SXBr7+p+O38QyJbgSbpZSAqt+1OXpidTY6EAvueXr9ye
dUXJl3DQQ1e/tLG+U3AjK5c9qcLlywGSwvQktedbgbqOcfsQgIoJbmcfPWK2nZEN
GavAR6ZenX7rmR3jlAsiu56u5gvrl0h6ZMhtEOY5/iNko2mbCbAK16s0/xL+8HiT
5ymcSuPj6KwzBVT99u2BT08uKjzZBIEoF6Kr8sDPQYZ2KGICVWT5XmPDnBuFIW7h
YQ7J6KauAeaObJmKNO21K4uMy1JdgGhu8KPasFMIVlEyDw+oSCWvTNAaqH590xMa
KunNk+8yY1Uh4gCof5LPEDsSKni2kLaYrjVB3376LkQc9le1RHeRBb2HDdcHYJNM
wg/thndS2YgNhclMmMQ0Y5ee3Y78UBtNlbt/5ZntUO3zaUj4cbMcfgT7tLd6niGQ
43eIezPbY4JsG142b4sV3DUtiRQsfqUi6I2ZY1VtbRNozSSWmDQI0wYEGt5Qc6uI
cFzcEu+xChwiH9jtA9pi2pX164oYkuOK+mGekp/SIOWphpnHV1Neq3Mt+wZOB+Me
ZWUKttRPpYoTKZlDRXhsucBOW5gXPA3PqR4W1siz1vhE+LWiJiNGtPPqIQn8UK9u
63pbcnDZYSzjFwLrt4UK7x96BMVDiavFGrTCEJVyj8SOcmvH8pZnBH7qDJ5ZRqto
eTc2Cs08fZINw2T1WWHbMWSHDuNYk7J26AKmjemh0eaEZtdZMCnrOd0pC9wevoEw
zQrZeHeRm0L/yjRqCdxF7hpygscbIRuXLT1j0lvS/W2fldqYzbp/Dg3X/Z/8w6QK
sl7SCfjBOTrCIfwsgrbxkfXdmC002JDso1/MfmXaAWtNXOyu3uahrZQmmUAQdx9u
zmIISD1tgBVsuMg+805vx7L1mdYAirLZryMZnyJBeGimCwNCERlnvWaxwqC2psrT
/jD5xU143huw3xUESMhYz+bjtSJB6tSKWlsNqRbdzbN61HVuDK9otk6VfXiUo05z
skJ5AHLsbMpqXUEe0OUiVFfRB/QZJPtTG6+QZ+LNjTpx77wE89kxbhmXCjgZhUQ2
vDXttReJwOUXHoO/1Zct/IF4E5+rOFIVCxRYwuuEBFTz6g6jrD0CUMTtJFadUQpT
On5rPMmaZLSZS0oxx7K7DwnXevZtxK+lDY6+ffYxOedojgBqs817SwGjtd78tQYx
cZoNooZmWQp58JViPRKx+mC3KkvTWQfmsslmCcbCpWa9qcw8u20654a/mGMqAfbO
pl4r8DsqMJeudr/I1R+FUSnddHo2t8T0r2kZzoZy/vjA0D/X2fc3tzk5DsL3v9yU
UmPMpqnrXNeoeZomz1WgCHhmlGYs+A5OcF9/SyE0+zF2reDrzjCKgumTk6E7JpXA
YW+ThEhyJ0ieDTB1b9k7jFaPEZUwyFTVnuqrc4E6TIGjxwP/Vb48/OC1E4uQVbPp
LTG7n199832MrZ1cRB5niHeHfgLEJmuQej6zI9P9/gFpc2Yukvv8vHyuzKbUfkyW
7eSS+34Jo+hQDCLG+C/hNsyWnZpu3YX6n3ZCo/8heyK1MuL4axUsA8cpVnX9puS8
pliQRrSpf/mEJOjyQfE3bKm+tWcDPB3ZAFpYowp1lb3sgII3TwVVgGVimwnJ+OW7
loD5vxrfw2zUIGCy3Z1OGjBX7e33Gd/oEVrl/8xCvyLfY9y+Tbv4S1nPUlst3vYs
rPsxx2AtY7wzqwomsy60U5RoAnnwvlPvIBseOxe1Th9NqCYwH97c4td1VER3LAUW
nNtmera6JX8pBl0CIfFMJ3LEcNo8CP+rkKtgvB81zTYve+wP76iTQ9iupbsqzaAU
aXjaYTsE38VVb5wYd6QuURT817XoYW/ViJCbI/kSvUv4APeJrXkT45twi3o/XP1O
+a+k4ujfJ4NXADKI1Tg8cUqLifvsW/Ik03x1iYXoBPLTiuBSo5+LCBX35PRee9cy
1+xxRNKY2frEFmCb2TGq+Rk4rkXEZVaU3ba3QST91UZ3QRQiWC0Gb9JC4sK5QR+Q
+eLQDpR4DCSZ3+4EwbFi/w1Av/xZWTJXTd4FeQlcKD+9VuCvA5fmKCoHUzEvHn4X
SF2VPwduM292Fca7Rd7rbbmzuyQUZ+XwT5GL8xED5K+ulakbU2wHOQXhn1kNbiAO
Z88X8VA3I82XhmFIW/oZF1hg1DdfpS5ufbKYNK3R876GWNZibaAqJCraijt1cAS5
sihlT7u4OXk2e3HCU/oNunoGir59OeqHhRvxcrSQbmFLXsgzJFQ0ZYq92mUcVDLe
AXhF7wiP2FCUIh5RsJ+dI+wAKkV7cmI52BBJm4WYyZQbBS+12vqPtd0kM4BQIYvK
Tykq7tyFAFNTSIMsBjoMisRqgeJojp1YZf6AUyuR+PC4hLzLP8TKnRHz0L1oPXQV
ElRu9ij9hP76i8q76KshcKRS3x3hRlKCzvRBVogqSPVNE5Eq3yFeybGb+3c1a/Ek
plL7c054s+NjrpKhRB4Ney3PI/PT9jbQs6j+cnmoLUmGRCHEEtfesOb82QK33NQZ
Q5B0cyU13qQmDO/Flmgi0DRXhw9+hROEnzC3zmGr3UFFvskhNltFCGSyLXhe3C9C
ZjstM5X6YU7dLVVjoaF2Bp+2BKVFI943ku3NYfKtsrxdKbyJ5W11m0bM2Mi0i3ms
TqzvbtzyDai+NEXQGlAC7mu6NnVZ85IP81GGYZd8p4l96JN9OJExOupQlXPuL1Bl
HiT5JzeudBf3iZy7hBO41aTLVXfr1MgsXkPpEKdeVqlEnYM33FJd3HRXVbC6W8Ly
wrGxWRXsM7fRz6/K/NpckUctW+i4TQkDmxAGjH+J+EX8B9UdDMoRcpyF3iTmhDC6
fW0c9KtUf0fmrD137bFIhGhNGTjrQDBGWdKulxeaeetMdFvLoiun8ogOBOviECs6
SeyoDQ4/n1PFPy55P1zCJDQ3qELMkewSYmc9pGT5AlFd3EThSY4EXafNPPdIASb6
x4G2PC/il5M1mzCscfe9SwSQu1cmTtO0utYf3rJ7xsJyA7nTnJqh1wqrJgXU3BRX
tM1/XjXLf8bfelrFH259RYnza2wVRAopPU2Fi/IzdXxuxfKIsV2Fnr0nZTjy40LU
PIvjcYfR9HAXqKIv/WDxdag93i8ZWW1tpOVkYqqDgjRmpy+je+msJPijAQuRRhPx
GzA1fVyu2YVe41rhFKgfIdKMwKGxRcxU0r+x8aOAYVhTL9WXWcLT5hCx3iRers5X
g25s5EjZaBDQ+S0acZRXdO8lRROp4tMFmI+UlXbrKfWSV4UJM6I+tB5zLB1VR4eV
N/oeBeiRIrEi0XNZ4SPtXWtzPmIqmRWOXfyB+Woij63HX5JS7CxQdukZZindGJJ8
D6Qy9flHhUV23AR6ut679b5ZaIfXu6wKlEK3fgIik7DYQryffbR/74tC/9bZi3RO
puU0pjr5ZrZ+QbywJi1cc6f7F67E4F1xbckbrCdRWfcGBcIxBkPKTVci9X5EjfAL
j9Aw7RHykdVJksyINHeVVblaG9Q8mz4qZ4xrtvQzta8bWSbnZdv7slX3BC66Ky/a
10e/4FF6BSA7p9uQNnPKw30fGyiw9ahYf1B6PQLbo0jmhpv2MbYE136nwmUlAYek
9aNy1qDdNkD9Mhq4EmtDTMwDF3IyTF3uRG2wKET7WBYUNr1UEeu8jYkomq/M8LZm
hwnr/ueJ3wPNWtbIC9JE/WtIx/lEt6fKHFze1LUcCtQ0jnU88I3QpsVvFBNi1qD+
UUwxVn2ua44Bq4G2dwOG5kYSS9oiOlKU/enVIlqm6uPdaWd6gFzNxYAN8cVLXGt+
G7QRDHbU+wZj9I7rUHm4k1BCquygC+yMapwfaz04jTUaW626hawSOVPb1s0GDRSn
MvXu0WjUqHxu6HTdg1lC8mAkv8oKOidHxzK5+bqbxgc2DZ+qsnjGZrXsDPdouB0y
cMXxBXdGazxuIVUXOZ1oKvPfe5AU+s96WlSFPF+1UyLbenWR5wq/qwqwgmNWiJTM
QzmEfaZwGoY93wPDb2A7A4H9agZ+Qzw6U8aMCBIB2vl4A5RkQp06YEt1rnMXa0MB
qDrZFbkKosmWZXvp0B8nxzzBHxjJBDDsbK/xfMWiyjHz+YkamRtZCC4sOFBOUZRc
RwvhDQ5gZWsLwLHBZCw9gp/+IcbkgH8wt3jVVe8qXQw0lKfYkofSz3aCbnKtoGyR
dmv8BmXPII8UwPmquBs+bqCaXnl8ElRxxSFjxWuPvJjeKNHmAv/LKP+smXczwt+m
Su0SzYnO+RAIW9sIMOgjsDSwWfYt6hZ7xPWgo/nmna4w4SlvYu0W0cuLsLSd4bnU
839S1SXYUIwQ2mRcjhmhqORIi6dFwvi7XWfbwxwY/FLGQi3aoHApSieIMl9YGcdt
deTbEd9zqyQo6BHbKKu5DfX+t/jLl7Tr22sPqMzO4HewyFjgWGvPBThQA98RITL/
mt0q7y9t9CS6Z/ZoKFMLE/n4a/ehfcgUTN+ODopbL4XbVP0q8fSeKWnfc1fhnt84
sitelj5hSq6l4q+pkBo1Ah0rkBAGzIm27yHO8oKYdrzExL8sFcXMJoQkgwT3hAvy
6FwjA5lOqeqO2JzFe4NsHQ0GD9fQLSm9pKutgpLLFGvhN1Gq6fhiZH66XqB+eLxZ
rPRCLQ57mWYX/cKT8AHhE6X8v5g7N9Q9+RwiGtnNrO4WC/RYnjXM5jljyfZWwrNT
FBnmS+MrxAexn9TF7PWCb3s9uIpwIAQPNkvSb9q70jl3n6S5zbBu7vWzoY3MSwp6
WtEowOz9Ebr7CRd+cPjSmre6AvQfFU5bDMbQ/1Y3OLlUtR2xzyRnRuMZeRVAt4hk
xvKntzTAY1YDZy//75p4I623KU+4gldMrLXO84meSULfCT0sk2LcyvxOyAnKEQzS
FL3L0QNr53B1HBrF+9Kp72yCvijRCt2Q0mipRazTCM9sE/isA2bgSXKaRbMlrBLL
tpvLUNa+klPz6vViddccgXAjD7wTvYdBcXnM0PXiX9nbRKDdM5ZZPKsl2lcRJOSg
O/5HRQoGAThjkv44ISQQ4iHFs+DC7k1M5RtS5niLkbnEMr90mg6idXDdb/d16tJw
U2/+eWwfAZc8OTgjB1ra0k3hRvN8VLhaLnDTMMdoq6Qxo16WjFyolGYzhtAotoWU
Ng+2ANyyDwc1f+REYLhsbgUC3CBE+pGzReIJTCqtjiGmhUHMt7K2r+Q0WzMD0wMH
5GUDaT8nL/LhEvtsNQ61zcHvPaNV17BxlSz30awdU6hXOXwO3cTegNml6mcX4yW0
88+z9zqFyqVp8kCSBD+ClOoxfqzp8wY3S6fRuPJBVB8dSVyychhJ5f4aXYDjfGxn
e3ghVHRyIor2hdrr0nwXIgLFcA4XxhinuI8iwnEM2eNX/GQ/enKo0jK/hRWZ1A3L
zuhp7mP7oVZceoZdouPpTfzren0QJlpX0wvIcj+h54IhCA0JQu9c7x5PoxQpm6x3
lwpxN9JU1xR0FCkxdwZdYvtj3BW8hynsZjJu+8VZSna7VjqFR/wBYEEJYLTLpbB7
zEyC94xMOctg+jFssB5NzopTCUyg4lBE6bKGRYMF3x69wWJJCZZ1ahmsIVYZZbmM
Om9vEHV0PE+jb0uNgmMH2YkBxU7yXzLljKj3KtVzjQkMnd/LItNAXXAznsLKNsXg
fmuwXtzYL1dOAJiOMzmTZBUWj4KuIz+GOTJ32BQyIEc+8OK26UNUwhQ0aOANdumC
yQU2MhK7dX7iTXKvqKcM+mahdPPsVwZP7OrdV/CaSP5Xgoqvm2f0dpo2X66pNkon
ybCRpb9bFCkbj1zqoo4DD96NHHfxTzGJuvbbChy5qIIeFjIvKRvMQBeG6F1P0LFa
pyz96/ddZEuBD34GTBJSj07yvQO9XJUiMBDdiYtxIOCgEpAU7IueIXFC497Xyghx
BRWOnZ5YS5+MOyV4Vib2z34v++sLF3njY6c/2n66bLbT3hRwVPe7Z2wE5T/gOwXM
sbsFSelHtb7GoDoRbxoGR/2b+5S3Imlw5Yumtf+UGVKaIhVTMzEW1voZX6zUmb3B
ZSpmZ9wgTiI/jx9sH9weHwbeaFKdEwuuFjJZLZrGH7BPjCoZH7Ed7ITuy8k+Lczg
SAfaZC3v6klr5IwUdOcbl/iHhPRlYm9PAjNAlBSz9T3Kc3wzFGEZwYeKfO5avt4c
eaQXbN9iqwfexw6q+S3l58oQRqjEHRdRkoWaWWLFdLtiPCbziDiOr1znOGMeUgLD
kSXTkcXn65J7lHKwyhoQnClNM2PBPpmDBN7C/9I+DXlQngssyfhW60X5FB2xcFz5
VtUY4wXHZsELSzEsFeGjlHfLHSrvoFImSQxNKF/lMa9XxIKF4bEDtAXDyDSOJ63H
Fu6kIKSzeiO0OnYMPjOARuF4XIXT1v3QzdLw7iKNKA9YMQ1D8p7wWJhoz0wAKYW9
BTvU6K+8I2HyIECTe0+lMlZ3NCnwxmFHzNhyMZ6t+J51bhcuge2dW7Jz17zDEM30
5Npyo0/Q34iGLdVc6YEL94PJ+95sh6pG7Iae9+5kuqIQmAR7GWEXi65XS4te2YWp
wZgEK19xHrTehS5U480yWzV2o+ZiOLV4zaZEumYRLbVdKaJv54hiaHU7Zjh/ffK0
2XaPgLV1EJS0AGBzX6upyBxHfVNWKZ1IdS2UsjcO7u/LkVeN0lF/jdOIfH17an5f
oe2F8vetYaldonTZVr1UNKfqZ+XMktydIDISkIzKfV3ytzHQhSJJkRch6qmeLNuN
lGuxmZCXYJaXYtjO0DCzLhbBP9hYeI27bWSwGy43Ehi1DIvD37TQZhC7MJD6NP52
ckTFgtX9N4bIWrXah9fnteVoFh3qnWLpA8gNnoo6lY7sRJ72kAnAbQnJLomUoy/C
9rmfBg7kjtlsst9bvLxHjopCGttnl+cWQarZTlwImiqak4GUP/H8A8u5VOYGjnXi
j3H/d9FtkG0J7llaN46LFyAOcqyL+So9vhfqRpQg2vEEVONPpUe35537kOVcELLq
EsRmx4+6XW84norVtbGaPpm4vI9OxsL6xj3KaZPWicJIhDWxavoKgCsh9ZpxyJ6T
SdYWgBN+Gt4G6L+VI44uncXstZsJbQfPJ3Kb0rsshuxvYNtp6NjUk/ricSJK9wQ4
+VbzgCFA9dkAQZDtcGwWabSoehTBkGW82xfoQz1XMfEbhAvwQg0VHfw8Z/AjOEg4
Lu0+IAnbHAkPdEv5pGY+UnNh1HyyHpPIhUId19Zwysbv12qOE65bYnZtVb3gmhT8
9XexcokpWNiQmQ9eYSV06peKsVt2OJZvhHQu8RKLOMYAp6Rf/OsdDcouRcVoI8TK
U7vuuPgUPvHs/lh/NosPvnLSpGHanf5w1ZEIpYZ7ux9rH0A+ew5/v2A83IVMFbQx
SeRm5aYPExkHONhU3pDex2dXWh6kJMGkI1meS2RAlXC9wMrdzHjlwBiVHBsqwlNj
/3e0zUJ3+yTfDJ+2wq4SbFjEuheuJPs4D0Abxab03X7IKj54GXVOyjT0CE62bevM
aTV/wA8V/+mbqKWsSMphiapb2+WKqhQV7nAWKri4LhYS1fKlLvimjRo0McUOkWBV
i1uOCv4l5EYAaKBdjPiGNKo3bB9ShfBNJmzoXAerzHnLnfzJyy/klyxp1GNBdbfU
BZXmxEqoNLJiX8V+6C/zkT59nW6HarzOparyMRoT9TU38rIGWpQ5A5iwLZ2h0lVM
DBw/FgrSHCGi575nP614CzkipSEOGS6EuJuRtS2dsX5wkSGnDIJ2BY1mQoi0GcZH
rIh6EVFB04+ZyW9uJcfh9AY4bDrEsgrg8w8/D0Zwq5DzXxtql0o1wx+kX0BujKUo
4gde0d+1D0YiGT7aULqpQOkvfZ4SOsamKe5RcLfDMe7eB92hKVIQ3IImGuASTgna
F2BjopH7tD3FvP5+GWkH8antz0valxXCNYgRe8I4Hn2cWFcXUO6jXa9gVf5P5uMN
nb89iuZpMAG9ujRz5CVSQwBhHOeZeNyOSohtA8F/iRm6/ZzbhrlPMtEu8Sabgzr8
ENZPkysVcrWQxa2r+jBIByfbQ4QB66DITfdHxDurX02RsqAOh8ppS1iSdAo6jU3M
5UceserZfW5Eu16p0FQl9kPsPpTI9m2F07j77CGZsJfPDaje/kWnszrIhSvFI/uJ
WDg1IngXbUBJC4068plg0P5eG96zIC9Lb35Vbqquc5qRzASSBIkFasDd63lZDa42
g4cMGtLEpH5Y21jSdHnIOHGhHTqYNoytEXO/e3BuQ9noUMdqqo0ErIKNNMK7Ou4o
UoBDgWUpaAuffPQNAzpCGSpvFs6YFoaI19DAmTstfH6fEIx0H3T5AylMcSD5XuLU
vbNwT0CQc7eO9yiKKpKi/JveasJGW6PgiBl6SSoaC94gPHqhVvbfrVQB/7AD5vM1
XSCQ+A4RxLHkONe8kCcLaP6VbvaZDOofVP5FtoIRtACW/0SyyDgrJ++teRbSAaBl
Oo3ZKnD/nn29M2G0ttWrpeOHNXjtUK9eiUcgZ6JHPDvjXGrtBpUyfJpVb/kmXhFV
6XEA7hIXTMYnvXzkd8RjLq76r6vOvZ4+YPlWYTv95Y7/QXUaqdG84E2ala55lt8g
rqjJLUv1mq2NrrBE2aP8z2lhf0sznlWGc3bcDEr/178JSD44Y4qYH184ooJlEulV
FKzSQeA7j4fJXpWU8eFZFJp1SIIbV4VPE+g6E1PkiJDI+PrP0qe7cBtEYnAvF1GC
n9nsxSxBPpvxhxMv5B3BaDkG2h760KUtya5RBg4OmDZ8SdVPU+224D9V8gOgrd38
CWzZlevXsa5EElXDi5fcB4dwYG9Q0t4iCSp/MqU97vWQr2J3IydwDqvl2T4GImR7
lRk7zYzaPi9FurL0AXrNyHCK1Iqfe3TnJ1A1pXEVla5M+zgHm7JTMTcI1iySfK4O
WUD1CmhlkKenWAQ2ttheGkFZszWmMDs8yPDfIvYd+3D3pFfZrtOVD38cif+ucYOS
9GhWYKfYAatoeKmppI4g7ybD7lLPO3gCNT3Q82g76tlz5bsT43v/zLprPpfAMmDA
6/JUlpndRVRW8N7LZm0Uf1MPAbEnSr9SbOD6YnPLUYxJ2vJ74UOVrNaPOK8MF/2n
NU1kuw9L5ftyreZtjJ7ftMvafjif7B5Cpog001FmR6YpSO1tJzQXP8StgUaTRi/g
sZcIhh0W+eG/wO7H2ohwCtdkueQ9Czq4//MUxjcr6uYYyd2EjovbA6o/bONHXFgb
MUHObIblTKYVPY3lyZXAGHwgVS6vba6D/2iuROeqK4iAlWS+E+q8dq81yRw8P07P
+OOBuXw2SVFtnVMeA5VZVltVGxhjzjxm/0HCWzA0WW4as0O07eKdKSLh2oWx1jNe
W/31Z1UI4YHI6FUmhg6d2NQgd/O/NLVISaxK2ikrWORzDb/aBwhnQzWdZZo5t0Dk
Fp5UivTeLEnC39Dii/UUIFH5jLGl0pK6IcKfDFX/AsX0OBjw5lfBjpGPCiyBdetk
67DPnVt69lJc7VfYUjoVKguhVSoX5T6gbLtRMq8jKv6LJvC+QNS5SwNmlLRrXaNL
QHrSoAQFiXWa/qLadXQr/f+JGDazuDAM12g2LtPFW4t+OB4q9wBgJSmse9kV/0vN
MIaBJ+4POsOiiLtCU7X2ljjIanOyJhv0h3WGS19HI0O7askndka7K4a3iiBW6e9t
herkAmVtmJ0j6ZYE+sWGXWn3dZ27Cjxq1PrCE2HvefTYlRr6eAnhrDi7AJH66WFW
AI2eTX8uVdviT5fIj2uXlNE/rTKDyayrAlNhjEYx60c2AhrlgqoblsTnQMrYrQtw
CNKZdAtSGP5mylArOFtG3C2l3GeHLThZlcI/8ajHnep7GUB0uzLIdx1KHxl59V3w
chCK+omwmz48aptvF86FREhyo6UKUKWu+ATWn6G1qMevZtAnTT6nmlGXvjuI0tm1
K9mhwsa+b7Rmc/9WahAbZ5ZLaY+6MzdFBnS57G9ocZEpdMkD5T6UArBh7KAvV3XU
fbaGDBjghCC+LRKrggOkX004XIfWzBswCb4eolp8jdw7ozJLg/fxjeIBmmgKMRs4
wU3Noy//hMLR7DnJcSieEO4Chxsgjeztcqqqf4FQVbeLSGj61uKJ7WDHZKOrTJRm
6Yf6oGMtcQKhJdZMf8qll15fo3jjkLfkqHDYshLOT8Gr/hIUL6y+9e9QNgB7AKvi
p7GAWqN8+o0JOMUvRskW72YWSw/t601AjxobwGt3SJhZ9cL5gxfp2K2h3X7O+uS7
rs9oHct+U+5+LKGnQmgJh+5w6/HywUtvrCGrMducMX/ScSIxH9N1kt8uKtdTJTN7
7PYOKvKEaeEEwtsTO5LqUBaSBYi/pFk6qalLNryCNM++KFUB11cEwpLHY1KnfhzV
xSB/V75Hc74P8oakYh+L0yJ7lqGBTzZlKQwXLhB8VCkAnBFBJxXqLapYJkqZag+1
ujOYqbTc/5r3xvMjpZRLLPuNj5o/mx8E0H2l8yE1ijSCDHulNo+MzMbzxtmCXBgR
PIAqz5Xd0Yp8FnyEvTPnzeFIhDjd6uN35hnzBzD6phWngVGwCYepbobP6iIl5HYG
Pg41UG/VE8RXGGrHkjJk/ZTSv4OAueFIAUU9EKdfHtIxqoVBtmCffIpGHzko0wyY
l5kqvBxOR74XSxGMJ/oJRfMpjaRHGVdYbEuWGS9JJbvjrdpFyb+GoNfQnThbUyKu
lxmGXobt1Ommvn3C7Y6JZT8+fcU2HwLo/0rxeMjQy934wx3t2v9EJc6fbJLzWX9V
4+dQfp47YDVV8rGQQUhLkZKmVQe4AWCz05e3TE3BIAfTKyjlFjYp9KvdBJNADCkt
JiCGoWWVxlAdVLz20+HAukBtVCh+kahF7wwjVLEJ6+AvGZsQaxtLN4VZjMdnUyc7
dgPwXRj4/FcBfKmqILJbQ6kzZa6CICVRye5iNrQGntmUkFQ8SMzt2ST91rq1RiRB
o26FrIXdAwxmpgaJMyEyshH9V4P9gYy9I2USoK89naDogmFqlUVLLwyhZapfmEVy
YF6WiYgUGdwkWzDVAjA5GcWhy7w8sAn+KOSO/H6Fp4Fl87e+ewt+J2hlbaaiqeth
GFWN/lnM1eRP+d1hfOrLgi4J+0a/poJAdHxMnTQoDfN7YP8T4Hlm0dHeUa9KaJOj
w52IEGwXYpjZz+c30Itn/Ixuhe/M4lovmmUVrJnEwfPnlx01I9fIivi9UlZHiWGH
wrB05scDAU6oXoUCGfzLp6gXQxOUbK9kP+Dnyc5b3sWDgbap+z+yVPb5FzV2i+/g
LKWDTHkYyORIInZHvDDYUB7avavhfByOnx3VYEKrzLbdyC91CIMNQRmLBi6UaqE+
brbB2S8P5kJ1w2dXA7txf4ULkeTT7aVaLInbZ8h+vhczk87K+zvmhsXsTEap38QC
KcSrTV/QkMIdDdJPwAf/nwWFaOceY2BIf+spQcY2vj50lqa3aNB++hSY05xafneW
y666WJeWfNCfxdfGFBFN0W7r5xU5djdQuN40acJlL7EkZ1YkqERvzOZWOpoqfvZ0
NpZ50+PCVSre5lHaD6R6JMjsEx3dtCFYZ8LSBfd8CUT/9bkwftFtjtDNKfsCR1RO
ir7kFVOvETxh0ARrfJh4sG375icvBBlVefueoTQJnUda9+7GsGzd7aJ2ULz/fooC
c0Ygcl9nqTz4sE2eRRtzPHHVu/4sFVH5NIW/7NGsgXsRuHxcfJtiy1TT99fSWVFT
qzKPCVHMQCCJO2gbt2U1fXo0XLZZ4AOeB5cxlnpq0cyPFaMCSjJ2QJ9zvsbTgk0s
KPswTI7Ewhsg0Zx6kmuuKjOAu3deDgxFiE6Vme5JP6yWqPVfSwqrBykU6oT7ekWi
q94C3zRAvTumM8vFy5kfzhp9Xq5wcfzM5+zzBrqIKpMTdG1qQPrfJtZmfV/fK+7b
fFpbVVabYceA9eFhN4nnATuIAZESGtnowu0yylFMuzud1Fxr26vHKSaZmOWbSL3s
QeVfP7yQOaH0otMRkY9g8SXEkuDF9haSHRZDq51S7uEr+JIK0jz5hz0NtjCMsex2
YM3e1U5QviDeyDcLVKNMpFW2kD7NI8pnryBe8cOmRu5GFWTiQmUA1jU4QX8K8q01
WWsRHCW+/QAPsdtNO/LME39uTGoF31ThmBpR559N4hOZlLe24oMkqcNTJZrmoO0r
dFdt36tNc7eGb1QJuJmIaLVUvDilLUufzNoNHQvgXlsMYyfUfPeIusLFzf5Yh0U5
IIX7+W/w8XMAOCrUXudjWMRaVRq1ip0Kn+o+wgaD3up9x/LPsYkjpBScwFBbT76g
qk/jvEitiHt1GSAMjVuSqCfWwuOTWdaObXP9N4N+BMHOxDENcQuFIKm7pDNvKqHV
Pw3FVFnE8FU8g7GdkUWthvc79nkwGJXomcGqu7A5WlOlFvyj0pVZPDKCXZVpXtC+
LzMvpDpOyZLyUAuAiyNvIB3vuvJ8LLcQVINgWhF6owttewqsXIQjmY5u6ZlW3AVp
1Gwvzm0VZZGplJLNm0+6pyCaacYHpGgcdYWmrGVLKbCnYg9Iie1RceUEhloZE9zp
25Eg/bCBmnfZSzgcoNMHP7Aw27nISvlgu8mcZFP4UMf/ok/CZ7P+JwC/m/C8tOc7
a3uM55zRXfcfs8Bnb8kOkSM4lf+vNdS6HaTPTp95XQ+VSusFJW2a/+cgqoDf4dAk
R02/bZft2NlbSlinn3+/MvnwTAHiz2bkVrwhMn1+dpIJ+nK4CTVPmCQpecgS4FEH
MiIT7wX065pi/2h/wLsjhLTel49f+dZODnrdgX13zSv9Z2aDZzYK9jfHrvqUDcUm
WjYHZxld5Z0b151FpGfbFoWgFby38wvMbO4+fY8/Gfu+h8Vj/EA0jg41ldNF9itO
87YahcBIgkU6weUP/9rJm6BgY/usOHAlWji1IT0TevKIo81eTwnts+Iuz/aaa6vg
5xmi+kUUKJO9tRm8DQVcl+BfxWp9gyUN0Dj8er0dG1lD4xJS7dT/gSwQZ+Ojl2qV
zDuJV6L5j0AjMK9u7wDJZhZtZneHAgOvietMqhsaaMSw9/Rg0INSTy826ZvrfjrW
ZIO0h2rVRFPKyTkhsUQBkQ/QMbCUsbvPO2yhHyVbMPeSezVSXLfe0vNHx+CsVPY3
A1k1BB6j95DYcRiRZ9oSimPaOqTHFQ8pHDFX8Iuc/YIz+l8eJc0MPplcAOwDav78
FZaXAuhBIDk1Bb3v96fS5e+XKRRABBg5mcEb4d+qaSNlqic/p5K0FRtWQWOxn/au
iKXjrDIQgrDAwM2MJZkjlHZi/9zN13yeX/YhlNDy+kKbwwxrsSbKT+6Fi20kWKEA
yo8pNPeJpJBgLqb6KQ9MiaZUFOH2OEM743n0v2GL11hhb8nNly/O5yvsP/Vl0XVj
Y1ieYNX5tDCtoclmaLixJ2vHbuIsngyu28g7/sTWLtSNXoaLWCfdsdcqSZJE4Vgz
61Zk3HsajwwloVGINHXuz4wWOW36wFrORbOGc9fVynWJaRqUcTMSAIKbDjDwnvp4
5dAT3VafGvul6ssqbd6nYbQeF8/kRw6djB9dPcswszWIZqx4KayBd3RPBGsYfVmI
wT8DbarV6lJe95z+Z9syExyklYcLNRIHpSNYQPiqMgm2tDB614Vi6aN9VOK21+FJ
hDXGL/ftwaadeSIRd7YGn8WupQcKzfLcS4ZQ288A24odki7vtvnWGlrT9WxbeMuS
l6bgMs8VAiEGnnAKZ6uz4PW+xd0z7Ek+szxzm64UV/p/nLDbOgwAj248CppqTrsE
+fVzuN77qp14zUa5GvUqfXSt3W0ZASIjTUpPZHFq71+uaIvrtflgQVqYhVcBLIol
d12xoqj1HXpjduFXEm/gcfkiKeTeyYTjFrXDyULmO2khguIV6nidsVktcDYKx9HI
893hubzNwHzfsFQ/syQ2+7ag1ZBFDWZCLL9eyiG4TSoXg1SwqR4jRJiuJL/zzyiY
FVmvk7jmvllEHruy0wEmK7KQjAa+/Qpmks0rfp29vPZTKz3F0UHNBMbzUz3LTYV+
tNbDEhYbnFZQHWVqSSmqFMs8fYRXQa+yWbsmrjynrNxmTFXFSgy2mlTkL+z+QUKV
rAEOpV2jex0e7zFuGCX7v1262w+Pa1+NxcWm6jLlXS/G+Zpz/UmBnTYU5SsMxmid
HCQFZybutz6GWhkb2A7S8Wzh2JMepadTayX7g7zbD/JOzD1latEqDIwP1iN7j44G
gFefcd80B15qJHQqh0YyZ/I6JQ4uqJebQqLABUoTW+m2DvgwPfyFEZp54uVHVd31
qrQ98wYsFQqlDqKz6NH5XyA/Yy5zDHEe3FNmCccz5vKino553APVgfmtickHkyIZ
5dZjTIEs1XsEj5vjFdeZgsSGf5LUUXlOnFUg9NZnXWtCnCrl4R8x4fjMQEXk/F7C
qiOmK6xRW1O9v6lKT/sZETz7bfQym4dX9jF5W5TSHWMORLKsZ3LoXka6ShNt41mV
7R5ZvBoPI6ypJiZP+tTeihqV95dlelau+xKlGalvP5KqNm0fRSEpDJDX1mWsehXA
SfqmCMdAHb4kyRmLT7TVniB3oygEyM9fRiFCxFdpcz/hY0uffeKP83Qq2Z6v/WIc
1V5OrcckKL/1LwA9IunlWlKRbFt4HnOvqXXZxVe+DgeaKCZRZdJN4DTkdqGEmWSY
MkfPO53n4iiKaDxDxlv1o9gguDUFXis6rTA6feBCoN7RW50kP1JC4LOCm79g+pmG
Dsgdc3Hah/9epjifknmbGN50cjRG1A4lluVr4LLI5/lUFQ99w937Z8n9Nji+sPVe
dE3dYs1nDlS+bSuiuVq8cUVFaW9stV0LYmpEJ+aITo2bnGePbOXMpK4ADR5rHgqm
u3uVk0xY97Tg9BHENdHlZiyf9crk8sykwNVnorVU2+WzHCxn9RdHWvhArVCh1q6j
Ddl5gAYwSZo0ViMIuxtW+zffIoXdXzxlpL7kFLFA6Lo26cSXpmkw21bvDL8MA6jE
NImpE+z2G6ET/kkM0SwNauTPMTq1sslY7p2oWC1fysbDg0m5uGJp21mv6TAlP7xj
RUO+jyULTBi9L1FIZbqXkLMr20PXFPkUv0ZPaS740fXobDHFEuuTeFKjD0CqpJIm
Q3s7IeVndMignMZAzOq+Sk6lsqln25Pgq8CCI4yGBuliHr15QhDQ1Z5DW2NFOoyG
9Gc66xwzKHRyP70Mg6D6HRCpxO2k121eUFqTMhdKteCDU7fLfaaeid4GWwJjRa2t
L03FfXH8sMHnA4cemVaviCR+u4H3p/wjF8hI+NyGW/ocTx78ximxcbND44PAp1eC
XpaXH8z7786i7buufkrp2FUjomiu4tb5vS49/bHkPkGoMk58K40vL1r9WCQs51Sm
InrxB0wivz6jttvf1BDGlLY+7vfymER+xdCwdr/HJ8Kw2bO9pQFJ8AlFSGIsHW8J
GbiIBN8jOl9lwVtdg0i2Aejg7cNUjf5QJX6U7ttqLyT+lBXv4rQCEWGg0x+JVYGU
b2jKnYnCxxy6O+9ji/V9YEgee4ihKTA96SdSMAFtaNTK/LIpODSd3roSeP4zIijV
eGVKnwMBlCVz4qv0FgesI7SMO2rA5Qt/16l2eEDuTeL8ATiI/ysftTA4mALB2IhH
aIDdOm+PUtau5RTL9Dq+PR7CDajEXFx9O/Xpw2h6oOyNqhfjWcy+JIBv8rACmoDl
n/wdLp2kOXfp8So6Eop6KN/aCJBQm+MaoE3Pyj0J/mnc0ym01/MqOtTXeJ4OlCm8
29wuk9R9Kmn0QL2LPfF8nSV5tSkAAp9Ig6Ab0Ph5mweICeLR53MsZAwsVqU8OU+Y
jvm6stSoRQ02ISkTmYRyfybEonpKLUJHVNUNepIyNXXB5ue0JQV/5o/iQPqk8xEE
NaloogZQBcPCI2qyTBwl8wvqbu0k50WUzAkgNdG3smv/MeOX172hIQdRT7An+Xx/
b5wDyidoMwL80Jl74famBRlUPC/6UAQwMb+OpJ7fPzBm0KfY+0kD+hB0rOnVDunu
3Gc5RmWu0CHTnlD/WkbPjhfBBVCBoaxNLsAlvMnfo2caQWyL5YyFVeMTFXX2D2pz
cfXm93e54/YYOKvNuKiGwEKumwg8TRgKU/KiXlS3zOHi5k/Q/xfEAwwt/lPQp0T0
f3cp6zuoL78XrfpnzBWTWbJzuTJyaYZQ5tAeFippg6b/XyCAfYIvr0HY18jaLgBP
TsWHNyO1qr0Y4u1saelqpOpYCpYArEgKysWPPh1CWi7BOWNussslmPPGKCOL5Pr6
F8cxVGSbbOQgoorNBXCVyXoJ1AlWduQSBoS/dZPGfBSEzPnhuZYlYsbz+Th0ITrJ
xgWZb+lH2GQv70Mg1n1SoczOVlCc+s3uzLF8Rd2aBk8THE3A9r2aFNWRF69TrsHr
KEPRZHc4iwZY0FKhtJLcnVjmuFtYyoyjoTq4/5mbR38u0koWLKbqX73x64QQUWdf
VDgHxPLW61yUwtotf4s8+OWI9vXvU0ssJ07hh20W9aL4CiSfba3pTPKizAP99cpm
GugdfQvhzwXbbycp5t2JuKUeQJ+7fpyzgLVzruH8eh1AlFb7vSDAov3xFc4wh21Y
PL3TCXdwMkAVMNiTQUVo+N4/kMeVTdLDJIs+OeblZHHSAR5CfrE1MeoJl5FzW5BL
n20XHJv3Mg9Ihrjwgo1+LfmJt8JsXZn4Qz+9Z0/hZ0r4wst556iBV2DMfCUCIB6N
WhntFJHuGinumi5qTyn2xwFBW0bFgAHNl2UhT/7IUuws5tg2mKAwcrY5wM7T/JFG
iPikZkShXbbo9+kpcj/iefii7jg7W9STEMB3KMYX1mwz05sJMOUkst5wia9z29aW
PXBsPNmVLXHGePSO17Xngu32dYbnMKv196xLhGbkL1wy6Z5LTjWUyCNCJNPTMZ2W
3lyRWbCx9+kbmCTcTZ9LIenHq4u2cPlwipfzJfvEQaUTf07k4cDLbtY+1gdes4Zo
Vk5ZMly81aKh3YqerKDgHD05ljnSEi/jj7IInJjOhbHnMKH1X6kRjeL7jI64DsiK
z/r4ySZ6a8arFVhXwaZCPfYh3W5ZjwazTQa8WI1YUnkZrvAIpvhs0uwEeeOUkzvo
B7VcdVemdrhDsRx6oJqMKGI9T85eVyHHCMMY7IgU2jAug+fo3QMr6FHnRj+MYtcA
zlBofQajIeLVq2QKvtI1+XxAbOsED2aw3TDiJsa0T3gNQ3dWpmnK0gL9prWNHK5n
Nbgt3BKnvTf0ccD4yV//hVOyIwx5nyF4FOK/SoqjfqkRKwWNnIOXKfqNko44zjjp
QPlX8HajzLK7JR5zKynHjpgbrZD1HvyybmlXZyr1wkKmoOBsDYR+ZqH5fJPk/vYz
dwqgol+Ir0n3ipgDZ4fSuTl9lLo5bo02VvGWyWgLes1KRYXAXQ6xsCJ/L9+9pXtA
7cuoM47mRpHeRYTV5GDvHidVf2OadXKxdJFEbB0hRTSUb3XLfXosnyKRp5rv7v+1
BflLjSVNQYd7DE92OX7hUlNqeeShv7Yqk53hwk7mGRqTu3PcYxJYqE3mhfvppUuz
ZR+Xrxlt7V27t24S0L+d5oabtrSh12SUwazz2LoF6ensx2o/CMrBrEjRaKs9Wd6W
6pOfOH8ibI5aZlhntWj8VSoDCRr0CMKM5VW/J7pk1UM2BriRW47suCv3fsZU2xbG
4nXBYtDYzieCDxswbvCgesw11bnFCf2hrl1ex0DJyreei5ZPuvZzaHifaOs9OMEg
oQVixJaxBx0dR2euz4ZkakPYI7SqAIPkXPtnuS9vUzLcGc/UiA13IqUnAWltwaln
gGHpaYElQkrmzv9sKcn261MOxMzq5xxQ3aZqNdgIM62ouIYb3UTvSEYmvlSXZlTP
UeRx/zT2Q37JRRvr0hrqd+oichdcbnp0T+UTbxQVB4ROPfrmmqUYoVcb/jlF4k8L
ixeDPgkEEDn5VvEpEAFH4E2Uyqe4hm19EuicNg7ALG0q8WLj6govuDKZ2fsfoqEv
syZDw8KO3nfh4I9+FFGtXwj40aLBtqahBSteHduKfRB3BtLXXhyXPDXR8MGmeYqY
sf+FBoSiM6XIFx6Q8kPz8+6OW2rrLkkpS8NVdWlbsMxGq5QKkhInqtAX7GFzVjSc
39u8WY9i71kJMvPR6XpEW25Axd0wngbguaepeJ8JIcPCUnGqx6fPhM4vZVwOk64y
r07I0X/ZqbLn7ilmdcrqwfvXVQnG0/pcKN9GKj5vROpLHoLrSF7pedcIgjVauDgG
2LIDojeY2VKMr5LiVC2uQLrE/7fgR+hLysfi6XurhCsHFAoyOMshhz/PaV+orWr7
lDKYTmh+D7l/oIaLlTGriEa2S9gktCkIYJY8mBuYUAzTRYjCbs0VjNs5Ox5YIdNy
2XFvc5ly3hohZezI/b5pLou4KZsIUR5AWHtnREXKIvtiY0bcmmTlfeRSeM0YBgP2
gi0CaLZtY2IEG3nhMF9GdFysvEnd/oGlRMnHJfSKegAU1LYmFgtzF5kdpTEY9AXf
tLBHRTr7kW0wcW+9WqDNKZi4nodZh+uXFnTnM0D4Txq9TV2XqqU9SjrCFyuKMmFt
YjIpIjFksYrThXNQvQDJx/dp9IZKT3Wwl1XH0xA8+UhhrHZybmEOPFF5Pp85G4wn
QHgcECS9M4HKjz8QBvzVSw73h+JvqZbTc9YF7GpxY1VVkkU43IcfFbHE89u/XC5M
JMU3MTM+LxC7In9gVddfuMVueiojzGOSuGWCYko77RAvkQDUsPgPijvcvEYD3Ilv
x04zP4sq804ZjtsONAO4M7We0AFGE/eE+1UyzDqL8Rft8r5rgO3RMf5Cq7mcDIzU
06uwNuu491yxvByD7JDz4u0Q2ZST/2szDvBquTlCXmual8WaSdK03FfxVYPAXmyx
Bs7VtYGa6kykJp+IqYMMS4jr2TAqXPTrYDTUtRWvvWjL94j/p7MRpQqN35r1DD8Y
wXFBul8qfAB1soCJjV4f8czEAVLR9aNH2eoEkxrlDvTTi8StN/QkcbJbYcnU078c
LtJ67AZ4zUEf4RDvPhBgD2Ejxv/BvxCxUwBe4MkrQ5p5BVWCGZ9EsviUvD0KToCB
BJ6MMeE6kGHlWiOF8aFsIKg/5W8LdHV7zUpFXeagnlDVKr4R2E0/63xc3O7migP2
Z2pHpqWpRbhnsdtnABt/YDO+LJgfJr7Jjkk6PlsKzAGzchIQx6aFTCkyFaSLhztD
U15H0VWX9TDIkrLm2k94i6KzbfHEiAi47rIunb460WyuA0UkNr/KxaPNbhoqRlbX
KTFQu9qMn/5kG8M+SXhyh4yC3i1gBFr+K25cjY1iJswBXEOO9LzBc5yjCUskTCQ5
4o83epZaGCUb5t6ntNulftXO7eBsCsXe/bvl16mpPADymyIIzQqyVbOZ+sPRP7qB
ovw19CeGKSdZ1DMTR7aXXTPG3vb9ZaU+IBcTQZ+8LBgptiKlNT8CeO0B2qYfF/nc
T0CvemvAVVI9TUrtGAbhjFVY3rCFwVa23D6SEacmQP2le0aLe9oBYHJl7iXqSBy3
JvvG1b66ALDiyGNqT41uX7qlwu7xVmyUMx5ZFtjf33TNnJQt0uI1VZsB6qtz3ga1
pklBxDmgY1X0/XOuJQprZJFhNLp7mvCQuHi9k5hJtuigSNGPnM6vHrSbAUK0/Fja
gjuEOgICUwGWXQ3aj9OqWKaa6CqII3sZJ7MEaG/sgYXIrEX7OXb0vn64Yu2ImH/w
fxbXXMFlkqhbffIT9kjmTlSnCIpuP1hpLB8yh7bSO/lcLrYArzq1dQighHJiZHAc
ljePi8OTP0ef1FcDcPS/zulCoGnHcf3FSG3ng8buWqLFKDKjqQY13OIl+nax34HL
lRlVbO4Q7UoCW+Izcxy9Jsyc0nIeCZ0sFFmiVKuPYwmc+f1ZsdPcQR8iKeo6JUhe
snnpyaEMWQ9xiOSa0kKsNuGdg6EywUrYbaNNa/+7bEhXizvSxfA8Sm4iwmy0t+1F
+ryDhS9myHcVUbhwHTrPGbK7/K0Ivummmv8z0+xLpKreLiadmenp0OiJnBPpw14I
oLmWoNqZKZiN0OhB787k3Yat5zWWJB/aJOjgrdukODXbngkunD25+HSvpodarE9R
srLEA6mNVbWpKsKKRjTNJolI0YfkV5lmkeqIITKOU0txP2yjKXEa60lfh0CUXZvy
KVI+1L3CYF134d9C5RE4yDGt8f2nT+hpAOO52ju9WSVRvpIqfdbxeWZqxrtx8gKW
m2rpp1BrjnGJ6uCrwIzbpVIuiolMip/9jvSDbXDxlgLuSMw7NDWAWKkFa3qvC426
GeztAZpqfMARsU2W+B6BNNVMqymgw55OzmpLzqbTF/Msuj2KZ1Jb4aARx5QnDHcl
cC8zVaUom3xXXOdXtKSNu1RD7rojHQd6CfxS3E8JW6AWJRoH78pD9T0p8yyI0Swq
lFdgnSX/1x7zmOowfjjqoWXK7GJyiKwMcPJcDPlTLk2AqrnDFAjA1GEpkNg5YbUc
kC4qqKBu91BfzIzS43RKpkjStm+vNCzNBf1sg8zhPdV6yI8DoFlCnAio1AWVbQB1
jo86MG6AbN8SIGGgxoOOCgKG4PABKDnd9r4U8cXQ+J6bf8Lp0BiibM/9nPy7Cu2w
Fy0NTDurGkq9eePIQVdzhYSiMp3n83mGNlPPqmu81kkQXcGpj08pKrz9qfywf9n1
/1befZkiVVA8agDrFYC5GBKhWAr+ujXSFirh0ahdtkPAP9udhmLi1eR7DU2CD64Q
8OiEfYnlh3+TeUuKCaWYRSrqAomxLw/m9eEyDj5PcVfPlG1itwOr6x41Eg/lGQiX
EJ2lchmdcLYgYGDf4RwEnpB/FsxTQGieXj3/Ny1xF3+NQNJlpKmYocXGdspoB33D
GNP6xUDxwuBbC49wzBh48h+cJc+Vzi8jhcI76Cqw9DthzK3egKcq022F1kmaN5CW
KJTqpZUClZGvazfi61CNT4oiMX1mugHVJnboGSdW5GmpL2jGV9YQEBcYx6Ev+t4+
6ti7y7Wd1Br0EPXcHKxJICHV9LUKBYQExDnNbn/mOhxIjneOw0A7e9Yi553duGHX
jIVsVrG4hbgGTfufmmehvRpGYQtlPgW2lQGpHwIiBhODpaIyb1d99YXEDTRQ6cmx
ytWncLHLLfvQTMMoWUCzfAzua3BteNoJ/eFKVx438h+W4C1qt+LsQfbVThPvkl3Z
Xvd/Pf1TfRPyihYuce1cKTfz+uu0FjzesvFY2vaIp10+dMMbkr+3z8e5Mj+FN4C6
eNhk9Ku21m5ObNDg/hHSyYcuZzKEUVKJQDCKvpUXSLsoLWqKApCPlWUdqVOPaGXt
zt0ypxZoxvcV/0SyYtFWhzblrtqiQfNzAAgldaiPO4OeD38ZeMohBuJ5ON06IYII
43rWH1PUPagRqYjXZzujRR05QllEXTuD/Fo5LTT0zLjRwwhFjS5jOV0PgoSfZ68X
QYvnKFPgw76ZIlKFywCLD79mgJjVDA/Ky5l3YEid9TPpdgp4hlQoURgFxmZzl7kq
r73OBI9VnTYkq3v2F0FP/8IzxaF5Rwvwf5ZNdft9tAJ0y08qF0rGSHOKRwOriMnK
IWx9pwD/bJZTHdbiAwtrba5LJKe8kPAym06ch5BtnfbvU7gniuMRURSGaIM2e7YS
tXyH0+W9j1BlfPqnW7gXnRpeYiTzSE0bVEXPFEaGD4F3Vqh9heXfUqK/JKF9RekA
BNPQp6Ek3wWSapr3ViA+aUZLK1MPCaImOLaCtSwz/iBizGXb78BuapnCa6Rds+Y5
OzHu+Ce77wJyPoEFR6IA4/yDwGLP9NfNU2LGis5wV8eFoH9FdK7JO15UOP9AzcL5
Jy3SV8+9+YCHZdvnB9793IyVtKLwOn0EfOS6sqQj8FdyJ5Sd7wrQ+19yrLT0lsvQ
Mk/7oMc5dzBT1wm14QeLFPhp38tsEmYxdjFMAu6vu3CMVBVH//1Iu5ApFkFNDLWN
cwni+6/5Aoy1q9YsM+BlOOvgRkbqQO8a5UwYUMiq0ZWNygP9qL76YdBqufGe9vdE
iAigkTl0GW55SR/MkOysrRxJxPB0v1ft1eIE8olmuUQVdxzXoLqMCSG9f5xVbjw4
UMsOM96katTlAQQDtazFnImWyIYCpFllTvx6pr2Y2zOrywJ9fQValeQkvmCqTae2
845yMTbknElZIwG4L45oYmMmwILh2bWgARWvV0DcfpTAidwOYOSf4kjgmPpLJ9Sw
oCn1UwdXpYlvQoBwb/K0nMk3jWlSnn4VahYPZ63K9giHRewMSo+68WeyQDQaFrQh
Fd9WQ5hrRMW6XxFXwv1+g5syM9BvpGFB/ogD6pIBeQuaPJ1X6FIzn+36GMmvK1bF
ncQ47/0pYNxz24p3HpI6AvgiIVuK+mT3YucR2PkPcYzbnuPT+c+TZjMQatb3SPgz
HRmvOlYRULumQ1JxFfFLexn3RoOqT90sfePudxVH7FCRdJoURDEBux/m31X93lrd
W2nexhssAzNnLcmyx26NyW38r9UzctSvXR76zLnXmflL2anrk2Dj+rZ7XwvrqA1I
b/i5CT1HtE/wMav6dcjnYOjKu1BZ8Iuriyor0YjDPIVeoQLiZUXYpjOZbcYvkduT
A1miKDeyT2R9S5zzJ2yic/sJ744pO+rxKm9YRiQAMxNSwMkZN10Hk8B3BCyi8gz3
tLNXRbgSfho9XbtV+niHQniyz0AZjQP2mbYKWoNZSAjJ2jrBVnTDx936JyoPMH1b
3syGbh+F3HpJDQZKzNnbcKJEJLn7vPLtPrRSJ2aYm+Cjyu6lqcgCiolreEcn4du2
+NR3nbnbKFxqIlbZ18ZBq1DEPB0o6uyYu/DKzH8c0FTqck6iSo9YkVRjg7LqoPUF
TQGNB8MzVamLh1QN3I/H5A3rvoMibZgM7F0zN/qTKmxieQWx4QiNoFo9AHo06bJF
DzXDVn7o1QxSA423UGb6m3FSDi+p5TdsMpo5trybATIYMAtsXuviuNl8Gw4uLG1Y
Jl9urPL3Z9ssTYvgRwNJGkgTDzVjpmX6e7ASn/Zu/jlwuSFqI65/OAAHFoqJtjin
9y4POAv162cX72Tj3VcPmRQwdXH17pat+zVsxa4phqgn+5/yBh9ASnCH+icVzpTF
nI6Vtw4xB43GYPWbDZCsFiJ+zwIgkeAG6a1IAn8xt14VG6XmTUnDqyD3dqtY9V5x
5kP0IK35TikfbiNv8N7BbxWTUL+Esqw9lxSuxxRxIHMFnKumrlQi+AUBz8fEPl29
3L1OqiT4kZmU9f45r2vGpDPqrz37teLpWrrghHAoHJp9bwj4rIPoykgnzuBpj3ps
n2b55nEwb9zuW5TdF0Ee5JXcoSgU9Bvbx2pC7GVRXKkf/v9D/NqJGbKXkJqDewQh
PilgDaOh3DpEHwpx+bYpGkHwpoKpKubu5hk4U3Pe4+F0i1hdE29Zl76daswPRBX5
rW9UcrqAeJHn57HJv0THE7lIpUnnL+kwqV7ds+VzL90vtLYtxaGhbqxWw9+RZpBT
uD8NdbcpCXcg4stOYMti73sXxDolts352kly2R3p9Vt9WHA0MpNdH/ksK/Bpw4PU
w3wRRB5JHmqHHasfaMxt/15OVcQii4wW8v0jIred61cEG6dpK3kMJ0Coe8m/Qknk
cmEz5fKWmK4EaEs9xbHTQSVXJBW8vKJ8O00yLi/4zcREKgTGEG5/RPpk1ojb+ZlG
vAKPvP430zImDRr+oSz25pr1faoeGONbFtF0CIx9dURymXHAL2Bcy/cWS3/IhIMn
NahD8Kv5CgUOtuQ5ODvxnhjPscu3c2TiHIG0+mpcMFw9DIz0bk+srwjwi1D5VWu9
2Af5aZtFHXmOYTK8U5Q0dGfGNFKNAd0P1EzCHj+1L+BmZNcPAbTtKbTPC4KllIAR
Uo6zYyHCezXVUiwJOERDEdkBzPQlG/0hy9tfr4ghioHDA7sdu1/B3eresFawkP5e
RflUlzq0F1n8l4/r4XiioVVJlgvze5cPVrW4UvdewsP3uYziZMMrgFEN9zFegqpB
SH5LgGWL32mY0AklNkrVnkBxM24b1WJn9kwJThTfVC6vtJFe8iH+3kRUCX+8x+Dl
OAZPzqSWK1FMk2tcD3UmIPR/nCbkJLtUzoMnBOqOAR/lUyqqQjekWdBHzYkrgrHE
OALs0Gn7cPYGXoYOBMx71ZRGer3TibHDRTa2qNALHUE2XiPAiOK/fYrZkDI87MB0
xtt0hEQwd7kjDrDmGiEnTmz+6oprKUruTJwWsxioQHFHQ10Sr7OWZcz5NWznxxYN
KhCBsoB2l8YchUE2q+usKLzb3EPth5HUOCHGK5NECGim3jccgwr7cVZBip0b2wmh
9ZfmNM37vlP3JmA2MF7l5DYL/adD1lF7wcxIxCPwA0K19DwazW+cwPaUKqxfzrfo
IaWQKfxRWErjNl1A+Wnps3D3jIukEJHApIhugy+m50PhCklO70F5s8XqKOkvzwiK
ayuq6p8lMWxtOAJ6n7t3g9SNEvfgVFcU6x1Pbob5+fPR6/oL4CggsnFXHuyewvJ9
0iKmnykavS3sGnK5OJA8KQasP6Uy7uGxBd+y3wLdUJ/gml3uXSdi8D9WR0vRXQhb
wUkJx7Tdqa+WIzHEf+EybmyQeNZSA44enZH3LDHiYtuehDuXs6LE6jb3XRW/WORH
fJqVy2cUOAO5WT0iWDnGZbqY3WNfRKcKkuomj3ZVfnRMyBe5TZRMik6v+1ZUSJ79
eezk8Hw8OI+TM4aBmJbWGRdj+NWNvsSYoVEa112LNEYrJIIaCZNPgr0FXsYg/gmX
QqWqWAmEozot72YWY2hfN6cI7ToZF8hXtK/TlSZ8tTsX5zLdoYTRRWUKmZtwMXVA
Jk+mtUizq37ynPULAsO18oOgWdXi/Y/LpxcC5eNFQWKDpD5R+B7Akw/6KDA48uZT
IxIllQ6OxWJ2EgTPWn9di76CMLfdY3hpT9uEKwbMrhSTg5MDhzlf/kVWHel623iz
Bvk5r+vtUsnWt2g1tIzMldv8pqyT3V6vA7Zg4sSRg3xVISf0YdLRA6JZHkLVBUOy
1lhqnHNwjIQk89942Wfoge9OxFtL/5WOQWH8+thtbtwXFJgNpT3eKvvmF3aR0Kkp
d8ywZZtJfGieeXewOMBk1jxTnYhqh0T6iep7Te0x8urenSVJtKym4ow8PRjIBpJK
Cl+lEudARSBEWGc6coNTBkxwj3WcmNPe+LI4zPZqXjKMbCHOea8sTFgx5ekqCoxG
y7GSyWSPFaYaV1wxbGn30SW2XG5wz+4V3LllzXYTU+p0nitm1xgJUWZf+zVXZUR7
tK4F+A1Mi/kVjQCj+ZL0H8F+qi6AXGYmeYnMBmnmvzBBtECIwKVqPHAB501GZRj7
dbYhoZ780GG2klj55g7FE5++GvJwjBI3xRFeniKXjX9QfndAWhjiQxaRkKeH3EL5
kdyNY6sn03MwRStX7Tt+lXJCViwN7XpXW8Qc0K/iacBOCHQx5deOtij9Dz76ieuT
o3hzAukPZZkAOiMLZvgygk79m3P7yUyh7rCSi0RWT9vtxSPa8PlVCnmRAih2Q+Vv
ngkEyLm5lGKh++N48JddPivKg4EvfrSLGwJS6iJnNf70vAaGCubM1i8ljBCiKO9E
xq/ad9Zarx6R6E4QA+0AnWzHE7+OTj/UU4ogcL/hfYPx4BV8bQvxyfGeKbhtnlm/
3HeFv0zkV51a6XhqFvlHX5pySFiV+DPBb79iBzqcsQQZ5JMb4BZLPrBu2Zd/0u8m
ETSAusr+mOlCDsXxPuPXL8A+VZLLyq2EOScPYYvwAqIBWrAvH3JyvShldKDO3e2u
Q3TWYMtC6d7W01W9uVaF+WUQwhAht3h53BKwf5bDMDohO7bCB+0gmHS6XGS9KqoU
nm8Pv57CFAYl8Uk2reOkq+ZIw03fPudCvK+/sEVsMVU0rhQ48VE+++dknIO4MIdS
uMbzmhm4Qbhm4ctAwftH5jao20qRQbxI90PEK8JxNny/9jUXV8HsiUWPgl010HV/
FK/sRCEdxEdytyP4w/9k5eA6AleGJrTH01euhJWxvGj8BX8wxZdnTUaLnOgMBQQB
lSUKr+gTHQf2vfTQYwnFU2unGb/H9I0UEwc/WFsnBJv0nQUAHoSCQ2wqeFxOQx/O
sBo/spaadofsxXPukP+3mf9yGZSAxJQxT29Ih8H1Qq8roIurec1QLye7mr57vshL
U+wrKrnAsdLgIHnaHaLESpQAo3NDn6BBsjNjFMz5fOsKG5UAAB23zlQbG9cxA93w
1qW4w0fTb7zNmbSAJLPeUncFkKwoXdg7lW9SEIMKjtgBNCKHivEpr9U25Tpu0i7/
F6mzFqvXeocN8W8i1msONysvFb2PRGdBY+/wZOx/1KHRldIaDYj+gB4tbqkfPc5V
utq3/gQEYcKZWfgO7B+08MOjrwpE79EQs3zO32w8VDoa9aCg9E/tbBM+pkJlDpLN
c/Gcop847OPdM8+8Mmb++MLBRUWHkLARGtbrsjzOC8jWcF/fpg+fvP7P6N/uGryQ
3XMtVT+OGhu8Rp9K56shm2F71zK+BtYKJns1q3SjBC9nZcAmhayFJhyFlY3lZTez
6h9q0mzE5WYrfV2jq7yn8CzRMo8UhlSNhtdX3joZplltaSx6G03OtvQEDQyfHY+J
vgQNYYioHDbgtDxz+Aq4sYXDWE8m4eE8bdgsuLkvghzyyCmcJ7+xfTPY8Pa+RNSv
quB7yHoyq4mFynKDLIx2KDCwJD6qV3WU8VkXQ+vQVSUSMopsOyWo82Npvc2kmWM3
8tMVg8Xt9XauC30wHCa0F8fVlwnrQbrENU/fR1rutGLTTcJ3HTB/3rkyfrN905ou
Vv616VKmfMFI9nxcn7YMC50gNBi3pXUAsLyWz8QIAgSdvXr3VWLGogrJtBfxVM4c
Y4UqfqwvW1J+tGIMbeYF3ZsfWKcPMD/UQQDWrE2U3L7nj7jcGib5lnS5IyMu8164
UsjagNnmeMKV/GpNBMKg4NnWPiwTid8H+fXZ9S7frnRrkFWhb+yMPoigEQWGLDME
UVxhvohLeB+652jN2S26a8P0QUazbkoeG/X1nJxf1j+Pa9ng/YwDpo/t1cDTOjhL
w0a03I6HUMMCgDFxYWvWGafAB/HNBbz637qUuYpOSAzK+ttOfktygOrnqKlOZVeD
TIRnzRc9hoPQGaFaFKIWaqsCY3MVSpeTvVJYiZecZX3mPzD6VoEhk0I+a6+NWE92
JYJINGJNmWwyIO+gB3uZY0hhLhIN21AE40TZpqfGOstzLUsol6QDRWX4tjdb0X4Q
50CIe6VpANLanaMjtz3O050yUJx1DKobOyQNCCB2UcGkPihA9np0fMV8nObODPCQ
FIFycfOOzFsTN7HbsLLSHiJ6DAYTeuddNxj5ING5ey6Be9Y8RtWi6knUeKGFo61M
APQYGB1c2aA3dp2XPpSQlMqQiJU4+41S+blUIWI+2+lfzDdARBfJDE0IzqTS76JK
dmdy4+d2U38vqFAGijDfiDu6x8m9TrXB9S3ib0r3ob8FDPB7wl+Q3+wpUsRqDj7j
+hYLtN0A2ElcjpukCe6xgBU79UnZcAtwsAksEOEPTbAQDoAUYupOl6l8hF9eL1eH
X+HybTgnBFMVujvE9xsJsNCCrfGOCEkMMLt4Hsgt803mqJJaM1tKtJNtysEcBx54
TfKyzJCQdrMIYXNeIBggDqOq9Tu4ohjgr2CQxEQewJKzLLrtzlLl9MbofECUqioH
3O/pAQINUp61XJPpeOKX452z7/nFLhfFzPOltKNln7mQITi6rjkNKkPPgbI9FgL/
xz8jcmxuXMwSmfUhZ7dIcZsLemgX7su4ut1FSD8xFiUY17a38sFOR3G6hlAcbDiA
rCwo4hYMTZ+TMb2WuiH3yWBodRyYIx3WJ5a6NoCSvUxvmADtPkNP7bvlEBMks8yu
v1ROMk407kF/+WXbyMpDUWuDxOeH997Fyk2YOU3k60kxpU4nDKdRo8TKkdK1ZTM2
L9tP/gMONF6PoYJ/UclfGwLW61EnBgrA4C+kXFlXsuJP8lbBHzS5twBPgOcJxOLl
RH5z9tkv9beYP2NmxDYzROorhKgbNqEfjWlEk5KSm8R3uLUUZJbYsX7xGYVdqo8z
rPfgPkxqA0ar+SGcZiEXPQv8TEqbb5w60Gdiy8tMW3TN4oFn7eOOMPw0FoINOl+h
+ucsm8DdmjcBFwZHUeA3yEcEOSLTv/QBdzq8jLjbMAxrlkjrhfOmhtWe6Gi3gDK5
XCzbFued7f1NVQdE9ZYS+B32TndZ/6NOM7TGjzkqwG32x4CLfFy2BM50dV5uHW1D
t7bRaee3erlLvkePPhnR65Ji2VwN6PFsiQxXtD7lXwSEWuNEJD2eaZ3T0wXsspyK
Kq15lQiUt9gPXXJSIBGY+JI3pdnZmpbIQD3MeW/dXHSy9ecZ97TFrYyqF+r4mIn1
pEsoIruWqV91bGRLCdndR/kQxSw+e/wgRu9sUd7VxGBTL8LUahmgFciv/jsanwLb
1vOt+FwZAjZAANKXjbXMfLzlo95BJCq562Vp34So+vfSp4apl2L8bdfCFW/RrCeM
ASWuJy0tJkoLcU+7J855xfb1d895PrU0So8a2vxnQEuhaZav9s5rbx4oP8wbPnhc
Y+Hl+vqWBG8Ef7Bj0zQoZO1PQnbgvbobIEatJtwrFDcsveFV1F/bigwjVS/89+iS
KAtee/oRMVqTD7uhAYuGX5P8hZkrNtbDLyocGZ8kTGWEhDVM57hb0Kq7eUgZ57Mn
YxmJ9WdYiM/9R8hDyjuMg6c3jc01c26lnjcqJDFUxcVa5oIz2cbOV2JN3olScXuY
WvhYWYZ7J0fyyX/OoiU6nHSm22JfK4e8/zV09ZMELRHk3xI73FJbXiMKBT814gwY
/YVWrvFSeidW4rS2EDjixeqFPQXc8FRmXPbjv6qdLWtuRyZ3LQ8Mipy0GS0C2oRo
MHNXZizU0Mpgkqjcw3iYEGrvGONqDM8BKSZVM3B2365pdNtUhswnGlgeDRUpf/1b
rXnIpXNChHwq/DG9AopQ9m1CWnAFzcKvjVtEHTscBogvi580FgVu3aD53JkHRvJK
aspQHTIfPhXZG3zUO2EUdZK8N/fSllLGp7Z0/FEaD5x1KWT4/1Mr+Qa5lQ200woN
YP2qeUtBcUpign3pnf9nbAwD+hsQPEL83bfoKEjOXhRGGYQliHfKvsVR29O9LS/I
MdnGT3nR5IByojRZ1zMbN3hKPPqii1He3ogW9We+jcqijksyPjkMeltT3x+7Cnt/
VCldmF+kBurQxNNlCtvk35cLvyieJ62PVFaYG5O8y4h1K7YFG6DilIvJpVHDlC/W
p1D9adoqrLBg3eD+iJ6SaZt6rtXOO/TIJV764h7rjIuFVUpdjRmNS4uUKHZzYiDw
lUN2HPNEMXOrm2+682tGFQ4oCY3jp1iSgEpv/znWPxIfj53vZYMJQD45h8vewRYY
jLLLlhWvdqhBWcwqdyP0HSbF3vIR+9+KI6+MNWKuU0+h2l4Z6JdHpA0IpgGPdU6L
49LXjGyMwPPHNr9B6yhGfJBol6hnFcQxRlOJ4+fjCviJ43tmiTgyTNMoMk010Zf3
j2prWa3G6nKxZzAYPmNhW/MEVGhKv1Va18qSyA7F9wHOFMXwEIRoU/0a8q5MYDvF
GErHE9JTEn/2eIK9vdc1EzbQ3PSXm8RWNOWabQU503iTr0HhYYgT4EYczlXj1dh5
hTPwN5KZOBK4RnnVMEJKXgOeQIU6Xi8306XiiJVUJQ+NtXglhCgOQm5q8Ry0BXr8
UH++outr0KoF9XR131ugGXtXJPnJC87VnaS3vwSZarYAKt5zl4lfUMykKv1yix/C
YlYfJEUOrrcDIW+ojPIN/GEyVMY1XQP2hy+q7qUJ/+znb1O8UY532hrqzozHUjVO
MWM1KgTjPBO9bboNms2L3yhdj0m5g/qExeGg3UDzg+Rf5qVffpbIzqzvyiDPVwBE
qRGLIJqcy9LH7kGeN1Sd+EnLDDpBRVX+w4ze+ggxY+zKab9UkzYMclgPPjEVjVGa
9nc3EmSacaa1gq1fDKd6wz237zjxIrnmfKs0U07z6dt08Tjl420mn3e/TZ2bKOqo
gIgQtzumLSDgbJPqxe1ZCLw/gacx25jF2hM8NTU2WtT42ti+9I/nAu3suokp7kIZ
kPvIB43R4owaS4DnkBbd6nHHh/qmfcO76TNIJSrHp1sjqGnlaoA1UJPxW5AbCgEC
EpXSmb7U7+sBNOKAGNGH+VQTJSYrBMou21M2yfoOS6Rn/b/nxKD/eb8Pt1avwaJq
QEvrJNCvT5622nIABdLolDNgiH5xohQMsRfBdkZltALnusJ5Y+7KiYQNgTnN9vW8
v62Sz6Zw8XHAa00eHNVKFO8fL52j+/rlfSXS3ApIYp+mon+NmBK02FlNhTtmAcfK
FIspMW3w4KGyLA4twc9+fJQebUQedRAywrqQ6sWtXNj10aVPOR7z523XcIZf3sFM
wdchu4HaM9eWDAioCQ1vYR51SawE74cElgkzVvWweqTYh3HPCMvkSsU714LwQUB2
J0R0aoWyssSlX4Q0skpQywweApW39hrTBDSz35hDcPXOO03Nj2wIUZDyr0v9lpKK
c3HqNdhM+wYnYOvZW7lxCogIip08Nse4CZr7hGvRhQOrc0m+KsrGkWVzlGyz05t8
iu2oHdvviWatgCA8Lj270s7AFgXu+UARzaVPmeEJljwSFHbYiPvgGxEA2d6Mn0wC
JZCydYgUOfHPj+257cn+tjZrzUfCWPdiFynF8e4StULhKoPtHvggJXChA/QJtmXv
AQxNnV5kMnA7wH0KMIfQbOj2Bg48kgw411/D1vL1QXYQCbDG6SJ4TR79mkRazSP7
pKp/LsqOrZppobZhMNSNn/ZmriAI6yAGio6rIIsh+Ru8WkNVTv/NJVxIU2ez8+7y
K5fAK4cnjkhZSpAj8ntMW/ERsCjd1d/HcRknjUkDyNRagtM/rutNmuHIpGEA5JpO
mB3+DtSZJEeMD9W423Pmh32T9sL00UAgo5QRNqNyQWzXl7ijypi9rZkHFF+nBzQY
hBJtkFbbGHuGPlz3XhJgsVxsOrgLC0VSPksoQEXJCF2AjgyvcliSk29RI7v1hZA5
BJkDQGg+vhde3x46oerqEp9NBMLfjBIXPxIVunqZh6Zp7mCJo4P9dnS8ivQufdmn
sqMmt+FcTlwaH8FcT5+UNMl4jZAk5Cob0bpMORO3n1i+qF0lP1MLImEB2FhGzeYc
Us8koTM2zObM+93yeR/Ux4twed1WlKBIrTpRxYlJMaWo00VjAAF+FNEGj1QJaVGr
jHlEI2/B5k54UTGZfRj4gUs2D0zVhFTzPoWc3XtlJmjSP8oYoAaL0gyawZAbog6X
x0rkzpRc/Gijbe2AUIS0DiRJL9jt/imMC1PwtzSZt2KBVpgHRNyM8tb3AsvW5nYx
pEXSRkDhhA3zoh6Ac7Oi1BTkGyl0nddvQ5de+PjrR5qlaqXplKdjkFTBb0HJg83h
PAQPUXfRLfixXyGR5a9aEq/FnQvkUZLaFajR1l6I1PNGKj0A98ENhQ1ISqDcwrcU
91/1Nd2l0+gJigLJ2CH0I90mdjjuq+my59cxd/jowR/vwcWB/ktRvyytsAIZGAdj
YJ4zdIfUFz0akUDFGN4F80lJvYKrsbf7ZIohCxd0jHkvxOd1+1jhEbKWJx7ulrnT
h8C+iEPYr/Y/nfWETm9TqTpF7EPhiO1kUNawmlOp2+2t+db4dhJBNb8gnAQqH0CA
JGqiu0DzKmsp2IFBdGFIqVxV6YoAVNjR5sFu7ja8JGWfy4qUyciluvyzLNPQLmL4
v/ogThUyVofh+lHiFfqVtCEMgGLKKgfcUn7qya6XQ7nn9LUZ6Hcop2VXUEkS0nD9
Obi1GaU2a01X9ff4QLaSWn5ydESDqZeFPctUQGl71acHei3wqT1SF2Nc/IVQ/5om
pfH10jSqfyMwJBdOPFERWrO8g4/b3nOn0VJAQ3e5R+2mELndSgMe+C6qtaq0KLLz
fyXfbqd40T6qWqZq8P1Bln3LnkyM64lHtRkAjAF2pZgrOwBebpsTm0JX+Q5l/H2C
0hSzTPWJcSd8UWpJGMbAuee3Q5J/RsixhZ/QgKTcYgtR4TaSJC71hpoQRasaeO5N
cp4OotYni5eNUN3JcvHBrXqExtUHUrxJrKno07njg4aah10+FTqeSHNCn+nF6r8b
8jcSaCxnL1DluADuf0qQEQcb2Q3+klpZENXXr4fA0OtbwUMnja9QBn7LPODP+tJg
L5IOSCKLx2fXI394plZkAfkG12dD828mxkO9++obP7sSaFnhFwDbcp+LXYTiNaLH
MXuovlYck1jMibAZpA+3DnN6wMkygIDNzQncSU1ibcIKGSK1GMQSDOl1A07U1d4l
zM4Nz93vJrr++yQjSITftLHCQkmqJLZcVIyraAlCKhmZxxFYER+mtaygL4T92qgJ
XTDGN3hMx59d10jiu359tBiAHvinZqAADMvzUyHvC6nTP/bzMV4KwgfDFPAatNVT
MZaf5vyMLk4206TqjKSiTeE88PL8Ufli+l9/4OGs82UWhgp4rdFXqb9SYphoxi+k
cBvGYNGD259srZdEIZa0xrVcP4SpscHrDD4F+JRcmx2NFuRT91b3Ev8lZuiH/499
T3LPsqy2Ln5ayacJsNvudRQ087klenP5gTVuPjQfoz7Jwmoiar8wt3n2FqrnDqdz
K2sRYorJR/WUlbA5vl25i5ZBpfT0r4GDkPC43CUttUkFZud0OJA2a/dcTcLVYASM
StfCfBMC4IeMO16SRHHk6pUjopgW/PFJ8wH8Y5UurEw974peC1BT2ugD2snAo2Bk
SwiopRkuNOEaqBDUBkiS/PFOH/SJFTXBch7AaAv3z/2tz+2Q+fndJfpw4aj4AiKD
c0ReJ49jymwqLlUKopH73drHaGKZC7qiKTNvpaEnpmLis+U93ds5qNi0jDJL3T8b
jmJS5TCV2mnsKl3Bc1eMq7ueBla0X6Ku2YR3+Q/vVdvBOMkEWIkW6iZL7p808Dt9
VtYp8of/WJ1tNJrQXWsPj5BUmX6pdSGG/+JSw+2VmyrfHd82Ysm0pW2W9o9Y0IJQ
vdUqxFs8TyqStmtqYli3S3bGkP83doQGJAea0Jq2ZFhm3cVWBODxC43mVNtNUWSe
HmdD2HPfcZjGIwbx4UHk/xWGHY/BukfIYX7hKxbOgvKYmAKH8JP9oNqAZT0wpKn7
Kw+OT6bADESZ4dgorqnwJPN4C+EEZmbjdodNTI5DGEwEpOSgURXa/wO8UVhPUmw1
IUmhbJlaDfxt5JZ3KShlzpts/AKVE29SbKtx5wOU3lTZNVTqMLcaGE8b86kQtIDg
h94DbLHbVylKJdi1N5lIsZBErLNqvk6EKzGNITuWfCZ2bU3LtEPS0utp4ahM3aIB
B5XDWAZJjyJvilYp6+6D8eNrrMPW++3v71kwQnmHFTR1qp3lzQ3tAwjrWTEVWYs2
8LlBmBUGhr0XDHvKXGk89WN3ETJpe1AIIBGyuLCvOXObR1Eva1KbZyzaCT0g8Zqh
K7i9RgLqNO48RsUjmZbW7eYvMkKmWPQDwg/MfnVb57Rf7stx1XAVzYqNSBCTTr5O
+9shdA9INHDtMTqm+gkBd338/WawGe6jBdfezx1uXls972OOnwpNGU2/E6xq6FtD
7tIteCY3mrsJSobU9n5WJA2z0lYab2lX5wgNlz0BMgVe/zJZbAEOuGv/CweL+n06
VqcSkuGx8CIJ+L5IzlqtlMTfX+58UyxDTWV59ICt1t9C/UOp/GLyGFZmdgNlI7rD
aI9yEmxwoBz4C58vNvOG9pui8tkOHHsQbal9GoJGb14gXAIMFcjQ/kC0Mme5kXe8
dnwi1LccdU4oBj0eNmu3fQPdqJBRRmZXnjqYjtLtFiq4QBHpZTuED5CRmv2FJwOr
JJYQRFg8dO4/W7REIsCDt2WpAXQ9dwWtrDemTbENxF5Ja9obR17cTCsekajVHCtS
gMbxajLpt002aQf9PgDGW4Z1uDWpEQE/J+HEPk02+q2f4MUoKFrPAjcyJGyLRToQ
iXJuFK8TkTdQgcjybrKyzCYl88mb5YZ+LIqRfo+aG6J+SkiSAaLbaVgMeREPxjlX
lRKI0FygaBkpozHVXOpcP16YpXy5In+MbWfTbMTr5vpQPITzFN9xeNFWHnrX8Z6D
I+WFW1TpX4DLsU6VRC0xSCdXNEA5Oqs89xEzc18FwZqjFYIq6RXu8VH0JbfPpPIm
zA4a9skf5Q3Q5Yhyxf4zM64dHgC5yoLYaf8oCcTV8HKI7iO/bJgniL9L22ZLD+Yt
rfgIWTW+hSfokrvwd2bq7K54hn6lWfmveJ204K5GNT42QyRQ5C/Doghwz+V9i2SB
GUE6nbSqvVHbb2QxhtCO2arxTapCG19FM7BxxfFby697Cicpm1aem9PWZ7egj3M4
oSJeTaZ7yvMVLvARM9ecQ5bA9FGN0X/2JdraflCiXwtFO9Q2rf/LYoiKZ8wmAG50
YPR/Uo7AxvwZs9YKdgVSYhGDi4zqWkkJoGBnxqIa74iXp7WqoSbwngySkYBX/EYY
Ns+chCGD11VsX6rEmb8VSOm9t9MofXq+24BJO4AKpJI+IWBWoHF1Xo5Gzm0uCMe3
tKqqRovxVzbLew3eRZ9ZvkkbehWgFRADnPN/p9BGOiPHCz1NOin8dPHS1wi1MHXV
n7HrcZrsIUy3m2rAVOa2f5M2hZ9d4qL0Hxy6cir39gFArG9jJvMoqkmupxdnpm3w
xsbp56WpzM8W69LR/lSNm1Od8oS+5kku8tUyPvwPiXgeSQlC2eYWDUGIj8LkzPxe
5ufqCgXeTa9DvZGOSxbaYUwMsnM76V2gPmxhlwhq5AreSGOjN4ihg4rfnKzZx8NO
0SEE0RCFEZw1EpSy2VDSgR9o4o1TsIL+HfpyxXGgO3GpmDiD9rHwF+p6GFZ/zLJj
4Nv+WzF5HefnguSZL0qWVk7jYlad+0DiXWu+LYAbGSWFjj+CBbT6dh6x478dvcYr
9KH+ZJhKCOsmm6+I5S0lBI+eGvAnzw/kPKkcEPZstFSBqApC6C4DpDeJ6BJ/XeL0
OIHzGpXbKpqcS7CnYG0TY3VdoftwcNoECw4qO+6ZlIk706vuxj6fsPwwZl1PnWlg
v7Lrd1lAxlNa43hm98p5EZqqliS86oYR25Dy9qGzIa7PDDjND3DTl3oxAZ/pN/jN
ufKJs8p5crizx6E/NvX15vO8zbM/sqjfbRRgyPyRQuE/89jmitGdMdnv0O8rpPeH
YWy9U6Bb2kPpdwt63yvbwGPBBE1vs2z0IkgdCoK9g1tbhHd7EAugfC039eCVmK3o
+kKxY7gB6gxVTXY4PBNUOp/RJiIknLqBzPgu7Th/wS45kFRc9VmtpYQry12g/psA
EqeWgJ3zh/+4rPsu679pAMgwyVPE8blKAcEBIFfxrHxWQhV10fxUJrY8L8SbP/c5
rmTrGN6FAsB8S7Ci52L2OuKxVz7l5rPkZx0uWZMoXIf9Es38uiJtkiABZiM8+yZx
HGg/aA+UVIqpfyGdoSzAs+nmkE/MiUOmdaz4DR4JngbHXfR0yrRP72KiUGGkGe2O
kgTOVFJZuANBl47GWng/7ygsOzEXoGFU0cmHf347+uFD/mMYkxEv2e8GsSXRiJ1m
FXFwmy5gbfnccs8sOoJdFfyd0/VPi9GgG8DPhSPhMbWcazoWs7nUX+LZ+t0awDBI
J6/jfxdg1hXFtyHil1c8fGcLMh2txQZtZukviljuSk0c6yX+GIbc5rIGo+SaCvD7
NmtNVnwSIDk4F7lndj8JzF81mo6nwFuHl/EQWIKIh4V/D9RAIAyYMHx5q4Z8LlTt
Y6pv7AyQ0H6thEMSRYmDatCvdCoeUd4rhHQhlJFJOgK9bJpDRGaq/pIBRR663LvF
K9uKyIacKt4rTGmlnjVmSSUxwXMhA0koxlGnml4yxl7cE7KJJnAPtG6AdVpfebcg
q0qv5G1pwDstVgjGvZ420pmbhjKIMKLqSDO08mrn3BiuMFwxeHdBuwCBtPYjGf4m
dEAWTeYYf3andzIM1/bvi780y7TP6WMET8XlC5VQCCm7q/CEnOmLLzuhsOIXiuA5
kEswtyPeBeQDgBje6KdzbSCCdE4SJCJTsr/zzooHa0H4YF8G2O5fytFcPsrLI1wW
G8vZHTVLzKQE7z+1Agbdeh6pKCOkKa2A/YuNM/WWJ/h5E5bXQtWQQd/UUSW+jEMV
IxCNxTli9207nxCZQ9TLhY07A3qNEHFVKWEB/wCH8c34ma8ZQl9gMk7gqgr2471a
UcHf2Wit36vdWqH3YFut2GPQsbJWOPaaPaT1HplFOPrFXktVMqUR+i4wm3fIIKEy
+0WykY4X72S64hhPfbxrhqlfpjp9I8HoGegVMlSuNJptKS2SSHmA9d9UgxIUJI+G
WpscwSZMCNG3QSIvRdHFoFr2TLc5HRcDmDotUKkSZMIN2aVBMui89vGXMcLBD9ik
BkEYkCfdmGlXmA5OvKRVefcc1trghXRaXQx78u2gAlb1lqFT7YY7VIwzzuexKD9i
EAjIz68uT4a5/uM9+IYOVREooVu5zcvZwjrPR1k5YDHIJaFams4zSh3wRahJ+jMj
rwer7IKPYpeE+dB1h2cIadX7TYwZnn9uQAwI7mrGK++fLeJqBk0xcwojOnkjdBwr
XfgyHENaMdX5PdjAju+tk0EkVLGfrX/uv0FNSkOfQXqWmqj+OeeqkxtLsVQHX7Hz
ed2ogI1AXLz9xxKD8q5P0ouLp8iOJ6WX/rj8yo4CEOs6rvHGRYlYJNL7dpnlcRpa
hSWArS+b2EUi+QLhaIRf2vby/+bC+yNStSMHTNK7eYCMruBjVf3J5ptVUPQmfPJT
F4n/3kXriFtMPpqsC4+UeHk04HsiIdbg6c6eUJ9F64+HtPszpdQokWCoDgSQkOy5
+R5mia6N7tbYCoMJIih9puGq8p3dfDwxBt1uxuWi+OHoSagN714UH6O7gK3kE0ys
gYXhkA1t2hGyWQVYkcVu5HsiRe8jQBh8JpIVn0uLVtx4rim0pijKadLzvH7L+cgQ
Xc3dvN4UWYj0hgkB6vfAcZW/3uyWVLZh6hX+SZzA73HsjBLEA1Au4EMmkctyjNKn
H8/uBFd24M8JWfFy/zg6ZsCMCwOUJOW+fcplgJQzfwfRkCJUKU2ENSpG4GtPMPee
vGFoWcalzK3Yz65fyY6RX0k3qXuLIQfmTsdZYil8+uIBMpPZOwj5aS6Gy0iJOQEc
CLdmzaXjam26D7bDvSlcjxzMUoX5/TUPFAoT8rujYf4gPpvGXjFq9KYqEla7vzHW
J2mQo2EDtXq0eD6rGnMNYnxlqee8/BTEhMJuORhVAYRIwW7SdtqzSCD/qWtjbz/3
OmC7H73QlzmVgCBFeGEH51Wd9ZH51MrXNYuLmukrCy9Tjav28FchrKzmz2sK3GBg
f/Gv5wAwOpLUoB0JoTgS0NVVJ65Wh12gDJSm4wmYHeiPPNG9o1ZwI/IqetUjfpwK
X6GWEgn9FzmHi60t/PatChdPsUxHnkCLBYBHV7LZZvfZvmrWuJRfZ7byac72dGNJ
fM7JQUaFkQ3SnDIR+fyYbyjUnSf9NqKhrkVZWf1e+nrSYmclFdlRsPTDjzWrKZVo
RHDsVo5FLE4HfONoSpVOQI0Br5iIy6am/FF2GJP28Z1Vv0OB+eJl89tjmUj/RRL0
XX7c4NY8M6hjGngoS8XHsg/v9TcYzKvFsvAsuEY+ADMecvkoSUkyVlfTTfe9EVSo
oQhgd7MHCYWRuoufakzG/bS5YR9Z1hSZ0hzVPHm8vMxgh81vHRHpWD3HE1Ipx3jg
IkAfL3cO+aAFTQanuakFcOR0eMH90b/PM0Wxf7fWE3LmUwWhdnH6MZ1VCus+0Fan
7zp4XSXC89btoF5P4nExXdN2i2+tanrtDRyvV/kFE9Dg3PZEWbWUQAt9psYDo6wq
8/3xvn2bQ0TwNFTbqXIKPe2RXYx5BhOWFsZ+WNrWxJDjYQJWMB2bz/di2YDL2LLD
ll+ZAza8KbQRIMri2liuidhCDBMLcClxmR1jK9lFvkV9wJedcBJvSb8yezJEc42R
iW1gZXxhq37c3GquTgkjzDB2cEODhLhA+c1TIt9mepoegF+OmUjUP0vrLbHr0Qaa
GMVbhWzulsJlrPRLW4jHNvNikY+aoc+fzXX99IKymAtTKVD2Bjd29+eJQ216b9Vz
fb+22F1306OKDgZzeL/swyFutwaXaIlLPS1ZXiYeI88cIA6sqW30EWDEfVnKkec0
eDzyAC6uWT0kl5jjxUVp905OWUb9Pu5E5wSxLJs4D3soStqhp1bafSwUYgMOqlD1
sZ87tYWUYroKWTdaSnZ3YMeJg6T4RiiZDbXIsmdtP3p3opr9ftrQO5cJWL4WvtWm
qV4oP12oUd3TEHftL9alNj+hdZesjDWMvmxpH6ce79sUcyLhKaMeN13H+NF8YFHK
JNcUY5rBSPpbzrLWUwNkL/+tRJhlEAmi9hxiaR5AMeJKJt9VGx2SLEDzFwHXXrXf
EfpBW+eLSLCcK7tSZNTjm9YpRQUcjf3esbh64zbARYJiNZ2nAm5y4Nrfr4vHFAnd
7BATZQtLxLMw0FzTOD0qW3FD9ZMR78KYx64xcB8vcmfYoBOxDFFrch0B6qWcGwAY
1FP9le6qckTWvuQWEv67eIQsrmsxruIPV5sxa4LP5+aCi9o8PI4VnN2gL2mj8Fz+
Xg9bnCWb66M6lC0+zoEiEhku1dZFEVsewAkpqPLud90j8q68WVFbYhP6OcF1IMfS
tfHqY8X81NHmEPYmE1RIX7oQylR25kuMH2k5ox1lDuY4/FIiO39nLm7DMCgSd7Bj
a7C6jpqE1D5KA18U6ao9ifCy3M/WSZ+BWSKnhaM2F4cxgTYSl/codwOGwihEL4ZJ
/k1PSVuffdKohkzJbTQ3swyImS1TkTLFhARlqHUTR+o6EspI/pxNs8uHpyfpf11b
OzWhGITCz1UW5RYwDol+Dz0BU9LtqXNXsQ06zrL1+81HHxeWhD5hebN/paN78957
NR5ave44KQcOqJW8p8JkygWtGFJBmBTz3TbTEwsLdiNGWrSwsUTwpfAHiO1ArvFd
LuQTy+7rXWr1MgDjujOQROWXxV0pYWezMEn7t0+/yDGsNYmLssDr2zS+uVHYOA9s
k+8t6IJWiV1qqD0pLQdEk7z/iJMGcLwACehDYXFob+ETUutm48HzESu8VEcf+M/y
tUOPyjBY3fqddyrbgdrIISUPAJzTqVmUAZ6uUZBYg2KMGAELjrB7bnOanxI/w4DY
8GEx1NC5MuKl9jElEyRfsRc14lqaLGfiHq26OmIhlEu73QWi+BnYIV4YKnfUrZto
swSqEA6BjRB+Z99JK3rznkuD/vBRGKnzwp1SZzqF1y/YjnGg4l3HHSlqADvXhN29
CZazdWwZHpxGcn/V/Kcj6uqKY9D/vI7DkPqoreSgY456wGMUY9I0MuHuXVJMHEVH
6A8PzKSEXTjE9Fc0nwPP3Y2xA5gloJS6x8grIBKASreX5FbVafQKUiAQhFCAm5OT
5yH62HAM0E5EGHVM/6i4e/lG6OADB6bn3MT8LkDmABC6eDFrHlbAWx3q0X1LT7Cy
emwbUkxYvkGWuBYUnPiw8K73+J5fSdO6JQbTThTDK0z4xjdca6GrN631dGdC30ri
5b04IRL3CTh4il03Ax2PnHMhdtkca5GYc2qKYb51AeIXLsDRVh2GZvZDkVLkVJR5
SI1Mu1CWxx7cgP+dryyxHvhSUyNkvpYxcpz52RfR7pZmYzb5+SCL9pcJGmyrKL90
wc0nBMWNsP2+mZo+tC8Urp+MHa6SlyBFv6Zb5gKO6hhDUZZXvhEyP6PeyOTDWylX
wjFtRR3sW3o0nWOwYSZ1tsfud/f6Ug/1hYZPqqaY04zu5I81oOFtJGJwQgJhdoQM
4F1QncdM/rQI2ErBW+9Aqvk1R7GMoOCE6eM03IFX1jIW0U02DYH6pTjLO0e+KmXS
B3ARvFNeQfq8Z7ml6E6BY/LKATN5uyeexCV6tCkmM2oEgSaWSukPo1KymlN88bQ3
ICgBHY1cUXzpQC+DDm9ZNGHcVAGnIEiL7EIgvtC4CpXh4ScYHaf7q6z7jYOLoSpo
Tcr25aulKTGftNHBNugTnee7eUwJqG8Ae6Ppo8fMGN0+GMhlJqJ5oC4smuWfE5rz
9D3f05KZCG0SxIPTiQ5Urx9Nly9ibv8Rd4ISeAtq/MlePltJrHmswAHLVdysSU/f
bKrfdfbki4PsijwfFDb1BQnbi5/FJsZe93iM0mp+JL1WTRGRInKOr0ekr7zK/5y7
xPD6ZBQApkIst51XsqrSTGNd3ekGAQOIlMZWStlmXWq+LaXLhH82e01DCM6B87hz
7ykdqhdes7LR/UAc8a0Dtp6/PWLm6w+AlrH8ODKOd9jN/I9eB5QIDF1jayjSekM+
u7syNg+GJSeAyXILAW/+iEtrWgR43PID8sWNS5Mo/cg1HBDgedleAGbb03177SAs
AlWfyRgGZ4Pilnxl9GwI8iigPpXPSklK/Z2hwNyCqaWI/lS/U39bg7pHvNMwOoFH
rm5BjlCofxxkO2pkvdDmvHOF/Y8aJvQ4QIXZGcQu17NlzS3f3ue9lT5ag8MdY1Wv
SLJW/Gr5zDbWCT89LUzYtxZTp1W/RyNBXit7mYikFQhg36rI0Bkp580v/ujMoHPv
48ikDADk7oOVC4qllHh5VccFPkdmCEJTSPBbitGytjpDHtLIZ91WC1xs9JclNutT
RRF/4KMiA5LFtmLS978B4UMToQxhjoTdv0Z2O9SYfSGRMSd4xc1PIUusSckBKT0D
/zSJPPnbbemgzpQriBsR3Jse8kPHLCqjDlvSHwjesRzFvBXmiQEFMQ7DZ7HuZ5oU
H7so2y22CvqjAr/2HwQbsG5KZ4HXufZXzAEZUlCVMyMbrE5YRSpIA7Y3+QHfTfPT
FPtqvsyGNZrgoligLOfrbpDP4MT9oOtFuPXNhb6ifHvhoZLmudEqc8T0DhBTa6zk
T8jgToET1eGJbMlekapJr9YVORoxMAtIZ/gAqOCZ/Gwm8ZOooW/v+8hWmq4Q4TWl
9EOSKk3wGqeaAH7eNsbTYG1fSm0ImoQkvl1f0CpNYNZyG1/kZZkgCFEUn0kGAXaK
GzMe2YOAt3+h99WX3SznBRylnZlwtaCCQRSeKOaUYE9+iDiTaD8rLiwvsjFbcwzt
8ALco9oC5qen/tQiAqtkvXOH2LCY242p8CKJFBiMuzit+Krax6UBYyJz7l3ozNvJ
9gpl05nZVcPE5BOFnnPFgVwLBEer9Adx8rYVjXqsG8/qOQwCyjTxAd6rMWSl/ZnO
SMZ0UQU7TI2P8zZ0DyXBhCmdb+C8zfMH+DQYqVNIrR8Tf+DospIAWm27cig1W+qb
wUHLWpq/e7et+EC0sSYhFhg8SNuPXJmnWqqzIl3N1PitUPMlndAq2M6SNacRzpFo
DIV3Hslv25k1pvfg6VL2R1Fg2kW9diL7z5wLf0+X+Z7yiy3LQYuiexUeKnyCLoYo
ghNDzNESiLYK6GomxB8UZQsda29pbWt/27cpB/yW/ND5ZGPIUJzSiN6iwHY/D2+i
jyGfTBsjJGA1824D5h7DTDT0W6VRWnGgaahuJTahmcLI6G3yptVztIx1Ql08+D1P
xJl+K1vhqlS+FWj0zNIN6s3hDI6lFWk8WJu97Atqhwo512QySOLSX0UdiKIuMhaK
64iOH8R+R/tlV4bnJxM5kWfELVL+O+L+XfXDwisKUDKpGKoRqodxsRPTuka08Ba/
4iTOrF3aSFZlAsY/lXg1zm0JPzv6d7gAk+1DqMiQizOsXsCzHAtf8cg1PFn06Tzn
AkBCLMEYXTtlDNF24uJ3vWesPFOfSSn1mcZDgwszKssHMVWzqj5nMk0ISCDNcKRy
d9vL5GM2aeZyKiqwVlPKGxL4kfm4Kl+ULlNDD+cZb7p8xEEPC6mcw1VGBVqJd225
Joiv2bRv77keiO7nCmDVdQVYvnqbWEp3IGmVORatYZhAd12Uevza+RHIZUdKk5oY
T8X9AlQ6cm0Ojhj7Qmrvubl4u5Nubvr13SxTvC3ecXGZtKgIy9jQlBVez41BGfex
2Qkclqib4DjNGc15JPM6BA6IOCqrm1yOvFK9wLhYWDDpQpMxpqqhp7/ytnVjkiWf
4feCVgAV0OLtesv1X0lFXM4rGCusivrZjK2L8hiR0h/F97TaMtIYAHLF8c4qM+ah
6TXeDKXc0d2WtYjw2tfrmQPhBS4+V6EQtjS6bK3OAK2UvLbanTztKWaO/ruAV7N7
f5cqhQBn3BhHHqfooaAS25Cy/zkwXUBPPp4yS88gov1R3Ec2wrK3ioY8y4qs3jAN
qRSOx7fOxFL0pfQDTPrLDWmwDjBiFK9w2bRqWNV0W+SSkkWs1KI8vdQ3Ufc0k+IR
EANG25QUFcf5yXVha+w7kKJQW7bkwRVhYgdAfAIb7517y/KuPwym5pypLo81WJOR
Y+t9RzqCdE4xb3j8my2Jb1xoLJ9DTupfq8lsLk3I3R5j53N7GfTvajIb3Tr3Tf/I
3sLM8iFYC6tsnQNJuSvno9evOpK/EUpJbliBpu7We4+bYWXi+LlDRhDGAYh9zcI3
BrVdpInnrsSZiX3vroHcGaNj74BgQ1uCG4Kt2wTdsq7C7YMnAfO9zoIcMWwdd6nP
F/7Zisbbky0dSk46S/13YURsNqlclaZBTGwlxG4un+qGE4jsTOxlPq3LwO07sRUy
bed07q3tupLoKZnSTjz39LAi0qAIDZQUcAiryrf3/QUbtVIywq8jV+ivBZZNA+Yf
ZZwS328zDx+NzVtj/97tCfyJxz/YCMBVxbrJmIGjnGTzJGMgGzAw788X6K0jJ3k8
lQqTTqsCCdc85oxJGtQsDUHrUcegVMkkUZbSr50DyOleNQLygMmFEJmAIYvsviPY
5xpcgpFVIRlZQZYNCBBr9d9/GSg+jAxdfMzpPrWXJd423b6oBCdnjXwsg+VbEeJw
v9mEanTc0xOx/Fq6PPMjcvwX9Ytiy2cggf8Eo/JBZASCTqED7qBwkx2ztAvK/VXG
M+8Zh1Yl+euGd/inIh4rrg8VbulsnZVQve4QB4Ka4NoY5zE8WfauOUxYZTxWoyoD
tIIBmNJh12o6K6qYB4rKvGOHGKjARYh6aVS8u59+OfWktj60+UJ8rIJxT9MfGbP3
lrGvlxwoP+a0U/ap8wulhE3PPOSPOn8q0tyuI9Jdceg54PLW6bv4+mk1z4g+rZLP
ZVDHEt1Nuu9yEZplJ/VQ5Xa/i6IKoYGWXF6O9x5s3tnJYBm77RzvT9y+BaLIgTw8
0dlsRHM0IDA+j3mVXIDFGgzCQ7dTg2A0MqHcrYp1XF8fgdMpMn40brdIqDOwaoPl
l+W6D+M/FwBWXRmDtW2QvhCZ1jnqP9z8Pocnq96D9eQPNR33MVcGk8xb5CpFFcVh
Fl0hpgDeDzul5a+zoN92zYSdDghHOdw0tBtUY1gY0L9xA9FF7KA8SOl4JpffiYaw
NAb1ALWsvc3pZk2J/0rYBFrIxwhb/4AncrtxcuTS6fDqaeR2E2wFRRUu1MB5/mhK
06h7glU5Azsaiczyo10dKlIQBPiDCiVbBH1E8EcBSzqxQ0/GjydqNMNDzFtzB30I
qwV5DIRE3Ely/21K2+MT3Af20jW0sf2WzFdVp1rblrpGsAQnitYAVBCcTw1++asn
IYF9h+7Q7sII1/ZE9uW1JZt78HClyI+ABmyhinakfL4E4I++k/rQGFRy3Y0a1fmZ
oApbHXjObo1VS7+mZwwFacBA1AZzs26C8Ey+ZyUoGxLQDIbVEcFoLfvrIC5nLzmX
yVz8QE9pl3PcVolOKynkF7MYEfVyE1yxBAlvpx+XIABcVi6nOZdGq2eUQyBD9RoJ
mBGhBLvYeYJRU5dtkprcz/Sk9ycsIuHX/sqjXrbunGVoR4J3Icbj25jfCM/qrqTJ
EuK7YLM8a+QMiJqwR5DDVXlVBjHwSB/FvL59a1WvvBWAVcAdgCIwXSuzDhfbnEd2
9+V7fiLcE8s1MDiBW/PMaLYOPXzQPUcsIYpr7UTVUSZU4jZXknEzG+W7MkVGRNm7
nG42H23WkAI4Ayq73B0s5TnBaqY4IoJG5Aw13QL9x4Oj0DMItPk3/THuZIW17f6p
KdXOq6zg6/kW59Lx1d14VNvT4tyFkRZzKIQVnssUR5AkOYHDgVhrETK8HQqLSceO
I59kYGB4Caqx81HUn6BBg+mUh/BLn8P/Fh2wp9+TTfGVBmGvGXqpSy069gvPNNT2
ZS4JvOHgVD/wMEcy8YzG8i8rLeg28i28JtzxYG+mpdtNB5k2wnxeeBwzsXS04xxC
C1S781WNOhUhEUnL7MPfe/YTMSzyKgCtSFKAwzbJJTvX/7FowAvG7STQYEPntiXP
pYMn9hM4UT3NL7fQeCf11lPQp9l6cxFmAxrafq6nlDGqbvkmYa2+MVJu/Uz3BTM4
M7XxAVn3nOyXsv9h35Vo/U0fY5EO56cWHJBmKqbMg/EGiC4RJrqU+xhBugsUktZx
mUfj1gN2H9KZa0Oqb+LvM992lcNiQg0g1WKvj+QQN1n82/+0E7aSFk5uWBl+I7Ps
EsRb93jPdoaIUB4muh2Kr2YkOeG0vZbMNpnVA9ynmsjGEZ995Q4Hu3xSd8IexHMk
Wn/GsaDecGTejdEfcXR9PpTfJUKCT+Y8fMj5Evm25JVh+QUbpwWpexjTfR6mqBD4
i5jzB8hkGXC89Ef0EwHlAlyCDFIDXIa8A+eeRdtuKjMpObs/JlLEnE7JKC168Hka
Eijs5t46cA9ZpMvM4zK5MBo6p6mHxE7U/Fa4Zj8Z8docmzWBD5Yn/IzqapmSRdaU
+2oSGNyLXk30tLfL9U7EqAmZzpGcC+wgqkFJRa2CEqG/snk/XdyC8ZaB2DREimtD
CTCBZnAwH4n1LhGsyQ+0MYu4OTmtqML8x6ZLLgZ5u8z25T3IykVEgjhoB6KwhYca
eLFnBdAepYMQjb3cxeyiYErc9daNLMFSjY1lRg+7uKmCHopSrAjbF5Us/IPoRguE
ljPRCXV5XQZrHRGNK5ycaI5HLICAhyW0pNgGV+YpdK2wNihDYYGKla+2JBAeCFsi
Xlk/xoOtX1WdwJL2hRRe2WT+DwmANXmfru/eJh8zeYp5+v+1lVz7yjW2lS+Cq5ew
trMUbmKQs1Jw2I7YRuHp7v10GGbuy7WCIBtpAKx1t/wvNift8zotX755P9IhICRr
wNsglZqRXX3NkYnxn+uwwYUuvVLGza93L5wR68aTxJi4xmbJpli2z/EPYTgOQTWq
nmumw7PqBkug5k6YAUxOeWwq6wC6F/YTPGgvYag7tOZQVb0RIWDyXmTAqzWu0E1A
VLC+GSuozIGN5MC6PXuKP4JoLMPRFDxJDcvlWOg+izi4QkSjAbrw3E+hFP3RxXCB
1//NB60aAyYN2Z/npLQHs05Bwwm/mp1dbCwS3i/dSl8Nu5a5BFa9xfmaohSfVqNW
QObhEUb2WEgvXw7S+eook0PVo1u9u1/31fjLXT1VfNN/qHJWF1AaBSYRPZG/4+kc
m7sYwxerrTLhPWrnFkQo3NXxwBzBUB/QnGu6T36UPs67KXntC0boEXPtTPdeCzVc
A8Mbfe3Wq1RXTGbCFNiiyBrMaZnBqi8fJlt7ta/5okkQRFIz+LwnV0B51E5vZGxj
BQVUbv7IrZ9N8d7G1rXGuFFaH7x30a4BziMmyUkZOVikDzA7i6hDnGsZzMB6N2UN
u8bbtCn1tY3M4HgjumCPrvvW5tBTwNVw722IzOUnppWY99GwL1GOMZycqbjNdlvG
1NtPRR30a/tl7LWiWNsEXK9bqchvvEbD9RkrsjTPKfwoukQnTMSkIexU6rWn8mYD
0afBtlfPIy/e371ZCUJ10HyI6ev4jNVxK3SVXp5M3P/VJ9tc7ISwRsoAexmeDqWj
ZQdLGzUvVgqWWcoVql2G6idtAQhlZyim+HHEOX+OdPbVa/eY522N3laHejtveYgi
LvFq1OwxTsierMnoBlNXgCf8vPG7lnGPpkwLCacd4xFszg61BQjCOlOZyFhIasYd
sjKyylFNGFCy29dHoMmAmGmdO5+3j7gRlboHiFp9ISpnA75WxM47ey5SJKzQIhfb
qDpgFkQ9pMnA1l/Frtq5aY0sGPzy7nBl06/nQ92bL+7W09GC6azTjoDF8qY+Np/P
WUMWuBGeimj+DHs6yHkcIhTuqbCxvDR4vlkEfVM4u6AylznSSItDwuXmbMIBaQXE
84VZcghNmn8cYgOmJ9trUb1IDUhotltZe82u6u/PIIrzX25qZd50ey/cLMZ6m2UJ
cN5KPjozf8wEf/fX0RDhNfTm+1fVCheNwb14yxfRWMRGJWcUEhdDfPeuS9sEOzf+
HCH36u/7sj2A2U158sJ1ioKczgfypBYij/0ZnEtsQf0KGsUDo+ybmg5Bszs8JKLW
HytLIkca1/DZYD6KHSZ0DI6hSTngwioTN3K387AntRSY49qsJQEyacAGPi9p80/q
DfyYzKpat3d0vCafpimYCMvKYILdfLguRTE7YIHvX7oxZdrHbSw3/ODbnRZh2Sa9
jZI7Edx5g+jgufJVKHXK1drCRBU4iMNf74q3jz66avm/ohvgWQky2SrwQmRA6o1g
f7PAnBPuv1cGo+k7V0k0KbkvVjawUELZW+mGhvMwF5s30iGDmP3+vQGXMnJlP30v
KlGhGNLGItTzh0RZCMs3scu2ps8OTVU3/0gmcKEYu2Zb6RPKPgCq5SELuF6O/Q9+
JnXFMTrzIEtmEMu22HoZE/VtloE6Rg943aawQH9ZAfdwna/50XiITrY7UHmS1H/K
tNRbBOO7IeQGo7lLuHnl0T/ET2RkhlwJoQeXG5ZDeNRTSNbrKZAAAq2atfRoKSUj
dMKs+Oh+DEGlrn4/ZN0/3AYZTPzFOLo/1LOzuLWoLPfPpSFX/NiEha0T2hn+N85N
UdBoC6u9xS9IL2eQ2fUJx4CRahxjIieoSgmrFSYPlfeteMm6DQpW+Ui6aQaUhn3/
4OwUOukbVilpHeSp+cyzO2wV9o2NbvQ/xbyWK687nRJnnqQ8R+EqFKFkpZ9jSnu+
RWNrVCYQfYw/Q7O4QF52q95GqTjGjoOVqsLE7KB+vK2zwrKLHbqwXHbfTHpm1l5+
i1JGq0lPN0vG4K6PYQLnTr5ObkSJT2RY1qEk5yUZFU9FYsKSic2LepPpCn558n09
CHd7PDQ2XoePixaGiSBzTukZom8O9WcQFGIA0IYns+T5GxHe4VVpj7sjpjNnupm0
UOz4T5zI9CsD4REgv6avu93hvFTgNHOBpNP90bUQ97Gxgy9bP/HuiIVTcWgc5cy6
A3Z/QcGFGZ/w0c4PfNnd4sqHrMkugVvZ3iwOrl1f9yj+HBCsDrCvuJwD76f8S78J
D9VMa3G4EeNkxzT7KgddF53eiPealNDT6qYFJ4NB54QmtUr/4Z8EyXIL18noWLhr
olHdVBDt21Rv3JV49pu3ln9attfKow0zDD/z15ELOKM1Pt/vUsOJJjMWR/znOpxT
8sfttsEG3CYi/SmxqdJNtp4SFE27sXQh0543GRw64AqhzK3C8UlKJRQNvKOj4/MU
Gf29Ujgr/1D+4By40xrMLsGwdWarBbs38mr8ScRYXBUrFx/BTzCcqLImE6qlqxOS
+Wdk471kx7fRR4IvjUV0+mGVITVWllEd9tiso8/XYrdLBPeu36CoqURsqJXY9Wwd
szN0HrXI1wjnsvow73l52q5BV1e7Hhjc0a4iEOYBjq579A7hpyaMOJCwr+jIKb/B
4j9uoLkUX9cYhF/TSL8PnmJ8QRCV118lRAg5pUC67jFi3jGfdzxXguJpAwRp4c+o
Lxj4TQ7DxOWVdPlcwzyCMyOICztROUwyFxhZ+RDa9B6hhGx5PhZzl+RfHQJzpab8
FudNLZUSmZchg3he7daNM+C++Ufun8KXz7XHGdHpNFrxqzKT3Mja8Ny/N5N3Kab+
Vc4CCQbduHSv4a0FzBECQN+cmFRIwaTbMtVRCH5mmGNo5i5/GO7kYFKunv3QsW0p
hZKPcWWrVYNu2u/HT4enDh+p1rWYt4B+f33kYD0ze8SPxmoQH9TZeXvjCyXCRr+5
c+rHDdfi70g2GfSsAJIVkMe1hsm0MI4S0ppYc7kYOvAxScsac8ubllmP/B531qTK
Lc2cLH/vn72kHIo98svDXXIrmyvKwe60vE3Bea7VE4GoW/IWqk6kDmnfIhgDQBsi
PAk6/949n4XFomn74ump3G6h9bTnXufMgNHqld1IaohoAMzEtrGDBTbdaVUe/73u
nCvmPRRP4f3A4SGawCYOle91QjAtwINWoOet/XmU7i6FG7fvoJj3DK2iKBlljzic
tvS3XIzpjhHVfiJE5brh8mrQT/DeclqznR/oOkzsIk2obqyv5v/+Vq/6vyKBG0+R
nys2NgfBASy/r7aNZBmOJGTH+0JGoY5mw/ilOHDIvOPJ2LehLAgltPcXlsr+BzAn
5E81i74M/rNnD7EJl1sL0JTnydBMb6+cAqgaCY3K2w+IRlAQQD/XQ3fHkGo3oTPs
PInzTUjmY+WVLswKescrFmhx8rfMffS2yf0fC7MNpNfTgGS2busquxRc+iupCZmm
2kD62q3Xfnku/nB3cUZt21QjHVNY1sWjDu3QX64inq6P2dqYcdyOTD1MgojUPwko
yL1YQwr8dNlRwMR7JMawL+un988D4tD+/jLlLDPCkLuv633xH+BcIuLT9hmqMB1T
NTu3j06U3egFEGFAUOU1M2Uo1rHy5XKEArmj2IiBPRJxWzSaP5uJ718U8o3YiOCx
uBW+VASljb3lqwmQMBd30jiOej7i5VQmtem45AfOHnMtZX5+6hB3CLrvxBxEJFD4
oizPB3uysbxMmZ79y361BZtR25H0bii5NnJpNXp+53IKA/e/CLDyLM0QCA/T4kfZ
cXFl1DjWse6zr+xnkSZQnTPOSGp6Ype3Nf8nKqTbQcNXRA+8HTVLR1P/oDhoakKY
nIXrqWg5TR4PYth4uPPnf0upSLrnbLDNWzh7J2dXrzBFleSTnyMoyah52pGYdpBr
gWa+hLuBT1YxkG2tcSJ2/ptUbzdtckkRaLMzLugBwf9x/JhMhSgY3SIY2h2KGDNv
uqwItu/nfsqzfX0N0J3bpxCEhHieUfGRT6mPGozNXlsuN5QXIsPI83IvG62w0PmK
LREzK/UfD6zo0rcT++FaoqgmD/VxrvHPFjDkPAaWjxg+vpd9GmHk/8ETDGeW5hqI
HT2XxdVjF6p9e/LooHfCv9j0CMw10C/z5UXY8Rnd16EaeaZ+aZmLmL4/anG96nkL
hByS7K1Zvoidn2DEJHAbxzjwjvkFo4KR2u+Fyw8xEn0mU0T8RI83m7hldBqAE0G7
N+smAOWyJp4oIR80c9Fvp2pYaQz4bbkHqmYfEY8d7k4vvfNn0rzUdFbC2E+2c4nt
jgZy51OqRIKbrLtK8q6BR37xku5eAQKuIOd9HOE8HUV6C3Ljgg+Vvigrcozlra81
W9A2E/467A+EC/XkYxaRn33/OjTy3iGqtSrotuRIHGeC1+o2JBVugv5LSVU/XdAg
6S6cY4ApAGrv9Z59BGcdYi4C44L5BKEwftzy2kiKSFZsxhHxbwO2cpxXohV0bF1H
XCadpWwloqsE8Rb9SASXxVpJvjQFs3WEZi709GD8iMN7y5TIFFllRhIQK5vQIQpD
pZ2mXNbl7JBryNg7x0JmJ76Rcm+970ZGcGI9Jt+4+IwO+iW6f91Lc1gC3BxYYD1T
sL2nfq5oDVX1D3QT814oa53gjStHP6ADBBROYXJqbkKqWb9cnRR4pul8MEj1HNTR
szt77n29jOxju8Z2JYyusNhRjXB4oOU+bnu3C7r4yC4WN9L6bpX1LupC88R1MLaL
wwid3vdPAxTnrstOF+2EHs0Q7McPdb9AeA85agrzZC07UQP6NdCaUepxbyo/oKSU
KTcd5+z56+b2oAUv2BN1vCczR7KN45Jgu11qdj/rcO6Vd0yMWSCgJ716H0kebBtM
IzllFw+H5mJ2HYAXM8JXvcr9e9AFtaqeykZibsqb8BY1OVoUIQfxJJHLE+P68ivV
JOkmOWVXZmmEGslhbQAEv+K9MdY4mE0pMk8tE94ssFVEicFnYcs5bbV5qjcYKG2I
Aijn+S8yKGRzGZh0PpdawF1aZINI9IXiSkkcJi7iJTDJKvbUsmPlmD20kZB1Euqr
rai8D0clptOztt9Di41BpNDWVHur/dsh2iPJJjOOD3/i3Nav9iR0UfvASelG4C6L
S6+6/S6z6leRNYEUPkQj1uCBIjuGEv/lbfKd5bAi0JSOaVoFzuOobY6IJsCwI57o
olT85nxJ57yrlHzs6Exs5Vrk/gPyDE1oiM+V3//TP76Rku9yyhrw/d/DTckaxZRU
qRDiIFXWxRi509ICYIUUpeiUFy8QT1i1WiBjoeEn+4UJADfpSr6etAVu2XLDl7EH
E+9PM2aA+eSvbtHteCftc1v500cvHcspU6YMdXcoWylfONjcFoO+r+JAxrgEclX2
z7yW+5H5p7dj/Y4xbcTMj8DuSp2F8CLr/djS8xeAHwgvncpAYMVBAUt+8jVGKmFe
Tw/1XvPfzsLQMFziEhx2CflLhlo11fez8ApjFbRqQVaGSOBOjse0WxaLzJyKKAY5
YtySU2ejra7l7qhei6gnvxCxeIPkQczpp4hE3k9OniZDwv6k9SDFPhOkuKMBi+UR
`protect end_protected
