localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTZNG_CHK = {
  {32'h4405adb8, 32'h444bf626} /* (31, 31, 31) {real, imag} */,
  {32'hc33947d5, 32'hc3070542} /* (31, 31, 30) {real, imag} */,
  {32'hc059f50f, 32'hc11e006d} /* (31, 31, 29) {real, imag} */,
  {32'h41e97e4d, 32'h4179d236} /* (31, 31, 28) {real, imag} */,
  {32'hc16f8cb4, 32'hc19a5db1} /* (31, 31, 27) {real, imag} */,
  {32'hc0a6d9e8, 32'hc14434ac} /* (31, 31, 26) {real, imag} */,
  {32'hbf46adf7, 32'h40b7705d} /* (31, 31, 25) {real, imag} */,
  {32'hc10c0492, 32'hbe293e34} /* (31, 31, 24) {real, imag} */,
  {32'hbe7b0c50, 32'hbfa6cd93} /* (31, 31, 23) {real, imag} */,
  {32'hc0a174a0, 32'hc004d2cd} /* (31, 31, 22) {real, imag} */,
  {32'hc0d14041, 32'h3f5e3097} /* (31, 31, 21) {real, imag} */,
  {32'hc0621ccf, 32'hbf87948f} /* (31, 31, 20) {real, imag} */,
  {32'h3f2e034e, 32'hbf172bc6} /* (31, 31, 19) {real, imag} */,
  {32'hc03ac907, 32'h3fd2971e} /* (31, 31, 18) {real, imag} */,
  {32'h400e7989, 32'h3e8dc66d} /* (31, 31, 17) {real, imag} */,
  {32'hbf012c87, 32'h3eb0fd6e} /* (31, 31, 16) {real, imag} */,
  {32'h3ea6d04a, 32'h3e9b3261} /* (31, 31, 15) {real, imag} */,
  {32'h3fcd27ac, 32'hbf22c772} /* (31, 31, 14) {real, imag} */,
  {32'hbf28da14, 32'h3ed6d99b} /* (31, 31, 13) {real, imag} */,
  {32'hbd427d46, 32'hbf6f415f} /* (31, 31, 12) {real, imag} */,
  {32'h40d1d4ce, 32'hc09a7b37} /* (31, 31, 11) {real, imag} */,
  {32'hbf8ff761, 32'h403afb85} /* (31, 31, 10) {real, imag} */,
  {32'h402bc7f7, 32'hc007357b} /* (31, 31, 9) {real, imag} */,
  {32'h40ea77af, 32'hc0ea43b7} /* (31, 31, 8) {real, imag} */,
  {32'hc017d079, 32'h4111a736} /* (31, 31, 7) {real, imag} */,
  {32'hc0845430, 32'h3dc1e6dc} /* (31, 31, 6) {real, imag} */,
  {32'hc0f80d9d, 32'hc1fc83b1} /* (31, 31, 5) {real, imag} */,
  {32'h418f91a2, 32'h41a2b5a5} /* (31, 31, 4) {real, imag} */,
  {32'h41621cac, 32'h410224ae} /* (31, 31, 3) {real, imag} */,
  {32'hc1ce3b51, 32'hc302df7d} /* (31, 31, 2) {real, imag} */,
  {32'hc2a80409, 32'h4416d8d6} /* (31, 31, 1) {real, imag} */,
  {32'h432eb4b6, 32'h44392af1} /* (31, 31, 0) {real, imag} */,
  {32'hc0a50780, 32'hc375fbf4} /* (31, 30, 31) {real, imag} */,
  {32'h3fab070e, 32'h42dd3cea} /* (31, 30, 30) {real, imag} */,
  {32'hc0590731, 32'h402281a9} /* (31, 30, 29) {real, imag} */,
  {32'hc153100e, 32'hc221904a} /* (31, 30, 28) {real, imag} */,
  {32'h41c99a66, 32'h41bcfbd2} /* (31, 30, 27) {real, imag} */,
  {32'h3f8d126f, 32'h408d7d53} /* (31, 30, 26) {real, imag} */,
  {32'hbfe4fe7e, 32'hc0974ea7} /* (31, 30, 25) {real, imag} */,
  {32'hc0136634, 32'hbe963717} /* (31, 30, 24) {real, imag} */,
  {32'h4068d29d, 32'h3dac41c5} /* (31, 30, 23) {real, imag} */,
  {32'h3f379520, 32'hbfa4baac} /* (31, 30, 22) {real, imag} */,
  {32'h40d15181, 32'hbed00a88} /* (31, 30, 21) {real, imag} */,
  {32'h3fc1d77e, 32'h3fcc5434} /* (31, 30, 20) {real, imag} */,
  {32'h3e79231f, 32'h3f2d7d20} /* (31, 30, 19) {real, imag} */,
  {32'h3f19226c, 32'h3fac12e0} /* (31, 30, 18) {real, imag} */,
  {32'hbe3828e9, 32'hbeff18f5} /* (31, 30, 17) {real, imag} */,
  {32'hbf0477ea, 32'h3f8195ac} /* (31, 30, 16) {real, imag} */,
  {32'h40250f7a, 32'hbf697eca} /* (31, 30, 15) {real, imag} */,
  {32'hc05871bf, 32'h3bed09ec} /* (31, 30, 14) {real, imag} */,
  {32'h3f172da3, 32'h40408e89} /* (31, 30, 13) {real, imag} */,
  {32'hbf1fc917, 32'hbfc8fc65} /* (31, 30, 12) {real, imag} */,
  {32'hc01c90d5, 32'h3f90f220} /* (31, 30, 11) {real, imag} */,
  {32'h400da93a, 32'h4030d079} /* (31, 30, 10) {real, imag} */,
  {32'h404b9db5, 32'hc015a8b2} /* (31, 30, 9) {real, imag} */,
  {32'hbfd155e6, 32'h3f5399b3} /* (31, 30, 8) {real, imag} */,
  {32'hc08b6286, 32'hc0ba04e2} /* (31, 30, 7) {real, imag} */,
  {32'hc07de68f, 32'h3fd86a91} /* (31, 30, 6) {real, imag} */,
  {32'hc0acfcf4, 32'h411da220} /* (31, 30, 5) {real, imag} */,
  {32'h41722c3e, 32'hc15751c0} /* (31, 30, 4) {real, imag} */,
  {32'h40e0cf33, 32'hbf9726d0} /* (31, 30, 3) {real, imag} */,
  {32'hc1c404b4, 32'h433dfba2} /* (31, 30, 2) {real, imag} */,
  {32'hc2618a05, 32'hc3cb743e} /* (31, 30, 1) {real, imag} */,
  {32'hc285841e, 32'hc34aebe0} /* (31, 30, 0) {real, imag} */,
  {32'h41f56310, 32'h41bafaa6} /* (31, 29, 31) {real, imag} */,
  {32'hc20a3ff3, 32'hc058c6da} /* (31, 29, 30) {real, imag} */,
  {32'hc05815b0, 32'hc0e3d64c} /* (31, 29, 29) {real, imag} */,
  {32'h409e1d60, 32'hc166a721} /* (31, 29, 28) {real, imag} */,
  {32'h3fdcc3eb, 32'h406cdbed} /* (31, 29, 27) {real, imag} */,
  {32'hc1099b50, 32'h40e2976f} /* (31, 29, 26) {real, imag} */,
  {32'hc0147cab, 32'hbfcce75d} /* (31, 29, 25) {real, imag} */,
  {32'h3f4a695e, 32'hbe2fd4c2} /* (31, 29, 24) {real, imag} */,
  {32'h40824be9, 32'hbfcf494b} /* (31, 29, 23) {real, imag} */,
  {32'hbf863e64, 32'h40172f33} /* (31, 29, 22) {real, imag} */,
  {32'hbfe3bb99, 32'h400fb292} /* (31, 29, 21) {real, imag} */,
  {32'h3fe3ca16, 32'h3efb83dd} /* (31, 29, 20) {real, imag} */,
  {32'hbe5fccb7, 32'h3f90e310} /* (31, 29, 19) {real, imag} */,
  {32'hbfd66753, 32'h3ec6802d} /* (31, 29, 18) {real, imag} */,
  {32'h3f8964d2, 32'h3ec77069} /* (31, 29, 17) {real, imag} */,
  {32'hbfaaa570, 32'h3da43bd3} /* (31, 29, 16) {real, imag} */,
  {32'h3fdc1770, 32'h402996f7} /* (31, 29, 15) {real, imag} */,
  {32'hbff14442, 32'hbf64b853} /* (31, 29, 14) {real, imag} */,
  {32'h3f0ba43b, 32'hbf1c3423} /* (31, 29, 13) {real, imag} */,
  {32'h3ec92e59, 32'hbeebc76e} /* (31, 29, 12) {real, imag} */,
  {32'hc005c1be, 32'h3f37f442} /* (31, 29, 11) {real, imag} */,
  {32'h405e795d, 32'hc043bee8} /* (31, 29, 10) {real, imag} */,
  {32'h3f879b70, 32'h3f8273ce} /* (31, 29, 9) {real, imag} */,
  {32'hc0a4e06e, 32'hc01438d0} /* (31, 29, 8) {real, imag} */,
  {32'h405b3196, 32'h3f994a0c} /* (31, 29, 7) {real, imag} */,
  {32'h400a7054, 32'hc05d7f5a} /* (31, 29, 6) {real, imag} */,
  {32'h409238b9, 32'hc0b11d43} /* (31, 29, 5) {real, imag} */,
  {32'h410533e4, 32'h4135567c} /* (31, 29, 4) {real, imag} */,
  {32'h40c34e79, 32'h3eda147a} /* (31, 29, 3) {real, imag} */,
  {32'hc22dba90, 32'h4208b6ca} /* (31, 29, 2) {real, imag} */,
  {32'h418db6d8, 32'hc23baebc} /* (31, 29, 1) {real, imag} */,
  {32'h3ffed618, 32'hc1415cf9} /* (31, 29, 0) {real, imag} */,
  {32'h4080ba3c, 32'h41e55f98} /* (31, 28, 31) {real, imag} */,
  {32'hc1be648c, 32'hc1d76d83} /* (31, 28, 30) {real, imag} */,
  {32'h41814fcb, 32'hc1321ad2} /* (31, 28, 29) {real, imag} */,
  {32'h41612e92, 32'hc095cb99} /* (31, 28, 28) {real, imag} */,
  {32'hc07946bc, 32'h3fba3d84} /* (31, 28, 27) {real, imag} */,
  {32'h403efcff, 32'h40c3cbde} /* (31, 28, 26) {real, imag} */,
  {32'hbe2ffc5f, 32'hbe487aaf} /* (31, 28, 25) {real, imag} */,
  {32'hc0aaeb2a, 32'hc0b1e5bd} /* (31, 28, 24) {real, imag} */,
  {32'h3f3cc9e2, 32'h3f9f90e3} /* (31, 28, 23) {real, imag} */,
  {32'hbfd289a8, 32'hbeceed64} /* (31, 28, 22) {real, imag} */,
  {32'hc083f46a, 32'hbfa28daf} /* (31, 28, 21) {real, imag} */,
  {32'h409ec28c, 32'h3fc3262d} /* (31, 28, 20) {real, imag} */,
  {32'h3f899e70, 32'h3ecb4847} /* (31, 28, 19) {real, imag} */,
  {32'hc04d7a1c, 32'hbf433794} /* (31, 28, 18) {real, imag} */,
  {32'hbe8a24b0, 32'hbf2e7925} /* (31, 28, 17) {real, imag} */,
  {32'h3f2985d7, 32'h3fae77c2} /* (31, 28, 16) {real, imag} */,
  {32'h3fa1ed52, 32'h3f3c3b56} /* (31, 28, 15) {real, imag} */,
  {32'hbfaa514c, 32'hbfcf95ad} /* (31, 28, 14) {real, imag} */,
  {32'hbee64a2a, 32'hc01c2c42} /* (31, 28, 13) {real, imag} */,
  {32'h3ff17d6c, 32'hbe3875cf} /* (31, 28, 12) {real, imag} */,
  {32'h3f8b48ef, 32'h4023b76e} /* (31, 28, 11) {real, imag} */,
  {32'hbf8e6661, 32'h3e064ef6} /* (31, 28, 10) {real, imag} */,
  {32'hc0270a20, 32'h3fe80d2c} /* (31, 28, 9) {real, imag} */,
  {32'hc110cfd6, 32'hc0921bb5} /* (31, 28, 8) {real, imag} */,
  {32'hbfb7549b, 32'h40cffe0b} /* (31, 28, 7) {real, imag} */,
  {32'h4091d70c, 32'hbf82f947} /* (31, 28, 6) {real, imag} */,
  {32'hbf435fcb, 32'hc0c3a4d3} /* (31, 28, 5) {real, imag} */,
  {32'h41158831, 32'h415843e9} /* (31, 28, 4) {real, imag} */,
  {32'hc03af72a, 32'hc0ba6b24} /* (31, 28, 3) {real, imag} */,
  {32'hc1dca5de, 32'hc2071833} /* (31, 28, 2) {real, imag} */,
  {32'h41d5ed1b, 32'hc078323f} /* (31, 28, 1) {real, imag} */,
  {32'h4146a760, 32'h41422e5c} /* (31, 28, 0) {real, imag} */,
  {32'hc1b22a28, 32'hc0e42970} /* (31, 27, 31) {real, imag} */,
  {32'h41ccb713, 32'h406f4438} /* (31, 27, 30) {real, imag} */,
  {32'h3ff1725d, 32'h3ef9ddc5} /* (31, 27, 29) {real, imag} */,
  {32'hc12c9a50, 32'hbf5efea8} /* (31, 27, 28) {real, imag} */,
  {32'h4015c1ba, 32'h40d4716e} /* (31, 27, 27) {real, imag} */,
  {32'h3fbce8f7, 32'hbfa8fd41} /* (31, 27, 26) {real, imag} */,
  {32'hc086d206, 32'hc07bd098} /* (31, 27, 25) {real, imag} */,
  {32'hbf568f22, 32'h3f9faa39} /* (31, 27, 24) {real, imag} */,
  {32'h4001d0c2, 32'hbfb513d3} /* (31, 27, 23) {real, imag} */,
  {32'h405915a5, 32'hbea3be6f} /* (31, 27, 22) {real, imag} */,
  {32'h3cdb3c01, 32'h3ffe8f55} /* (31, 27, 21) {real, imag} */,
  {32'hbfbbf870, 32'hbedf1e7d} /* (31, 27, 20) {real, imag} */,
  {32'h3f87685c, 32'h3f25df9a} /* (31, 27, 19) {real, imag} */,
  {32'h400a9a3f, 32'h3f11baf4} /* (31, 27, 18) {real, imag} */,
  {32'hbfe9e9cd, 32'h3fb7fca5} /* (31, 27, 17) {real, imag} */,
  {32'hbece53ad, 32'h3f4c4bed} /* (31, 27, 16) {real, imag} */,
  {32'hbfa7cd4e, 32'h3e797c2a} /* (31, 27, 15) {real, imag} */,
  {32'hc057bda1, 32'hc014a430} /* (31, 27, 14) {real, imag} */,
  {32'h3fab88fd, 32'hbf938f3b} /* (31, 27, 13) {real, imag} */,
  {32'h3e2f5e7b, 32'hbfd05a73} /* (31, 27, 12) {real, imag} */,
  {32'hbff60355, 32'h3eeb03bd} /* (31, 27, 11) {real, imag} */,
  {32'hbf9a132b, 32'hbbed0b6e} /* (31, 27, 10) {real, imag} */,
  {32'h3bfcc686, 32'h3f8532a3} /* (31, 27, 9) {real, imag} */,
  {32'hc071ed45, 32'hbfb8235a} /* (31, 27, 8) {real, imag} */,
  {32'h3fe81a00, 32'hc001856e} /* (31, 27, 7) {real, imag} */,
  {32'h40524e1d, 32'h401f3e23} /* (31, 27, 6) {real, imag} */,
  {32'h405feff4, 32'h40c76489} /* (31, 27, 5) {real, imag} */,
  {32'h404c158b, 32'h3fabf1b0} /* (31, 27, 4) {real, imag} */,
  {32'hbff953b3, 32'h3f5f9430} /* (31, 27, 3) {real, imag} */,
  {32'h407f630c, 32'h417451df} /* (31, 27, 2) {real, imag} */,
  {32'hbfc6fcba, 32'hc1ba6d4e} /* (31, 27, 1) {real, imag} */,
  {32'hc13ae3c2, 32'hc10a3851} /* (31, 27, 0) {real, imag} */,
  {32'hc058cc7e, 32'h3fec3245} /* (31, 26, 31) {real, imag} */,
  {32'hc0de9241, 32'hc0218deb} /* (31, 26, 30) {real, imag} */,
  {32'h4002a5e3, 32'hc0a02d2b} /* (31, 26, 29) {real, imag} */,
  {32'h401ff486, 32'h40083027} /* (31, 26, 28) {real, imag} */,
  {32'hbde99d7e, 32'hc030e0d1} /* (31, 26, 27) {real, imag} */,
  {32'h3dce4676, 32'hc06078bd} /* (31, 26, 26) {real, imag} */,
  {32'h404c5ec8, 32'h3fb7a113} /* (31, 26, 25) {real, imag} */,
  {32'h3d6a9425, 32'h3f15ac45} /* (31, 26, 24) {real, imag} */,
  {32'h407ccc96, 32'hc07fee99} /* (31, 26, 23) {real, imag} */,
  {32'h3f4ffa8e, 32'h40473037} /* (31, 26, 22) {real, imag} */,
  {32'h3edb90a8, 32'h403eca24} /* (31, 26, 21) {real, imag} */,
  {32'hbfff588c, 32'hbd0f3424} /* (31, 26, 20) {real, imag} */,
  {32'h3d68b3ec, 32'hbf7315c3} /* (31, 26, 19) {real, imag} */,
  {32'hbfa0d9be, 32'hbe52ab43} /* (31, 26, 18) {real, imag} */,
  {32'hbff8022d, 32'h3f1a4bf9} /* (31, 26, 17) {real, imag} */,
  {32'h3f89e255, 32'hbee28903} /* (31, 26, 16) {real, imag} */,
  {32'hbfcb168a, 32'hbf9cc199} /* (31, 26, 15) {real, imag} */,
  {32'h3ee36f8d, 32'hbf5e414f} /* (31, 26, 14) {real, imag} */,
  {32'h4006202b, 32'h401f55a8} /* (31, 26, 13) {real, imag} */,
  {32'hbe1af801, 32'hc02634e2} /* (31, 26, 12) {real, imag} */,
  {32'hbf469b5f, 32'h403f9ce4} /* (31, 26, 11) {real, imag} */,
  {32'hbdc43537, 32'h3f12d3af} /* (31, 26, 10) {real, imag} */,
  {32'hbfeec62b, 32'h40768424} /* (31, 26, 9) {real, imag} */,
  {32'h401080e0, 32'hc06530d6} /* (31, 26, 8) {real, imag} */,
  {32'h3f96787c, 32'hbfa0b8e5} /* (31, 26, 7) {real, imag} */,
  {32'h3f5503d7, 32'h402df677} /* (31, 26, 6) {real, imag} */,
  {32'h404727b2, 32'h406e5f86} /* (31, 26, 5) {real, imag} */,
  {32'hc07015b6, 32'hbf030fa1} /* (31, 26, 4) {real, imag} */,
  {32'h40754371, 32'h3f7e4ab9} /* (31, 26, 3) {real, imag} */,
  {32'hc0c015f3, 32'h3db64700} /* (31, 26, 2) {real, imag} */,
  {32'hc05d0c51, 32'hc0662491} /* (31, 26, 1) {real, imag} */,
  {32'h40e9f4dd, 32'h40526f8b} /* (31, 26, 0) {real, imag} */,
  {32'h4130aa83, 32'h4061b55e} /* (31, 25, 31) {real, imag} */,
  {32'hc0e0ad80, 32'hc06fde6f} /* (31, 25, 30) {real, imag} */,
  {32'hbf9ea797, 32'hc0314e01} /* (31, 25, 29) {real, imag} */,
  {32'h400e8ee2, 32'h3deb0e5d} /* (31, 25, 28) {real, imag} */,
  {32'h4079b545, 32'h3f858ecf} /* (31, 25, 27) {real, imag} */,
  {32'hbfd6aba3, 32'hbfe7b85e} /* (31, 25, 26) {real, imag} */,
  {32'h401528b8, 32'h3fe6a6ea} /* (31, 25, 25) {real, imag} */,
  {32'h3f6c39bc, 32'hbfcd7291} /* (31, 25, 24) {real, imag} */,
  {32'h40b6da70, 32'hbfa0b8ae} /* (31, 25, 23) {real, imag} */,
  {32'h3ff546cb, 32'h407459a1} /* (31, 25, 22) {real, imag} */,
  {32'hbf7bca81, 32'h402363fa} /* (31, 25, 21) {real, imag} */,
  {32'hc00b14c1, 32'hbefae141} /* (31, 25, 20) {real, imag} */,
  {32'hbe6a14c2, 32'hc049cdcb} /* (31, 25, 19) {real, imag} */,
  {32'hbf0f9621, 32'h3fc535a3} /* (31, 25, 18) {real, imag} */,
  {32'h3e4a8f08, 32'hbddee26a} /* (31, 25, 17) {real, imag} */,
  {32'h3fa09cf0, 32'hbf0139c8} /* (31, 25, 16) {real, imag} */,
  {32'h3f4d2ac3, 32'hbf154163} /* (31, 25, 15) {real, imag} */,
  {32'hbf8bcba3, 32'h3f903ad9} /* (31, 25, 14) {real, imag} */,
  {32'h3f764e5a, 32'h3eb4b5f8} /* (31, 25, 13) {real, imag} */,
  {32'hbf850c4c, 32'h3f9f8f57} /* (31, 25, 12) {real, imag} */,
  {32'h3f06a278, 32'hbf798add} /* (31, 25, 11) {real, imag} */,
  {32'h3fb78b39, 32'h3fe88e17} /* (31, 25, 10) {real, imag} */,
  {32'hc037a0b8, 32'hc0aef25e} /* (31, 25, 9) {real, imag} */,
  {32'hbf5f8b88, 32'hbf8ea523} /* (31, 25, 8) {real, imag} */,
  {32'hbf8bb162, 32'h3f82daaf} /* (31, 25, 7) {real, imag} */,
  {32'h3fe99f3a, 32'hbecd0f71} /* (31, 25, 6) {real, imag} */,
  {32'h3eb11e4c, 32'h3ee2d6f3} /* (31, 25, 5) {real, imag} */,
  {32'hc045ff83, 32'hbf530ac8} /* (31, 25, 4) {real, imag} */,
  {32'h3f8b6e18, 32'hc069308f} /* (31, 25, 3) {real, imag} */,
  {32'hc0c410b0, 32'hc0c58bb1} /* (31, 25, 2) {real, imag} */,
  {32'h3f5195d5, 32'h409dc796} /* (31, 25, 1) {real, imag} */,
  {32'h40fd9587, 32'h401b2a8b} /* (31, 25, 0) {real, imag} */,
  {32'hc0aa3801, 32'hc0a0fa9c} /* (31, 24, 31) {real, imag} */,
  {32'h40367e84, 32'h41037261} /* (31, 24, 30) {real, imag} */,
  {32'hbedec9e5, 32'hbe8e00d5} /* (31, 24, 29) {real, imag} */,
  {32'hc09cc120, 32'hc0cde85c} /* (31, 24, 28) {real, imag} */,
  {32'h40629544, 32'h3f90bb22} /* (31, 24, 27) {real, imag} */,
  {32'hc086f6f7, 32'hbfcb36d0} /* (31, 24, 26) {real, imag} */,
  {32'h40416878, 32'hbfbafdc3} /* (31, 24, 25) {real, imag} */,
  {32'h405ccb28, 32'h404c7dae} /* (31, 24, 24) {real, imag} */,
  {32'h3ff8efe3, 32'hbfaaf990} /* (31, 24, 23) {real, imag} */,
  {32'h3f7a487e, 32'h3febe1b4} /* (31, 24, 22) {real, imag} */,
  {32'hbfdf5dd4, 32'hbfcac007} /* (31, 24, 21) {real, imag} */,
  {32'hbf2f5895, 32'h3fd5f43c} /* (31, 24, 20) {real, imag} */,
  {32'h4020f0d6, 32'hbf5a1f2e} /* (31, 24, 19) {real, imag} */,
  {32'hbe8ad6a5, 32'hbdb78bc7} /* (31, 24, 18) {real, imag} */,
  {32'h3f8f3828, 32'hbfc6edc1} /* (31, 24, 17) {real, imag} */,
  {32'h3f932648, 32'h3fba007e} /* (31, 24, 16) {real, imag} */,
  {32'h3f5efda2, 32'hc008c90d} /* (31, 24, 15) {real, imag} */,
  {32'hbdb58dd1, 32'h4043946a} /* (31, 24, 14) {real, imag} */,
  {32'h3e86e151, 32'hbf5c5204} /* (31, 24, 13) {real, imag} */,
  {32'h3e20c76a, 32'h3fc6a66a} /* (31, 24, 12) {real, imag} */,
  {32'h3fae5eae, 32'h3ef80a72} /* (31, 24, 11) {real, imag} */,
  {32'h3fca3d71, 32'h3fec697e} /* (31, 24, 10) {real, imag} */,
  {32'hbf122d7e, 32'h3fbf6728} /* (31, 24, 9) {real, imag} */,
  {32'hbf0d9b54, 32'hc05627f4} /* (31, 24, 8) {real, imag} */,
  {32'h4014936d, 32'hc03044c4} /* (31, 24, 7) {real, imag} */,
  {32'h401eef85, 32'h3f94e423} /* (31, 24, 6) {real, imag} */,
  {32'hc00b83e8, 32'h41267ab1} /* (31, 24, 5) {real, imag} */,
  {32'h3fc812ed, 32'h3fc6c3b7} /* (31, 24, 4) {real, imag} */,
  {32'h3f8a314a, 32'hbfca0f8c} /* (31, 24, 3) {real, imag} */,
  {32'h3fcfe120, 32'h40ad4816} /* (31, 24, 2) {real, imag} */,
  {32'hc0e4bf63, 32'hc12190c1} /* (31, 24, 1) {real, imag} */,
  {32'hc08b7462, 32'hc08cebb7} /* (31, 24, 0) {real, imag} */,
  {32'h40927803, 32'h4007e91f} /* (31, 23, 31) {real, imag} */,
  {32'hc022b7ec, 32'h408af764} /* (31, 23, 30) {real, imag} */,
  {32'h3eb8022d, 32'h3f81821c} /* (31, 23, 29) {real, imag} */,
  {32'h403e0bdb, 32'hbf6a0a8b} /* (31, 23, 28) {real, imag} */,
  {32'hc0641535, 32'hc045ab8a} /* (31, 23, 27) {real, imag} */,
  {32'h3e7bb245, 32'hc0728afd} /* (31, 23, 26) {real, imag} */,
  {32'h404177b4, 32'h3f626274} /* (31, 23, 25) {real, imag} */,
  {32'h3f99e880, 32'hbdc7827d} /* (31, 23, 24) {real, imag} */,
  {32'h3ed54fad, 32'hbef0398b} /* (31, 23, 23) {real, imag} */,
  {32'hbf504fe9, 32'h3f93e724} /* (31, 23, 22) {real, imag} */,
  {32'hc00f7c54, 32'h3f1ba66b} /* (31, 23, 21) {real, imag} */,
  {32'h3f0eb261, 32'hbf8a9177} /* (31, 23, 20) {real, imag} */,
  {32'hbc2360d4, 32'h3f875a84} /* (31, 23, 19) {real, imag} */,
  {32'hc011ea36, 32'hbf87a171} /* (31, 23, 18) {real, imag} */,
  {32'hbef96ccc, 32'hc0403b1d} /* (31, 23, 17) {real, imag} */,
  {32'h404788e9, 32'h3e7b48b1} /* (31, 23, 16) {real, imag} */,
  {32'h402397ad, 32'h3faf1e95} /* (31, 23, 15) {real, imag} */,
  {32'hbe9410e9, 32'hbfcf9d71} /* (31, 23, 14) {real, imag} */,
  {32'hc01e491d, 32'hbfaeccc7} /* (31, 23, 13) {real, imag} */,
  {32'h3fdaef10, 32'h3f3ac462} /* (31, 23, 12) {real, imag} */,
  {32'h3e66ccf0, 32'h3fa36655} /* (31, 23, 11) {real, imag} */,
  {32'hbf834740, 32'h3f5fbddf} /* (31, 23, 10) {real, imag} */,
  {32'hbf9eda83, 32'h4010208c} /* (31, 23, 9) {real, imag} */,
  {32'hbfe0cbdc, 32'h3fbbc197} /* (31, 23, 8) {real, imag} */,
  {32'hbefc61ea, 32'hbe572340} /* (31, 23, 7) {real, imag} */,
  {32'hbf92ea80, 32'h40876faa} /* (31, 23, 6) {real, imag} */,
  {32'h3fa00ff2, 32'hc0673690} /* (31, 23, 5) {real, imag} */,
  {32'hbf1e17e8, 32'h3f83740a} /* (31, 23, 4) {real, imag} */,
  {32'hc049536b, 32'h3e28a974} /* (31, 23, 3) {real, imag} */,
  {32'hbf5e64ef, 32'h3e077887} /* (31, 23, 2) {real, imag} */,
  {32'h3feab4c5, 32'hc0557dc7} /* (31, 23, 1) {real, imag} */,
  {32'hc0e05343, 32'hc02f6bc9} /* (31, 23, 0) {real, imag} */,
  {32'h3ff86b9c, 32'h4053ba7a} /* (31, 22, 31) {real, imag} */,
  {32'hc08b10db, 32'h3f146348} /* (31, 22, 30) {real, imag} */,
  {32'h3fe8f4e2, 32'hbc188db3} /* (31, 22, 29) {real, imag} */,
  {32'h40483d5b, 32'hbf837128} /* (31, 22, 28) {real, imag} */,
  {32'hc06f0cb9, 32'h405dc255} /* (31, 22, 27) {real, imag} */,
  {32'h3fe3c034, 32'h3f9cbbe1} /* (31, 22, 26) {real, imag} */,
  {32'h401f594c, 32'hbd71f007} /* (31, 22, 25) {real, imag} */,
  {32'h3e47a747, 32'h400b7553} /* (31, 22, 24) {real, imag} */,
  {32'h3f5d4a88, 32'hbaeefa4e} /* (31, 22, 23) {real, imag} */,
  {32'hbfadaef9, 32'hc00ca718} /* (31, 22, 22) {real, imag} */,
  {32'hbff06e71, 32'h4023b567} /* (31, 22, 21) {real, imag} */,
  {32'h3dfbe87a, 32'h3ff78e78} /* (31, 22, 20) {real, imag} */,
  {32'h3e4be579, 32'hbef33953} /* (31, 22, 19) {real, imag} */,
  {32'h3ed4fd4f, 32'hbf17a100} /* (31, 22, 18) {real, imag} */,
  {32'h4022017d, 32'h3f291cf3} /* (31, 22, 17) {real, imag} */,
  {32'h3f6e457a, 32'hbf36445a} /* (31, 22, 16) {real, imag} */,
  {32'hbf90b800, 32'h3fccbb57} /* (31, 22, 15) {real, imag} */,
  {32'hbf2817bf, 32'hbf0571a1} /* (31, 22, 14) {real, imag} */,
  {32'h402fa7b5, 32'hbfa22842} /* (31, 22, 13) {real, imag} */,
  {32'hbeeee40b, 32'hc0568f1c} /* (31, 22, 12) {real, imag} */,
  {32'hc046052b, 32'h3fff85a5} /* (31, 22, 11) {real, imag} */,
  {32'h3fe9afc7, 32'hbe80e91a} /* (31, 22, 10) {real, imag} */,
  {32'hc01da3a3, 32'h4004b322} /* (31, 22, 9) {real, imag} */,
  {32'h3f02d428, 32'h3f6cc8aa} /* (31, 22, 8) {real, imag} */,
  {32'h3f711ce8, 32'h3ef4d81f} /* (31, 22, 7) {real, imag} */,
  {32'h4004154f, 32'h402d5da7} /* (31, 22, 6) {real, imag} */,
  {32'h40841d70, 32'h3ee6d711} /* (31, 22, 5) {real, imag} */,
  {32'h4007395e, 32'h4029f354} /* (31, 22, 4) {real, imag} */,
  {32'h3fb9257a, 32'hc03af9b5} /* (31, 22, 3) {real, imag} */,
  {32'hc0780fa5, 32'hc0748377} /* (31, 22, 2) {real, imag} */,
  {32'h40383bde, 32'h3ff3419e} /* (31, 22, 1) {real, imag} */,
  {32'h3f87df4f, 32'h3f76ce24} /* (31, 22, 0) {real, imag} */,
  {32'hc09ad55e, 32'hbfecabb5} /* (31, 21, 31) {real, imag} */,
  {32'h40419d4e, 32'hc012050c} /* (31, 21, 30) {real, imag} */,
  {32'h3f8fc082, 32'hbf832640} /* (31, 21, 29) {real, imag} */,
  {32'hc0037859, 32'h3f834568} /* (31, 21, 28) {real, imag} */,
  {32'h3fb04ea7, 32'hbf4cbff6} /* (31, 21, 27) {real, imag} */,
  {32'hbf8dfe58, 32'h3ff32a04} /* (31, 21, 26) {real, imag} */,
  {32'hbd9e9074, 32'h3f607380} /* (31, 21, 25) {real, imag} */,
  {32'h3e81d1f1, 32'h3fd3d129} /* (31, 21, 24) {real, imag} */,
  {32'hbf8f6823, 32'h3f292a38} /* (31, 21, 23) {real, imag} */,
  {32'hbfa4ffdc, 32'hc03a709f} /* (31, 21, 22) {real, imag} */,
  {32'hbf3dd551, 32'hc01c7065} /* (31, 21, 21) {real, imag} */,
  {32'hbde2ca78, 32'h3dc8e9d0} /* (31, 21, 20) {real, imag} */,
  {32'hbfcd8d40, 32'h3eca8e77} /* (31, 21, 19) {real, imag} */,
  {32'h3f565db2, 32'h3f0d8b98} /* (31, 21, 18) {real, imag} */,
  {32'hbf4d43cd, 32'h3fb6c910} /* (31, 21, 17) {real, imag} */,
  {32'h3f852f3a, 32'h3d0b5d9d} /* (31, 21, 16) {real, imag} */,
  {32'h3efc86d5, 32'h3f74eb7a} /* (31, 21, 15) {real, imag} */,
  {32'hbf1397f7, 32'h3d01140d} /* (31, 21, 14) {real, imag} */,
  {32'hbf34e7ff, 32'hbe8b16fc} /* (31, 21, 13) {real, imag} */,
  {32'h3f7d20e4, 32'h3f5834bb} /* (31, 21, 12) {real, imag} */,
  {32'h3f835bfe, 32'h40008c23} /* (31, 21, 11) {real, imag} */,
  {32'hc016e5a9, 32'hbf920683} /* (31, 21, 10) {real, imag} */,
  {32'hbe377a29, 32'hc003977a} /* (31, 21, 9) {real, imag} */,
  {32'hbec17e94, 32'h3eafcf2c} /* (31, 21, 8) {real, imag} */,
  {32'hbf177472, 32'hc07d9559} /* (31, 21, 7) {real, imag} */,
  {32'h3f710ad3, 32'hbea186ca} /* (31, 21, 6) {real, imag} */,
  {32'hbe3154de, 32'h405a8b84} /* (31, 21, 5) {real, imag} */,
  {32'h3f67b5b8, 32'h3eb3606f} /* (31, 21, 4) {real, imag} */,
  {32'h3e581771, 32'hc021ad13} /* (31, 21, 3) {real, imag} */,
  {32'h4072ac32, 32'h406711e1} /* (31, 21, 2) {real, imag} */,
  {32'hbf2f07d3, 32'hc0a56eac} /* (31, 21, 1) {real, imag} */,
  {32'hc081f377, 32'hbe83a5ce} /* (31, 21, 0) {real, imag} */,
  {32'hc0281452, 32'h3fc841a0} /* (31, 20, 31) {real, imag} */,
  {32'h3f5c0785, 32'h3f8aff8b} /* (31, 20, 30) {real, imag} */,
  {32'h3ea80f8a, 32'hc0210cde} /* (31, 20, 29) {real, imag} */,
  {32'hbf6a199e, 32'hbea85265} /* (31, 20, 28) {real, imag} */,
  {32'hbd708314, 32'h401bec0c} /* (31, 20, 27) {real, imag} */,
  {32'h3f8c940c, 32'hbd18770e} /* (31, 20, 26) {real, imag} */,
  {32'hbf518937, 32'hbfe428e3} /* (31, 20, 25) {real, imag} */,
  {32'hc01b1edf, 32'hbd126bdd} /* (31, 20, 24) {real, imag} */,
  {32'h401b1a7b, 32'h4087fdda} /* (31, 20, 23) {real, imag} */,
  {32'hbebd38b6, 32'h4049d19e} /* (31, 20, 22) {real, imag} */,
  {32'hc00d171c, 32'h3fa6fcf1} /* (31, 20, 21) {real, imag} */,
  {32'hbf0e85d5, 32'hbf242ca9} /* (31, 20, 20) {real, imag} */,
  {32'hbe385614, 32'hbfd9d3b7} /* (31, 20, 19) {real, imag} */,
  {32'h3e4ecdc5, 32'hbf0c97af} /* (31, 20, 18) {real, imag} */,
  {32'hbf1f00aa, 32'hbfb4b894} /* (31, 20, 17) {real, imag} */,
  {32'hbf312fc1, 32'h3ceb4557} /* (31, 20, 16) {real, imag} */,
  {32'hbf804afc, 32'hbfd67960} /* (31, 20, 15) {real, imag} */,
  {32'h3f318f27, 32'h3f7f0be5} /* (31, 20, 14) {real, imag} */,
  {32'hbef14f25, 32'hbf29a2af} /* (31, 20, 13) {real, imag} */,
  {32'hbfcabdf1, 32'hbf221f17} /* (31, 20, 12) {real, imag} */,
  {32'h3fcf6b8a, 32'hbe8e3d54} /* (31, 20, 11) {real, imag} */,
  {32'h40060663, 32'h3e97fe70} /* (31, 20, 10) {real, imag} */,
  {32'h3f2dc7ec, 32'hc03b4397} /* (31, 20, 9) {real, imag} */,
  {32'hc02e5013, 32'h3f6dba1f} /* (31, 20, 8) {real, imag} */,
  {32'hc03c82a4, 32'h404243f2} /* (31, 20, 7) {real, imag} */,
  {32'hbf3edac1, 32'hbddf9a73} /* (31, 20, 6) {real, imag} */,
  {32'h3faa9b83, 32'hbfbf59ae} /* (31, 20, 5) {real, imag} */,
  {32'h3ddcfd07, 32'hbf75bbb1} /* (31, 20, 4) {real, imag} */,
  {32'h3ec55d64, 32'h40069a28} /* (31, 20, 3) {real, imag} */,
  {32'hbdcf253f, 32'hbef2144c} /* (31, 20, 2) {real, imag} */,
  {32'h402be7f6, 32'h405be44d} /* (31, 20, 1) {real, imag} */,
  {32'h3fe85382, 32'hbf21c761} /* (31, 20, 0) {real, imag} */,
  {32'h40844eaa, 32'h400205b5} /* (31, 19, 31) {real, imag} */,
  {32'hbedc0e59, 32'h400635d4} /* (31, 19, 30) {real, imag} */,
  {32'h3f7b1889, 32'hbfcedea3} /* (31, 19, 29) {real, imag} */,
  {32'hbe97d612, 32'hbdc89d0d} /* (31, 19, 28) {real, imag} */,
  {32'hbe1d7700, 32'hbea377a5} /* (31, 19, 27) {real, imag} */,
  {32'hc0390e8f, 32'h4006f539} /* (31, 19, 26) {real, imag} */,
  {32'hbead4c9a, 32'hbfee9c78} /* (31, 19, 25) {real, imag} */,
  {32'hc04aee14, 32'hc004d974} /* (31, 19, 24) {real, imag} */,
  {32'hbfa36183, 32'hbe19e99d} /* (31, 19, 23) {real, imag} */,
  {32'hbf74ef1e, 32'hbf1b483e} /* (31, 19, 22) {real, imag} */,
  {32'h3f0b9ea0, 32'hbedcabef} /* (31, 19, 21) {real, imag} */,
  {32'h3ef6d26f, 32'hbf4c55f8} /* (31, 19, 20) {real, imag} */,
  {32'h401d2eff, 32'h3fc5e022} /* (31, 19, 19) {real, imag} */,
  {32'h400b426b, 32'hc00093c4} /* (31, 19, 18) {real, imag} */,
  {32'hbfc5d692, 32'h3fd0a0e1} /* (31, 19, 17) {real, imag} */,
  {32'h3d573b05, 32'hbfc8c1ed} /* (31, 19, 16) {real, imag} */,
  {32'hbee31729, 32'h3f58676c} /* (31, 19, 15) {real, imag} */,
  {32'h3eaede22, 32'hbe35d315} /* (31, 19, 14) {real, imag} */,
  {32'hbf844687, 32'h3f654d37} /* (31, 19, 13) {real, imag} */,
  {32'hbfe70951, 32'hc0264706} /* (31, 19, 12) {real, imag} */,
  {32'hbfc37fdc, 32'hbeadc67a} /* (31, 19, 11) {real, imag} */,
  {32'hbfa0868a, 32'h3fcb0574} /* (31, 19, 10) {real, imag} */,
  {32'hbf008dea, 32'hc05baede} /* (31, 19, 9) {real, imag} */,
  {32'h3f29cf4f, 32'h3d9045fe} /* (31, 19, 8) {real, imag} */,
  {32'hbfe0116e, 32'h3f22d718} /* (31, 19, 7) {real, imag} */,
  {32'h40438ab0, 32'h3f945489} /* (31, 19, 6) {real, imag} */,
  {32'hbfa0e682, 32'hc0448c96} /* (31, 19, 5) {real, imag} */,
  {32'h3feb8fbe, 32'h3f0c2d0e} /* (31, 19, 4) {real, imag} */,
  {32'h3fbccd12, 32'hbe596391} /* (31, 19, 3) {real, imag} */,
  {32'h4063bfe1, 32'h40155108} /* (31, 19, 2) {real, imag} */,
  {32'hc095af5f, 32'h3ffb872f} /* (31, 19, 1) {real, imag} */,
  {32'h3fd5a783, 32'hbf70286c} /* (31, 19, 0) {real, imag} */,
  {32'hc076de31, 32'h3ff22aa6} /* (31, 18, 31) {real, imag} */,
  {32'h3f5f58fe, 32'h3ecbeb24} /* (31, 18, 30) {real, imag} */,
  {32'hbf10b1c4, 32'hc002c461} /* (31, 18, 29) {real, imag} */,
  {32'hbfce6a82, 32'hbf44bc23} /* (31, 18, 28) {real, imag} */,
  {32'h40565eb0, 32'h3ddf41ba} /* (31, 18, 27) {real, imag} */,
  {32'h4015912a, 32'hc01af90c} /* (31, 18, 26) {real, imag} */,
  {32'hc0175c19, 32'hbf5ad9bd} /* (31, 18, 25) {real, imag} */,
  {32'hbf3dc827, 32'hbe88e968} /* (31, 18, 24) {real, imag} */,
  {32'h3e15e754, 32'hbf33df29} /* (31, 18, 23) {real, imag} */,
  {32'hbfe7c218, 32'hbee777cd} /* (31, 18, 22) {real, imag} */,
  {32'h3eb88052, 32'hbfb3d030} /* (31, 18, 21) {real, imag} */,
  {32'h3e9112c0, 32'hbf5aa8a4} /* (31, 18, 20) {real, imag} */,
  {32'hbfa59bd5, 32'hbebac522} /* (31, 18, 19) {real, imag} */,
  {32'h400ef1e0, 32'h3e57b842} /* (31, 18, 18) {real, imag} */,
  {32'h3fa800cd, 32'h3d83b4f4} /* (31, 18, 17) {real, imag} */,
  {32'h3f11de77, 32'hbe7237cc} /* (31, 18, 16) {real, imag} */,
  {32'hbe831669, 32'hbee3ac8e} /* (31, 18, 15) {real, imag} */,
  {32'hbf4d13da, 32'hbf9d1270} /* (31, 18, 14) {real, imag} */,
  {32'hbf6d719b, 32'h3f87c7bf} /* (31, 18, 13) {real, imag} */,
  {32'hbd98c70f, 32'h40113816} /* (31, 18, 12) {real, imag} */,
  {32'h3f5ebc46, 32'h3fd11bc5} /* (31, 18, 11) {real, imag} */,
  {32'h3e45186e, 32'hbe99809b} /* (31, 18, 10) {real, imag} */,
  {32'hbfd2dc28, 32'hbf926134} /* (31, 18, 9) {real, imag} */,
  {32'h3d34b848, 32'h3f37f462} /* (31, 18, 8) {real, imag} */,
  {32'hbf706505, 32'hbe05660d} /* (31, 18, 7) {real, imag} */,
  {32'hbebe1b96, 32'h3f7e3aa6} /* (31, 18, 6) {real, imag} */,
  {32'h3f835cbe, 32'hbfc09175} /* (31, 18, 5) {real, imag} */,
  {32'h3f2b2b68, 32'hbfbd7477} /* (31, 18, 4) {real, imag} */,
  {32'h3f3dfc67, 32'h3e90c3c5} /* (31, 18, 3) {real, imag} */,
  {32'h3d992927, 32'h3fa37dca} /* (31, 18, 2) {real, imag} */,
  {32'hc08be964, 32'h3fb1996a} /* (31, 18, 1) {real, imag} */,
  {32'hc0228f13, 32'h4032571e} /* (31, 18, 0) {real, imag} */,
  {32'h40113d7b, 32'hbe6c9b0d} /* (31, 17, 31) {real, imag} */,
  {32'hbfcd813e, 32'hbf933277} /* (31, 17, 30) {real, imag} */,
  {32'hbf513254, 32'h4002e7cb} /* (31, 17, 29) {real, imag} */,
  {32'h3f6f33c2, 32'hbeeb684a} /* (31, 17, 28) {real, imag} */,
  {32'hbf1fc5b7, 32'hbf40de12} /* (31, 17, 27) {real, imag} */,
  {32'h3f3acfa1, 32'hbf0814ce} /* (31, 17, 26) {real, imag} */,
  {32'h3f0e39d7, 32'hbf7a8231} /* (31, 17, 25) {real, imag} */,
  {32'hbfcecff6, 32'h3fa30fbb} /* (31, 17, 24) {real, imag} */,
  {32'hbfb2d781, 32'h3f488efb} /* (31, 17, 23) {real, imag} */,
  {32'hbc85630a, 32'h3f95419f} /* (31, 17, 22) {real, imag} */,
  {32'h3d6426e1, 32'h3e94d071} /* (31, 17, 21) {real, imag} */,
  {32'hbda750aa, 32'h3f03a6ab} /* (31, 17, 20) {real, imag} */,
  {32'hbfcbe16a, 32'h3f94b9ff} /* (31, 17, 19) {real, imag} */,
  {32'hbea8d9f1, 32'hbeef1dc6} /* (31, 17, 18) {real, imag} */,
  {32'hbddd7fd4, 32'hbf69ced5} /* (31, 17, 17) {real, imag} */,
  {32'h3fc1cdec, 32'h3f45b93d} /* (31, 17, 16) {real, imag} */,
  {32'hbec5f17f, 32'hbe11d6ab} /* (31, 17, 15) {real, imag} */,
  {32'h3e5514cf, 32'h3f0a4226} /* (31, 17, 14) {real, imag} */,
  {32'hbf8c6498, 32'h3f9a2591} /* (31, 17, 13) {real, imag} */,
  {32'h3f015bae, 32'hbff5b649} /* (31, 17, 12) {real, imag} */,
  {32'h402c9471, 32'hc0350bed} /* (31, 17, 11) {real, imag} */,
  {32'hbfd73cc1, 32'hc051650b} /* (31, 17, 10) {real, imag} */,
  {32'hbdebb25d, 32'hbed0b2ea} /* (31, 17, 9) {real, imag} */,
  {32'hbe3afc1b, 32'hbde7e8a3} /* (31, 17, 8) {real, imag} */,
  {32'h3db0f2fd, 32'hc00e383e} /* (31, 17, 7) {real, imag} */,
  {32'h3fb615ab, 32'h3e08fa40} /* (31, 17, 6) {real, imag} */,
  {32'h3fc23fef, 32'h40014e71} /* (31, 17, 5) {real, imag} */,
  {32'h3f2636eb, 32'h3ffe5f3e} /* (31, 17, 4) {real, imag} */,
  {32'hbe83e5a8, 32'h3fad6794} /* (31, 17, 3) {real, imag} */,
  {32'hbf3ab295, 32'h3db1cbce} /* (31, 17, 2) {real, imag} */,
  {32'h3e412b34, 32'h3f56f2fc} /* (31, 17, 1) {real, imag} */,
  {32'h3f100cee, 32'h3f8016d5} /* (31, 17, 0) {real, imag} */,
  {32'h3f9085fe, 32'hbed3b0e6} /* (31, 16, 31) {real, imag} */,
  {32'hbf307ae3, 32'h3f11e38a} /* (31, 16, 30) {real, imag} */,
  {32'hbf6da3c7, 32'hbeb481a6} /* (31, 16, 29) {real, imag} */,
  {32'hbf1512c6, 32'hbf3b1cea} /* (31, 16, 28) {real, imag} */,
  {32'hbf5b1f2b, 32'h3ecfbc1b} /* (31, 16, 27) {real, imag} */,
  {32'hbf890f30, 32'h3de5e854} /* (31, 16, 26) {real, imag} */,
  {32'hbe4d37c2, 32'h3f2e36cf} /* (31, 16, 25) {real, imag} */,
  {32'h3fad19c6, 32'h3f92073d} /* (31, 16, 24) {real, imag} */,
  {32'h3fd406f6, 32'hbdda1ae2} /* (31, 16, 23) {real, imag} */,
  {32'hbc9c7f25, 32'hbefbf6f1} /* (31, 16, 22) {real, imag} */,
  {32'h3fc3a467, 32'h3f74089e} /* (31, 16, 21) {real, imag} */,
  {32'hbf1695d1, 32'h3fa75c2e} /* (31, 16, 20) {real, imag} */,
  {32'h3f95b8b3, 32'h3f68c66b} /* (31, 16, 19) {real, imag} */,
  {32'h3f8bcd92, 32'hbe9ef901} /* (31, 16, 18) {real, imag} */,
  {32'hc007b5ae, 32'h3ff2fa12} /* (31, 16, 17) {real, imag} */,
  {32'h3f1392e1, 32'h3ed7fdcd} /* (31, 16, 16) {real, imag} */,
  {32'hbd87c77d, 32'h3f8c80bb} /* (31, 16, 15) {real, imag} */,
  {32'hbf6de832, 32'hbfee736c} /* (31, 16, 14) {real, imag} */,
  {32'hbfbd17c6, 32'h3f4ef2ed} /* (31, 16, 13) {real, imag} */,
  {32'h3fafd41b, 32'hbd11291e} /* (31, 16, 12) {real, imag} */,
  {32'hbfa36618, 32'hbf730f3b} /* (31, 16, 11) {real, imag} */,
  {32'h3b61ff91, 32'h3faddc8c} /* (31, 16, 10) {real, imag} */,
  {32'hbfb42fb1, 32'hbdaac685} /* (31, 16, 9) {real, imag} */,
  {32'hbe519ca3, 32'hbff58a40} /* (31, 16, 8) {real, imag} */,
  {32'hbf2b9441, 32'h3fa1184c} /* (31, 16, 7) {real, imag} */,
  {32'h3fd937b4, 32'hbf7fef36} /* (31, 16, 6) {real, imag} */,
  {32'h3e21a2fe, 32'h3e96422e} /* (31, 16, 5) {real, imag} */,
  {32'h3eaa0ed8, 32'hbe027f0b} /* (31, 16, 4) {real, imag} */,
  {32'h3fd80838, 32'hbf2d16d4} /* (31, 16, 3) {real, imag} */,
  {32'h3f475e26, 32'hc0258797} /* (31, 16, 2) {real, imag} */,
  {32'h3f818d20, 32'hbef86f0a} /* (31, 16, 1) {real, imag} */,
  {32'hbe79f132, 32'h3ea9a70e} /* (31, 16, 0) {real, imag} */,
  {32'hbffdbb20, 32'hbfbd54aa} /* (31, 15, 31) {real, imag} */,
  {32'h3f1c99b3, 32'hbe98287c} /* (31, 15, 30) {real, imag} */,
  {32'h3f4e7403, 32'hbcf6c35b} /* (31, 15, 29) {real, imag} */,
  {32'hbfd64d13, 32'h3f2d804b} /* (31, 15, 28) {real, imag} */,
  {32'h3f75a701, 32'hbec1e93a} /* (31, 15, 27) {real, imag} */,
  {32'h40422c14, 32'h3f80769a} /* (31, 15, 26) {real, imag} */,
  {32'hbf1f985c, 32'hbf61908e} /* (31, 15, 25) {real, imag} */,
  {32'h401b9d7d, 32'h3dd138f0} /* (31, 15, 24) {real, imag} */,
  {32'hbf31f466, 32'hc01a7d58} /* (31, 15, 23) {real, imag} */,
  {32'h3fef9670, 32'h3f907e41} /* (31, 15, 22) {real, imag} */,
  {32'h3f068662, 32'hbf8d4ded} /* (31, 15, 21) {real, imag} */,
  {32'h3de5b477, 32'h3f81fe94} /* (31, 15, 20) {real, imag} */,
  {32'h3f68760e, 32'hbfbccfa3} /* (31, 15, 19) {real, imag} */,
  {32'hbf2a57ec, 32'hbf73b83f} /* (31, 15, 18) {real, imag} */,
  {32'hbd02e3f1, 32'h3e217ad9} /* (31, 15, 17) {real, imag} */,
  {32'hbeb0d866, 32'hbf3c11a3} /* (31, 15, 16) {real, imag} */,
  {32'hbe4b9c02, 32'h3e97d001} /* (31, 15, 15) {real, imag} */,
  {32'hbfeae86e, 32'h3f8c8087} /* (31, 15, 14) {real, imag} */,
  {32'h3e05868a, 32'h3f986e1d} /* (31, 15, 13) {real, imag} */,
  {32'hbf9b9b8d, 32'h3eba8858} /* (31, 15, 12) {real, imag} */,
  {32'h3f8ce65b, 32'hbfbc80e1} /* (31, 15, 11) {real, imag} */,
  {32'h3f213c95, 32'hbe94319a} /* (31, 15, 10) {real, imag} */,
  {32'hbf19ccfc, 32'h3fb9f420} /* (31, 15, 9) {real, imag} */,
  {32'hbfd179ef, 32'hc0203834} /* (31, 15, 8) {real, imag} */,
  {32'h3ee012ab, 32'hbf7c804b} /* (31, 15, 7) {real, imag} */,
  {32'h3dd490f4, 32'h3f672149} /* (31, 15, 6) {real, imag} */,
  {32'hbfdd1932, 32'hbe9c9b8e} /* (31, 15, 5) {real, imag} */,
  {32'h3f3e935e, 32'hbf0466b2} /* (31, 15, 4) {real, imag} */,
  {32'hbf3bcaa4, 32'h3eb76db7} /* (31, 15, 3) {real, imag} */,
  {32'hbe8d62db, 32'h3ebbc0cb} /* (31, 15, 2) {real, imag} */,
  {32'hbec3162a, 32'h3f08169a} /* (31, 15, 1) {real, imag} */,
  {32'hc01b169f, 32'hbec713ee} /* (31, 15, 0) {real, imag} */,
  {32'h402cbae6, 32'hc0014c0f} /* (31, 14, 31) {real, imag} */,
  {32'hbf669dd1, 32'h3f955736} /* (31, 14, 30) {real, imag} */,
  {32'hbef711bf, 32'hc0033f55} /* (31, 14, 29) {real, imag} */,
  {32'hbe4d7cf6, 32'hbfe78d14} /* (31, 14, 28) {real, imag} */,
  {32'hbf6727ff, 32'h3e5e2dc6} /* (31, 14, 27) {real, imag} */,
  {32'hbfb78726, 32'hbdbb57e1} /* (31, 14, 26) {real, imag} */,
  {32'h3f86b93e, 32'h3e6473d6} /* (31, 14, 25) {real, imag} */,
  {32'h3ff71bce, 32'h404948d8} /* (31, 14, 24) {real, imag} */,
  {32'hc02a21f9, 32'hbf8d07e0} /* (31, 14, 23) {real, imag} */,
  {32'h3da57182, 32'hbeb2b789} /* (31, 14, 22) {real, imag} */,
  {32'h3e8298a4, 32'h400b21af} /* (31, 14, 21) {real, imag} */,
  {32'h3b47e049, 32'hbfd21971} /* (31, 14, 20) {real, imag} */,
  {32'h3fe8829c, 32'h3ed19077} /* (31, 14, 19) {real, imag} */,
  {32'h3e0fab20, 32'hbdbc912d} /* (31, 14, 18) {real, imag} */,
  {32'hc0083aae, 32'hbe2d26a8} /* (31, 14, 17) {real, imag} */,
  {32'h3f68e0b7, 32'hbfc29364} /* (31, 14, 16) {real, imag} */,
  {32'hbeb253d9, 32'h3f8c1b00} /* (31, 14, 15) {real, imag} */,
  {32'hbfa46a65, 32'hc0046b4a} /* (31, 14, 14) {real, imag} */,
  {32'h3faf9b77, 32'h3f14bd06} /* (31, 14, 13) {real, imag} */,
  {32'hbfd51c94, 32'h3e95d55b} /* (31, 14, 12) {real, imag} */,
  {32'hbe9401dd, 32'hc0171320} /* (31, 14, 11) {real, imag} */,
  {32'hbfd71641, 32'hbc69f29b} /* (31, 14, 10) {real, imag} */,
  {32'h40211688, 32'h3d5cf583} /* (31, 14, 9) {real, imag} */,
  {32'hbe8f17ba, 32'hbf4cf01b} /* (31, 14, 8) {real, imag} */,
  {32'hbfa2f7e4, 32'h3fe8b479} /* (31, 14, 7) {real, imag} */,
  {32'hbf025edb, 32'h3fbf652f} /* (31, 14, 6) {real, imag} */,
  {32'hbfe0fabd, 32'hbf307440} /* (31, 14, 5) {real, imag} */,
  {32'hc00270c8, 32'h3f2973c7} /* (31, 14, 4) {real, imag} */,
  {32'h3fcb772f, 32'hbd4b9d6f} /* (31, 14, 3) {real, imag} */,
  {32'hbf0b8032, 32'h3f81b975} /* (31, 14, 2) {real, imag} */,
  {32'h4072e479, 32'h3fb1aecb} /* (31, 14, 1) {real, imag} */,
  {32'h4015d953, 32'hbf9cc1a7} /* (31, 14, 0) {real, imag} */,
  {32'hc00cf4b2, 32'hc0360934} /* (31, 13, 31) {real, imag} */,
  {32'hbf6bea67, 32'h3f93e232} /* (31, 13, 30) {real, imag} */,
  {32'hbf46de87, 32'h3f609c20} /* (31, 13, 29) {real, imag} */,
  {32'hbe957ee5, 32'hbf0cbb5e} /* (31, 13, 28) {real, imag} */,
  {32'h3ecc777f, 32'hbf5e0468} /* (31, 13, 27) {real, imag} */,
  {32'h40665c13, 32'hbf9c669f} /* (31, 13, 26) {real, imag} */,
  {32'h3ffb223b, 32'h4082d8db} /* (31, 13, 25) {real, imag} */,
  {32'h3f3ba730, 32'h3fe67f4d} /* (31, 13, 24) {real, imag} */,
  {32'hbf86d0c5, 32'hbf93ddb4} /* (31, 13, 23) {real, imag} */,
  {32'h3fd93500, 32'hc0158e9c} /* (31, 13, 22) {real, imag} */,
  {32'hbe61a32b, 32'h3e8311f3} /* (31, 13, 21) {real, imag} */,
  {32'hbf9b5291, 32'hbe9c4a0a} /* (31, 13, 20) {real, imag} */,
  {32'hbf294d70, 32'hbd134101} /* (31, 13, 19) {real, imag} */,
  {32'hbf7dc642, 32'hbfdfa624} /* (31, 13, 18) {real, imag} */,
  {32'hbeab23b5, 32'hbfbb2c7f} /* (31, 13, 17) {real, imag} */,
  {32'hbed0a384, 32'hbf4b93f5} /* (31, 13, 16) {real, imag} */,
  {32'h3faf6e2e, 32'hbf4c4b95} /* (31, 13, 15) {real, imag} */,
  {32'hbf9dab7c, 32'h3d63623e} /* (31, 13, 14) {real, imag} */,
  {32'hc032bfcf, 32'h3f7cccbf} /* (31, 13, 13) {real, imag} */,
  {32'h3fa0af57, 32'h3f88de2e} /* (31, 13, 12) {real, imag} */,
  {32'h3f101259, 32'h3ffb9515} /* (31, 13, 11) {real, imag} */,
  {32'hbfc7a384, 32'hbfe3f73f} /* (31, 13, 10) {real, imag} */,
  {32'h3fe6fe05, 32'hc01548fe} /* (31, 13, 9) {real, imag} */,
  {32'hbef6b690, 32'hbf5f7b52} /* (31, 13, 8) {real, imag} */,
  {32'h3e3c90cc, 32'hbf06602a} /* (31, 13, 7) {real, imag} */,
  {32'h3f1e9206, 32'hbf3bfbd2} /* (31, 13, 6) {real, imag} */,
  {32'hbfe14f29, 32'h40322daa} /* (31, 13, 5) {real, imag} */,
  {32'hc02ef729, 32'hbeb4365e} /* (31, 13, 4) {real, imag} */,
  {32'h3fa7fcde, 32'hbfcc9b00} /* (31, 13, 3) {real, imag} */,
  {32'hbda9de6a, 32'h3f794a6e} /* (31, 13, 2) {real, imag} */,
  {32'h402f5fe5, 32'h4030c423} /* (31, 13, 1) {real, imag} */,
  {32'hbff01b4e, 32'hbea75fae} /* (31, 13, 0) {real, imag} */,
  {32'h407382be, 32'h3fb82010} /* (31, 12, 31) {real, imag} */,
  {32'h3db1c527, 32'h3e849477} /* (31, 12, 30) {real, imag} */,
  {32'hbf8b32d2, 32'hbeceaf9c} /* (31, 12, 29) {real, imag} */,
  {32'hbf6263f8, 32'h3fc1f4bd} /* (31, 12, 28) {real, imag} */,
  {32'h3ec8c9c5, 32'h4040cb53} /* (31, 12, 27) {real, imag} */,
  {32'h3d704fc2, 32'hc070b2fa} /* (31, 12, 26) {real, imag} */,
  {32'h3e0b26df, 32'hbdbdd786} /* (31, 12, 25) {real, imag} */,
  {32'h3fa219bb, 32'hbfa9efa6} /* (31, 12, 24) {real, imag} */,
  {32'h3e3b45da, 32'hbfa5b396} /* (31, 12, 23) {real, imag} */,
  {32'h3ff2d38f, 32'hbf9156c1} /* (31, 12, 22) {real, imag} */,
  {32'h4023c2d9, 32'h402266fe} /* (31, 12, 21) {real, imag} */,
  {32'h3fedd6db, 32'h40229ff0} /* (31, 12, 20) {real, imag} */,
  {32'hbf8f6302, 32'hbf84dca6} /* (31, 12, 19) {real, imag} */,
  {32'hc022a534, 32'h3f616e5c} /* (31, 12, 18) {real, imag} */,
  {32'h3f6619c7, 32'h3fc8841b} /* (31, 12, 17) {real, imag} */,
  {32'hbe1362a6, 32'h3ff35833} /* (31, 12, 16) {real, imag} */,
  {32'h3e9fef79, 32'h3eab0d4c} /* (31, 12, 15) {real, imag} */,
  {32'hbf797fe9, 32'hbf580c88} /* (31, 12, 14) {real, imag} */,
  {32'h3f1bb97e, 32'hbf33e980} /* (31, 12, 13) {real, imag} */,
  {32'hbf2dd5ea, 32'h3fd902e8} /* (31, 12, 12) {real, imag} */,
  {32'h3d6a8969, 32'hbfb5874e} /* (31, 12, 11) {real, imag} */,
  {32'hbfb97606, 32'hc02f62e0} /* (31, 12, 10) {real, imag} */,
  {32'hbd69cbdf, 32'hbfb57a88} /* (31, 12, 9) {real, imag} */,
  {32'hbf9342e4, 32'h3fedecb5} /* (31, 12, 8) {real, imag} */,
  {32'hbf351fa4, 32'h3f81da52} /* (31, 12, 7) {real, imag} */,
  {32'h3ed34790, 32'h3f7da26e} /* (31, 12, 6) {real, imag} */,
  {32'h4004b40c, 32'hbdae78e1} /* (31, 12, 5) {real, imag} */,
  {32'hbefdcfd1, 32'h40101e32} /* (31, 12, 4) {real, imag} */,
  {32'h40190d68, 32'hbe8ad0d2} /* (31, 12, 3) {real, imag} */,
  {32'hbfeba609, 32'h3eb78c4f} /* (31, 12, 2) {real, imag} */,
  {32'h3fd6b639, 32'h3f37ee69} /* (31, 12, 1) {real, imag} */,
  {32'hc09d0661, 32'hc05715cd} /* (31, 12, 0) {real, imag} */,
  {32'h40a493c2, 32'hc0483920} /* (31, 11, 31) {real, imag} */,
  {32'hc034fd9d, 32'h3fefbf6d} /* (31, 11, 30) {real, imag} */,
  {32'hbfdc56ce, 32'hbf41a365} /* (31, 11, 29) {real, imag} */,
  {32'hbdee9fc7, 32'hbe368694} /* (31, 11, 28) {real, imag} */,
  {32'hc04cdea8, 32'h40488b06} /* (31, 11, 27) {real, imag} */,
  {32'hbf04b0fa, 32'h40a18fd0} /* (31, 11, 26) {real, imag} */,
  {32'h3f63b330, 32'h3d1f410a} /* (31, 11, 25) {real, imag} */,
  {32'h3f860255, 32'h40671f87} /* (31, 11, 24) {real, imag} */,
  {32'hbf86ec8d, 32'h3fa9ad8f} /* (31, 11, 23) {real, imag} */,
  {32'hbf2a2131, 32'h3fc9852b} /* (31, 11, 22) {real, imag} */,
  {32'hbeaafb00, 32'hbcdc6ca8} /* (31, 11, 21) {real, imag} */,
  {32'hbe84a8b7, 32'h3fcecd1f} /* (31, 11, 20) {real, imag} */,
  {32'h3e0d22ec, 32'hbef86db1} /* (31, 11, 19) {real, imag} */,
  {32'hc02e2546, 32'hbe4cec1e} /* (31, 11, 18) {real, imag} */,
  {32'h3f6dcaa7, 32'hbf711393} /* (31, 11, 17) {real, imag} */,
  {32'h3f54e978, 32'h3fd7e4fb} /* (31, 11, 16) {real, imag} */,
  {32'hbdc7c23f, 32'h3e198f9f} /* (31, 11, 15) {real, imag} */,
  {32'h3f73d978, 32'hbd10fd8f} /* (31, 11, 14) {real, imag} */,
  {32'hbf8eef61, 32'h3ebf1a05} /* (31, 11, 13) {real, imag} */,
  {32'h4066e3c7, 32'hc00935ff} /* (31, 11, 12) {real, imag} */,
  {32'h3f50bb0c, 32'h3d8b16ac} /* (31, 11, 11) {real, imag} */,
  {32'hbffcd3fa, 32'hbef088a4} /* (31, 11, 10) {real, imag} */,
  {32'h4021fbdc, 32'h3f5055c7} /* (31, 11, 9) {real, imag} */,
  {32'hbebe1c1a, 32'hbe9d3c00} /* (31, 11, 8) {real, imag} */,
  {32'h3f400336, 32'hbfe81d6b} /* (31, 11, 7) {real, imag} */,
  {32'hbea25769, 32'h4038d41f} /* (31, 11, 6) {real, imag} */,
  {32'hbf836dd4, 32'h3f20dc90} /* (31, 11, 5) {real, imag} */,
  {32'h4055d6d1, 32'h3ecf1599} /* (31, 11, 4) {real, imag} */,
  {32'h3f0aa5f2, 32'h3fbfb9d7} /* (31, 11, 3) {real, imag} */,
  {32'hc089599e, 32'h3f313a2a} /* (31, 11, 2) {real, imag} */,
  {32'h40bedc32, 32'hbfccc3ec} /* (31, 11, 1) {real, imag} */,
  {32'h406a26be, 32'hc0535263} /* (31, 11, 0) {real, imag} */,
  {32'hc05d0fb1, 32'h3e3dfefe} /* (31, 10, 31) {real, imag} */,
  {32'h408bde3d, 32'hbfa8c1db} /* (31, 10, 30) {real, imag} */,
  {32'hbe452f11, 32'h3fba2053} /* (31, 10, 29) {real, imag} */,
  {32'hbe3b261b, 32'h3f95466b} /* (31, 10, 28) {real, imag} */,
  {32'hbe2de58e, 32'hbe1b7526} /* (31, 10, 27) {real, imag} */,
  {32'h3e1555a5, 32'hbd39978e} /* (31, 10, 26) {real, imag} */,
  {32'hbf90c833, 32'hc031e12a} /* (31, 10, 25) {real, imag} */,
  {32'hc01802ec, 32'hbf8f1919} /* (31, 10, 24) {real, imag} */,
  {32'h3f28ff38, 32'hbf05ef27} /* (31, 10, 23) {real, imag} */,
  {32'hbfbdf5fc, 32'h3f067274} /* (31, 10, 22) {real, imag} */,
  {32'hbff9eabb, 32'hbf3816d6} /* (31, 10, 21) {real, imag} */,
  {32'hbeefda1f, 32'h4010059e} /* (31, 10, 20) {real, imag} */,
  {32'h3f04105b, 32'hbfac391a} /* (31, 10, 19) {real, imag} */,
  {32'h3fa8bbe4, 32'hbfddc73c} /* (31, 10, 18) {real, imag} */,
  {32'h3e779b25, 32'h3f3ff222} /* (31, 10, 17) {real, imag} */,
  {32'h3f3cf0ec, 32'hbec17661} /* (31, 10, 16) {real, imag} */,
  {32'h3f35b320, 32'h3e8ec475} /* (31, 10, 15) {real, imag} */,
  {32'h3fab335f, 32'hbe7d7e79} /* (31, 10, 14) {real, imag} */,
  {32'h3fa52b4c, 32'hbee5f5ee} /* (31, 10, 13) {real, imag} */,
  {32'h3f91022e, 32'h3e759bf4} /* (31, 10, 12) {real, imag} */,
  {32'hbef0eb05, 32'h3ed4e984} /* (31, 10, 11) {real, imag} */,
  {32'h3f19270c, 32'hbfb484d6} /* (31, 10, 10) {real, imag} */,
  {32'h3ee5c44c, 32'h406614ab} /* (31, 10, 9) {real, imag} */,
  {32'h3f069ad1, 32'hc0264a68} /* (31, 10, 8) {real, imag} */,
  {32'h3f92b86a, 32'hbeb08718} /* (31, 10, 7) {real, imag} */,
  {32'hbda456c8, 32'hbf6e1c7c} /* (31, 10, 6) {real, imag} */,
  {32'h3fd5ea44, 32'h4052bc3c} /* (31, 10, 5) {real, imag} */,
  {32'hbfc08022, 32'h401761ff} /* (31, 10, 4) {real, imag} */,
  {32'h3f7d441a, 32'h3f66f25a} /* (31, 10, 3) {real, imag} */,
  {32'h3ebab4e9, 32'h40460128} /* (31, 10, 2) {real, imag} */,
  {32'hc02f4fed, 32'h403a3ddf} /* (31, 10, 1) {real, imag} */,
  {32'hc04b00eb, 32'hc035e07c} /* (31, 10, 0) {real, imag} */,
  {32'hc036eeb4, 32'hc042bffc} /* (31, 9, 31) {real, imag} */,
  {32'h410c94f4, 32'h3fe34491} /* (31, 9, 30) {real, imag} */,
  {32'hc0af2c39, 32'hbf042b04} /* (31, 9, 29) {real, imag} */,
  {32'h4006569f, 32'h4032d870} /* (31, 9, 28) {real, imag} */,
  {32'h3b9f5322, 32'hbe4e7deb} /* (31, 9, 27) {real, imag} */,
  {32'h404f7ec0, 32'h4066db77} /* (31, 9, 26) {real, imag} */,
  {32'hbde78b33, 32'hbf9f11fe} /* (31, 9, 25) {real, imag} */,
  {32'hbf5538db, 32'hc0837560} /* (31, 9, 24) {real, imag} */,
  {32'h3ed15b5c, 32'hc04549fd} /* (31, 9, 23) {real, imag} */,
  {32'h3f6b771b, 32'h3f9fef8c} /* (31, 9, 22) {real, imag} */,
  {32'h4015d319, 32'hbf5c0df1} /* (31, 9, 21) {real, imag} */,
  {32'hc011f9e6, 32'hbf88c66e} /* (31, 9, 20) {real, imag} */,
  {32'hc03468c5, 32'h3e31d07e} /* (31, 9, 19) {real, imag} */,
  {32'h3feade6b, 32'h3fc3e7c2} /* (31, 9, 18) {real, imag} */,
  {32'hbfcbe414, 32'hc01323e9} /* (31, 9, 17) {real, imag} */,
  {32'h3fa36f1b, 32'h3c12efba} /* (31, 9, 16) {real, imag} */,
  {32'hc0203cf3, 32'hbfc6898d} /* (31, 9, 15) {real, imag} */,
  {32'hbfb15442, 32'h3f45b389} /* (31, 9, 14) {real, imag} */,
  {32'h3f9beece, 32'hbdafef2d} /* (31, 9, 13) {real, imag} */,
  {32'h40080c20, 32'h3ce14c5d} /* (31, 9, 12) {real, imag} */,
  {32'h3f626ab5, 32'hbf3919e5} /* (31, 9, 11) {real, imag} */,
  {32'h401ca27c, 32'hbda0535b} /* (31, 9, 10) {real, imag} */,
  {32'hc095a14c, 32'hc0008bb4} /* (31, 9, 9) {real, imag} */,
  {32'h403bf4e9, 32'hc05e7c3e} /* (31, 9, 8) {real, imag} */,
  {32'hbf850ade, 32'hc016490c} /* (31, 9, 7) {real, imag} */,
  {32'hbf51f932, 32'h3f8f0f40} /* (31, 9, 6) {real, imag} */,
  {32'h40937619, 32'hbfc52b0f} /* (31, 9, 5) {real, imag} */,
  {32'h404224fc, 32'hc01a7b20} /* (31, 9, 4) {real, imag} */,
  {32'hc0da4716, 32'h40959960} /* (31, 9, 3) {real, imag} */,
  {32'h4084a20a, 32'hc07a483d} /* (31, 9, 2) {real, imag} */,
  {32'hc0a50389, 32'h3fe12bc7} /* (31, 9, 1) {real, imag} */,
  {32'hc035798d, 32'hbf0ba218} /* (31, 9, 0) {real, imag} */,
  {32'h40f77750, 32'hc17d5cf5} /* (31, 8, 31) {real, imag} */,
  {32'hbf558af0, 32'h40c2d984} /* (31, 8, 30) {real, imag} */,
  {32'hbfd1c0e0, 32'hbefcf5f0} /* (31, 8, 29) {real, imag} */,
  {32'hc06afd8d, 32'h3ebee1e7} /* (31, 8, 28) {real, imag} */,
  {32'h3eeebc28, 32'h411b8949} /* (31, 8, 27) {real, imag} */,
  {32'hbc980722, 32'h3fecb148} /* (31, 8, 26) {real, imag} */,
  {32'hc007ec91, 32'hbd08c4b5} /* (31, 8, 25) {real, imag} */,
  {32'h3f2ec070, 32'h408017f8} /* (31, 8, 24) {real, imag} */,
  {32'h402324b4, 32'hbfaacd16} /* (31, 8, 23) {real, imag} */,
  {32'hbfc1453c, 32'hc043ea12} /* (31, 8, 22) {real, imag} */,
  {32'hbf24fe94, 32'hbf305a18} /* (31, 8, 21) {real, imag} */,
  {32'hbeaf9f0d, 32'hc008dc47} /* (31, 8, 20) {real, imag} */,
  {32'h3dce2417, 32'h3f2bb6f9} /* (31, 8, 19) {real, imag} */,
  {32'h3e608ecf, 32'h3fbd7cce} /* (31, 8, 18) {real, imag} */,
  {32'h4001ac78, 32'h3f59cd53} /* (31, 8, 17) {real, imag} */,
  {32'hc011db6a, 32'hbf50b664} /* (31, 8, 16) {real, imag} */,
  {32'h3f81926d, 32'h3ec3a324} /* (31, 8, 15) {real, imag} */,
  {32'hbf803946, 32'h3ef7b605} /* (31, 8, 14) {real, imag} */,
  {32'h3ff700bc, 32'hbfcecc69} /* (31, 8, 13) {real, imag} */,
  {32'hbfda68a7, 32'h3f9741be} /* (31, 8, 12) {real, imag} */,
  {32'hbffb15b0, 32'hbfb6159a} /* (31, 8, 11) {real, imag} */,
  {32'h401383f9, 32'h3eeeb6f8} /* (31, 8, 10) {real, imag} */,
  {32'hc0268734, 32'hbe2ea78f} /* (31, 8, 9) {real, imag} */,
  {32'hc01a5cfc, 32'h40301769} /* (31, 8, 8) {real, imag} */,
  {32'hc017e22d, 32'hc0831359} /* (31, 8, 7) {real, imag} */,
  {32'hc04c072f, 32'hbf0e3375} /* (31, 8, 6) {real, imag} */,
  {32'hbd98e0c1, 32'h4037683f} /* (31, 8, 5) {real, imag} */,
  {32'h407f7b55, 32'hc01de680} /* (31, 8, 4) {real, imag} */,
  {32'h3e94e96b, 32'h3f62f008} /* (31, 8, 3) {real, imag} */,
  {32'hbedd2a7a, 32'h413f2f4f} /* (31, 8, 2) {real, imag} */,
  {32'h409012a4, 32'hc124ce92} /* (31, 8, 1) {real, imag} */,
  {32'h3fffbc67, 32'hc060332b} /* (31, 8, 0) {real, imag} */,
  {32'hc0ab4394, 32'h41203d89} /* (31, 7, 31) {real, imag} */,
  {32'hc0080fce, 32'h405bfd5a} /* (31, 7, 30) {real, imag} */,
  {32'hc0137a9c, 32'hc05140fe} /* (31, 7, 29) {real, imag} */,
  {32'hc0424b77, 32'hc0747af2} /* (31, 7, 28) {real, imag} */,
  {32'h3eb273fb, 32'h3f52edd4} /* (31, 7, 27) {real, imag} */,
  {32'h403c520d, 32'h3fd370ab} /* (31, 7, 26) {real, imag} */,
  {32'h4012c406, 32'h4065e631} /* (31, 7, 25) {real, imag} */,
  {32'h4025c705, 32'hbff4c3bd} /* (31, 7, 24) {real, imag} */,
  {32'h3fa75486, 32'hc0a63d7e} /* (31, 7, 23) {real, imag} */,
  {32'hc0355e50, 32'h3dd94058} /* (31, 7, 22) {real, imag} */,
  {32'hc012f2d6, 32'h3fe528ed} /* (31, 7, 21) {real, imag} */,
  {32'h3e49120b, 32'h3f655fed} /* (31, 7, 20) {real, imag} */,
  {32'hbfe64dcf, 32'h3f6f94d1} /* (31, 7, 19) {real, imag} */,
  {32'h3ecf1fec, 32'h3fad74e2} /* (31, 7, 18) {real, imag} */,
  {32'hbfbf52db, 32'h3f55f455} /* (31, 7, 17) {real, imag} */,
  {32'hbfa603f2, 32'hbff2c167} /* (31, 7, 16) {real, imag} */,
  {32'h3fe334b9, 32'hbfab317c} /* (31, 7, 15) {real, imag} */,
  {32'h3f9100bf, 32'hc0059e95} /* (31, 7, 14) {real, imag} */,
  {32'hbf67930d, 32'h3e843c66} /* (31, 7, 13) {real, imag} */,
  {32'h3fcb3157, 32'hc0320b20} /* (31, 7, 12) {real, imag} */,
  {32'hbf8d8f81, 32'h403f7d9e} /* (31, 7, 11) {real, imag} */,
  {32'h3e8d7b52, 32'h408b38b0} /* (31, 7, 10) {real, imag} */,
  {32'h3f811bec, 32'h3fc4bcc0} /* (31, 7, 9) {real, imag} */,
  {32'h3fb15b5a, 32'h3fa52b02} /* (31, 7, 8) {real, imag} */,
  {32'hbf02dbd2, 32'h3f8daa93} /* (31, 7, 7) {real, imag} */,
  {32'h3fba4c78, 32'h4053653b} /* (31, 7, 6) {real, imag} */,
  {32'h3ff03f72, 32'h408d2d3a} /* (31, 7, 5) {real, imag} */,
  {32'hc0a3fc5c, 32'hc0bfb318} /* (31, 7, 4) {real, imag} */,
  {32'h3fa8c72e, 32'hc084a4db} /* (31, 7, 3) {real, imag} */,
  {32'h409433c2, 32'hbfecd3dd} /* (31, 7, 2) {real, imag} */,
  {32'hc0865ac8, 32'hc0b5f1bd} /* (31, 7, 1) {real, imag} */,
  {32'h3e033c9c, 32'hbf3c350a} /* (31, 7, 0) {real, imag} */,
  {32'hc02e5067, 32'h41095004} /* (31, 6, 31) {real, imag} */,
  {32'h3f33a0fe, 32'h40c54a3c} /* (31, 6, 30) {real, imag} */,
  {32'h40a5628d, 32'h40291bc8} /* (31, 6, 29) {real, imag} */,
  {32'h3f611383, 32'hc041d314} /* (31, 6, 28) {real, imag} */,
  {32'hbf5dfc92, 32'h402dbc61} /* (31, 6, 27) {real, imag} */,
  {32'h3cb29b46, 32'h405d5fd4} /* (31, 6, 26) {real, imag} */,
  {32'h4053a2da, 32'h4053606d} /* (31, 6, 25) {real, imag} */,
  {32'h3fa3ec49, 32'h3ff8f65f} /* (31, 6, 24) {real, imag} */,
  {32'hbfefbe55, 32'hbf8004d0} /* (31, 6, 23) {real, imag} */,
  {32'hbf2ec3b3, 32'h3fba202c} /* (31, 6, 22) {real, imag} */,
  {32'hbf542c75, 32'hbf1cda0f} /* (31, 6, 21) {real, imag} */,
  {32'hbe9479e9, 32'hbf85b5e9} /* (31, 6, 20) {real, imag} */,
  {32'hc07e97b6, 32'hbf8c37c4} /* (31, 6, 19) {real, imag} */,
  {32'h3f75d0cc, 32'h3fd7f082} /* (31, 6, 18) {real, imag} */,
  {32'hbecc838c, 32'hbf7999ed} /* (31, 6, 17) {real, imag} */,
  {32'h3fafc11b, 32'hc029d477} /* (31, 6, 16) {real, imag} */,
  {32'hbe605592, 32'hbe7d11d8} /* (31, 6, 15) {real, imag} */,
  {32'hbf730fde, 32'h3fd07ff5} /* (31, 6, 14) {real, imag} */,
  {32'hbf9f8af4, 32'h3f721ec0} /* (31, 6, 13) {real, imag} */,
  {32'hc026e127, 32'hbe9630f1} /* (31, 6, 12) {real, imag} */,
  {32'h3f34880e, 32'h3ff2110c} /* (31, 6, 11) {real, imag} */,
  {32'h40880b00, 32'h3fc0de55} /* (31, 6, 10) {real, imag} */,
  {32'h3fa8c8fa, 32'hc0020797} /* (31, 6, 9) {real, imag} */,
  {32'h40164ffd, 32'h3ff44446} /* (31, 6, 8) {real, imag} */,
  {32'h3f120f4c, 32'h40791f53} /* (31, 6, 7) {real, imag} */,
  {32'hc0c3b93f, 32'h402948fd} /* (31, 6, 6) {real, imag} */,
  {32'h40416002, 32'h4068641a} /* (31, 6, 5) {real, imag} */,
  {32'h4040c5e2, 32'hc07a7709} /* (31, 6, 4) {real, imag} */,
  {32'hc0c8e7f2, 32'hc0a5019b} /* (31, 6, 3) {real, imag} */,
  {32'hc03e7dfe, 32'hc113bc74} /* (31, 6, 2) {real, imag} */,
  {32'hc087e8dd, 32'h3f7b487c} /* (31, 6, 1) {real, imag} */,
  {32'h40079cb4, 32'hc01d0230} /* (31, 6, 0) {real, imag} */,
  {32'hc0d7eb7e, 32'hc209fd83} /* (31, 5, 31) {real, imag} */,
  {32'h40096907, 32'h40f4ab44} /* (31, 5, 30) {real, imag} */,
  {32'hc09bba7b, 32'hc1231e52} /* (31, 5, 29) {real, imag} */,
  {32'h3fc77e5d, 32'hc083d14c} /* (31, 5, 28) {real, imag} */,
  {32'hbfc9c2ad, 32'h402d131a} /* (31, 5, 27) {real, imag} */,
  {32'hbeb9ae1c, 32'hc04ac8c2} /* (31, 5, 26) {real, imag} */,
  {32'hc01607b3, 32'h3f8c333d} /* (31, 5, 25) {real, imag} */,
  {32'h40839c46, 32'h408521e5} /* (31, 5, 24) {real, imag} */,
  {32'hbf4e4e91, 32'hbfb49a44} /* (31, 5, 23) {real, imag} */,
  {32'h3f00bc85, 32'h3ea48cfa} /* (31, 5, 22) {real, imag} */,
  {32'hbee9e59a, 32'h3ffd3401} /* (31, 5, 21) {real, imag} */,
  {32'h3fe3c4f1, 32'hc058b754} /* (31, 5, 20) {real, imag} */,
  {32'h3edd3926, 32'hbf01fc3a} /* (31, 5, 19) {real, imag} */,
  {32'h3f18c3a2, 32'hbf8ffebb} /* (31, 5, 18) {real, imag} */,
  {32'hbfec6098, 32'hbb9fb68b} /* (31, 5, 17) {real, imag} */,
  {32'hbb1f4c75, 32'h3f0aa8da} /* (31, 5, 16) {real, imag} */,
  {32'h3d2fbc86, 32'h3e96f1f1} /* (31, 5, 15) {real, imag} */,
  {32'hbfaf1175, 32'hbfacdc48} /* (31, 5, 14) {real, imag} */,
  {32'h3edcbdcc, 32'h3fd8b700} /* (31, 5, 13) {real, imag} */,
  {32'hbfec6c1f, 32'h4043077e} /* (31, 5, 12) {real, imag} */,
  {32'hc0859cf4, 32'h3f95e244} /* (31, 5, 11) {real, imag} */,
  {32'hc0251677, 32'hbf08976c} /* (31, 5, 10) {real, imag} */,
  {32'hbfe1144a, 32'h404f1cc2} /* (31, 5, 9) {real, imag} */,
  {32'hc00cbfa6, 32'hbfd4ce88} /* (31, 5, 8) {real, imag} */,
  {32'h3f81447a, 32'hc0c2487e} /* (31, 5, 7) {real, imag} */,
  {32'hbfc9a6d9, 32'hbad4afe7} /* (31, 5, 6) {real, imag} */,
  {32'hc02d4540, 32'h3fe3e8c9} /* (31, 5, 5) {real, imag} */,
  {32'h4078abcb, 32'hbf247139} /* (31, 5, 4) {real, imag} */,
  {32'hc09b04c9, 32'hc096f027} /* (31, 5, 3) {real, imag} */,
  {32'hc149838f, 32'h412e51e9} /* (31, 5, 2) {real, imag} */,
  {32'h41b323c8, 32'hc1694fe3} /* (31, 5, 1) {real, imag} */,
  {32'h4185105b, 32'hc1935b84} /* (31, 5, 0) {real, imag} */,
  {32'hc1ffdd89, 32'h419af120} /* (31, 4, 31) {real, imag} */,
  {32'h41962fc0, 32'hc198500d} /* (31, 4, 30) {real, imag} */,
  {32'hbf7ec318, 32'h40ce076f} /* (31, 4, 29) {real, imag} */,
  {32'hbf941fb1, 32'h4110a117} /* (31, 4, 28) {real, imag} */,
  {32'hc04a9d28, 32'hc033df8d} /* (31, 4, 27) {real, imag} */,
  {32'h3eaed6ac, 32'hc088a1b8} /* (31, 4, 26) {real, imag} */,
  {32'hbf449144, 32'hc013b834} /* (31, 4, 25) {real, imag} */,
  {32'hbed370e1, 32'hc04699dc} /* (31, 4, 24) {real, imag} */,
  {32'hbfbde391, 32'h404c37b0} /* (31, 4, 23) {real, imag} */,
  {32'h4053fbf8, 32'hbf236671} /* (31, 4, 22) {real, imag} */,
  {32'h4038f6a4, 32'h3fc26fbb} /* (31, 4, 21) {real, imag} */,
  {32'hbf83541f, 32'h3e79f3df} /* (31, 4, 20) {real, imag} */,
  {32'hbe74f736, 32'h3d95eefc} /* (31, 4, 19) {real, imag} */,
  {32'h3f423fa8, 32'hbfa52da9} /* (31, 4, 18) {real, imag} */,
  {32'h3f63682b, 32'hbdeb48e5} /* (31, 4, 17) {real, imag} */,
  {32'hbd311964, 32'h3e9a6b5c} /* (31, 4, 16) {real, imag} */,
  {32'hbffd382e, 32'hbe076b7d} /* (31, 4, 15) {real, imag} */,
  {32'h4009636c, 32'h4043b2ba} /* (31, 4, 14) {real, imag} */,
  {32'h3fc18595, 32'hbf676f87} /* (31, 4, 13) {real, imag} */,
  {32'hc04adafa, 32'hbfd3cb34} /* (31, 4, 12) {real, imag} */,
  {32'h409ee958, 32'h40573855} /* (31, 4, 11) {real, imag} */,
  {32'hbf4cdf4c, 32'hbf0d5328} /* (31, 4, 10) {real, imag} */,
  {32'hbd2faf67, 32'h3f6259d6} /* (31, 4, 9) {real, imag} */,
  {32'h40334fcb, 32'h3e91bf1f} /* (31, 4, 8) {real, imag} */,
  {32'h4028620d, 32'h406a9dd5} /* (31, 4, 7) {real, imag} */,
  {32'h408835b6, 32'h404c9d00} /* (31, 4, 6) {real, imag} */,
  {32'h412cd2c8, 32'hc05fd2a8} /* (31, 4, 5) {real, imag} */,
  {32'hc14baf62, 32'hc0bf47f6} /* (31, 4, 4) {real, imag} */,
  {32'hc0f1dc53, 32'h3d2c52e7} /* (31, 4, 3) {real, imag} */,
  {32'h416296ad, 32'hc1e646ec} /* (31, 4, 2) {real, imag} */,
  {32'hc1a40cb3, 32'h424b03c4} /* (31, 4, 1) {real, imag} */,
  {32'h41591b99, 32'h41c60966} /* (31, 4, 0) {real, imag} */,
  {32'hc1dcd3c0, 32'hc1e98d21} /* (31, 3, 31) {real, imag} */,
  {32'h4232533d, 32'h3ea2e905} /* (31, 3, 30) {real, imag} */,
  {32'h40b5caa4, 32'hc0271096} /* (31, 3, 29) {real, imag} */,
  {32'hc0fbe03a, 32'h41649e61} /* (31, 3, 28) {real, imag} */,
  {32'hbf7a25c9, 32'hc12c52a2} /* (31, 3, 27) {real, imag} */,
  {32'hbf2a284e, 32'hc0169c76} /* (31, 3, 26) {real, imag} */,
  {32'hbfe349ad, 32'hbf9b4af4} /* (31, 3, 25) {real, imag} */,
  {32'h3f7be866, 32'h40863b2b} /* (31, 3, 24) {real, imag} */,
  {32'h3fd15431, 32'hbf6ba67a} /* (31, 3, 23) {real, imag} */,
  {32'h4039d039, 32'h4034e648} /* (31, 3, 22) {real, imag} */,
  {32'hbf9c2d66, 32'h3e89aaad} /* (31, 3, 21) {real, imag} */,
  {32'hc006d944, 32'h3de46237} /* (31, 3, 20) {real, imag} */,
  {32'hbf2340ad, 32'h40076875} /* (31, 3, 19) {real, imag} */,
  {32'h3f5252d7, 32'hc006bde9} /* (31, 3, 18) {real, imag} */,
  {32'hbdd3a65f, 32'hbe82cdb3} /* (31, 3, 17) {real, imag} */,
  {32'hbf0b18cc, 32'hc00b49d0} /* (31, 3, 16) {real, imag} */,
  {32'hbe9736fd, 32'hbf72194d} /* (31, 3, 15) {real, imag} */,
  {32'h3ffac8d9, 32'h40a8032a} /* (31, 3, 14) {real, imag} */,
  {32'hbeae5878, 32'hbedbc459} /* (31, 3, 13) {real, imag} */,
  {32'h3f7821e0, 32'h3e82d4c7} /* (31, 3, 12) {real, imag} */,
  {32'hbf359e7c, 32'hbfe4a69f} /* (31, 3, 11) {real, imag} */,
  {32'hbf6d8af1, 32'hc00f2aee} /* (31, 3, 10) {real, imag} */,
  {32'h40449654, 32'h407082b6} /* (31, 3, 9) {real, imag} */,
  {32'hc00adf51, 32'h3fb08c70} /* (31, 3, 8) {real, imag} */,
  {32'h40512162, 32'hc027c274} /* (31, 3, 7) {real, imag} */,
  {32'hc04fd972, 32'hbf03e6bd} /* (31, 3, 6) {real, imag} */,
  {32'hc0c8180d, 32'h3ff635ec} /* (31, 3, 5) {real, imag} */,
  {32'hc0824e77, 32'hc11d1293} /* (31, 3, 4) {real, imag} */,
  {32'hc0afe47e, 32'hc1499d63} /* (31, 3, 3) {real, imag} */,
  {32'h41991450, 32'h3eb04014} /* (31, 3, 2) {real, imag} */,
  {32'hc1fd1b4e, 32'h427592a6} /* (31, 3, 1) {real, imag} */,
  {32'h4090b3f6, 32'hc14b4f84} /* (31, 3, 0) {real, imag} */,
  {32'hc1d1658e, 32'hc3be0ad6} /* (31, 2, 31) {real, imag} */,
  {32'h42967d5a, 32'h432231dd} /* (31, 2, 30) {real, imag} */,
  {32'hc1b2542c, 32'hc1032ab9} /* (31, 2, 29) {real, imag} */,
  {32'hc19bc397, 32'hc021b15a} /* (31, 2, 28) {real, imag} */,
  {32'h41248f9c, 32'h418cce9a} /* (31, 2, 27) {real, imag} */,
  {32'h4066d6b6, 32'h40842024} /* (31, 2, 26) {real, imag} */,
  {32'h3faa2123, 32'h3f9e8617} /* (31, 2, 25) {real, imag} */,
  {32'h40d7a494, 32'h41013c1b} /* (31, 2, 24) {real, imag} */,
  {32'h3ed092ea, 32'hc0962649} /* (31, 2, 23) {real, imag} */,
  {32'hbe41a295, 32'hbf745af2} /* (31, 2, 22) {real, imag} */,
  {32'h3f074bd4, 32'hbfa03e0e} /* (31, 2, 21) {real, imag} */,
  {32'h3ed309c2, 32'h400e74a5} /* (31, 2, 20) {real, imag} */,
  {32'h40125f90, 32'hbf9ba7e8} /* (31, 2, 19) {real, imag} */,
  {32'h4006ab3e, 32'hbf2c8dd2} /* (31, 2, 18) {real, imag} */,
  {32'h3e4ca095, 32'h3f8a50e5} /* (31, 2, 17) {real, imag} */,
  {32'h3f46cfb2, 32'h3f59ea01} /* (31, 2, 16) {real, imag} */,
  {32'h3f22aa12, 32'hbf7b38cc} /* (31, 2, 15) {real, imag} */,
  {32'hbe4ceadd, 32'hbed984e4} /* (31, 2, 14) {real, imag} */,
  {32'hbe921cb7, 32'hc013b4f0} /* (31, 2, 13) {real, imag} */,
  {32'h3e2d14dd, 32'h3f6a9b87} /* (31, 2, 12) {real, imag} */,
  {32'hc08e23c1, 32'h401c2de0} /* (31, 2, 11) {real, imag} */,
  {32'h3f72c956, 32'hbfec808d} /* (31, 2, 10) {real, imag} */,
  {32'hbf300945, 32'hbf1966f0} /* (31, 2, 9) {real, imag} */,
  {32'hc0c4a3b8, 32'h411381e9} /* (31, 2, 8) {real, imag} */,
  {32'h409c2598, 32'hc059de92} /* (31, 2, 7) {real, imag} */,
  {32'hc00efc93, 32'hc03166a0} /* (31, 2, 6) {real, imag} */,
  {32'hc138aa0b, 32'h41a988e3} /* (31, 2, 5) {real, imag} */,
  {32'h40997199, 32'hc191f598} /* (31, 2, 4) {real, imag} */,
  {32'hc1b29041, 32'hc0c0787d} /* (31, 2, 3) {real, imag} */,
  {32'h4214d5ee, 32'h42f14415} /* (31, 2, 2) {real, imag} */,
  {32'hc28ed767, 32'hc33e6304} /* (31, 2, 1) {real, imag} */,
  {32'h41042068, 32'hc3624196} /* (31, 2, 0) {real, imag} */,
  {32'h4344c965, 32'h4407fd22} /* (31, 1, 31) {real, imag} */,
  {32'hc11b89ec, 32'hc2e5de86} /* (31, 1, 30) {real, imag} */,
  {32'h409e9d0a, 32'hc0f53094} /* (31, 1, 29) {real, imag} */,
  {32'hc19fbc62, 32'h420de9c4} /* (31, 1, 28) {real, imag} */,
  {32'hc075fc07, 32'hc1ea5854} /* (31, 1, 27) {real, imag} */,
  {32'hc124507e, 32'h400cf5e9} /* (31, 1, 26) {real, imag} */,
  {32'h3f2b8969, 32'hc080824f} /* (31, 1, 25) {real, imag} */,
  {32'h3dd47b1f, 32'hc0924b6c} /* (31, 1, 24) {real, imag} */,
  {32'hbf5fd1f8, 32'hc052c65b} /* (31, 1, 23) {real, imag} */,
  {32'hc0ca7963, 32'hbdd5e25f} /* (31, 1, 22) {real, imag} */,
  {32'hc0569840, 32'hc0b538bc} /* (31, 1, 21) {real, imag} */,
  {32'h402fa83a, 32'h4009ea39} /* (31, 1, 20) {real, imag} */,
  {32'hbf8a6cf8, 32'hbfebc496} /* (31, 1, 19) {real, imag} */,
  {32'hc09b8aef, 32'hc02bf1ce} /* (31, 1, 18) {real, imag} */,
  {32'hbe2dce92, 32'hbeb0c51c} /* (31, 1, 17) {real, imag} */,
  {32'hbfb0b248, 32'h3e97b39a} /* (31, 1, 16) {real, imag} */,
  {32'hbf694cc0, 32'h3f5228da} /* (31, 1, 15) {real, imag} */,
  {32'h400b8735, 32'hbff3a28a} /* (31, 1, 14) {real, imag} */,
  {32'h3f567d6d, 32'h3f0f7361} /* (31, 1, 13) {real, imag} */,
  {32'h40644c9e, 32'h3fdf108e} /* (31, 1, 12) {real, imag} */,
  {32'h40c7ea4c, 32'hc0658ced} /* (31, 1, 11) {real, imag} */,
  {32'h3f890c71, 32'hbcf948e1} /* (31, 1, 10) {real, imag} */,
  {32'hc079e560, 32'hbffce1a2} /* (31, 1, 9) {real, imag} */,
  {32'h411ba76c, 32'hc0e0464c} /* (31, 1, 8) {real, imag} */,
  {32'hc0f30270, 32'h4109ff6e} /* (31, 1, 7) {real, imag} */,
  {32'h4033a287, 32'hc0563815} /* (31, 1, 6) {real, imag} */,
  {32'h40b8e41b, 32'hc1bde69e} /* (31, 1, 5) {real, imag} */,
  {32'h40710768, 32'h40b73d3c} /* (31, 1, 4) {real, imag} */,
  {32'h4199b3d9, 32'hc11cdff7} /* (31, 1, 3) {real, imag} */,
  {32'h431af7b3, 32'hc3604a4c} /* (31, 1, 2) {real, imag} */,
  {32'hc3aa13d4, 32'h444b82a2} /* (31, 1, 1) {real, imag} */,
  {32'hc1c9a61e, 32'h44599db9} /* (31, 1, 0) {real, imag} */,
  {32'h43f8eeaf, 32'h43f2ee9e} /* (31, 0, 31) {real, imag} */,
  {32'hc2c83a22, 32'hc1b9a883} /* (31, 0, 30) {real, imag} */,
  {32'h40b9f1d8, 32'hc10688cd} /* (31, 0, 29) {real, imag} */,
  {32'hc10f78d7, 32'hc134bfd9} /* (31, 0, 28) {real, imag} */,
  {32'h3eb178f7, 32'hc1b2c9b5} /* (31, 0, 27) {real, imag} */,
  {32'hbe569a77, 32'h40900d4c} /* (31, 0, 26) {real, imag} */,
  {32'hbe5e227a, 32'hbf6ba998} /* (31, 0, 25) {real, imag} */,
  {32'hc122d2b2, 32'hbf5f2e60} /* (31, 0, 24) {real, imag} */,
  {32'hbfb50995, 32'hbd9071fb} /* (31, 0, 23) {real, imag} */,
  {32'h3ef0d534, 32'h3f4db9d7} /* (31, 0, 22) {real, imag} */,
  {32'hbf40ada2, 32'hc00bc104} /* (31, 0, 21) {real, imag} */,
  {32'hbfaf02d5, 32'h3eed8bee} /* (31, 0, 20) {real, imag} */,
  {32'h3eba03a0, 32'h3f9207e4} /* (31, 0, 19) {real, imag} */,
  {32'hbf9c77e3, 32'hbfab8ca8} /* (31, 0, 18) {real, imag} */,
  {32'h3f7c92f4, 32'hc018ee15} /* (31, 0, 17) {real, imag} */,
  {32'hbf1bb697, 32'hc02b344d} /* (31, 0, 16) {real, imag} */,
  {32'hbed34cd7, 32'hbc1599da} /* (31, 0, 15) {real, imag} */,
  {32'h40829427, 32'hbec200ee} /* (31, 0, 14) {real, imag} */,
  {32'hbf05cd0b, 32'h3fc0526f} /* (31, 0, 13) {real, imag} */,
  {32'hbf8195f2, 32'h3f41d5af} /* (31, 0, 12) {real, imag} */,
  {32'h3e720b74, 32'hc0afa305} /* (31, 0, 11) {real, imag} */,
  {32'h40542e0e, 32'hc0163344} /* (31, 0, 10) {real, imag} */,
  {32'h3f56a504, 32'h3eaf3d27} /* (31, 0, 9) {real, imag} */,
  {32'h4086b665, 32'h40009ca8} /* (31, 0, 8) {real, imag} */,
  {32'hc0a4ec6a, 32'hbf407311} /* (31, 0, 7) {real, imag} */,
  {32'h40282af0, 32'hbf1f976d} /* (31, 0, 6) {real, imag} */,
  {32'h40766113, 32'hc1647cd2} /* (31, 0, 5) {real, imag} */,
  {32'h4119f0b6, 32'hc0984cf1} /* (31, 0, 4) {real, imag} */,
  {32'h40e92c10, 32'h40b1590d} /* (31, 0, 3) {real, imag} */,
  {32'h42a5062c, 32'hc2aaf1e8} /* (31, 0, 2) {real, imag} */,
  {32'hc3b5ba3a, 32'h441220bc} /* (31, 0, 1) {real, imag} */,
  {32'h42ad3089, 32'h4470e74f} /* (31, 0, 0) {real, imag} */,
  {32'hc4101db2, 32'hc4259730} /* (30, 31, 31) {real, imag} */,
  {32'h438094da, 32'h43321858} /* (30, 31, 30) {real, imag} */,
  {32'hc15e74e7, 32'h415d584f} /* (30, 31, 29) {real, imag} */,
  {32'hc1f3bc94, 32'hc171ecc8} /* (30, 31, 28) {real, imag} */,
  {32'h41deaa82, 32'h41ed0171} /* (30, 31, 27) {real, imag} */,
  {32'h40b49222, 32'h3f0ef6cc} /* (30, 31, 26) {real, imag} */,
  {32'hc10a7bb7, 32'hc0660183} /* (30, 31, 25) {real, imag} */,
  {32'h4195e005, 32'h40258639} /* (30, 31, 24) {real, imag} */,
  {32'h3e8c5ffe, 32'hbf251469} /* (30, 31, 23) {real, imag} */,
  {32'h40972715, 32'h405577cd} /* (30, 31, 22) {real, imag} */,
  {32'h40d4e124, 32'h3f2db7d1} /* (30, 31, 21) {real, imag} */,
  {32'h4023af26, 32'hbdb2de06} /* (30, 31, 20) {real, imag} */,
  {32'hbffeae5d, 32'hc092e7f4} /* (30, 31, 19) {real, imag} */,
  {32'h4089e5d6, 32'hc02b9ee3} /* (30, 31, 18) {real, imag} */,
  {32'hbec74663, 32'h3fb32487} /* (30, 31, 17) {real, imag} */,
  {32'hbf83b9c4, 32'h3c452f02} /* (30, 31, 16) {real, imag} */,
  {32'hbc8e9d8b, 32'h3eb72f54} /* (30, 31, 15) {real, imag} */,
  {32'hc07d6086, 32'h3cee3d61} /* (30, 31, 14) {real, imag} */,
  {32'hbf8d1f42, 32'hbfe3a8a2} /* (30, 31, 13) {real, imag} */,
  {32'hbf91004d, 32'hbe975261} /* (30, 31, 12) {real, imag} */,
  {32'hc01b7283, 32'h4128e89c} /* (30, 31, 11) {real, imag} */,
  {32'hc076eec8, 32'hc03ea4ce} /* (30, 31, 10) {real, imag} */,
  {32'hc0d06433, 32'h40a1773a} /* (30, 31, 9) {real, imag} */,
  {32'hc0a7e4eb, 32'h40f9ef3a} /* (30, 31, 8) {real, imag} */,
  {32'h40393b16, 32'hc0fa62ca} /* (30, 31, 7) {real, imag} */,
  {32'h40cd96a8, 32'h412d74c5} /* (30, 31, 6) {real, imag} */,
  {32'h4140e774, 32'h424ccf86} /* (30, 31, 5) {real, imag} */,
  {32'hc1ef9c2f, 32'hc1a61ab4} /* (30, 31, 4) {real, imag} */,
  {32'hc18b5e36, 32'hbef0691d} /* (30, 31, 3) {real, imag} */,
  {32'h4182779c, 32'h433b15b1} /* (30, 31, 2) {real, imag} */,
  {32'h41c4e950, 32'hc4068a5c} /* (30, 31, 1) {real, imag} */,
  {32'hc3392074, 32'hc40d4f55} /* (30, 31, 0) {real, imag} */,
  {32'hc06c0445, 32'h438e9193} /* (30, 30, 31) {real, imag} */,
  {32'h41508195, 32'hc3389c33} /* (30, 30, 30) {real, imag} */,
  {32'h40a3258e, 32'h408fdef4} /* (30, 30, 29) {real, imag} */,
  {32'h420753db, 32'h4240b24b} /* (30, 30, 28) {real, imag} */,
  {32'hc20a4c56, 32'hc1863c08} /* (30, 30, 27) {real, imag} */,
  {32'hbfe854dd, 32'hc08d9de9} /* (30, 30, 26) {real, imag} */,
  {32'h3f1c0eb5, 32'h4082a530} /* (30, 30, 25) {real, imag} */,
  {32'hc0f6d6f1, 32'hc0bf46f4} /* (30, 30, 24) {real, imag} */,
  {32'hbf71539b, 32'h402f79f4} /* (30, 30, 23) {real, imag} */,
  {32'h4001e860, 32'h4080d7d0} /* (30, 30, 22) {real, imag} */,
  {32'hc0f430c6, 32'hbff0ecf6} /* (30, 30, 21) {real, imag} */,
  {32'h3f2b1183, 32'hbf54a96f} /* (30, 30, 20) {real, imag} */,
  {32'h3e850304, 32'hbd7b589b} /* (30, 30, 19) {real, imag} */,
  {32'hc07e05c3, 32'hbf055f9c} /* (30, 30, 18) {real, imag} */,
  {32'hbeb622ac, 32'h4029f31c} /* (30, 30, 17) {real, imag} */,
  {32'h3f027bee, 32'h3f9f59a4} /* (30, 30, 16) {real, imag} */,
  {32'hc02a7867, 32'hbd21f263} /* (30, 30, 15) {real, imag} */,
  {32'h404b2c9a, 32'hc03714ee} /* (30, 30, 14) {real, imag} */,
  {32'hbfa333ba, 32'hbe5b3062} /* (30, 30, 13) {real, imag} */,
  {32'hc02f2d66, 32'h4044eadf} /* (30, 30, 12) {real, imag} */,
  {32'h40d793ef, 32'hc0cf1038} /* (30, 30, 11) {real, imag} */,
  {32'hbfb2b7f5, 32'hbe2f4c53} /* (30, 30, 10) {real, imag} */,
  {32'hc0629fca, 32'hc01dc65f} /* (30, 30, 9) {real, imag} */,
  {32'h411c647d, 32'hc0f24b1f} /* (30, 30, 8) {real, imag} */,
  {32'hc123b7aa, 32'h413e340a} /* (30, 30, 7) {real, imag} */,
  {32'h400fa093, 32'hc106bdf4} /* (30, 30, 6) {real, imag} */,
  {32'h4115c006, 32'hc21209b1} /* (30, 30, 5) {real, imag} */,
  {32'hc2144f00, 32'h419ebd67} /* (30, 30, 4) {real, imag} */,
  {32'h413993e9, 32'h402f159a} /* (30, 30, 3) {real, imag} */,
  {32'h41b0175f, 32'hc3675454} /* (30, 30, 2) {real, imag} */,
  {32'h42e44b9b, 32'h43e66b07} /* (30, 30, 1) {real, imag} */,
  {32'h42a9df32, 32'h434c8af2} /* (30, 30, 0) {real, imag} */,
  {32'hc236ad6f, 32'hc1ec813b} /* (30, 29, 31) {real, imag} */,
  {32'h4267b321, 32'hbf6fec37} /* (30, 29, 30) {real, imag} */,
  {32'hbfe61e01, 32'h40f037cf} /* (30, 29, 29) {real, imag} */,
  {32'hc0022452, 32'h404c88ea} /* (30, 29, 28) {real, imag} */,
  {32'hc0ee4e4f, 32'hc128e4bb} /* (30, 29, 27) {real, imag} */,
  {32'hc06a24fb, 32'h40ab177a} /* (30, 29, 26) {real, imag} */,
  {32'hc0071bfc, 32'hc01f9fa9} /* (30, 29, 25) {real, imag} */,
  {32'h40b0cbef, 32'h3f668333} /* (30, 29, 24) {real, imag} */,
  {32'hbfae8848, 32'h401bd7e2} /* (30, 29, 23) {real, imag} */,
  {32'h4025c4f6, 32'h408c9c69} /* (30, 29, 22) {real, imag} */,
  {32'hbfe1a2cc, 32'hc091394e} /* (30, 29, 21) {real, imag} */,
  {32'h3f3c8752, 32'hbf0ee040} /* (30, 29, 20) {real, imag} */,
  {32'h3fa44cbe, 32'hbf24fe37} /* (30, 29, 19) {real, imag} */,
  {32'h403c6233, 32'hbf0d8472} /* (30, 29, 18) {real, imag} */,
  {32'h3e95bfb2, 32'h3e0f53a6} /* (30, 29, 17) {real, imag} */,
  {32'hc00e7b81, 32'hbe2a1814} /* (30, 29, 16) {real, imag} */,
  {32'hbd35b7e3, 32'h3f2cd7fc} /* (30, 29, 15) {real, imag} */,
  {32'hbea1592c, 32'hbe2f88b1} /* (30, 29, 14) {real, imag} */,
  {32'hbeb58590, 32'h4003fffc} /* (30, 29, 13) {real, imag} */,
  {32'hbf3c9cc2, 32'h3f177697} /* (30, 29, 12) {real, imag} */,
  {32'hbfc7d9f5, 32'h406de4f2} /* (30, 29, 11) {real, imag} */,
  {32'hc0a91d20, 32'hc01148db} /* (30, 29, 10) {real, imag} */,
  {32'hc0aadeca, 32'hc00b87e7} /* (30, 29, 9) {real, imag} */,
  {32'h40aba62d, 32'hbdb8d9c4} /* (30, 29, 8) {real, imag} */,
  {32'hbdf0c3e7, 32'hc0a249d9} /* (30, 29, 7) {real, imag} */,
  {32'hc096839a, 32'hbf5ae6e3} /* (30, 29, 6) {real, imag} */,
  {32'h40222ddc, 32'h413a6e7c} /* (30, 29, 5) {real, imag} */,
  {32'hc168e66a, 32'hc177c4a0} /* (30, 29, 4) {real, imag} */,
  {32'hc0b1d76b, 32'h3ed3156f} /* (30, 29, 3) {real, imag} */,
  {32'h4231fed4, 32'hc2705097} /* (30, 29, 2) {real, imag} */,
  {32'hc1882d18, 32'h4286fa98} /* (30, 29, 1) {real, imag} */,
  {32'hc0d00007, 32'h40591057} /* (30, 29, 0) {real, imag} */,
  {32'hc2029c05, 32'hc28c1420} /* (30, 28, 31) {real, imag} */,
  {32'h4223e130, 32'h41e534a5} /* (30, 28, 30) {real, imag} */,
  {32'hc01e7dd8, 32'hc0d147ee} /* (30, 28, 29) {real, imag} */,
  {32'hc13891ad, 32'hc0c41e17} /* (30, 28, 28) {real, imag} */,
  {32'h40f80ab1, 32'hc02964dd} /* (30, 28, 27) {real, imag} */,
  {32'h3e138acb, 32'h402ea893} /* (30, 28, 26) {real, imag} */,
  {32'hbea03c27, 32'hc05d341d} /* (30, 28, 25) {real, imag} */,
  {32'h40bdeeae, 32'hbe113cdc} /* (30, 28, 24) {real, imag} */,
  {32'h3f8da545, 32'hbecb32f8} /* (30, 28, 23) {real, imag} */,
  {32'hc026b2c3, 32'h3fde8d7e} /* (30, 28, 22) {real, imag} */,
  {32'hbdf5a8a0, 32'h3e33810d} /* (30, 28, 21) {real, imag} */,
  {32'h40780b6c, 32'h4002b7bc} /* (30, 28, 20) {real, imag} */,
  {32'h3e8edc62, 32'hbfce630c} /* (30, 28, 19) {real, imag} */,
  {32'h3ff2fbc1, 32'hbe3c0b9e} /* (30, 28, 18) {real, imag} */,
  {32'h3f8217db, 32'h3fbee9ee} /* (30, 28, 17) {real, imag} */,
  {32'h3f61ed2b, 32'h3f6bc1da} /* (30, 28, 16) {real, imag} */,
  {32'hc032094c, 32'hbeab797b} /* (30, 28, 15) {real, imag} */,
  {32'h3f199c76, 32'h3f0d89cf} /* (30, 28, 14) {real, imag} */,
  {32'h3ce79ce5, 32'h3dbfd9d3} /* (30, 28, 13) {real, imag} */,
  {32'h3fea8b98, 32'h3f08cd6d} /* (30, 28, 12) {real, imag} */,
  {32'hc057ea9f, 32'h40e54ae2} /* (30, 28, 11) {real, imag} */,
  {32'h3fc5ff71, 32'hc0763dec} /* (30, 28, 10) {real, imag} */,
  {32'hc0436d89, 32'hc02f2b8f} /* (30, 28, 9) {real, imag} */,
  {32'hbe74efa5, 32'h409558ab} /* (30, 28, 8) {real, imag} */,
  {32'hc02834fd, 32'hbe561384} /* (30, 28, 7) {real, imag} */,
  {32'hc0b1319c, 32'hc063b132} /* (30, 28, 6) {real, imag} */,
  {32'hc0437c1f, 32'h4103c120} /* (30, 28, 5) {real, imag} */,
  {32'hc08bf3ec, 32'hc186f7d9} /* (30, 28, 4) {real, imag} */,
  {32'h3f0dc41a, 32'h3fca41d4} /* (30, 28, 3) {real, imag} */,
  {32'h42056b8e, 32'h41d47a65} /* (30, 28, 2) {real, imag} */,
  {32'hc22100bd, 32'hc158cb75} /* (30, 28, 1) {real, imag} */,
  {32'hc0e6cae1, 32'hc164deb8} /* (30, 28, 0) {real, imag} */,
  {32'h41e55b7c, 32'h41d6dbc5} /* (30, 27, 31) {real, imag} */,
  {32'hc1032788, 32'hc066c6c3} /* (30, 27, 30) {real, imag} */,
  {32'h407f3888, 32'h3fbd380d} /* (30, 27, 29) {real, imag} */,
  {32'h40d0eb07, 32'h409d4fcb} /* (30, 27, 28) {real, imag} */,
  {32'hc178083c, 32'hc1528df3} /* (30, 27, 27) {real, imag} */,
  {32'hc04d3532, 32'h4087f054} /* (30, 27, 26) {real, imag} */,
  {32'h401d0abf, 32'hbe1539b8} /* (30, 27, 25) {real, imag} */,
  {32'hc09eda4b, 32'hc03a9c8b} /* (30, 27, 24) {real, imag} */,
  {32'h3f38bee6, 32'hc008e1d3} /* (30, 27, 23) {real, imag} */,
  {32'hbe846cea, 32'h4042ae19} /* (30, 27, 22) {real, imag} */,
  {32'hc09a86b1, 32'hbf6f4cd9} /* (30, 27, 21) {real, imag} */,
  {32'hbfc6e97a, 32'hc0395d3a} /* (30, 27, 20) {real, imag} */,
  {32'h3fa781d6, 32'h3f916e84} /* (30, 27, 19) {real, imag} */,
  {32'hbfa2d2ee, 32'h400c3b95} /* (30, 27, 18) {real, imag} */,
  {32'hbfc1c7bd, 32'h3fbd16c8} /* (30, 27, 17) {real, imag} */,
  {32'h3ece6f24, 32'hbe83ad69} /* (30, 27, 16) {real, imag} */,
  {32'h4004d570, 32'hbed95fef} /* (30, 27, 15) {real, imag} */,
  {32'h4030b8aa, 32'hc01527bd} /* (30, 27, 14) {real, imag} */,
  {32'hbfd83f11, 32'h3f04cc68} /* (30, 27, 13) {real, imag} */,
  {32'hbfb33d31, 32'hbdfcf8d0} /* (30, 27, 12) {real, imag} */,
  {32'h3f728b52, 32'hc0cd0e8d} /* (30, 27, 11) {real, imag} */,
  {32'h3fbe7311, 32'hc0575d63} /* (30, 27, 10) {real, imag} */,
  {32'hc0044ac7, 32'h3f1fd613} /* (30, 27, 9) {real, imag} */,
  {32'h40062f23, 32'hc08db10c} /* (30, 27, 8) {real, imag} */,
  {32'hbfaabacc, 32'h3decf768} /* (30, 27, 7) {real, imag} */,
  {32'h4023dbed, 32'hbfa1c822} /* (30, 27, 6) {real, imag} */,
  {32'h408db01e, 32'hc1309096} /* (30, 27, 5) {real, imag} */,
  {32'hc0d86bdf, 32'h40a1507a} /* (30, 27, 4) {real, imag} */,
  {32'hbf7a62fd, 32'hc0a326cb} /* (30, 27, 3) {real, imag} */,
  {32'hc07ca3ca, 32'hc178ce92} /* (30, 27, 2) {real, imag} */,
  {32'h4184c940, 32'h422cd933} /* (30, 27, 1) {real, imag} */,
  {32'h419be0a5, 32'h41f47949} /* (30, 27, 0) {real, imag} */,
  {32'h40238bd0, 32'h40626806} /* (30, 26, 31) {real, imag} */,
  {32'h409c197e, 32'hc101e3d7} /* (30, 26, 30) {real, imag} */,
  {32'hc080c0d5, 32'hc02c802b} /* (30, 26, 29) {real, imag} */,
  {32'h3f539fc9, 32'hbfd635a2} /* (30, 26, 28) {real, imag} */,
  {32'h3fa1cc06, 32'hbff49ab2} /* (30, 26, 27) {real, imag} */,
  {32'hc029fed6, 32'hc0365bf5} /* (30, 26, 26) {real, imag} */,
  {32'h3ffad705, 32'h3f785683} /* (30, 26, 25) {real, imag} */,
  {32'hbfe1e2a0, 32'hc0707d6f} /* (30, 26, 24) {real, imag} */,
  {32'h4012321f, 32'hbfd9d84b} /* (30, 26, 23) {real, imag} */,
  {32'h3e9df42b, 32'h408041fe} /* (30, 26, 22) {real, imag} */,
  {32'hbf3c6d95, 32'hbff9dc8c} /* (30, 26, 21) {real, imag} */,
  {32'h3f346531, 32'h3f9fd1fa} /* (30, 26, 20) {real, imag} */,
  {32'hc037e0fd, 32'hbf7c8ae1} /* (30, 26, 19) {real, imag} */,
  {32'h3f267245, 32'h3fdefdf0} /* (30, 26, 18) {real, imag} */,
  {32'h3f1625de, 32'hbe80581e} /* (30, 26, 17) {real, imag} */,
  {32'hbf606ef8, 32'hbecd8e21} /* (30, 26, 16) {real, imag} */,
  {32'h3e6907f6, 32'h3f259052} /* (30, 26, 15) {real, imag} */,
  {32'h3ead0d58, 32'h3e52d7f9} /* (30, 26, 14) {real, imag} */,
  {32'h3fb8331e, 32'h3e67160f} /* (30, 26, 13) {real, imag} */,
  {32'hbf15bcf3, 32'hbfbf2ee7} /* (30, 26, 12) {real, imag} */,
  {32'hc006ebfd, 32'hc0142b5a} /* (30, 26, 11) {real, imag} */,
  {32'h3e920a76, 32'hbf65d316} /* (30, 26, 10) {real, imag} */,
  {32'hbf06f21d, 32'hbdff462b} /* (30, 26, 9) {real, imag} */,
  {32'hc03f8c37, 32'hbfd0db2f} /* (30, 26, 8) {real, imag} */,
  {32'hbef86617, 32'h3fb44006} /* (30, 26, 7) {real, imag} */,
  {32'hc00cb8f6, 32'hbf0ff9e0} /* (30, 26, 6) {real, imag} */,
  {32'hc01e9d42, 32'h40170f2b} /* (30, 26, 5) {real, imag} */,
  {32'hc017f02a, 32'hc00ecb35} /* (30, 26, 4) {real, imag} */,
  {32'h3f60b55b, 32'h40179db9} /* (30, 26, 3) {real, imag} */,
  {32'hc051de7a, 32'hc0a1caec} /* (30, 26, 2) {real, imag} */,
  {32'h404bb3b6, 32'hc0277838} /* (30, 26, 1) {real, imag} */,
  {32'hc06274b9, 32'h40494e40} /* (30, 26, 0) {real, imag} */,
  {32'hc1167e39, 32'hc0a44690} /* (30, 25, 31) {real, imag} */,
  {32'h40274e72, 32'h3f530a15} /* (30, 25, 30) {real, imag} */,
  {32'h4037e9fa, 32'h41004d3a} /* (30, 25, 29) {real, imag} */,
  {32'hc00d6311, 32'h3e05ba3f} /* (30, 25, 28) {real, imag} */,
  {32'h4022c710, 32'h404a8afc} /* (30, 25, 27) {real, imag} */,
  {32'hbfc98102, 32'h3ef89af1} /* (30, 25, 26) {real, imag} */,
  {32'hbec72a5c, 32'hc0d30df8} /* (30, 25, 25) {real, imag} */,
  {32'h3f03472b, 32'h40235838} /* (30, 25, 24) {real, imag} */,
  {32'hbf5ae840, 32'h4027a841} /* (30, 25, 23) {real, imag} */,
  {32'h3f3c43fa, 32'hbf84fd2b} /* (30, 25, 22) {real, imag} */,
  {32'h402175b8, 32'hc04ce749} /* (30, 25, 21) {real, imag} */,
  {32'h3f9f5592, 32'hbf92480d} /* (30, 25, 20) {real, imag} */,
  {32'h3e45a926, 32'h3f4caef3} /* (30, 25, 19) {real, imag} */,
  {32'hbd576c77, 32'hbfc76369} /* (30, 25, 18) {real, imag} */,
  {32'h3fb87925, 32'hbf5959ad} /* (30, 25, 17) {real, imag} */,
  {32'hbe857fd8, 32'hbf0095ee} /* (30, 25, 16) {real, imag} */,
  {32'h3da4052b, 32'h3f3d2c56} /* (30, 25, 15) {real, imag} */,
  {32'hc038e7a0, 32'h3f4912eb} /* (30, 25, 14) {real, imag} */,
  {32'hbdf28afb, 32'hbfca0434} /* (30, 25, 13) {real, imag} */,
  {32'hbfdfe10c, 32'h3efba5af} /* (30, 25, 12) {real, imag} */,
  {32'h3fb0f6f3, 32'hc08eb314} /* (30, 25, 11) {real, imag} */,
  {32'hbeaa7cf2, 32'h3f8681e6} /* (30, 25, 10) {real, imag} */,
  {32'h408182b7, 32'hbf21fd47} /* (30, 25, 9) {real, imag} */,
  {32'h4008b29b, 32'h3e8c398b} /* (30, 25, 8) {real, imag} */,
  {32'hc00d0b7e, 32'h3eb9f4ec} /* (30, 25, 7) {real, imag} */,
  {32'h3f02cfbb, 32'h3f682430} /* (30, 25, 6) {real, imag} */,
  {32'h3fb26ac5, 32'h4027bce3} /* (30, 25, 5) {real, imag} */,
  {32'hbf8ba9ce, 32'h3eae69d9} /* (30, 25, 4) {real, imag} */,
  {32'hbfcb3b67, 32'hbc1a4fd3} /* (30, 25, 3) {real, imag} */,
  {32'h408f15c2, 32'h4065677e} /* (30, 25, 2) {real, imag} */,
  {32'hbf31d5e5, 32'hc0d6cb0f} /* (30, 25, 1) {real, imag} */,
  {32'hc0902899, 32'hc0dbe2db} /* (30, 25, 0) {real, imag} */,
  {32'h41289ab7, 32'h40c029c6} /* (30, 24, 31) {real, imag} */,
  {32'hc0ad8628, 32'hc0f40b15} /* (30, 24, 30) {real, imag} */,
  {32'hc089f15e, 32'hc02564b9} /* (30, 24, 29) {real, imag} */,
  {32'h40473fe4, 32'h40c0d3a0} /* (30, 24, 28) {real, imag} */,
  {32'hbffa1cf2, 32'hc0adffa5} /* (30, 24, 27) {real, imag} */,
  {32'h3bf8e284, 32'h3e6ad753} /* (30, 24, 26) {real, imag} */,
  {32'hc090ba36, 32'hc00de5ba} /* (30, 24, 25) {real, imag} */,
  {32'h4056f660, 32'hbe8fb5fa} /* (30, 24, 24) {real, imag} */,
  {32'h40218c45, 32'h3f9f36f7} /* (30, 24, 23) {real, imag} */,
  {32'hbea13ce6, 32'hbf2268e3} /* (30, 24, 22) {real, imag} */,
  {32'hc013c0dc, 32'hbf42146b} /* (30, 24, 21) {real, imag} */,
  {32'hbfcd36b5, 32'hbeb02dd2} /* (30, 24, 20) {real, imag} */,
  {32'hbf662476, 32'hbd59a64b} /* (30, 24, 19) {real, imag} */,
  {32'h3f250ecc, 32'hbf59cca0} /* (30, 24, 18) {real, imag} */,
  {32'h3f874e11, 32'h3fc5b43c} /* (30, 24, 17) {real, imag} */,
  {32'hbfea807a, 32'hbfbd26e9} /* (30, 24, 16) {real, imag} */,
  {32'hbd30e27d, 32'hbf31edd0} /* (30, 24, 15) {real, imag} */,
  {32'h3fd47777, 32'hbf506108} /* (30, 24, 14) {real, imag} */,
  {32'h3e9ea54d, 32'h3fbc711c} /* (30, 24, 13) {real, imag} */,
  {32'hbff72724, 32'hbfb2ee79} /* (30, 24, 12) {real, imag} */,
  {32'h3fc694bd, 32'hc00b5e85} /* (30, 24, 11) {real, imag} */,
  {32'hc002f45a, 32'h3f59c352} /* (30, 24, 10) {real, imag} */,
  {32'h40397b0b, 32'hbf6b4a8f} /* (30, 24, 9) {real, imag} */,
  {32'hc05e7ebf, 32'hc0bb1f41} /* (30, 24, 8) {real, imag} */,
  {32'h409cf4d5, 32'hbf3138e0} /* (30, 24, 7) {real, imag} */,
  {32'hc08aa8c3, 32'hbf60e139} /* (30, 24, 6) {real, imag} */,
  {32'hbf906945, 32'hc01cccc6} /* (30, 24, 5) {real, imag} */,
  {32'h3d775cf6, 32'hbf67e0b4} /* (30, 24, 4) {real, imag} */,
  {32'h3ff43654, 32'h4079815b} /* (30, 24, 3) {real, imag} */,
  {32'hc0de3753, 32'hc1726839} /* (30, 24, 2) {real, imag} */,
  {32'h4154b7ac, 32'h41a9e599} /* (30, 24, 1) {real, imag} */,
  {32'h40deb631, 32'h40a83d2b} /* (30, 24, 0) {real, imag} */,
  {32'hc028eaae, 32'hc0d2b6a8} /* (30, 23, 31) {real, imag} */,
  {32'h40460be4, 32'hc07fc8d5} /* (30, 23, 30) {real, imag} */,
  {32'hbfa4ff1f, 32'h3f855fa1} /* (30, 23, 29) {real, imag} */,
  {32'hc01d3f72, 32'h3fafa453} /* (30, 23, 28) {real, imag} */,
  {32'hc04c6bcd, 32'h3fc2a556} /* (30, 23, 27) {real, imag} */,
  {32'h3f199939, 32'h3f0617c5} /* (30, 23, 26) {real, imag} */,
  {32'hbfb42236, 32'h4004d0bd} /* (30, 23, 25) {real, imag} */,
  {32'hbf18b5e1, 32'hbece7eb5} /* (30, 23, 24) {real, imag} */,
  {32'h40358163, 32'h3fa2e287} /* (30, 23, 23) {real, imag} */,
  {32'hc06db83e, 32'h403877aa} /* (30, 23, 22) {real, imag} */,
  {32'hbfb954fa, 32'hbf68b539} /* (30, 23, 21) {real, imag} */,
  {32'hbf9d1d6d, 32'h3e1da932} /* (30, 23, 20) {real, imag} */,
  {32'h3fd913c2, 32'hbf81c364} /* (30, 23, 19) {real, imag} */,
  {32'hc022b762, 32'hbf0320cb} /* (30, 23, 18) {real, imag} */,
  {32'h3f2416ef, 32'hbf20d197} /* (30, 23, 17) {real, imag} */,
  {32'hbf80ebe6, 32'hbf754af4} /* (30, 23, 16) {real, imag} */,
  {32'h3f89dd3d, 32'h40137581} /* (30, 23, 15) {real, imag} */,
  {32'h40497aa0, 32'h3fbb4ae7} /* (30, 23, 14) {real, imag} */,
  {32'hbe8daafd, 32'hc02c120f} /* (30, 23, 13) {real, imag} */,
  {32'h3f78b39c, 32'h401b27c7} /* (30, 23, 12) {real, imag} */,
  {32'h3e945fae, 32'h3fd5e613} /* (30, 23, 11) {real, imag} */,
  {32'hbef11a1d, 32'h3f3f43d8} /* (30, 23, 10) {real, imag} */,
  {32'hc01b239b, 32'hc01b133e} /* (30, 23, 9) {real, imag} */,
  {32'h400725ae, 32'h4021748e} /* (30, 23, 8) {real, imag} */,
  {32'h3f862c69, 32'hbfc58c72} /* (30, 23, 7) {real, imag} */,
  {32'h4011be92, 32'hbf85e969} /* (30, 23, 6) {real, imag} */,
  {32'h3f36d268, 32'h40d82942} /* (30, 23, 5) {real, imag} */,
  {32'hbfb61e3f, 32'hbf5cc55e} /* (30, 23, 4) {real, imag} */,
  {32'hc0256bd3, 32'hc04505af} /* (30, 23, 3) {real, imag} */,
  {32'h40daef62, 32'hc0c21e1c} /* (30, 23, 2) {real, imag} */,
  {32'hc08d956f, 32'h40fe74a5} /* (30, 23, 1) {real, imag} */,
  {32'h3fe6aa3a, 32'h3fa10770} /* (30, 23, 0) {real, imag} */,
  {32'hc055e24b, 32'hc0c04817} /* (30, 22, 31) {real, imag} */,
  {32'h40ca3399, 32'h3f7cf704} /* (30, 22, 30) {real, imag} */,
  {32'hbe5499ed, 32'h3fefe13c} /* (30, 22, 29) {real, imag} */,
  {32'hc05fddc0, 32'h3fe1eb4a} /* (30, 22, 28) {real, imag} */,
  {32'h3be6d593, 32'hbf7fb755} /* (30, 22, 27) {real, imag} */,
  {32'h3fd5329b, 32'h4017534f} /* (30, 22, 26) {real, imag} */,
  {32'h3f19e2df, 32'hc09b6fca} /* (30, 22, 25) {real, imag} */,
  {32'hc0199f4c, 32'hbfe61655} /* (30, 22, 24) {real, imag} */,
  {32'h401789b3, 32'hc052604d} /* (30, 22, 23) {real, imag} */,
  {32'h409eae66, 32'h3ff19a02} /* (30, 22, 22) {real, imag} */,
  {32'h3e2c0539, 32'hc0165883} /* (30, 22, 21) {real, imag} */,
  {32'hc0656dbf, 32'hbf05e75c} /* (30, 22, 20) {real, imag} */,
  {32'h40165474, 32'h3fe402ac} /* (30, 22, 19) {real, imag} */,
  {32'h3f34b0e5, 32'h3ec45672} /* (30, 22, 18) {real, imag} */,
  {32'hc01b9be4, 32'h3fa3ff80} /* (30, 22, 17) {real, imag} */,
  {32'hbfd7c82d, 32'hbd7250b7} /* (30, 22, 16) {real, imag} */,
  {32'hbffc6049, 32'hbfd17e7b} /* (30, 22, 15) {real, imag} */,
  {32'h4000c9de, 32'h3f560d0f} /* (30, 22, 14) {real, imag} */,
  {32'h3fff0565, 32'h4004c592} /* (30, 22, 13) {real, imag} */,
  {32'hbfb4301e, 32'h3ff7e4cf} /* (30, 22, 12) {real, imag} */,
  {32'hc01d897c, 32'h3fa9fcc3} /* (30, 22, 11) {real, imag} */,
  {32'hbdda7a25, 32'hc03ec3da} /* (30, 22, 10) {real, imag} */,
  {32'hc03c32e3, 32'hc006a7fd} /* (30, 22, 9) {real, imag} */,
  {32'h40226636, 32'h3f62f228} /* (30, 22, 8) {real, imag} */,
  {32'hbd483500, 32'h3f1892b8} /* (30, 22, 7) {real, imag} */,
  {32'h3fa67089, 32'hc012ed46} /* (30, 22, 6) {real, imag} */,
  {32'h3f27d14f, 32'h404970a9} /* (30, 22, 5) {real, imag} */,
  {32'h3f7eaa66, 32'hbfef38a1} /* (30, 22, 4) {real, imag} */,
  {32'hbf83bf4a, 32'hc0860765} /* (30, 22, 3) {real, imag} */,
  {32'h408cb370, 32'h3efde828} /* (30, 22, 2) {real, imag} */,
  {32'hc0e89c19, 32'hc014e960} /* (30, 22, 1) {real, imag} */,
  {32'hbfa41854, 32'hbffee284} /* (30, 22, 0) {real, imag} */,
  {32'h41166d0e, 32'h3e7daeec} /* (30, 21, 31) {real, imag} */,
  {32'hc1029f2a, 32'h407d0d03} /* (30, 21, 30) {real, imag} */,
  {32'hc059715e, 32'hc0122ab5} /* (30, 21, 29) {real, imag} */,
  {32'hbf28cb1d, 32'h3f99c103} /* (30, 21, 28) {real, imag} */,
  {32'hbfcc48e4, 32'h3eb7c760} /* (30, 21, 27) {real, imag} */,
  {32'h3fc02eab, 32'h3f46f7be} /* (30, 21, 26) {real, imag} */,
  {32'h3e305409, 32'h3ffd4f3e} /* (30, 21, 25) {real, imag} */,
  {32'h3ed51a4a, 32'hbfaf05c1} /* (30, 21, 24) {real, imag} */,
  {32'hc00cf8c0, 32'hc086a73a} /* (30, 21, 23) {real, imag} */,
  {32'h402ffe7e, 32'hbb180c4c} /* (30, 21, 22) {real, imag} */,
  {32'hbfde87e3, 32'h4088ccaa} /* (30, 21, 21) {real, imag} */,
  {32'hbfebb5b5, 32'hc0036bba} /* (30, 21, 20) {real, imag} */,
  {32'h3f60d02c, 32'h3fa747bb} /* (30, 21, 19) {real, imag} */,
  {32'h3e84ae6e, 32'hc03fd7fb} /* (30, 21, 18) {real, imag} */,
  {32'h3f9f6b74, 32'hbf166674} /* (30, 21, 17) {real, imag} */,
  {32'hbf279864, 32'h3f92f11b} /* (30, 21, 16) {real, imag} */,
  {32'h3df9183f, 32'hbeaf0472} /* (30, 21, 15) {real, imag} */,
  {32'h3fe48f97, 32'h4008f1cc} /* (30, 21, 14) {real, imag} */,
  {32'hc0024b73, 32'h3fdc7722} /* (30, 21, 13) {real, imag} */,
  {32'hc0016e2d, 32'hbf873c1f} /* (30, 21, 12) {real, imag} */,
  {32'hbf1a43b3, 32'hc02a7ae5} /* (30, 21, 11) {real, imag} */,
  {32'h3f97c63e, 32'h3f742f40} /* (30, 21, 10) {real, imag} */,
  {32'h4023b5a1, 32'h401dc97a} /* (30, 21, 9) {real, imag} */,
  {32'hbe6cc9f7, 32'h3f71f8de} /* (30, 21, 8) {real, imag} */,
  {32'h3fdb5843, 32'hbeb255f4} /* (30, 21, 7) {real, imag} */,
  {32'h4035ff47, 32'hc008ef82} /* (30, 21, 6) {real, imag} */,
  {32'hbf10a447, 32'h3f3a1691} /* (30, 21, 5) {real, imag} */,
  {32'hbff18544, 32'hbfc52931} /* (30, 21, 4) {real, imag} */,
  {32'h3dc8369d, 32'hc0174600} /* (30, 21, 3) {real, imag} */,
  {32'hc097ba39, 32'hc0bdb837} /* (30, 21, 2) {real, imag} */,
  {32'h40aeaf72, 32'h409553f5} /* (30, 21, 1) {real, imag} */,
  {32'h4121d09a, 32'h41115250} /* (30, 21, 0) {real, imag} */,
  {32'h3f2d7aa5, 32'hbffd3363} /* (30, 20, 31) {real, imag} */,
  {32'hbf10ce1c, 32'h3fad2953} /* (30, 20, 30) {real, imag} */,
  {32'hbfd2457b, 32'hc06dc6dc} /* (30, 20, 29) {real, imag} */,
  {32'hbf257e10, 32'h3fe19a1e} /* (30, 20, 28) {real, imag} */,
  {32'hbf3b984a, 32'h403ea07e} /* (30, 20, 27) {real, imag} */,
  {32'h3ff0e87e, 32'h3fbe53b7} /* (30, 20, 26) {real, imag} */,
  {32'hbe2c4b4f, 32'h3dc432d0} /* (30, 20, 25) {real, imag} */,
  {32'h404a452c, 32'h40538745} /* (30, 20, 24) {real, imag} */,
  {32'h3f75a34d, 32'h3ed05fd0} /* (30, 20, 23) {real, imag} */,
  {32'hbf805a4c, 32'hc042b7c7} /* (30, 20, 22) {real, imag} */,
  {32'h3f5f4ba3, 32'hbfa1c197} /* (30, 20, 21) {real, imag} */,
  {32'hbfed576a, 32'h3fb68ee0} /* (30, 20, 20) {real, imag} */,
  {32'h3ff531d8, 32'hbf9aedee} /* (30, 20, 19) {real, imag} */,
  {32'hbf62b5d7, 32'h3ff69330} /* (30, 20, 18) {real, imag} */,
  {32'hbf0189ff, 32'h3f60a596} /* (30, 20, 17) {real, imag} */,
  {32'hbd3d68a9, 32'hbf63e5b6} /* (30, 20, 16) {real, imag} */,
  {32'hbfafabda, 32'h3fce57c0} /* (30, 20, 15) {real, imag} */,
  {32'hbcb80cfa, 32'hbff0b890} /* (30, 20, 14) {real, imag} */,
  {32'hc0072257, 32'h3d3942a2} /* (30, 20, 13) {real, imag} */,
  {32'hbf87a7ba, 32'h3e2ea960} /* (30, 20, 12) {real, imag} */,
  {32'h3f1e3824, 32'h3f728698} /* (30, 20, 11) {real, imag} */,
  {32'hbfa0ca4b, 32'hbfe53003} /* (30, 20, 10) {real, imag} */,
  {32'h3ecd4d3c, 32'hbcbbbd92} /* (30, 20, 9) {real, imag} */,
  {32'h401f4d75, 32'hbe6b58fd} /* (30, 20, 8) {real, imag} */,
  {32'hc001c4bd, 32'h3f8a893b} /* (30, 20, 7) {real, imag} */,
  {32'h3fee84ea, 32'h404239ad} /* (30, 20, 6) {real, imag} */,
  {32'hbf9a5334, 32'hbfe84c42} /* (30, 20, 5) {real, imag} */,
  {32'hbe86f8e4, 32'h3f363068} /* (30, 20, 4) {real, imag} */,
  {32'h3fcd2e63, 32'h4081f2fe} /* (30, 20, 3) {real, imag} */,
  {32'h3f600548, 32'hc01a4eb5} /* (30, 20, 2) {real, imag} */,
  {32'hbf51c6c6, 32'hbfc55aaf} /* (30, 20, 1) {real, imag} */,
  {32'hbf7bfbb2, 32'hbe700dbf} /* (30, 20, 0) {real, imag} */,
  {32'hbfc53271, 32'h3eb9a809} /* (30, 19, 31) {real, imag} */,
  {32'hbfb6d199, 32'h3f14cf3d} /* (30, 19, 30) {real, imag} */,
  {32'hbd64f06c, 32'h3f0a2adb} /* (30, 19, 29) {real, imag} */,
  {32'hbf948cb3, 32'h3fdcf08a} /* (30, 19, 28) {real, imag} */,
  {32'hc00a1492, 32'h3dd1c659} /* (30, 19, 27) {real, imag} */,
  {32'h3f8de987, 32'h3f8c99a5} /* (30, 19, 26) {real, imag} */,
  {32'hbdd70d4c, 32'hc073100a} /* (30, 19, 25) {real, imag} */,
  {32'h3eaa56c2, 32'h3fc8ab17} /* (30, 19, 24) {real, imag} */,
  {32'h3ed75885, 32'h3e2f0b51} /* (30, 19, 23) {real, imag} */,
  {32'hbea494ea, 32'hbeded19e} /* (30, 19, 22) {real, imag} */,
  {32'h3f5e4a31, 32'hbf753208} /* (30, 19, 21) {real, imag} */,
  {32'h3e3a3e03, 32'h403085b7} /* (30, 19, 20) {real, imag} */,
  {32'hbeb81d64, 32'hbfa151b2} /* (30, 19, 19) {real, imag} */,
  {32'hbea9eae6, 32'hc04c2600} /* (30, 19, 18) {real, imag} */,
  {32'h3edb208e, 32'h3eade901} /* (30, 19, 17) {real, imag} */,
  {32'h3f1c5c45, 32'hbea8beff} /* (30, 19, 16) {real, imag} */,
  {32'hbe994fc6, 32'hbf9f8d6b} /* (30, 19, 15) {real, imag} */,
  {32'hbd837598, 32'h3fb323c2} /* (30, 19, 14) {real, imag} */,
  {32'hbf00f903, 32'h3f23f217} /* (30, 19, 13) {real, imag} */,
  {32'h3f251e72, 32'hbf11f805} /* (30, 19, 12) {real, imag} */,
  {32'hbd15af26, 32'hbe223007} /* (30, 19, 11) {real, imag} */,
  {32'hbea8a7bb, 32'h3fa629ad} /* (30, 19, 10) {real, imag} */,
  {32'hbfaf0d8c, 32'h3da2993d} /* (30, 19, 9) {real, imag} */,
  {32'hbf192290, 32'hbf8897a3} /* (30, 19, 8) {real, imag} */,
  {32'h3ff1cfb7, 32'h3f846642} /* (30, 19, 7) {real, imag} */,
  {32'hbf1ff56d, 32'hbe846584} /* (30, 19, 6) {real, imag} */,
  {32'hbf91f709, 32'h3f1f2254} /* (30, 19, 5) {real, imag} */,
  {32'h3ee560b9, 32'hbf45e288} /* (30, 19, 4) {real, imag} */,
  {32'hbf684ed6, 32'hbd915c11} /* (30, 19, 3) {real, imag} */,
  {32'h4016249b, 32'hbfda266c} /* (30, 19, 2) {real, imag} */,
  {32'h3d87f1c7, 32'h3f94acf3} /* (30, 19, 1) {real, imag} */,
  {32'h3ea36205, 32'hbfcf19ae} /* (30, 19, 0) {real, imag} */,
  {32'h4071b038, 32'hbf406ef5} /* (30, 18, 31) {real, imag} */,
  {32'hc06c1028, 32'hbe8b2706} /* (30, 18, 30) {real, imag} */,
  {32'hbf8fe52f, 32'h3dce051e} /* (30, 18, 29) {real, imag} */,
  {32'h40648148, 32'h40796f1b} /* (30, 18, 28) {real, imag} */,
  {32'hbf888358, 32'h3e8c922d} /* (30, 18, 27) {real, imag} */,
  {32'hbfb11a5c, 32'hbe0df049} /* (30, 18, 26) {real, imag} */,
  {32'h4029df99, 32'h3efd6d1a} /* (30, 18, 25) {real, imag} */,
  {32'hbf671e1c, 32'h3f3f2154} /* (30, 18, 24) {real, imag} */,
  {32'hbf4be799, 32'h3f4be052} /* (30, 18, 23) {real, imag} */,
  {32'h3c60277b, 32'h3ebb346d} /* (30, 18, 22) {real, imag} */,
  {32'h3fc3bf37, 32'h4024d126} /* (30, 18, 21) {real, imag} */,
  {32'h3f3512f6, 32'hbdf1ad91} /* (30, 18, 20) {real, imag} */,
  {32'h3f6ee5ad, 32'h3e206ed3} /* (30, 18, 19) {real, imag} */,
  {32'h3f93e4fb, 32'h3f124506} /* (30, 18, 18) {real, imag} */,
  {32'h3f9cc3d5, 32'h3fac8da3} /* (30, 18, 17) {real, imag} */,
  {32'h3f3c6ac0, 32'hbf84fc21} /* (30, 18, 16) {real, imag} */,
  {32'h3f51c217, 32'hbfd05436} /* (30, 18, 15) {real, imag} */,
  {32'hbf569975, 32'hbdbd897a} /* (30, 18, 14) {real, imag} */,
  {32'h3f993cb2, 32'hc02a1f5c} /* (30, 18, 13) {real, imag} */,
  {32'h400eed84, 32'h3f08801f} /* (30, 18, 12) {real, imag} */,
  {32'h3f01c0b1, 32'h3f806591} /* (30, 18, 11) {real, imag} */,
  {32'hbf7a8ea2, 32'h3e9ff295} /* (30, 18, 10) {real, imag} */,
  {32'h3f60ef85, 32'h3f155e4f} /* (30, 18, 9) {real, imag} */,
  {32'h3e862827, 32'hbfa64f07} /* (30, 18, 8) {real, imag} */,
  {32'h3dc90418, 32'hbfbddf0e} /* (30, 18, 7) {real, imag} */,
  {32'h40920ed7, 32'h3eff3c88} /* (30, 18, 6) {real, imag} */,
  {32'hc011dcb3, 32'hbe5c4feb} /* (30, 18, 5) {real, imag} */,
  {32'h400f191e, 32'hbf16e86f} /* (30, 18, 4) {real, imag} */,
  {32'hbfa73ed6, 32'h400448b9} /* (30, 18, 3) {real, imag} */,
  {32'hc0856d79, 32'hbfe3a18f} /* (30, 18, 2) {real, imag} */,
  {32'h4095b446, 32'h404728ae} /* (30, 18, 1) {real, imag} */,
  {32'h40679b7a, 32'hbf12f625} /* (30, 18, 0) {real, imag} */,
  {32'hc0275bc6, 32'h400bd609} /* (30, 17, 31) {real, imag} */,
  {32'h3ffdff6d, 32'h3fd64126} /* (30, 17, 30) {real, imag} */,
  {32'hbeb9abda, 32'hbfb41cb9} /* (30, 17, 29) {real, imag} */,
  {32'h400921f4, 32'h3ee9a74a} /* (30, 17, 28) {real, imag} */,
  {32'hbe8f61ef, 32'hbf4c832f} /* (30, 17, 27) {real, imag} */,
  {32'hc089e295, 32'h3e6af85e} /* (30, 17, 26) {real, imag} */,
  {32'h4025073f, 32'h3fbfd775} /* (30, 17, 25) {real, imag} */,
  {32'hbf9d4eda, 32'hbed8f8de} /* (30, 17, 24) {real, imag} */,
  {32'h3f738082, 32'h3ec75fb0} /* (30, 17, 23) {real, imag} */,
  {32'hbda8d4c4, 32'h3fcd6ddb} /* (30, 17, 22) {real, imag} */,
  {32'h3fb281e5, 32'hbfb785a1} /* (30, 17, 21) {real, imag} */,
  {32'h400b4d36, 32'hbedb924e} /* (30, 17, 20) {real, imag} */,
  {32'h3ec18d89, 32'h3f3b481f} /* (30, 17, 19) {real, imag} */,
  {32'hbf302cb2, 32'hbf1c0c3e} /* (30, 17, 18) {real, imag} */,
  {32'h3f99762f, 32'h3f4db926} /* (30, 17, 17) {real, imag} */,
  {32'hbeb61216, 32'h3f190227} /* (30, 17, 16) {real, imag} */,
  {32'h3e61fc98, 32'hbebf007a} /* (30, 17, 15) {real, imag} */,
  {32'hbf1dc105, 32'hbed29d0c} /* (30, 17, 14) {real, imag} */,
  {32'hbf290bf8, 32'h3f98aea4} /* (30, 17, 13) {real, imag} */,
  {32'h3f4dbaf0, 32'h3e99a59d} /* (30, 17, 12) {real, imag} */,
  {32'h3f8a79e4, 32'hbe42fda9} /* (30, 17, 11) {real, imag} */,
  {32'h3fe98f3b, 32'hbfbefbe2} /* (30, 17, 10) {real, imag} */,
  {32'h3fd241c1, 32'hbff9c11c} /* (30, 17, 9) {real, imag} */,
  {32'h3f87ed2e, 32'hbf26f9ca} /* (30, 17, 8) {real, imag} */,
  {32'h3e0da0c3, 32'hbef5fb57} /* (30, 17, 7) {real, imag} */,
  {32'hc0237e66, 32'hbeea66a0} /* (30, 17, 6) {real, imag} */,
  {32'h3f7893a9, 32'h3ed54d85} /* (30, 17, 5) {real, imag} */,
  {32'hbe973e0f, 32'hbf219783} /* (30, 17, 4) {real, imag} */,
  {32'h3fa055cc, 32'hc02e91d4} /* (30, 17, 3) {real, imag} */,
  {32'h3f499053, 32'h3fbaadcf} /* (30, 17, 2) {real, imag} */,
  {32'hbf87beba, 32'h3fc0b241} /* (30, 17, 1) {real, imag} */,
  {32'hbfd39531, 32'h3f2f58f4} /* (30, 17, 0) {real, imag} */,
  {32'h3d2a8ef2, 32'hbf0b27ee} /* (30, 16, 31) {real, imag} */,
  {32'hbf95846a, 32'h3f2e5dc4} /* (30, 16, 30) {real, imag} */,
  {32'hbf6ee17e, 32'hbf35a41e} /* (30, 16, 29) {real, imag} */,
  {32'h3fd1cd1f, 32'hbff36b99} /* (30, 16, 28) {real, imag} */,
  {32'h3f9b1824, 32'hbe8661d1} /* (30, 16, 27) {real, imag} */,
  {32'h3f64b4d5, 32'h3f2a2c1d} /* (30, 16, 26) {real, imag} */,
  {32'hbe67cc25, 32'h3dd75498} /* (30, 16, 25) {real, imag} */,
  {32'hbed7b09e, 32'hbf75ec2b} /* (30, 16, 24) {real, imag} */,
  {32'h3f3e7f8d, 32'hbf8ae11f} /* (30, 16, 23) {real, imag} */,
  {32'h3fe4ca01, 32'hbf200283} /* (30, 16, 22) {real, imag} */,
  {32'hbf93c723, 32'hbe9a27bf} /* (30, 16, 21) {real, imag} */,
  {32'hbd400c2e, 32'h3fb1e9be} /* (30, 16, 20) {real, imag} */,
  {32'hbfa0d6a2, 32'h4036ebde} /* (30, 16, 19) {real, imag} */,
  {32'h3e19b8b7, 32'hbe5f7184} /* (30, 16, 18) {real, imag} */,
  {32'hbfc3e2ff, 32'hc005a201} /* (30, 16, 17) {real, imag} */,
  {32'hbeb8eca6, 32'hbf6609bd} /* (30, 16, 16) {real, imag} */,
  {32'hbf153aa6, 32'hbf8245c7} /* (30, 16, 15) {real, imag} */,
  {32'h3f903413, 32'hbf51521f} /* (30, 16, 14) {real, imag} */,
  {32'hbf96c174, 32'h3e11cd9d} /* (30, 16, 13) {real, imag} */,
  {32'hbeefe73a, 32'hbe9dae99} /* (30, 16, 12) {real, imag} */,
  {32'h3fb2a05e, 32'hbf80d188} /* (30, 16, 11) {real, imag} */,
  {32'hbd22b248, 32'hc03f956f} /* (30, 16, 10) {real, imag} */,
  {32'h3f50a68f, 32'h3eff9adf} /* (30, 16, 9) {real, imag} */,
  {32'h3fdce25e, 32'h3f813f15} /* (30, 16, 8) {real, imag} */,
  {32'hbf1dec47, 32'hbf59efa8} /* (30, 16, 7) {real, imag} */,
  {32'hbfe45997, 32'hbefe6e89} /* (30, 16, 6) {real, imag} */,
  {32'hbf5b97de, 32'hbf9021bf} /* (30, 16, 5) {real, imag} */,
  {32'h3dbce757, 32'hbe844ff9} /* (30, 16, 4) {real, imag} */,
  {32'h3f535c47, 32'h3e216b3d} /* (30, 16, 3) {real, imag} */,
  {32'hbe9b09e2, 32'hbc23c428} /* (30, 16, 2) {real, imag} */,
  {32'hbfc11956, 32'h3fb36792} /* (30, 16, 1) {real, imag} */,
  {32'hbfbd63ef, 32'h3f1c93f1} /* (30, 16, 0) {real, imag} */,
  {32'h408264ae, 32'h3fa46882} /* (30, 15, 31) {real, imag} */,
  {32'hc03989f2, 32'h3e4cdd42} /* (30, 15, 30) {real, imag} */,
  {32'h3d090f9b, 32'hbf5f4cc2} /* (30, 15, 29) {real, imag} */,
  {32'hbe63ec37, 32'hc0137263} /* (30, 15, 28) {real, imag} */,
  {32'h3f9b2e0d, 32'hbc8f4fce} /* (30, 15, 27) {real, imag} */,
  {32'h3f8fe955, 32'hbf9b4580} /* (30, 15, 26) {real, imag} */,
  {32'hbe52aa6a, 32'h3f8f971e} /* (30, 15, 25) {real, imag} */,
  {32'h3f8426c4, 32'hbf1f4ffd} /* (30, 15, 24) {real, imag} */,
  {32'hbf308bb1, 32'h3ee0ce75} /* (30, 15, 23) {real, imag} */,
  {32'h3fe2f660, 32'h3efbe3af} /* (30, 15, 22) {real, imag} */,
  {32'hbf1913e5, 32'hbf5c19cd} /* (30, 15, 21) {real, imag} */,
  {32'hbead762c, 32'hbdd9efe1} /* (30, 15, 20) {real, imag} */,
  {32'hbeb83b4f, 32'hbe4f7675} /* (30, 15, 19) {real, imag} */,
  {32'h3ede5885, 32'h4021e01a} /* (30, 15, 18) {real, imag} */,
  {32'hbf7ea8cd, 32'hc016321b} /* (30, 15, 17) {real, imag} */,
  {32'h3e8b3d63, 32'h3fb1706e} /* (30, 15, 16) {real, imag} */,
  {32'hbf962a58, 32'h3d634a7c} /* (30, 15, 15) {real, imag} */,
  {32'hc0514631, 32'hbf54ac0d} /* (30, 15, 14) {real, imag} */,
  {32'h3e36842d, 32'hbd841183} /* (30, 15, 13) {real, imag} */,
  {32'hbf378cbe, 32'h4001e98b} /* (30, 15, 12) {real, imag} */,
  {32'h3eca1e25, 32'hbffb9fad} /* (30, 15, 11) {real, imag} */,
  {32'h3fc862b8, 32'h3fb6139f} /* (30, 15, 10) {real, imag} */,
  {32'h3fd13bc1, 32'hbe38cfb0} /* (30, 15, 9) {real, imag} */,
  {32'hbf64a18c, 32'hbf6f5abd} /* (30, 15, 8) {real, imag} */,
  {32'h3b52da9e, 32'hc036722c} /* (30, 15, 7) {real, imag} */,
  {32'h3fcee70e, 32'h3fdd1bcb} /* (30, 15, 6) {real, imag} */,
  {32'hbf2c1aa8, 32'hbf832976} /* (30, 15, 5) {real, imag} */,
  {32'h3fb129a9, 32'h40048c79} /* (30, 15, 4) {real, imag} */,
  {32'hbec63898, 32'h3df43195} /* (30, 15, 3) {real, imag} */,
  {32'hc01d685a, 32'hbf1035ad} /* (30, 15, 2) {real, imag} */,
  {32'h3fed4cc6, 32'hbf86f184} /* (30, 15, 1) {real, imag} */,
  {32'h403cc802, 32'h3fc9221a} /* (30, 15, 0) {real, imag} */,
  {32'hc0819833, 32'h40940d7e} /* (30, 14, 31) {real, imag} */,
  {32'h3fc5d93d, 32'hc04e9c1d} /* (30, 14, 30) {real, imag} */,
  {32'h3ffcbf43, 32'h3f919b54} /* (30, 14, 29) {real, imag} */,
  {32'hc04ac1a3, 32'h40ae0cff} /* (30, 14, 28) {real, imag} */,
  {32'hbe4f082e, 32'hbfdb740a} /* (30, 14, 27) {real, imag} */,
  {32'h3f874b47, 32'hbf8b94cf} /* (30, 14, 26) {real, imag} */,
  {32'hbf5f0621, 32'hbd9115b9} /* (30, 14, 25) {real, imag} */,
  {32'h3fce23ee, 32'hc05d582c} /* (30, 14, 24) {real, imag} */,
  {32'h3e00b2ee, 32'h3f72030c} /* (30, 14, 23) {real, imag} */,
  {32'h3ed4d428, 32'hbf67edb7} /* (30, 14, 22) {real, imag} */,
  {32'hbd267e65, 32'hbf0e2d65} /* (30, 14, 21) {real, imag} */,
  {32'hbf97c1fe, 32'h3e374f27} /* (30, 14, 20) {real, imag} */,
  {32'h3fbdb3f7, 32'h3ffd256c} /* (30, 14, 19) {real, imag} */,
  {32'h3fc2d00f, 32'h3ecef339} /* (30, 14, 18) {real, imag} */,
  {32'h3f46311f, 32'hbf8a90e7} /* (30, 14, 17) {real, imag} */,
  {32'hbfcc525d, 32'hbeabfa8d} /* (30, 14, 16) {real, imag} */,
  {32'hbe3b1b0d, 32'h3f809acd} /* (30, 14, 15) {real, imag} */,
  {32'h3f9f1164, 32'hbf95fc4f} /* (30, 14, 14) {real, imag} */,
  {32'hc00baa15, 32'hbd9bafc8} /* (30, 14, 13) {real, imag} */,
  {32'h3fe3501d, 32'h3fc89809} /* (30, 14, 12) {real, imag} */,
  {32'h3f986ef5, 32'h3eabe36b} /* (30, 14, 11) {real, imag} */,
  {32'hbf970306, 32'hc0235455} /* (30, 14, 10) {real, imag} */,
  {32'h3e375f59, 32'hc020995b} /* (30, 14, 9) {real, imag} */,
  {32'h3f84a796, 32'hbf227935} /* (30, 14, 8) {real, imag} */,
  {32'h3f8c4433, 32'hbe91bfd9} /* (30, 14, 7) {real, imag} */,
  {32'h40144aac, 32'hbf7e1e67} /* (30, 14, 6) {real, imag} */,
  {32'h3fb93c7f, 32'h3fd757a5} /* (30, 14, 5) {real, imag} */,
  {32'h3ce1a10c, 32'h3fbe9973} /* (30, 14, 4) {real, imag} */,
  {32'h3f34918f, 32'hbe1f1117} /* (30, 14, 3) {real, imag} */,
  {32'h3ef7e8ab, 32'h3f999573} /* (30, 14, 2) {real, imag} */,
  {32'hc039f520, 32'hbfbd2dc4} /* (30, 14, 1) {real, imag} */,
  {32'hc051c253, 32'hbfd38a5d} /* (30, 14, 0) {real, imag} */,
  {32'h3f167f77, 32'hbf6fd0d9} /* (30, 13, 31) {real, imag} */,
  {32'h3c3a7e8b, 32'hbf0c9e01} /* (30, 13, 30) {real, imag} */,
  {32'hbf8d9f0f, 32'hbe9a720f} /* (30, 13, 29) {real, imag} */,
  {32'h3f9c36c9, 32'hc04fb744} /* (30, 13, 28) {real, imag} */,
  {32'h3ed760a5, 32'hc0181080} /* (30, 13, 27) {real, imag} */,
  {32'hc0663078, 32'hc06e35a3} /* (30, 13, 26) {real, imag} */,
  {32'hc0017bf5, 32'hbd811f65} /* (30, 13, 25) {real, imag} */,
  {32'hbf7225a6, 32'h3f8acfb0} /* (30, 13, 24) {real, imag} */,
  {32'h3fb63967, 32'hbf90f324} /* (30, 13, 23) {real, imag} */,
  {32'h3f558019, 32'hc0164741} /* (30, 13, 22) {real, imag} */,
  {32'h3c0fa1fb, 32'h3fabf2aa} /* (30, 13, 21) {real, imag} */,
  {32'h400af863, 32'hbe0c32f9} /* (30, 13, 20) {real, imag} */,
  {32'h3e020355, 32'h3e8d346d} /* (30, 13, 19) {real, imag} */,
  {32'h400ca525, 32'h3fbd6807} /* (30, 13, 18) {real, imag} */,
  {32'hbe207fe6, 32'h3f53daef} /* (30, 13, 17) {real, imag} */,
  {32'h4009719f, 32'hba8a8aa1} /* (30, 13, 16) {real, imag} */,
  {32'h3f6e3d1f, 32'hbe981ea9} /* (30, 13, 15) {real, imag} */,
  {32'hbf808ba9, 32'hc04d7bd5} /* (30, 13, 14) {real, imag} */,
  {32'h3e7955c6, 32'hbf3691ce} /* (30, 13, 13) {real, imag} */,
  {32'hbfde8cd1, 32'hbf82afc9} /* (30, 13, 12) {real, imag} */,
  {32'hbf6a1753, 32'h3f2181c4} /* (30, 13, 11) {real, imag} */,
  {32'hbf2594ea, 32'h3d415764} /* (30, 13, 10) {real, imag} */,
  {32'h3fad5921, 32'h3f7f5e28} /* (30, 13, 9) {real, imag} */,
  {32'hc001d2f1, 32'h3ed6ba79} /* (30, 13, 8) {real, imag} */,
  {32'hbf98f65e, 32'hc07fcefa} /* (30, 13, 7) {real, imag} */,
  {32'hbfa33dcf, 32'h4000a268} /* (30, 13, 6) {real, imag} */,
  {32'hbf347e71, 32'h40105b3c} /* (30, 13, 5) {real, imag} */,
  {32'h3fad63c0, 32'hc01a8e24} /* (30, 13, 4) {real, imag} */,
  {32'hbf18dde4, 32'h3efe5ffa} /* (30, 13, 3) {real, imag} */,
  {32'hbe4aa8c2, 32'h3f85c364} /* (30, 13, 2) {real, imag} */,
  {32'h4027c2bf, 32'hc08de4f8} /* (30, 13, 1) {real, imag} */,
  {32'h4024e6a6, 32'hbf62951e} /* (30, 13, 0) {real, imag} */,
  {32'h4041e90d, 32'h3f45d973} /* (30, 12, 31) {real, imag} */,
  {32'h400f9ab1, 32'hbe4e5192} /* (30, 12, 30) {real, imag} */,
  {32'hbdd920d6, 32'h3f1023bb} /* (30, 12, 29) {real, imag} */,
  {32'hbf0ce45a, 32'hbece7084} /* (30, 12, 28) {real, imag} */,
  {32'h3f49aed2, 32'h3fd5a8cc} /* (30, 12, 27) {real, imag} */,
  {32'hbfaa89f7, 32'hbfaee495} /* (30, 12, 26) {real, imag} */,
  {32'hbe22386b, 32'hbdfd29f3} /* (30, 12, 25) {real, imag} */,
  {32'h40144552, 32'h3f9416e1} /* (30, 12, 24) {real, imag} */,
  {32'hc0404ab5, 32'h3fec11f4} /* (30, 12, 23) {real, imag} */,
  {32'hbf45576f, 32'hbf480a09} /* (30, 12, 22) {real, imag} */,
  {32'h3db5c9d1, 32'h3e4f6297} /* (30, 12, 21) {real, imag} */,
  {32'h3f48252b, 32'h404e2a35} /* (30, 12, 20) {real, imag} */,
  {32'h3f803f17, 32'hbeb969b8} /* (30, 12, 19) {real, imag} */,
  {32'hbed449eb, 32'h3fea7604} /* (30, 12, 18) {real, imag} */,
  {32'hc016a76f, 32'h3f903f42} /* (30, 12, 17) {real, imag} */,
  {32'hbea27dd6, 32'h3d5e071b} /* (30, 12, 16) {real, imag} */,
  {32'h3e3b7ffe, 32'hbe7717d1} /* (30, 12, 15) {real, imag} */,
  {32'hbf184a9e, 32'h403ebb59} /* (30, 12, 14) {real, imag} */,
  {32'hbfeb9f85, 32'hbfe3d686} /* (30, 12, 13) {real, imag} */,
  {32'hc01ad6b7, 32'h3f96e081} /* (30, 12, 12) {real, imag} */,
  {32'h3f8367aa, 32'hbfa6ada0} /* (30, 12, 11) {real, imag} */,
  {32'h3f7b2998, 32'hc02d0035} /* (30, 12, 10) {real, imag} */,
  {32'hbf166e1a, 32'h40b0ba38} /* (30, 12, 9) {real, imag} */,
  {32'h3f10e1b9, 32'hbf3cd8d9} /* (30, 12, 8) {real, imag} */,
  {32'hbf97ea64, 32'h3f315d5e} /* (30, 12, 7) {real, imag} */,
  {32'h3dc9fff4, 32'hc024c2fd} /* (30, 12, 6) {real, imag} */,
  {32'h3d5ab544, 32'hbfb682e5} /* (30, 12, 5) {real, imag} */,
  {32'hbfa1da36, 32'hbfc38145} /* (30, 12, 4) {real, imag} */,
  {32'h4003f506, 32'hbfd5646f} /* (30, 12, 3) {real, imag} */,
  {32'hbfef002e, 32'hbe60a826} /* (30, 12, 2) {real, imag} */,
  {32'h3f830da1, 32'h3f64442d} /* (30, 12, 1) {real, imag} */,
  {32'hc0188b30, 32'hc03abde7} /* (30, 12, 0) {real, imag} */,
  {32'hc0d83fd2, 32'h40fd7c8f} /* (30, 11, 31) {real, imag} */,
  {32'h40161f93, 32'hc000055f} /* (30, 11, 30) {real, imag} */,
  {32'hbfc382f3, 32'hc080ca19} /* (30, 11, 29) {real, imag} */,
  {32'h4051feca, 32'h3d1ed3b3} /* (30, 11, 28) {real, imag} */,
  {32'h401b59f1, 32'hc042d322} /* (30, 11, 27) {real, imag} */,
  {32'h3f9909d3, 32'h403abf95} /* (30, 11, 26) {real, imag} */,
  {32'hbfbbf7e2, 32'hbf2a9c4d} /* (30, 11, 25) {real, imag} */,
  {32'hbe152fa2, 32'hc071c05e} /* (30, 11, 24) {real, imag} */,
  {32'h3f52bea4, 32'hbfa3ae8f} /* (30, 11, 23) {real, imag} */,
  {32'h3fd1c944, 32'h3fad667b} /* (30, 11, 22) {real, imag} */,
  {32'h3f653a69, 32'hc05f38dd} /* (30, 11, 21) {real, imag} */,
  {32'hbf9a3255, 32'h3fc54290} /* (30, 11, 20) {real, imag} */,
  {32'hbf361a24, 32'hbe8c92ac} /* (30, 11, 19) {real, imag} */,
  {32'h3e85e50a, 32'hbe683e83} /* (30, 11, 18) {real, imag} */,
  {32'h401df63e, 32'h3ef08ec5} /* (30, 11, 17) {real, imag} */,
  {32'hc02c0bcf, 32'h3fb3676b} /* (30, 11, 16) {real, imag} */,
  {32'hbea223ca, 32'hbeca8b92} /* (30, 11, 15) {real, imag} */,
  {32'hbf2afb14, 32'h3f77d69a} /* (30, 11, 14) {real, imag} */,
  {32'h3f86bad5, 32'h3d590e49} /* (30, 11, 13) {real, imag} */,
  {32'hc06e3e5c, 32'hbc23d8d9} /* (30, 11, 12) {real, imag} */,
  {32'h3ff61c0f, 32'hbff6a365} /* (30, 11, 11) {real, imag} */,
  {32'h405ad45e, 32'hc0c3f160} /* (30, 11, 10) {real, imag} */,
  {32'hbfc0ad53, 32'hbffce433} /* (30, 11, 9) {real, imag} */,
  {32'h406546bd, 32'hbe96d5c4} /* (30, 11, 8) {real, imag} */,
  {32'hbef1ead0, 32'hc00c3875} /* (30, 11, 7) {real, imag} */,
  {32'h3fe2611d, 32'h400a8cb7} /* (30, 11, 6) {real, imag} */,
  {32'h408e3ba2, 32'hc00511be} /* (30, 11, 5) {real, imag} */,
  {32'hbfb8da4c, 32'hbfbc551d} /* (30, 11, 4) {real, imag} */,
  {32'hbf2e1987, 32'hc01023f8} /* (30, 11, 3) {real, imag} */,
  {32'h40b6f6bf, 32'hbf54f47d} /* (30, 11, 2) {real, imag} */,
  {32'hc11634fd, 32'h40a70247} /* (30, 11, 1) {real, imag} */,
  {32'hc087d318, 32'h41142422} /* (30, 11, 0) {real, imag} */,
  {32'h40edf53b, 32'h4010c10c} /* (30, 10, 31) {real, imag} */,
  {32'hbf36eab4, 32'hc01f84ca} /* (30, 10, 30) {real, imag} */,
  {32'h404154b9, 32'hbfc513ca} /* (30, 10, 29) {real, imag} */,
  {32'hbfda24c3, 32'hbf0077d1} /* (30, 10, 28) {real, imag} */,
  {32'hbf330c93, 32'h405e96a0} /* (30, 10, 27) {real, imag} */,
  {32'hbf1edca7, 32'h4017460f} /* (30, 10, 26) {real, imag} */,
  {32'h3ffee535, 32'h40080e2b} /* (30, 10, 25) {real, imag} */,
  {32'hbf9ed3a4, 32'h403843ca} /* (30, 10, 24) {real, imag} */,
  {32'h3db9be4b, 32'h3d8e55e5} /* (30, 10, 23) {real, imag} */,
  {32'hbfaebed2, 32'hbfd1c02f} /* (30, 10, 22) {real, imag} */,
  {32'hc0624645, 32'hbfcf80a3} /* (30, 10, 21) {real, imag} */,
  {32'hbf1e2bd6, 32'h3ea57529} /* (30, 10, 20) {real, imag} */,
  {32'h401def0d, 32'hbf13c16c} /* (30, 10, 19) {real, imag} */,
  {32'h3fed0775, 32'hbf879a89} /* (30, 10, 18) {real, imag} */,
  {32'h3f6a7b94, 32'hbfd81380} /* (30, 10, 17) {real, imag} */,
  {32'h3fe302b1, 32'h4003d098} /* (30, 10, 16) {real, imag} */,
  {32'h3f0261cc, 32'h3f3e72b9} /* (30, 10, 15) {real, imag} */,
  {32'hbff030f7, 32'hbee4d820} /* (30, 10, 14) {real, imag} */,
  {32'hbfa26805, 32'hc016608f} /* (30, 10, 13) {real, imag} */,
  {32'hc01e31c8, 32'h3f7a67c0} /* (30, 10, 12) {real, imag} */,
  {32'h3f7926ce, 32'h40032794} /* (30, 10, 11) {real, imag} */,
  {32'h4011b23f, 32'h3ff5dc9c} /* (30, 10, 10) {real, imag} */,
  {32'hbd8b9551, 32'hc003df4f} /* (30, 10, 9) {real, imag} */,
  {32'hc01bd342, 32'h3fc24fb5} /* (30, 10, 8) {real, imag} */,
  {32'hbf81f3c4, 32'hbf318ace} /* (30, 10, 7) {real, imag} */,
  {32'hbea6e9ce, 32'hc087ab9c} /* (30, 10, 6) {real, imag} */,
  {32'hbec3f03b, 32'hc0234dca} /* (30, 10, 5) {real, imag} */,
  {32'h402ce9c2, 32'hbffac0c9} /* (30, 10, 4) {real, imag} */,
  {32'h3f9bda61, 32'hbf89f92e} /* (30, 10, 3) {real, imag} */,
  {32'hc0524f54, 32'h40c8bcf9} /* (30, 10, 2) {real, imag} */,
  {32'h402067ee, 32'hc0af85d4} /* (30, 10, 1) {real, imag} */,
  {32'h401e1d87, 32'hbed9ff22} /* (30, 10, 0) {real, imag} */,
  {32'h403cc6c1, 32'h40d871fc} /* (30, 9, 31) {real, imag} */,
  {32'hc0e5553c, 32'h3f9546d4} /* (30, 9, 30) {real, imag} */,
  {32'h4042ff08, 32'hbe2cbe72} /* (30, 9, 29) {real, imag} */,
  {32'h3fe8f894, 32'hc013d56a} /* (30, 9, 28) {real, imag} */,
  {32'hbfd18ba2, 32'h3e82b654} /* (30, 9, 27) {real, imag} */,
  {32'h4072dca3, 32'h4004fa01} /* (30, 9, 26) {real, imag} */,
  {32'h3f5b71b7, 32'hbf441f96} /* (30, 9, 25) {real, imag} */,
  {32'hbf96fcc7, 32'h3fa6bdf0} /* (30, 9, 24) {real, imag} */,
  {32'h3ff1bb0f, 32'hbfb7a355} /* (30, 9, 23) {real, imag} */,
  {32'hc00697b3, 32'h407cea2f} /* (30, 9, 22) {real, imag} */,
  {32'h3fc2820a, 32'h40333c39} /* (30, 9, 21) {real, imag} */,
  {32'hc0586504, 32'hc02dfbdd} /* (30, 9, 20) {real, imag} */,
  {32'hbf639d48, 32'hc07a5b1d} /* (30, 9, 19) {real, imag} */,
  {32'h3f6fac7e, 32'hc01a3bdf} /* (30, 9, 18) {real, imag} */,
  {32'h3fc0eefd, 32'hbed820ee} /* (30, 9, 17) {real, imag} */,
  {32'h3fdbb862, 32'h3f1a24b7} /* (30, 9, 16) {real, imag} */,
  {32'hbfae2354, 32'h3f8fb503} /* (30, 9, 15) {real, imag} */,
  {32'hbf1b88f5, 32'hbfdb43b0} /* (30, 9, 14) {real, imag} */,
  {32'h4027ea93, 32'h4024e155} /* (30, 9, 13) {real, imag} */,
  {32'hbefb7c7f, 32'hbf7dcb42} /* (30, 9, 12) {real, imag} */,
  {32'hc0434cfd, 32'hbe5fee32} /* (30, 9, 11) {real, imag} */,
  {32'hbf957808, 32'h4058f46d} /* (30, 9, 10) {real, imag} */,
  {32'h3fe4181b, 32'hbf7fcba9} /* (30, 9, 9) {real, imag} */,
  {32'hc0a95a81, 32'h3f35b6fe} /* (30, 9, 8) {real, imag} */,
  {32'h3fb0cd85, 32'hbd8a4d7d} /* (30, 9, 7) {real, imag} */,
  {32'h3f1b2971, 32'hbfe8a3f1} /* (30, 9, 6) {real, imag} */,
  {32'h404371d9, 32'hc01c770e} /* (30, 9, 5) {real, imag} */,
  {32'h40b4c74b, 32'h3e9b86a6} /* (30, 9, 4) {real, imag} */,
  {32'hc0efe04f, 32'h3fff1d3a} /* (30, 9, 3) {real, imag} */,
  {32'hc0bdf112, 32'h3ec35aff} /* (30, 9, 2) {real, imag} */,
  {32'h40dae08a, 32'hc0d349c8} /* (30, 9, 1) {real, imag} */,
  {32'h3f80f19a, 32'hbb8ff004} /* (30, 9, 0) {real, imag} */,
  {32'hc14b4257, 32'h41d1e713} /* (30, 8, 31) {real, imag} */,
  {32'hc0446717, 32'hc14d5f80} /* (30, 8, 30) {real, imag} */,
  {32'hc0aec216, 32'hbfa60cd1} /* (30, 8, 29) {real, imag} */,
  {32'hc00cdcc6, 32'h3f7c7aef} /* (30, 8, 28) {real, imag} */,
  {32'h4028d0d0, 32'hc0051b57} /* (30, 8, 27) {real, imag} */,
  {32'h3dcd6d0a, 32'h40822c24} /* (30, 8, 26) {real, imag} */,
  {32'hc08317a4, 32'h3fd22a32} /* (30, 8, 25) {real, imag} */,
  {32'hbfd0148f, 32'hbfb0463e} /* (30, 8, 24) {real, imag} */,
  {32'hbcc6f69c, 32'h4043fa8b} /* (30, 8, 23) {real, imag} */,
  {32'h3be8df56, 32'hc0d389f4} /* (30, 8, 22) {real, imag} */,
  {32'hbf37e79f, 32'hc0676381} /* (30, 8, 21) {real, imag} */,
  {32'hbd5ad07f, 32'hc02eb31a} /* (30, 8, 20) {real, imag} */,
  {32'h3f5aaa70, 32'hbcb30945} /* (30, 8, 19) {real, imag} */,
  {32'h3f6958db, 32'hbdc5f7eb} /* (30, 8, 18) {real, imag} */,
  {32'h3fe17cab, 32'hbf4f63af} /* (30, 8, 17) {real, imag} */,
  {32'hbf35f79b, 32'h3e14305f} /* (30, 8, 16) {real, imag} */,
  {32'hbec4b6de, 32'h3e1429a9} /* (30, 8, 15) {real, imag} */,
  {32'h3e963049, 32'h3c35f2d2} /* (30, 8, 14) {real, imag} */,
  {32'h3f6df20d, 32'h3e4e80a3} /* (30, 8, 13) {real, imag} */,
  {32'h3fe7d96a, 32'h3f9b98c4} /* (30, 8, 12) {real, imag} */,
  {32'h3ffea7ee, 32'hbfc87bd5} /* (30, 8, 11) {real, imag} */,
  {32'hc05fd871, 32'hbc836b41} /* (30, 8, 10) {real, imag} */,
  {32'hbf0bf646, 32'h3dace64b} /* (30, 8, 9) {real, imag} */,
  {32'h400b8f47, 32'hc01068ad} /* (30, 8, 8) {real, imag} */,
  {32'hc050fe38, 32'hbf7923c6} /* (30, 8, 7) {real, imag} */,
  {32'h3fadc060, 32'hc04ac2b4} /* (30, 8, 6) {real, imag} */,
  {32'h40cf66e5, 32'hc0a13f24} /* (30, 8, 5) {real, imag} */,
  {32'hc00541e7, 32'h40c45195} /* (30, 8, 4) {real, imag} */,
  {32'h3f44582d, 32'h3f07b39f} /* (30, 8, 3) {real, imag} */,
  {32'h4086c307, 32'hc0c036a3} /* (30, 8, 2) {real, imag} */,
  {32'hc103c893, 32'h414d30fa} /* (30, 8, 1) {real, imag} */,
  {32'hc0141188, 32'h41585f96} /* (30, 8, 0) {real, imag} */,
  {32'h409d099d, 32'hc06de482} /* (30, 7, 31) {real, imag} */,
  {32'hbfb05b43, 32'h3fa0895a} /* (30, 7, 30) {real, imag} */,
  {32'hbf317449, 32'hbfe9fd1c} /* (30, 7, 29) {real, imag} */,
  {32'hbfc8589e, 32'h40588919} /* (30, 7, 28) {real, imag} */,
  {32'h3f60cf7f, 32'h3f8cecab} /* (30, 7, 27) {real, imag} */,
  {32'h3fcb83ca, 32'hbf2d80c7} /* (30, 7, 26) {real, imag} */,
  {32'hbe940ca3, 32'hbfcd007a} /* (30, 7, 25) {real, imag} */,
  {32'hbfb65369, 32'h40390a79} /* (30, 7, 24) {real, imag} */,
  {32'hc002b430, 32'h3f9fed16} /* (30, 7, 23) {real, imag} */,
  {32'h3fa5b05d, 32'hbfb79661} /* (30, 7, 22) {real, imag} */,
  {32'hbe9c68da, 32'h3eaa2c27} /* (30, 7, 21) {real, imag} */,
  {32'hbeebc2a7, 32'hbf6be4c8} /* (30, 7, 20) {real, imag} */,
  {32'h3fe53981, 32'hc0b639a8} /* (30, 7, 19) {real, imag} */,
  {32'h3fa5eeb8, 32'h40365c4e} /* (30, 7, 18) {real, imag} */,
  {32'hbf633a9a, 32'h40132e0c} /* (30, 7, 17) {real, imag} */,
  {32'h404db097, 32'h3fd9263f} /* (30, 7, 16) {real, imag} */,
  {32'hbf02a778, 32'hbfa4d687} /* (30, 7, 15) {real, imag} */,
  {32'h3f0ee549, 32'hbf91924d} /* (30, 7, 14) {real, imag} */,
  {32'hc02cd315, 32'hbe46d0db} /* (30, 7, 13) {real, imag} */,
  {32'h3f1c0a62, 32'h3e7f6c42} /* (30, 7, 12) {real, imag} */,
  {32'h3e4d70cb, 32'hc0094139} /* (30, 7, 11) {real, imag} */,
  {32'h3e93d9f0, 32'h3fe76b22} /* (30, 7, 10) {real, imag} */,
  {32'hc02007eb, 32'h3f4b65de} /* (30, 7, 9) {real, imag} */,
  {32'hc021cd31, 32'hc035456d} /* (30, 7, 8) {real, imag} */,
  {32'hbf44fa0e, 32'hbe35d3fe} /* (30, 7, 7) {real, imag} */,
  {32'hc09f42e2, 32'hbfdf6b29} /* (30, 7, 6) {real, imag} */,
  {32'hc08c1e31, 32'h405dc5dd} /* (30, 7, 5) {real, imag} */,
  {32'hbe8e4c8c, 32'h4000cd59} /* (30, 7, 4) {real, imag} */,
  {32'hbf971acd, 32'hc045bb99} /* (30, 7, 3) {real, imag} */,
  {32'hbff72b1a, 32'hbe8c437b} /* (30, 7, 2) {real, imag} */,
  {32'h4116344d, 32'hc09cb3fa} /* (30, 7, 1) {real, imag} */,
  {32'h410132a3, 32'hc07580f2} /* (30, 7, 0) {real, imag} */,
  {32'hc0ab581b, 32'h40cfaf15} /* (30, 6, 31) {real, imag} */,
  {32'hbeeca322, 32'hc07cd97b} /* (30, 6, 30) {real, imag} */,
  {32'hbfb39035, 32'hc0934042} /* (30, 6, 29) {real, imag} */,
  {32'hc1082d4b, 32'h3f7ffdf3} /* (30, 6, 28) {real, imag} */,
  {32'h3e42bb59, 32'hbfedf71c} /* (30, 6, 27) {real, imag} */,
  {32'h40dfd167, 32'hc0285a08} /* (30, 6, 26) {real, imag} */,
  {32'h3ee0afa2, 32'hbf74096a} /* (30, 6, 25) {real, imag} */,
  {32'h40533e14, 32'hbf8a23d2} /* (30, 6, 24) {real, imag} */,
  {32'hbf38d4c1, 32'hc0868cf5} /* (30, 6, 23) {real, imag} */,
  {32'h3f4552a2, 32'hbf204697} /* (30, 6, 22) {real, imag} */,
  {32'h3fb2f880, 32'hc01c30e8} /* (30, 6, 21) {real, imag} */,
  {32'hbfde9023, 32'h3fe520e5} /* (30, 6, 20) {real, imag} */,
  {32'hbf269f85, 32'hbff8603c} /* (30, 6, 19) {real, imag} */,
  {32'hbd3554cf, 32'hbfe6bcef} /* (30, 6, 18) {real, imag} */,
  {32'h3f7ecd65, 32'hbf383201} /* (30, 6, 17) {real, imag} */,
  {32'h40104f9c, 32'h3f26f9d3} /* (30, 6, 16) {real, imag} */,
  {32'hbf8b6022, 32'hbf22f123} /* (30, 6, 15) {real, imag} */,
  {32'hbf81ecea, 32'hbef75bfa} /* (30, 6, 14) {real, imag} */,
  {32'h3f341a9e, 32'hbf8d1a94} /* (30, 6, 13) {real, imag} */,
  {32'h3f9d4690, 32'hbe14d980} /* (30, 6, 12) {real, imag} */,
  {32'h3f891814, 32'hc0145d13} /* (30, 6, 11) {real, imag} */,
  {32'hbf9152c7, 32'h3ec5c348} /* (30, 6, 10) {real, imag} */,
  {32'hc038f59b, 32'h401ac9e3} /* (30, 6, 9) {real, imag} */,
  {32'hbfac4e54, 32'hc04f757f} /* (30, 6, 8) {real, imag} */,
  {32'h3f89ed43, 32'hbf0d0a17} /* (30, 6, 7) {real, imag} */,
  {32'hbff1eee6, 32'hbd583b31} /* (30, 6, 6) {real, imag} */,
  {32'hc00ea5dc, 32'hc0c639e6} /* (30, 6, 5) {real, imag} */,
  {32'hc02423f4, 32'h402631ea} /* (30, 6, 4) {real, imag} */,
  {32'h40a52d29, 32'h400ab742} /* (30, 6, 3) {real, imag} */,
  {32'h400ba8e4, 32'hc0df54e4} /* (30, 6, 2) {real, imag} */,
  {32'hbfbbbb74, 32'h3f383793} /* (30, 6, 1) {real, imag} */,
  {32'h400ee842, 32'hc01f88dd} /* (30, 6, 0) {real, imag} */,
  {32'hbfb52aa4, 32'h42430ab8} /* (30, 5, 31) {real, imag} */,
  {32'hc0d6a900, 32'hc16ce489} /* (30, 5, 30) {real, imag} */,
  {32'hc0828427, 32'h403ae6bd} /* (30, 5, 29) {real, imag} */,
  {32'h41263bef, 32'h3fa41740} /* (30, 5, 28) {real, imag} */,
  {32'h41018ed1, 32'hc10c01f0} /* (30, 5, 27) {real, imag} */,
  {32'hc05e7122, 32'hc03d15bd} /* (30, 5, 26) {real, imag} */,
  {32'hc046458f, 32'h4053e3f9} /* (30, 5, 25) {real, imag} */,
  {32'hc077c079, 32'hbfca8aad} /* (30, 5, 24) {real, imag} */,
  {32'h3f05603b, 32'h3db55d5a} /* (30, 5, 23) {real, imag} */,
  {32'hbf22efd5, 32'hc0bf93dd} /* (30, 5, 22) {real, imag} */,
  {32'hc0703673, 32'hbf9069a8} /* (30, 5, 21) {real, imag} */,
  {32'hbf4d7003, 32'hbf3ac034} /* (30, 5, 20) {real, imag} */,
  {32'h3f98e479, 32'hc001d2a9} /* (30, 5, 19) {real, imag} */,
  {32'hbfd9c08a, 32'h3fc23917} /* (30, 5, 18) {real, imag} */,
  {32'hbecabed2, 32'h3e3e83b4} /* (30, 5, 17) {real, imag} */,
  {32'hc0167def, 32'h3f800322} /* (30, 5, 16) {real, imag} */,
  {32'h400d84ed, 32'hbe52e36d} /* (30, 5, 15) {real, imag} */,
  {32'h403e4f88, 32'h3f5918c9} /* (30, 5, 14) {real, imag} */,
  {32'h3fe19cd7, 32'h400646dc} /* (30, 5, 13) {real, imag} */,
  {32'h3faa924b, 32'hbf9ba8a7} /* (30, 5, 12) {real, imag} */,
  {32'h4081403c, 32'h3f89dce2} /* (30, 5, 11) {real, imag} */,
  {32'hbf83f3f3, 32'h3f1ff5e1} /* (30, 5, 10) {real, imag} */,
  {32'h3faf5049, 32'hbf2c3552} /* (30, 5, 9) {real, imag} */,
  {32'h3ef73f07, 32'h401c649f} /* (30, 5, 8) {real, imag} */,
  {32'hbfdfe2be, 32'h400fa790} /* (30, 5, 7) {real, imag} */,
  {32'h40733d33, 32'hc0061f0e} /* (30, 5, 6) {real, imag} */,
  {32'hbf5fd5a8, 32'hc108ab9a} /* (30, 5, 5) {real, imag} */,
  {32'hc0546cb6, 32'hc0041a87} /* (30, 5, 4) {real, imag} */,
  {32'hc09490dc, 32'h40a33c4e} /* (30, 5, 3) {real, imag} */,
  {32'h41377ad8, 32'hc12bb034} /* (30, 5, 2) {real, imag} */,
  {32'hc20d9a00, 32'h4223aa24} /* (30, 5, 1) {real, imag} */,
  {32'hc10f778f, 32'h420a52cb} /* (30, 5, 0) {real, imag} */,
  {32'h42275d2f, 32'hc209eaa5} /* (30, 4, 31) {real, imag} */,
  {32'hc1ffefef, 32'h4225b0ce} /* (30, 4, 30) {real, imag} */,
  {32'hbf980553, 32'h3fd32861} /* (30, 4, 29) {real, imag} */,
  {32'h40011c6a, 32'hc1370ca3} /* (30, 4, 28) {real, imag} */,
  {32'h40850ebc, 32'h414b986a} /* (30, 4, 27) {real, imag} */,
  {32'h40c46e43, 32'hbfa9b31c} /* (30, 4, 26) {real, imag} */,
  {32'hbffd56c5, 32'h3e103e98} /* (30, 4, 25) {real, imag} */,
  {32'hbfc32460, 32'h4000d33f} /* (30, 4, 24) {real, imag} */,
  {32'hc0969cb8, 32'hbff274a8} /* (30, 4, 23) {real, imag} */,
  {32'hbfc0efa1, 32'hbf114708} /* (30, 4, 22) {real, imag} */,
  {32'h40838147, 32'h40a21e4c} /* (30, 4, 21) {real, imag} */,
  {32'hc08f4a4b, 32'hc0598d7b} /* (30, 4, 20) {real, imag} */,
  {32'hbf14a898, 32'hbf43133f} /* (30, 4, 19) {real, imag} */,
  {32'hbdb29236, 32'h406b5298} /* (30, 4, 18) {real, imag} */,
  {32'hbf166b92, 32'hc00cfca8} /* (30, 4, 17) {real, imag} */,
  {32'hbe6985b0, 32'hbfbcbfad} /* (30, 4, 16) {real, imag} */,
  {32'h402cc952, 32'h3f6760dc} /* (30, 4, 15) {real, imag} */,
  {32'hc079075d, 32'h3fb7d87d} /* (30, 4, 14) {real, imag} */,
  {32'h3eb27d7d, 32'h3e1a6413} /* (30, 4, 13) {real, imag} */,
  {32'h3ee5f52b, 32'hbfe99149} /* (30, 4, 12) {real, imag} */,
  {32'hbfbb2b8e, 32'hbf137266} /* (30, 4, 11) {real, imag} */,
  {32'h40a54489, 32'h3ffc9286} /* (30, 4, 10) {real, imag} */,
  {32'h4011c8dc, 32'h3faba89a} /* (30, 4, 9) {real, imag} */,
  {32'hc0899c17, 32'h40baa25c} /* (30, 4, 8) {real, imag} */,
  {32'h401474ef, 32'hc051069c} /* (30, 4, 7) {real, imag} */,
  {32'h3f0c4fe9, 32'h3f966e0c} /* (30, 4, 6) {real, imag} */,
  {32'hc1498394, 32'h40347a7c} /* (30, 4, 5) {real, imag} */,
  {32'h3f828e05, 32'h40566f0e} /* (30, 4, 4) {real, imag} */,
  {32'h404ed4f1, 32'hc03bda0a} /* (30, 4, 3) {real, imag} */,
  {32'hc1dfbd95, 32'h424e6be5} /* (30, 4, 2) {real, imag} */,
  {32'h4175143c, 32'hc2a5023a} /* (30, 4, 1) {real, imag} */,
  {32'h3ee369fa, 32'hc1ebd48a} /* (30, 4, 0) {real, imag} */,
  {32'h425b74d8, 32'h42638df0} /* (30, 3, 31) {real, imag} */,
  {32'hc24c371c, 32'hc14b8448} /* (30, 3, 30) {real, imag} */,
  {32'h3fd87d79, 32'hc05f7f8b} /* (30, 3, 29) {real, imag} */,
  {32'h4102690d, 32'hc1558dd1} /* (30, 3, 28) {real, imag} */,
  {32'h408a97f6, 32'h40dc955f} /* (30, 3, 27) {real, imag} */,
  {32'h4090069a, 32'hc0891573} /* (30, 3, 26) {real, imag} */,
  {32'hbd82f28d, 32'hbf968ceb} /* (30, 3, 25) {real, imag} */,
  {32'hc0d38e5a, 32'h408d7dfe} /* (30, 3, 24) {real, imag} */,
  {32'h3ff02b19, 32'hbe488e19} /* (30, 3, 23) {real, imag} */,
  {32'h40b0f982, 32'hbff7436a} /* (30, 3, 22) {real, imag} */,
  {32'hbe7d8f60, 32'h3d64b515} /* (30, 3, 21) {real, imag} */,
  {32'hbfbbaf96, 32'h403f77c3} /* (30, 3, 20) {real, imag} */,
  {32'hc08e5650, 32'h3f91cf40} /* (30, 3, 19) {real, imag} */,
  {32'hc010b8a6, 32'hbf84f826} /* (30, 3, 18) {real, imag} */,
  {32'h3f0f198c, 32'hbec7404d} /* (30, 3, 17) {real, imag} */,
  {32'hbf7850ed, 32'h3d733db1} /* (30, 3, 16) {real, imag} */,
  {32'h3eee5477, 32'hbfccc76a} /* (30, 3, 15) {real, imag} */,
  {32'hc01fe22e, 32'h3f9e4649} /* (30, 3, 14) {real, imag} */,
  {32'hbf811ef4, 32'hbe9f15a9} /* (30, 3, 13) {real, imag} */,
  {32'hbf51984e, 32'h400f0d6e} /* (30, 3, 12) {real, imag} */,
  {32'h3fd3017f, 32'hc0280b06} /* (30, 3, 11) {real, imag} */,
  {32'h3f0e56ae, 32'h3e71b180} /* (30, 3, 10) {real, imag} */,
  {32'h3ed00f30, 32'hbe83ec3c} /* (30, 3, 9) {real, imag} */,
  {32'hbebe3edd, 32'hc0880148} /* (30, 3, 8) {real, imag} */,
  {32'h40b2bb25, 32'hc02a185c} /* (30, 3, 7) {real, imag} */,
  {32'h401c68de, 32'h3e548867} /* (30, 3, 6) {real, imag} */,
  {32'h3f16ca90, 32'h4026b9c5} /* (30, 3, 5) {real, imag} */,
  {32'h413d366f, 32'h4198c15d} /* (30, 3, 4) {real, imag} */,
  {32'h415fa31a, 32'hc097a24d} /* (30, 3, 3) {real, imag} */,
  {32'hc24dc073, 32'h414ebf45} /* (30, 3, 2) {real, imag} */,
  {32'h420f5519, 32'hc28b2aea} /* (30, 3, 1) {real, imag} */,
  {32'hc130fc6f, 32'h3fb71427} /* (30, 3, 0) {real, imag} */,
  {32'h42b01dd2, 32'h43ddbab4} /* (30, 2, 31) {real, imag} */,
  {32'hc2f4b5f1, 32'hc359f467} /* (30, 2, 30) {real, imag} */,
  {32'h410f371c, 32'h3febe84c} /* (30, 2, 29) {real, imag} */,
  {32'h42170128, 32'h41905b99} /* (30, 2, 28) {real, imag} */,
  {32'hc1cb41b3, 32'hc1581812} /* (30, 2, 27) {real, imag} */,
  {32'hc02f33ca, 32'hc0a7683c} /* (30, 2, 26) {real, imag} */,
  {32'h413d7688, 32'h40001b9d} /* (30, 2, 25) {real, imag} */,
  {32'hc1b859c7, 32'hc12fa83a} /* (30, 2, 24) {real, imag} */,
  {32'hbf5f8718, 32'hc009e7fb} /* (30, 2, 23) {real, imag} */,
  {32'h40046152, 32'hbe7d2a0e} /* (30, 2, 22) {real, imag} */,
  {32'hc1194fd8, 32'hbf5c6638} /* (30, 2, 21) {real, imag} */,
  {32'hbea260df, 32'h4075d5ec} /* (30, 2, 20) {real, imag} */,
  {32'hbd67eb86, 32'hbf392de4} /* (30, 2, 19) {real, imag} */,
  {32'hc040907e, 32'hc00c3f86} /* (30, 2, 18) {real, imag} */,
  {32'h4088cfe2, 32'hbefa9d54} /* (30, 2, 17) {real, imag} */,
  {32'h3fa4594b, 32'hc0082653} /* (30, 2, 16) {real, imag} */,
  {32'hbf6e0795, 32'h3fdc31f2} /* (30, 2, 15) {real, imag} */,
  {32'h40ae8274, 32'hbfd6e77e} /* (30, 2, 14) {real, imag} */,
  {32'hbee2b415, 32'h3f8e3691} /* (30, 2, 13) {real, imag} */,
  {32'h3e5a3e1b, 32'h3fc3c554} /* (30, 2, 12) {real, imag} */,
  {32'h40c2724c, 32'hc03d34a1} /* (30, 2, 11) {real, imag} */,
  {32'hc056f322, 32'h40ac9f26} /* (30, 2, 10) {real, imag} */,
  {32'hc0361ebd, 32'h3fdad88c} /* (30, 2, 9) {real, imag} */,
  {32'h41054c07, 32'hc163ceec} /* (30, 2, 8) {real, imag} */,
  {32'h400b45ac, 32'h4069f3c3} /* (30, 2, 7) {real, imag} */,
  {32'h3cea1769, 32'h4086813e} /* (30, 2, 6) {real, imag} */,
  {32'h41e1e526, 32'hc1e8055c} /* (30, 2, 5) {real, imag} */,
  {32'h406a5d3b, 32'h4218f3d9} /* (30, 2, 4) {real, imag} */,
  {32'h40588da8, 32'hc048bf4e} /* (30, 2, 3) {real, imag} */,
  {32'hc2c3eebb, 32'hc30de680} /* (30, 2, 2) {real, imag} */,
  {32'h42b31a1f, 32'h4373a611} /* (30, 2, 1) {real, imag} */,
  {32'h40e32513, 32'h437acf45} /* (30, 2, 0) {real, imag} */,
  {32'hc363a405, 32'hc3ffa953} /* (30, 1, 31) {real, imag} */,
  {32'h41cb8a6c, 32'h4307b885} /* (30, 1, 30) {real, imag} */,
  {32'h41356100, 32'h41a7a084} /* (30, 1, 29) {real, imag} */,
  {32'h41c155f6, 32'hc24df572} /* (30, 1, 28) {real, imag} */,
  {32'h41823857, 32'h42740455} /* (30, 1, 27) {real, imag} */,
  {32'h41409e32, 32'h40be798d} /* (30, 1, 26) {real, imag} */,
  {32'hc0a5e6b7, 32'hc093b168} /* (30, 1, 25) {real, imag} */,
  {32'h4127ee15, 32'h40afc6a7} /* (30, 1, 24) {real, imag} */,
  {32'hbee60919, 32'h4067ab3a} /* (30, 1, 23) {real, imag} */,
  {32'h3f098a48, 32'hbeb21c95} /* (30, 1, 22) {real, imag} */,
  {32'h411efae8, 32'h40b5b8a4} /* (30, 1, 21) {real, imag} */,
  {32'hbf024f6d, 32'h3f1a84bd} /* (30, 1, 20) {real, imag} */,
  {32'h3dfb848c, 32'h405320f9} /* (30, 1, 19) {real, imag} */,
  {32'h40915d2f, 32'hbf826d14} /* (30, 1, 18) {real, imag} */,
  {32'hbd1fdad1, 32'h3ea4843d} /* (30, 1, 17) {real, imag} */,
  {32'h3f04ee2a, 32'hbf65538a} /* (30, 1, 16) {real, imag} */,
  {32'h4016b34f, 32'h3f9f0ffb} /* (30, 1, 15) {real, imag} */,
  {32'hc0a2af1c, 32'hbfe25a27} /* (30, 1, 14) {real, imag} */,
  {32'h3f18767d, 32'hbfab01c8} /* (30, 1, 13) {real, imag} */,
  {32'hbefb618f, 32'hbfd6b4cd} /* (30, 1, 12) {real, imag} */,
  {32'hc0812554, 32'h40ad2f43} /* (30, 1, 11) {real, imag} */,
  {32'h3fa39e56, 32'h408111d6} /* (30, 1, 10) {real, imag} */,
  {32'hbfc18ac4, 32'h3f2e0329} /* (30, 1, 9) {real, imag} */,
  {32'hc17bcab0, 32'h412bbe0e} /* (30, 1, 8) {real, imag} */,
  {32'h40d2f533, 32'hc0ab4cf5} /* (30, 1, 7) {real, imag} */,
  {32'h3f136497, 32'h403b6f8e} /* (30, 1, 6) {real, imag} */,
  {32'hc11c1686, 32'h4200ba84} /* (30, 1, 5) {real, imag} */,
  {32'h4184de41, 32'hc0132bcb} /* (30, 1, 4) {real, imag} */,
  {32'h408f793e, 32'h41b34366} /* (30, 1, 3) {real, imag} */,
  {32'hc32b295f, 32'h4383799c} /* (30, 1, 2) {real, imag} */,
  {32'h43750664, 32'hc44999dc} /* (30, 1, 1) {real, imag} */,
  {32'hc2afa8fc, 32'hc41443e2} /* (30, 1, 0) {real, imag} */,
  {32'hc3c36af0, 32'hc3a7593f} /* (30, 0, 31) {real, imag} */,
  {32'h42eeccbe, 32'h4229bd12} /* (30, 0, 30) {real, imag} */,
  {32'h415f0961, 32'h419a76a0} /* (30, 0, 29) {real, imag} */,
  {32'h4155c923, 32'h3fcb0799} /* (30, 0, 28) {real, imag} */,
  {32'h40a975c8, 32'h41d4565e} /* (30, 0, 27) {real, imag} */,
  {32'hc09510c4, 32'h40338645} /* (30, 0, 26) {real, imag} */,
  {32'hc1802800, 32'h403ca201} /* (30, 0, 25) {real, imag} */,
  {32'h414aaaf1, 32'hc010aea1} /* (30, 0, 24) {real, imag} */,
  {32'h3fd1e90f, 32'h4085a126} /* (30, 0, 23) {real, imag} */,
  {32'h40200834, 32'hc00fe783} /* (30, 0, 22) {real, imag} */,
  {32'h404f99ba, 32'hbe829f24} /* (30, 0, 21) {real, imag} */,
  {32'h400e87a5, 32'h3fa5e5d4} /* (30, 0, 20) {real, imag} */,
  {32'hc01b6059, 32'h40158a47} /* (30, 0, 19) {real, imag} */,
  {32'hbf513d6f, 32'hbf1e8120} /* (30, 0, 18) {real, imag} */,
  {32'h3f2b66b0, 32'hbe88768f} /* (30, 0, 17) {real, imag} */,
  {32'hbf22ff31, 32'h3f595a4f} /* (30, 0, 16) {real, imag} */,
  {32'h3f98a979, 32'hbfddf0aa} /* (30, 0, 15) {real, imag} */,
  {32'hbf6fa3d0, 32'h3e38170d} /* (30, 0, 14) {real, imag} */,
  {32'h3ff47b1d, 32'h3f723380} /* (30, 0, 13) {real, imag} */,
  {32'h407182b2, 32'hc0956e94} /* (30, 0, 12) {real, imag} */,
  {32'hbf4a8bc6, 32'h405b4cde} /* (30, 0, 11) {real, imag} */,
  {32'hbfadbb07, 32'h404d6fa9} /* (30, 0, 10) {real, imag} */,
  {32'h3e9bea89, 32'h40538dc6} /* (30, 0, 9) {real, imag} */,
  {32'hc10566f5, 32'h3f0b4d1d} /* (30, 0, 8) {real, imag} */,
  {32'h4048b250, 32'hc01dd484} /* (30, 0, 7) {real, imag} */,
  {32'hbf925047, 32'h40b5e02c} /* (30, 0, 6) {real, imag} */,
  {32'h40a57bae, 32'h41e2251c} /* (30, 0, 5) {real, imag} */,
  {32'hc1fcdbb5, 32'hbfe29442} /* (30, 0, 4) {real, imag} */,
  {32'h3f6de1f0, 32'h418b0cfa} /* (30, 0, 3) {real, imag} */,
  {32'hc2dd8506, 32'h42c375da} /* (30, 0, 2) {real, imag} */,
  {32'h43625fb0, 32'hc3ddd790} /* (30, 0, 1) {real, imag} */,
  {32'hc2d25a25, 32'hc3eb6535} /* (30, 0, 0) {real, imag} */,
  {32'hc305191c, 32'hc312a991} /* (29, 31, 31) {real, imag} */,
  {32'h428de949, 32'h4236a51c} /* (29, 31, 30) {real, imag} */,
  {32'h4193d282, 32'hc10acee1} /* (29, 31, 29) {real, imag} */,
  {32'h3fb9c2f0, 32'hc112524c} /* (29, 31, 28) {real, imag} */,
  {32'h410bd82b, 32'h415ef585} /* (29, 31, 27) {real, imag} */,
  {32'hc0bfab25, 32'h4087bef7} /* (29, 31, 26) {real, imag} */,
  {32'hc05c90f7, 32'h40c03355} /* (29, 31, 25) {real, imag} */,
  {32'h40c1d97f, 32'h3f086677} /* (29, 31, 24) {real, imag} */,
  {32'h40a6e3db, 32'hbf186961} /* (29, 31, 23) {real, imag} */,
  {32'hbfcb5f66, 32'h40aabdd2} /* (29, 31, 22) {real, imag} */,
  {32'h40a92429, 32'h3f813282} /* (29, 31, 21) {real, imag} */,
  {32'h3fa44955, 32'hbfb4bb7b} /* (29, 31, 20) {real, imag} */,
  {32'hc090fd2b, 32'h3fb65adf} /* (29, 31, 19) {real, imag} */,
  {32'h3fac38ab, 32'hc0214903} /* (29, 31, 18) {real, imag} */,
  {32'hbe779aa0, 32'h3fa174b7} /* (29, 31, 17) {real, imag} */,
  {32'h3fc807aa, 32'hbf869e0c} /* (29, 31, 16) {real, imag} */,
  {32'hbf3c2eb6, 32'h3fb3cac4} /* (29, 31, 15) {real, imag} */,
  {32'hc03cb5ad, 32'h3e6c8d9a} /* (29, 31, 14) {real, imag} */,
  {32'hc0054d15, 32'hbeddf50e} /* (29, 31, 13) {real, imag} */,
  {32'hc00139ae, 32'hc004f27e} /* (29, 31, 12) {real, imag} */,
  {32'hbefa3260, 32'h4077ab16} /* (29, 31, 11) {real, imag} */,
  {32'h40029cc3, 32'hc0245fd5} /* (29, 31, 10) {real, imag} */,
  {32'h3fa8c932, 32'h3f75c066} /* (29, 31, 9) {real, imag} */,
  {32'hc0489e6d, 32'h40bc6647} /* (29, 31, 8) {real, imag} */,
  {32'h40eed908, 32'hbff1df49} /* (29, 31, 7) {real, imag} */,
  {32'hbfb12724, 32'h405b4a53} /* (29, 31, 6) {real, imag} */,
  {32'h40eaa911, 32'h41a48fdb} /* (29, 31, 5) {real, imag} */,
  {32'hc17a3ebd, 32'hc17a5bdf} /* (29, 31, 4) {real, imag} */,
  {32'hc09296ea, 32'h418fe05d} /* (29, 31, 3) {real, imag} */,
  {32'h41a54c6d, 32'h41ea1b89} /* (29, 31, 2) {real, imag} */,
  {32'hc156cbdc, 32'hc309411e} /* (29, 31, 1) {real, imag} */,
  {32'hc239a83e, 32'hc2edf486} /* (29, 31, 0) {real, imag} */,
  {32'h3e0edecd, 32'h42797067} /* (29, 30, 31) {real, imag} */,
  {32'hbf461e4e, 32'hc237bc33} /* (29, 30, 30) {real, imag} */,
  {32'hc09c3ece, 32'h40a52078} /* (29, 30, 29) {real, imag} */,
  {32'h410ddbb4, 32'h40ed8c99} /* (29, 30, 28) {real, imag} */,
  {32'hc0978e0e, 32'hc1031486} /* (29, 30, 27) {real, imag} */,
  {32'h3f2677fd, 32'h3faa731c} /* (29, 30, 26) {real, imag} */,
  {32'h4061550d, 32'h3fe4fa8b} /* (29, 30, 25) {real, imag} */,
  {32'hbe725135, 32'h3d92f1a9} /* (29, 30, 24) {real, imag} */,
  {32'hc0261f69, 32'hbf82e819} /* (29, 30, 23) {real, imag} */,
  {32'h401a2f6b, 32'h401010a1} /* (29, 30, 22) {real, imag} */,
  {32'hbfdeb1e8, 32'hbf332e49} /* (29, 30, 21) {real, imag} */,
  {32'h401b2741, 32'h3ff88e6f} /* (29, 30, 20) {real, imag} */,
  {32'hbe1a92ea, 32'hbf26b3a5} /* (29, 30, 19) {real, imag} */,
  {32'hbdfbab29, 32'h3f637d52} /* (29, 30, 18) {real, imag} */,
  {32'hbd9e4d98, 32'h3fc6489a} /* (29, 30, 17) {real, imag} */,
  {32'h3d0b7e42, 32'hbfb3f94a} /* (29, 30, 16) {real, imag} */,
  {32'hbfa64b0d, 32'h3e9da80f} /* (29, 30, 15) {real, imag} */,
  {32'h3eeeddca, 32'h3f0555ec} /* (29, 30, 14) {real, imag} */,
  {32'h40139edf, 32'hbf484c37} /* (29, 30, 13) {real, imag} */,
  {32'hbf70da12, 32'hc0154323} /* (29, 30, 12) {real, imag} */,
  {32'h402646cc, 32'h4023e261} /* (29, 30, 11) {real, imag} */,
  {32'hc0ae287e, 32'h3f3287fb} /* (29, 30, 10) {real, imag} */,
  {32'hc00d2dab, 32'hbfff3ef1} /* (29, 30, 9) {real, imag} */,
  {32'h3ff86345, 32'hc0ba86e4} /* (29, 30, 8) {real, imag} */,
  {32'h3eb6a0e3, 32'hbe167ddd} /* (29, 30, 7) {real, imag} */,
  {32'h3fe8e697, 32'hbff13430} /* (29, 30, 6) {real, imag} */,
  {32'h40b3d60d, 32'hc11e1b0e} /* (29, 30, 5) {real, imag} */,
  {32'hc13f49f0, 32'h409d3dd2} /* (29, 30, 4) {real, imag} */,
  {32'h3f2497ba, 32'h40ffd906} /* (29, 30, 3) {real, imag} */,
  {32'hc122bd67, 32'hc285d676} /* (29, 30, 2) {real, imag} */,
  {32'h42350981, 32'h42fa7b46} /* (29, 30, 1) {real, imag} */,
  {32'h41eb9fff, 32'h422de765} /* (29, 30, 0) {real, imag} */,
  {32'hc1672ddb, 32'hc0348f70} /* (29, 29, 31) {real, imag} */,
  {32'h4152d32d, 32'hc14c7491} /* (29, 29, 30) {real, imag} */,
  {32'hbffe0a78, 32'hc1013dbd} /* (29, 29, 29) {real, imag} */,
  {32'hc08dd30f, 32'h415fc88b} /* (29, 29, 28) {real, imag} */,
  {32'hc02a8370, 32'hc0c94701} /* (29, 29, 27) {real, imag} */,
  {32'h4097c6df, 32'hc01c03b8} /* (29, 29, 26) {real, imag} */,
  {32'hc07f4c49, 32'h4020f3c7} /* (29, 29, 25) {real, imag} */,
  {32'h3ef1d2cc, 32'hc02680b9} /* (29, 29, 24) {real, imag} */,
  {32'hc086b745, 32'h3e8ef1ab} /* (29, 29, 23) {real, imag} */,
  {32'h400b7aaf, 32'hbfd4571a} /* (29, 29, 22) {real, imag} */,
  {32'h3e49adc0, 32'hbffb1ec5} /* (29, 29, 21) {real, imag} */,
  {32'h401b7461, 32'hc0219d5d} /* (29, 29, 20) {real, imag} */,
  {32'h3f66ab3b, 32'hbfccf8bc} /* (29, 29, 19) {real, imag} */,
  {32'h3ef6bd0a, 32'h3fb405c4} /* (29, 29, 18) {real, imag} */,
  {32'hbfd4efd5, 32'h3f40fcbe} /* (29, 29, 17) {real, imag} */,
  {32'h3ff78287, 32'h3fb2d139} /* (29, 29, 16) {real, imag} */,
  {32'h40067646, 32'hbf8dbb0a} /* (29, 29, 15) {real, imag} */,
  {32'h4017f213, 32'hbf846594} /* (29, 29, 14) {real, imag} */,
  {32'hc0997ba9, 32'hbf4cafc6} /* (29, 29, 13) {real, imag} */,
  {32'h3f978cfa, 32'hbf26c8b3} /* (29, 29, 12) {real, imag} */,
  {32'h3e83226d, 32'h3e5b57ca} /* (29, 29, 11) {real, imag} */,
  {32'hbfc6dcc2, 32'h401b7a6c} /* (29, 29, 10) {real, imag} */,
  {32'hc0874862, 32'hbf309b80} /* (29, 29, 9) {real, imag} */,
  {32'h4124b160, 32'hbfe6d2ea} /* (29, 29, 8) {real, imag} */,
  {32'hc018a876, 32'h40dbf8b8} /* (29, 29, 7) {real, imag} */,
  {32'h40bd73a7, 32'hbcb8ac42} /* (29, 29, 6) {real, imag} */,
  {32'h405402ad, 32'h400d712c} /* (29, 29, 5) {real, imag} */,
  {32'hc0900e9d, 32'hbeaceec9} /* (29, 29, 4) {real, imag} */,
  {32'hbeaf6fb8, 32'h3ed57494} /* (29, 29, 3) {real, imag} */,
  {32'h3f9367d1, 32'hc12c782d} /* (29, 29, 2) {real, imag} */,
  {32'hc08c98ce, 32'h41b50186} /* (29, 29, 1) {real, imag} */,
  {32'hc05308e2, 32'h4168914e} /* (29, 29, 0) {real, imag} */,
  {32'hc16327ba, 32'hc18e6c47} /* (29, 28, 31) {real, imag} */,
  {32'h419e7eed, 32'h4108a5d4} /* (29, 28, 30) {real, imag} */,
  {32'h40cbbe5d, 32'h405685f9} /* (29, 28, 29) {real, imag} */,
  {32'hc11c79da, 32'hc0b4e4e0} /* (29, 28, 28) {real, imag} */,
  {32'h40cfad1b, 32'h3fc22649} /* (29, 28, 27) {real, imag} */,
  {32'hbdf96e97, 32'hc02e5f4d} /* (29, 28, 26) {real, imag} */,
  {32'h405a0273, 32'h3d3c5b72} /* (29, 28, 25) {real, imag} */,
  {32'h403b200c, 32'h405720fb} /* (29, 28, 24) {real, imag} */,
  {32'h4038f582, 32'h3f09a6ff} /* (29, 28, 23) {real, imag} */,
  {32'hc047901e, 32'hbf639236} /* (29, 28, 22) {real, imag} */,
  {32'h400c31b2, 32'hbfb0f8f9} /* (29, 28, 21) {real, imag} */,
  {32'hbd17ee89, 32'h3f8463df} /* (29, 28, 20) {real, imag} */,
  {32'h3f1e239e, 32'h3ee2b1df} /* (29, 28, 19) {real, imag} */,
  {32'h40050d63, 32'h3faa71fb} /* (29, 28, 18) {real, imag} */,
  {32'h3f1b672b, 32'h401ba190} /* (29, 28, 17) {real, imag} */,
  {32'h3e1d6b4e, 32'hbd9cf8ce} /* (29, 28, 16) {real, imag} */,
  {32'h3f41a6c4, 32'hbf669b9f} /* (29, 28, 15) {real, imag} */,
  {32'h3f0e5ad8, 32'h3f4d64ed} /* (29, 28, 14) {real, imag} */,
  {32'h3e5eeefc, 32'hbf3b27fa} /* (29, 28, 13) {real, imag} */,
  {32'h3f87c16d, 32'hbfb85295} /* (29, 28, 12) {real, imag} */,
  {32'hbf717df2, 32'h4003cf8a} /* (29, 28, 11) {real, imag} */,
  {32'hbfc9cf76, 32'hc00c2427} /* (29, 28, 10) {real, imag} */,
  {32'hbdf4fc27, 32'h3fc6245d} /* (29, 28, 9) {real, imag} */,
  {32'h400b8e5d, 32'h3f11cf15} /* (29, 28, 8) {real, imag} */,
  {32'h402e92fa, 32'h3fd45ca4} /* (29, 28, 7) {real, imag} */,
  {32'hbfaeadc4, 32'h4088e21a} /* (29, 28, 6) {real, imag} */,
  {32'h3e98ca41, 32'h40e00290} /* (29, 28, 5) {real, imag} */,
  {32'hbd57e5e4, 32'hc0aa5fc9} /* (29, 28, 4) {real, imag} */,
  {32'hc098c676, 32'hbfd71129} /* (29, 28, 3) {real, imag} */,
  {32'h415e52e1, 32'h41308ece} /* (29, 28, 2) {real, imag} */,
  {32'hc18c773f, 32'hc125908f} /* (29, 28, 1) {real, imag} */,
  {32'hc08fda18, 32'hc1bf6cb2} /* (29, 28, 0) {real, imag} */,
  {32'h41a2e425, 32'h410092fa} /* (29, 27, 31) {real, imag} */,
  {32'hbfb6d6cb, 32'hc0ea0352} /* (29, 27, 30) {real, imag} */,
  {32'hc0818064, 32'h3f64a0f2} /* (29, 27, 29) {real, imag} */,
  {32'hbf849c7c, 32'h3fa770f0} /* (29, 27, 28) {real, imag} */,
  {32'hc0d57fcd, 32'h4086c11d} /* (29, 27, 27) {real, imag} */,
  {32'h3fc0ca1f, 32'hc02f167c} /* (29, 27, 26) {real, imag} */,
  {32'h408b521f, 32'hbeefd78e} /* (29, 27, 25) {real, imag} */,
  {32'hbf9fa26f, 32'hc00d12f9} /* (29, 27, 24) {real, imag} */,
  {32'h4027f69c, 32'hbff97103} /* (29, 27, 23) {real, imag} */,
  {32'hc012e072, 32'hc01b205e} /* (29, 27, 22) {real, imag} */,
  {32'h3ebda071, 32'h4018e76f} /* (29, 27, 21) {real, imag} */,
  {32'h3fa898e7, 32'hc01745fc} /* (29, 27, 20) {real, imag} */,
  {32'h3e8bdf78, 32'h3e093580} /* (29, 27, 19) {real, imag} */,
  {32'hc012ba9f, 32'h3e3a3257} /* (29, 27, 18) {real, imag} */,
  {32'hbf078f01, 32'hbeceb292} /* (29, 27, 17) {real, imag} */,
  {32'hbf4077c7, 32'hc01105e6} /* (29, 27, 16) {real, imag} */,
  {32'hbd4551f2, 32'hbf855491} /* (29, 27, 15) {real, imag} */,
  {32'hbfbdf442, 32'hbf995e5f} /* (29, 27, 14) {real, imag} */,
  {32'h40413538, 32'h3e9df0c6} /* (29, 27, 13) {real, imag} */,
  {32'h3fd6e36a, 32'h3f3d41fd} /* (29, 27, 12) {real, imag} */,
  {32'h3fcc7169, 32'hbfd27998} /* (29, 27, 11) {real, imag} */,
  {32'hbfc9a999, 32'h3e614d9c} /* (29, 27, 10) {real, imag} */,
  {32'h3fc33f49, 32'h3f81d43a} /* (29, 27, 9) {real, imag} */,
  {32'h406540c7, 32'h4029490a} /* (29, 27, 8) {real, imag} */,
  {32'hc0af9a51, 32'h3ff4604d} /* (29, 27, 7) {real, imag} */,
  {32'hc04ee3ed, 32'h3fc699b2} /* (29, 27, 6) {real, imag} */,
  {32'hbfc373a5, 32'hc0dec2c2} /* (29, 27, 5) {real, imag} */,
  {32'h3f2f2677, 32'h400f3bb8} /* (29, 27, 4) {real, imag} */,
  {32'hbf224813, 32'hc0ac12f7} /* (29, 27, 3) {real, imag} */,
  {32'hc05ba367, 32'hc1290779} /* (29, 27, 2) {real, imag} */,
  {32'h40cf63af, 32'h41b550d2} /* (29, 27, 1) {real, imag} */,
  {32'h40e0630f, 32'h413cbcad} /* (29, 27, 0) {real, imag} */,
  {32'hbe3b6f49, 32'h40b73fb9} /* (29, 26, 31) {real, imag} */,
  {32'h3feb47b3, 32'h40d209da} /* (29, 26, 30) {real, imag} */,
  {32'h40497701, 32'h3f894c1d} /* (29, 26, 29) {real, imag} */,
  {32'hbf99900a, 32'hbef7e6b0} /* (29, 26, 28) {real, imag} */,
  {32'hc000b00f, 32'h3e4e020f} /* (29, 26, 27) {real, imag} */,
  {32'hc024436a, 32'hbf7c6631} /* (29, 26, 26) {real, imag} */,
  {32'hc0f4274b, 32'hc08b2ab0} /* (29, 26, 25) {real, imag} */,
  {32'h3f9de225, 32'h400cd59b} /* (29, 26, 24) {real, imag} */,
  {32'hbf63524f, 32'h3e45e47a} /* (29, 26, 23) {real, imag} */,
  {32'hbf417089, 32'h3fb04aae} /* (29, 26, 22) {real, imag} */,
  {32'hbf894c35, 32'hbf80bf34} /* (29, 26, 21) {real, imag} */,
  {32'hc056c37d, 32'hbf8de583} /* (29, 26, 20) {real, imag} */,
  {32'hbf9b96e4, 32'hbef45485} /* (29, 26, 19) {real, imag} */,
  {32'h3f1bf115, 32'h3e365f7d} /* (29, 26, 18) {real, imag} */,
  {32'hbf368527, 32'h3fcd4995} /* (29, 26, 17) {real, imag} */,
  {32'hbfb1ced6, 32'h3f502797} /* (29, 26, 16) {real, imag} */,
  {32'h3f3a6790, 32'h3f90e7a5} /* (29, 26, 15) {real, imag} */,
  {32'hc02b2552, 32'hbf522f3f} /* (29, 26, 14) {real, imag} */,
  {32'h400cf67c, 32'hbf648ea2} /* (29, 26, 13) {real, imag} */,
  {32'h4024d7d3, 32'h3f9a1cd0} /* (29, 26, 12) {real, imag} */,
  {32'h3f899e2c, 32'hbf8ebbc8} /* (29, 26, 11) {real, imag} */,
  {32'h3f0abd42, 32'h405eeb20} /* (29, 26, 10) {real, imag} */,
  {32'hbda36846, 32'hc0d11e32} /* (29, 26, 9) {real, imag} */,
  {32'h3e29e194, 32'h3f1586cd} /* (29, 26, 8) {real, imag} */,
  {32'hc0348af6, 32'h3fc0acd3} /* (29, 26, 7) {real, imag} */,
  {32'h40243e8d, 32'hc0863a4d} /* (29, 26, 6) {real, imag} */,
  {32'h3f99d84c, 32'h4095512a} /* (29, 26, 5) {real, imag} */,
  {32'hbe49cc70, 32'h3f8d9687} /* (29, 26, 4) {real, imag} */,
  {32'hbf499fb3, 32'h3ee6bc7d} /* (29, 26, 3) {real, imag} */,
  {32'h3ff5cfb9, 32'h404b9900} /* (29, 26, 2) {real, imag} */,
  {32'hc0544b3e, 32'h403439f2} /* (29, 26, 1) {real, imag} */,
  {32'h3fedd97d, 32'hc06ec828} /* (29, 26, 0) {real, imag} */,
  {32'hbe8e2bbc, 32'hbfa5f9aa} /* (29, 25, 31) {real, imag} */,
  {32'h4022ae4b, 32'h3fe65434} /* (29, 25, 30) {real, imag} */,
  {32'h404dea96, 32'hbfbd2870} /* (29, 25, 29) {real, imag} */,
  {32'hc07e78ad, 32'hc05afbcf} /* (29, 25, 28) {real, imag} */,
  {32'h405e7499, 32'hc02c37ef} /* (29, 25, 27) {real, imag} */,
  {32'h3f45aaec, 32'hbf8842ac} /* (29, 25, 26) {real, imag} */,
  {32'hbfc72b43, 32'h3f867dbf} /* (29, 25, 25) {real, imag} */,
  {32'h3f1f4136, 32'h3f879f5b} /* (29, 25, 24) {real, imag} */,
  {32'hc02b0197, 32'h3caec191} /* (29, 25, 23) {real, imag} */,
  {32'h40980f9c, 32'hbf89e9b3} /* (29, 25, 22) {real, imag} */,
  {32'hbf12d479, 32'hbf8f16c2} /* (29, 25, 21) {real, imag} */,
  {32'h3f8d7aa6, 32'h3ed1681e} /* (29, 25, 20) {real, imag} */,
  {32'h40079594, 32'h3f173295} /* (29, 25, 19) {real, imag} */,
  {32'hc0080ea3, 32'hbefe3aca} /* (29, 25, 18) {real, imag} */,
  {32'h4001665c, 32'hbe00aacf} /* (29, 25, 17) {real, imag} */,
  {32'h3e6fb714, 32'hbf16de8e} /* (29, 25, 16) {real, imag} */,
  {32'h3fe77170, 32'h3f7008dc} /* (29, 25, 15) {real, imag} */,
  {32'h3f207332, 32'hc03f1754} /* (29, 25, 14) {real, imag} */,
  {32'h3f9f2459, 32'hc078ad53} /* (29, 25, 13) {real, imag} */,
  {32'hc026796d, 32'h3fcde374} /* (29, 25, 12) {real, imag} */,
  {32'hc01714f8, 32'hbe723c75} /* (29, 25, 11) {real, imag} */,
  {32'hbff4a5ff, 32'hbbc9904c} /* (29, 25, 10) {real, imag} */,
  {32'h3e81c838, 32'h3fefcd7e} /* (29, 25, 9) {real, imag} */,
  {32'hbfa6a23e, 32'hbf81f8de} /* (29, 25, 8) {real, imag} */,
  {32'h3fd1cdc7, 32'h3f9a509d} /* (29, 25, 7) {real, imag} */,
  {32'h3f07a552, 32'hc06d30f5} /* (29, 25, 6) {real, imag} */,
  {32'h3f17a4f5, 32'h3f93c984} /* (29, 25, 5) {real, imag} */,
  {32'h401bb393, 32'hc04f664a} /* (29, 25, 4) {real, imag} */,
  {32'h3f840823, 32'hc01138c7} /* (29, 25, 3) {real, imag} */,
  {32'h3d8f0b8d, 32'h3de1614d} /* (29, 25, 2) {real, imag} */,
  {32'h3fd75b98, 32'h3fda3262} /* (29, 25, 1) {real, imag} */,
  {32'h3f2151c2, 32'hc0905de5} /* (29, 25, 0) {real, imag} */,
  {32'h408656ba, 32'h3eaaa2b5} /* (29, 24, 31) {real, imag} */,
  {32'hbf4a5e6e, 32'hc05bd5ac} /* (29, 24, 30) {real, imag} */,
  {32'hc08efb8f, 32'h403d6df5} /* (29, 24, 29) {real, imag} */,
  {32'h3f9b0c69, 32'hc08436d0} /* (29, 24, 28) {real, imag} */,
  {32'hbf2ebb89, 32'h402e15c6} /* (29, 24, 27) {real, imag} */,
  {32'h3d7353f4, 32'hbfe13940} /* (29, 24, 26) {real, imag} */,
  {32'hc054d775, 32'h3ee8c705} /* (29, 24, 25) {real, imag} */,
  {32'hc09623d0, 32'h3f775233} /* (29, 24, 24) {real, imag} */,
  {32'h3f7b1c18, 32'h402a4d01} /* (29, 24, 23) {real, imag} */,
  {32'hbeaf0e6a, 32'hc09ec0de} /* (29, 24, 22) {real, imag} */,
  {32'hc09be87a, 32'h406c9191} /* (29, 24, 21) {real, imag} */,
  {32'h3f916923, 32'h3fafee2d} /* (29, 24, 20) {real, imag} */,
  {32'hbfe143a3, 32'hbe332f46} /* (29, 24, 19) {real, imag} */,
  {32'h3e496e5a, 32'h3f35f8dd} /* (29, 24, 18) {real, imag} */,
  {32'h3e0a31e8, 32'h3f345b05} /* (29, 24, 17) {real, imag} */,
  {32'hbf9199b0, 32'hbdf53c33} /* (29, 24, 16) {real, imag} */,
  {32'h3e871995, 32'h3fdf8de8} /* (29, 24, 15) {real, imag} */,
  {32'h3f4b61be, 32'h3f5892fb} /* (29, 24, 14) {real, imag} */,
  {32'h3fefbdfa, 32'hbf3d6fc5} /* (29, 24, 13) {real, imag} */,
  {32'hbec61305, 32'hbecb3cf0} /* (29, 24, 12) {real, imag} */,
  {32'hc01854f0, 32'h3fc5c7c6} /* (29, 24, 11) {real, imag} */,
  {32'hbe979af9, 32'hbfe478e7} /* (29, 24, 10) {real, imag} */,
  {32'h3fb102fe, 32'hbcf84efa} /* (29, 24, 9) {real, imag} */,
  {32'h3fa92dbc, 32'h3f25fbaa} /* (29, 24, 8) {real, imag} */,
  {32'h408f2518, 32'h40020a47} /* (29, 24, 7) {real, imag} */,
  {32'h4072f5cd, 32'h3f832d9a} /* (29, 24, 6) {real, imag} */,
  {32'hbea48db3, 32'h3f1f061c} /* (29, 24, 5) {real, imag} */,
  {32'hbf5a648c, 32'hbf95de39} /* (29, 24, 4) {real, imag} */,
  {32'hbfcf7554, 32'h3fc25c17} /* (29, 24, 3) {real, imag} */,
  {32'hbda6c9d5, 32'hc0a9084a} /* (29, 24, 2) {real, imag} */,
  {32'h407042a5, 32'h40bcee6f} /* (29, 24, 1) {real, imag} */,
  {32'h402d1bdd, 32'h4087f2e5} /* (29, 24, 0) {real, imag} */,
  {32'hbf39ddb7, 32'hc0da730a} /* (29, 23, 31) {real, imag} */,
  {32'hc0043b2d, 32'h3f153de8} /* (29, 23, 30) {real, imag} */,
  {32'h3f5575b1, 32'h3fdcc5c0} /* (29, 23, 29) {real, imag} */,
  {32'hbf379ba9, 32'hc0032a00} /* (29, 23, 28) {real, imag} */,
  {32'hc0863403, 32'h3fb4941f} /* (29, 23, 27) {real, imag} */,
  {32'hbff98d5a, 32'h3fb336fd} /* (29, 23, 26) {real, imag} */,
  {32'h3fc1f29c, 32'h3f19495f} /* (29, 23, 25) {real, imag} */,
  {32'h3ee45f1b, 32'hbfaa9888} /* (29, 23, 24) {real, imag} */,
  {32'h3ed8e5ad, 32'h3ffdec9b} /* (29, 23, 23) {real, imag} */,
  {32'h3fe736ac, 32'hc029a599} /* (29, 23, 22) {real, imag} */,
  {32'h3fbd1c22, 32'hbefe1ad8} /* (29, 23, 21) {real, imag} */,
  {32'h3f3a9bc0, 32'h3ee4a463} /* (29, 23, 20) {real, imag} */,
  {32'hbfcbf6a4, 32'h3f8a4f78} /* (29, 23, 19) {real, imag} */,
  {32'hbfda4ee0, 32'h3ef2e015} /* (29, 23, 18) {real, imag} */,
  {32'hbe928ee1, 32'hbeb68f9f} /* (29, 23, 17) {real, imag} */,
  {32'hbef68c41, 32'hbeeaa077} /* (29, 23, 16) {real, imag} */,
  {32'hbf2f84fb, 32'h3d726d33} /* (29, 23, 15) {real, imag} */,
  {32'h3ff94224, 32'hbf46c065} /* (29, 23, 14) {real, imag} */,
  {32'hbf9a3517, 32'h408433a9} /* (29, 23, 13) {real, imag} */,
  {32'h3f526379, 32'h40221241} /* (29, 23, 12) {real, imag} */,
  {32'hbfcc039c, 32'hc000eef6} /* (29, 23, 11) {real, imag} */,
  {32'h3fbc68d5, 32'hbff47aa6} /* (29, 23, 10) {real, imag} */,
  {32'h3f87ea77, 32'h3fa5c48a} /* (29, 23, 9) {real, imag} */,
  {32'hbf1d90e8, 32'hbf3dbfb0} /* (29, 23, 8) {real, imag} */,
  {32'hc00df3f1, 32'h3f0c6194} /* (29, 23, 7) {real, imag} */,
  {32'hbf91c9d5, 32'h404ea6b2} /* (29, 23, 6) {real, imag} */,
  {32'h404762b9, 32'h403e6069} /* (29, 23, 5) {real, imag} */,
  {32'h3fd97e89, 32'h40b617ab} /* (29, 23, 4) {real, imag} */,
  {32'hc09e1285, 32'hbfc16734} /* (29, 23, 3) {real, imag} */,
  {32'h4040c6d4, 32'hbf4f3770} /* (29, 23, 2) {real, imag} */,
  {32'hc00d905c, 32'h4087c143} /* (29, 23, 1) {real, imag} */,
  {32'h3fce5bf5, 32'h3f9e872c} /* (29, 23, 0) {real, imag} */,
  {32'hc0763e19, 32'hbf1fc4f5} /* (29, 22, 31) {real, imag} */,
  {32'h403af073, 32'hc0137a86} /* (29, 22, 30) {real, imag} */,
  {32'h40470e3c, 32'h3ffb6932} /* (29, 22, 29) {real, imag} */,
  {32'h3d219c9a, 32'hbdf66766} /* (29, 22, 28) {real, imag} */,
  {32'h3f245149, 32'h404ff351} /* (29, 22, 27) {real, imag} */,
  {32'h3fb749c1, 32'h4094dd39} /* (29, 22, 26) {real, imag} */,
  {32'h3f25c5c0, 32'h3fe5a3ae} /* (29, 22, 25) {real, imag} */,
  {32'hc02481a5, 32'h3deca734} /* (29, 22, 24) {real, imag} */,
  {32'h3f807290, 32'h3f2e9e8e} /* (29, 22, 23) {real, imag} */,
  {32'hbfb4aed6, 32'h401acd7b} /* (29, 22, 22) {real, imag} */,
  {32'hbd18f747, 32'h3f5270f4} /* (29, 22, 21) {real, imag} */,
  {32'hc0108dca, 32'hbdf0e7a6} /* (29, 22, 20) {real, imag} */,
  {32'hbf2cb94a, 32'hc04dd813} /* (29, 22, 19) {real, imag} */,
  {32'hbf740269, 32'h3ee35052} /* (29, 22, 18) {real, imag} */,
  {32'h3ff8d4bd, 32'hbf896060} /* (29, 22, 17) {real, imag} */,
  {32'h3f129543, 32'h3f64da3b} /* (29, 22, 16) {real, imag} */,
  {32'hbf8a868a, 32'h3f437d3f} /* (29, 22, 15) {real, imag} */,
  {32'h3ecce083, 32'hbebd89ec} /* (29, 22, 14) {real, imag} */,
  {32'hbfc5b79a, 32'h3f9f00e1} /* (29, 22, 13) {real, imag} */,
  {32'h3e8b8882, 32'hc0818ec6} /* (29, 22, 12) {real, imag} */,
  {32'hc0556e64, 32'hc0768a08} /* (29, 22, 11) {real, imag} */,
  {32'h4007c179, 32'h4026aedb} /* (29, 22, 10) {real, imag} */,
  {32'hbf945c1f, 32'h40695d60} /* (29, 22, 9) {real, imag} */,
  {32'h40afa642, 32'hbee22a6b} /* (29, 22, 8) {real, imag} */,
  {32'h3eac2612, 32'h3d96c174} /* (29, 22, 7) {real, imag} */,
  {32'hbf3a619f, 32'h3e8bc337} /* (29, 22, 6) {real, imag} */,
  {32'h3f8a7ec3, 32'hbf852291} /* (29, 22, 5) {real, imag} */,
  {32'hbf39d105, 32'hbf5c28cd} /* (29, 22, 4) {real, imag} */,
  {32'hbf9759b0, 32'hbf33d793} /* (29, 22, 3) {real, imag} */,
  {32'h4041e4bf, 32'hc0381928} /* (29, 22, 2) {real, imag} */,
  {32'hbe0b72db, 32'hbf0df828} /* (29, 22, 1) {real, imag} */,
  {32'hc01d8daa, 32'h40dce454} /* (29, 22, 0) {real, imag} */,
  {32'h4077a877, 32'hbfc7e879} /* (29, 21, 31) {real, imag} */,
  {32'hc0829c46, 32'hbf5af039} /* (29, 21, 30) {real, imag} */,
  {32'h3f907739, 32'h3f5a2d09} /* (29, 21, 29) {real, imag} */,
  {32'h3f8231e7, 32'h4005576d} /* (29, 21, 28) {real, imag} */,
  {32'hbe43a040, 32'hbf960ea0} /* (29, 21, 27) {real, imag} */,
  {32'hbf64711c, 32'h402ed046} /* (29, 21, 26) {real, imag} */,
  {32'h40519300, 32'hbfb6ecf2} /* (29, 21, 25) {real, imag} */,
  {32'hbe447e93, 32'h3f9000ba} /* (29, 21, 24) {real, imag} */,
  {32'hbf5420a8, 32'h3f8a26e1} /* (29, 21, 23) {real, imag} */,
  {32'hc02b6683, 32'hc017f3aa} /* (29, 21, 22) {real, imag} */,
  {32'hc03e036c, 32'h3ea95202} /* (29, 21, 21) {real, imag} */,
  {32'hbf9a147e, 32'hbe006371} /* (29, 21, 20) {real, imag} */,
  {32'h3fe7faa7, 32'h4003b30d} /* (29, 21, 19) {real, imag} */,
  {32'h3eab5090, 32'h400307e0} /* (29, 21, 18) {real, imag} */,
  {32'hbf7a69dc, 32'h3f420dba} /* (29, 21, 17) {real, imag} */,
  {32'hbdd9e18c, 32'h3e0e9955} /* (29, 21, 16) {real, imag} */,
  {32'hbda4ca61, 32'h3e07e2a6} /* (29, 21, 15) {real, imag} */,
  {32'h4033c2fe, 32'hc0421c84} /* (29, 21, 14) {real, imag} */,
  {32'hbd91b779, 32'hbf940a93} /* (29, 21, 13) {real, imag} */,
  {32'h3f0f5f87, 32'hbf0eebf7} /* (29, 21, 12) {real, imag} */,
  {32'h408cbb0c, 32'hbf936635} /* (29, 21, 11) {real, imag} */,
  {32'hbec7e146, 32'h4029aa4f} /* (29, 21, 10) {real, imag} */,
  {32'hbe9edb48, 32'h3ff62f2b} /* (29, 21, 9) {real, imag} */,
  {32'hbf17e641, 32'h40480bab} /* (29, 21, 8) {real, imag} */,
  {32'hc08289e0, 32'hbf37cdb0} /* (29, 21, 7) {real, imag} */,
  {32'hc00bbac0, 32'h3f58fdda} /* (29, 21, 6) {real, imag} */,
  {32'hbf12a33a, 32'hbe66d25b} /* (29, 21, 5) {real, imag} */,
  {32'hbfc137d5, 32'h3f0a4870} /* (29, 21, 4) {real, imag} */,
  {32'hbfeb2d86, 32'hc04e5477} /* (29, 21, 3) {real, imag} */,
  {32'hbffc5481, 32'hbfee7920} /* (29, 21, 2) {real, imag} */,
  {32'h4096aabb, 32'h3ece73a9} /* (29, 21, 1) {real, imag} */,
  {32'h3faec751, 32'h3f110f10} /* (29, 21, 0) {real, imag} */,
  {32'h3ee9496f, 32'h400bf4ed} /* (29, 20, 31) {real, imag} */,
  {32'h3f949b8d, 32'h3de5c5d7} /* (29, 20, 30) {real, imag} */,
  {32'h3dc080d8, 32'h3fef6603} /* (29, 20, 29) {real, imag} */,
  {32'h408a27cb, 32'hbe0d931a} /* (29, 20, 28) {real, imag} */,
  {32'hc043de2d, 32'hbfe83c4d} /* (29, 20, 27) {real, imag} */,
  {32'h3d944ea3, 32'hbd32f524} /* (29, 20, 26) {real, imag} */,
  {32'h3f778bfe, 32'h40178742} /* (29, 20, 25) {real, imag} */,
  {32'hbfbc94ee, 32'h3fb1069e} /* (29, 20, 24) {real, imag} */,
  {32'h3e2e8886, 32'hbfd3bf81} /* (29, 20, 23) {real, imag} */,
  {32'h3fb9e2ac, 32'h3f74d70d} /* (29, 20, 22) {real, imag} */,
  {32'hbf244c9e, 32'hbfb00dcf} /* (29, 20, 21) {real, imag} */,
  {32'h3e7e2b02, 32'hc09001c2} /* (29, 20, 20) {real, imag} */,
  {32'h3e63cb5f, 32'hbfac2cbf} /* (29, 20, 19) {real, imag} */,
  {32'h3f80c4ad, 32'hbae2bab3} /* (29, 20, 18) {real, imag} */,
  {32'hbf827b91, 32'h3e3e616e} /* (29, 20, 17) {real, imag} */,
  {32'h3f751ed5, 32'h3fbf36ed} /* (29, 20, 16) {real, imag} */,
  {32'h3fecb634, 32'hc03d43e5} /* (29, 20, 15) {real, imag} */,
  {32'h3e7babab, 32'h3ecfd3ec} /* (29, 20, 14) {real, imag} */,
  {32'hbf06c8bb, 32'h4080263b} /* (29, 20, 13) {real, imag} */,
  {32'h3fac99f8, 32'h3f4ecb9d} /* (29, 20, 12) {real, imag} */,
  {32'h3f5734dd, 32'hbfdf2ac9} /* (29, 20, 11) {real, imag} */,
  {32'hbf23c813, 32'hbf0e59ca} /* (29, 20, 10) {real, imag} */,
  {32'h3f29e8d7, 32'hbfb43cbe} /* (29, 20, 9) {real, imag} */,
  {32'hc011dcbd, 32'h3fa999db} /* (29, 20, 8) {real, imag} */,
  {32'h3e42de42, 32'h3f22ba8a} /* (29, 20, 7) {real, imag} */,
  {32'h3c8077d1, 32'hc039f8b7} /* (29, 20, 6) {real, imag} */,
  {32'hbfcddf7c, 32'h40295be0} /* (29, 20, 5) {real, imag} */,
  {32'hbfa65484, 32'hbf6b65cc} /* (29, 20, 4) {real, imag} */,
  {32'hbfe2ef4f, 32'h3f8351af} /* (29, 20, 3) {real, imag} */,
  {32'h3ff9b196, 32'h3fa824c2} /* (29, 20, 2) {real, imag} */,
  {32'hbc63d6f1, 32'hbf8ae325} /* (29, 20, 1) {real, imag} */,
  {32'h3e67fde9, 32'hbec4bc0b} /* (29, 20, 0) {real, imag} */,
  {32'hbf1bb909, 32'h3f99834d} /* (29, 19, 31) {real, imag} */,
  {32'h402fbbcf, 32'h3f9e735c} /* (29, 19, 30) {real, imag} */,
  {32'hbe77af20, 32'h3da1dd58} /* (29, 19, 29) {real, imag} */,
  {32'h3f6935a5, 32'hc0061f4c} /* (29, 19, 28) {real, imag} */,
  {32'h3f8f3b1f, 32'h40074401} /* (29, 19, 27) {real, imag} */,
  {32'hbf9896b1, 32'hc01929f1} /* (29, 19, 26) {real, imag} */,
  {32'h3f554613, 32'hbf8d4464} /* (29, 19, 25) {real, imag} */,
  {32'hbf5b99bd, 32'h3f30192f} /* (29, 19, 24) {real, imag} */,
  {32'h3ecba86f, 32'h3e20fcf6} /* (29, 19, 23) {real, imag} */,
  {32'h4000b2f3, 32'hbf875e64} /* (29, 19, 22) {real, imag} */,
  {32'hc028fa43, 32'h40403bad} /* (29, 19, 21) {real, imag} */,
  {32'hc01866ed, 32'h3f287d6c} /* (29, 19, 20) {real, imag} */,
  {32'h3f480b55, 32'hbf5dd4cf} /* (29, 19, 19) {real, imag} */,
  {32'h3f620b19, 32'hbedb4a93} /* (29, 19, 18) {real, imag} */,
  {32'hbee1f1ff, 32'hbfe4848b} /* (29, 19, 17) {real, imag} */,
  {32'h3f6ecf5a, 32'hbfaf8b91} /* (29, 19, 16) {real, imag} */,
  {32'h3f605dae, 32'h3f959e22} /* (29, 19, 15) {real, imag} */,
  {32'hbf1ac461, 32'h3e883e90} /* (29, 19, 14) {real, imag} */,
  {32'hbfee7941, 32'hc0237bc9} /* (29, 19, 13) {real, imag} */,
  {32'hbfc48bf5, 32'h3f9b2433} /* (29, 19, 12) {real, imag} */,
  {32'h3fd72bd4, 32'hbf1351d3} /* (29, 19, 11) {real, imag} */,
  {32'h3f5a7621, 32'h3e0039f8} /* (29, 19, 10) {real, imag} */,
  {32'hbf30919a, 32'hbfae6bea} /* (29, 19, 9) {real, imag} */,
  {32'h3fc8984f, 32'h3f115164} /* (29, 19, 8) {real, imag} */,
  {32'h3fc3b785, 32'hbf3f196e} /* (29, 19, 7) {real, imag} */,
  {32'h402deeca, 32'h3f51bd96} /* (29, 19, 6) {real, imag} */,
  {32'h3e320476, 32'h3ea922f5} /* (29, 19, 5) {real, imag} */,
  {32'h3f32866b, 32'h3f4e7484} /* (29, 19, 4) {real, imag} */,
  {32'hbfb2c330, 32'hbd7d7eb3} /* (29, 19, 3) {real, imag} */,
  {32'hc0494ed7, 32'hbedee00b} /* (29, 19, 2) {real, imag} */,
  {32'h3ee91e81, 32'h3ea7b2e1} /* (29, 19, 1) {real, imag} */,
  {32'hbf5977df, 32'hbfbcf13b} /* (29, 19, 0) {real, imag} */,
  {32'h3f673561, 32'hbf1a3c4e} /* (29, 18, 31) {real, imag} */,
  {32'hc03a8403, 32'hbf289af3} /* (29, 18, 30) {real, imag} */,
  {32'hbed08289, 32'h3f83168c} /* (29, 18, 29) {real, imag} */,
  {32'h3f7ecba1, 32'h3ff2303a} /* (29, 18, 28) {real, imag} */,
  {32'hc02449b0, 32'h3fd512b8} /* (29, 18, 27) {real, imag} */,
  {32'hbf1c6b34, 32'h401bf9dc} /* (29, 18, 26) {real, imag} */,
  {32'hbf02c8a5, 32'hc01e70f1} /* (29, 18, 25) {real, imag} */,
  {32'hbf51cc45, 32'hbe579328} /* (29, 18, 24) {real, imag} */,
  {32'h3fafd817, 32'h3ef1a359} /* (29, 18, 23) {real, imag} */,
  {32'hbdbb3b8c, 32'hc02717d6} /* (29, 18, 22) {real, imag} */,
  {32'hbe754814, 32'h3fa3b26f} /* (29, 18, 21) {real, imag} */,
  {32'h3e8061bc, 32'h3fcdd507} /* (29, 18, 20) {real, imag} */,
  {32'hc0058451, 32'hbfa56953} /* (29, 18, 19) {real, imag} */,
  {32'hbf620dfb, 32'h3e4c9218} /* (29, 18, 18) {real, imag} */,
  {32'h3f26a8e0, 32'hbf0a8ec2} /* (29, 18, 17) {real, imag} */,
  {32'hbe9e9381, 32'h3f239fde} /* (29, 18, 16) {real, imag} */,
  {32'hc00966a3, 32'h3fe83a17} /* (29, 18, 15) {real, imag} */,
  {32'hbe8972f2, 32'h3ebee70b} /* (29, 18, 14) {real, imag} */,
  {32'hc00438fa, 32'hc0023de7} /* (29, 18, 13) {real, imag} */,
  {32'h3fde4a4e, 32'h3dbc5896} /* (29, 18, 12) {real, imag} */,
  {32'hbc7913de, 32'hc023f77c} /* (29, 18, 11) {real, imag} */,
  {32'h4008c0c8, 32'hbf3b67f7} /* (29, 18, 10) {real, imag} */,
  {32'hbfbd0880, 32'hbfd68714} /* (29, 18, 9) {real, imag} */,
  {32'h3fee803e, 32'hbf4fefa6} /* (29, 18, 8) {real, imag} */,
  {32'h3fc05634, 32'hbee1a1a3} /* (29, 18, 7) {real, imag} */,
  {32'h3f2b225b, 32'h3f6cd580} /* (29, 18, 6) {real, imag} */,
  {32'hbff85413, 32'hbf4368e3} /* (29, 18, 5) {real, imag} */,
  {32'h3f50a0ab, 32'h3f3db0b2} /* (29, 18, 4) {real, imag} */,
  {32'hbe8df4b0, 32'h3ebb022d} /* (29, 18, 3) {real, imag} */,
  {32'hbff33bd2, 32'hbf850070} /* (29, 18, 2) {real, imag} */,
  {32'h401a4490, 32'hbf42ce48} /* (29, 18, 1) {real, imag} */,
  {32'h3ee24657, 32'h3f1f3b1d} /* (29, 18, 0) {real, imag} */,
  {32'hbfc2ee23, 32'hbf8d7b80} /* (29, 17, 31) {real, imag} */,
  {32'h4082c94f, 32'hbf6eb0c0} /* (29, 17, 30) {real, imag} */,
  {32'h3cb5cdad, 32'hbf80074e} /* (29, 17, 29) {real, imag} */,
  {32'hbf011f08, 32'h3fb17fde} /* (29, 17, 28) {real, imag} */,
  {32'hbff032f4, 32'hbfa4a978} /* (29, 17, 27) {real, imag} */,
  {32'h3f7522f6, 32'h3e0ebe80} /* (29, 17, 26) {real, imag} */,
  {32'hbf3f90e2, 32'h3f3b91f3} /* (29, 17, 25) {real, imag} */,
  {32'hbf905e43, 32'hbdfaf710} /* (29, 17, 24) {real, imag} */,
  {32'h3e9f04b7, 32'hbfb4a5ef} /* (29, 17, 23) {real, imag} */,
  {32'hbf5639d0, 32'h3ef3feb7} /* (29, 17, 22) {real, imag} */,
  {32'h3e036e4c, 32'hc042f3fb} /* (29, 17, 21) {real, imag} */,
  {32'h3f49c3cc, 32'h3e09c72b} /* (29, 17, 20) {real, imag} */,
  {32'h3f9d2975, 32'h3fa3ad7d} /* (29, 17, 19) {real, imag} */,
  {32'h3dfb7a8b, 32'hbfbb5699} /* (29, 17, 18) {real, imag} */,
  {32'h3ed5d220, 32'h3eb511e7} /* (29, 17, 17) {real, imag} */,
  {32'hbfa85a60, 32'hbed881c4} /* (29, 17, 16) {real, imag} */,
  {32'h3f8695b4, 32'hbf10414c} /* (29, 17, 15) {real, imag} */,
  {32'hbed8e380, 32'hbfadb8fc} /* (29, 17, 14) {real, imag} */,
  {32'hbfa951ee, 32'hbe4fcd1f} /* (29, 17, 13) {real, imag} */,
  {32'hbf1f3c3d, 32'h3fe33c5e} /* (29, 17, 12) {real, imag} */,
  {32'h400569f4, 32'h3ec98163} /* (29, 17, 11) {real, imag} */,
  {32'hc07f57c6, 32'h401840e3} /* (29, 17, 10) {real, imag} */,
  {32'h3ef70fc1, 32'h3f49e99c} /* (29, 17, 9) {real, imag} */,
  {32'hbfacdaf1, 32'hbf1fdcd8} /* (29, 17, 8) {real, imag} */,
  {32'hbe3b8c07, 32'hbfbe9a41} /* (29, 17, 7) {real, imag} */,
  {32'hbfb5b1a1, 32'h3f8059d0} /* (29, 17, 6) {real, imag} */,
  {32'h3decdbae, 32'hbd9d0677} /* (29, 17, 5) {real, imag} */,
  {32'hbf488ad2, 32'hbebd3558} /* (29, 17, 4) {real, imag} */,
  {32'hbf7865ce, 32'hbf50679c} /* (29, 17, 3) {real, imag} */,
  {32'h40275438, 32'hbf2c5b78} /* (29, 17, 2) {real, imag} */,
  {32'hbfa762a9, 32'hbf44c9df} /* (29, 17, 1) {real, imag} */,
  {32'hbd32f800, 32'hbf0b13ee} /* (29, 17, 0) {real, imag} */,
  {32'hbe4a68b7, 32'h3f58ef6f} /* (29, 16, 31) {real, imag} */,
  {32'h3f34fe48, 32'h3ebb495d} /* (29, 16, 30) {real, imag} */,
  {32'hbfaae10f, 32'hbef2c36b} /* (29, 16, 29) {real, imag} */,
  {32'hbf94dd90, 32'h3fb97693} /* (29, 16, 28) {real, imag} */,
  {32'h3e79a41e, 32'hbf2ca988} /* (29, 16, 27) {real, imag} */,
  {32'h3e048498, 32'hbf483315} /* (29, 16, 26) {real, imag} */,
  {32'hbf4bb3fd, 32'h3ed5f114} /* (29, 16, 25) {real, imag} */,
  {32'h3f631e0b, 32'h3f4bce93} /* (29, 16, 24) {real, imag} */,
  {32'h3e544c41, 32'h3e16fd9a} /* (29, 16, 23) {real, imag} */,
  {32'hbd307ada, 32'h3e816f4d} /* (29, 16, 22) {real, imag} */,
  {32'hc0347a74, 32'hbecdf961} /* (29, 16, 21) {real, imag} */,
  {32'hbfa2127d, 32'hbee32dde} /* (29, 16, 20) {real, imag} */,
  {32'hbf4f9155, 32'hbf535912} /* (29, 16, 19) {real, imag} */,
  {32'h3f849911, 32'h3fab3f16} /* (29, 16, 18) {real, imag} */,
  {32'h3fd4d416, 32'h3e6a4452} /* (29, 16, 17) {real, imag} */,
  {32'h3e5e0899, 32'h3ee978f8} /* (29, 16, 16) {real, imag} */,
  {32'hbe8b0286, 32'h3ed385fa} /* (29, 16, 15) {real, imag} */,
  {32'h3faf79b2, 32'hbf3c4d7d} /* (29, 16, 14) {real, imag} */,
  {32'h3eb1b425, 32'hbf38d2d8} /* (29, 16, 13) {real, imag} */,
  {32'hbee98c1d, 32'hbf93ebec} /* (29, 16, 12) {real, imag} */,
  {32'hbf2e79b3, 32'h3f5c1159} /* (29, 16, 11) {real, imag} */,
  {32'hbf56aa10, 32'hbfd2987f} /* (29, 16, 10) {real, imag} */,
  {32'h3e978e9d, 32'hbee1c9b7} /* (29, 16, 9) {real, imag} */,
  {32'h3ff273fa, 32'h3fb763eb} /* (29, 16, 8) {real, imag} */,
  {32'hbf94058c, 32'hbf97ba66} /* (29, 16, 7) {real, imag} */,
  {32'h3e37ba2f, 32'h3f3c45c2} /* (29, 16, 6) {real, imag} */,
  {32'h3f0f254c, 32'h3f23846e} /* (29, 16, 5) {real, imag} */,
  {32'h3ec708bf, 32'h3db2de16} /* (29, 16, 4) {real, imag} */,
  {32'h3f8d257f, 32'hbfd14f91} /* (29, 16, 3) {real, imag} */,
  {32'h3e79f529, 32'h3ca8bed9} /* (29, 16, 2) {real, imag} */,
  {32'hbe44ba32, 32'h3dd32852} /* (29, 16, 1) {real, imag} */,
  {32'h3f4c1dc6, 32'h3fd43828} /* (29, 16, 0) {real, imag} */,
  {32'h404a11c4, 32'h3fd1936a} /* (29, 15, 31) {real, imag} */,
  {32'hbf3e848b, 32'hbeccc229} /* (29, 15, 30) {real, imag} */,
  {32'hc02b689f, 32'hbf89eef1} /* (29, 15, 29) {real, imag} */,
  {32'hbf1ee632, 32'h3e9b7c50} /* (29, 15, 28) {real, imag} */,
  {32'h3fb46db7, 32'h3d88787a} /* (29, 15, 27) {real, imag} */,
  {32'h3f765d32, 32'h3dded79f} /* (29, 15, 26) {real, imag} */,
  {32'h3f9fe945, 32'h3dbe7ecf} /* (29, 15, 25) {real, imag} */,
  {32'h3fa218fd, 32'hbda36cdc} /* (29, 15, 24) {real, imag} */,
  {32'h3f98b4b5, 32'h3e9b3de1} /* (29, 15, 23) {real, imag} */,
  {32'h3fa9427d, 32'h3f8bd9aa} /* (29, 15, 22) {real, imag} */,
  {32'hbf8b92f3, 32'h400242c2} /* (29, 15, 21) {real, imag} */,
  {32'hbfab9f40, 32'hc00c82d5} /* (29, 15, 20) {real, imag} */,
  {32'hbfdf5e4d, 32'hc0164642} /* (29, 15, 19) {real, imag} */,
  {32'hbfb0dd9d, 32'hbf9330a6} /* (29, 15, 18) {real, imag} */,
  {32'h3f42097b, 32'hbf5a7f06} /* (29, 15, 17) {real, imag} */,
  {32'hbff056f1, 32'hbe5b9e7f} /* (29, 15, 16) {real, imag} */,
  {32'hbf0541a3, 32'hbe4fddc1} /* (29, 15, 15) {real, imag} */,
  {32'hbb8b218b, 32'h40245f10} /* (29, 15, 14) {real, imag} */,
  {32'h3db821e8, 32'hbec0e8d2} /* (29, 15, 13) {real, imag} */,
  {32'hbf3ce433, 32'h3f171a69} /* (29, 15, 12) {real, imag} */,
  {32'hbb37cefe, 32'h3e16330e} /* (29, 15, 11) {real, imag} */,
  {32'hbfb53341, 32'hbf9f9211} /* (29, 15, 10) {real, imag} */,
  {32'h3e812acb, 32'h3fa267fd} /* (29, 15, 9) {real, imag} */,
  {32'hbf674865, 32'h3fa55e4b} /* (29, 15, 8) {real, imag} */,
  {32'h3f82c651, 32'h3f202b01} /* (29, 15, 7) {real, imag} */,
  {32'hbed4ea9e, 32'h3f5440ac} /* (29, 15, 6) {real, imag} */,
  {32'h3f64e83c, 32'hbf7f9281} /* (29, 15, 5) {real, imag} */,
  {32'hbe523f73, 32'h3fd5dda8} /* (29, 15, 4) {real, imag} */,
  {32'hbf26fa04, 32'hbedf2b3d} /* (29, 15, 3) {real, imag} */,
  {32'hbf309309, 32'hbef0af2b} /* (29, 15, 2) {real, imag} */,
  {32'h3f2390a4, 32'hbf373077} /* (29, 15, 1) {real, imag} */,
  {32'hbfded959, 32'hbf5c665c} /* (29, 15, 0) {real, imag} */,
  {32'hc04ebba2, 32'h3ffe631a} /* (29, 14, 31) {real, imag} */,
  {32'hbe93bb90, 32'hc030c050} /* (29, 14, 30) {real, imag} */,
  {32'hbfcf9644, 32'h3f167e11} /* (29, 14, 29) {real, imag} */,
  {32'hbe411eb4, 32'h3fa0a940} /* (29, 14, 28) {real, imag} */,
  {32'hbce7ddff, 32'hbdd08929} /* (29, 14, 27) {real, imag} */,
  {32'hbf9723d5, 32'hbe0fabe7} /* (29, 14, 26) {real, imag} */,
  {32'h4017085d, 32'hbf6831ce} /* (29, 14, 25) {real, imag} */,
  {32'hbf8007c4, 32'hc0536366} /* (29, 14, 24) {real, imag} */,
  {32'h3f16703a, 32'h3f9e327c} /* (29, 14, 23) {real, imag} */,
  {32'h3f525efa, 32'h3fdc9aa5} /* (29, 14, 22) {real, imag} */,
  {32'hc0600f28, 32'h3ee6ca44} /* (29, 14, 21) {real, imag} */,
  {32'hbe7d80fa, 32'h3f1d1d64} /* (29, 14, 20) {real, imag} */,
  {32'h3fb0006f, 32'h3faced48} /* (29, 14, 19) {real, imag} */,
  {32'hbf2e56e3, 32'h3fa2c76c} /* (29, 14, 18) {real, imag} */,
  {32'h3e97cb20, 32'h3f5023ff} /* (29, 14, 17) {real, imag} */,
  {32'h3fce004a, 32'h3e8820b0} /* (29, 14, 16) {real, imag} */,
  {32'hbf51acef, 32'h3f5022c9} /* (29, 14, 15) {real, imag} */,
  {32'hbfa021c1, 32'hbfac7201} /* (29, 14, 14) {real, imag} */,
  {32'h3fd3d4ef, 32'h3fafd71a} /* (29, 14, 13) {real, imag} */,
  {32'h3fae3eae, 32'hbf7ef999} /* (29, 14, 12) {real, imag} */,
  {32'h3f2fd6e0, 32'h40473a73} /* (29, 14, 11) {real, imag} */,
  {32'h3fc123bd, 32'h40211f79} /* (29, 14, 10) {real, imag} */,
  {32'hc07526b9, 32'h3f7e1eb6} /* (29, 14, 9) {real, imag} */,
  {32'h402a0056, 32'hbf165bac} /* (29, 14, 8) {real, imag} */,
  {32'h3f881e06, 32'h3f122bfb} /* (29, 14, 7) {real, imag} */,
  {32'hbeb7135e, 32'h3f067c63} /* (29, 14, 6) {real, imag} */,
  {32'h3fdb78cf, 32'h3da9545f} /* (29, 14, 5) {real, imag} */,
  {32'hbfa16c17, 32'h3e3eba11} /* (29, 14, 4) {real, imag} */,
  {32'hbed6ef37, 32'h3f3bcf4c} /* (29, 14, 3) {real, imag} */,
  {32'hbeb32c97, 32'hbfc5c6bb} /* (29, 14, 2) {real, imag} */,
  {32'hc00e0096, 32'hbf00e6a2} /* (29, 14, 1) {real, imag} */,
  {32'hc037dfcf, 32'hbf431e85} /* (29, 14, 0) {real, imag} */,
  {32'h40588c99, 32'hbff38cc2} /* (29, 13, 31) {real, imag} */,
  {32'h3e73835b, 32'h3f3499c3} /* (29, 13, 30) {real, imag} */,
  {32'h3fc609b4, 32'h3f847545} /* (29, 13, 29) {real, imag} */,
  {32'hbfc0001d, 32'h3f300a04} /* (29, 13, 28) {real, imag} */,
  {32'hbe8d18e7, 32'hbfb4f2e4} /* (29, 13, 27) {real, imag} */,
  {32'hbf5716c7, 32'hbfcb4fca} /* (29, 13, 26) {real, imag} */,
  {32'hbf7ce6c1, 32'h3f51049e} /* (29, 13, 25) {real, imag} */,
  {32'hbdf55df3, 32'h3f9ee859} /* (29, 13, 24) {real, imag} */,
  {32'h4077de13, 32'hc01efdbb} /* (29, 13, 23) {real, imag} */,
  {32'hbfdbf469, 32'h3f42aed8} /* (29, 13, 22) {real, imag} */,
  {32'hbf83214b, 32'hc0123cc2} /* (29, 13, 21) {real, imag} */,
  {32'hbf9710bb, 32'h3ee328be} /* (29, 13, 20) {real, imag} */,
  {32'hbeea7738, 32'hc01bf43a} /* (29, 13, 19) {real, imag} */,
  {32'h3f61f0fa, 32'hbeb82a6f} /* (29, 13, 18) {real, imag} */,
  {32'hbe5d751e, 32'hbef5d5bf} /* (29, 13, 17) {real, imag} */,
  {32'hbd9884a2, 32'hbfb8f4f5} /* (29, 13, 16) {real, imag} */,
  {32'hbf804f3b, 32'hbf1b8258} /* (29, 13, 15) {real, imag} */,
  {32'hbf40f0a1, 32'hbefba9d5} /* (29, 13, 14) {real, imag} */,
  {32'hbe8b9889, 32'hbfe2658d} /* (29, 13, 13) {real, imag} */,
  {32'hbfdc1b19, 32'hbe41f404} /* (29, 13, 12) {real, imag} */,
  {32'hbd455834, 32'h3e20ac2c} /* (29, 13, 11) {real, imag} */,
  {32'hbf74b723, 32'hbf4c333b} /* (29, 13, 10) {real, imag} */,
  {32'h3ff39d05, 32'h40267260} /* (29, 13, 9) {real, imag} */,
  {32'hc0307939, 32'hc065370e} /* (29, 13, 8) {real, imag} */,
  {32'h3ea529e5, 32'h3f899e6f} /* (29, 13, 7) {real, imag} */,
  {32'h3f32ba70, 32'hbf9cba1e} /* (29, 13, 6) {real, imag} */,
  {32'hbf59be1e, 32'hbeb1c8d4} /* (29, 13, 5) {real, imag} */,
  {32'hbf4d9128, 32'hbe3e4c90} /* (29, 13, 4) {real, imag} */,
  {32'hbf724e0e, 32'hbffff77d} /* (29, 13, 3) {real, imag} */,
  {32'hc03ac04e, 32'h3f46256e} /* (29, 13, 2) {real, imag} */,
  {32'hbe63a0f1, 32'h3e429669} /* (29, 13, 1) {real, imag} */,
  {32'hbf5c9b6f, 32'hbfb20ddb} /* (29, 13, 0) {real, imag} */,
  {32'hc01a98ae, 32'hc024b903} /* (29, 12, 31) {real, imag} */,
  {32'hc01433f8, 32'hbfc00f3e} /* (29, 12, 30) {real, imag} */,
  {32'h40863b71, 32'h3fdf89a9} /* (29, 12, 29) {real, imag} */,
  {32'h3f110b75, 32'h3eb5c29a} /* (29, 12, 28) {real, imag} */,
  {32'hbbdaf5d3, 32'h3eb109ab} /* (29, 12, 27) {real, imag} */,
  {32'hbec063de, 32'h3f26b9cf} /* (29, 12, 26) {real, imag} */,
  {32'h4067f208, 32'h3fc4a26d} /* (29, 12, 25) {real, imag} */,
  {32'h3d17670b, 32'hbf12a7d8} /* (29, 12, 24) {real, imag} */,
  {32'h3f2f721d, 32'h405b3252} /* (29, 12, 23) {real, imag} */,
  {32'hbd8f1fe1, 32'h3f2c8057} /* (29, 12, 22) {real, imag} */,
  {32'h3f966488, 32'h3fca9487} /* (29, 12, 21) {real, imag} */,
  {32'h3ee9985c, 32'h3e593939} /* (29, 12, 20) {real, imag} */,
  {32'hc03ca1eb, 32'h40164ade} /* (29, 12, 19) {real, imag} */,
  {32'h3f28f55b, 32'hbf458025} /* (29, 12, 18) {real, imag} */,
  {32'h3e36d29a, 32'hbfa18dbc} /* (29, 12, 17) {real, imag} */,
  {32'h3d946752, 32'h3e89e6c8} /* (29, 12, 16) {real, imag} */,
  {32'h3de4178f, 32'hc013ce90} /* (29, 12, 15) {real, imag} */,
  {32'h3ee22726, 32'h3fc8d36a} /* (29, 12, 14) {real, imag} */,
  {32'hbf87e13c, 32'h3ff92bfa} /* (29, 12, 13) {real, imag} */,
  {32'h3fc27083, 32'h401a3065} /* (29, 12, 12) {real, imag} */,
  {32'hbfd70437, 32'h3e8ec548} /* (29, 12, 11) {real, imag} */,
  {32'h4013ee33, 32'h3e03e858} /* (29, 12, 10) {real, imag} */,
  {32'h3d377092, 32'hbd26edaf} /* (29, 12, 9) {real, imag} */,
  {32'h4037589b, 32'hbe205053} /* (29, 12, 8) {real, imag} */,
  {32'hc0b931d4, 32'h402bfbf4} /* (29, 12, 7) {real, imag} */,
  {32'h3f9f1f45, 32'hbeed64bd} /* (29, 12, 6) {real, imag} */,
  {32'h3fcb5d26, 32'h3f205133} /* (29, 12, 5) {real, imag} */,
  {32'h3f04ee13, 32'hbf54018f} /* (29, 12, 4) {real, imag} */,
  {32'hbc15d4b2, 32'hbf213b10} /* (29, 12, 3) {real, imag} */,
  {32'h3ec8e986, 32'h4004f041} /* (29, 12, 2) {real, imag} */,
  {32'h3f0c58b2, 32'hbf892c06} /* (29, 12, 1) {real, imag} */,
  {32'h3febec95, 32'h3fb93cb3} /* (29, 12, 0) {real, imag} */,
  {32'hbf8f65e5, 32'h3fb766ee} /* (29, 11, 31) {real, imag} */,
  {32'h400acfb2, 32'hc095caf1} /* (29, 11, 30) {real, imag} */,
  {32'h3e9b52a0, 32'hbf685c64} /* (29, 11, 29) {real, imag} */,
  {32'hc04967a3, 32'hc03ebd41} /* (29, 11, 28) {real, imag} */,
  {32'h4011d379, 32'h3fca5d9e} /* (29, 11, 27) {real, imag} */,
  {32'hbfae1640, 32'h40094f11} /* (29, 11, 26) {real, imag} */,
  {32'hc02dd570, 32'h40077429} /* (29, 11, 25) {real, imag} */,
  {32'h401fb101, 32'h4041ab36} /* (29, 11, 24) {real, imag} */,
  {32'h3e675383, 32'h400ba37c} /* (29, 11, 23) {real, imag} */,
  {32'h3f86bdd3, 32'h3f641b1e} /* (29, 11, 22) {real, imag} */,
  {32'hbf504858, 32'hc0344af2} /* (29, 11, 21) {real, imag} */,
  {32'h3f706995, 32'hbf6c161d} /* (29, 11, 20) {real, imag} */,
  {32'hbfb255dc, 32'hbede9ee0} /* (29, 11, 19) {real, imag} */,
  {32'hc0217535, 32'hbf259d26} /* (29, 11, 18) {real, imag} */,
  {32'h3f8c2c92, 32'h3feb7d36} /* (29, 11, 17) {real, imag} */,
  {32'h3dee8838, 32'hbd2ddb5f} /* (29, 11, 16) {real, imag} */,
  {32'hbf3f051a, 32'hbfc05928} /* (29, 11, 15) {real, imag} */,
  {32'hc05626b4, 32'h400667ef} /* (29, 11, 14) {real, imag} */,
  {32'h3feba3b4, 32'h3f02890c} /* (29, 11, 13) {real, imag} */,
  {32'hbec3e153, 32'h402b8f5a} /* (29, 11, 12) {real, imag} */,
  {32'hc002dc43, 32'hbe1838a6} /* (29, 11, 11) {real, imag} */,
  {32'h40139faa, 32'hbea676c2} /* (29, 11, 10) {real, imag} */,
  {32'h3f23a9af, 32'hbfacb08a} /* (29, 11, 9) {real, imag} */,
  {32'hbd089bcc, 32'h3edb3540} /* (29, 11, 8) {real, imag} */,
  {32'hbe390945, 32'h3f24491b} /* (29, 11, 7) {real, imag} */,
  {32'h401fcbd3, 32'hc0429d41} /* (29, 11, 6) {real, imag} */,
  {32'hbfc5391b, 32'h3fbdb286} /* (29, 11, 5) {real, imag} */,
  {32'h403000f7, 32'hbe8ab97c} /* (29, 11, 4) {real, imag} */,
  {32'h406166c6, 32'hbea38925} /* (29, 11, 3) {real, imag} */,
  {32'h403619c6, 32'hbfa46289} /* (29, 11, 2) {real, imag} */,
  {32'hc05ece4f, 32'h3fe6b75e} /* (29, 11, 1) {real, imag} */,
  {32'hc05bfe06, 32'h4005d76c} /* (29, 11, 0) {real, imag} */,
  {32'h4068891e, 32'hbfd882d4} /* (29, 10, 31) {real, imag} */,
  {32'hc0ba47c1, 32'h4093c12e} /* (29, 10, 30) {real, imag} */,
  {32'hbd01198b, 32'hc02c7112} /* (29, 10, 29) {real, imag} */,
  {32'h3fdf16f1, 32'hc0c857b5} /* (29, 10, 28) {real, imag} */,
  {32'hc05bf3f1, 32'hbf6aafcb} /* (29, 10, 27) {real, imag} */,
  {32'hbe7c455b, 32'h3f035924} /* (29, 10, 26) {real, imag} */,
  {32'hc09e3d94, 32'hbe9e0f11} /* (29, 10, 25) {real, imag} */,
  {32'h401fd116, 32'h3f3b227e} /* (29, 10, 24) {real, imag} */,
  {32'hbfa0efef, 32'h3f01b3e3} /* (29, 10, 23) {real, imag} */,
  {32'hbf11ae5e, 32'hbfb0424e} /* (29, 10, 22) {real, imag} */,
  {32'h40616794, 32'h3f9fa4d2} /* (29, 10, 21) {real, imag} */,
  {32'hbe1199da, 32'hbfc98058} /* (29, 10, 20) {real, imag} */,
  {32'hbf9151e2, 32'h3c58370a} /* (29, 10, 19) {real, imag} */,
  {32'hc0448abf, 32'hbfdeee58} /* (29, 10, 18) {real, imag} */,
  {32'hbf398aff, 32'h3e1a7346} /* (29, 10, 17) {real, imag} */,
  {32'hbfb1e1b7, 32'hbe969af5} /* (29, 10, 16) {real, imag} */,
  {32'hbf5809b8, 32'h3f476f28} /* (29, 10, 15) {real, imag} */,
  {32'h3fb0e7f7, 32'hbfcafbbc} /* (29, 10, 14) {real, imag} */,
  {32'h40371cb5, 32'h40878ab1} /* (29, 10, 13) {real, imag} */,
  {32'hbedaf5d2, 32'hbfd68117} /* (29, 10, 12) {real, imag} */,
  {32'hbf0ed199, 32'hc0006cb9} /* (29, 10, 11) {real, imag} */,
  {32'h3fd00c92, 32'h3e43d882} /* (29, 10, 10) {real, imag} */,
  {32'h3ff701fe, 32'h405076fd} /* (29, 10, 9) {real, imag} */,
  {32'h3ed2e8d2, 32'hbfcfad12} /* (29, 10, 8) {real, imag} */,
  {32'hc050fbc9, 32'h3f6627d3} /* (29, 10, 7) {real, imag} */,
  {32'hc00afb57, 32'hbe93fa92} /* (29, 10, 6) {real, imag} */,
  {32'hc018eecf, 32'h40103dbd} /* (29, 10, 5) {real, imag} */,
  {32'hbf0cec6c, 32'h40901a8e} /* (29, 10, 4) {real, imag} */,
  {32'h40b6edaa, 32'h4068460f} /* (29, 10, 3) {real, imag} */,
  {32'h4056c07d, 32'h3e3d80d4} /* (29, 10, 2) {real, imag} */,
  {32'hbfcf2c1c, 32'h3e8f0960} /* (29, 10, 1) {real, imag} */,
  {32'h4019aa3c, 32'hc00fb0c7} /* (29, 10, 0) {real, imag} */,
  {32'h40d30aea, 32'h403317cf} /* (29, 9, 31) {real, imag} */,
  {32'hbfe81209, 32'h3f9983e8} /* (29, 9, 30) {real, imag} */,
  {32'h3fd4f7ff, 32'hbf18b9e0} /* (29, 9, 29) {real, imag} */,
  {32'h400bd30b, 32'h3fb355f8} /* (29, 9, 28) {real, imag} */,
  {32'hc08b7cb2, 32'h3ff506f6} /* (29, 9, 27) {real, imag} */,
  {32'h3f26fda4, 32'h3fedf074} /* (29, 9, 26) {real, imag} */,
  {32'h3dc88c71, 32'h3e878877} /* (29, 9, 25) {real, imag} */,
  {32'hbff66746, 32'hbdc05568} /* (29, 9, 24) {real, imag} */,
  {32'h402313f7, 32'h3f05fc8a} /* (29, 9, 23) {real, imag} */,
  {32'hbfa4a644, 32'h3e7df0a9} /* (29, 9, 22) {real, imag} */,
  {32'hc0000967, 32'h3f9d3222} /* (29, 9, 21) {real, imag} */,
  {32'hbda82ec8, 32'hc0500d4d} /* (29, 9, 20) {real, imag} */,
  {32'h408071ec, 32'h3ff1b9c8} /* (29, 9, 19) {real, imag} */,
  {32'hbf05f899, 32'h3f81fe11} /* (29, 9, 18) {real, imag} */,
  {32'h3f75cd59, 32'hc043e2b8} /* (29, 9, 17) {real, imag} */,
  {32'h3e8e6524, 32'hbfadc811} /* (29, 9, 16) {real, imag} */,
  {32'h40261193, 32'hbf163843} /* (29, 9, 15) {real, imag} */,
  {32'h3f6751d8, 32'hbfd1a2cf} /* (29, 9, 14) {real, imag} */,
  {32'hbff6497d, 32'hbf8c1629} /* (29, 9, 13) {real, imag} */,
  {32'h3c73b8ad, 32'hc021f5a8} /* (29, 9, 12) {real, imag} */,
  {32'hbf1b4cae, 32'hc008ef81} /* (29, 9, 11) {real, imag} */,
  {32'h3ff00d24, 32'h3fb95e19} /* (29, 9, 10) {real, imag} */,
  {32'h3eb7562a, 32'hbd246c66} /* (29, 9, 9) {real, imag} */,
  {32'hc023b575, 32'h3fce6c6d} /* (29, 9, 8) {real, imag} */,
  {32'hbf8ab9dd, 32'hc03d4cc5} /* (29, 9, 7) {real, imag} */,
  {32'hc0205876, 32'hbeef2ffd} /* (29, 9, 6) {real, imag} */,
  {32'h40025dde, 32'hbed854b6} /* (29, 9, 5) {real, imag} */,
  {32'hbfe2dd39, 32'h3f2bdc69} /* (29, 9, 4) {real, imag} */,
  {32'hbe9a7d33, 32'hbca68d07} /* (29, 9, 3) {real, imag} */,
  {32'hbd462a9f, 32'h40193ff0} /* (29, 9, 2) {real, imag} */,
  {32'hc02db620, 32'hc03d5a47} /* (29, 9, 1) {real, imag} */,
  {32'h3fbd1da9, 32'hbfffc696} /* (29, 9, 0) {real, imag} */,
  {32'h3f239ee9, 32'h4120d26f} /* (29, 8, 31) {real, imag} */,
  {32'h3f2408b6, 32'hc1052180} /* (29, 8, 30) {real, imag} */,
  {32'hc0d78b74, 32'hbf5a018d} /* (29, 8, 29) {real, imag} */,
  {32'h4050ef37, 32'h3fe6d226} /* (29, 8, 28) {real, imag} */,
  {32'hc0047e8f, 32'h4057981a} /* (29, 8, 27) {real, imag} */,
  {32'hbecd92d3, 32'h3f9cf727} /* (29, 8, 26) {real, imag} */,
  {32'h3f267825, 32'h40276162} /* (29, 8, 25) {real, imag} */,
  {32'hc027f2c8, 32'h3f06dda0} /* (29, 8, 24) {real, imag} */,
  {32'h3f7af86b, 32'h40a6cd17} /* (29, 8, 23) {real, imag} */,
  {32'h3fda9f9e, 32'hbf189195} /* (29, 8, 22) {real, imag} */,
  {32'hbf2e7e65, 32'h40151356} /* (29, 8, 21) {real, imag} */,
  {32'hbfa2d17d, 32'h3f4492a0} /* (29, 8, 20) {real, imag} */,
  {32'h3f7fbff1, 32'hbfc8e866} /* (29, 8, 19) {real, imag} */,
  {32'h3ed197cf, 32'hbf5231a9} /* (29, 8, 18) {real, imag} */,
  {32'h3fd43ab4, 32'h3eef01a9} /* (29, 8, 17) {real, imag} */,
  {32'hbed5d46e, 32'hbe92e09a} /* (29, 8, 16) {real, imag} */,
  {32'hc05556e2, 32'h3eb0ca37} /* (29, 8, 15) {real, imag} */,
  {32'h3f674755, 32'hbf9aa3e4} /* (29, 8, 14) {real, imag} */,
  {32'hc0192f1c, 32'hbf0b64f5} /* (29, 8, 13) {real, imag} */,
  {32'hbdd03108, 32'hbff91c23} /* (29, 8, 12) {real, imag} */,
  {32'h40a1dbf7, 32'hbf8fab7f} /* (29, 8, 11) {real, imag} */,
  {32'hbf1b6b9c, 32'h4099d531} /* (29, 8, 10) {real, imag} */,
  {32'hc04647a1, 32'hbfd53ee6} /* (29, 8, 9) {real, imag} */,
  {32'h3feaccaf, 32'h3ff7a712} /* (29, 8, 8) {real, imag} */,
  {32'h4065981d, 32'h3fdfa151} /* (29, 8, 7) {real, imag} */,
  {32'h405a6f54, 32'h3fa9b800} /* (29, 8, 6) {real, imag} */,
  {32'h3ed1ad44, 32'hc0acbf54} /* (29, 8, 5) {real, imag} */,
  {32'hbf7b7c0d, 32'hbfa2c5ea} /* (29, 8, 4) {real, imag} */,
  {32'h4023808f, 32'hc06aaa5a} /* (29, 8, 3) {real, imag} */,
  {32'h404b968b, 32'h400846c9} /* (29, 8, 2) {real, imag} */,
  {32'hc0a9e787, 32'h40a03b31} /* (29, 8, 1) {real, imag} */,
  {32'hbd176c8a, 32'h407c3f61} /* (29, 8, 0) {real, imag} */,
  {32'h3f8b9872, 32'hc087f436} /* (29, 7, 31) {real, imag} */,
  {32'h3e031459, 32'hbfc25400} /* (29, 7, 30) {real, imag} */,
  {32'h408793fd, 32'h403eeb1a} /* (29, 7, 29) {real, imag} */,
  {32'h40a21fcc, 32'h407aab26} /* (29, 7, 28) {real, imag} */,
  {32'hc003fea2, 32'hbfddff3f} /* (29, 7, 27) {real, imag} */,
  {32'h3f5f808a, 32'h3fbda42b} /* (29, 7, 26) {real, imag} */,
  {32'h3f01d1d1, 32'h40adf394} /* (29, 7, 25) {real, imag} */,
  {32'hbeeaf237, 32'h3fb04e84} /* (29, 7, 24) {real, imag} */,
  {32'hbf8b0bec, 32'hbf8efeea} /* (29, 7, 23) {real, imag} */,
  {32'hbffc3631, 32'h3f77eb87} /* (29, 7, 22) {real, imag} */,
  {32'h3facb872, 32'hc014ec57} /* (29, 7, 21) {real, imag} */,
  {32'h3e0fea22, 32'h405d6e45} /* (29, 7, 20) {real, imag} */,
  {32'h3f9f1402, 32'hbf107ce9} /* (29, 7, 19) {real, imag} */,
  {32'hbf9b1fd8, 32'hbfa3b318} /* (29, 7, 18) {real, imag} */,
  {32'hbea4098e, 32'h4033a229} /* (29, 7, 17) {real, imag} */,
  {32'hbffc8f02, 32'hbf66c8e7} /* (29, 7, 16) {real, imag} */,
  {32'h3f6c6876, 32'h3fb1085b} /* (29, 7, 15) {real, imag} */,
  {32'hbeecfead, 32'h3ee8a575} /* (29, 7, 14) {real, imag} */,
  {32'h3f25a7ea, 32'h3ff95b86} /* (29, 7, 13) {real, imag} */,
  {32'hbf891ff0, 32'hbfba7cf5} /* (29, 7, 12) {real, imag} */,
  {32'h3fd30c5b, 32'h3f5b5700} /* (29, 7, 11) {real, imag} */,
  {32'hc01f4648, 32'hc0102a09} /* (29, 7, 10) {real, imag} */,
  {32'h3fd55819, 32'hbfefc7f3} /* (29, 7, 9) {real, imag} */,
  {32'h3f616f30, 32'h40bad4d6} /* (29, 7, 8) {real, imag} */,
  {32'hbfa46db7, 32'h3f1b823b} /* (29, 7, 7) {real, imag} */,
  {32'hc0390e10, 32'hbff8addf} /* (29, 7, 6) {real, imag} */,
  {32'hc04c39d2, 32'hbfcd3a61} /* (29, 7, 5) {real, imag} */,
  {32'h4003a2d5, 32'hc04a54eb} /* (29, 7, 4) {real, imag} */,
  {32'h3f94e39a, 32'h400e2e11} /* (29, 7, 3) {real, imag} */,
  {32'hc0c581cd, 32'hc02708de} /* (29, 7, 2) {real, imag} */,
  {32'h40979fb9, 32'hc0da823d} /* (29, 7, 1) {real, imag} */,
  {32'h3ff0c19f, 32'hc0f16b33} /* (29, 7, 0) {real, imag} */,
  {32'h3fbd0033, 32'h3f8526ed} /* (29, 6, 31) {real, imag} */,
  {32'h3fa4570c, 32'h3f691bea} /* (29, 6, 30) {real, imag} */,
  {32'h407f5110, 32'h3fa67f5c} /* (29, 6, 29) {real, imag} */,
  {32'h400783f1, 32'hc06afb2d} /* (29, 6, 28) {real, imag} */,
  {32'h400f3c84, 32'hbf91377d} /* (29, 6, 27) {real, imag} */,
  {32'hbfb8f00c, 32'hbeabd345} /* (29, 6, 26) {real, imag} */,
  {32'h401c1439, 32'hc099b8ed} /* (29, 6, 25) {real, imag} */,
  {32'hbfb2a01c, 32'h3f374b37} /* (29, 6, 24) {real, imag} */,
  {32'hbf5d426d, 32'h3ed07e43} /* (29, 6, 23) {real, imag} */,
  {32'hbe124e47, 32'hc06a1d05} /* (29, 6, 22) {real, imag} */,
  {32'h3ee92302, 32'hbf1fff3f} /* (29, 6, 21) {real, imag} */,
  {32'hbf6d70de, 32'h3fa8dd03} /* (29, 6, 20) {real, imag} */,
  {32'hc014850c, 32'h404d6778} /* (29, 6, 19) {real, imag} */,
  {32'h3fb5906f, 32'h3eea608c} /* (29, 6, 18) {real, imag} */,
  {32'h3fe410c2, 32'h3f5f6214} /* (29, 6, 17) {real, imag} */,
  {32'hbeb56cbf, 32'h3f22c8a3} /* (29, 6, 16) {real, imag} */,
  {32'h3db04820, 32'h3f6b353f} /* (29, 6, 15) {real, imag} */,
  {32'hbfb9712d, 32'h3fba2898} /* (29, 6, 14) {real, imag} */,
  {32'hbfe44311, 32'h3e989ca2} /* (29, 6, 13) {real, imag} */,
  {32'h3eb05a8b, 32'hbe4aa71a} /* (29, 6, 12) {real, imag} */,
  {32'hbfff8106, 32'hc0819498} /* (29, 6, 11) {real, imag} */,
  {32'h3eebc1fb, 32'h3e0095f1} /* (29, 6, 10) {real, imag} */,
  {32'hc08f3d36, 32'h405a82a9} /* (29, 6, 9) {real, imag} */,
  {32'h407e06ba, 32'hbfad576e} /* (29, 6, 8) {real, imag} */,
  {32'hc067987d, 32'hc07a6bf3} /* (29, 6, 7) {real, imag} */,
  {32'h40058633, 32'hc0b41a1f} /* (29, 6, 6) {real, imag} */,
  {32'h3ff69762, 32'hbf55db08} /* (29, 6, 5) {real, imag} */,
  {32'h40641de8, 32'hbfcae0a0} /* (29, 6, 4) {real, imag} */,
  {32'h3fbc5b66, 32'hbe95a4fa} /* (29, 6, 3) {real, imag} */,
  {32'hc011bdef, 32'h40108219} /* (29, 6, 2) {real, imag} */,
  {32'hbe510fc5, 32'h40805452} /* (29, 6, 1) {real, imag} */,
  {32'h40296a32, 32'h408b4469} /* (29, 6, 0) {real, imag} */,
  {32'hbfa53227, 32'h415f877d} /* (29, 5, 31) {real, imag} */,
  {32'hc104dcb9, 32'hc0d7ca2a} /* (29, 5, 30) {real, imag} */,
  {32'hbf4bedf7, 32'hbfa76212} /* (29, 5, 29) {real, imag} */,
  {32'h4042e185, 32'h4087bcf0} /* (29, 5, 28) {real, imag} */,
  {32'hc09f7f55, 32'hc0c9d929} /* (29, 5, 27) {real, imag} */,
  {32'h3faa53cc, 32'h3fa0d492} /* (29, 5, 26) {real, imag} */,
  {32'h4065f808, 32'h3f62a152} /* (29, 5, 25) {real, imag} */,
  {32'h4018534e, 32'hc05473d5} /* (29, 5, 24) {real, imag} */,
  {32'h3f95e49e, 32'h3f4bca09} /* (29, 5, 23) {real, imag} */,
  {32'hc0009519, 32'hbef07d34} /* (29, 5, 22) {real, imag} */,
  {32'hbed9d6fd, 32'hbfc56f45} /* (29, 5, 21) {real, imag} */,
  {32'hbf7f3e07, 32'h3f052055} /* (29, 5, 20) {real, imag} */,
  {32'h3f80ea06, 32'h3f964e86} /* (29, 5, 19) {real, imag} */,
  {32'hbf8e5633, 32'h3fc5ef5e} /* (29, 5, 18) {real, imag} */,
  {32'h3f740595, 32'hbf7e7b2a} /* (29, 5, 17) {real, imag} */,
  {32'hbf294277, 32'h3ea059ab} /* (29, 5, 16) {real, imag} */,
  {32'h3eaadfd5, 32'hbfe665ec} /* (29, 5, 15) {real, imag} */,
  {32'h3f694081, 32'h3e9836f1} /* (29, 5, 14) {real, imag} */,
  {32'h402050d3, 32'hbeeb67fe} /* (29, 5, 13) {real, imag} */,
  {32'hbf819448, 32'h3f8a5e8b} /* (29, 5, 12) {real, imag} */,
  {32'hbfbea8f2, 32'hbf27930c} /* (29, 5, 11) {real, imag} */,
  {32'hbf295958, 32'h401c97ca} /* (29, 5, 10) {real, imag} */,
  {32'h3eadb976, 32'h40054f4c} /* (29, 5, 9) {real, imag} */,
  {32'hbf1600ea, 32'h3ed4f729} /* (29, 5, 8) {real, imag} */,
  {32'h400f4e6f, 32'hc0843d78} /* (29, 5, 7) {real, imag} */,
  {32'hbffcbf33, 32'hbf854e73} /* (29, 5, 6) {real, imag} */,
  {32'h410c5983, 32'hc07e87c5} /* (29, 5, 5) {real, imag} */,
  {32'hc04e22fb, 32'h4080e270} /* (29, 5, 4) {real, imag} */,
  {32'hbed3f32b, 32'h4016d08d} /* (29, 5, 3) {real, imag} */,
  {32'h402ee25d, 32'hc0a42b00} /* (29, 5, 2) {real, imag} */,
  {32'hc118768c, 32'h4107a8d0} /* (29, 5, 1) {real, imag} */,
  {32'h409b5e1d, 32'h418c1f9a} /* (29, 5, 0) {real, imag} */,
  {32'h41450b21, 32'hc0dd6827} /* (29, 4, 31) {real, imag} */,
  {32'hc158e69e, 32'h4195de58} /* (29, 4, 30) {real, imag} */,
  {32'h3e7d10e7, 32'h3ce4c7f9} /* (29, 4, 29) {real, imag} */,
  {32'h400593b5, 32'hc00b72cf} /* (29, 4, 28) {real, imag} */,
  {32'hc033fb9b, 32'hbf7602bf} /* (29, 4, 27) {real, imag} */,
  {32'h40a2ae10, 32'hbee800ba} /* (29, 4, 26) {real, imag} */,
  {32'h404ddeff, 32'hbffd5c1d} /* (29, 4, 25) {real, imag} */,
  {32'hbeb0e402, 32'h40169c1d} /* (29, 4, 24) {real, imag} */,
  {32'h402815ff, 32'hc02f1676} /* (29, 4, 23) {real, imag} */,
  {32'hc0157474, 32'hc043f5ce} /* (29, 4, 22) {real, imag} */,
  {32'hc004e689, 32'h4014e404} /* (29, 4, 21) {real, imag} */,
  {32'hbf0ec1c5, 32'hbf996950} /* (29, 4, 20) {real, imag} */,
  {32'h3f8f9288, 32'hbf60340f} /* (29, 4, 19) {real, imag} */,
  {32'hbf74cb8f, 32'h403ff773} /* (29, 4, 18) {real, imag} */,
  {32'hbf15e826, 32'h3f027613} /* (29, 4, 17) {real, imag} */,
  {32'h3c0576be, 32'h3f76f8bc} /* (29, 4, 16) {real, imag} */,
  {32'h3fb7c8b5, 32'hbee34892} /* (29, 4, 15) {real, imag} */,
  {32'h3fe9f432, 32'h3ede3477} /* (29, 4, 14) {real, imag} */,
  {32'hbf1a3be3, 32'hc02275e9} /* (29, 4, 13) {real, imag} */,
  {32'hbf103123, 32'h3e511a02} /* (29, 4, 12) {real, imag} */,
  {32'hc01f68dd, 32'hbf745f9f} /* (29, 4, 11) {real, imag} */,
  {32'hbf2d1e44, 32'h4087b9b3} /* (29, 4, 10) {real, imag} */,
  {32'hbfaa4fc4, 32'h3fb510a6} /* (29, 4, 9) {real, imag} */,
  {32'hbfe27f1f, 32'hc00f6193} /* (29, 4, 8) {real, imag} */,
  {32'hbeaab2ff, 32'hc0dbef37} /* (29, 4, 7) {real, imag} */,
  {32'h402f992b, 32'hc08da8fa} /* (29, 4, 6) {real, imag} */,
  {32'h4080a58e, 32'hc0053475} /* (29, 4, 5) {real, imag} */,
  {32'h407c800b, 32'hbe1ab0b3} /* (29, 4, 4) {real, imag} */,
  {32'hc0007116, 32'h40b68917} /* (29, 4, 3) {real, imag} */,
  {32'hc0fd30dc, 32'h4197ed6d} /* (29, 4, 2) {real, imag} */,
  {32'h414f1384, 32'hc1f5161b} /* (29, 4, 1) {real, imag} */,
  {32'h412b451a, 32'hc0aaf819} /* (29, 4, 0) {real, imag} */,
  {32'h415b38a8, 32'h41d60566} /* (29, 3, 31) {real, imag} */,
  {32'hc1a5cc30, 32'hc0fba628} /* (29, 3, 30) {real, imag} */,
  {32'h3f4f8cb4, 32'hbf69a11a} /* (29, 3, 29) {real, imag} */,
  {32'h3f89ea0f, 32'hc09f186d} /* (29, 3, 28) {real, imag} */,
  {32'hc1006436, 32'h410f77e1} /* (29, 3, 27) {real, imag} */,
  {32'h3fc79d13, 32'hbf4a3453} /* (29, 3, 26) {real, imag} */,
  {32'h40bce19d, 32'h3ed36b08} /* (29, 3, 25) {real, imag} */,
  {32'hc003d391, 32'h40702555} /* (29, 3, 24) {real, imag} */,
  {32'h4028500d, 32'hc07ba9a5} /* (29, 3, 23) {real, imag} */,
  {32'hc0aabc6e, 32'hbfa031c5} /* (29, 3, 22) {real, imag} */,
  {32'h4035dbf5, 32'h3fe29b29} /* (29, 3, 21) {real, imag} */,
  {32'hbf9758b0, 32'hbf61e54c} /* (29, 3, 20) {real, imag} */,
  {32'h3fb1cfbb, 32'h3d24e6c0} /* (29, 3, 19) {real, imag} */,
  {32'h3f190b0c, 32'hbe465fa9} /* (29, 3, 18) {real, imag} */,
  {32'hbffa7a1c, 32'hbf5ce193} /* (29, 3, 17) {real, imag} */,
  {32'h3f88ed77, 32'h3f7b076b} /* (29, 3, 16) {real, imag} */,
  {32'h3f52faae, 32'hbf3b20ca} /* (29, 3, 15) {real, imag} */,
  {32'hbff9de2e, 32'hbf932d03} /* (29, 3, 14) {real, imag} */,
  {32'hbfd59ab9, 32'h3f6c7aac} /* (29, 3, 13) {real, imag} */,
  {32'h4005a478, 32'h40694227} /* (29, 3, 12) {real, imag} */,
  {32'hbe431877, 32'h3fe62129} /* (29, 3, 11) {real, imag} */,
  {32'h3fde6473, 32'h4056cb2f} /* (29, 3, 10) {real, imag} */,
  {32'h3f8ae3f0, 32'hc017846f} /* (29, 3, 9) {real, imag} */,
  {32'hc022cca5, 32'h40908aab} /* (29, 3, 8) {real, imag} */,
  {32'h40a92bba, 32'h3cb01ffc} /* (29, 3, 7) {real, imag} */,
  {32'hbdb91586, 32'h4035e84b} /* (29, 3, 6) {real, imag} */,
  {32'hc0c7a80a, 32'hbf8df81d} /* (29, 3, 5) {real, imag} */,
  {32'h40f5b294, 32'h3f84e2cc} /* (29, 3, 4) {real, imag} */,
  {32'h4040e80e, 32'hc0c09d7a} /* (29, 3, 3) {real, imag} */,
  {32'hc1ebd41e, 32'hbf29d3a3} /* (29, 3, 2) {real, imag} */,
  {32'h3f2d62c8, 32'hc1b9b95b} /* (29, 3, 1) {real, imag} */,
  {32'hc05d9b3d, 32'h40b2ffd9} /* (29, 3, 0) {real, imag} */,
  {32'h4194c473, 32'h42e58a99} /* (29, 2, 31) {real, imag} */,
  {32'hc2245837, 32'hc22f4217} /* (29, 2, 30) {real, imag} */,
  {32'h40d874a9, 32'hbf54f58e} /* (29, 2, 29) {real, imag} */,
  {32'h41236e3b, 32'h3f8aa78f} /* (29, 2, 28) {real, imag} */,
  {32'hc08e76cd, 32'hc0f8e770} /* (29, 2, 27) {real, imag} */,
  {32'h40030d2b, 32'hc0c94930} /* (29, 2, 26) {real, imag} */,
  {32'hbf91f0e0, 32'hc088e116} /* (29, 2, 25) {real, imag} */,
  {32'hc058ce96, 32'hc0da5840} /* (29, 2, 24) {real, imag} */,
  {32'hbfc83ae4, 32'hbf9dff91} /* (29, 2, 23) {real, imag} */,
  {32'hbf1db8d3, 32'h3f146883} /* (29, 2, 22) {real, imag} */,
  {32'hbfa0103a, 32'h3f0af5da} /* (29, 2, 21) {real, imag} */,
  {32'hbf48e669, 32'h3f3e4c58} /* (29, 2, 20) {real, imag} */,
  {32'hbf9b560e, 32'hbf045551} /* (29, 2, 19) {real, imag} */,
  {32'hc03b4e11, 32'hbf558f5c} /* (29, 2, 18) {real, imag} */,
  {32'hbf3f620b, 32'hc002edbe} /* (29, 2, 17) {real, imag} */,
  {32'h3d967779, 32'h3aa137b0} /* (29, 2, 16) {real, imag} */,
  {32'h3dc549cb, 32'h3e923cf3} /* (29, 2, 15) {real, imag} */,
  {32'h3f843619, 32'h4007737c} /* (29, 2, 14) {real, imag} */,
  {32'hbf5c8aa6, 32'h3f1a5cb9} /* (29, 2, 13) {real, imag} */,
  {32'h3ecf1a0f, 32'h3fa54d67} /* (29, 2, 12) {real, imag} */,
  {32'h4015fd27, 32'hc07da490} /* (29, 2, 11) {real, imag} */,
  {32'hbf50ca93, 32'h403b9e7d} /* (29, 2, 10) {real, imag} */,
  {32'h4058f7ed, 32'hc0918067} /* (29, 2, 9) {real, imag} */,
  {32'hc0c72788, 32'hc0a376ad} /* (29, 2, 8) {real, imag} */,
  {32'hc0b61a4a, 32'h40806ffc} /* (29, 2, 7) {real, imag} */,
  {32'hbfbe2f5c, 32'hc0578355} /* (29, 2, 6) {real, imag} */,
  {32'hc0f5717c, 32'hc116a8c5} /* (29, 2, 5) {real, imag} */,
  {32'h400ef944, 32'h41cc64b1} /* (29, 2, 4) {real, imag} */,
  {32'h407676ce, 32'hc08a4197} /* (29, 2, 3) {real, imag} */,
  {32'hc1ecc9da, 32'hc246c764} /* (29, 2, 2) {real, imag} */,
  {32'h41c9b592, 32'h428a68f0} /* (29, 2, 1) {real, imag} */,
  {32'hc09bbc3f, 32'h4298f038} /* (29, 2, 0) {real, imag} */,
  {32'hc287da1a, 32'hc2a18326} /* (29, 1, 31) {real, imag} */,
  {32'h4112c960, 32'h421f2440} /* (29, 1, 30) {real, imag} */,
  {32'hc110ec6c, 32'h4091a928} /* (29, 1, 29) {real, imag} */,
  {32'h405ceea8, 32'hc13ac18d} /* (29, 1, 28) {real, imag} */,
  {32'h412ee02a, 32'h4155195a} /* (29, 1, 27) {real, imag} */,
  {32'hbe3b91d1, 32'h40576db5} /* (29, 1, 26) {real, imag} */,
  {32'hbf92f272, 32'hc0f12eed} /* (29, 1, 25) {real, imag} */,
  {32'h40316663, 32'h407ed12c} /* (29, 1, 24) {real, imag} */,
  {32'h3e370693, 32'hc088d0c7} /* (29, 1, 23) {real, imag} */,
  {32'h401e0688, 32'h3f957027} /* (29, 1, 22) {real, imag} */,
  {32'h409b5841, 32'h40dc4b6c} /* (29, 1, 21) {real, imag} */,
  {32'hbef65b42, 32'hbf3cebfd} /* (29, 1, 20) {real, imag} */,
  {32'hbf0c5dcf, 32'hbfbd4055} /* (29, 1, 19) {real, imag} */,
  {32'h406f70d3, 32'h40025a78} /* (29, 1, 18) {real, imag} */,
  {32'h3f1630a9, 32'hbf0da003} /* (29, 1, 17) {real, imag} */,
  {32'h3f07853d, 32'h3fd6b7cb} /* (29, 1, 16) {real, imag} */,
  {32'h3ff6b0f8, 32'h3e2a66f6} /* (29, 1, 15) {real, imag} */,
  {32'hc08126ce, 32'h3f74d79c} /* (29, 1, 14) {real, imag} */,
  {32'h3f254958, 32'h3f0f8a12} /* (29, 1, 13) {real, imag} */,
  {32'h3f9648a7, 32'h3f96d530} /* (29, 1, 12) {real, imag} */,
  {32'hbf872020, 32'h3fbabbee} /* (29, 1, 11) {real, imag} */,
  {32'h3ee34bf7, 32'hbd6088e0} /* (29, 1, 10) {real, imag} */,
  {32'h4020d2df, 32'h3f17818a} /* (29, 1, 9) {real, imag} */,
  {32'hc0a729fe, 32'hbdb36117} /* (29, 1, 8) {real, imag} */,
  {32'h3ff0c035, 32'hc05f6f85} /* (29, 1, 7) {real, imag} */,
  {32'h40484aee, 32'h40844f2f} /* (29, 1, 6) {real, imag} */,
  {32'hc10fb5df, 32'h418ea5a3} /* (29, 1, 5) {real, imag} */,
  {32'hc090f8dd, 32'hc16d854f} /* (29, 1, 4) {real, imag} */,
  {32'h41946661, 32'h41927a72} /* (29, 1, 3) {real, imag} */,
  {32'hc21431e3, 32'h42934ac6} /* (29, 1, 2) {real, imag} */,
  {32'h41ffaae4, 32'hc339b71d} /* (29, 1, 1) {real, imag} */,
  {32'hc187b308, 32'hc2f1e859} /* (29, 1, 0) {real, imag} */,
  {32'hc28e7e07, 32'hc289abac} /* (29, 0, 31) {real, imag} */,
  {32'h41a48bbe, 32'h40572dd9} /* (29, 0, 30) {real, imag} */,
  {32'hc131d470, 32'h41984692} /* (29, 0, 29) {real, imag} */,
  {32'h412f7f39, 32'h3ff187ea} /* (29, 0, 28) {real, imag} */,
  {32'h416a7091, 32'h4133b17c} /* (29, 0, 27) {real, imag} */,
  {32'hc10fe016, 32'hc01d2c13} /* (29, 0, 26) {real, imag} */,
  {32'hc0c2bbe2, 32'h40db86dd} /* (29, 0, 25) {real, imag} */,
  {32'h408531ba, 32'h3f826c82} /* (29, 0, 24) {real, imag} */,
  {32'h3f6ef582, 32'h3fc5057f} /* (29, 0, 23) {real, imag} */,
  {32'h40960c17, 32'hc036364e} /* (29, 0, 22) {real, imag} */,
  {32'h4014b00d, 32'hbf8f131d} /* (29, 0, 21) {real, imag} */,
  {32'hc0831a9d, 32'hbe2dfe7c} /* (29, 0, 20) {real, imag} */,
  {32'hbf27a437, 32'hc04c0374} /* (29, 0, 19) {real, imag} */,
  {32'h3fdf6a58, 32'hc0585fcc} /* (29, 0, 18) {real, imag} */,
  {32'hbfd09e88, 32'hbf0cadb8} /* (29, 0, 17) {real, imag} */,
  {32'hbecafaff, 32'h3fad3113} /* (29, 0, 16) {real, imag} */,
  {32'hbf10ad08, 32'h3fa08fc0} /* (29, 0, 15) {real, imag} */,
  {32'h3e9bce9e, 32'h3ff4208b} /* (29, 0, 14) {real, imag} */,
  {32'hbe83853f, 32'h3f41b6b2} /* (29, 0, 13) {real, imag} */,
  {32'h3ff2d6c4, 32'hc0179a91} /* (29, 0, 12) {real, imag} */,
  {32'hbeb31e99, 32'h401efc6a} /* (29, 0, 11) {real, imag} */,
  {32'h3fadff49, 32'hc0196d95} /* (29, 0, 10) {real, imag} */,
  {32'h3f60c307, 32'hc04d9cd9} /* (29, 0, 9) {real, imag} */,
  {32'hc08369a4, 32'hc01527fe} /* (29, 0, 8) {real, imag} */,
  {32'h4085c387, 32'hc02ef542} /* (29, 0, 7) {real, imag} */,
  {32'hc08cb2df, 32'h4027c2ac} /* (29, 0, 6) {real, imag} */,
  {32'h4092e3ce, 32'h414aeba8} /* (29, 0, 5) {real, imag} */,
  {32'hc17286fd, 32'h3f8b7f3e} /* (29, 0, 4) {real, imag} */,
  {32'hc16924d5, 32'h400e3985} /* (29, 0, 3) {real, imag} */,
  {32'hc1b61ee2, 32'h41b35bfc} /* (29, 0, 2) {real, imag} */,
  {32'h4269be17, 32'hc2acb596} /* (29, 0, 1) {real, imag} */,
  {32'hc1f2f479, 32'hc2797e12} /* (29, 0, 0) {real, imag} */,
  {32'hc2a2aa6d, 32'hc2805593} /* (28, 31, 31) {real, imag} */,
  {32'h4273320d, 32'h417c37e8} /* (28, 31, 30) {real, imag} */,
  {32'hc009aebc, 32'h412060b2} /* (28, 31, 29) {real, imag} */,
  {32'hc0012445, 32'h3f3de2c2} /* (28, 31, 28) {real, imag} */,
  {32'h413448a3, 32'h40e0e8ab} /* (28, 31, 27) {real, imag} */,
  {32'h409c706f, 32'hc044e51c} /* (28, 31, 26) {real, imag} */,
  {32'hbf6cce40, 32'h3e876091} /* (28, 31, 25) {real, imag} */,
  {32'h40d90411, 32'h3ea579ca} /* (28, 31, 24) {real, imag} */,
  {32'h40147b07, 32'hc03d9252} /* (28, 31, 23) {real, imag} */,
  {32'hbfde5996, 32'h400a8812} /* (28, 31, 22) {real, imag} */,
  {32'h402b2cad, 32'h3f4b5145} /* (28, 31, 21) {real, imag} */,
  {32'hbd4c28e7, 32'h4022a943} /* (28, 31, 20) {real, imag} */,
  {32'hbf4f52d2, 32'h3f112b16} /* (28, 31, 19) {real, imag} */,
  {32'h3e6d7d40, 32'hbfbc7029} /* (28, 31, 18) {real, imag} */,
  {32'hbfe7244e, 32'h3fcfdb2c} /* (28, 31, 17) {real, imag} */,
  {32'h3ff1b942, 32'hbf59a416} /* (28, 31, 16) {real, imag} */,
  {32'hbf3b3760, 32'h3eb46be6} /* (28, 31, 15) {real, imag} */,
  {32'hc064db7c, 32'hbe8ab14c} /* (28, 31, 14) {real, imag} */,
  {32'hbfcf6a6a, 32'hbf2647fc} /* (28, 31, 13) {real, imag} */,
  {32'h40939630, 32'hbfaca6e8} /* (28, 31, 12) {real, imag} */,
  {32'hc10e6297, 32'h40b68869} /* (28, 31, 11) {real, imag} */,
  {32'h3f0a3475, 32'hbfd88f48} /* (28, 31, 10) {real, imag} */,
  {32'h3e9aa20a, 32'hbef528e8} /* (28, 31, 9) {real, imag} */,
  {32'hc04b0976, 32'h40d8bdd4} /* (28, 31, 8) {real, imag} */,
  {32'h4098dac9, 32'hbf511f23} /* (28, 31, 7) {real, imag} */,
  {32'hc08b297c, 32'hc04fa4d0} /* (28, 31, 6) {real, imag} */,
  {32'h40f7fd93, 32'h419d40e3} /* (28, 31, 5) {real, imag} */,
  {32'hc033a82e, 32'hc14c6779} /* (28, 31, 4) {real, imag} */,
  {32'hbf616836, 32'hc0f36c88} /* (28, 31, 3) {real, imag} */,
  {32'h413ecfd2, 32'h41e14199} /* (28, 31, 2) {real, imag} */,
  {32'hc0391f02, 32'hc2848756} /* (28, 31, 1) {real, imag} */,
  {32'hc242fdcf, 32'hc2655ace} /* (28, 31, 0) {real, imag} */,
  {32'h40f21c1a, 32'h422f8b17} /* (28, 30, 31) {real, imag} */,
  {32'hbed63da6, 32'hc2090cdb} /* (28, 30, 30) {real, imag} */,
  {32'h404847a9, 32'h40ced8c3} /* (28, 30, 29) {real, imag} */,
  {32'hbff383fd, 32'h4117c94b} /* (28, 30, 28) {real, imag} */,
  {32'hc0f3c0ef, 32'hc10248da} /* (28, 30, 27) {real, imag} */,
  {32'hc0321fd8, 32'h3f8f70a1} /* (28, 30, 26) {real, imag} */,
  {32'h4056e43c, 32'h3f1b3850} /* (28, 30, 25) {real, imag} */,
  {32'hc056644a, 32'hc0c53aa0} /* (28, 30, 24) {real, imag} */,
  {32'hc03f6dea, 32'hbf6339b5} /* (28, 30, 23) {real, imag} */,
  {32'h3d0dd17a, 32'h400a8a19} /* (28, 30, 22) {real, imag} */,
  {32'hc0310ebe, 32'hbe58f34c} /* (28, 30, 21) {real, imag} */,
  {32'h3e6f6f84, 32'h400a52ec} /* (28, 30, 20) {real, imag} */,
  {32'h3ed39cea, 32'h3f75867f} /* (28, 30, 19) {real, imag} */,
  {32'hbff52692, 32'hc0379659} /* (28, 30, 18) {real, imag} */,
  {32'hbf7fa5d2, 32'h3f826fab} /* (28, 30, 17) {real, imag} */,
  {32'hbfc8505e, 32'hbf8b2399} /* (28, 30, 16) {real, imag} */,
  {32'hbea6b8e9, 32'h39dc551e} /* (28, 30, 15) {real, imag} */,
  {32'h3f2910be, 32'h3e89bcd4} /* (28, 30, 14) {real, imag} */,
  {32'h3e47920c, 32'hbea5855f} /* (28, 30, 13) {real, imag} */,
  {32'hbfc33504, 32'h3f8c2fa4} /* (28, 30, 12) {real, imag} */,
  {32'h40658017, 32'hc03530f2} /* (28, 30, 11) {real, imag} */,
  {32'hc08d7904, 32'hbf3de555} /* (28, 30, 10) {real, imag} */,
  {32'h400a6410, 32'hbf82cc7e} /* (28, 30, 9) {real, imag} */,
  {32'h3fdc27e3, 32'hc0fc2d8d} /* (28, 30, 8) {real, imag} */,
  {32'h3f43795b, 32'h400b0930} /* (28, 30, 7) {real, imag} */,
  {32'hc02c7ab4, 32'h4034fd57} /* (28, 30, 6) {real, imag} */,
  {32'h404ea0ce, 32'hc1065381} /* (28, 30, 5) {real, imag} */,
  {32'hc08cb6ee, 32'h41529b05} /* (28, 30, 4) {real, imag} */,
  {32'h40618cda, 32'h41168dc2} /* (28, 30, 3) {real, imag} */,
  {32'hc13c128f, 32'hc2468722} /* (28, 30, 2) {real, imag} */,
  {32'h4202aeb2, 32'h4295499b} /* (28, 30, 1) {real, imag} */,
  {32'h41b0c404, 32'h421e4bbc} /* (28, 30, 0) {real, imag} */,
  {32'hc17761d3, 32'h3fb4b744} /* (28, 29, 31) {real, imag} */,
  {32'h410ff4b0, 32'h3f99ecb4} /* (28, 29, 30) {real, imag} */,
  {32'hc0e2339b, 32'hbe63cc90} /* (28, 29, 29) {real, imag} */,
  {32'h4028bb93, 32'h3f06a61d} /* (28, 29, 28) {real, imag} */,
  {32'h3fe0ef12, 32'hc07193af} /* (28, 29, 27) {real, imag} */,
  {32'h3f929d97, 32'hc0b067e5} /* (28, 29, 26) {real, imag} */,
  {32'hc0b1e5a5, 32'hc0a86f08} /* (28, 29, 25) {real, imag} */,
  {32'h3e835fa0, 32'h3e929c85} /* (28, 29, 24) {real, imag} */,
  {32'h3fe227be, 32'h40051c41} /* (28, 29, 23) {real, imag} */,
  {32'hbf6e16c2, 32'h404c1b17} /* (28, 29, 22) {real, imag} */,
  {32'h3e015fbf, 32'hbfda031e} /* (28, 29, 21) {real, imag} */,
  {32'h3dc3bf9c, 32'h4020503d} /* (28, 29, 20) {real, imag} */,
  {32'hc02418d1, 32'hbf262597} /* (28, 29, 19) {real, imag} */,
  {32'hbf138d5c, 32'hbfc152f7} /* (28, 29, 18) {real, imag} */,
  {32'hbed0a859, 32'hbea95d13} /* (28, 29, 17) {real, imag} */,
  {32'hbe8c67a4, 32'hc0009711} /* (28, 29, 16) {real, imag} */,
  {32'hbfd16e68, 32'h403001d0} /* (28, 29, 15) {real, imag} */,
  {32'h3fb702e4, 32'hbfc5adf0} /* (28, 29, 14) {real, imag} */,
  {32'h40022d2b, 32'hbf6e8a9c} /* (28, 29, 13) {real, imag} */,
  {32'hc06e3c89, 32'hc006bace} /* (28, 29, 12) {real, imag} */,
  {32'h3fbd8b15, 32'h4064362b} /* (28, 29, 11) {real, imag} */,
  {32'hbf87a913, 32'hc00b4825} /* (28, 29, 10) {real, imag} */,
  {32'hc08cd733, 32'hbe8523d7} /* (28, 29, 9) {real, imag} */,
  {32'h3f4781fc, 32'hbfca1226} /* (28, 29, 8) {real, imag} */,
  {32'h3ffa16f1, 32'h4005e67a} /* (28, 29, 7) {real, imag} */,
  {32'h3d5a7b3c, 32'h3fbb473b} /* (28, 29, 6) {real, imag} */,
  {32'h402fe671, 32'hc08da99c} /* (28, 29, 5) {real, imag} */,
  {32'hc036eac3, 32'h4054920d} /* (28, 29, 4) {real, imag} */,
  {32'h3fec68c3, 32'hc0a2d561} /* (28, 29, 3) {real, imag} */,
  {32'h415dd7c4, 32'hc1242df6} /* (28, 29, 2) {real, imag} */,
  {32'h3fdc962d, 32'h4195b01c} /* (28, 29, 1) {real, imag} */,
  {32'h3fe52126, 32'h3f8d7d16} /* (28, 29, 0) {real, imag} */,
  {32'hc17f0f95, 32'hc1c55b5a} /* (28, 28, 31) {real, imag} */,
  {32'h41708f1e, 32'h4082c799} /* (28, 28, 30) {real, imag} */,
  {32'hc0213521, 32'hc09431cd} /* (28, 28, 29) {real, imag} */,
  {32'hc08b4c23, 32'h3f9bcfa0} /* (28, 28, 28) {real, imag} */,
  {32'h3df37b9b, 32'h3f3abe2d} /* (28, 28, 27) {real, imag} */,
  {32'h40493917, 32'h4069414b} /* (28, 28, 26) {real, imag} */,
  {32'hc044de01, 32'hbf873b32} /* (28, 28, 25) {real, imag} */,
  {32'h40122a80, 32'h3df0d213} /* (28, 28, 24) {real, imag} */,
  {32'h404ad63d, 32'hc03cc251} /* (28, 28, 23) {real, imag} */,
  {32'h3f47164e, 32'h3fceeec5} /* (28, 28, 22) {real, imag} */,
  {32'h3ff49769, 32'hbf285f7b} /* (28, 28, 21) {real, imag} */,
  {32'hbf0fa309, 32'h3efc582a} /* (28, 28, 20) {real, imag} */,
  {32'h406ce146, 32'hbf73d46b} /* (28, 28, 19) {real, imag} */,
  {32'h3f4d997b, 32'h3f7aa0a6} /* (28, 28, 18) {real, imag} */,
  {32'h3f15d200, 32'h3d099f7a} /* (28, 28, 17) {real, imag} */,
  {32'h3ee2f0bd, 32'h3efb5d21} /* (28, 28, 16) {real, imag} */,
  {32'hbf94d277, 32'h3eadb9c8} /* (28, 28, 15) {real, imag} */,
  {32'hbefddd7d, 32'hbf38e123} /* (28, 28, 14) {real, imag} */,
  {32'hbfc89136, 32'hc03a7128} /* (28, 28, 13) {real, imag} */,
  {32'h3acd0892, 32'hbf59c098} /* (28, 28, 12) {real, imag} */,
  {32'h3fce843c, 32'h4003daa3} /* (28, 28, 11) {real, imag} */,
  {32'hbf93486b, 32'hbf8f6941} /* (28, 28, 10) {real, imag} */,
  {32'h4063e850, 32'h3fdb589a} /* (28, 28, 9) {real, imag} */,
  {32'hbf686f11, 32'h3f8aa181} /* (28, 28, 8) {real, imag} */,
  {32'hc07aa49a, 32'h3e1775a2} /* (28, 28, 7) {real, imag} */,
  {32'h4022a9ca, 32'hc0301058} /* (28, 28, 6) {real, imag} */,
  {32'hbe838c20, 32'h40a0ff43} /* (28, 28, 5) {real, imag} */,
  {32'hc1474531, 32'hc0e2b654} /* (28, 28, 4) {real, imag} */,
  {32'hc04cbbe0, 32'h40a030b9} /* (28, 28, 3) {real, imag} */,
  {32'h414abae3, 32'hc0369d72} /* (28, 28, 2) {real, imag} */,
  {32'hc174f041, 32'hc12dee90} /* (28, 28, 1) {real, imag} */,
  {32'hc0db90c1, 32'hc062319f} /* (28, 28, 0) {real, imag} */,
  {32'h41425323, 32'h40b0aa2b} /* (28, 27, 31) {real, imag} */,
  {32'hc094879a, 32'hc08c62be} /* (28, 27, 30) {real, imag} */,
  {32'hc0746d4c, 32'hbf59642e} /* (28, 27, 29) {real, imag} */,
  {32'hc039dd74, 32'hbfae8f0b} /* (28, 27, 28) {real, imag} */,
  {32'h3cd622be, 32'hbf396928} /* (28, 27, 27) {real, imag} */,
  {32'hbfc3a1d2, 32'hc0f18960} /* (28, 27, 26) {real, imag} */,
  {32'h3fb1c5f8, 32'h3e9a601d} /* (28, 27, 25) {real, imag} */,
  {32'h3f241ad8, 32'h403a7b93} /* (28, 27, 24) {real, imag} */,
  {32'hc031be0e, 32'h3e931244} /* (28, 27, 23) {real, imag} */,
  {32'h3ee65f48, 32'h408a34b3} /* (28, 27, 22) {real, imag} */,
  {32'hbfc93fe1, 32'hbf059275} /* (28, 27, 21) {real, imag} */,
  {32'h3e98f05f, 32'hbe6faaf9} /* (28, 27, 20) {real, imag} */,
  {32'h3ff2028b, 32'h3e8f6aab} /* (28, 27, 19) {real, imag} */,
  {32'h3f0bcf74, 32'h3eaf5479} /* (28, 27, 18) {real, imag} */,
  {32'h3edd8c4d, 32'h3e65d09a} /* (28, 27, 17) {real, imag} */,
  {32'h3f687a3d, 32'h3ecc82c3} /* (28, 27, 16) {real, imag} */,
  {32'hbf2c3805, 32'hbc955d1e} /* (28, 27, 15) {real, imag} */,
  {32'h3f6a543c, 32'hbfa86e68} /* (28, 27, 14) {real, imag} */,
  {32'h4087d218, 32'h3f573a3a} /* (28, 27, 13) {real, imag} */,
  {32'h3dc9a26b, 32'h401e3010} /* (28, 27, 12) {real, imag} */,
  {32'hbf91d970, 32'hc011ef71} /* (28, 27, 11) {real, imag} */,
  {32'hbf18d197, 32'h3f2528de} /* (28, 27, 10) {real, imag} */,
  {32'h3fd4f557, 32'h3f81a135} /* (28, 27, 9) {real, imag} */,
  {32'hbf767709, 32'h3fed0b80} /* (28, 27, 8) {real, imag} */,
  {32'hc073f349, 32'h408d0571} /* (28, 27, 7) {real, imag} */,
  {32'hbf01d6e2, 32'h3e0bbbdf} /* (28, 27, 6) {real, imag} */,
  {32'hc002ad9a, 32'hc098a706} /* (28, 27, 5) {real, imag} */,
  {32'h40be5549, 32'h401f5275} /* (28, 27, 4) {real, imag} */,
  {32'h401b2a21, 32'h3f2e7c37} /* (28, 27, 3) {real, imag} */,
  {32'hbef3f08f, 32'hc02a723c} /* (28, 27, 2) {real, imag} */,
  {32'h4016f3b3, 32'h410013c3} /* (28, 27, 1) {real, imag} */,
  {32'h40dde50e, 32'h40c1c34a} /* (28, 27, 0) {real, imag} */,
  {32'hbf870635, 32'h403be1cd} /* (28, 26, 31) {real, imag} */,
  {32'hc0584f04, 32'h409755f6} /* (28, 26, 30) {real, imag} */,
  {32'h3ebd04bb, 32'hbfd1c5e1} /* (28, 26, 29) {real, imag} */,
  {32'h3fe13c31, 32'h3f01e0f1} /* (28, 26, 28) {real, imag} */,
  {32'h3fe89a5d, 32'hbfba08ac} /* (28, 26, 27) {real, imag} */,
  {32'hbe4a8a10, 32'h407b7110} /* (28, 26, 26) {real, imag} */,
  {32'hbd7878f6, 32'h3fd2741a} /* (28, 26, 25) {real, imag} */,
  {32'h3f9ab373, 32'hbff48743} /* (28, 26, 24) {real, imag} */,
  {32'h402138d3, 32'h3fbe7e35} /* (28, 26, 23) {real, imag} */,
  {32'hbf1d800e, 32'hc005c35c} /* (28, 26, 22) {real, imag} */,
  {32'hc0194e3e, 32'h3f5dcfd7} /* (28, 26, 21) {real, imag} */,
  {32'hbfc2014f, 32'hbffff70a} /* (28, 26, 20) {real, imag} */,
  {32'hbf20c614, 32'h3fdadb42} /* (28, 26, 19) {real, imag} */,
  {32'hbfa47b83, 32'hbf77401b} /* (28, 26, 18) {real, imag} */,
  {32'h3c8c41c0, 32'hbf7b5302} /* (28, 26, 17) {real, imag} */,
  {32'h3f0038f6, 32'hbcc65452} /* (28, 26, 16) {real, imag} */,
  {32'h3f9da833, 32'hbeca6984} /* (28, 26, 15) {real, imag} */,
  {32'h3f2a8b39, 32'hbe67a37a} /* (28, 26, 14) {real, imag} */,
  {32'h3f84dab4, 32'h3fcf3d8b} /* (28, 26, 13) {real, imag} */,
  {32'h3e171f0d, 32'h40972812} /* (28, 26, 12) {real, imag} */,
  {32'h401a7ff6, 32'h3fd43620} /* (28, 26, 11) {real, imag} */,
  {32'hbfb15884, 32'h408e39b6} /* (28, 26, 10) {real, imag} */,
  {32'h4039ed8b, 32'h3f1d8bab} /* (28, 26, 9) {real, imag} */,
  {32'h406dfb40, 32'h3f987903} /* (28, 26, 8) {real, imag} */,
  {32'hbe940f9d, 32'hc0302897} /* (28, 26, 7) {real, imag} */,
  {32'hbffadc81, 32'hbfc5a99d} /* (28, 26, 6) {real, imag} */,
  {32'hc03b7bd0, 32'h3f28cafd} /* (28, 26, 5) {real, imag} */,
  {32'hc016d383, 32'hc043559b} /* (28, 26, 4) {real, imag} */,
  {32'hbf113567, 32'h400b1602} /* (28, 26, 3) {real, imag} */,
  {32'hc0c505f6, 32'hc065ac28} /* (28, 26, 2) {real, imag} */,
  {32'hc0872809, 32'hbdaf95a4} /* (28, 26, 1) {real, imag} */,
  {32'hc00e91e8, 32'h409b6666} /* (28, 26, 0) {real, imag} */,
  {32'hc10b524d, 32'h3f61f465} /* (28, 25, 31) {real, imag} */,
  {32'h40b1c70e, 32'hbe9990e9} /* (28, 25, 30) {real, imag} */,
  {32'hc0313c59, 32'h3fe8d68c} /* (28, 25, 29) {real, imag} */,
  {32'hbf0e68e3, 32'h40204f41} /* (28, 25, 28) {real, imag} */,
  {32'hbfbf5d6f, 32'hc09e6d43} /* (28, 25, 27) {real, imag} */,
  {32'hc0a87f67, 32'hc01df0d8} /* (28, 25, 26) {real, imag} */,
  {32'h40a2e4f3, 32'h400a6e7e} /* (28, 25, 25) {real, imag} */,
  {32'hbdbe2c17, 32'hbfec7ae2} /* (28, 25, 24) {real, imag} */,
  {32'h3fa7ce63, 32'h3f034421} /* (28, 25, 23) {real, imag} */,
  {32'hc06ce5d0, 32'hc0369534} /* (28, 25, 22) {real, imag} */,
  {32'h400bfb3c, 32'h4010a173} /* (28, 25, 21) {real, imag} */,
  {32'hbf4bccf6, 32'h3f8eea51} /* (28, 25, 20) {real, imag} */,
  {32'h3fca2df4, 32'h3d45506f} /* (28, 25, 19) {real, imag} */,
  {32'h400d307c, 32'hbfce0ddd} /* (28, 25, 18) {real, imag} */,
  {32'hbf9531ad, 32'h3f939686} /* (28, 25, 17) {real, imag} */,
  {32'h3ff9ade5, 32'h3f8e4a98} /* (28, 25, 16) {real, imag} */,
  {32'h3fbdd93d, 32'h3f626fad} /* (28, 25, 15) {real, imag} */,
  {32'hbfaa8fc9, 32'hbd3e15a9} /* (28, 25, 14) {real, imag} */,
  {32'hbede77dd, 32'h406392e0} /* (28, 25, 13) {real, imag} */,
  {32'h40068999, 32'hc007e3f5} /* (28, 25, 12) {real, imag} */,
  {32'hbed3432b, 32'h3ebbb186} /* (28, 25, 11) {real, imag} */,
  {32'hbefbcde7, 32'h3ea8b1b9} /* (28, 25, 10) {real, imag} */,
  {32'h406ea534, 32'hc0165a6d} /* (28, 25, 9) {real, imag} */,
  {32'hbed279eb, 32'h3f7ecc48} /* (28, 25, 8) {real, imag} */,
  {32'hc011806b, 32'h40268217} /* (28, 25, 7) {real, imag} */,
  {32'hc02ec76e, 32'h3fa9fb9b} /* (28, 25, 6) {real, imag} */,
  {32'hbf2c604b, 32'h40c52dcc} /* (28, 25, 5) {real, imag} */,
  {32'h400203f5, 32'hc03bd5d9} /* (28, 25, 4) {real, imag} */,
  {32'hc0179b29, 32'hc03000ad} /* (28, 25, 3) {real, imag} */,
  {32'h401228c5, 32'h4080f5ec} /* (28, 25, 2) {real, imag} */,
  {32'h3f90a002, 32'hc0a49773} /* (28, 25, 1) {real, imag} */,
  {32'hc037cb8f, 32'hc05ad442} /* (28, 25, 0) {real, imag} */,
  {32'h4132a3a2, 32'h406ef32a} /* (28, 24, 31) {real, imag} */,
  {32'hc07eff2f, 32'hc0b830a9} /* (28, 24, 30) {real, imag} */,
  {32'hbf5d449a, 32'hbf7b6921} /* (28, 24, 29) {real, imag} */,
  {32'h40901f6d, 32'hbfbfcfd5} /* (28, 24, 28) {real, imag} */,
  {32'hc00db859, 32'h40ce739c} /* (28, 24, 27) {real, imag} */,
  {32'hc0668c5a, 32'h3fab1618} /* (28, 24, 26) {real, imag} */,
  {32'h407bfadd, 32'hc0560785} /* (28, 24, 25) {real, imag} */,
  {32'hbf118345, 32'h3db97a45} /* (28, 24, 24) {real, imag} */,
  {32'h3fd5fefe, 32'h3efaaeb8} /* (28, 24, 23) {real, imag} */,
  {32'hbfde9834, 32'hbefc46e9} /* (28, 24, 22) {real, imag} */,
  {32'hbf918368, 32'hbf8c270f} /* (28, 24, 21) {real, imag} */,
  {32'hc001f06b, 32'h40747d13} /* (28, 24, 20) {real, imag} */,
  {32'hc00d94f4, 32'hbf538ab9} /* (28, 24, 19) {real, imag} */,
  {32'h4036db56, 32'h3f7a0b2c} /* (28, 24, 18) {real, imag} */,
  {32'h40088128, 32'h3e79a066} /* (28, 24, 17) {real, imag} */,
  {32'hbe84735b, 32'h3ff4517c} /* (28, 24, 16) {real, imag} */,
  {32'hbd695a67, 32'hbe10608d} /* (28, 24, 15) {real, imag} */,
  {32'hbf845fe0, 32'h3d4f1088} /* (28, 24, 14) {real, imag} */,
  {32'hbfe04118, 32'hbf60cebe} /* (28, 24, 13) {real, imag} */,
  {32'hbe1c7c19, 32'hbff19bb2} /* (28, 24, 12) {real, imag} */,
  {32'hc03d1744, 32'hc050333e} /* (28, 24, 11) {real, imag} */,
  {32'h3f9c2a37, 32'h3fad1e9d} /* (28, 24, 10) {real, imag} */,
  {32'h402a56b7, 32'hc00bf837} /* (28, 24, 9) {real, imag} */,
  {32'h4002310a, 32'hbe753c80} /* (28, 24, 8) {real, imag} */,
  {32'h40375430, 32'h403d33ad} /* (28, 24, 7) {real, imag} */,
  {32'h3ea194b5, 32'hc013ad3a} /* (28, 24, 6) {real, imag} */,
  {32'h40490168, 32'hc094a619} /* (28, 24, 5) {real, imag} */,
  {32'h4083a5cf, 32'h401cd06c} /* (28, 24, 4) {real, imag} */,
  {32'hc084bf9e, 32'hc0c966e2} /* (28, 24, 3) {real, imag} */,
  {32'hc04fdc1b, 32'hc093aa16} /* (28, 24, 2) {real, imag} */,
  {32'h40f9bfbb, 32'h40e9cc1c} /* (28, 24, 1) {real, imag} */,
  {32'h40024a59, 32'h3f877adf} /* (28, 24, 0) {real, imag} */,
  {32'hc0c542a9, 32'h3f942ea8} /* (28, 23, 31) {real, imag} */,
  {32'h400f13c1, 32'h3fa468f9} /* (28, 23, 30) {real, imag} */,
  {32'hc087a579, 32'hbff3817a} /* (28, 23, 29) {real, imag} */,
  {32'hbfa59298, 32'hc00a7a3b} /* (28, 23, 28) {real, imag} */,
  {32'hbf3f8367, 32'hbf5da665} /* (28, 23, 27) {real, imag} */,
  {32'h40b7a914, 32'h408475b6} /* (28, 23, 26) {real, imag} */,
  {32'hbe887da2, 32'hc0528a84} /* (28, 23, 25) {real, imag} */,
  {32'hc07c17be, 32'hc03aab6b} /* (28, 23, 24) {real, imag} */,
  {32'hbf8ecb38, 32'hbfc6d569} /* (28, 23, 23) {real, imag} */,
  {32'h401d0f85, 32'hbf7ec0bc} /* (28, 23, 22) {real, imag} */,
  {32'h3f09735b, 32'hbf80f578} /* (28, 23, 21) {real, imag} */,
  {32'h3f6b93c6, 32'hc02148d5} /* (28, 23, 20) {real, imag} */,
  {32'h3fc2f901, 32'hbf8748f0} /* (28, 23, 19) {real, imag} */,
  {32'hbf7fff97, 32'h3f862180} /* (28, 23, 18) {real, imag} */,
  {32'h3fa69a84, 32'hbe7fda12} /* (28, 23, 17) {real, imag} */,
  {32'h3f8eed85, 32'h3f26cba1} /* (28, 23, 16) {real, imag} */,
  {32'h3f184cf4, 32'h3fb4b63d} /* (28, 23, 15) {real, imag} */,
  {32'hbeb4a93e, 32'h3f530304} /* (28, 23, 14) {real, imag} */,
  {32'hbf2a1f84, 32'h3f223627} /* (28, 23, 13) {real, imag} */,
  {32'hbd971eb5, 32'hbed9bfc1} /* (28, 23, 12) {real, imag} */,
  {32'h40616539, 32'hbee6d828} /* (28, 23, 11) {real, imag} */,
  {32'hbf1c5928, 32'hbfbe1b9e} /* (28, 23, 10) {real, imag} */,
  {32'h3ff3c38a, 32'hbdbb7700} /* (28, 23, 9) {real, imag} */,
  {32'h401775cd, 32'h3f3b3853} /* (28, 23, 8) {real, imag} */,
  {32'h3ff1a975, 32'h3fcf9a28} /* (28, 23, 7) {real, imag} */,
  {32'hbf2fcd1f, 32'h3e9750b0} /* (28, 23, 6) {real, imag} */,
  {32'h3ffe6500, 32'h3fd562d7} /* (28, 23, 5) {real, imag} */,
  {32'hc0cac31e, 32'hc0447286} /* (28, 23, 4) {real, imag} */,
  {32'h3ed68390, 32'h3fc4b25e} /* (28, 23, 3) {real, imag} */,
  {32'h40166f44, 32'hc023ce49} /* (28, 23, 2) {real, imag} */,
  {32'h3f94f384, 32'h401fe32c} /* (28, 23, 1) {real, imag} */,
  {32'hbfdf855f, 32'h40029399} /* (28, 23, 0) {real, imag} */,
  {32'h3ea86129, 32'hbe38cfc1} /* (28, 22, 31) {real, imag} */,
  {32'h409cbc3d, 32'hbea44f25} /* (28, 22, 30) {real, imag} */,
  {32'h40327463, 32'h3fe43631} /* (28, 22, 29) {real, imag} */,
  {32'h3fd4ca0a, 32'h40243aae} /* (28, 22, 28) {real, imag} */,
  {32'h3fce53e6, 32'hbfcaffed} /* (28, 22, 27) {real, imag} */,
  {32'hbfdcf3c7, 32'hc00e56f2} /* (28, 22, 26) {real, imag} */,
  {32'hc008f060, 32'h3ed97695} /* (28, 22, 25) {real, imag} */,
  {32'h4049b0f1, 32'h404f4612} /* (28, 22, 24) {real, imag} */,
  {32'h40909e3e, 32'h401a416b} /* (28, 22, 23) {real, imag} */,
  {32'hbf963542, 32'h3d4d6542} /* (28, 22, 22) {real, imag} */,
  {32'hbfbcb373, 32'hbf073de9} /* (28, 22, 21) {real, imag} */,
  {32'hc0130e31, 32'hbfc8d618} /* (28, 22, 20) {real, imag} */,
  {32'hbe47f782, 32'hbfa482a1} /* (28, 22, 19) {real, imag} */,
  {32'hbf6e0ee6, 32'h3ff4cbc4} /* (28, 22, 18) {real, imag} */,
  {32'hc03c24fd, 32'hbe6f738d} /* (28, 22, 17) {real, imag} */,
  {32'hbf3c4ba9, 32'h3f90d99b} /* (28, 22, 16) {real, imag} */,
  {32'h3f1eb52e, 32'hbd2296a3} /* (28, 22, 15) {real, imag} */,
  {32'hbe73be23, 32'hbf96c78f} /* (28, 22, 14) {real, imag} */,
  {32'h3eb80f8e, 32'hbf5ce9e6} /* (28, 22, 13) {real, imag} */,
  {32'h3f872626, 32'hc0009178} /* (28, 22, 12) {real, imag} */,
  {32'h40269995, 32'h3fc1863e} /* (28, 22, 11) {real, imag} */,
  {32'hbed04182, 32'h3e512868} /* (28, 22, 10) {real, imag} */,
  {32'h3fc1f4fb, 32'h40b84927} /* (28, 22, 9) {real, imag} */,
  {32'h3f3b9b4c, 32'h3dd93fbe} /* (28, 22, 8) {real, imag} */,
  {32'hbfef55d0, 32'hc011a2fc} /* (28, 22, 7) {real, imag} */,
  {32'hc052101f, 32'hc02ee1d2} /* (28, 22, 6) {real, imag} */,
  {32'hbf91f6f5, 32'hbf578439} /* (28, 22, 5) {real, imag} */,
  {32'hbf0c2bb8, 32'hbe4bb2cf} /* (28, 22, 4) {real, imag} */,
  {32'h4017d97b, 32'h3f366b18} /* (28, 22, 3) {real, imag} */,
  {32'h3fda92f9, 32'hc08d9ae1} /* (28, 22, 2) {real, imag} */,
  {32'hc0005cad, 32'h400627b2} /* (28, 22, 1) {real, imag} */,
  {32'hc054d540, 32'h3e371ff7} /* (28, 22, 0) {real, imag} */,
  {32'h40c4f597, 32'h3ee0def7} /* (28, 21, 31) {real, imag} */,
  {32'h3f2a8bae, 32'h4090e89b} /* (28, 21, 30) {real, imag} */,
  {32'h407219de, 32'hbed2fdb1} /* (28, 21, 29) {real, imag} */,
  {32'hbde7de12, 32'hbf3621ee} /* (28, 21, 28) {real, imag} */,
  {32'hc08dadab, 32'h3fc8faf0} /* (28, 21, 27) {real, imag} */,
  {32'hbf35661e, 32'h4006d69f} /* (28, 21, 26) {real, imag} */,
  {32'hbf6db495, 32'h3f33a646} /* (28, 21, 25) {real, imag} */,
  {32'hbfc0710c, 32'hbf72b120} /* (28, 21, 24) {real, imag} */,
  {32'hbfa176fe, 32'hbfb0bf3e} /* (28, 21, 23) {real, imag} */,
  {32'hbf3438c4, 32'hc0605f69} /* (28, 21, 22) {real, imag} */,
  {32'h3fbac362, 32'h3ec6f49a} /* (28, 21, 21) {real, imag} */,
  {32'h3cba5a73, 32'hbd0167f2} /* (28, 21, 20) {real, imag} */,
  {32'hc021da80, 32'hbf246f60} /* (28, 21, 19) {real, imag} */,
  {32'hc00a2132, 32'h3fb66002} /* (28, 21, 18) {real, imag} */,
  {32'h3f2627b6, 32'hc01232d7} /* (28, 21, 17) {real, imag} */,
  {32'h3f8cec99, 32'h3f99b96d} /* (28, 21, 16) {real, imag} */,
  {32'hbfc589fc, 32'h3f3ecad1} /* (28, 21, 15) {real, imag} */,
  {32'h3f74bc0c, 32'hbfc3120b} /* (28, 21, 14) {real, imag} */,
  {32'hc04fcb4b, 32'h3ff1e093} /* (28, 21, 13) {real, imag} */,
  {32'hc037db67, 32'hc08292dd} /* (28, 21, 12) {real, imag} */,
  {32'hbfe79f49, 32'h3f2e9dae} /* (28, 21, 11) {real, imag} */,
  {32'h40466326, 32'h3f41948e} /* (28, 21, 10) {real, imag} */,
  {32'hc00263a9, 32'hbf942af2} /* (28, 21, 9) {real, imag} */,
  {32'h3edb81f1, 32'hc027934f} /* (28, 21, 8) {real, imag} */,
  {32'hbea05ad5, 32'h3ff3b3f2} /* (28, 21, 7) {real, imag} */,
  {32'h40077799, 32'h3f744a58} /* (28, 21, 6) {real, imag} */,
  {32'h3e497105, 32'h3f7572ce} /* (28, 21, 5) {real, imag} */,
  {32'h3fdc3e72, 32'h3e560e89} /* (28, 21, 4) {real, imag} */,
  {32'hbfa6b8fc, 32'hbfcadd48} /* (28, 21, 3) {real, imag} */,
  {32'hc0861605, 32'h3fbec722} /* (28, 21, 2) {real, imag} */,
  {32'h40240363, 32'h3f850734} /* (28, 21, 1) {real, imag} */,
  {32'h3fe3816e, 32'h3f50b365} /* (28, 21, 0) {real, imag} */,
  {32'hbee8cee5, 32'h3f0ae55e} /* (28, 20, 31) {real, imag} */,
  {32'h3fb774e4, 32'h401b53b4} /* (28, 20, 30) {real, imag} */,
  {32'hbf90858b, 32'h3f8ea72a} /* (28, 20, 29) {real, imag} */,
  {32'h3fdf9347, 32'hbf946c9a} /* (28, 20, 28) {real, imag} */,
  {32'hbf852eeb, 32'hbd06574a} /* (28, 20, 27) {real, imag} */,
  {32'hbc3e84f3, 32'hc002bc8d} /* (28, 20, 26) {real, imag} */,
  {32'hbffe9a14, 32'hc02ce580} /* (28, 20, 25) {real, imag} */,
  {32'hc00fffcc, 32'h4025d88e} /* (28, 20, 24) {real, imag} */,
  {32'hc088eacb, 32'hbd97ce63} /* (28, 20, 23) {real, imag} */,
  {32'hbfbcf0f3, 32'h3f2330dd} /* (28, 20, 22) {real, imag} */,
  {32'hbf99036f, 32'h401aa869} /* (28, 20, 21) {real, imag} */,
  {32'h3fbd91ce, 32'h3f6e707b} /* (28, 20, 20) {real, imag} */,
  {32'hc058fdfb, 32'hbeee7a83} /* (28, 20, 19) {real, imag} */,
  {32'h3e9b48bb, 32'hbf98a939} /* (28, 20, 18) {real, imag} */,
  {32'h3f55c58d, 32'hbf309354} /* (28, 20, 17) {real, imag} */,
  {32'hbe964693, 32'hbeb3a858} /* (28, 20, 16) {real, imag} */,
  {32'h3eef6f5d, 32'hbe6644e1} /* (28, 20, 15) {real, imag} */,
  {32'h40626763, 32'h3fef22a7} /* (28, 20, 14) {real, imag} */,
  {32'hbe78b5c1, 32'hbf934bfd} /* (28, 20, 13) {real, imag} */,
  {32'hbf552a95, 32'h40302acb} /* (28, 20, 12) {real, imag} */,
  {32'h3bbadd0d, 32'hc01a1c67} /* (28, 20, 11) {real, imag} */,
  {32'h3f586bce, 32'hc078b071} /* (28, 20, 10) {real, imag} */,
  {32'hbfbcc756, 32'hbfdde237} /* (28, 20, 9) {real, imag} */,
  {32'hbf78c178, 32'hbe8ca19c} /* (28, 20, 8) {real, imag} */,
  {32'h3e7b1165, 32'hbfd58dc4} /* (28, 20, 7) {real, imag} */,
  {32'h40779d32, 32'h4010010f} /* (28, 20, 6) {real, imag} */,
  {32'h3fa5ec41, 32'h404a4e62} /* (28, 20, 5) {real, imag} */,
  {32'h3f7c320e, 32'hbedc4408} /* (28, 20, 4) {real, imag} */,
  {32'h3f42e556, 32'hbf82ff4a} /* (28, 20, 3) {real, imag} */,
  {32'h3ef65f3d, 32'hbf86f31e} /* (28, 20, 2) {real, imag} */,
  {32'hbffc1300, 32'h402dc558} /* (28, 20, 1) {real, imag} */,
  {32'hbfafaf59, 32'h3f5bf710} /* (28, 20, 0) {real, imag} */,
  {32'hbf0e1e0f, 32'hc050aff7} /* (28, 19, 31) {real, imag} */,
  {32'h3fb96083, 32'hbfc575ea} /* (28, 19, 30) {real, imag} */,
  {32'hbf1ff6c6, 32'hbf80295a} /* (28, 19, 29) {real, imag} */,
  {32'hbf62b581, 32'hbfaed179} /* (28, 19, 28) {real, imag} */,
  {32'h3cadb9ef, 32'h40055e28} /* (28, 19, 27) {real, imag} */,
  {32'h3f028175, 32'hc013c14d} /* (28, 19, 26) {real, imag} */,
  {32'h3d8b5bc7, 32'hbfc0aa81} /* (28, 19, 25) {real, imag} */,
  {32'h3f0f6814, 32'h4084fc28} /* (28, 19, 24) {real, imag} */,
  {32'h3f7a5be0, 32'hbfa86078} /* (28, 19, 23) {real, imag} */,
  {32'h40218688, 32'h3fbdd1bb} /* (28, 19, 22) {real, imag} */,
  {32'hbe9f51ec, 32'hbfe79158} /* (28, 19, 21) {real, imag} */,
  {32'hbf064ecb, 32'h3ee8d718} /* (28, 19, 20) {real, imag} */,
  {32'hc030a9ad, 32'h3f8f6d84} /* (28, 19, 19) {real, imag} */,
  {32'hbf9b55bb, 32'hbf9daa51} /* (28, 19, 18) {real, imag} */,
  {32'hbe772da3, 32'h3e353280} /* (28, 19, 17) {real, imag} */,
  {32'hbf27cf22, 32'hbdf7ec96} /* (28, 19, 16) {real, imag} */,
  {32'h3f9c8e31, 32'h3f288f64} /* (28, 19, 15) {real, imag} */,
  {32'hbfe522f8, 32'h3f5e7995} /* (28, 19, 14) {real, imag} */,
  {32'h4042099e, 32'hbe289413} /* (28, 19, 13) {real, imag} */,
  {32'h3fb17dbc, 32'hc018ef63} /* (28, 19, 12) {real, imag} */,
  {32'h3ee85fa3, 32'h3f3ec0ee} /* (28, 19, 11) {real, imag} */,
  {32'hbee0fcef, 32'hbedf8e08} /* (28, 19, 10) {real, imag} */,
  {32'h3fde985b, 32'h3f9cd431} /* (28, 19, 9) {real, imag} */,
  {32'hbfc082c6, 32'hbf1ab088} /* (28, 19, 8) {real, imag} */,
  {32'hbfb1c963, 32'hc0068f93} /* (28, 19, 7) {real, imag} */,
  {32'h401fb089, 32'hbf1e214c} /* (28, 19, 6) {real, imag} */,
  {32'h40141f80, 32'h3da45921} /* (28, 19, 5) {real, imag} */,
  {32'h3f78986a, 32'hc015b7f5} /* (28, 19, 4) {real, imag} */,
  {32'hbf1ecc27, 32'hbfc87f04} /* (28, 19, 3) {real, imag} */,
  {32'hbf1d4bd3, 32'h4016b9e6} /* (28, 19, 2) {real, imag} */,
  {32'hbf65a805, 32'hbff3f9d9} /* (28, 19, 1) {real, imag} */,
  {32'hc0425d6b, 32'h3fe00a38} /* (28, 19, 0) {real, imag} */,
  {32'h40120b7d, 32'hbf98c784} /* (28, 18, 31) {real, imag} */,
  {32'hbfcc131c, 32'h403b753b} /* (28, 18, 30) {real, imag} */,
  {32'hbf39dee9, 32'hbec0741f} /* (28, 18, 29) {real, imag} */,
  {32'h4004934f, 32'h3ec8a8a7} /* (28, 18, 28) {real, imag} */,
  {32'hbf6b610f, 32'h3e07c57b} /* (28, 18, 27) {real, imag} */,
  {32'h3f346962, 32'hbfb2f3de} /* (28, 18, 26) {real, imag} */,
  {32'hbfa0eee2, 32'h3fbebaf4} /* (28, 18, 25) {real, imag} */,
  {32'h3f3ad753, 32'hbff10793} /* (28, 18, 24) {real, imag} */,
  {32'hbedd9ac7, 32'h3fd1f8a1} /* (28, 18, 23) {real, imag} */,
  {32'h3eb7f41c, 32'h3cefc3b4} /* (28, 18, 22) {real, imag} */,
  {32'h3f8bd469, 32'h3fbb5965} /* (28, 18, 21) {real, imag} */,
  {32'hbd977b99, 32'hbf9d261e} /* (28, 18, 20) {real, imag} */,
  {32'hbe66f262, 32'hbe86946a} /* (28, 18, 19) {real, imag} */,
  {32'hbf866575, 32'hbfad2587} /* (28, 18, 18) {real, imag} */,
  {32'hbe022f65, 32'h3f97ca49} /* (28, 18, 17) {real, imag} */,
  {32'hbe5e5c07, 32'hbf9c8951} /* (28, 18, 16) {real, imag} */,
  {32'h3f6c66c8, 32'hbf4480bf} /* (28, 18, 15) {real, imag} */,
  {32'hbed61d58, 32'hc01dd523} /* (28, 18, 14) {real, imag} */,
  {32'h3f1d784c, 32'h404af479} /* (28, 18, 13) {real, imag} */,
  {32'hc01cc6df, 32'h3ee0d517} /* (28, 18, 12) {real, imag} */,
  {32'h3e568f5f, 32'h3fa77a38} /* (28, 18, 11) {real, imag} */,
  {32'hbdbb1c14, 32'h40111c92} /* (28, 18, 10) {real, imag} */,
  {32'hbe109740, 32'hbf85c466} /* (28, 18, 9) {real, imag} */,
  {32'h4006a048, 32'h3fc98b95} /* (28, 18, 8) {real, imag} */,
  {32'h3fd8eca4, 32'hbfcd1dbc} /* (28, 18, 7) {real, imag} */,
  {32'h3f936fc2, 32'hbf4bcd87} /* (28, 18, 6) {real, imag} */,
  {32'hbf429b73, 32'hbf99c2f2} /* (28, 18, 5) {real, imag} */,
  {32'h3f3f8812, 32'h3fb52800} /* (28, 18, 4) {real, imag} */,
  {32'h3df86fb8, 32'h3efed998} /* (28, 18, 3) {real, imag} */,
  {32'h3ea12fab, 32'hbedc24e4} /* (28, 18, 2) {real, imag} */,
  {32'h406aaa4d, 32'h3cc1166d} /* (28, 18, 1) {real, imag} */,
  {32'h3f1919b1, 32'hbf808e9d} /* (28, 18, 0) {real, imag} */,
  {32'hc0280c4c, 32'hbf7324ec} /* (28, 17, 31) {real, imag} */,
  {32'h3fa858cf, 32'hbf1f03ce} /* (28, 17, 30) {real, imag} */,
  {32'hbfbe30fe, 32'hbf9ebfcb} /* (28, 17, 29) {real, imag} */,
  {32'h3eb495c8, 32'hbfeaef46} /* (28, 17, 28) {real, imag} */,
  {32'h401137b3, 32'h3f613839} /* (28, 17, 27) {real, imag} */,
  {32'h3fb8d515, 32'hbe82569d} /* (28, 17, 26) {real, imag} */,
  {32'h3c9643d8, 32'h3fe3e0e6} /* (28, 17, 25) {real, imag} */,
  {32'h3ea2a18d, 32'h3efc9787} /* (28, 17, 24) {real, imag} */,
  {32'h3f151b3b, 32'h3fc36ca2} /* (28, 17, 23) {real, imag} */,
  {32'h3ee306df, 32'hbf27ed57} /* (28, 17, 22) {real, imag} */,
  {32'hc0368fb0, 32'hbf6474a6} /* (28, 17, 21) {real, imag} */,
  {32'hbf903a61, 32'hbfb553b8} /* (28, 17, 20) {real, imag} */,
  {32'hbd5395de, 32'h3e1762d0} /* (28, 17, 19) {real, imag} */,
  {32'h3f961a3c, 32'hbdb313d7} /* (28, 17, 18) {real, imag} */,
  {32'hbea641d3, 32'hbe640677} /* (28, 17, 17) {real, imag} */,
  {32'h3e0acbf8, 32'hbf65d9f9} /* (28, 17, 16) {real, imag} */,
  {32'h3f409de2, 32'h3f167e35} /* (28, 17, 15) {real, imag} */,
  {32'hbe6842a6, 32'hbf457f54} /* (28, 17, 14) {real, imag} */,
  {32'hbf73d121, 32'hbf3d37b4} /* (28, 17, 13) {real, imag} */,
  {32'h3f87d565, 32'h3eb2f728} /* (28, 17, 12) {real, imag} */,
  {32'hc04aa4cd, 32'hbebac52c} /* (28, 17, 11) {real, imag} */,
  {32'h401e2b6b, 32'h3f894a5b} /* (28, 17, 10) {real, imag} */,
  {32'h402cf4dd, 32'h3fb6b210} /* (28, 17, 9) {real, imag} */,
  {32'h40055808, 32'h405cbc06} /* (28, 17, 8) {real, imag} */,
  {32'h40135186, 32'hbee14e64} /* (28, 17, 7) {real, imag} */,
  {32'hbed24904, 32'hbfe19913} /* (28, 17, 6) {real, imag} */,
  {32'hbdbafa89, 32'h3e7414e9} /* (28, 17, 5) {real, imag} */,
  {32'hbfd98c37, 32'h3fb5c1c8} /* (28, 17, 4) {real, imag} */,
  {32'hbffec727, 32'h3f46a8ca} /* (28, 17, 3) {real, imag} */,
  {32'hbbe311d7, 32'hbfdaf243} /* (28, 17, 2) {real, imag} */,
  {32'hbf87b66a, 32'hbefe4a66} /* (28, 17, 1) {real, imag} */,
  {32'hbf3a5c64, 32'h3e20f418} /* (28, 17, 0) {real, imag} */,
  {32'h3f80c595, 32'hbdcc2d01} /* (28, 16, 31) {real, imag} */,
  {32'h3e42b288, 32'hbf7ec8a6} /* (28, 16, 30) {real, imag} */,
  {32'hbfbf0126, 32'h3ddf52d8} /* (28, 16, 29) {real, imag} */,
  {32'h3ec8e32e, 32'h3ff0ef53} /* (28, 16, 28) {real, imag} */,
  {32'hbf9d87b4, 32'hbf84030d} /* (28, 16, 27) {real, imag} */,
  {32'h3f56260f, 32'h3fd88531} /* (28, 16, 26) {real, imag} */,
  {32'h3f7db075, 32'h3efd1ba0} /* (28, 16, 25) {real, imag} */,
  {32'hbecb4894, 32'h3f22b414} /* (28, 16, 24) {real, imag} */,
  {32'hbf398267, 32'hbee7af6c} /* (28, 16, 23) {real, imag} */,
  {32'hbfa080e5, 32'hbd167db6} /* (28, 16, 22) {real, imag} */,
  {32'hbea221ad, 32'hbfb4d365} /* (28, 16, 21) {real, imag} */,
  {32'hbf88156e, 32'h3f0def1b} /* (28, 16, 20) {real, imag} */,
  {32'h4081afce, 32'hbd3b0c5a} /* (28, 16, 19) {real, imag} */,
  {32'hbeed59e9, 32'hbf80281e} /* (28, 16, 18) {real, imag} */,
  {32'hbf7ede65, 32'hbee7d674} /* (28, 16, 17) {real, imag} */,
  {32'h3fe78f22, 32'h3e1ab163} /* (28, 16, 16) {real, imag} */,
  {32'hbec9877e, 32'hbf0025e6} /* (28, 16, 15) {real, imag} */,
  {32'hbf725fc5, 32'hbf20023e} /* (28, 16, 14) {real, imag} */,
  {32'hbf4c0294, 32'hbfd08ae6} /* (28, 16, 13) {real, imag} */,
  {32'h3ef5c42d, 32'h3f0f674e} /* (28, 16, 12) {real, imag} */,
  {32'h3f8ce44b, 32'hbed93c86} /* (28, 16, 11) {real, imag} */,
  {32'hbf396cf8, 32'hbf0e0552} /* (28, 16, 10) {real, imag} */,
  {32'hbfdab5c0, 32'hbf46d0d0} /* (28, 16, 9) {real, imag} */,
  {32'hbed18232, 32'hbfe10177} /* (28, 16, 8) {real, imag} */,
  {32'hbf1b103a, 32'hbf7b277d} /* (28, 16, 7) {real, imag} */,
  {32'h3e9da2f0, 32'hbf97e984} /* (28, 16, 6) {real, imag} */,
  {32'hc01ec4fc, 32'h3e0bfe47} /* (28, 16, 5) {real, imag} */,
  {32'hbe801ac5, 32'h3fcb0508} /* (28, 16, 4) {real, imag} */,
  {32'h3f2903c2, 32'hbf9093d9} /* (28, 16, 3) {real, imag} */,
  {32'h3f28950c, 32'h3f570baa} /* (28, 16, 2) {real, imag} */,
  {32'h3f8bdc65, 32'hbe5370ba} /* (28, 16, 1) {real, imag} */,
  {32'h3eed3bdf, 32'hc00b8bd5} /* (28, 16, 0) {real, imag} */,
  {32'h3e5a6c8d, 32'hbf060890} /* (28, 15, 31) {real, imag} */,
  {32'h3ee56730, 32'hbeffec71} /* (28, 15, 30) {real, imag} */,
  {32'h3d848438, 32'hc039de8b} /* (28, 15, 29) {real, imag} */,
  {32'h3f63d961, 32'h3f19b2ff} /* (28, 15, 28) {real, imag} */,
  {32'h3fc3441b, 32'hbe2c2713} /* (28, 15, 27) {real, imag} */,
  {32'h3f327ca8, 32'h4024a8df} /* (28, 15, 26) {real, imag} */,
  {32'hbec7a204, 32'h3f89ccdb} /* (28, 15, 25) {real, imag} */,
  {32'hbf3065bf, 32'hc0016621} /* (28, 15, 24) {real, imag} */,
  {32'h3e5f8b0b, 32'hbf688ebb} /* (28, 15, 23) {real, imag} */,
  {32'hbe418edc, 32'hbe99a965} /* (28, 15, 22) {real, imag} */,
  {32'hbf8012fb, 32'hbc47e3f0} /* (28, 15, 21) {real, imag} */,
  {32'h403a495f, 32'h3ecd2344} /* (28, 15, 20) {real, imag} */,
  {32'hbf9b01ae, 32'h4036f703} /* (28, 15, 19) {real, imag} */,
  {32'h3f5526f6, 32'h3f821958} /* (28, 15, 18) {real, imag} */,
  {32'h3e2a55a6, 32'hbfff8c82} /* (28, 15, 17) {real, imag} */,
  {32'hbf122511, 32'hbe048ea5} /* (28, 15, 16) {real, imag} */,
  {32'h3f8b5662, 32'hbf0a91bf} /* (28, 15, 15) {real, imag} */,
  {32'h4001c6a2, 32'h3e763e3b} /* (28, 15, 14) {real, imag} */,
  {32'h3f91208b, 32'h3f22029b} /* (28, 15, 13) {real, imag} */,
  {32'hbfc733b5, 32'hc0115872} /* (28, 15, 12) {real, imag} */,
  {32'h404229c2, 32'hbfa0d16e} /* (28, 15, 11) {real, imag} */,
  {32'hbf0e2b04, 32'h3d0994f6} /* (28, 15, 10) {real, imag} */,
  {32'hbf3f8b0a, 32'hbf3f2702} /* (28, 15, 9) {real, imag} */,
  {32'hbf7745af, 32'hbff7a638} /* (28, 15, 8) {real, imag} */,
  {32'hbf196f37, 32'h3ffc4fae} /* (28, 15, 7) {real, imag} */,
  {32'hbf82e25e, 32'h3f10b3a4} /* (28, 15, 6) {real, imag} */,
  {32'hbf0a152e, 32'h3fad6811} /* (28, 15, 5) {real, imag} */,
  {32'h3ed3c0ac, 32'h3f3dac7a} /* (28, 15, 4) {real, imag} */,
  {32'hbf3ecba7, 32'h400aa8f8} /* (28, 15, 3) {real, imag} */,
  {32'h3e59ecb7, 32'h3e6440db} /* (28, 15, 2) {real, imag} */,
  {32'h3fc3e42c, 32'hbfc2cb7c} /* (28, 15, 1) {real, imag} */,
  {32'hbf08f434, 32'h3fba38b5} /* (28, 15, 0) {real, imag} */,
  {32'hc03c3619, 32'h3e7b98e0} /* (28, 14, 31) {real, imag} */,
  {32'h3f56b248, 32'h3f09a328} /* (28, 14, 30) {real, imag} */,
  {32'h3eb087c5, 32'h3f4a781b} /* (28, 14, 29) {real, imag} */,
  {32'h3fb08d51, 32'hbed99a26} /* (28, 14, 28) {real, imag} */,
  {32'hbf0ff506, 32'h3e44634e} /* (28, 14, 27) {real, imag} */,
  {32'h4049f721, 32'hc029a84b} /* (28, 14, 26) {real, imag} */,
  {32'hc0086ae4, 32'hbca2f146} /* (28, 14, 25) {real, imag} */,
  {32'hbfd0d80c, 32'h3fb14802} /* (28, 14, 24) {real, imag} */,
  {32'h3f605405, 32'h3f1c6036} /* (28, 14, 23) {real, imag} */,
  {32'h3f592577, 32'h3fe4b1a7} /* (28, 14, 22) {real, imag} */,
  {32'hbf6df43c, 32'h3f4a3cee} /* (28, 14, 21) {real, imag} */,
  {32'h3fa61d56, 32'h3f7ec496} /* (28, 14, 20) {real, imag} */,
  {32'h3fae4ff7, 32'hbf3577d2} /* (28, 14, 19) {real, imag} */,
  {32'hbf592ffd, 32'h3fc0e1fe} /* (28, 14, 18) {real, imag} */,
  {32'hbefd2816, 32'h3f967e08} /* (28, 14, 17) {real, imag} */,
  {32'hbef04334, 32'h3f2a949e} /* (28, 14, 16) {real, imag} */,
  {32'hbfe3c94a, 32'hbfbf7c80} /* (28, 14, 15) {real, imag} */,
  {32'h3eb626c5, 32'h3e86404b} /* (28, 14, 14) {real, imag} */,
  {32'hbf4c7723, 32'hba48f653} /* (28, 14, 13) {real, imag} */,
  {32'hbedcaa5c, 32'h3b0eee0e} /* (28, 14, 12) {real, imag} */,
  {32'h3fad8327, 32'hbefa426b} /* (28, 14, 11) {real, imag} */,
  {32'hc0860799, 32'hc00489ba} /* (28, 14, 10) {real, imag} */,
  {32'h3e49b43e, 32'hbfa1dd08} /* (28, 14, 9) {real, imag} */,
  {32'hc00bd9ee, 32'hbfb58b4f} /* (28, 14, 8) {real, imag} */,
  {32'h3fa76325, 32'h3ef3c4a4} /* (28, 14, 7) {real, imag} */,
  {32'h4004e3e8, 32'hbf86bcbb} /* (28, 14, 6) {real, imag} */,
  {32'h3fca4511, 32'hbe05e599} /* (28, 14, 5) {real, imag} */,
  {32'h3fb010b0, 32'h3fb3d69d} /* (28, 14, 4) {real, imag} */,
  {32'h3e68014d, 32'hbf598c1b} /* (28, 14, 3) {real, imag} */,
  {32'h3fa3cd07, 32'hc016d243} /* (28, 14, 2) {real, imag} */,
  {32'h3fca307f, 32'h3fbdda2e} /* (28, 14, 1) {real, imag} */,
  {32'hc005dcf7, 32'h3fb4b309} /* (28, 14, 0) {real, imag} */,
  {32'h3f688ae3, 32'h3e3dc453} /* (28, 13, 31) {real, imag} */,
  {32'hbfaccff6, 32'h4000a4f2} /* (28, 13, 30) {real, imag} */,
  {32'h400f4878, 32'h3df6281b} /* (28, 13, 29) {real, imag} */,
  {32'hbea29449, 32'hbdda5533} /* (28, 13, 28) {real, imag} */,
  {32'h3f8141f3, 32'h3f1408c6} /* (28, 13, 27) {real, imag} */,
  {32'h3e1c28c6, 32'hbeefc298} /* (28, 13, 26) {real, imag} */,
  {32'hbdab9ef6, 32'h400014be} /* (28, 13, 25) {real, imag} */,
  {32'h3f73c722, 32'h3ef1a336} /* (28, 13, 24) {real, imag} */,
  {32'hbfa7f3cf, 32'hbea60e71} /* (28, 13, 23) {real, imag} */,
  {32'hc062d755, 32'h3e1e31f1} /* (28, 13, 22) {real, imag} */,
  {32'hc04d0ace, 32'hbfa85cf0} /* (28, 13, 21) {real, imag} */,
  {32'h3f27f2e7, 32'hbfacb6c2} /* (28, 13, 20) {real, imag} */,
  {32'hbfe6bcb7, 32'h3ff972b2} /* (28, 13, 19) {real, imag} */,
  {32'hbd266330, 32'h4035c5fe} /* (28, 13, 18) {real, imag} */,
  {32'h3f4429b5, 32'h40079742} /* (28, 13, 17) {real, imag} */,
  {32'h3fb101cf, 32'hbfa4a6c9} /* (28, 13, 16) {real, imag} */,
  {32'h3cac67e2, 32'h3fc7db63} /* (28, 13, 15) {real, imag} */,
  {32'hbf102b24, 32'hbf152220} /* (28, 13, 14) {real, imag} */,
  {32'h3f3f18fb, 32'hbe6f160f} /* (28, 13, 13) {real, imag} */,
  {32'hbf5dde6c, 32'h3f941aa6} /* (28, 13, 12) {real, imag} */,
  {32'hbf88ba7f, 32'h3f088d20} /* (28, 13, 11) {real, imag} */,
  {32'h40131133, 32'h402efde6} /* (28, 13, 10) {real, imag} */,
  {32'hbfad25c9, 32'hbe5592be} /* (28, 13, 9) {real, imag} */,
  {32'h40294e46, 32'hbfb07ec8} /* (28, 13, 8) {real, imag} */,
  {32'h3ee2c745, 32'h3fc1ff86} /* (28, 13, 7) {real, imag} */,
  {32'h3fffb60f, 32'hbe7dc6a3} /* (28, 13, 6) {real, imag} */,
  {32'hbe67c916, 32'h4029b02b} /* (28, 13, 5) {real, imag} */,
  {32'hc00c3bdd, 32'hc0302fe4} /* (28, 13, 4) {real, imag} */,
  {32'h3fc24f4e, 32'h3fa47113} /* (28, 13, 3) {real, imag} */,
  {32'hc00da3dc, 32'hbf36a67a} /* (28, 13, 2) {real, imag} */,
  {32'hbef4a09f, 32'hbfca3657} /* (28, 13, 1) {real, imag} */,
  {32'h40045fad, 32'hbe991342} /* (28, 13, 0) {real, imag} */,
  {32'hbfa8047c, 32'h3ef544d3} /* (28, 12, 31) {real, imag} */,
  {32'h40bc88b1, 32'hbe268ad9} /* (28, 12, 30) {real, imag} */,
  {32'hbe27ba99, 32'hbff2296a} /* (28, 12, 29) {real, imag} */,
  {32'hbf755ca4, 32'hbf000153} /* (28, 12, 28) {real, imag} */,
  {32'hbfbbe502, 32'hc0897102} /* (28, 12, 27) {real, imag} */,
  {32'h3f7f1770, 32'hbf345bd5} /* (28, 12, 26) {real, imag} */,
  {32'h3f9e3dd2, 32'h3fee0a6d} /* (28, 12, 25) {real, imag} */,
  {32'hc04e99ef, 32'hbeed9636} /* (28, 12, 24) {real, imag} */,
  {32'h3e8816dc, 32'h3fdefc0e} /* (28, 12, 23) {real, imag} */,
  {32'h3e3f72ee, 32'h4062eba9} /* (28, 12, 22) {real, imag} */,
  {32'hbf8dd9c4, 32'hc0870963} /* (28, 12, 21) {real, imag} */,
  {32'hbf3aabaa, 32'h3fda90ef} /* (28, 12, 20) {real, imag} */,
  {32'h3efeeb6c, 32'h3f9adfa3} /* (28, 12, 19) {real, imag} */,
  {32'hbf82f9b1, 32'h3fe4f536} /* (28, 12, 18) {real, imag} */,
  {32'hbf821d3a, 32'hc0069c22} /* (28, 12, 17) {real, imag} */,
  {32'h3e37ef9b, 32'hbf34faff} /* (28, 12, 16) {real, imag} */,
  {32'hbf67c15b, 32'h3fc19cb2} /* (28, 12, 15) {real, imag} */,
  {32'hbecf1ed3, 32'h3fae31a9} /* (28, 12, 14) {real, imag} */,
  {32'hc013395a, 32'hbd89b6b4} /* (28, 12, 13) {real, imag} */,
  {32'hbe6fa3bd, 32'hbfca008a} /* (28, 12, 12) {real, imag} */,
  {32'h3f67886f, 32'h3f1a4157} /* (28, 12, 11) {real, imag} */,
  {32'h3edee188, 32'h3f05d50b} /* (28, 12, 10) {real, imag} */,
  {32'hbe28b58f, 32'hc00019a5} /* (28, 12, 9) {real, imag} */,
  {32'h400f024b, 32'h3ff883ce} /* (28, 12, 8) {real, imag} */,
  {32'h3f739bd8, 32'hbf188815} /* (28, 12, 7) {real, imag} */,
  {32'h3eab286a, 32'hbf2544bb} /* (28, 12, 6) {real, imag} */,
  {32'h3ef08dde, 32'h4019db4d} /* (28, 12, 5) {real, imag} */,
  {32'hbea3befb, 32'hbfa656d9} /* (28, 12, 4) {real, imag} */,
  {32'hc0042199, 32'hbf5184f1} /* (28, 12, 3) {real, imag} */,
  {32'h3d949bd2, 32'hbbee8f8e} /* (28, 12, 2) {real, imag} */,
  {32'h3fdcc14b, 32'hbf74f1d0} /* (28, 12, 1) {real, imag} */,
  {32'h3fb6509d, 32'h3f696db0} /* (28, 12, 0) {real, imag} */,
  {32'h3e8e9075, 32'h402e9585} /* (28, 11, 31) {real, imag} */,
  {32'h409380a9, 32'hbfb45ca5} /* (28, 11, 30) {real, imag} */,
  {32'h3f9d6471, 32'h3ff2dbb8} /* (28, 11, 29) {real, imag} */,
  {32'h3eaa5dea, 32'h3edd1316} /* (28, 11, 28) {real, imag} */,
  {32'hbf66046e, 32'hc053d3b8} /* (28, 11, 27) {real, imag} */,
  {32'h400d1ccf, 32'hbf8bb339} /* (28, 11, 26) {real, imag} */,
  {32'hbf6abe51, 32'h4014c4ec} /* (28, 11, 25) {real, imag} */,
  {32'h3f954a1a, 32'h3f63330c} /* (28, 11, 24) {real, imag} */,
  {32'h3fd9ee66, 32'hbf8666b2} /* (28, 11, 23) {real, imag} */,
  {32'hbfc42222, 32'h4008b443} /* (28, 11, 22) {real, imag} */,
  {32'h3f460a39, 32'hbf961da7} /* (28, 11, 21) {real, imag} */,
  {32'h3f361cfc, 32'h3d976a36} /* (28, 11, 20) {real, imag} */,
  {32'hbfadf3d0, 32'hbedcdb93} /* (28, 11, 19) {real, imag} */,
  {32'h3fa259a1, 32'h3db93eac} /* (28, 11, 18) {real, imag} */,
  {32'hbf753314, 32'h3f3db492} /* (28, 11, 17) {real, imag} */,
  {32'h4002c145, 32'h3f8097bc} /* (28, 11, 16) {real, imag} */,
  {32'h3f46a2fc, 32'h3ebaa2ea} /* (28, 11, 15) {real, imag} */,
  {32'hbf1eaf87, 32'h3e5fe6a5} /* (28, 11, 14) {real, imag} */,
  {32'hbdc93c18, 32'hc004bc1d} /* (28, 11, 13) {real, imag} */,
  {32'h3f889bbf, 32'hbf68d333} /* (28, 11, 12) {real, imag} */,
  {32'h3f410f8f, 32'h3fccda4c} /* (28, 11, 11) {real, imag} */,
  {32'hc02e8fb9, 32'h3fe48fbe} /* (28, 11, 10) {real, imag} */,
  {32'hbf6393ad, 32'hbe6df008} /* (28, 11, 9) {real, imag} */,
  {32'hbfc44395, 32'h3fda59d4} /* (28, 11, 8) {real, imag} */,
  {32'hbfaae917, 32'hbfeacbf7} /* (28, 11, 7) {real, imag} */,
  {32'h3fd26cdd, 32'h3ee3638e} /* (28, 11, 6) {real, imag} */,
  {32'h3fa39311, 32'hbfde37c0} /* (28, 11, 5) {real, imag} */,
  {32'h3eb89dd4, 32'h3fae0401} /* (28, 11, 4) {real, imag} */,
  {32'hc04f1c07, 32'hc036eb5b} /* (28, 11, 3) {real, imag} */,
  {32'h40c0dc4f, 32'hbf9f0f44} /* (28, 11, 2) {real, imag} */,
  {32'hc0051d94, 32'h3f35ab0a} /* (28, 11, 1) {real, imag} */,
  {32'hc07c47e9, 32'h3ff5a1a6} /* (28, 11, 0) {real, imag} */,
  {32'hbf99d3ba, 32'hbffec947} /* (28, 10, 31) {real, imag} */,
  {32'hc0091ea6, 32'h4093b8e5} /* (28, 10, 30) {real, imag} */,
  {32'hc034a9ae, 32'hc0302868} /* (28, 10, 29) {real, imag} */,
  {32'hc0151e2f, 32'hbfac7fd1} /* (28, 10, 28) {real, imag} */,
  {32'hbea40b57, 32'hbec7b3d3} /* (28, 10, 27) {real, imag} */,
  {32'hbf293d1a, 32'hbf000ad2} /* (28, 10, 26) {real, imag} */,
  {32'h3f87ae71, 32'hbfa1859e} /* (28, 10, 25) {real, imag} */,
  {32'hbf615943, 32'hbf1e4c1e} /* (28, 10, 24) {real, imag} */,
  {32'h3fe45b1b, 32'hc0060b1c} /* (28, 10, 23) {real, imag} */,
  {32'hbf7a2359, 32'h3d5f644c} /* (28, 10, 22) {real, imag} */,
  {32'hbf7be1d6, 32'h3f10d108} /* (28, 10, 21) {real, imag} */,
  {32'h3e43960d, 32'hc00e7aaf} /* (28, 10, 20) {real, imag} */,
  {32'h3f4f3e3a, 32'hbf4fc331} /* (28, 10, 19) {real, imag} */,
  {32'hbf81e910, 32'hbeb8b617} /* (28, 10, 18) {real, imag} */,
  {32'hbdc11fc4, 32'h3f3bfa82} /* (28, 10, 17) {real, imag} */,
  {32'hbfb34f4c, 32'h3fe62484} /* (28, 10, 16) {real, imag} */,
  {32'hbf53aca8, 32'hbfa70d84} /* (28, 10, 15) {real, imag} */,
  {32'hbf8fd182, 32'h3f951148} /* (28, 10, 14) {real, imag} */,
  {32'h4094ce2b, 32'hbfbe7ced} /* (28, 10, 13) {real, imag} */,
  {32'h401cf79e, 32'h3f285c0f} /* (28, 10, 12) {real, imag} */,
  {32'hbfd038b9, 32'hc00faeac} /* (28, 10, 11) {real, imag} */,
  {32'h3f986544, 32'h3e7c278b} /* (28, 10, 10) {real, imag} */,
  {32'h3f80cba6, 32'hc0156a34} /* (28, 10, 9) {real, imag} */,
  {32'hbdc5bafa, 32'h3b55281d} /* (28, 10, 8) {real, imag} */,
  {32'h405249a1, 32'hc020cc01} /* (28, 10, 7) {real, imag} */,
  {32'h3d09571e, 32'h40255b6e} /* (28, 10, 6) {real, imag} */,
  {32'hbff9839d, 32'h3f916e3a} /* (28, 10, 5) {real, imag} */,
  {32'hbfef864e, 32'hbfc31565} /* (28, 10, 4) {real, imag} */,
  {32'hbdff1f40, 32'h3fa06c05} /* (28, 10, 3) {real, imag} */,
  {32'hc016a007, 32'h40274b08} /* (28, 10, 2) {real, imag} */,
  {32'h3f259192, 32'hc07db59b} /* (28, 10, 1) {real, imag} */,
  {32'h40543155, 32'h4084879a} /* (28, 10, 0) {real, imag} */,
  {32'h3fbbb751, 32'hc007a556} /* (28, 9, 31) {real, imag} */,
  {32'hc0bce4e9, 32'hbf8af65f} /* (28, 9, 30) {real, imag} */,
  {32'hbf9496ca, 32'h40534b9f} /* (28, 9, 29) {real, imag} */,
  {32'h406fcb32, 32'hbfda2b9e} /* (28, 9, 28) {real, imag} */,
  {32'h3ff2e5b3, 32'h406b8948} /* (28, 9, 27) {real, imag} */,
  {32'h40218bdc, 32'hc0508525} /* (28, 9, 26) {real, imag} */,
  {32'hbfe17dfe, 32'hc049886b} /* (28, 9, 25) {real, imag} */,
  {32'h3f005ee1, 32'hbf4ca706} /* (28, 9, 24) {real, imag} */,
  {32'hbf74748f, 32'hbe477d9d} /* (28, 9, 23) {real, imag} */,
  {32'h4090b68a, 32'h3f8359d2} /* (28, 9, 22) {real, imag} */,
  {32'h3fed58ce, 32'h40447b56} /* (28, 9, 21) {real, imag} */,
  {32'h3f3b92c7, 32'hc0220a1a} /* (28, 9, 20) {real, imag} */,
  {32'hbf56aca9, 32'hbde6a04d} /* (28, 9, 19) {real, imag} */,
  {32'hbe6ef564, 32'h3fd7ff4c} /* (28, 9, 18) {real, imag} */,
  {32'hbf2b41e4, 32'h3fa67a0e} /* (28, 9, 17) {real, imag} */,
  {32'h3e915dde, 32'h3f8e01cd} /* (28, 9, 16) {real, imag} */,
  {32'hbf4532a5, 32'hbeed04ee} /* (28, 9, 15) {real, imag} */,
  {32'hbdc00a17, 32'hbf973ca5} /* (28, 9, 14) {real, imag} */,
  {32'h401be979, 32'h3cb8ef85} /* (28, 9, 13) {real, imag} */,
  {32'h3f725ddc, 32'hbf7acc24} /* (28, 9, 12) {real, imag} */,
  {32'hc0075137, 32'hbfac046c} /* (28, 9, 11) {real, imag} */,
  {32'hbfe8a169, 32'h4007d171} /* (28, 9, 10) {real, imag} */,
  {32'h3d9430b5, 32'hc00bcfb2} /* (28, 9, 9) {real, imag} */,
  {32'h4018d338, 32'hbdedf27e} /* (28, 9, 8) {real, imag} */,
  {32'hbfe355d0, 32'hbf824fe0} /* (28, 9, 7) {real, imag} */,
  {32'hbf56308f, 32'h3f59e19c} /* (28, 9, 6) {real, imag} */,
  {32'hc02b0222, 32'hc07571a4} /* (28, 9, 5) {real, imag} */,
  {32'h403f20da, 32'hbfb4ae58} /* (28, 9, 4) {real, imag} */,
  {32'hbe9245e5, 32'h3e3ce781} /* (28, 9, 3) {real, imag} */,
  {32'hbfdbd98d, 32'h4096984e} /* (28, 9, 2) {real, imag} */,
  {32'h3fc08a5b, 32'hbed8ee8e} /* (28, 9, 1) {real, imag} */,
  {32'h3fe3ee44, 32'hbffe17a8} /* (28, 9, 0) {real, imag} */,
  {32'hc033ada7, 32'h41181725} /* (28, 8, 31) {real, imag} */,
  {32'hc06295a1, 32'hc0e2f547} /* (28, 8, 30) {real, imag} */,
  {32'h3f8464f7, 32'hc0250a53} /* (28, 8, 29) {real, imag} */,
  {32'hbe4fb669, 32'h3f1d7811} /* (28, 8, 28) {real, imag} */,
  {32'h3f9d2b4a, 32'hbe8ca92a} /* (28, 8, 27) {real, imag} */,
  {32'hc043b5d4, 32'hc07685ee} /* (28, 8, 26) {real, imag} */,
  {32'h3ee6ec84, 32'h3f9d4f38} /* (28, 8, 25) {real, imag} */,
  {32'hc086a581, 32'hc001bf7e} /* (28, 8, 24) {real, imag} */,
  {32'h400f1b12, 32'h3f828a35} /* (28, 8, 23) {real, imag} */,
  {32'h3f9e9d57, 32'hc08b57d8} /* (28, 8, 22) {real, imag} */,
  {32'hbf381b0a, 32'hbfae6ac5} /* (28, 8, 21) {real, imag} */,
  {32'hbf895bd7, 32'h40bf00b4} /* (28, 8, 20) {real, imag} */,
  {32'hbf96b5df, 32'h3da91710} /* (28, 8, 19) {real, imag} */,
  {32'hbf950cb7, 32'h3f5445c4} /* (28, 8, 18) {real, imag} */,
  {32'h3e9fa726, 32'hbf55fb8d} /* (28, 8, 17) {real, imag} */,
  {32'h3f21b1c1, 32'h3e6cb8fa} /* (28, 8, 16) {real, imag} */,
  {32'h3ef7686a, 32'hbf6e726a} /* (28, 8, 15) {real, imag} */,
  {32'hbfaa325b, 32'hbf67f300} /* (28, 8, 14) {real, imag} */,
  {32'hbf11cd46, 32'hbf3e4a05} /* (28, 8, 13) {real, imag} */,
  {32'hbe4050e7, 32'h4044ac53} /* (28, 8, 12) {real, imag} */,
  {32'h3e3c9fa6, 32'h3e530964} /* (28, 8, 11) {real, imag} */,
  {32'h3fb29765, 32'h3f84ad9b} /* (28, 8, 10) {real, imag} */,
  {32'h3fd64dd1, 32'h3fbd6146} /* (28, 8, 9) {real, imag} */,
  {32'h3f8547c9, 32'hc0693079} /* (28, 8, 8) {real, imag} */,
  {32'h3f9bd4c6, 32'h403654c3} /* (28, 8, 7) {real, imag} */,
  {32'h3f8e1766, 32'hbfe3016d} /* (28, 8, 6) {real, imag} */,
  {32'h3fc5b72a, 32'h4071f2cf} /* (28, 8, 5) {real, imag} */,
  {32'hbf343a0c, 32'h40081829} /* (28, 8, 4) {real, imag} */,
  {32'hc0915586, 32'hbf168c9c} /* (28, 8, 3) {real, imag} */,
  {32'h40759d92, 32'hc0060cd3} /* (28, 8, 2) {real, imag} */,
  {32'hc00d24a4, 32'h4101b241} /* (28, 8, 1) {real, imag} */,
  {32'hc06ad888, 32'h410a298c} /* (28, 8, 0) {real, imag} */,
  {32'hc0211cb3, 32'h3faf36b2} /* (28, 7, 31) {real, imag} */,
  {32'h407bc3b4, 32'hbf875e90} /* (28, 7, 30) {real, imag} */,
  {32'hbf62fb5e, 32'hbf417e5a} /* (28, 7, 29) {real, imag} */,
  {32'hc0190a04, 32'h4093e1ff} /* (28, 7, 28) {real, imag} */,
  {32'hc007cc51, 32'hbf0b0101} /* (28, 7, 27) {real, imag} */,
  {32'h4044163c, 32'h3fee0c64} /* (28, 7, 26) {real, imag} */,
  {32'hbe6c13f1, 32'hbf85f4a6} /* (28, 7, 25) {real, imag} */,
  {32'h40b99d2b, 32'hbef1ebdd} /* (28, 7, 24) {real, imag} */,
  {32'hbf83a962, 32'hbff1c73d} /* (28, 7, 23) {real, imag} */,
  {32'h3d7dce85, 32'h3f820ad8} /* (28, 7, 22) {real, imag} */,
  {32'hbfd1b067, 32'hbf15c220} /* (28, 7, 21) {real, imag} */,
  {32'hc05927d5, 32'h3f7b78ed} /* (28, 7, 20) {real, imag} */,
  {32'h3f3ec830, 32'hc002aa3f} /* (28, 7, 19) {real, imag} */,
  {32'hbf9fdfcf, 32'hbfea44b2} /* (28, 7, 18) {real, imag} */,
  {32'h3f65dd1f, 32'hbfe18916} /* (28, 7, 17) {real, imag} */,
  {32'hbfbae3ba, 32'hbf921620} /* (28, 7, 16) {real, imag} */,
  {32'hbf65ee18, 32'h3ea89a25} /* (28, 7, 15) {real, imag} */,
  {32'h3ffbd4cc, 32'h3f9ae7e2} /* (28, 7, 14) {real, imag} */,
  {32'h401700f1, 32'hbe3d275e} /* (28, 7, 13) {real, imag} */,
  {32'hbfad2662, 32'h3f5561c5} /* (28, 7, 12) {real, imag} */,
  {32'h4042ee7e, 32'h3f89b3fc} /* (28, 7, 11) {real, imag} */,
  {32'h3f7fe3ed, 32'hbf6e7884} /* (28, 7, 10) {real, imag} */,
  {32'hc0113eae, 32'h400496dc} /* (28, 7, 9) {real, imag} */,
  {32'hbea5d736, 32'h3fa83128} /* (28, 7, 8) {real, imag} */,
  {32'hbf5c6220, 32'hc02cd9e2} /* (28, 7, 7) {real, imag} */,
  {32'hbfc54346, 32'hbef1bc8f} /* (28, 7, 6) {real, imag} */,
  {32'hbed8f2e5, 32'hc08304b8} /* (28, 7, 5) {real, imag} */,
  {32'h4093fb78, 32'h401a5ccd} /* (28, 7, 4) {real, imag} */,
  {32'hbfa4ad75, 32'h404ad35f} /* (28, 7, 3) {real, imag} */,
  {32'hc0c04ffe, 32'hc0f9d384} /* (28, 7, 2) {real, imag} */,
  {32'hbfc898a5, 32'h3eb47eea} /* (28, 7, 1) {real, imag} */,
  {32'h3f7cb4d9, 32'hbf47fbc3} /* (28, 7, 0) {real, imag} */,
  {32'h40a5fd73, 32'h3f349049} /* (28, 6, 31) {real, imag} */,
  {32'hc0d9d2fe, 32'hbfaef098} /* (28, 6, 30) {real, imag} */,
  {32'hc049b4a2, 32'hbfb0f998} /* (28, 6, 29) {real, imag} */,
  {32'h3fce4fd9, 32'h40a1a0c0} /* (28, 6, 28) {real, imag} */,
  {32'h40b14066, 32'h3f36719a} /* (28, 6, 27) {real, imag} */,
  {32'hc01f36e7, 32'h40cd044a} /* (28, 6, 26) {real, imag} */,
  {32'h3fdba8df, 32'h3f9f811d} /* (28, 6, 25) {real, imag} */,
  {32'h3f0211f4, 32'hc09c2a86} /* (28, 6, 24) {real, imag} */,
  {32'hbfb2c32b, 32'h3f520d4a} /* (28, 6, 23) {real, imag} */,
  {32'hc0110ce3, 32'h3fa5667a} /* (28, 6, 22) {real, imag} */,
  {32'h3e6cd0c5, 32'h4075163b} /* (28, 6, 21) {real, imag} */,
  {32'h3da30289, 32'h3fb2fd23} /* (28, 6, 20) {real, imag} */,
  {32'hbfa14995, 32'h3f3d3efb} /* (28, 6, 19) {real, imag} */,
  {32'h3f34962f, 32'hc002696c} /* (28, 6, 18) {real, imag} */,
  {32'hbfaaf57a, 32'h3fcba35d} /* (28, 6, 17) {real, imag} */,
  {32'h3e03923d, 32'h3f2037fe} /* (28, 6, 16) {real, imag} */,
  {32'h3f8667fd, 32'h3ee1b908} /* (28, 6, 15) {real, imag} */,
  {32'h3ffdaa5e, 32'h3fe7c17f} /* (28, 6, 14) {real, imag} */,
  {32'hbf9b09f6, 32'hc0307474} /* (28, 6, 13) {real, imag} */,
  {32'hbc91c8fe, 32'hbd590fbf} /* (28, 6, 12) {real, imag} */,
  {32'h4014f598, 32'h3d655cf5} /* (28, 6, 11) {real, imag} */,
  {32'hbed0f436, 32'h3f8c1334} /* (28, 6, 10) {real, imag} */,
  {32'h40886f94, 32'hbc419dbb} /* (28, 6, 9) {real, imag} */,
  {32'h3fb4d835, 32'hbfa88c20} /* (28, 6, 8) {real, imag} */,
  {32'hbd6a3f72, 32'h3f83627d} /* (28, 6, 7) {real, imag} */,
  {32'h3f8ab697, 32'h40ac9ac2} /* (28, 6, 6) {real, imag} */,
  {32'h4008468b, 32'h402fddb2} /* (28, 6, 5) {real, imag} */,
  {32'h4067b802, 32'hbf3f83c2} /* (28, 6, 4) {real, imag} */,
  {32'hbf3c757f, 32'h400b8af5} /* (28, 6, 3) {real, imag} */,
  {32'h4003a936, 32'hbf0573b5} /* (28, 6, 2) {real, imag} */,
  {32'h404bd348, 32'h40ca37ce} /* (28, 6, 1) {real, imag} */,
  {32'hc07b48ec, 32'hc06f52a1} /* (28, 6, 0) {real, imag} */,
  {32'h4190779a, 32'h417d56a4} /* (28, 5, 31) {real, imag} */,
  {32'hc013a504, 32'hc0f7df37} /* (28, 5, 30) {real, imag} */,
  {32'h3e0df25f, 32'h4040e73f} /* (28, 5, 29) {real, imag} */,
  {32'hbfd0d1df, 32'hbfd49da7} /* (28, 5, 28) {real, imag} */,
  {32'hc0090f67, 32'hc05cf097} /* (28, 5, 27) {real, imag} */,
  {32'h3f9cfacd, 32'h408d0954} /* (28, 5, 26) {real, imag} */,
  {32'hc086ab95, 32'h40057588} /* (28, 5, 25) {real, imag} */,
  {32'h401641df, 32'h3ff2230d} /* (28, 5, 24) {real, imag} */,
  {32'hbf9a1513, 32'hbfeebc8c} /* (28, 5, 23) {real, imag} */,
  {32'hbd8d0dce, 32'hbe6c5352} /* (28, 5, 22) {real, imag} */,
  {32'hbfdad2b2, 32'hc0642c35} /* (28, 5, 21) {real, imag} */,
  {32'hbea1c70c, 32'hbf1075dc} /* (28, 5, 20) {real, imag} */,
  {32'h3ff7d555, 32'hbf71547f} /* (28, 5, 19) {real, imag} */,
  {32'hbf79296e, 32'hbf5d4b3e} /* (28, 5, 18) {real, imag} */,
  {32'hc003fafc, 32'hbe527bda} /* (28, 5, 17) {real, imag} */,
  {32'h3de246a6, 32'h3f5ff73d} /* (28, 5, 16) {real, imag} */,
  {32'h3ed1cb8e, 32'h3df3d72e} /* (28, 5, 15) {real, imag} */,
  {32'h3e1a312a, 32'h3f2289cd} /* (28, 5, 14) {real, imag} */,
  {32'hc00d7367, 32'h3fc30b93} /* (28, 5, 13) {real, imag} */,
  {32'hbfb35aeb, 32'h40032483} /* (28, 5, 12) {real, imag} */,
  {32'hbf80a6a5, 32'h3fc6c642} /* (28, 5, 11) {real, imag} */,
  {32'h3d86f96f, 32'hbfb6e87d} /* (28, 5, 10) {real, imag} */,
  {32'hbfa30339, 32'h3f3e5da0} /* (28, 5, 9) {real, imag} */,
  {32'h3f776bf0, 32'h3ec6960d} /* (28, 5, 8) {real, imag} */,
  {32'hc071abe9, 32'h3f16fa45} /* (28, 5, 7) {real, imag} */,
  {32'h3ffe57af, 32'hc0869a9c} /* (28, 5, 6) {real, imag} */,
  {32'h40765dfa, 32'h3fa7e5ad} /* (28, 5, 5) {real, imag} */,
  {32'hc00a00a7, 32'h408a66ea} /* (28, 5, 4) {real, imag} */,
  {32'hbf62f4c1, 32'hc0973345} /* (28, 5, 3) {real, imag} */,
  {32'h40cd7f53, 32'hc0f3b139} /* (28, 5, 2) {real, imag} */,
  {32'hc0ea40ea, 32'h419535ba} /* (28, 5, 1) {real, imag} */,
  {32'hc0086bf0, 32'h41494cfd} /* (28, 5, 0) {real, imag} */,
  {32'h408e88b4, 32'hc13490eb} /* (28, 4, 31) {real, imag} */,
  {32'hc06b3588, 32'h40e44e7e} /* (28, 4, 30) {real, imag} */,
  {32'h404aa862, 32'hc0e699af} /* (28, 4, 29) {real, imag} */,
  {32'h40419bd6, 32'hc1312b4f} /* (28, 4, 28) {real, imag} */,
  {32'h3e60b2d4, 32'h40e4b1be} /* (28, 4, 27) {real, imag} */,
  {32'h3fc8d40f, 32'hbfa9dc95} /* (28, 4, 26) {real, imag} */,
  {32'hbf2132df, 32'h401500bc} /* (28, 4, 25) {real, imag} */,
  {32'h40596cd9, 32'hbe8e15df} /* (28, 4, 24) {real, imag} */,
  {32'hbf1c108f, 32'h3f4f27e3} /* (28, 4, 23) {real, imag} */,
  {32'hbf898d35, 32'h3e88198c} /* (28, 4, 22) {real, imag} */,
  {32'hbfb527e4, 32'h405f8d07} /* (28, 4, 21) {real, imag} */,
  {32'h3cb7e85c, 32'h3de5e575} /* (28, 4, 20) {real, imag} */,
  {32'hbfc0032f, 32'h3f3abadf} /* (28, 4, 19) {real, imag} */,
  {32'h408c5787, 32'hc02c4799} /* (28, 4, 18) {real, imag} */,
  {32'h3e2aa35c, 32'hc018b69e} /* (28, 4, 17) {real, imag} */,
  {32'h3ed289c6, 32'h3f07dae8} /* (28, 4, 16) {real, imag} */,
  {32'h3fbd7c0d, 32'hbe24e5dd} /* (28, 4, 15) {real, imag} */,
  {32'hbf96e9aa, 32'h3e6292da} /* (28, 4, 14) {real, imag} */,
  {32'hc03d947f, 32'h3fe8381f} /* (28, 4, 13) {real, imag} */,
  {32'h3fc9e7ee, 32'hbea7d92e} /* (28, 4, 12) {real, imag} */,
  {32'h3fe48a25, 32'hbf42d7c4} /* (28, 4, 11) {real, imag} */,
  {32'h40bc5284, 32'h3f6fab6e} /* (28, 4, 10) {real, imag} */,
  {32'hbe0baf7a, 32'hbcd3abdb} /* (28, 4, 9) {real, imag} */,
  {32'hbeca6dc6, 32'h3f9f8fc5} /* (28, 4, 8) {real, imag} */,
  {32'h3fc16cc6, 32'hbf977432} /* (28, 4, 7) {real, imag} */,
  {32'hbfb7eced, 32'hbf09694d} /* (28, 4, 6) {real, imag} */,
  {32'hc1020aac, 32'h3f89661c} /* (28, 4, 5) {real, imag} */,
  {32'hbce8de18, 32'hbf81e48f} /* (28, 4, 4) {real, imag} */,
  {32'hc0410f25, 32'h4028b712} /* (28, 4, 3) {real, imag} */,
  {32'hc16e7d42, 32'h4179cf63} /* (28, 4, 2) {real, imag} */,
  {32'h40a15b95, 32'hc1b065c4} /* (28, 4, 1) {real, imag} */,
  {32'h40a1d8c4, 32'hc17c9e3a} /* (28, 4, 0) {real, imag} */,
  {32'h41d2b196, 32'h412aff60} /* (28, 3, 31) {real, imag} */,
  {32'hc186eb88, 32'h3ebe6c21} /* (28, 3, 30) {real, imag} */,
  {32'h40f4506e, 32'hbe069131} /* (28, 3, 29) {real, imag} */,
  {32'hbda3f672, 32'hc037d2a5} /* (28, 3, 28) {real, imag} */,
  {32'h404c7d1a, 32'h40046f1e} /* (28, 3, 27) {real, imag} */,
  {32'hc082049d, 32'h4048f17b} /* (28, 3, 26) {real, imag} */,
  {32'hc08f357f, 32'hc007a2b1} /* (28, 3, 25) {real, imag} */,
  {32'hc0bfdd3c, 32'h405eba9f} /* (28, 3, 24) {real, imag} */,
  {32'hc050ea24, 32'h3edc8c1e} /* (28, 3, 23) {real, imag} */,
  {32'h3e92aeaf, 32'hbeb7e8ee} /* (28, 3, 22) {real, imag} */,
  {32'h3fc76b7b, 32'h3e575774} /* (28, 3, 21) {real, imag} */,
  {32'hbf522cae, 32'hbdae6340} /* (28, 3, 20) {real, imag} */,
  {32'h400624bc, 32'hbf88f456} /* (28, 3, 19) {real, imag} */,
  {32'h3ef2723d, 32'h3f7fe4c0} /* (28, 3, 18) {real, imag} */,
  {32'h40372d01, 32'h3e775184} /* (28, 3, 17) {real, imag} */,
  {32'hbf683918, 32'h3e9a769e} /* (28, 3, 16) {real, imag} */,
  {32'h3e46ea41, 32'h3f875574} /* (28, 3, 15) {real, imag} */,
  {32'h3e252ff7, 32'hbf64ae63} /* (28, 3, 14) {real, imag} */,
  {32'hbe59bacd, 32'hbf974f89} /* (28, 3, 13) {real, imag} */,
  {32'h3e298183, 32'h3f705d2e} /* (28, 3, 12) {real, imag} */,
  {32'h4017a4c9, 32'hbe43c503} /* (28, 3, 11) {real, imag} */,
  {32'hbfe8ce6e, 32'h40401d89} /* (28, 3, 10) {real, imag} */,
  {32'h3e7dbd14, 32'h40474690} /* (28, 3, 9) {real, imag} */,
  {32'h3eeacea7, 32'hc0666f30} /* (28, 3, 8) {real, imag} */,
  {32'hc0dc7eec, 32'hbff1c779} /* (28, 3, 7) {real, imag} */,
  {32'hc05ecff1, 32'h404bc3a7} /* (28, 3, 6) {real, imag} */,
  {32'hc04292dd, 32'hc08f6722} /* (28, 3, 5) {real, imag} */,
  {32'hc0dc7505, 32'h408ecc45} /* (28, 3, 4) {real, imag} */,
  {32'h4070aadc, 32'hc12a09aa} /* (28, 3, 3) {real, imag} */,
  {32'hc12a4cb1, 32'h413675b7} /* (28, 3, 2) {real, imag} */,
  {32'h4126716e, 32'hc1ee3c59} /* (28, 3, 1) {real, imag} */,
  {32'h41336d8d, 32'hbfd50841} /* (28, 3, 0) {real, imag} */,
  {32'h41847eef, 32'h4299b604} /* (28, 2, 31) {real, imag} */,
  {32'hc1be7cca, 32'hc237fb5b} /* (28, 2, 30) {real, imag} */,
  {32'h406d31cc, 32'h40b9549b} /* (28, 2, 29) {real, imag} */,
  {32'h414b7da9, 32'h41037185} /* (28, 2, 28) {real, imag} */,
  {32'hbfc36d5f, 32'h400c0275} /* (28, 2, 27) {real, imag} */,
  {32'h3e0b00fd, 32'hbe84a4e7} /* (28, 2, 26) {real, imag} */,
  {32'hbf54daa7, 32'h4040ca0e} /* (28, 2, 25) {real, imag} */,
  {32'hc087c7f0, 32'hc093bbe7} /* (28, 2, 24) {real, imag} */,
  {32'h4011f205, 32'h4069d4b3} /* (28, 2, 23) {real, imag} */,
  {32'h405b96e1, 32'hc00b9834} /* (28, 2, 22) {real, imag} */,
  {32'hc04ab0f1, 32'hc0006b50} /* (28, 2, 21) {real, imag} */,
  {32'h3f9c8fb1, 32'hbfa5037d} /* (28, 2, 20) {real, imag} */,
  {32'h3fe25252, 32'hbccc0ea2} /* (28, 2, 19) {real, imag} */,
  {32'hc0392a72, 32'h3fe9e4d1} /* (28, 2, 18) {real, imag} */,
  {32'h3ea5eba1, 32'hbec08774} /* (28, 2, 17) {real, imag} */,
  {32'hbfffdf68, 32'h3fe9bf47} /* (28, 2, 16) {real, imag} */,
  {32'h3fc5a361, 32'h3fa0233c} /* (28, 2, 15) {real, imag} */,
  {32'h3e077e67, 32'hc013ca58} /* (28, 2, 14) {real, imag} */,
  {32'h3f78674e, 32'h3efef6ef} /* (28, 2, 13) {real, imag} */,
  {32'hbfab0afe, 32'hbd164d32} /* (28, 2, 12) {real, imag} */,
  {32'h400fb283, 32'hc09889f8} /* (28, 2, 11) {real, imag} */,
  {32'h3f54dd40, 32'hbfb26a98} /* (28, 2, 10) {real, imag} */,
  {32'h3ff7d26a, 32'hbf821546} /* (28, 2, 9) {real, imag} */,
  {32'hbe46dd04, 32'hc0694703} /* (28, 2, 8) {real, imag} */,
  {32'hc04c536e, 32'h40412846} /* (28, 2, 7) {real, imag} */,
  {32'h40a4b623, 32'h3fb86729} /* (28, 2, 6) {real, imag} */,
  {32'hbe9a6503, 32'hc15e1578} /* (28, 2, 5) {real, imag} */,
  {32'h41397d6a, 32'h416014e9} /* (28, 2, 4) {real, imag} */,
  {32'hbfec2131, 32'hc0476acc} /* (28, 2, 3) {real, imag} */,
  {32'hc128dc08, 32'hc1ad4b29} /* (28, 2, 2) {real, imag} */,
  {32'h41540e86, 32'h4229ffb7} /* (28, 2, 1) {real, imag} */,
  {32'h40bddd35, 32'h422f47c3} /* (28, 2, 0) {real, imag} */,
  {32'hc1f846e9, 32'hc297ad61} /* (28, 1, 31) {real, imag} */,
  {32'h3f86e60b, 32'h41ead033} /* (28, 1, 30) {real, imag} */,
  {32'h40782d77, 32'hc01fddc9} /* (28, 1, 29) {real, imag} */,
  {32'hc078edbc, 32'hc0b0b6e9} /* (28, 1, 28) {real, imag} */,
  {32'h414e30bd, 32'h41608355} /* (28, 1, 27) {real, imag} */,
  {32'hbe31e5bb, 32'h40781325} /* (28, 1, 26) {real, imag} */,
  {32'hbfeb043e, 32'h3fe931bb} /* (28, 1, 25) {real, imag} */,
  {32'h40814e4e, 32'h402646a6} /* (28, 1, 24) {real, imag} */,
  {32'h3fa937a6, 32'h3fef9820} /* (28, 1, 23) {real, imag} */,
  {32'hc0823008, 32'hc08b7f47} /* (28, 1, 22) {real, imag} */,
  {32'h40d54d63, 32'hbf7b1802} /* (28, 1, 21) {real, imag} */,
  {32'hbf2544dc, 32'hbfe95c1e} /* (28, 1, 20) {real, imag} */,
  {32'h3f94715b, 32'h3fe70035} /* (28, 1, 19) {real, imag} */,
  {32'h3c4986f2, 32'h4081babf} /* (28, 1, 18) {real, imag} */,
  {32'hbfba89d8, 32'hbd7e8d30} /* (28, 1, 17) {real, imag} */,
  {32'hbfceb193, 32'h3eee13dd} /* (28, 1, 16) {real, imag} */,
  {32'hbeff0de6, 32'h3f3f81bf} /* (28, 1, 15) {real, imag} */,
  {32'hc0484c0c, 32'hbf4a479a} /* (28, 1, 14) {real, imag} */,
  {32'h3e972fce, 32'hbe4cc2f4} /* (28, 1, 13) {real, imag} */,
  {32'hbdd0917f, 32'hc04048e9} /* (28, 1, 12) {real, imag} */,
  {32'hc03dc3b7, 32'h3f7687af} /* (28, 1, 11) {real, imag} */,
  {32'hbf42b01e, 32'hbeaacc9d} /* (28, 1, 10) {real, imag} */,
  {32'h400ef6bf, 32'hc0868bec} /* (28, 1, 9) {real, imag} */,
  {32'hc0b37989, 32'h4088a5be} /* (28, 1, 8) {real, imag} */,
  {32'h40927df3, 32'hc03ce5d6} /* (28, 1, 7) {real, imag} */,
  {32'h3fb848df, 32'h409bbce7} /* (28, 1, 6) {real, imag} */,
  {32'h3ecf40a8, 32'h41172f38} /* (28, 1, 5) {real, imag} */,
  {32'h40be14b6, 32'hc101d080} /* (28, 1, 4) {real, imag} */,
  {32'h4071ea86, 32'h40fa3c9f} /* (28, 1, 3) {real, imag} */,
  {32'hc1c317df, 32'h425ee6e3} /* (28, 1, 2) {real, imag} */,
  {32'h40e7006a, 32'hc2e4c5b8} /* (28, 1, 1) {real, imag} */,
  {32'hc1c80f1d, 32'hc26f6af6} /* (28, 1, 0) {real, imag} */,
  {32'hc25be04b, 32'hc202f6bb} /* (28, 0, 31) {real, imag} */,
  {32'h418b47f7, 32'hbfdbe539} /* (28, 0, 30) {real, imag} */,
  {32'h40967372, 32'h411ba78e} /* (28, 0, 29) {real, imag} */,
  {32'h4047d27e, 32'hc0905c56} /* (28, 0, 28) {real, imag} */,
  {32'h3efd30e6, 32'h40d831b1} /* (28, 0, 27) {real, imag} */,
  {32'hbfcfaba1, 32'h404bc282} /* (28, 0, 26) {real, imag} */,
  {32'hc0a99bc5, 32'h3fd59e07} /* (28, 0, 25) {real, imag} */,
  {32'h4087034b, 32'h3f1312f6} /* (28, 0, 24) {real, imag} */,
  {32'h40a0f3b0, 32'hc0311608} /* (28, 0, 23) {real, imag} */,
  {32'hba70eff8, 32'h4072353f} /* (28, 0, 22) {real, imag} */,
  {32'h40190d63, 32'h3fb221e0} /* (28, 0, 21) {real, imag} */,
  {32'hbe2ade7a, 32'h3ee71309} /* (28, 0, 20) {real, imag} */,
  {32'hbea3a473, 32'h403d9d20} /* (28, 0, 19) {real, imag} */,
  {32'h3fd3de62, 32'h3ee5505b} /* (28, 0, 18) {real, imag} */,
  {32'h3f5f462e, 32'h3ef13711} /* (28, 0, 17) {real, imag} */,
  {32'h3f99023b, 32'h3ef26135} /* (28, 0, 16) {real, imag} */,
  {32'hbfcd545c, 32'hbf2c61e7} /* (28, 0, 15) {real, imag} */,
  {32'hc084a11f, 32'h3f923215} /* (28, 0, 14) {real, imag} */,
  {32'hbe99f321, 32'hbe4554b0} /* (28, 0, 13) {real, imag} */,
  {32'h3f550d7c, 32'h3e4384fe} /* (28, 0, 12) {real, imag} */,
  {32'h3f0467b7, 32'h40978442} /* (28, 0, 11) {real, imag} */,
  {32'h4042ef8d, 32'h3f6b0428} /* (28, 0, 10) {real, imag} */,
  {32'hc09478e6, 32'h40be9dcc} /* (28, 0, 9) {real, imag} */,
  {32'hbfe685ad, 32'h403bcf93} /* (28, 0, 8) {real, imag} */,
  {32'h40a9dbd3, 32'hc04be6d4} /* (28, 0, 7) {real, imag} */,
  {32'h405a41ca, 32'hbd32855c} /* (28, 0, 6) {real, imag} */,
  {32'h40ecbeb1, 32'h41014cc7} /* (28, 0, 5) {real, imag} */,
  {32'hc0475a4e, 32'h40a7bf94} /* (28, 0, 4) {real, imag} */,
  {32'h3f91e829, 32'hc0b50e8f} /* (28, 0, 3) {real, imag} */,
  {32'hc18101bc, 32'h404ddff0} /* (28, 0, 2) {real, imag} */,
  {32'h419928ba, 32'hc2766e9a} /* (28, 0, 1) {real, imag} */,
  {32'hc1c0d8dc, 32'hc2292b7d} /* (28, 0, 0) {real, imag} */,
  {32'h41f0874a, 32'h413b802b} /* (27, 31, 31) {real, imag} */,
  {32'hc1c3a727, 32'hc1362d5a} /* (27, 31, 30) {real, imag} */,
  {32'hbfb3d9f7, 32'h404ff685} /* (27, 31, 29) {real, imag} */,
  {32'h4018f32d, 32'h408c1844} /* (27, 31, 28) {real, imag} */,
  {32'hc0607d42, 32'hbc802d18} /* (27, 31, 27) {real, imag} */,
  {32'h40025ce8, 32'h3f495afd} /* (27, 31, 26) {real, imag} */,
  {32'h3f4948e3, 32'hc03d81ec} /* (27, 31, 25) {real, imag} */,
  {32'hc014941d, 32'h3fd30dd7} /* (27, 31, 24) {real, imag} */,
  {32'hc04e1db6, 32'h3f6ad560} /* (27, 31, 23) {real, imag} */,
  {32'h400626f2, 32'hbefdd859} /* (27, 31, 22) {real, imag} */,
  {32'hc04d1370, 32'h3f5dfee8} /* (27, 31, 21) {real, imag} */,
  {32'h3e0aee17, 32'hc027db4c} /* (27, 31, 20) {real, imag} */,
  {32'hbeb92a98, 32'hbcc8b997} /* (27, 31, 19) {real, imag} */,
  {32'hbf3373a9, 32'h3f8a30ac} /* (27, 31, 18) {real, imag} */,
  {32'hbdb1ecd5, 32'h3f2fe896} /* (27, 31, 17) {real, imag} */,
  {32'hbf801fb0, 32'h3dc45d4a} /* (27, 31, 16) {real, imag} */,
  {32'hc004e58c, 32'hbf2f0935} /* (27, 31, 15) {real, imag} */,
  {32'h409e1ee8, 32'h3f9b1a93} /* (27, 31, 14) {real, imag} */,
  {32'hbeec0151, 32'h3e577fa0} /* (27, 31, 13) {real, imag} */,
  {32'hbfc5472d, 32'h3f14f934} /* (27, 31, 12) {real, imag} */,
  {32'h3fb7df63, 32'hbff775b8} /* (27, 31, 11) {real, imag} */,
  {32'h4005cc47, 32'hbfb53b23} /* (27, 31, 10) {real, imag} */,
  {32'h3f5f104f, 32'h3fc50179} /* (27, 31, 9) {real, imag} */,
  {32'hbfd81ed3, 32'hc036b250} /* (27, 31, 8) {real, imag} */,
  {32'hbfd91ea6, 32'h3ef8bb81} /* (27, 31, 7) {real, imag} */,
  {32'hbfcb4d0b, 32'h3f4bff48} /* (27, 31, 6) {real, imag} */,
  {32'hc0c948a1, 32'hc09b7a59} /* (27, 31, 5) {real, imag} */,
  {32'h40c3c742, 32'hbf60b2ec} /* (27, 31, 4) {real, imag} */,
  {32'h3ffed1bc, 32'hc07cfbf3} /* (27, 31, 3) {real, imag} */,
  {32'hc057f2af, 32'hc02372a3} /* (27, 31, 2) {real, imag} */,
  {32'h41122117, 32'h41b0298d} /* (27, 31, 1) {real, imag} */,
  {32'h41459674, 32'h419a32ba} /* (27, 31, 0) {real, imag} */,
  {32'hc093818b, 32'hc13a6913} /* (27, 30, 31) {real, imag} */,
  {32'h404f8a8b, 32'h41a00a3f} /* (27, 30, 30) {real, imag} */,
  {32'hbfedf73f, 32'hc105c269} /* (27, 30, 29) {real, imag} */,
  {32'hc10634bc, 32'hbfed488a} /* (27, 30, 28) {real, imag} */,
  {32'h4100a4de, 32'h3f6c5326} /* (27, 30, 27) {real, imag} */,
  {32'hc017585c, 32'hc03f7f11} /* (27, 30, 26) {real, imag} */,
  {32'h3e06d04c, 32'hc081bd4c} /* (27, 30, 25) {real, imag} */,
  {32'h401c05ae, 32'h402c3680} /* (27, 30, 24) {real, imag} */,
  {32'hc007738b, 32'h3fab94ef} /* (27, 30, 23) {real, imag} */,
  {32'h3eaabd67, 32'h3fd53c84} /* (27, 30, 22) {real, imag} */,
  {32'h3fbb3e14, 32'h3fca6bc1} /* (27, 30, 21) {real, imag} */,
  {32'hbf22afa0, 32'hbeded270} /* (27, 30, 20) {real, imag} */,
  {32'hbe2310a7, 32'h3d322e36} /* (27, 30, 19) {real, imag} */,
  {32'h3f213394, 32'h3ee044e4} /* (27, 30, 18) {real, imag} */,
  {32'h3e0cbd60, 32'hbc72ed7d} /* (27, 30, 17) {real, imag} */,
  {32'hbfa54b41, 32'hbfd7d883} /* (27, 30, 16) {real, imag} */,
  {32'h40470f29, 32'h3f30cd4a} /* (27, 30, 15) {real, imag} */,
  {32'hbfb3f172, 32'h3e99989e} /* (27, 30, 14) {real, imag} */,
  {32'h3e3bade1, 32'hbfa6613f} /* (27, 30, 13) {real, imag} */,
  {32'hbf99e90d, 32'h4046f0dc} /* (27, 30, 12) {real, imag} */,
  {32'h3f9764fa, 32'hbe0c1de5} /* (27, 30, 11) {real, imag} */,
  {32'hbfd269ff, 32'h3fe6cbec} /* (27, 30, 10) {real, imag} */,
  {32'h3f908d58, 32'h4017a708} /* (27, 30, 9) {real, imag} */,
  {32'h3e39bfc9, 32'hc0821c3b} /* (27, 30, 8) {real, imag} */,
  {32'hc0079ac3, 32'hc0025595} /* (27, 30, 7) {real, imag} */,
  {32'h3f33072a, 32'h406a7b7a} /* (27, 30, 6) {real, imag} */,
  {32'h4073739d, 32'h4105d7a4} /* (27, 30, 5) {real, imag} */,
  {32'h40f84785, 32'hc0c819f0} /* (27, 30, 4) {real, imag} */,
  {32'hc038effb, 32'hc0a97526} /* (27, 30, 3) {real, imag} */,
  {32'h4097097e, 32'h41cf2c64} /* (27, 30, 2) {real, imag} */,
  {32'hc136e0ad, 32'hc1fb6439} /* (27, 30, 1) {real, imag} */,
  {32'hc008cb01, 32'hbfd00d3f} /* (27, 30, 0) {real, imag} */,
  {32'h41a1700a, 32'h3f8d8ff1} /* (27, 29, 31) {real, imag} */,
  {32'hc0c3df69, 32'hc065fbcb} /* (27, 29, 30) {real, imag} */,
  {32'h40b09664, 32'h3ece51df} /* (27, 29, 29) {real, imag} */,
  {32'h3e04b724, 32'hc0a2c8c7} /* (27, 29, 28) {real, imag} */,
  {32'h40c70d87, 32'h401f3264} /* (27, 29, 27) {real, imag} */,
  {32'h3e3670a5, 32'hc06f508c} /* (27, 29, 26) {real, imag} */,
  {32'hbf0c92a6, 32'hbdcea0f7} /* (27, 29, 25) {real, imag} */,
  {32'h401c83ce, 32'h3f5cbf02} /* (27, 29, 24) {real, imag} */,
  {32'h3e8afb8d, 32'h3e9b9b31} /* (27, 29, 23) {real, imag} */,
  {32'h4004257d, 32'h3f16f761} /* (27, 29, 22) {real, imag} */,
  {32'h3f6862d5, 32'h3f81f1d3} /* (27, 29, 21) {real, imag} */,
  {32'h3fd09b47, 32'h40737cc2} /* (27, 29, 20) {real, imag} */,
  {32'h3f8b2bcd, 32'hbf012f23} /* (27, 29, 19) {real, imag} */,
  {32'h402ec3d2, 32'hbe33bd40} /* (27, 29, 18) {real, imag} */,
  {32'hbfcad96b, 32'hbf37486f} /* (27, 29, 17) {real, imag} */,
  {32'hbf905fad, 32'hbfd3d5e1} /* (27, 29, 16) {real, imag} */,
  {32'hbe0006cd, 32'hbfbaec90} /* (27, 29, 15) {real, imag} */,
  {32'hc01c5a30, 32'hbb737b2c} /* (27, 29, 14) {real, imag} */,
  {32'h3fadbfd4, 32'h3fbe038d} /* (27, 29, 13) {real, imag} */,
  {32'hbe3718b0, 32'h3ff9d36a} /* (27, 29, 12) {real, imag} */,
  {32'h3f95a72e, 32'h3e940fa9} /* (27, 29, 11) {real, imag} */,
  {32'h3fa56779, 32'h3ff95acc} /* (27, 29, 10) {real, imag} */,
  {32'h40163d8f, 32'hc019e6b1} /* (27, 29, 9) {real, imag} */,
  {32'hbfce2121, 32'hc00a8a83} /* (27, 29, 8) {real, imag} */,
  {32'h3cb6057a, 32'hc06b8ee1} /* (27, 29, 7) {real, imag} */,
  {32'hc02cc475, 32'h4034d93e} /* (27, 29, 6) {real, imag} */,
  {32'hbf131618, 32'hc08f01f5} /* (27, 29, 5) {real, imag} */,
  {32'h3fde757e, 32'h3f3c18d0} /* (27, 29, 4) {real, imag} */,
  {32'h3f72a659, 32'hc097a7c7} /* (27, 29, 3) {real, imag} */,
  {32'hc064c0c9, 32'h4060ef6b} /* (27, 29, 2) {real, imag} */,
  {32'hc113464c, 32'hbf850d83} /* (27, 29, 1) {real, imag} */,
  {32'hc0be0f01, 32'hc04e89a2} /* (27, 29, 0) {real, imag} */,
  {32'h40d167ae, 32'h4011a9c7} /* (27, 28, 31) {real, imag} */,
  {32'hc1104b52, 32'hc011871f} /* (27, 28, 30) {real, imag} */,
  {32'h3c847f3f, 32'hbfdda250} /* (27, 28, 29) {real, imag} */,
  {32'hc005bdb6, 32'hbfca8684} /* (27, 28, 28) {real, imag} */,
  {32'hbf728cb8, 32'hbf53e868} /* (27, 28, 27) {real, imag} */,
  {32'hc09d94e5, 32'hbeb312c1} /* (27, 28, 26) {real, imag} */,
  {32'h3f58d8c9, 32'h3f79e9b4} /* (27, 28, 25) {real, imag} */,
  {32'hbfb6185f, 32'hbe06a849} /* (27, 28, 24) {real, imag} */,
  {32'hbfed25d4, 32'h40276d15} /* (27, 28, 23) {real, imag} */,
  {32'hbf184884, 32'h3f7bdc25} /* (27, 28, 22) {real, imag} */,
  {32'h3fc6a016, 32'hbfbf70c6} /* (27, 28, 21) {real, imag} */,
  {32'h3f077251, 32'hbfbbb9bd} /* (27, 28, 20) {real, imag} */,
  {32'h4035cc54, 32'h3f323201} /* (27, 28, 19) {real, imag} */,
  {32'hc02c2cdc, 32'hbfa0875f} /* (27, 28, 18) {real, imag} */,
  {32'hbec9cb55, 32'h3f669be9} /* (27, 28, 17) {real, imag} */,
  {32'h3e2445be, 32'h3f409260} /* (27, 28, 16) {real, imag} */,
  {32'hbecceedd, 32'hbfdc2dbd} /* (27, 28, 15) {real, imag} */,
  {32'hbebd6b4f, 32'hbecdab2f} /* (27, 28, 14) {real, imag} */,
  {32'h3ddbf666, 32'hbffdff5c} /* (27, 28, 13) {real, imag} */,
  {32'hbed2ea8a, 32'hbf85115f} /* (27, 28, 12) {real, imag} */,
  {32'hbf1d5bd1, 32'hc0025c36} /* (27, 28, 11) {real, imag} */,
  {32'h3e837953, 32'h3f9e4f82} /* (27, 28, 10) {real, imag} */,
  {32'hbfbf75bb, 32'hbf94de1d} /* (27, 28, 9) {real, imag} */,
  {32'hbfef9a82, 32'hc0024658} /* (27, 28, 8) {real, imag} */,
  {32'h401f2b4d, 32'hc0a3e6ef} /* (27, 28, 7) {real, imag} */,
  {32'h3f21a316, 32'h40d3b4f0} /* (27, 28, 6) {real, imag} */,
  {32'h40823a65, 32'h3fdce113} /* (27, 28, 5) {real, imag} */,
  {32'h40a1dd7a, 32'h40956ca2} /* (27, 28, 4) {real, imag} */,
  {32'hbf6512a6, 32'h3f549fd3} /* (27, 28, 3) {real, imag} */,
  {32'hc12ccdc3, 32'h410117d8} /* (27, 28, 2) {real, imag} */,
  {32'h402fd995, 32'h3ee1e5cb} /* (27, 28, 1) {real, imag} */,
  {32'h41312030, 32'h4035a22a} /* (27, 28, 0) {real, imag} */,
  {32'hc0f4dcc6, 32'hc0c1b4ae} /* (27, 27, 31) {real, imag} */,
  {32'hc0909846, 32'hbef19a38} /* (27, 27, 30) {real, imag} */,
  {32'hbf503096, 32'hbf88b712} /* (27, 27, 29) {real, imag} */,
  {32'hbd5fa857, 32'h40974581} /* (27, 27, 28) {real, imag} */,
  {32'h3fea0327, 32'h401b0258} /* (27, 27, 27) {real, imag} */,
  {32'h40664fe6, 32'h3e561a66} /* (27, 27, 26) {real, imag} */,
  {32'h40652a28, 32'hbfffcab4} /* (27, 27, 25) {real, imag} */,
  {32'hbee496a6, 32'hbde6a6af} /* (27, 27, 24) {real, imag} */,
  {32'hbfa9e7a7, 32'h3ea1c918} /* (27, 27, 23) {real, imag} */,
  {32'hbe4f32f7, 32'hbe832ddd} /* (27, 27, 22) {real, imag} */,
  {32'h40033778, 32'hbf1d0c8a} /* (27, 27, 21) {real, imag} */,
  {32'hbfc683a0, 32'h3ec2022a} /* (27, 27, 20) {real, imag} */,
  {32'hbfafe74d, 32'hbff7d59f} /* (27, 27, 19) {real, imag} */,
  {32'hbfc1a4a4, 32'hc0200d61} /* (27, 27, 18) {real, imag} */,
  {32'h3f4b842b, 32'h3f16d0f2} /* (27, 27, 17) {real, imag} */,
  {32'hbefc070f, 32'h3ebdf3eb} /* (27, 27, 16) {real, imag} */,
  {32'hbecab523, 32'hbf043559} /* (27, 27, 15) {real, imag} */,
  {32'hbfa71920, 32'h3ce9454c} /* (27, 27, 14) {real, imag} */,
  {32'h3c8257ef, 32'hbfa27efc} /* (27, 27, 13) {real, imag} */,
  {32'h3ec27b29, 32'h3f28fde9} /* (27, 27, 12) {real, imag} */,
  {32'hbecef7eb, 32'h3ffa7f68} /* (27, 27, 11) {real, imag} */,
  {32'h400e096f, 32'hbfc3376d} /* (27, 27, 10) {real, imag} */,
  {32'h3fcadd4b, 32'hc01fa993} /* (27, 27, 9) {real, imag} */,
  {32'h4078f31b, 32'h40595302} /* (27, 27, 8) {real, imag} */,
  {32'h402c385e, 32'h3e910810} /* (27, 27, 7) {real, imag} */,
  {32'h3ee1a944, 32'hc0262d57} /* (27, 27, 6) {real, imag} */,
  {32'hbf0739ee, 32'h3fb27c4c} /* (27, 27, 5) {real, imag} */,
  {32'hc04d8572, 32'hbf024562} /* (27, 27, 4) {real, imag} */,
  {32'h4050b7a0, 32'hc0217033} /* (27, 27, 3) {real, imag} */,
  {32'h40281f28, 32'h3e885dee} /* (27, 27, 2) {real, imag} */,
  {32'hc0272efd, 32'hc01246b0} /* (27, 27, 1) {real, imag} */,
  {32'hc1122386, 32'hc07b6cf7} /* (27, 27, 0) {real, imag} */,
  {32'hc0b84561, 32'h3ed7c82b} /* (27, 26, 31) {real, imag} */,
  {32'h403a9f94, 32'hbfc82ef9} /* (27, 26, 30) {real, imag} */,
  {32'hbeb7cc61, 32'h40412712} /* (27, 26, 29) {real, imag} */,
  {32'hbfc5c414, 32'hbf9e479f} /* (27, 26, 28) {real, imag} */,
  {32'hc03b5608, 32'hbe4eec0a} /* (27, 26, 27) {real, imag} */,
  {32'h40510580, 32'h403a86c0} /* (27, 26, 26) {real, imag} */,
  {32'hbfe249bf, 32'h3e6ffc0f} /* (27, 26, 25) {real, imag} */,
  {32'h403fe0e8, 32'hc01c6eb1} /* (27, 26, 24) {real, imag} */,
  {32'h3f6d8a42, 32'hbe880aa6} /* (27, 26, 23) {real, imag} */,
  {32'h40909daa, 32'h3fe10b9c} /* (27, 26, 22) {real, imag} */,
  {32'hbda0fdb6, 32'h40612fbc} /* (27, 26, 21) {real, imag} */,
  {32'h3f1d57c3, 32'hbf63911a} /* (27, 26, 20) {real, imag} */,
  {32'hbf925132, 32'h400a0770} /* (27, 26, 19) {real, imag} */,
  {32'h3f1b3d98, 32'h3ec87fb9} /* (27, 26, 18) {real, imag} */,
  {32'hbf98fccc, 32'h3e426bc2} /* (27, 26, 17) {real, imag} */,
  {32'h3ea5105e, 32'hc0410c77} /* (27, 26, 16) {real, imag} */,
  {32'hbf6e1eb2, 32'h403a6208} /* (27, 26, 15) {real, imag} */,
  {32'hc0446eb9, 32'h3dfe8523} /* (27, 26, 14) {real, imag} */,
  {32'hbf84bad3, 32'h3ed76af8} /* (27, 26, 13) {real, imag} */,
  {32'h3fabd762, 32'hbfd1a2d4} /* (27, 26, 12) {real, imag} */,
  {32'h3fc543ac, 32'h3f1fd771} /* (27, 26, 11) {real, imag} */,
  {32'h3f116813, 32'h3f8d8c2b} /* (27, 26, 10) {real, imag} */,
  {32'h3fd8386f, 32'h3f2a26f6} /* (27, 26, 9) {real, imag} */,
  {32'h3f8921ea, 32'h3f4f8e42} /* (27, 26, 8) {real, imag} */,
  {32'hc01f10c4, 32'h3d6f3431} /* (27, 26, 7) {real, imag} */,
  {32'hbf764cb1, 32'h3f05d391} /* (27, 26, 6) {real, imag} */,
  {32'h3f418cc0, 32'h3eecbbf2} /* (27, 26, 5) {real, imag} */,
  {32'hbfc8e110, 32'hc0649cfb} /* (27, 26, 4) {real, imag} */,
  {32'h3e6f5746, 32'h3f51ff86} /* (27, 26, 3) {real, imag} */,
  {32'h3fb37722, 32'h404f20e0} /* (27, 26, 2) {real, imag} */,
  {32'h3f1ae0b8, 32'hc0b3aa13} /* (27, 26, 1) {real, imag} */,
  {32'h3f20dc05, 32'h3fc0e2b4} /* (27, 26, 0) {real, imag} */,
  {32'h40e38bbf, 32'h405d41b7} /* (27, 25, 31) {real, imag} */,
  {32'hc04a77ee, 32'hbfcbc35b} /* (27, 25, 30) {real, imag} */,
  {32'h402bee61, 32'h3f7c0ab8} /* (27, 25, 29) {real, imag} */,
  {32'hbef6e11f, 32'hc093ade1} /* (27, 25, 28) {real, imag} */,
  {32'hbfc528cc, 32'h400afc01} /* (27, 25, 27) {real, imag} */,
  {32'h402c0ae2, 32'hc0a96982} /* (27, 25, 26) {real, imag} */,
  {32'hc0878dfb, 32'h3eb40064} /* (27, 25, 25) {real, imag} */,
  {32'hc03e6fef, 32'hc01102e8} /* (27, 25, 24) {real, imag} */,
  {32'h4046c4df, 32'h3f9cb95d} /* (27, 25, 23) {real, imag} */,
  {32'h3f632e9e, 32'h3f26b4b5} /* (27, 25, 22) {real, imag} */,
  {32'h3f0aca99, 32'hc07f2085} /* (27, 25, 21) {real, imag} */,
  {32'h3f08916d, 32'h3db71cc2} /* (27, 25, 20) {real, imag} */,
  {32'h4024690b, 32'hbf77fc15} /* (27, 25, 19) {real, imag} */,
  {32'hbdf25361, 32'h3f608bb5} /* (27, 25, 18) {real, imag} */,
  {32'h3d62b7de, 32'h3f8718ba} /* (27, 25, 17) {real, imag} */,
  {32'hbfdf2bee, 32'h3f128fbc} /* (27, 25, 16) {real, imag} */,
  {32'h3f96d2d2, 32'hbfe88aac} /* (27, 25, 15) {real, imag} */,
  {32'hbfe687e5, 32'hbfac1dbd} /* (27, 25, 14) {real, imag} */,
  {32'hc022efd2, 32'h3fad5e61} /* (27, 25, 13) {real, imag} */,
  {32'h3f2ed021, 32'hc01ae579} /* (27, 25, 12) {real, imag} */,
  {32'hc001cdb3, 32'h4021d753} /* (27, 25, 11) {real, imag} */,
  {32'hbf9ade38, 32'hbff5d54a} /* (27, 25, 10) {real, imag} */,
  {32'hbf698581, 32'hc0828555} /* (27, 25, 9) {real, imag} */,
  {32'h4090bf8b, 32'h408804c1} /* (27, 25, 8) {real, imag} */,
  {32'h40b898cf, 32'hc035fbcf} /* (27, 25, 7) {real, imag} */,
  {32'h3fbbc27a, 32'hbde26aa3} /* (27, 25, 6) {real, imag} */,
  {32'h407b4371, 32'hbe0cc8a0} /* (27, 25, 5) {real, imag} */,
  {32'hbf42f68e, 32'hbf87126e} /* (27, 25, 4) {real, imag} */,
  {32'hbfdbcada, 32'h404daef7} /* (27, 25, 3) {real, imag} */,
  {32'hbf8fc1ff, 32'h3f8627ea} /* (27, 25, 2) {real, imag} */,
  {32'hbd4bd0c0, 32'h405ec0af} /* (27, 25, 1) {real, imag} */,
  {32'hc01f65cc, 32'hbed500df} /* (27, 25, 0) {real, imag} */,
  {32'hc01cef36, 32'hbeba0d0e} /* (27, 24, 31) {real, imag} */,
  {32'hc017bb41, 32'h3f7d76b0} /* (27, 24, 30) {real, imag} */,
  {32'h3d54cad2, 32'h3fc152b0} /* (27, 24, 29) {real, imag} */,
  {32'hc05c5d2c, 32'hbfa2d2e7} /* (27, 24, 28) {real, imag} */,
  {32'hbfa80aad, 32'hbea94e13} /* (27, 24, 27) {real, imag} */,
  {32'hc0277f0f, 32'hbfcbc753} /* (27, 24, 26) {real, imag} */,
  {32'h3fa54d06, 32'h3f811eb5} /* (27, 24, 25) {real, imag} */,
  {32'h3e0fcca6, 32'hbf9b61e9} /* (27, 24, 24) {real, imag} */,
  {32'h3fe93622, 32'hbf63d655} /* (27, 24, 23) {real, imag} */,
  {32'hbfc56cbb, 32'hbfa446b6} /* (27, 24, 22) {real, imag} */,
  {32'h3f885d6d, 32'h401fa70e} /* (27, 24, 21) {real, imag} */,
  {32'hbfb9a342, 32'hbe8673a1} /* (27, 24, 20) {real, imag} */,
  {32'hbebee095, 32'h3f826334} /* (27, 24, 19) {real, imag} */,
  {32'h4021a876, 32'h3e34b07b} /* (27, 24, 18) {real, imag} */,
  {32'h3dc903a1, 32'h3de9a344} /* (27, 24, 17) {real, imag} */,
  {32'h3f870503, 32'hbfc88c85} /* (27, 24, 16) {real, imag} */,
  {32'hbf4c0a7e, 32'hbfe0441e} /* (27, 24, 15) {real, imag} */,
  {32'hbfb0ee06, 32'hbf93f940} /* (27, 24, 14) {real, imag} */,
  {32'hbf67f26d, 32'hbfc0c93e} /* (27, 24, 13) {real, imag} */,
  {32'h3fd292fb, 32'hbfdd6393} /* (27, 24, 12) {real, imag} */,
  {32'h3f77e49b, 32'h404d86b0} /* (27, 24, 11) {real, imag} */,
  {32'hc057e571, 32'hc021db4f} /* (27, 24, 10) {real, imag} */,
  {32'hbe6f3d14, 32'h400061da} /* (27, 24, 9) {real, imag} */,
  {32'h408c3f64, 32'h405a3a91} /* (27, 24, 8) {real, imag} */,
  {32'h408a7d9d, 32'h3f1e5827} /* (27, 24, 7) {real, imag} */,
  {32'hbf91f928, 32'h402b1978} /* (27, 24, 6) {real, imag} */,
  {32'h3fbc4363, 32'hbf68de19} /* (27, 24, 5) {real, imag} */,
  {32'hbfcb0572, 32'hbfa8ad70} /* (27, 24, 4) {real, imag} */,
  {32'h3f89a3af, 32'h3fdec7b5} /* (27, 24, 3) {real, imag} */,
  {32'h3fce8ef6, 32'hbeb33a66} /* (27, 24, 2) {real, imag} */,
  {32'hbfee2973, 32'hc0a0dfab} /* (27, 24, 1) {real, imag} */,
  {32'hc0516c3f, 32'hbeb3b691} /* (27, 24, 0) {real, imag} */,
  {32'hbfc6cb47, 32'hc03c9fe1} /* (27, 23, 31) {real, imag} */,
  {32'h3f83ff41, 32'h40462b80} /* (27, 23, 30) {real, imag} */,
  {32'h3fc606b8, 32'h4045b338} /* (27, 23, 29) {real, imag} */,
  {32'h404026a1, 32'h3f340ccf} /* (27, 23, 28) {real, imag} */,
  {32'h3fc24979, 32'hbe46bd8c} /* (27, 23, 27) {real, imag} */,
  {32'hbf5c842a, 32'hc0449b4d} /* (27, 23, 26) {real, imag} */,
  {32'h40490474, 32'hbfff9c75} /* (27, 23, 25) {real, imag} */,
  {32'hbf37efeb, 32'h3ef6272c} /* (27, 23, 24) {real, imag} */,
  {32'h3da16d77, 32'h3e81f1fa} /* (27, 23, 23) {real, imag} */,
  {32'hbfbb6337, 32'h3ef38df4} /* (27, 23, 22) {real, imag} */,
  {32'h3f6f426e, 32'h3f291b72} /* (27, 23, 21) {real, imag} */,
  {32'h3fa6bc4e, 32'hbeb6ea12} /* (27, 23, 20) {real, imag} */,
  {32'hbf6ea113, 32'h3f92a2ad} /* (27, 23, 19) {real, imag} */,
  {32'h3fe0f21e, 32'h3f6e37f5} /* (27, 23, 18) {real, imag} */,
  {32'hc01f9b3c, 32'h403942f4} /* (27, 23, 17) {real, imag} */,
  {32'h3fe898a1, 32'hbf94b62a} /* (27, 23, 16) {real, imag} */,
  {32'hc013e270, 32'hbfa35734} /* (27, 23, 15) {real, imag} */,
  {32'hbf2f1d76, 32'h400f1755} /* (27, 23, 14) {real, imag} */,
  {32'h3f111837, 32'hbfe97a9c} /* (27, 23, 13) {real, imag} */,
  {32'hc01a8be7, 32'hbfabb8e5} /* (27, 23, 12) {real, imag} */,
  {32'h4050c463, 32'hc00f0951} /* (27, 23, 11) {real, imag} */,
  {32'h4058406a, 32'hc00b3912} /* (27, 23, 10) {real, imag} */,
  {32'hbfa04efc, 32'hbe985573} /* (27, 23, 9) {real, imag} */,
  {32'hbf1a746c, 32'hbe930b38} /* (27, 23, 8) {real, imag} */,
  {32'hbf09a3fe, 32'h3f0acad6} /* (27, 23, 7) {real, imag} */,
  {32'hc06f1d8e, 32'h4006f92e} /* (27, 23, 6) {real, imag} */,
  {32'hc0336e72, 32'hc00f84ad} /* (27, 23, 5) {real, imag} */,
  {32'hbec2bb50, 32'h3ff906ae} /* (27, 23, 4) {real, imag} */,
  {32'hbee01ea8, 32'hbfa148ed} /* (27, 23, 3) {real, imag} */,
  {32'hc05c621c, 32'hbf61d454} /* (27, 23, 2) {real, imag} */,
  {32'h40abc1b7, 32'hc01ce76e} /* (27, 23, 1) {real, imag} */,
  {32'hc03370e3, 32'hbeed0818} /* (27, 23, 0) {real, imag} */,
  {32'h40539100, 32'h3fcba251} /* (27, 22, 31) {real, imag} */,
  {32'h3fd59a25, 32'hbe115172} /* (27, 22, 30) {real, imag} */,
  {32'hbfa62d74, 32'h3eb64c4c} /* (27, 22, 29) {real, imag} */,
  {32'h3f8643f3, 32'h3ee4817b} /* (27, 22, 28) {real, imag} */,
  {32'h3ecea807, 32'hc0300066} /* (27, 22, 27) {real, imag} */,
  {32'hbff4988d, 32'h401c594d} /* (27, 22, 26) {real, imag} */,
  {32'hbf444414, 32'hbe862679} /* (27, 22, 25) {real, imag} */,
  {32'h40670953, 32'hbf8294ac} /* (27, 22, 24) {real, imag} */,
  {32'hc0385d8a, 32'h4020fef0} /* (27, 22, 23) {real, imag} */,
  {32'hbfd8e992, 32'h403d3ec2} /* (27, 22, 22) {real, imag} */,
  {32'h400e2585, 32'h3fa85ae8} /* (27, 22, 21) {real, imag} */,
  {32'hbf212563, 32'hbf4ddfad} /* (27, 22, 20) {real, imag} */,
  {32'hc039bb14, 32'hbe0d027e} /* (27, 22, 19) {real, imag} */,
  {32'h3ea89044, 32'h3cd4cada} /* (27, 22, 18) {real, imag} */,
  {32'hbe84dacf, 32'hc047cca7} /* (27, 22, 17) {real, imag} */,
  {32'h3f803f66, 32'h404a80ff} /* (27, 22, 16) {real, imag} */,
  {32'hbeeeeb59, 32'h3e1f1827} /* (27, 22, 15) {real, imag} */,
  {32'h3f751cb9, 32'hbef832ee} /* (27, 22, 14) {real, imag} */,
  {32'h3fcf4747, 32'hc0146463} /* (27, 22, 13) {real, imag} */,
  {32'hc00c7958, 32'h3e403587} /* (27, 22, 12) {real, imag} */,
  {32'h3f2d385e, 32'hbe83c52b} /* (27, 22, 11) {real, imag} */,
  {32'hbf5257ea, 32'h3f334998} /* (27, 22, 10) {real, imag} */,
  {32'hbf06d8ce, 32'hc0198881} /* (27, 22, 9) {real, imag} */,
  {32'hbe8bc86e, 32'h4001cae0} /* (27, 22, 8) {real, imag} */,
  {32'h3fe7fced, 32'hbe95b110} /* (27, 22, 7) {real, imag} */,
  {32'hbe2f80b5, 32'h3e4e9b7d} /* (27, 22, 6) {real, imag} */,
  {32'hbede51ce, 32'hbf17ddb3} /* (27, 22, 5) {real, imag} */,
  {32'h40245036, 32'hc00fa842} /* (27, 22, 4) {real, imag} */,
  {32'h3f628772, 32'h40454d46} /* (27, 22, 3) {real, imag} */,
  {32'hbe249ea4, 32'h3fa481a2} /* (27, 22, 2) {real, imag} */,
  {32'hc051ab04, 32'hbf0131c8} /* (27, 22, 1) {real, imag} */,
  {32'h40a09d74, 32'hc0630413} /* (27, 22, 0) {real, imag} */,
  {32'hbfee2c20, 32'h3fe016db} /* (27, 21, 31) {real, imag} */,
  {32'hbf9329b7, 32'h3f831c0c} /* (27, 21, 30) {real, imag} */,
  {32'h3cd5c127, 32'h3d2d495d} /* (27, 21, 29) {real, imag} */,
  {32'hbe9c77fb, 32'hbff002b3} /* (27, 21, 28) {real, imag} */,
  {32'h3fa11385, 32'hbe039194} /* (27, 21, 27) {real, imag} */,
  {32'h402ff600, 32'h4013e432} /* (27, 21, 26) {real, imag} */,
  {32'hbfa1e2bc, 32'h3f1d4dae} /* (27, 21, 25) {real, imag} */,
  {32'h3e2bff6f, 32'hbf507e74} /* (27, 21, 24) {real, imag} */,
  {32'hbc6a7e41, 32'h409f9c6b} /* (27, 21, 23) {real, imag} */,
  {32'hc04cba86, 32'h3f5c0d4c} /* (27, 21, 22) {real, imag} */,
  {32'h3f3d226f, 32'hc0916bad} /* (27, 21, 21) {real, imag} */,
  {32'h3f3f1553, 32'h3e76daea} /* (27, 21, 20) {real, imag} */,
  {32'h3fcfe771, 32'hbf4b7a9e} /* (27, 21, 19) {real, imag} */,
  {32'h3f8c76a5, 32'hbe0a75b0} /* (27, 21, 18) {real, imag} */,
  {32'hbf6d71a8, 32'h4038ae65} /* (27, 21, 17) {real, imag} */,
  {32'h3f61d80d, 32'h3ead965d} /* (27, 21, 16) {real, imag} */,
  {32'h3f5bb3e5, 32'hbf47ec73} /* (27, 21, 15) {real, imag} */,
  {32'hbf97b6d0, 32'h401db7cf} /* (27, 21, 14) {real, imag} */,
  {32'h3fe51997, 32'h3c94d058} /* (27, 21, 13) {real, imag} */,
  {32'h3fca881c, 32'hbf802ca8} /* (27, 21, 12) {real, imag} */,
  {32'h3edbaf5f, 32'h4005f873} /* (27, 21, 11) {real, imag} */,
  {32'h3f7714d4, 32'h3e7ada90} /* (27, 21, 10) {real, imag} */,
  {32'h3f818db5, 32'h3e6f3c5b} /* (27, 21, 9) {real, imag} */,
  {32'hc013f3ff, 32'h3e567170} /* (27, 21, 8) {real, imag} */,
  {32'hbfdc3560, 32'h3efdf25a} /* (27, 21, 7) {real, imag} */,
  {32'hbf48f719, 32'h3fe0e37d} /* (27, 21, 6) {real, imag} */,
  {32'h40479bd2, 32'hbd9af95c} /* (27, 21, 5) {real, imag} */,
  {32'hbfde736b, 32'hbfdf34d9} /* (27, 21, 4) {real, imag} */,
  {32'hbec97f4e, 32'h3fb41a08} /* (27, 21, 3) {real, imag} */,
  {32'h3fc94a29, 32'hc023bd4d} /* (27, 21, 2) {real, imag} */,
  {32'h4017d5e3, 32'hbec488b1} /* (27, 21, 1) {real, imag} */,
  {32'hc02204ea, 32'hc01cdce3} /* (27, 21, 0) {real, imag} */,
  {32'h3fbe8eca, 32'h3ecda98e} /* (27, 20, 31) {real, imag} */,
  {32'hbf6b018f, 32'hbfc44c6b} /* (27, 20, 30) {real, imag} */,
  {32'hbe415c79, 32'hbf117062} /* (27, 20, 29) {real, imag} */,
  {32'hbf496fd9, 32'h3f4e93a7} /* (27, 20, 28) {real, imag} */,
  {32'hbd8a3259, 32'h402f83f1} /* (27, 20, 27) {real, imag} */,
  {32'hc00533b6, 32'h3e8a66b0} /* (27, 20, 26) {real, imag} */,
  {32'h4039ac44, 32'hc002e359} /* (27, 20, 25) {real, imag} */,
  {32'h3f0029f4, 32'hbf9f5f8c} /* (27, 20, 24) {real, imag} */,
  {32'h3f9a10b0, 32'hbf5d4e92} /* (27, 20, 23) {real, imag} */,
  {32'h3ec00ed7, 32'h3f07758a} /* (27, 20, 22) {real, imag} */,
  {32'hc0520705, 32'hbfd98205} /* (27, 20, 21) {real, imag} */,
  {32'hbfb74f4b, 32'h3e52b13f} /* (27, 20, 20) {real, imag} */,
  {32'h3c6b81df, 32'h3fe0cb13} /* (27, 20, 19) {real, imag} */,
  {32'h3fd5ad9e, 32'hc01835d3} /* (27, 20, 18) {real, imag} */,
  {32'h3f0557b2, 32'hbdf189f7} /* (27, 20, 17) {real, imag} */,
  {32'h3ec41525, 32'h3ecccb72} /* (27, 20, 16) {real, imag} */,
  {32'h3f3ca4de, 32'hc02e0353} /* (27, 20, 15) {real, imag} */,
  {32'hbe6a2e64, 32'h3f8ae92c} /* (27, 20, 14) {real, imag} */,
  {32'h3f3ff40f, 32'hbf51d6c7} /* (27, 20, 13) {real, imag} */,
  {32'h3f862225, 32'hbd6527c5} /* (27, 20, 12) {real, imag} */,
  {32'h3e95204c, 32'h401f2b56} /* (27, 20, 11) {real, imag} */,
  {32'hbfdf3f0c, 32'h3efd44dd} /* (27, 20, 10) {real, imag} */,
  {32'h3fd0fb73, 32'h40018b83} /* (27, 20, 9) {real, imag} */,
  {32'h4034fad4, 32'hbfd05d66} /* (27, 20, 8) {real, imag} */,
  {32'h3ebff6b9, 32'hbfc718af} /* (27, 20, 7) {real, imag} */,
  {32'hbfa13b05, 32'hbfee11f9} /* (27, 20, 6) {real, imag} */,
  {32'h400900bb, 32'hbfaa7226} /* (27, 20, 5) {real, imag} */,
  {32'hbf8c6c8a, 32'h3fb1fafc} /* (27, 20, 4) {real, imag} */,
  {32'hbf5b0193, 32'h3fe863aa} /* (27, 20, 3) {real, imag} */,
  {32'hbff82369, 32'h40057cfb} /* (27, 20, 2) {real, imag} */,
  {32'hbfb9a7f7, 32'h3f3c284e} /* (27, 20, 1) {real, imag} */,
  {32'h4020fad2, 32'h3f983e67} /* (27, 20, 0) {real, imag} */,
  {32'hbfad07e9, 32'hbf9c1afd} /* (27, 19, 31) {real, imag} */,
  {32'h3e74479b, 32'h3fa0795d} /* (27, 19, 30) {real, imag} */,
  {32'h4011aa42, 32'hbf640024} /* (27, 19, 29) {real, imag} */,
  {32'h3ecc0e99, 32'hbf020344} /* (27, 19, 28) {real, imag} */,
  {32'h3fd4213e, 32'h3e1bc280} /* (27, 19, 27) {real, imag} */,
  {32'hbfbf2f28, 32'hbfdaf5d3} /* (27, 19, 26) {real, imag} */,
  {32'h3fad94e0, 32'hbe5707d1} /* (27, 19, 25) {real, imag} */,
  {32'h3fb4c84a, 32'h4030b606} /* (27, 19, 24) {real, imag} */,
  {32'h3f98e492, 32'hbf005669} /* (27, 19, 23) {real, imag} */,
  {32'h3d6d70a5, 32'h3f91bf6d} /* (27, 19, 22) {real, imag} */,
  {32'h3f8a97dc, 32'hbf36b6db} /* (27, 19, 21) {real, imag} */,
  {32'hbedc322c, 32'hbfcd0a86} /* (27, 19, 20) {real, imag} */,
  {32'hbfe4263f, 32'h3f8fb466} /* (27, 19, 19) {real, imag} */,
  {32'hbf01c955, 32'h409b55ad} /* (27, 19, 18) {real, imag} */,
  {32'h3f09fecd, 32'hbf92e69c} /* (27, 19, 17) {real, imag} */,
  {32'h3da4954b, 32'h3ee3a2ca} /* (27, 19, 16) {real, imag} */,
  {32'h3f975547, 32'hbe9d70ce} /* (27, 19, 15) {real, imag} */,
  {32'hbfb3ad3d, 32'hbfd32c24} /* (27, 19, 14) {real, imag} */,
  {32'hbd62c332, 32'h3ea56690} /* (27, 19, 13) {real, imag} */,
  {32'h3fe3f62c, 32'h3f013d3e} /* (27, 19, 12) {real, imag} */,
  {32'hc01aa770, 32'hc00f59bc} /* (27, 19, 11) {real, imag} */,
  {32'h3ff1c1b4, 32'hc08ec3a7} /* (27, 19, 10) {real, imag} */,
  {32'hbfc96116, 32'h405836e5} /* (27, 19, 9) {real, imag} */,
  {32'h3f179cb0, 32'h3ea9b76a} /* (27, 19, 8) {real, imag} */,
  {32'h3fd82137, 32'h400f5e48} /* (27, 19, 7) {real, imag} */,
  {32'h4006cd13, 32'hbefcb7da} /* (27, 19, 6) {real, imag} */,
  {32'hc0238465, 32'h3fc4aead} /* (27, 19, 5) {real, imag} */,
  {32'h3e3ada87, 32'h3f9f2377} /* (27, 19, 4) {real, imag} */,
  {32'h4028577e, 32'hbf772884} /* (27, 19, 3) {real, imag} */,
  {32'hbe3ae9fc, 32'hbfba0139} /* (27, 19, 2) {real, imag} */,
  {32'h3e8a999b, 32'h3fda5709} /* (27, 19, 1) {real, imag} */,
  {32'hc0087b36, 32'hc0136a0c} /* (27, 19, 0) {real, imag} */,
  {32'hc032010f, 32'hbf0fbe3a} /* (27, 18, 31) {real, imag} */,
  {32'h40512989, 32'hbf93e7de} /* (27, 18, 30) {real, imag} */,
  {32'h3f46f243, 32'h3eabd956} /* (27, 18, 29) {real, imag} */,
  {32'hc0162f48, 32'h3f97068e} /* (27, 18, 28) {real, imag} */,
  {32'h3e08dec3, 32'hc019c64c} /* (27, 18, 27) {real, imag} */,
  {32'h3ea59b4e, 32'hbfa64bd1} /* (27, 18, 26) {real, imag} */,
  {32'hbebd436d, 32'hbfa7c023} /* (27, 18, 25) {real, imag} */,
  {32'h3fe8be4d, 32'hbf837988} /* (27, 18, 24) {real, imag} */,
  {32'hbeba3c6c, 32'hc03c90cc} /* (27, 18, 23) {real, imag} */,
  {32'h3f9c9100, 32'hbfcd32cd} /* (27, 18, 22) {real, imag} */,
  {32'hc02d05d1, 32'h402595b7} /* (27, 18, 21) {real, imag} */,
  {32'h40098b50, 32'h3fc17466} /* (27, 18, 20) {real, imag} */,
  {32'h3f9d8633, 32'hbfbe0e67} /* (27, 18, 19) {real, imag} */,
  {32'h3ee50b9b, 32'h3fdd43a5} /* (27, 18, 18) {real, imag} */,
  {32'hbf9bc091, 32'h3f269a77} /* (27, 18, 17) {real, imag} */,
  {32'h3f40e3a9, 32'hbfd1ac27} /* (27, 18, 16) {real, imag} */,
  {32'h3fcfeb1a, 32'h402f3dcf} /* (27, 18, 15) {real, imag} */,
  {32'h3ed9ea0d, 32'h3fdb0cc8} /* (27, 18, 14) {real, imag} */,
  {32'h3e8d1fcd, 32'h3e95c01e} /* (27, 18, 13) {real, imag} */,
  {32'h3d43a662, 32'h400a4167} /* (27, 18, 12) {real, imag} */,
  {32'h4014ce64, 32'h3f392ac0} /* (27, 18, 11) {real, imag} */,
  {32'hbfefd602, 32'hbf6c0f28} /* (27, 18, 10) {real, imag} */,
  {32'h3f3f994b, 32'hbff5d793} /* (27, 18, 9) {real, imag} */,
  {32'hbfac8f5b, 32'h3fd3bf51} /* (27, 18, 8) {real, imag} */,
  {32'hc03533a0, 32'h402e4ff3} /* (27, 18, 7) {real, imag} */,
  {32'hc01df9ee, 32'hbf7054c6} /* (27, 18, 6) {real, imag} */,
  {32'hc04774cf, 32'h3efb3592} /* (27, 18, 5) {real, imag} */,
  {32'hbf7c4ff5, 32'hbed16666} /* (27, 18, 4) {real, imag} */,
  {32'hbfc1e97b, 32'hbf937552} /* (27, 18, 3) {real, imag} */,
  {32'hbeb0cd0b, 32'hbef222e8} /* (27, 18, 2) {real, imag} */,
  {32'hbf942db1, 32'hbeb29ac0} /* (27, 18, 1) {real, imag} */,
  {32'h3f7647c4, 32'hbfbf52f9} /* (27, 18, 0) {real, imag} */,
  {32'h3fafb58e, 32'hbf11e280} /* (27, 17, 31) {real, imag} */,
  {32'hbf822b48, 32'h3f12f6ac} /* (27, 17, 30) {real, imag} */,
  {32'hbf28fd6b, 32'hbd43fc18} /* (27, 17, 29) {real, imag} */,
  {32'h3f3c26e5, 32'hbe748840} /* (27, 17, 28) {real, imag} */,
  {32'h3eb7008d, 32'hbf26e790} /* (27, 17, 27) {real, imag} */,
  {32'h3df30846, 32'h3f36a2cf} /* (27, 17, 26) {real, imag} */,
  {32'h3eedfe4a, 32'h3bb84b36} /* (27, 17, 25) {real, imag} */,
  {32'hc030d357, 32'hbd27467d} /* (27, 17, 24) {real, imag} */,
  {32'hbe9651e6, 32'hbe9468b6} /* (27, 17, 23) {real, imag} */,
  {32'h40340cf0, 32'h3ff90c07} /* (27, 17, 22) {real, imag} */,
  {32'h3edfe4c8, 32'hbf76ddc1} /* (27, 17, 21) {real, imag} */,
  {32'hbf0bf606, 32'hc03b39e3} /* (27, 17, 20) {real, imag} */,
  {32'h3f80c508, 32'hbfc231b9} /* (27, 17, 19) {real, imag} */,
  {32'h3e5c7b59, 32'hbfd90a45} /* (27, 17, 18) {real, imag} */,
  {32'h3f505a21, 32'hbf63f3a4} /* (27, 17, 17) {real, imag} */,
  {32'hbf9e2443, 32'hc016650c} /* (27, 17, 16) {real, imag} */,
  {32'h3fcddc9f, 32'h3fa6af97} /* (27, 17, 15) {real, imag} */,
  {32'hbfdc3959, 32'h3e0a7f8f} /* (27, 17, 14) {real, imag} */,
  {32'hc003eea9, 32'h3f7df29e} /* (27, 17, 13) {real, imag} */,
  {32'h3f29167c, 32'h3dc82eac} /* (27, 17, 12) {real, imag} */,
  {32'h3ea4cc4a, 32'h3ee74c0d} /* (27, 17, 11) {real, imag} */,
  {32'h3fbd5660, 32'hbfe17856} /* (27, 17, 10) {real, imag} */,
  {32'h3f7c5297, 32'hbe077448} /* (27, 17, 9) {real, imag} */,
  {32'hc026de24, 32'h3e81d4b1} /* (27, 17, 8) {real, imag} */,
  {32'hbfe0749c, 32'h3eea7c07} /* (27, 17, 7) {real, imag} */,
  {32'hbe72c29d, 32'hbf6386b5} /* (27, 17, 6) {real, imag} */,
  {32'hc00ef763, 32'hbf2d0dcc} /* (27, 17, 5) {real, imag} */,
  {32'hbee080a4, 32'h3f266e4a} /* (27, 17, 4) {real, imag} */,
  {32'h3c571ccc, 32'h3e714429} /* (27, 17, 3) {real, imag} */,
  {32'hbea57944, 32'hc05748c3} /* (27, 17, 2) {real, imag} */,
  {32'hbf1f4a4f, 32'h3efa6754} /* (27, 17, 1) {real, imag} */,
  {32'h402cafd7, 32'hc063f311} /* (27, 17, 0) {real, imag} */,
  {32'hbf747d8b, 32'hbf4fe89b} /* (27, 16, 31) {real, imag} */,
  {32'hbf6f8795, 32'h3f4f1682} /* (27, 16, 30) {real, imag} */,
  {32'hbe3f42da, 32'hbfb3e0e6} /* (27, 16, 29) {real, imag} */,
  {32'h3e9ac01c, 32'h3eb448d7} /* (27, 16, 28) {real, imag} */,
  {32'hbd803875, 32'hbe424207} /* (27, 16, 27) {real, imag} */,
  {32'hbf5220cb, 32'hbe3fec29} /* (27, 16, 26) {real, imag} */,
  {32'h3f462552, 32'hbf3540c3} /* (27, 16, 25) {real, imag} */,
  {32'h3f16d58e, 32'h3f2ecbed} /* (27, 16, 24) {real, imag} */,
  {32'h3fcdafa5, 32'hbff4bcbc} /* (27, 16, 23) {real, imag} */,
  {32'hbf0b72f7, 32'h3fb5b82f} /* (27, 16, 22) {real, imag} */,
  {32'h3fc5b3f1, 32'h3f88631c} /* (27, 16, 21) {real, imag} */,
  {32'h3f3354fa, 32'hbe1cb779} /* (27, 16, 20) {real, imag} */,
  {32'h3f74bb90, 32'hbebb313b} /* (27, 16, 19) {real, imag} */,
  {32'hbf378ce3, 32'hbfa0da6e} /* (27, 16, 18) {real, imag} */,
  {32'hbd0dc93a, 32'h3f7f4540} /* (27, 16, 17) {real, imag} */,
  {32'hbf55ca0a, 32'h3fda67d5} /* (27, 16, 16) {real, imag} */,
  {32'h3f11a220, 32'hbcbea816} /* (27, 16, 15) {real, imag} */,
  {32'h3ef7bf25, 32'hbee23ad0} /* (27, 16, 14) {real, imag} */,
  {32'hc02e8748, 32'h3e172af4} /* (27, 16, 13) {real, imag} */,
  {32'hc076b2ee, 32'hbf8a6c35} /* (27, 16, 12) {real, imag} */,
  {32'hbf70482f, 32'h3f7b03df} /* (27, 16, 11) {real, imag} */,
  {32'h3fa2d87b, 32'h3f9a2c78} /* (27, 16, 10) {real, imag} */,
  {32'hbd7b1d81, 32'hbdbc97da} /* (27, 16, 9) {real, imag} */,
  {32'hbe256b50, 32'hc03644ac} /* (27, 16, 8) {real, imag} */,
  {32'h3f0816e6, 32'h3e52b0a0} /* (27, 16, 7) {real, imag} */,
  {32'h3e523392, 32'h3dded9aa} /* (27, 16, 6) {real, imag} */,
  {32'h3d6d4a89, 32'hbf856c50} /* (27, 16, 5) {real, imag} */,
  {32'hbf421cd5, 32'hbfa42fbd} /* (27, 16, 4) {real, imag} */,
  {32'h3e3d0c71, 32'h3fa41233} /* (27, 16, 3) {real, imag} */,
  {32'h3881167f, 32'hbdf0ab10} /* (27, 16, 2) {real, imag} */,
  {32'h3d800434, 32'hbf18b804} /* (27, 16, 1) {real, imag} */,
  {32'h3f21364b, 32'hbb816a99} /* (27, 16, 0) {real, imag} */,
  {32'hc003050b, 32'hbe46e20e} /* (27, 15, 31) {real, imag} */,
  {32'hbe0dfde1, 32'hbf3f53df} /* (27, 15, 30) {real, imag} */,
  {32'hbf131738, 32'hbecee514} /* (27, 15, 29) {real, imag} */,
  {32'h3ea76196, 32'h3f3454c9} /* (27, 15, 28) {real, imag} */,
  {32'h3dc4fe2e, 32'hbe782fc5} /* (27, 15, 27) {real, imag} */,
  {32'hbe94ae1f, 32'hbfbd9c14} /* (27, 15, 26) {real, imag} */,
  {32'hbfc41e23, 32'h3f1bb780} /* (27, 15, 25) {real, imag} */,
  {32'h3c840ad9, 32'hbd8f1982} /* (27, 15, 24) {real, imag} */,
  {32'hbf91aa07, 32'h3f5efc56} /* (27, 15, 23) {real, imag} */,
  {32'hbfb0865f, 32'hbf79abde} /* (27, 15, 22) {real, imag} */,
  {32'h3f0ecb66, 32'hbdad275e} /* (27, 15, 21) {real, imag} */,
  {32'hbfa84386, 32'hbf133e6f} /* (27, 15, 20) {real, imag} */,
  {32'hbee89856, 32'hbfd10549} /* (27, 15, 19) {real, imag} */,
  {32'hc004ebae, 32'hc01bf860} /* (27, 15, 18) {real, imag} */,
  {32'h3e407555, 32'hbda0f4e5} /* (27, 15, 17) {real, imag} */,
  {32'h3fc65ea4, 32'h3f8f236f} /* (27, 15, 16) {real, imag} */,
  {32'hbeed27b9, 32'h3f076289} /* (27, 15, 15) {real, imag} */,
  {32'hbf3233b3, 32'hbc8fe803} /* (27, 15, 14) {real, imag} */,
  {32'h3f68ec5f, 32'h3d60ed97} /* (27, 15, 13) {real, imag} */,
  {32'hbdee3616, 32'hbf8a9baf} /* (27, 15, 12) {real, imag} */,
  {32'h3ea5ba1a, 32'h40270535} /* (27, 15, 11) {real, imag} */,
  {32'h3f84d324, 32'h3f464d45} /* (27, 15, 10) {real, imag} */,
  {32'hbf43dc07, 32'hbf80c5fd} /* (27, 15, 9) {real, imag} */,
  {32'h40098117, 32'h3f23d31e} /* (27, 15, 8) {real, imag} */,
  {32'hbfeb535f, 32'h3eeb29a9} /* (27, 15, 7) {real, imag} */,
  {32'hbfa46434, 32'hc010f8cc} /* (27, 15, 6) {real, imag} */,
  {32'h406e160c, 32'hbe381dbe} /* (27, 15, 5) {real, imag} */,
  {32'hbfae0b34, 32'hbf69fc8b} /* (27, 15, 4) {real, imag} */,
  {32'h3ee99e9c, 32'hbdb37548} /* (27, 15, 3) {real, imag} */,
  {32'hbf0f7d1d, 32'h3fbdce1a} /* (27, 15, 2) {real, imag} */,
  {32'hbd8a66e3, 32'h40031d5c} /* (27, 15, 1) {real, imag} */,
  {32'h3cfd026f, 32'h3ed856f7} /* (27, 15, 0) {real, imag} */,
  {32'hbd2446c6, 32'hc04b67f8} /* (27, 14, 31) {real, imag} */,
  {32'hbf68fffc, 32'h3fd0de96} /* (27, 14, 30) {real, imag} */,
  {32'h3f1ffd36, 32'h3f3793bf} /* (27, 14, 29) {real, imag} */,
  {32'hbf4cbbcf, 32'h405017fb} /* (27, 14, 28) {real, imag} */,
  {32'hbefd831f, 32'h3e4bf915} /* (27, 14, 27) {real, imag} */,
  {32'h401778ad, 32'h4029776e} /* (27, 14, 26) {real, imag} */,
  {32'hc02d2c78, 32'h3f8b4d74} /* (27, 14, 25) {real, imag} */,
  {32'hbfc8f6ff, 32'hc007fae2} /* (27, 14, 24) {real, imag} */,
  {32'h3f40d98f, 32'hbf2bcfd2} /* (27, 14, 23) {real, imag} */,
  {32'h3f718fe8, 32'hc06fe94e} /* (27, 14, 22) {real, imag} */,
  {32'h3fa5b91f, 32'h3ca42698} /* (27, 14, 21) {real, imag} */,
  {32'h3f35441c, 32'h403e1220} /* (27, 14, 20) {real, imag} */,
  {32'h3f9392ec, 32'h3fb8035a} /* (27, 14, 19) {real, imag} */,
  {32'hbfa15d40, 32'h3f05c707} /* (27, 14, 18) {real, imag} */,
  {32'h3f26bb51, 32'hbf55f0e5} /* (27, 14, 17) {real, imag} */,
  {32'hbf13dc09, 32'h3e5093b3} /* (27, 14, 16) {real, imag} */,
  {32'h3fa3687b, 32'h40096edf} /* (27, 14, 15) {real, imag} */,
  {32'hbf034b87, 32'hbee92175} /* (27, 14, 14) {real, imag} */,
  {32'h3fb11e7b, 32'hbf2f909e} /* (27, 14, 13) {real, imag} */,
  {32'h3f6433ed, 32'h40680cc3} /* (27, 14, 12) {real, imag} */,
  {32'h3fd95279, 32'hbf583309} /* (27, 14, 11) {real, imag} */,
  {32'h4085aabf, 32'h401ebd1f} /* (27, 14, 10) {real, imag} */,
  {32'hc02a7f1f, 32'hbf4637e7} /* (27, 14, 9) {real, imag} */,
  {32'hbf1df981, 32'hbd2b3a26} /* (27, 14, 8) {real, imag} */,
  {32'h3f895c5d, 32'h3edb605d} /* (27, 14, 7) {real, imag} */,
  {32'h3ef94f67, 32'hbeeac5e3} /* (27, 14, 6) {real, imag} */,
  {32'h3fdf4870, 32'h3c11d1b2} /* (27, 14, 5) {real, imag} */,
  {32'hbeff8478, 32'h3f1f2e1b} /* (27, 14, 4) {real, imag} */,
  {32'h3fa1b1ca, 32'h404ed7bb} /* (27, 14, 3) {real, imag} */,
  {32'h3c630062, 32'hc06216cb} /* (27, 14, 2) {real, imag} */,
  {32'hbec1d39b, 32'h3f677abd} /* (27, 14, 1) {real, imag} */,
  {32'h3e9abafa, 32'hbf8bce1e} /* (27, 14, 0) {real, imag} */,
  {32'h3fc53417, 32'h3f2eddc6} /* (27, 13, 31) {real, imag} */,
  {32'h3f0de3d6, 32'h3f339c2d} /* (27, 13, 30) {real, imag} */,
  {32'hbff8d255, 32'hbe403044} /* (27, 13, 29) {real, imag} */,
  {32'h403c642f, 32'hbebac3d7} /* (27, 13, 28) {real, imag} */,
  {32'hc08cfcd4, 32'h3f51fe2d} /* (27, 13, 27) {real, imag} */,
  {32'h3ee30f62, 32'h3e317e98} /* (27, 13, 26) {real, imag} */,
  {32'hbf4d9e14, 32'hbfa1cf32} /* (27, 13, 25) {real, imag} */,
  {32'hc0199763, 32'h3f612b74} /* (27, 13, 24) {real, imag} */,
  {32'hbfff00f3, 32'hc0004707} /* (27, 13, 23) {real, imag} */,
  {32'h402d6d13, 32'h3faffebe} /* (27, 13, 22) {real, imag} */,
  {32'hc006e756, 32'hbe9a4d89} /* (27, 13, 21) {real, imag} */,
  {32'hbec45608, 32'hbff36cea} /* (27, 13, 20) {real, imag} */,
  {32'h3f0df1be, 32'hc0279810} /* (27, 13, 19) {real, imag} */,
  {32'h3eebf40d, 32'hbfc430e3} /* (27, 13, 18) {real, imag} */,
  {32'hbfc6592c, 32'h3f691dc9} /* (27, 13, 17) {real, imag} */,
  {32'h3ff6ca54, 32'h3f84d977} /* (27, 13, 16) {real, imag} */,
  {32'hbf0fb343, 32'hc006bcbf} /* (27, 13, 15) {real, imag} */,
  {32'hbfb04eb0, 32'hbedfe41b} /* (27, 13, 14) {real, imag} */,
  {32'h3f00d326, 32'hbfa659fa} /* (27, 13, 13) {real, imag} */,
  {32'hbeeb3d57, 32'h3e8a1290} /* (27, 13, 12) {real, imag} */,
  {32'h40336db6, 32'h40010629} /* (27, 13, 11) {real, imag} */,
  {32'h3f565a8a, 32'hbf4a1cd5} /* (27, 13, 10) {real, imag} */,
  {32'h3fa88a6d, 32'h40434a5f} /* (27, 13, 9) {real, imag} */,
  {32'h3ef36f94, 32'h3d4cb3f6} /* (27, 13, 8) {real, imag} */,
  {32'h40457e48, 32'h4024bd87} /* (27, 13, 7) {real, imag} */,
  {32'hbfd699b0, 32'hbf8ff6ec} /* (27, 13, 6) {real, imag} */,
  {32'h3fd84010, 32'h3fa13fca} /* (27, 13, 5) {real, imag} */,
  {32'hbfe34d10, 32'h3ed0cf67} /* (27, 13, 4) {real, imag} */,
  {32'hbfc477c0, 32'h3f8da572} /* (27, 13, 3) {real, imag} */,
  {32'h3f5355ca, 32'hbfb5206e} /* (27, 13, 2) {real, imag} */,
  {32'hbec99177, 32'h3e987a26} /* (27, 13, 1) {real, imag} */,
  {32'hc00233ee, 32'h3e154b6e} /* (27, 13, 0) {real, imag} */,
  {32'h3f6cb9fd, 32'h3ff0a08c} /* (27, 12, 31) {real, imag} */,
  {32'hbe61dbdd, 32'hbe8b2bee} /* (27, 12, 30) {real, imag} */,
  {32'h3fed27ef, 32'hbf8c739c} /* (27, 12, 29) {real, imag} */,
  {32'hc073cf27, 32'hc030c764} /* (27, 12, 28) {real, imag} */,
  {32'hbf766380, 32'h3ff1e2fe} /* (27, 12, 27) {real, imag} */,
  {32'h4018846c, 32'hbf4a4877} /* (27, 12, 26) {real, imag} */,
  {32'h3ee6b39a, 32'h40647faf} /* (27, 12, 25) {real, imag} */,
  {32'hbed49f0a, 32'hbf0a6c4b} /* (27, 12, 24) {real, imag} */,
  {32'h40566376, 32'h3fb33bdb} /* (27, 12, 23) {real, imag} */,
  {32'hbfa5fc4a, 32'h3fb93d80} /* (27, 12, 22) {real, imag} */,
  {32'h3fde74b9, 32'h3ff76a7d} /* (27, 12, 21) {real, imag} */,
  {32'h3e8308d4, 32'hbcda7e9c} /* (27, 12, 20) {real, imag} */,
  {32'hc017ba11, 32'h3f0c9d01} /* (27, 12, 19) {real, imag} */,
  {32'hc0102707, 32'hbf6ee016} /* (27, 12, 18) {real, imag} */,
  {32'hbfbc7b50, 32'h3fa8037f} /* (27, 12, 17) {real, imag} */,
  {32'h3f1e630f, 32'hbf78794e} /* (27, 12, 16) {real, imag} */,
  {32'h3f072c7e, 32'h3f3208a8} /* (27, 12, 15) {real, imag} */,
  {32'hbeb3db66, 32'hbf188428} /* (27, 12, 14) {real, imag} */,
  {32'hbf9a1caa, 32'h3e8e85bd} /* (27, 12, 13) {real, imag} */,
  {32'h3f99093f, 32'hc046d039} /* (27, 12, 12) {real, imag} */,
  {32'hbecbf366, 32'h3f8c0ae2} /* (27, 12, 11) {real, imag} */,
  {32'h3f5b9abb, 32'h40441966} /* (27, 12, 10) {real, imag} */,
  {32'hbf64a03b, 32'h402d76cb} /* (27, 12, 9) {real, imag} */,
  {32'h3f8ba5a8, 32'hbf24c5f9} /* (27, 12, 8) {real, imag} */,
  {32'h3c96aae1, 32'hbe7cc52b} /* (27, 12, 7) {real, imag} */,
  {32'hc043896a, 32'hbb1057d2} /* (27, 12, 6) {real, imag} */,
  {32'hc031db2d, 32'h4016cefd} /* (27, 12, 5) {real, imag} */,
  {32'h4011dacd, 32'h3fc7fb4b} /* (27, 12, 4) {real, imag} */,
  {32'hbf771c42, 32'hbf047229} /* (27, 12, 3) {real, imag} */,
  {32'h3f017388, 32'h3fb20dcf} /* (27, 12, 2) {real, imag} */,
  {32'h3fec3568, 32'h3fede6dc} /* (27, 12, 1) {real, imag} */,
  {32'h3fffa6b6, 32'h3f83da9b} /* (27, 12, 0) {real, imag} */,
  {32'hbd4f2ca0, 32'hc04d1ce8} /* (27, 11, 31) {real, imag} */,
  {32'hbf04d3d9, 32'hbf9805c1} /* (27, 11, 30) {real, imag} */,
  {32'h3f60776d, 32'hbeb71427} /* (27, 11, 29) {real, imag} */,
  {32'hbfa41bf3, 32'hc0249dd5} /* (27, 11, 28) {real, imag} */,
  {32'hbf8e103d, 32'h4084e02b} /* (27, 11, 27) {real, imag} */,
  {32'hbe125a4e, 32'h3f4e80b6} /* (27, 11, 26) {real, imag} */,
  {32'h3d16777c, 32'hc091ea22} /* (27, 11, 25) {real, imag} */,
  {32'hbd925911, 32'h4007e676} /* (27, 11, 24) {real, imag} */,
  {32'h3f835bf0, 32'h3fe13111} /* (27, 11, 23) {real, imag} */,
  {32'hbf32661f, 32'h3eeebbfe} /* (27, 11, 22) {real, imag} */,
  {32'h3f808ba7, 32'h3feee766} /* (27, 11, 21) {real, imag} */,
  {32'h3ef47941, 32'h3e1503a8} /* (27, 11, 20) {real, imag} */,
  {32'h40374aab, 32'hbfe0200a} /* (27, 11, 19) {real, imag} */,
  {32'h404361ca, 32'h3fa56707} /* (27, 11, 18) {real, imag} */,
  {32'hbf90a454, 32'hbd12eea5} /* (27, 11, 17) {real, imag} */,
  {32'hbe0aaa25, 32'hc01cb5e9} /* (27, 11, 16) {real, imag} */,
  {32'hbf38874f, 32'h40132243} /* (27, 11, 15) {real, imag} */,
  {32'hbf893eeb, 32'h400b5439} /* (27, 11, 14) {real, imag} */,
  {32'hbf9c5260, 32'hc02e9ae5} /* (27, 11, 13) {real, imag} */,
  {32'hc0180ddc, 32'h3e628dcc} /* (27, 11, 12) {real, imag} */,
  {32'h3ef763fd, 32'hc023d47a} /* (27, 11, 11) {real, imag} */,
  {32'hc0535fce, 32'hc055ea4f} /* (27, 11, 10) {real, imag} */,
  {32'h3ebf331c, 32'hc0301d27} /* (27, 11, 9) {real, imag} */,
  {32'hbf80ac3a, 32'h3ed259d9} /* (27, 11, 8) {real, imag} */,
  {32'h3f1f8b64, 32'hbdcb4795} /* (27, 11, 7) {real, imag} */,
  {32'h3f64ccad, 32'h3cf147bb} /* (27, 11, 6) {real, imag} */,
  {32'hc009222b, 32'hbf284b67} /* (27, 11, 5) {real, imag} */,
  {32'h409ea013, 32'hbf00c09f} /* (27, 11, 4) {real, imag} */,
  {32'h3f8bc9ee, 32'hbfa7b1ca} /* (27, 11, 3) {real, imag} */,
  {32'hbf8e85de, 32'hbfda826f} /* (27, 11, 2) {real, imag} */,
  {32'h3fab1855, 32'hbdea4e0c} /* (27, 11, 1) {real, imag} */,
  {32'h3f8239f4, 32'hc065110e} /* (27, 11, 0) {real, imag} */,
  {32'hc046147a, 32'h3fd58e0a} /* (27, 10, 31) {real, imag} */,
  {32'hbe2e4f19, 32'hbfbfe55a} /* (27, 10, 30) {real, imag} */,
  {32'hbfdf3c7b, 32'hbf299875} /* (27, 10, 29) {real, imag} */,
  {32'h3fd9b4ae, 32'hbfb12229} /* (27, 10, 28) {real, imag} */,
  {32'h40291ab7, 32'hbf300d66} /* (27, 10, 27) {real, imag} */,
  {32'hbfb0461a, 32'hbe36d040} /* (27, 10, 26) {real, imag} */,
  {32'h3fbf170e, 32'hc022114a} /* (27, 10, 25) {real, imag} */,
  {32'hc002424f, 32'h3f636df5} /* (27, 10, 24) {real, imag} */,
  {32'hbf759a5e, 32'h40093e0c} /* (27, 10, 23) {real, imag} */,
  {32'h40346a3f, 32'hc006702d} /* (27, 10, 22) {real, imag} */,
  {32'hbe349673, 32'h403b1da1} /* (27, 10, 21) {real, imag} */,
  {32'h3f7530c5, 32'h3f7f6d4b} /* (27, 10, 20) {real, imag} */,
  {32'h3e21e46c, 32'h3f9feadb} /* (27, 10, 19) {real, imag} */,
  {32'hbea7dff0, 32'hbedfcad1} /* (27, 10, 18) {real, imag} */,
  {32'h3f943218, 32'hc03f2a7e} /* (27, 10, 17) {real, imag} */,
  {32'hbe0ac5f7, 32'h3ee5adf6} /* (27, 10, 16) {real, imag} */,
  {32'h3c54781e, 32'h3fb38557} /* (27, 10, 15) {real, imag} */,
  {32'h3f306f3a, 32'h3ea2eab7} /* (27, 10, 14) {real, imag} */,
  {32'h3ff82404, 32'hbf1c13a9} /* (27, 10, 13) {real, imag} */,
  {32'hc06d6841, 32'hbf3c72b5} /* (27, 10, 12) {real, imag} */,
  {32'h40018e37, 32'hbfa66817} /* (27, 10, 11) {real, imag} */,
  {32'hbe7cd5b5, 32'h3eeaf798} /* (27, 10, 10) {real, imag} */,
  {32'h3f0fac16, 32'h3dcb4e38} /* (27, 10, 9) {real, imag} */,
  {32'hbf179172, 32'hc013f253} /* (27, 10, 8) {real, imag} */,
  {32'h40826f7e, 32'h3fee9773} /* (27, 10, 7) {real, imag} */,
  {32'hc05314f3, 32'hbf2a4d29} /* (27, 10, 6) {real, imag} */,
  {32'h3f6e1fc0, 32'hbf3c50cf} /* (27, 10, 5) {real, imag} */,
  {32'hbf45891e, 32'h400b2fa3} /* (27, 10, 4) {real, imag} */,
  {32'hc04f1fe4, 32'h407ebaca} /* (27, 10, 3) {real, imag} */,
  {32'hc045f8eb, 32'hc04bb80e} /* (27, 10, 2) {real, imag} */,
  {32'h4070e1c2, 32'h4041a511} /* (27, 10, 1) {real, imag} */,
  {32'hbff015df, 32'h40268bc1} /* (27, 10, 0) {real, imag} */,
  {32'hbfe24110, 32'h4002e75b} /* (27, 9, 31) {real, imag} */,
  {32'h3fc644ec, 32'h40553d71} /* (27, 9, 30) {real, imag} */,
  {32'h401c687a, 32'h3e41c2a0} /* (27, 9, 29) {real, imag} */,
  {32'hc0032d92, 32'hc078ea99} /* (27, 9, 28) {real, imag} */,
  {32'hbf202c70, 32'hc053a9a6} /* (27, 9, 27) {real, imag} */,
  {32'hc05027b7, 32'hc08230ce} /* (27, 9, 26) {real, imag} */,
  {32'h4017a41c, 32'h400bda81} /* (27, 9, 25) {real, imag} */,
  {32'h3f942f7e, 32'hc00020de} /* (27, 9, 24) {real, imag} */,
  {32'h4028d329, 32'h3fc651ea} /* (27, 9, 23) {real, imag} */,
  {32'h3f502d83, 32'h3e8563ee} /* (27, 9, 22) {real, imag} */,
  {32'hc0453144, 32'hbffeb768} /* (27, 9, 21) {real, imag} */,
  {32'h3f9cb88f, 32'h3f088a0c} /* (27, 9, 20) {real, imag} */,
  {32'h3f705267, 32'h3fa00a1e} /* (27, 9, 19) {real, imag} */,
  {32'hbf44332c, 32'hbf266de2} /* (27, 9, 18) {real, imag} */,
  {32'h40905394, 32'h3f85a276} /* (27, 9, 17) {real, imag} */,
  {32'hc09056ce, 32'h3f6b4aa8} /* (27, 9, 16) {real, imag} */,
  {32'hbf062c23, 32'hbff8cc56} /* (27, 9, 15) {real, imag} */,
  {32'h3fe0369c, 32'hbf3911ef} /* (27, 9, 14) {real, imag} */,
  {32'h401193df, 32'h3f92e5af} /* (27, 9, 13) {real, imag} */,
  {32'hbfcc486b, 32'h3eeae6ae} /* (27, 9, 12) {real, imag} */,
  {32'hbec6535d, 32'h408a14b7} /* (27, 9, 11) {real, imag} */,
  {32'hbe406c9c, 32'hbf6f3394} /* (27, 9, 10) {real, imag} */,
  {32'hbfaa981b, 32'h4016483c} /* (27, 9, 9) {real, imag} */,
  {32'hbfb44cd8, 32'hbf471c6b} /* (27, 9, 8) {real, imag} */,
  {32'hbfd85180, 32'hbf77d8d2} /* (27, 9, 7) {real, imag} */,
  {32'h3f44b2fa, 32'hbffdaa94} /* (27, 9, 6) {real, imag} */,
  {32'h40882a84, 32'h4030df36} /* (27, 9, 5) {real, imag} */,
  {32'hc04b0959, 32'h3ee3ad60} /* (27, 9, 4) {real, imag} */,
  {32'hbf23b245, 32'hc083808a} /* (27, 9, 3) {real, imag} */,
  {32'hbf532417, 32'h401bdff9} /* (27, 9, 2) {real, imag} */,
  {32'h3ec7d51a, 32'hbcdd3235} /* (27, 9, 1) {real, imag} */,
  {32'hbf16f9e4, 32'h3f181959} /* (27, 9, 0) {real, imag} */,
  {32'h3fb3496f, 32'hc0e3aac5} /* (27, 8, 31) {real, imag} */,
  {32'hbf4f1e09, 32'h40474cc4} /* (27, 8, 30) {real, imag} */,
  {32'h40abb0cd, 32'h3f78abd3} /* (27, 8, 29) {real, imag} */,
  {32'hc04e51e0, 32'h402ad5c7} /* (27, 8, 28) {real, imag} */,
  {32'h408564d6, 32'hbf84a23e} /* (27, 8, 27) {real, imag} */,
  {32'hbf1d3044, 32'h3ff8701f} /* (27, 8, 26) {real, imag} */,
  {32'hbe7d66ea, 32'hbfb5af90} /* (27, 8, 25) {real, imag} */,
  {32'h409b4674, 32'h402d7a92} /* (27, 8, 24) {real, imag} */,
  {32'h40125a82, 32'h3f455dc4} /* (27, 8, 23) {real, imag} */,
  {32'hbeca444a, 32'h3fbb2755} /* (27, 8, 22) {real, imag} */,
  {32'hbda298e0, 32'hbf2ff646} /* (27, 8, 21) {real, imag} */,
  {32'hc01ff298, 32'hbfa3cac9} /* (27, 8, 20) {real, imag} */,
  {32'h3fa1e5d6, 32'h3f9f3a02} /* (27, 8, 19) {real, imag} */,
  {32'hbf0c2630, 32'hbf3c2ac0} /* (27, 8, 18) {real, imag} */,
  {32'hbf9441cb, 32'h3ed41270} /* (27, 8, 17) {real, imag} */,
  {32'hbfd6e331, 32'h3e510f03} /* (27, 8, 16) {real, imag} */,
  {32'h40039008, 32'hbf328b9a} /* (27, 8, 15) {real, imag} */,
  {32'hbe235597, 32'hbf0132f4} /* (27, 8, 14) {real, imag} */,
  {32'h3f306094, 32'hbf37a66b} /* (27, 8, 13) {real, imag} */,
  {32'h4011a9e5, 32'hc0054996} /* (27, 8, 12) {real, imag} */,
  {32'h40a48e5a, 32'h3fa562e8} /* (27, 8, 11) {real, imag} */,
  {32'hc08487ff, 32'hc06251f1} /* (27, 8, 10) {real, imag} */,
  {32'hbfd5a14b, 32'hbfe75ba6} /* (27, 8, 9) {real, imag} */,
  {32'hbfce4d9f, 32'h3f787213} /* (27, 8, 8) {real, imag} */,
  {32'hc0380f4a, 32'h3d25b993} /* (27, 8, 7) {real, imag} */,
  {32'h404b2687, 32'hc052268c} /* (27, 8, 6) {real, imag} */,
  {32'hbf9a6e9e, 32'hbf31b8a3} /* (27, 8, 5) {real, imag} */,
  {32'hc0154ed6, 32'hbf7d92c0} /* (27, 8, 4) {real, imag} */,
  {32'hc02440a0, 32'h4058e83f} /* (27, 8, 3) {real, imag} */,
  {32'h3fe11007, 32'h40067ed2} /* (27, 8, 2) {real, imag} */,
  {32'hbe788339, 32'hbe67282a} /* (27, 8, 1) {real, imag} */,
  {32'h3ef4ce51, 32'hc07c5a6d} /* (27, 8, 0) {real, imag} */,
  {32'h3eeed053, 32'hc03c1047} /* (27, 7, 31) {real, imag} */,
  {32'h40ad7551, 32'hbf05d6b1} /* (27, 7, 30) {real, imag} */,
  {32'h4018f901, 32'hc017b318} /* (27, 7, 29) {real, imag} */,
  {32'hbf3e9330, 32'h4021d07b} /* (27, 7, 28) {real, imag} */,
  {32'hbbb0cb30, 32'hc006984c} /* (27, 7, 27) {real, imag} */,
  {32'hc0053779, 32'hbe882c43} /* (27, 7, 26) {real, imag} */,
  {32'hc0214c0c, 32'hbf5e018f} /* (27, 7, 25) {real, imag} */,
  {32'h404d0c11, 32'hbf73713d} /* (27, 7, 24) {real, imag} */,
  {32'h3f5c08a1, 32'hbfb952a5} /* (27, 7, 23) {real, imag} */,
  {32'hbee8f595, 32'h3faf993a} /* (27, 7, 22) {real, imag} */,
  {32'h40119f08, 32'hc0548cba} /* (27, 7, 21) {real, imag} */,
  {32'h400b12c9, 32'h400a363e} /* (27, 7, 20) {real, imag} */,
  {32'hbfa8aa49, 32'h4041f33f} /* (27, 7, 19) {real, imag} */,
  {32'h3e6a62ff, 32'hbc698fbc} /* (27, 7, 18) {real, imag} */,
  {32'h3d4c65fa, 32'h401656d2} /* (27, 7, 17) {real, imag} */,
  {32'hc05751a2, 32'h3dfdc26e} /* (27, 7, 16) {real, imag} */,
  {32'h3fb60222, 32'h3ff66af9} /* (27, 7, 15) {real, imag} */,
  {32'h3fe1e8fe, 32'h3fa42c9b} /* (27, 7, 14) {real, imag} */,
  {32'h3fafde29, 32'h3e4b4162} /* (27, 7, 13) {real, imag} */,
  {32'h3fd7be94, 32'hbfb70916} /* (27, 7, 12) {real, imag} */,
  {32'hbf2ab465, 32'hc01de006} /* (27, 7, 11) {real, imag} */,
  {32'hbf3bc1c1, 32'hbd075f86} /* (27, 7, 10) {real, imag} */,
  {32'h3bd5b41d, 32'hbe8c52b9} /* (27, 7, 9) {real, imag} */,
  {32'h3fa3b06d, 32'hbf9bd9e7} /* (27, 7, 8) {real, imag} */,
  {32'hc0169c4f, 32'hbe07855a} /* (27, 7, 7) {real, imag} */,
  {32'hbfae8b6e, 32'hbed81cad} /* (27, 7, 6) {real, imag} */,
  {32'h3f2f0650, 32'h40083c63} /* (27, 7, 5) {real, imag} */,
  {32'h3fd34ece, 32'hc0006f9f} /* (27, 7, 4) {real, imag} */,
  {32'h3fed553e, 32'h4029dcf3} /* (27, 7, 3) {real, imag} */,
  {32'h40a3b2ba, 32'hc04ef264} /* (27, 7, 2) {real, imag} */,
  {32'hbfc4b3da, 32'h4086646e} /* (27, 7, 1) {real, imag} */,
  {32'hc0020a27, 32'h4080b46c} /* (27, 7, 0) {real, imag} */,
  {32'hc0bb4b55, 32'hc081f36d} /* (27, 6, 31) {real, imag} */,
  {32'hc02e3f92, 32'h3f2342c0} /* (27, 6, 30) {real, imag} */,
  {32'hc096f727, 32'hbedb3d77} /* (27, 6, 29) {real, imag} */,
  {32'h4026d152, 32'hbe8d984f} /* (27, 6, 28) {real, imag} */,
  {32'h40ddab85, 32'h3f52dc1c} /* (27, 6, 27) {real, imag} */,
  {32'h40437847, 32'h4025f2d6} /* (27, 6, 26) {real, imag} */,
  {32'h3fd94627, 32'hc081368e} /* (27, 6, 25) {real, imag} */,
  {32'hbf81ccc7, 32'hbf82fd5b} /* (27, 6, 24) {real, imag} */,
  {32'hbff40f35, 32'h3da50418} /* (27, 6, 23) {real, imag} */,
  {32'h40846292, 32'h3f8e5ae1} /* (27, 6, 22) {real, imag} */,
  {32'hbf91532d, 32'h3decd91e} /* (27, 6, 21) {real, imag} */,
  {32'h3f8e30b4, 32'hbe9ca189} /* (27, 6, 20) {real, imag} */,
  {32'h3f8cf68e, 32'hbf89c0ae} /* (27, 6, 19) {real, imag} */,
  {32'hbed9f72d, 32'hbf52516b} /* (27, 6, 18) {real, imag} */,
  {32'hbfb75c59, 32'hbfd77077} /* (27, 6, 17) {real, imag} */,
  {32'h3f19bf7c, 32'hbf20c466} /* (27, 6, 16) {real, imag} */,
  {32'h3fd9cd71, 32'h3fdfab86} /* (27, 6, 15) {real, imag} */,
  {32'hbf6d01c5, 32'hc04d98aa} /* (27, 6, 14) {real, imag} */,
  {32'h3d4d75b2, 32'hbf68b209} /* (27, 6, 13) {real, imag} */,
  {32'hc01845d5, 32'hbf899229} /* (27, 6, 12) {real, imag} */,
  {32'h401f3757, 32'h3fbe0315} /* (27, 6, 11) {real, imag} */,
  {32'hbe93be9a, 32'h3f5afcac} /* (27, 6, 10) {real, imag} */,
  {32'hc0882f43, 32'h3e1a63f7} /* (27, 6, 9) {real, imag} */,
  {32'h405607b1, 32'h40ac1ec9} /* (27, 6, 8) {real, imag} */,
  {32'hbf983560, 32'hc0245e4e} /* (27, 6, 7) {real, imag} */,
  {32'h3faba6b1, 32'hc0618351} /* (27, 6, 6) {real, imag} */,
  {32'h3f46fcec, 32'hc082aee8} /* (27, 6, 5) {real, imag} */,
  {32'hbfad30ee, 32'hbfd4e0b6} /* (27, 6, 4) {real, imag} */,
  {32'h3fcb9bf1, 32'h3fd1e184} /* (27, 6, 3) {real, imag} */,
  {32'h3f2015d5, 32'h3cb9a8cd} /* (27, 6, 2) {real, imag} */,
  {32'hc0a71829, 32'hbfe58fd8} /* (27, 6, 1) {real, imag} */,
  {32'h3f9b8565, 32'hc0b65cb7} /* (27, 6, 0) {real, imag} */,
  {32'h402e0763, 32'hc0e47694} /* (27, 5, 31) {real, imag} */,
  {32'h40e04304, 32'h40caa814} /* (27, 5, 30) {real, imag} */,
  {32'hc09e9e35, 32'h408b27d3} /* (27, 5, 29) {real, imag} */,
  {32'hbec4796c, 32'h4006750a} /* (27, 5, 28) {real, imag} */,
  {32'h40a64ae3, 32'hbf645568} /* (27, 5, 27) {real, imag} */,
  {32'h3fbd669f, 32'hc0017847} /* (27, 5, 26) {real, imag} */,
  {32'hbef1bdb8, 32'hc03f7d86} /* (27, 5, 25) {real, imag} */,
  {32'hbf6bb8d8, 32'hbe0c72fc} /* (27, 5, 24) {real, imag} */,
  {32'hc0221747, 32'h3f967fd6} /* (27, 5, 23) {real, imag} */,
  {32'h3f38dd2c, 32'h3ea246a1} /* (27, 5, 22) {real, imag} */,
  {32'h3ecd6be8, 32'h3f0888ac} /* (27, 5, 21) {real, imag} */,
  {32'h3fe3e395, 32'hbf530f71} /* (27, 5, 20) {real, imag} */,
  {32'h3f4ae9e3, 32'hbecbe975} /* (27, 5, 19) {real, imag} */,
  {32'h3fc87c99, 32'h3ff4d531} /* (27, 5, 18) {real, imag} */,
  {32'h3f627bb8, 32'h3f154524} /* (27, 5, 17) {real, imag} */,
  {32'h3fc2b545, 32'hbf8274f3} /* (27, 5, 16) {real, imag} */,
  {32'hbf9815e2, 32'hbd3c0c47} /* (27, 5, 15) {real, imag} */,
  {32'hc002687f, 32'hbe81e47a} /* (27, 5, 14) {real, imag} */,
  {32'h3e5dffe2, 32'h3fe6923d} /* (27, 5, 13) {real, imag} */,
  {32'h40265e21, 32'hc063ac2b} /* (27, 5, 12) {real, imag} */,
  {32'h3f01d9ad, 32'h3aa9764a} /* (27, 5, 11) {real, imag} */,
  {32'h40028719, 32'h404b8737} /* (27, 5, 10) {real, imag} */,
  {32'h3f8d666e, 32'h3fc54d96} /* (27, 5, 9) {real, imag} */,
  {32'hbf11f288, 32'hc06e393d} /* (27, 5, 8) {real, imag} */,
  {32'h3fdaf5f4, 32'hc0001acf} /* (27, 5, 7) {real, imag} */,
  {32'hbf075d88, 32'h408f49a9} /* (27, 5, 6) {real, imag} */,
  {32'h400f7287, 32'h4064ae49} /* (27, 5, 5) {real, imag} */,
  {32'h3ea3e1e5, 32'hbf306ac2} /* (27, 5, 4) {real, imag} */,
  {32'h3fb4ad8d, 32'hbf4e50af} /* (27, 5, 3) {real, imag} */,
  {32'hbf90a631, 32'h4023b676} /* (27, 5, 2) {real, imag} */,
  {32'hc11ac09a, 32'hc0fc55fb} /* (27, 5, 1) {real, imag} */,
  {32'hc09603b5, 32'hc02a6ebb} /* (27, 5, 0) {real, imag} */,
  {32'hc107038a, 32'h409d7308} /* (27, 4, 31) {real, imag} */,
  {32'h408fa855, 32'hc09a1b25} /* (27, 4, 30) {real, imag} */,
  {32'h3f8742c5, 32'hc097b284} /* (27, 4, 29) {real, imag} */,
  {32'hc0200b31, 32'h40c356a9} /* (27, 4, 28) {real, imag} */,
  {32'hbf00df38, 32'hbfdcec75} /* (27, 4, 27) {real, imag} */,
  {32'hc01add25, 32'hc02bb02e} /* (27, 4, 26) {real, imag} */,
  {32'h3f3acb9e, 32'h4030dfde} /* (27, 4, 25) {real, imag} */,
  {32'hc0469bcb, 32'hc0386780} /* (27, 4, 24) {real, imag} */,
  {32'hbf60b185, 32'hc0376772} /* (27, 4, 23) {real, imag} */,
  {32'h40459902, 32'h3fd1c407} /* (27, 4, 22) {real, imag} */,
  {32'h3d5de636, 32'h3e9f9b6d} /* (27, 4, 21) {real, imag} */,
  {32'hbfb824da, 32'hbf5900cf} /* (27, 4, 20) {real, imag} */,
  {32'hbf1b8849, 32'hc004eb2a} /* (27, 4, 19) {real, imag} */,
  {32'hbf6df517, 32'h3f1c8534} /* (27, 4, 18) {real, imag} */,
  {32'h4008ceb7, 32'hbd1ecb70} /* (27, 4, 17) {real, imag} */,
  {32'h3f2e4e5d, 32'h3fec6afd} /* (27, 4, 16) {real, imag} */,
  {32'hbf586f08, 32'hbff66f32} /* (27, 4, 15) {real, imag} */,
  {32'hbedf2730, 32'hc0387066} /* (27, 4, 14) {real, imag} */,
  {32'h3f4fb661, 32'h3d790902} /* (27, 4, 13) {real, imag} */,
  {32'h3d58b60f, 32'h3f949e16} /* (27, 4, 12) {real, imag} */,
  {32'hbfd88994, 32'h3f9e343f} /* (27, 4, 11) {real, imag} */,
  {32'hc0277fba, 32'hbd9492cd} /* (27, 4, 10) {real, imag} */,
  {32'h4020881a, 32'h3fb9f7c4} /* (27, 4, 9) {real, imag} */,
  {32'h3f09d70c, 32'h3f894a95} /* (27, 4, 8) {real, imag} */,
  {32'h3f588417, 32'hbd366576} /* (27, 4, 7) {real, imag} */,
  {32'h3f217938, 32'h40b5d367} /* (27, 4, 6) {real, imag} */,
  {32'h400c33ef, 32'hc00a9010} /* (27, 4, 5) {real, imag} */,
  {32'hbe6709e5, 32'h3fc4be96} /* (27, 4, 4) {real, imag} */,
  {32'hbfefce2f, 32'hc0691709} /* (27, 4, 3) {real, imag} */,
  {32'hc0b2ce47, 32'hc10f0c40} /* (27, 4, 2) {real, imag} */,
  {32'hbdd0dbce, 32'h4148be4f} /* (27, 4, 1) {real, imag} */,
  {32'h4033948a, 32'hc0bef1c9} /* (27, 4, 0) {real, imag} */,
  {32'hc166aef6, 32'hc0414338} /* (27, 3, 31) {real, imag} */,
  {32'h4125b26e, 32'h40a16882} /* (27, 3, 30) {real, imag} */,
  {32'h40408634, 32'hbfc1ad07} /* (27, 3, 29) {real, imag} */,
  {32'h408c3375, 32'h4099fe23} /* (27, 3, 28) {real, imag} */,
  {32'hc057d16d, 32'hc099f7ff} /* (27, 3, 27) {real, imag} */,
  {32'hc06b7706, 32'h3fc648d3} /* (27, 3, 26) {real, imag} */,
  {32'h3fc8e2c0, 32'hc01fca64} /* (27, 3, 25) {real, imag} */,
  {32'h4052654c, 32'hc0b6088c} /* (27, 3, 24) {real, imag} */,
  {32'h4064cb4c, 32'h3f0ed7ff} /* (27, 3, 23) {real, imag} */,
  {32'hc069cb85, 32'h3fec087f} /* (27, 3, 22) {real, imag} */,
  {32'h3de76713, 32'h3f3fcdbe} /* (27, 3, 21) {real, imag} */,
  {32'hbffcdf3b, 32'hbf1257e2} /* (27, 3, 20) {real, imag} */,
  {32'h3fb75ce3, 32'h3ffd8a3e} /* (27, 3, 19) {real, imag} */,
  {32'h4002a637, 32'hbfa0c9f3} /* (27, 3, 18) {real, imag} */,
  {32'h3fcedf2a, 32'h3eccac7f} /* (27, 3, 17) {real, imag} */,
  {32'hbf1179e7, 32'h3f486f0e} /* (27, 3, 16) {real, imag} */,
  {32'hbfb13587, 32'hbf9ffe99} /* (27, 3, 15) {real, imag} */,
  {32'hbff6e634, 32'hbf6cb042} /* (27, 3, 14) {real, imag} */,
  {32'hbdc33c44, 32'hbfc9ed6c} /* (27, 3, 13) {real, imag} */,
  {32'h3fab9341, 32'h4072a760} /* (27, 3, 12) {real, imag} */,
  {32'h3ec3eef8, 32'h3f5a83fb} /* (27, 3, 11) {real, imag} */,
  {32'hbfa37384, 32'hbf537098} /* (27, 3, 10) {real, imag} */,
  {32'hbe95d50a, 32'hc0840704} /* (27, 3, 9) {real, imag} */,
  {32'hbfed8ecc, 32'hc0253476} /* (27, 3, 8) {real, imag} */,
  {32'hc01f906b, 32'h40ba0525} /* (27, 3, 7) {real, imag} */,
  {32'h409c0eea, 32'hc0a6b752} /* (27, 3, 6) {real, imag} */,
  {32'hbeb857db, 32'h406bee5c} /* (27, 3, 5) {real, imag} */,
  {32'hc0593fcc, 32'h3f376669} /* (27, 3, 4) {real, imag} */,
  {32'h3ee62d79, 32'hbebee5d6} /* (27, 3, 3) {real, imag} */,
  {32'h40bceed7, 32'hc098f1f8} /* (27, 3, 2) {real, imag} */,
  {32'hc0568e65, 32'h40c03f11} /* (27, 3, 1) {real, imag} */,
  {32'h40c7d274, 32'h40e61689} /* (27, 3, 0) {real, imag} */,
  {32'hc1a82d7f, 32'hc1c7bc0f} /* (27, 2, 31) {real, imag} */,
  {32'h41162c06, 32'h4158debb} /* (27, 2, 30) {real, imag} */,
  {32'hc10b551f, 32'hc0c6d987} /* (27, 2, 29) {real, imag} */,
  {32'hc0f8113a, 32'hbfaa624d} /* (27, 2, 28) {real, imag} */,
  {32'h402c482e, 32'h3f94c0cc} /* (27, 2, 27) {real, imag} */,
  {32'h40c4968c, 32'h3f73ad20} /* (27, 2, 26) {real, imag} */,
  {32'hc0c699f9, 32'h3fd28b11} /* (27, 2, 25) {real, imag} */,
  {32'h409ae812, 32'hbd72b0d9} /* (27, 2, 24) {real, imag} */,
  {32'h408144c1, 32'hc026f217} /* (27, 2, 23) {real, imag} */,
  {32'h3f6e2f07, 32'hbe807e23} /* (27, 2, 22) {real, imag} */,
  {32'h3fbe1424, 32'hc00aa8dc} /* (27, 2, 21) {real, imag} */,
  {32'h3f52c271, 32'h3e40a0eb} /* (27, 2, 20) {real, imag} */,
  {32'h3e98d62b, 32'hbfe45646} /* (27, 2, 19) {real, imag} */,
  {32'h3f5c026b, 32'hbfdb7718} /* (27, 2, 18) {real, imag} */,
  {32'hbf3da239, 32'h3fdb4bd5} /* (27, 2, 17) {real, imag} */,
  {32'h3ee1cc05, 32'hbf6279c4} /* (27, 2, 16) {real, imag} */,
  {32'h3f1eebc2, 32'hbe96032d} /* (27, 2, 15) {real, imag} */,
  {32'h400ff890, 32'h4017f52d} /* (27, 2, 14) {real, imag} */,
  {32'hbfbffae9, 32'h3e670592} /* (27, 2, 13) {real, imag} */,
  {32'hbd7cce16, 32'hbf377f67} /* (27, 2, 12) {real, imag} */,
  {32'hbeabc85a, 32'hbda4229a} /* (27, 2, 11) {real, imag} */,
  {32'h3fa17119, 32'hbf7ca388} /* (27, 2, 10) {real, imag} */,
  {32'hbfc42388, 32'hbf87605b} /* (27, 2, 9) {real, imag} */,
  {32'h3f10ba7f, 32'hc02f5192} /* (27, 2, 8) {real, imag} */,
  {32'hc027a38e, 32'hbfe5d850} /* (27, 2, 7) {real, imag} */,
  {32'h40508184, 32'hc03df438} /* (27, 2, 6) {real, imag} */,
  {32'hc0567007, 32'h40e2ed8a} /* (27, 2, 5) {real, imag} */,
  {32'hc01541ec, 32'hc0b22f88} /* (27, 2, 4) {real, imag} */,
  {32'h3f0e996d, 32'h3f4d643d} /* (27, 2, 3) {real, imag} */,
  {32'h413d996e, 32'h41975b94} /* (27, 2, 2) {real, imag} */,
  {32'hc11282a5, 32'hc1938103} /* (27, 2, 1) {real, imag} */,
  {32'h408f6436, 32'hc1d11684} /* (27, 2, 0) {real, imag} */,
  {32'h41da5ff9, 32'h419094fc} /* (27, 1, 31) {real, imag} */,
  {32'hc0e75f58, 32'hc0ea406e} /* (27, 1, 30) {real, imag} */,
  {32'h402ad420, 32'h3ff72679} /* (27, 1, 29) {real, imag} */,
  {32'h409b6c95, 32'h3e5219cc} /* (27, 1, 28) {real, imag} */,
  {32'hc11d150a, 32'hc0adf41d} /* (27, 1, 27) {real, imag} */,
  {32'hbfdd9fcb, 32'hba02e6c4} /* (27, 1, 26) {real, imag} */,
  {32'hbf168fc2, 32'h40dc7c6e} /* (27, 1, 25) {real, imag} */,
  {32'hc0735bea, 32'hc000afaa} /* (27, 1, 24) {real, imag} */,
  {32'hbf2c7b1b, 32'h3e36ccf8} /* (27, 1, 23) {real, imag} */,
  {32'h3f310329, 32'h3ebb188b} /* (27, 1, 22) {real, imag} */,
  {32'hbfb3cb61, 32'hbe486256} /* (27, 1, 21) {real, imag} */,
  {32'hbf294eac, 32'h400e3b14} /* (27, 1, 20) {real, imag} */,
  {32'h3eef630c, 32'hbf0b56b3} /* (27, 1, 19) {real, imag} */,
  {32'h3e44b447, 32'hbfdd867e} /* (27, 1, 18) {real, imag} */,
  {32'h3e38d079, 32'hbfad38c6} /* (27, 1, 17) {real, imag} */,
  {32'h3f7377e9, 32'h3ecec20d} /* (27, 1, 16) {real, imag} */,
  {32'hbf6d8895, 32'hbff7cc2c} /* (27, 1, 15) {real, imag} */,
  {32'h3fd33820, 32'h40286d7f} /* (27, 1, 14) {real, imag} */,
  {32'h3fd97a92, 32'h3fd8e425} /* (27, 1, 13) {real, imag} */,
  {32'h3f327c75, 32'h3f28ada2} /* (27, 1, 12) {real, imag} */,
  {32'hbecfac62, 32'hc03b0c96} /* (27, 1, 11) {real, imag} */,
  {32'h3e617b9a, 32'hbea7a5d4} /* (27, 1, 10) {real, imag} */,
  {32'hbf51b2b5, 32'hbff66049} /* (27, 1, 9) {real, imag} */,
  {32'h3f96c8fb, 32'hc0ef1ee6} /* (27, 1, 8) {real, imag} */,
  {32'h405a8f36, 32'h4082c89c} /* (27, 1, 7) {real, imag} */,
  {32'h405d669e, 32'hbdc0627e} /* (27, 1, 6) {real, imag} */,
  {32'hbfc70060, 32'hc018e11d} /* (27, 1, 5) {real, imag} */,
  {32'hbfb114fa, 32'h4079456f} /* (27, 1, 4) {real, imag} */,
  {32'hbd4191cf, 32'hc12f0c18} /* (27, 1, 3) {real, imag} */,
  {32'h412302a0, 32'hc1a09a80} /* (27, 1, 2) {real, imag} */,
  {32'h3f566ac7, 32'h420fff4d} /* (27, 1, 1) {real, imag} */,
  {32'h4119c833, 32'h41f9609c} /* (27, 1, 0) {real, imag} */,
  {32'h41bf434e, 32'h406a13f0} /* (27, 0, 31) {real, imag} */,
  {32'hc155d1fa, 32'hc08f3c4a} /* (27, 0, 30) {real, imag} */,
  {32'h4014e698, 32'hc0c71ffa} /* (27, 0, 29) {real, imag} */,
  {32'h3f5f5806, 32'hbec6de7a} /* (27, 0, 28) {real, imag} */,
  {32'h3fd4f815, 32'hbf82b3d8} /* (27, 0, 27) {real, imag} */,
  {32'h400b9005, 32'hbf77f103} /* (27, 0, 26) {real, imag} */,
  {32'hbfddc9c2, 32'hbfd3b395} /* (27, 0, 25) {real, imag} */,
  {32'hc06d38ef, 32'hc00658f4} /* (27, 0, 24) {real, imag} */,
  {32'hbffd0919, 32'h3fac93ef} /* (27, 0, 23) {real, imag} */,
  {32'hc063744f, 32'hbe8423e7} /* (27, 0, 22) {real, imag} */,
  {32'hbf7722d3, 32'h3f264e94} /* (27, 0, 21) {real, imag} */,
  {32'h3fb3ff8e, 32'h4033920e} /* (27, 0, 20) {real, imag} */,
  {32'h4018a80e, 32'h400d4a76} /* (27, 0, 19) {real, imag} */,
  {32'hbf4d7535, 32'hbfcdcc67} /* (27, 0, 18) {real, imag} */,
  {32'hbe1f8122, 32'hbecd5c71} /* (27, 0, 17) {real, imag} */,
  {32'h40203f1d, 32'h3f2dbd3d} /* (27, 0, 16) {real, imag} */,
  {32'hbddbc3a8, 32'hbfa05ea2} /* (27, 0, 15) {real, imag} */,
  {32'h402e143d, 32'hbec36a3e} /* (27, 0, 14) {real, imag} */,
  {32'h3ea1555c, 32'hbfb35a7a} /* (27, 0, 13) {real, imag} */,
  {32'hbe8342f9, 32'h4078eb62} /* (27, 0, 12) {real, imag} */,
  {32'hbe4f03d4, 32'hc0286376} /* (27, 0, 11) {real, imag} */,
  {32'hc046c0e9, 32'h3f664861} /* (27, 0, 10) {real, imag} */,
  {32'hc0862a32, 32'h3eb7f0c6} /* (27, 0, 9) {real, imag} */,
  {32'h3f697f93, 32'h40b1186f} /* (27, 0, 8) {real, imag} */,
  {32'hbfc4af65, 32'h40100ce9} /* (27, 0, 7) {real, imag} */,
  {32'hc001eb1b, 32'h3f98fbe5} /* (27, 0, 6) {real, imag} */,
  {32'h3ee28906, 32'hc1039572} /* (27, 0, 5) {real, imag} */,
  {32'h3f7e5061, 32'hc0b994c0} /* (27, 0, 4) {real, imag} */,
  {32'hc09d2a03, 32'h3fe69f80} /* (27, 0, 3) {real, imag} */,
  {32'h408e1be2, 32'hc0ebf752} /* (27, 0, 2) {real, imag} */,
  {32'h3ebdfd1d, 32'h41dc1fd6} /* (27, 0, 1) {real, imag} */,
  {32'h402bf908, 32'h41a493ea} /* (27, 0, 0) {real, imag} */,
  {32'h40254c21, 32'hc010b9cb} /* (26, 31, 31) {real, imag} */,
  {32'hc0a165ba, 32'hbfd8d645} /* (26, 31, 30) {real, imag} */,
  {32'hbfddd0c4, 32'hbfc5c2f0} /* (26, 31, 29) {real, imag} */,
  {32'h405ef213, 32'hbeee749f} /* (26, 31, 28) {real, imag} */,
  {32'h3fd042bf, 32'hbf547200} /* (26, 31, 27) {real, imag} */,
  {32'hbfdc08f6, 32'h3f86795b} /* (26, 31, 26) {real, imag} */,
  {32'hc00cdb3f, 32'h3f047097} /* (26, 31, 25) {real, imag} */,
  {32'hbfe38f38, 32'hbdea8ccb} /* (26, 31, 24) {real, imag} */,
  {32'h3d8ea803, 32'hbe844276} /* (26, 31, 23) {real, imag} */,
  {32'hbeca6573, 32'h3f457d48} /* (26, 31, 22) {real, imag} */,
  {32'hbfcf6ced, 32'hbf841dee} /* (26, 31, 21) {real, imag} */,
  {32'hbfe927c5, 32'h3fbe7e27} /* (26, 31, 20) {real, imag} */,
  {32'hbf94b634, 32'hc092b145} /* (26, 31, 19) {real, imag} */,
  {32'h3dc3d062, 32'h406662a7} /* (26, 31, 18) {real, imag} */,
  {32'h3f630e27, 32'hbf20c22e} /* (26, 31, 17) {real, imag} */,
  {32'hbf970166, 32'hbb70d60b} /* (26, 31, 16) {real, imag} */,
  {32'h3f50d2f5, 32'hbed5c50a} /* (26, 31, 15) {real, imag} */,
  {32'h40553579, 32'hbf45d2db} /* (26, 31, 14) {real, imag} */,
  {32'hbf274220, 32'hbf4c7075} /* (26, 31, 13) {real, imag} */,
  {32'h4003492a, 32'hc060efa2} /* (26, 31, 12) {real, imag} */,
  {32'hc0244862, 32'hbeb538b9} /* (26, 31, 11) {real, imag} */,
  {32'h405cc29b, 32'hbf831b1f} /* (26, 31, 10) {real, imag} */,
  {32'hc031aec7, 32'h4022b2d0} /* (26, 31, 9) {real, imag} */,
  {32'hbda22654, 32'h4077f0bf} /* (26, 31, 8) {real, imag} */,
  {32'hbf8a8852, 32'h3e42121d} /* (26, 31, 7) {real, imag} */,
  {32'h402c43b9, 32'h3fec328e} /* (26, 31, 6) {real, imag} */,
  {32'h3f17178b, 32'h3eaf24de} /* (26, 31, 5) {real, imag} */,
  {32'h409a9625, 32'hc08eb14c} /* (26, 31, 4) {real, imag} */,
  {32'hbfc7890e, 32'h409daa5a} /* (26, 31, 3) {real, imag} */,
  {32'hbfa02e9b, 32'h402730e6} /* (26, 31, 2) {real, imag} */,
  {32'hc00d659d, 32'h3ffdb69d} /* (26, 31, 1) {real, imag} */,
  {32'h40da89fd, 32'h40ada06d} /* (26, 31, 0) {real, imag} */,
  {32'hc094fde1, 32'hc00574d0} /* (26, 30, 31) {real, imag} */,
  {32'hc021b009, 32'h408f9777} /* (26, 30, 30) {real, imag} */,
  {32'h408ed09f, 32'h4097124e} /* (26, 30, 29) {real, imag} */,
  {32'h3f45075f, 32'hc045920f} /* (26, 30, 28) {real, imag} */,
  {32'hc07814a4, 32'hc029bbc2} /* (26, 30, 27) {real, imag} */,
  {32'h40174786, 32'hc021126d} /* (26, 30, 26) {real, imag} */,
  {32'hc01384c3, 32'hc02ac462} /* (26, 30, 25) {real, imag} */,
  {32'h40337ebb, 32'hbfc2ca4a} /* (26, 30, 24) {real, imag} */,
  {32'hc00260d3, 32'h3cea575b} /* (26, 30, 23) {real, imag} */,
  {32'hbf3c4a28, 32'h3f5a84b0} /* (26, 30, 22) {real, imag} */,
  {32'hbd780b4c, 32'hbf00bad3} /* (26, 30, 21) {real, imag} */,
  {32'hbf9ddb82, 32'hc00b93bc} /* (26, 30, 20) {real, imag} */,
  {32'hbebaee0e, 32'hbf3ee320} /* (26, 30, 19) {real, imag} */,
  {32'h3e1f833e, 32'h3fc1092a} /* (26, 30, 18) {real, imag} */,
  {32'h3d608073, 32'hbf3c1301} /* (26, 30, 17) {real, imag} */,
  {32'h3f0bec93, 32'hbf2fe88e} /* (26, 30, 16) {real, imag} */,
  {32'h3f17f216, 32'h3df3b102} /* (26, 30, 15) {real, imag} */,
  {32'hbe659c17, 32'hbed4bd46} /* (26, 30, 14) {real, imag} */,
  {32'h3f64a396, 32'h3f1596ac} /* (26, 30, 13) {real, imag} */,
  {32'h3e956e2b, 32'hc00327d7} /* (26, 30, 12) {real, imag} */,
  {32'hbf45b2b5, 32'h404cd1b1} /* (26, 30, 11) {real, imag} */,
  {32'h3d3d5e44, 32'h402df3d3} /* (26, 30, 10) {real, imag} */,
  {32'hbe91cc60, 32'hc063b0f8} /* (26, 30, 9) {real, imag} */,
  {32'hc086f4a6, 32'hc072a58f} /* (26, 30, 8) {real, imag} */,
  {32'h408d016f, 32'h3f2f1e01} /* (26, 30, 7) {real, imag} */,
  {32'hc0540ec3, 32'hbf08e127} /* (26, 30, 6) {real, imag} */,
  {32'hc00519da, 32'hc051c7be} /* (26, 30, 5) {real, imag} */,
  {32'hc0732384, 32'h40bbbcdd} /* (26, 30, 4) {real, imag} */,
  {32'hc08aa37f, 32'h3f8961d1} /* (26, 30, 3) {real, imag} */,
  {32'h40111794, 32'h3f6a094c} /* (26, 30, 2) {real, imag} */,
  {32'h4177f004, 32'hbf45dfa0} /* (26, 30, 1) {real, imag} */,
  {32'hc04bb2ad, 32'h40d9123d} /* (26, 30, 0) {real, imag} */,
  {32'h409e1ac8, 32'h409c9657} /* (26, 29, 31) {real, imag} */,
  {32'h40818f2c, 32'hbe64e367} /* (26, 29, 30) {real, imag} */,
  {32'hc0ac7eaf, 32'hc0363480} /* (26, 29, 29) {real, imag} */,
  {32'h400ea393, 32'h3f3af0db} /* (26, 29, 28) {real, imag} */,
  {32'h3f4b099e, 32'h40cde56b} /* (26, 29, 27) {real, imag} */,
  {32'hbfcaa794, 32'hbf076948} /* (26, 29, 26) {real, imag} */,
  {32'hbfac9b5f, 32'h3f5467b3} /* (26, 29, 25) {real, imag} */,
  {32'hbfb15f48, 32'h3eb4a96e} /* (26, 29, 24) {real, imag} */,
  {32'hbf4e15d5, 32'h3f320b60} /* (26, 29, 23) {real, imag} */,
  {32'hbd9430d8, 32'h3f17bf8b} /* (26, 29, 22) {real, imag} */,
  {32'hbd84e2fa, 32'h3ff69bc3} /* (26, 29, 21) {real, imag} */,
  {32'hc0029e8b, 32'h3ee2df02} /* (26, 29, 20) {real, imag} */,
  {32'h3de224b2, 32'h3f45a578} /* (26, 29, 19) {real, imag} */,
  {32'h3f460090, 32'h4040bb10} /* (26, 29, 18) {real, imag} */,
  {32'hbd1e3d90, 32'hbf5faab7} /* (26, 29, 17) {real, imag} */,
  {32'h4000a010, 32'hbfb2bfb8} /* (26, 29, 16) {real, imag} */,
  {32'h3ef2480e, 32'hbf8a7ea8} /* (26, 29, 15) {real, imag} */,
  {32'hbdfc664c, 32'h3fc8e794} /* (26, 29, 14) {real, imag} */,
  {32'h3fd21d92, 32'hbee0d861} /* (26, 29, 13) {real, imag} */,
  {32'hbfddb37b, 32'hbf16d481} /* (26, 29, 12) {real, imag} */,
  {32'h400a163a, 32'hc09ee6fa} /* (26, 29, 11) {real, imag} */,
  {32'h3edaa3b0, 32'h4083f50e} /* (26, 29, 10) {real, imag} */,
  {32'h3fb52286, 32'h40256647} /* (26, 29, 9) {real, imag} */,
  {32'h3eb0fa07, 32'h3e07b6b6} /* (26, 29, 8) {real, imag} */,
  {32'h3e975dd1, 32'h40629c63} /* (26, 29, 7) {real, imag} */,
  {32'h3fa31404, 32'hc0420fb4} /* (26, 29, 6) {real, imag} */,
  {32'hbe90aad0, 32'h3faeb037} /* (26, 29, 5) {real, imag} */,
  {32'h3f74e174, 32'hbfb99042} /* (26, 29, 4) {real, imag} */,
  {32'h3f62ba39, 32'hbf8e6837} /* (26, 29, 3) {real, imag} */,
  {32'h4039cad5, 32'h4036926a} /* (26, 29, 2) {real, imag} */,
  {32'h4003a051, 32'hc0db2f83} /* (26, 29, 1) {real, imag} */,
  {32'hbfe5c67b, 32'hc06f525c} /* (26, 29, 0) {real, imag} */,
  {32'h408c4afe, 32'hbfd16813} /* (26, 28, 31) {real, imag} */,
  {32'hbfd45848, 32'hc0060e3e} /* (26, 28, 30) {real, imag} */,
  {32'hc04fc698, 32'h40d783f5} /* (26, 28, 29) {real, imag} */,
  {32'h3fdc2c2b, 32'h4028e9bc} /* (26, 28, 28) {real, imag} */,
  {32'h3f65fc91, 32'hc0012ccc} /* (26, 28, 27) {real, imag} */,
  {32'h3f88ae55, 32'h3fe1c387} /* (26, 28, 26) {real, imag} */,
  {32'hc03e9322, 32'h3da085d5} /* (26, 28, 25) {real, imag} */,
  {32'hc0245e40, 32'hbec46166} /* (26, 28, 24) {real, imag} */,
  {32'hc0950b40, 32'hc00c2721} /* (26, 28, 23) {real, imag} */,
  {32'h4017486a, 32'h3f5bb70d} /* (26, 28, 22) {real, imag} */,
  {32'h3fdf4300, 32'hbf132931} /* (26, 28, 21) {real, imag} */,
  {32'hbf97d385, 32'hbe5315fc} /* (26, 28, 20) {real, imag} */,
  {32'hbeecfcd8, 32'h3eeb253e} /* (26, 28, 19) {real, imag} */,
  {32'hbd641b5b, 32'hbe087ced} /* (26, 28, 18) {real, imag} */,
  {32'h3ec6baa1, 32'hbf298374} /* (26, 28, 17) {real, imag} */,
  {32'h3ee8d7ce, 32'h3fb067e6} /* (26, 28, 16) {real, imag} */,
  {32'hc003b0e1, 32'h3d593a13} /* (26, 28, 15) {real, imag} */,
  {32'h3e50d875, 32'h3e495b8d} /* (26, 28, 14) {real, imag} */,
  {32'h3fb50ce1, 32'hc031ca38} /* (26, 28, 13) {real, imag} */,
  {32'h401e087c, 32'hbf516b46} /* (26, 28, 12) {real, imag} */,
  {32'hc02b9eae, 32'hbf96eb80} /* (26, 28, 11) {real, imag} */,
  {32'h401ea21c, 32'hc000137f} /* (26, 28, 10) {real, imag} */,
  {32'hbff4d61d, 32'hc07d1a78} /* (26, 28, 9) {real, imag} */,
  {32'h3fad1275, 32'h3fab780a} /* (26, 28, 8) {real, imag} */,
  {32'hc057ab43, 32'hbfa53ff3} /* (26, 28, 7) {real, imag} */,
  {32'hbcee8db6, 32'h40904e26} /* (26, 28, 6) {real, imag} */,
  {32'h4007c61c, 32'h40108763} /* (26, 28, 5) {real, imag} */,
  {32'hc0993046, 32'hc08de49c} /* (26, 28, 4) {real, imag} */,
  {32'h3f31c94d, 32'h40d09fc5} /* (26, 28, 3) {real, imag} */,
  {32'h3dad635a, 32'h3f0cf19e} /* (26, 28, 2) {real, imag} */,
  {32'h3e2b9e70, 32'hc0694071} /* (26, 28, 1) {real, imag} */,
  {32'h40796794, 32'h3fd6a601} /* (26, 28, 0) {real, imag} */,
  {32'h4067b859, 32'h406af89b} /* (26, 27, 31) {real, imag} */,
  {32'hbfbf8687, 32'h408ac48e} /* (26, 27, 30) {real, imag} */,
  {32'hbf06a079, 32'hbd372c5d} /* (26, 27, 29) {real, imag} */,
  {32'h4006fad8, 32'hbfc51e82} /* (26, 27, 28) {real, imag} */,
  {32'h3f5c9302, 32'h3f524488} /* (26, 27, 27) {real, imag} */,
  {32'h3f7cdaa0, 32'h3e0fa616} /* (26, 27, 26) {real, imag} */,
  {32'h3fed661f, 32'hc0922340} /* (26, 27, 25) {real, imag} */,
  {32'hbf89d831, 32'h3ec66967} /* (26, 27, 24) {real, imag} */,
  {32'hbec5d478, 32'h408d1901} /* (26, 27, 23) {real, imag} */,
  {32'hc057289c, 32'hbff8f978} /* (26, 27, 22) {real, imag} */,
  {32'h3ffa659c, 32'hbee53f81} /* (26, 27, 21) {real, imag} */,
  {32'hc06c0f0b, 32'h3e8a40fe} /* (26, 27, 20) {real, imag} */,
  {32'h40298669, 32'hbf84df96} /* (26, 27, 19) {real, imag} */,
  {32'h3e609241, 32'hbf6e2563} /* (26, 27, 18) {real, imag} */,
  {32'hbc39cecd, 32'hc005cc26} /* (26, 27, 17) {real, imag} */,
  {32'hc0515bef, 32'h3faa0599} /* (26, 27, 16) {real, imag} */,
  {32'hbed6e592, 32'h401f99f7} /* (26, 27, 15) {real, imag} */,
  {32'h3fa837c3, 32'h3e9be891} /* (26, 27, 14) {real, imag} */,
  {32'h3d87cd45, 32'h3f4600d6} /* (26, 27, 13) {real, imag} */,
  {32'h3fc2c72e, 32'h40155204} /* (26, 27, 12) {real, imag} */,
  {32'hc03564fc, 32'h4053665b} /* (26, 27, 11) {real, imag} */,
  {32'h3ba9ee3b, 32'h3fcecced} /* (26, 27, 10) {real, imag} */,
  {32'hbfa2d56b, 32'h4019b1dc} /* (26, 27, 9) {real, imag} */,
  {32'hc05553a0, 32'h3f99a487} /* (26, 27, 8) {real, imag} */,
  {32'hbfe8ec74, 32'h3fc71690} /* (26, 27, 7) {real, imag} */,
  {32'hbfe5678a, 32'hbe84dbb4} /* (26, 27, 6) {real, imag} */,
  {32'h3f9ed637, 32'h400f332f} /* (26, 27, 5) {real, imag} */,
  {32'h3e554d58, 32'hc0f401f8} /* (26, 27, 4) {real, imag} */,
  {32'hc0b0fc94, 32'hc0204bbc} /* (26, 27, 3) {real, imag} */,
  {32'h408baa81, 32'hbdf9e99a} /* (26, 27, 2) {real, imag} */,
  {32'h3f3b570a, 32'hbfa61197} /* (26, 27, 1) {real, imag} */,
  {32'hc0a5ff76, 32'hc00cf3cd} /* (26, 27, 0) {real, imag} */,
  {32'h3faa677d, 32'hc0009b89} /* (26, 26, 31) {real, imag} */,
  {32'h3f40747d, 32'hbfe58c61} /* (26, 26, 30) {real, imag} */,
  {32'h3f652bc5, 32'h4037b723} /* (26, 26, 29) {real, imag} */,
  {32'hc00136ed, 32'h401ce551} /* (26, 26, 28) {real, imag} */,
  {32'hbf9e28c8, 32'hc09f3e10} /* (26, 26, 27) {real, imag} */,
  {32'hbf6b6f7a, 32'hbfc556d9} /* (26, 26, 26) {real, imag} */,
  {32'h40114447, 32'h40df1fa6} /* (26, 26, 25) {real, imag} */,
  {32'hc0377333, 32'h3fa7f883} /* (26, 26, 24) {real, imag} */,
  {32'h402dfd9c, 32'h4004a85a} /* (26, 26, 23) {real, imag} */,
  {32'hc0977cdf, 32'hc08c6e64} /* (26, 26, 22) {real, imag} */,
  {32'hbfde75c1, 32'hbe7ac317} /* (26, 26, 21) {real, imag} */,
  {32'h3e3fe59e, 32'h3f4049a4} /* (26, 26, 20) {real, imag} */,
  {32'h3fc8a97a, 32'h3eaf817f} /* (26, 26, 19) {real, imag} */,
  {32'hbf5238cf, 32'hbf5c9230} /* (26, 26, 18) {real, imag} */,
  {32'hbfa7e70e, 32'hbfa0b9ce} /* (26, 26, 17) {real, imag} */,
  {32'hbe93a315, 32'hc025a53d} /* (26, 26, 16) {real, imag} */,
  {32'h3fcbe06d, 32'h3f36d20a} /* (26, 26, 15) {real, imag} */,
  {32'hbf1b1d84, 32'hc0605020} /* (26, 26, 14) {real, imag} */,
  {32'hbe7793a8, 32'h40002282} /* (26, 26, 13) {real, imag} */,
  {32'hc01c9ce9, 32'h40739c27} /* (26, 26, 12) {real, imag} */,
  {32'h3fd0943b, 32'hbfb1554a} /* (26, 26, 11) {real, imag} */,
  {32'h3e6664ea, 32'hbea287c6} /* (26, 26, 10) {real, imag} */,
  {32'hc0764b54, 32'hbf2f4879} /* (26, 26, 9) {real, imag} */,
  {32'h3f920603, 32'hbe884d98} /* (26, 26, 8) {real, imag} */,
  {32'h4006d6a2, 32'h3fd2e224} /* (26, 26, 7) {real, imag} */,
  {32'h3f1744d3, 32'h3f6add00} /* (26, 26, 6) {real, imag} */,
  {32'h401c4a3d, 32'h403ba499} /* (26, 26, 5) {real, imag} */,
  {32'h401a30bb, 32'hc06574e7} /* (26, 26, 4) {real, imag} */,
  {32'h3fec65f6, 32'h3f3ef286} /* (26, 26, 3) {real, imag} */,
  {32'hc0b8876e, 32'h401ff751} /* (26, 26, 2) {real, imag} */,
  {32'hbf6c405a, 32'h3f6497c5} /* (26, 26, 1) {real, imag} */,
  {32'hbf1908b5, 32'h40595e66} /* (26, 26, 0) {real, imag} */,
  {32'h3f1d0cae, 32'h3fddd69a} /* (26, 25, 31) {real, imag} */,
  {32'hc06abe98, 32'hc00a08c2} /* (26, 25, 30) {real, imag} */,
  {32'h40cda99a, 32'hbfd4dcc3} /* (26, 25, 29) {real, imag} */,
  {32'h40e1cb89, 32'h3fa81189} /* (26, 25, 28) {real, imag} */,
  {32'hc015fa14, 32'hbeef3a1f} /* (26, 25, 27) {real, imag} */,
  {32'h3e901b9b, 32'hbf6e4e26} /* (26, 25, 26) {real, imag} */,
  {32'hbe077fe5, 32'hbdb4d627} /* (26, 25, 25) {real, imag} */,
  {32'hbfeb9576, 32'h3fa7ac6c} /* (26, 25, 24) {real, imag} */,
  {32'h401b37c6, 32'h3ef01082} /* (26, 25, 23) {real, imag} */,
  {32'h405b7d15, 32'h400624bb} /* (26, 25, 22) {real, imag} */,
  {32'hc032baf8, 32'h3e9a5d9f} /* (26, 25, 21) {real, imag} */,
  {32'hc01c73d2, 32'h3faa3ea6} /* (26, 25, 20) {real, imag} */,
  {32'hc01539cd, 32'hbda27fd2} /* (26, 25, 19) {real, imag} */,
  {32'hbfe55b7b, 32'h40087eac} /* (26, 25, 18) {real, imag} */,
  {32'hc01fac40, 32'h400fc751} /* (26, 25, 17) {real, imag} */,
  {32'h3f8bc452, 32'hbfd897c7} /* (26, 25, 16) {real, imag} */,
  {32'hc07b2d16, 32'hbf64ab32} /* (26, 25, 15) {real, imag} */,
  {32'hbd915c9d, 32'hbe35d4de} /* (26, 25, 14) {real, imag} */,
  {32'h3f67505f, 32'hbf6af4aa} /* (26, 25, 13) {real, imag} */,
  {32'hbfd46c0c, 32'h3f98f295} /* (26, 25, 12) {real, imag} */,
  {32'h40886654, 32'h3f3e7491} /* (26, 25, 11) {real, imag} */,
  {32'h4000b0e4, 32'hbe8ffa3e} /* (26, 25, 10) {real, imag} */,
  {32'hbff55c28, 32'h3e8a5d77} /* (26, 25, 9) {real, imag} */,
  {32'hc008d310, 32'hbdf059c9} /* (26, 25, 8) {real, imag} */,
  {32'h40a1982b, 32'h3f359295} /* (26, 25, 7) {real, imag} */,
  {32'h3edbccf1, 32'hc056a618} /* (26, 25, 6) {real, imag} */,
  {32'hc02406f5, 32'h40338707} /* (26, 25, 5) {real, imag} */,
  {32'h40630b8f, 32'h3f1fe4e8} /* (26, 25, 4) {real, imag} */,
  {32'h3ff36b32, 32'hc0088079} /* (26, 25, 3) {real, imag} */,
  {32'h4074d4ba, 32'h40a6e606} /* (26, 25, 2) {real, imag} */,
  {32'h3fc324c6, 32'hc0b210e1} /* (26, 25, 1) {real, imag} */,
  {32'hc0135aa7, 32'h40ba7ca0} /* (26, 25, 0) {real, imag} */,
  {32'hbfaf2cd4, 32'hc07a0d19} /* (26, 24, 31) {real, imag} */,
  {32'h3e5620ff, 32'hbfbc79a3} /* (26, 24, 30) {real, imag} */,
  {32'hbf978c2b, 32'h40269671} /* (26, 24, 29) {real, imag} */,
  {32'hc089f3b5, 32'h3f9be7d7} /* (26, 24, 28) {real, imag} */,
  {32'hc025376b, 32'h3e1fef39} /* (26, 24, 27) {real, imag} */,
  {32'hbf4c1b81, 32'hc00d3d7e} /* (26, 24, 26) {real, imag} */,
  {32'h401e9261, 32'h3dd0774a} /* (26, 24, 25) {real, imag} */,
  {32'h4004a31f, 32'h401e0f5a} /* (26, 24, 24) {real, imag} */,
  {32'h3f31eade, 32'hbfffbab3} /* (26, 24, 23) {real, imag} */,
  {32'hc003d8d9, 32'h3f19c529} /* (26, 24, 22) {real, imag} */,
  {32'hbf47e9dc, 32'h3fa32ca7} /* (26, 24, 21) {real, imag} */,
  {32'h3f7d154a, 32'h4067c5d5} /* (26, 24, 20) {real, imag} */,
  {32'hbec3c69c, 32'hc0925b33} /* (26, 24, 19) {real, imag} */,
  {32'hc004c6f0, 32'hbe7809d0} /* (26, 24, 18) {real, imag} */,
  {32'h3ded34e9, 32'h3f6f47ad} /* (26, 24, 17) {real, imag} */,
  {32'h3eca2b8b, 32'h3f4338cd} /* (26, 24, 16) {real, imag} */,
  {32'h3f630c4b, 32'hbf5c30c6} /* (26, 24, 15) {real, imag} */,
  {32'hbf985a73, 32'h3eacc059} /* (26, 24, 14) {real, imag} */,
  {32'hc00af6a5, 32'h400df1db} /* (26, 24, 13) {real, imag} */,
  {32'hbde3d9b7, 32'h3f798e3c} /* (26, 24, 12) {real, imag} */,
  {32'hbfa750ad, 32'h3f2746f3} /* (26, 24, 11) {real, imag} */,
  {32'hbfba8024, 32'hbff5484a} /* (26, 24, 10) {real, imag} */,
  {32'h405e4209, 32'h408cf861} /* (26, 24, 9) {real, imag} */,
  {32'h3f1aca0c, 32'hc0256bef} /* (26, 24, 8) {real, imag} */,
  {32'hbf2a19bd, 32'h3ffd715d} /* (26, 24, 7) {real, imag} */,
  {32'hbfe63b45, 32'hc08d0b30} /* (26, 24, 6) {real, imag} */,
  {32'hc066521e, 32'h4008485e} /* (26, 24, 5) {real, imag} */,
  {32'hc0388e5e, 32'h404764a2} /* (26, 24, 4) {real, imag} */,
  {32'hbfcd5d8f, 32'hc0507b88} /* (26, 24, 3) {real, imag} */,
  {32'h400b176a, 32'h3fb3371c} /* (26, 24, 2) {real, imag} */,
  {32'h3ea1b563, 32'hc026e9af} /* (26, 24, 1) {real, imag} */,
  {32'h3ec5eb66, 32'h3f4bc3cc} /* (26, 24, 0) {real, imag} */,
  {32'hbf20550a, 32'hbe3efe72} /* (26, 23, 31) {real, imag} */,
  {32'h40641196, 32'hbe4053c9} /* (26, 23, 30) {real, imag} */,
  {32'h40754288, 32'hc000d935} /* (26, 23, 29) {real, imag} */,
  {32'hbfdba76f, 32'h3fac408b} /* (26, 23, 28) {real, imag} */,
  {32'h3f177b88, 32'hbfba4309} /* (26, 23, 27) {real, imag} */,
  {32'h3f1e1dcc, 32'hbfd2a41a} /* (26, 23, 26) {real, imag} */,
  {32'h40778d07, 32'h404d752e} /* (26, 23, 25) {real, imag} */,
  {32'h3f8db2d6, 32'hbe70adc2} /* (26, 23, 24) {real, imag} */,
  {32'h408bbaec, 32'h3fb75de9} /* (26, 23, 23) {real, imag} */,
  {32'hbe867f2b, 32'h3e363727} /* (26, 23, 22) {real, imag} */,
  {32'h3e0d6009, 32'hbff3ecf1} /* (26, 23, 21) {real, imag} */,
  {32'h3fee31c3, 32'h3e585e73} /* (26, 23, 20) {real, imag} */,
  {32'h3fd8c8d7, 32'hbfad7993} /* (26, 23, 19) {real, imag} */,
  {32'h3d2837fd, 32'h40653f65} /* (26, 23, 18) {real, imag} */,
  {32'h40116019, 32'hbeb4dd5c} /* (26, 23, 17) {real, imag} */,
  {32'h3f21a260, 32'hbec5552d} /* (26, 23, 16) {real, imag} */,
  {32'h3f880573, 32'hbfa25030} /* (26, 23, 15) {real, imag} */,
  {32'h3eea3c57, 32'h3f70ced5} /* (26, 23, 14) {real, imag} */,
  {32'hbf310ad0, 32'h400259e5} /* (26, 23, 13) {real, imag} */,
  {32'hbfe18918, 32'hc00dfee2} /* (26, 23, 12) {real, imag} */,
  {32'h3f27e291, 32'h3fb72aab} /* (26, 23, 11) {real, imag} */,
  {32'hc05120f2, 32'h3f528d3b} /* (26, 23, 10) {real, imag} */,
  {32'h3f9745db, 32'h3ee3b0ea} /* (26, 23, 9) {real, imag} */,
  {32'h404e8bf4, 32'hbe4c9b3b} /* (26, 23, 8) {real, imag} */,
  {32'h3f5086da, 32'hc0886732} /* (26, 23, 7) {real, imag} */,
  {32'h3f41c6dd, 32'hbf0010b3} /* (26, 23, 6) {real, imag} */,
  {32'h4050453b, 32'hbfc32053} /* (26, 23, 5) {real, imag} */,
  {32'hbf41ef51, 32'hbda394f7} /* (26, 23, 4) {real, imag} */,
  {32'hc0923c50, 32'hc007525c} /* (26, 23, 3) {real, imag} */,
  {32'hbd522cc1, 32'h40876fdc} /* (26, 23, 2) {real, imag} */,
  {32'hbf9dd291, 32'hbffc7194} /* (26, 23, 1) {real, imag} */,
  {32'hbe992be7, 32'hc0e18d71} /* (26, 23, 0) {real, imag} */,
  {32'h3ef6d77d, 32'hc0017ade} /* (26, 22, 31) {real, imag} */,
  {32'hbea63c9a, 32'h3dfa37a3} /* (26, 22, 30) {real, imag} */,
  {32'hbd03211b, 32'hbf996a0a} /* (26, 22, 29) {real, imag} */,
  {32'h40811e0a, 32'hbf68e049} /* (26, 22, 28) {real, imag} */,
  {32'h3f7bcbec, 32'h4044e55c} /* (26, 22, 27) {real, imag} */,
  {32'h4013b9a3, 32'hc03fcedf} /* (26, 22, 26) {real, imag} */,
  {32'hbfe0a6a8, 32'hbf9a4e30} /* (26, 22, 25) {real, imag} */,
  {32'h3f85db20, 32'hc001ed28} /* (26, 22, 24) {real, imag} */,
  {32'hbf82f6c9, 32'h4023aaca} /* (26, 22, 23) {real, imag} */,
  {32'h3f1d23ec, 32'h3e277789} /* (26, 22, 22) {real, imag} */,
  {32'hc0774731, 32'hc02ce653} /* (26, 22, 21) {real, imag} */,
  {32'hbfd900c7, 32'h40181ce5} /* (26, 22, 20) {real, imag} */,
  {32'h40432b93, 32'hbfbc4587} /* (26, 22, 19) {real, imag} */,
  {32'hc03ff4a9, 32'hc00476b6} /* (26, 22, 18) {real, imag} */,
  {32'hbeb42c24, 32'h3f465244} /* (26, 22, 17) {real, imag} */,
  {32'h3f44890e, 32'hbdbaa56c} /* (26, 22, 16) {real, imag} */,
  {32'h3f5d68e8, 32'hc06cd765} /* (26, 22, 15) {real, imag} */,
  {32'h3f40c29a, 32'h3cd04858} /* (26, 22, 14) {real, imag} */,
  {32'hbf2bdd08, 32'h4005e02f} /* (26, 22, 13) {real, imag} */,
  {32'hbf5e6c0d, 32'h400eb868} /* (26, 22, 12) {real, imag} */,
  {32'hbf817183, 32'h3ff27ea5} /* (26, 22, 11) {real, imag} */,
  {32'h3fe1ddfc, 32'hc05075b9} /* (26, 22, 10) {real, imag} */,
  {32'h3fa6e25a, 32'hbfe1ebed} /* (26, 22, 9) {real, imag} */,
  {32'h3c757c37, 32'h4005b9ef} /* (26, 22, 8) {real, imag} */,
  {32'hc0367c75, 32'hbf969aed} /* (26, 22, 7) {real, imag} */,
  {32'hbfd7ade7, 32'h3f791533} /* (26, 22, 6) {real, imag} */,
  {32'hbf90ba6f, 32'hc02edf8f} /* (26, 22, 5) {real, imag} */,
  {32'hbf9400ea, 32'h401af297} /* (26, 22, 4) {real, imag} */,
  {32'hc03d4a07, 32'hbf5b3529} /* (26, 22, 3) {real, imag} */,
  {32'h3f23cb6d, 32'hbf3fed04} /* (26, 22, 2) {real, imag} */,
  {32'hbf8785c5, 32'hc011c163} /* (26, 22, 1) {real, imag} */,
  {32'h3f6e59db, 32'h4004ea7d} /* (26, 22, 0) {real, imag} */,
  {32'hbf038ff5, 32'hbf2a517b} /* (26, 21, 31) {real, imag} */,
  {32'h40505a04, 32'hbfc20c6f} /* (26, 21, 30) {real, imag} */,
  {32'h3f9d2159, 32'h40254345} /* (26, 21, 29) {real, imag} */,
  {32'hbfe3986a, 32'hbf498b18} /* (26, 21, 28) {real, imag} */,
  {32'h3ebe83b6, 32'hbfe378dd} /* (26, 21, 27) {real, imag} */,
  {32'h3f558e34, 32'hbfbbc2e2} /* (26, 21, 26) {real, imag} */,
  {32'hc040561c, 32'h40076d76} /* (26, 21, 25) {real, imag} */,
  {32'hbf777948, 32'hbf2aa832} /* (26, 21, 24) {real, imag} */,
  {32'h3ddf5117, 32'h3f69f1b6} /* (26, 21, 23) {real, imag} */,
  {32'hbf4ae3ad, 32'h3fb35790} /* (26, 21, 22) {real, imag} */,
  {32'hbeb01961, 32'hbf93bdc1} /* (26, 21, 21) {real, imag} */,
  {32'h3fc2aecf, 32'hbfd21616} /* (26, 21, 20) {real, imag} */,
  {32'hbeaa298a, 32'hc00c538c} /* (26, 21, 19) {real, imag} */,
  {32'hbde40550, 32'hbfc52922} /* (26, 21, 18) {real, imag} */,
  {32'h402e4454, 32'h3e26c7c2} /* (26, 21, 17) {real, imag} */,
  {32'hbe73cdbf, 32'hc009f769} /* (26, 21, 16) {real, imag} */,
  {32'hbf8cea31, 32'h4023b7d8} /* (26, 21, 15) {real, imag} */,
  {32'h3f691425, 32'hc0212d42} /* (26, 21, 14) {real, imag} */,
  {32'h3fa32567, 32'h3f77df1b} /* (26, 21, 13) {real, imag} */,
  {32'hbfd371f0, 32'hbfeb0f70} /* (26, 21, 12) {real, imag} */,
  {32'hc0462074, 32'h3fb099f6} /* (26, 21, 11) {real, imag} */,
  {32'h3f7eadef, 32'h4026a3f6} /* (26, 21, 10) {real, imag} */,
  {32'h3f8d18a0, 32'hbfaf40de} /* (26, 21, 9) {real, imag} */,
  {32'h3ff643f7, 32'hc00149fe} /* (26, 21, 8) {real, imag} */,
  {32'hc0118f2e, 32'hc029e430} /* (26, 21, 7) {real, imag} */,
  {32'h3fd8b5e3, 32'h408ff45e} /* (26, 21, 6) {real, imag} */,
  {32'hc08830e8, 32'h3f9cb904} /* (26, 21, 5) {real, imag} */,
  {32'hbf42ba99, 32'hbfaac074} /* (26, 21, 4) {real, imag} */,
  {32'h3ead7971, 32'hbd8bf1b2} /* (26, 21, 3) {real, imag} */,
  {32'h3f192d92, 32'h40263abf} /* (26, 21, 2) {real, imag} */,
  {32'h3eee10cd, 32'h40627459} /* (26, 21, 1) {real, imag} */,
  {32'h3fe4870c, 32'hc008d44d} /* (26, 21, 0) {real, imag} */,
  {32'hc00c9537, 32'h3f298ab3} /* (26, 20, 31) {real, imag} */,
  {32'h3f4c1ddd, 32'hbec5d8af} /* (26, 20, 30) {real, imag} */,
  {32'hbddc0b06, 32'hbdb7873a} /* (26, 20, 29) {real, imag} */,
  {32'hc0058252, 32'h3f3c84f8} /* (26, 20, 28) {real, imag} */,
  {32'h403c5d32, 32'hbe8f7e59} /* (26, 20, 27) {real, imag} */,
  {32'hbfbce0c3, 32'h3f006f9b} /* (26, 20, 26) {real, imag} */,
  {32'hbf073c36, 32'hc0039a42} /* (26, 20, 25) {real, imag} */,
  {32'hbf2e173e, 32'hbd2ae7eb} /* (26, 20, 24) {real, imag} */,
  {32'h3ebc2b87, 32'h3e7bfba7} /* (26, 20, 23) {real, imag} */,
  {32'h3f092773, 32'h4081fccf} /* (26, 20, 22) {real, imag} */,
  {32'h3fdbeaef, 32'hbfc560e4} /* (26, 20, 21) {real, imag} */,
  {32'hbf6318af, 32'hbf913d9f} /* (26, 20, 20) {real, imag} */,
  {32'h401195aa, 32'h3fa1f89e} /* (26, 20, 19) {real, imag} */,
  {32'hbea2cd98, 32'hbd9752d2} /* (26, 20, 18) {real, imag} */,
  {32'h3daf6fd4, 32'hbf39d966} /* (26, 20, 17) {real, imag} */,
  {32'hbf53b9e7, 32'hbdf1a81f} /* (26, 20, 16) {real, imag} */,
  {32'hbedba813, 32'hc001d1fa} /* (26, 20, 15) {real, imag} */,
  {32'h3fa2108f, 32'hc009ca51} /* (26, 20, 14) {real, imag} */,
  {32'h4038b87a, 32'hc00397ff} /* (26, 20, 13) {real, imag} */,
  {32'h3f922ec0, 32'hbe8480ce} /* (26, 20, 12) {real, imag} */,
  {32'hbf7df7b5, 32'h3ec2286f} /* (26, 20, 11) {real, imag} */,
  {32'h403a7efc, 32'hbfa8f06d} /* (26, 20, 10) {real, imag} */,
  {32'h3fcbc3ec, 32'h3e58ce91} /* (26, 20, 9) {real, imag} */,
  {32'h3fc3012f, 32'h3f9aac2c} /* (26, 20, 8) {real, imag} */,
  {32'h3fc7e1ac, 32'hc057a324} /* (26, 20, 7) {real, imag} */,
  {32'h3f72289c, 32'h401fb4d1} /* (26, 20, 6) {real, imag} */,
  {32'h3fa9ca0f, 32'hbf76d525} /* (26, 20, 5) {real, imag} */,
  {32'h3df04810, 32'hbfcd5b49} /* (26, 20, 4) {real, imag} */,
  {32'hbf6d6874, 32'h3e60f095} /* (26, 20, 3) {real, imag} */,
  {32'hc060e4bc, 32'h3fd6b9b0} /* (26, 20, 2) {real, imag} */,
  {32'hbfc0440b, 32'hbeabe591} /* (26, 20, 1) {real, imag} */,
  {32'hbfceacd1, 32'h3f25738f} /* (26, 20, 0) {real, imag} */,
  {32'h3e9be9d1, 32'h4016e70f} /* (26, 19, 31) {real, imag} */,
  {32'hbff8bdfd, 32'h3e058189} /* (26, 19, 30) {real, imag} */,
  {32'hc002fd50, 32'h3ea51556} /* (26, 19, 29) {real, imag} */,
  {32'h40179cde, 32'hbec6d125} /* (26, 19, 28) {real, imag} */,
  {32'hc0381fc7, 32'h3fd8b0af} /* (26, 19, 27) {real, imag} */,
  {32'hbf683461, 32'hc00f1574} /* (26, 19, 26) {real, imag} */,
  {32'hc0320e5d, 32'h4006b8d9} /* (26, 19, 25) {real, imag} */,
  {32'h3f290e11, 32'hbfce0f40} /* (26, 19, 24) {real, imag} */,
  {32'h3f125029, 32'h3e612b79} /* (26, 19, 23) {real, imag} */,
  {32'hbe3365d9, 32'hbffde375} /* (26, 19, 22) {real, imag} */,
  {32'hbf715124, 32'hbe29a128} /* (26, 19, 21) {real, imag} */,
  {32'hc011d3c7, 32'h401761e4} /* (26, 19, 20) {real, imag} */,
  {32'h3f83b336, 32'h3fd65d88} /* (26, 19, 19) {real, imag} */,
  {32'h3fda6630, 32'hc0c13e60} /* (26, 19, 18) {real, imag} */,
  {32'h3f3916c9, 32'h401029ac} /* (26, 19, 17) {real, imag} */,
  {32'hbebd3ea8, 32'h3fe2f582} /* (26, 19, 16) {real, imag} */,
  {32'h3f1c93c8, 32'hbdf462de} /* (26, 19, 15) {real, imag} */,
  {32'h3fb7e5a6, 32'hbf0bcfed} /* (26, 19, 14) {real, imag} */,
  {32'hc04a8a81, 32'h3f679101} /* (26, 19, 13) {real, imag} */,
  {32'h3f381e14, 32'h3fec833a} /* (26, 19, 12) {real, imag} */,
  {32'h3fc9481e, 32'hc00c3ed6} /* (26, 19, 11) {real, imag} */,
  {32'hbde94372, 32'hbefe1bfb} /* (26, 19, 10) {real, imag} */,
  {32'h3efe2e66, 32'h3feecee2} /* (26, 19, 9) {real, imag} */,
  {32'h3f3a2df7, 32'h3e0db93a} /* (26, 19, 8) {real, imag} */,
  {32'hbcade284, 32'h3f55eb01} /* (26, 19, 7) {real, imag} */,
  {32'hc0276e1c, 32'h3fb14633} /* (26, 19, 6) {real, imag} */,
  {32'h3f9c4bc2, 32'h3fcb2067} /* (26, 19, 5) {real, imag} */,
  {32'h3e2a8c3b, 32'h3f660c32} /* (26, 19, 4) {real, imag} */,
  {32'h3ff77fbe, 32'h3d812b2b} /* (26, 19, 3) {real, imag} */,
  {32'hbe76248d, 32'hbf7b9ad3} /* (26, 19, 2) {real, imag} */,
  {32'h401ca526, 32'h40376a08} /* (26, 19, 1) {real, imag} */,
  {32'hbe2aea41, 32'h3f5e9988} /* (26, 19, 0) {real, imag} */,
  {32'hbef688cf, 32'h3ef2ee15} /* (26, 18, 31) {real, imag} */,
  {32'h3fc2b17d, 32'hbf4ea1a1} /* (26, 18, 30) {real, imag} */,
  {32'h3f400449, 32'h3eb77228} /* (26, 18, 29) {real, imag} */,
  {32'hbf349af8, 32'hbdf6a3ac} /* (26, 18, 28) {real, imag} */,
  {32'h3fa69792, 32'hc04a0da1} /* (26, 18, 27) {real, imag} */,
  {32'hc033066e, 32'hbf55ecec} /* (26, 18, 26) {real, imag} */,
  {32'h3f448e4d, 32'h3f0b3899} /* (26, 18, 25) {real, imag} */,
  {32'hbeba69d1, 32'hc02da327} /* (26, 18, 24) {real, imag} */,
  {32'h3fbc7d27, 32'hbf2abefe} /* (26, 18, 23) {real, imag} */,
  {32'h3f981212, 32'hbfcbf117} /* (26, 18, 22) {real, imag} */,
  {32'hbf68e93a, 32'hbf6da19f} /* (26, 18, 21) {real, imag} */,
  {32'hbf7709fa, 32'hbf81690c} /* (26, 18, 20) {real, imag} */,
  {32'hbf4b0c1f, 32'hbf5eaaa8} /* (26, 18, 19) {real, imag} */,
  {32'h40071fb9, 32'hbf7ee161} /* (26, 18, 18) {real, imag} */,
  {32'hbeb2e298, 32'h3f87adff} /* (26, 18, 17) {real, imag} */,
  {32'hbf3e5208, 32'hbfb33f8a} /* (26, 18, 16) {real, imag} */,
  {32'h3f0b1f49, 32'hbf965de3} /* (26, 18, 15) {real, imag} */,
  {32'hbfb52932, 32'h4020bf4e} /* (26, 18, 14) {real, imag} */,
  {32'hc00eea61, 32'h3faa7d5e} /* (26, 18, 13) {real, imag} */,
  {32'hbfe977f1, 32'h3fb125c6} /* (26, 18, 12) {real, imag} */,
  {32'h3f1b2bc9, 32'hc029c36b} /* (26, 18, 11) {real, imag} */,
  {32'hbf9439b6, 32'h3f183f97} /* (26, 18, 10) {real, imag} */,
  {32'h3f952fa4, 32'h3fdf0b84} /* (26, 18, 9) {real, imag} */,
  {32'hc03b5feb, 32'h3fcc43e4} /* (26, 18, 8) {real, imag} */,
  {32'hbf2fba6f, 32'h3e0f1b6d} /* (26, 18, 7) {real, imag} */,
  {32'hbd1fe17a, 32'hc04c42a4} /* (26, 18, 6) {real, imag} */,
  {32'hbec1a9af, 32'hbf5bf4b6} /* (26, 18, 5) {real, imag} */,
  {32'hbd1ab65e, 32'hbf803288} /* (26, 18, 4) {real, imag} */,
  {32'hbf29fe59, 32'hbe89bcc9} /* (26, 18, 3) {real, imag} */,
  {32'hbe55e0ee, 32'hc00051b0} /* (26, 18, 2) {real, imag} */,
  {32'hc028ee9c, 32'h3f6561e9} /* (26, 18, 1) {real, imag} */,
  {32'hc00b42a1, 32'hbff6ec47} /* (26, 18, 0) {real, imag} */,
  {32'hbf5982d9, 32'h3f570e0c} /* (26, 17, 31) {real, imag} */,
  {32'hbd504e96, 32'hbead53e2} /* (26, 17, 30) {real, imag} */,
  {32'h40319c8e, 32'hbdd2aa9a} /* (26, 17, 29) {real, imag} */,
  {32'hbfe33081, 32'hbfddd7f2} /* (26, 17, 28) {real, imag} */,
  {32'h3cc4560f, 32'h3fc64234} /* (26, 17, 27) {real, imag} */,
  {32'hbdc57d2f, 32'hbf38738e} /* (26, 17, 26) {real, imag} */,
  {32'h3f45cc8a, 32'h4000760d} /* (26, 17, 25) {real, imag} */,
  {32'hbfbac3f3, 32'h3fb89c13} /* (26, 17, 24) {real, imag} */,
  {32'hc02d3103, 32'hbfffccb4} /* (26, 17, 23) {real, imag} */,
  {32'h3fcdba1b, 32'hc02c493d} /* (26, 17, 22) {real, imag} */,
  {32'hc00440b5, 32'hbdda8ea2} /* (26, 17, 21) {real, imag} */,
  {32'h3ea2aa1a, 32'hbd94c268} /* (26, 17, 20) {real, imag} */,
  {32'h3f3d1716, 32'hbf9e4fbe} /* (26, 17, 19) {real, imag} */,
  {32'hbf2da467, 32'h3f7620fd} /* (26, 17, 18) {real, imag} */,
  {32'h3d0b1cbf, 32'h3fb77db6} /* (26, 17, 17) {real, imag} */,
  {32'h3f932be9, 32'hbf409762} /* (26, 17, 16) {real, imag} */,
  {32'hbf3acb9a, 32'hbe65a00f} /* (26, 17, 15) {real, imag} */,
  {32'hc00fa6b2, 32'h3f37226b} /* (26, 17, 14) {real, imag} */,
  {32'hbe94eac7, 32'hc010c9d9} /* (26, 17, 13) {real, imag} */,
  {32'hbe7f5604, 32'hbd8302ac} /* (26, 17, 12) {real, imag} */,
  {32'hc0341d61, 32'h3ebdc9d7} /* (26, 17, 11) {real, imag} */,
  {32'hbef5bbac, 32'h3f6d7ac8} /* (26, 17, 10) {real, imag} */,
  {32'h3e94d305, 32'h3f45c660} /* (26, 17, 9) {real, imag} */,
  {32'hc04217eb, 32'h400eb1b3} /* (26, 17, 8) {real, imag} */,
  {32'h3fa0197c, 32'h4015222a} /* (26, 17, 7) {real, imag} */,
  {32'h3fbfb7a8, 32'hbfc9581e} /* (26, 17, 6) {real, imag} */,
  {32'hbfc2348e, 32'h3fdaac1e} /* (26, 17, 5) {real, imag} */,
  {32'h3e3837b7, 32'hbf9e54db} /* (26, 17, 4) {real, imag} */,
  {32'h3e6f0adc, 32'h400d5533} /* (26, 17, 3) {real, imag} */,
  {32'h3f61a2ad, 32'hbf8dbb7f} /* (26, 17, 2) {real, imag} */,
  {32'h3f7d0699, 32'h3fc13c5e} /* (26, 17, 1) {real, imag} */,
  {32'h401fd2ae, 32'hbf6d758d} /* (26, 17, 0) {real, imag} */,
  {32'h3b086186, 32'h3f831dc3} /* (26, 16, 31) {real, imag} */,
  {32'h3dd3e79e, 32'hbf763cb5} /* (26, 16, 30) {real, imag} */,
  {32'h3f1efb02, 32'h3f0e6195} /* (26, 16, 29) {real, imag} */,
  {32'hbffb8f4f, 32'hbdc571fa} /* (26, 16, 28) {real, imag} */,
  {32'hbf680666, 32'hbfbb4748} /* (26, 16, 27) {real, imag} */,
  {32'hbec1dbcb, 32'h3f78dbbb} /* (26, 16, 26) {real, imag} */,
  {32'h3e1e94ae, 32'h3ea21f18} /* (26, 16, 25) {real, imag} */,
  {32'hbe1ef30b, 32'h3e16fff3} /* (26, 16, 24) {real, imag} */,
  {32'hbf694e32, 32'hbf8be399} /* (26, 16, 23) {real, imag} */,
  {32'hbde653c5, 32'h3ffa72ea} /* (26, 16, 22) {real, imag} */,
  {32'h3e894f2a, 32'hbeeb3811} /* (26, 16, 21) {real, imag} */,
  {32'hbf8f14e2, 32'hbfafb8dd} /* (26, 16, 20) {real, imag} */,
  {32'h3fb39c2a, 32'h3f513fd9} /* (26, 16, 19) {real, imag} */,
  {32'h3fa611b0, 32'h40313ba3} /* (26, 16, 18) {real, imag} */,
  {32'hbecbcf9d, 32'h3f1ce9d1} /* (26, 16, 17) {real, imag} */,
  {32'h3e6d240d, 32'h3f93f0e0} /* (26, 16, 16) {real, imag} */,
  {32'h4008dee3, 32'hbf87d890} /* (26, 16, 15) {real, imag} */,
  {32'h3fc366ef, 32'h3fe4bef3} /* (26, 16, 14) {real, imag} */,
  {32'h3f8226ca, 32'hbeac4c09} /* (26, 16, 13) {real, imag} */,
  {32'h3fd8bb47, 32'hbe24ed12} /* (26, 16, 12) {real, imag} */,
  {32'h3eee18f4, 32'hbfa1bb8f} /* (26, 16, 11) {real, imag} */,
  {32'h3e9a932f, 32'hbd11b5bd} /* (26, 16, 10) {real, imag} */,
  {32'h3e8794ef, 32'hbd5d73cc} /* (26, 16, 9) {real, imag} */,
  {32'h3f68e110, 32'h3f77f78a} /* (26, 16, 8) {real, imag} */,
  {32'h3e8ce073, 32'h3f21d4f5} /* (26, 16, 7) {real, imag} */,
  {32'hbeffb8fe, 32'hbf9a68cb} /* (26, 16, 6) {real, imag} */,
  {32'hbf4567b9, 32'h3f7bb584} /* (26, 16, 5) {real, imag} */,
  {32'hbf419a01, 32'h3de68fde} /* (26, 16, 4) {real, imag} */,
  {32'h3f7f6698, 32'hbed273fc} /* (26, 16, 3) {real, imag} */,
  {32'h3f52bab8, 32'hbee2161a} /* (26, 16, 2) {real, imag} */,
  {32'h3f04af00, 32'h3f234812} /* (26, 16, 1) {real, imag} */,
  {32'h3ed7c19c, 32'hbebed2fa} /* (26, 16, 0) {real, imag} */,
  {32'hbf119c35, 32'hbe265ed7} /* (26, 15, 31) {real, imag} */,
  {32'hc0873980, 32'hbf1f1471} /* (26, 15, 30) {real, imag} */,
  {32'h3f994a48, 32'hbffe731f} /* (26, 15, 29) {real, imag} */,
  {32'h3fe1e99a, 32'h3e1c870c} /* (26, 15, 28) {real, imag} */,
  {32'hbfb069b5, 32'h3f4e7655} /* (26, 15, 27) {real, imag} */,
  {32'hbea643d8, 32'hbf62c195} /* (26, 15, 26) {real, imag} */,
  {32'hbfb71c6f, 32'hbfc984f0} /* (26, 15, 25) {real, imag} */,
  {32'hbf380e44, 32'h3fe63b13} /* (26, 15, 24) {real, imag} */,
  {32'h3dbebc79, 32'h3f2d760d} /* (26, 15, 23) {real, imag} */,
  {32'hc02a7f44, 32'h4009b310} /* (26, 15, 22) {real, imag} */,
  {32'h3b7ae2f8, 32'hbe251ab8} /* (26, 15, 21) {real, imag} */,
  {32'hbe8942a7, 32'hbf5ebf31} /* (26, 15, 20) {real, imag} */,
  {32'hbfbbddab, 32'h3fae14a1} /* (26, 15, 19) {real, imag} */,
  {32'h3fc56e47, 32'h3f13f363} /* (26, 15, 18) {real, imag} */,
  {32'h4004be78, 32'h3f29917d} /* (26, 15, 17) {real, imag} */,
  {32'hc054a131, 32'hbefdb083} /* (26, 15, 16) {real, imag} */,
  {32'hbe89eddc, 32'h3faf980b} /* (26, 15, 15) {real, imag} */,
  {32'h3e98cc4c, 32'hc00fb219} /* (26, 15, 14) {real, imag} */,
  {32'hbf88480a, 32'h3fe22591} /* (26, 15, 13) {real, imag} */,
  {32'h3f9baa6a, 32'h3f608416} /* (26, 15, 12) {real, imag} */,
  {32'hbf2edd01, 32'hbfd6cb25} /* (26, 15, 11) {real, imag} */,
  {32'hbf6ba6b5, 32'h3ad3ba65} /* (26, 15, 10) {real, imag} */,
  {32'h3fc6191b, 32'hbf3ee991} /* (26, 15, 9) {real, imag} */,
  {32'h3d5f333c, 32'hbf7e0439} /* (26, 15, 8) {real, imag} */,
  {32'h3e998e6b, 32'hbf417655} /* (26, 15, 7) {real, imag} */,
  {32'hc015095b, 32'h3f925327} /* (26, 15, 6) {real, imag} */,
  {32'hbf8829d2, 32'h3fa5aee1} /* (26, 15, 5) {real, imag} */,
  {32'hbfb273c1, 32'hbfa061b2} /* (26, 15, 4) {real, imag} */,
  {32'hbef575d9, 32'hbe44200e} /* (26, 15, 3) {real, imag} */,
  {32'h4042ac02, 32'hc0016be9} /* (26, 15, 2) {real, imag} */,
  {32'h3f2d8816, 32'hbe8a03c2} /* (26, 15, 1) {real, imag} */,
  {32'hbfecfbd8, 32'h3e519dbd} /* (26, 15, 0) {real, imag} */,
  {32'h3e9fd9d4, 32'hbfcc7d70} /* (26, 14, 31) {real, imag} */,
  {32'hbf042e7c, 32'hbeb00279} /* (26, 14, 30) {real, imag} */,
  {32'h3f5c2e80, 32'h4044a5aa} /* (26, 14, 29) {real, imag} */,
  {32'hc04bc63a, 32'hbedd9599} /* (26, 14, 28) {real, imag} */,
  {32'hbdd0a57f, 32'hbf6b59b7} /* (26, 14, 27) {real, imag} */,
  {32'h400fed4f, 32'hbfe8e88d} /* (26, 14, 26) {real, imag} */,
  {32'h402e623d, 32'hbf6587ef} /* (26, 14, 25) {real, imag} */,
  {32'h3c859e7c, 32'hbfcb151f} /* (26, 14, 24) {real, imag} */,
  {32'hbeccdaf9, 32'hbfd5014c} /* (26, 14, 23) {real, imag} */,
  {32'hc002c641, 32'hc030c47c} /* (26, 14, 22) {real, imag} */,
  {32'h3f5dd10c, 32'hbe4fb6ef} /* (26, 14, 21) {real, imag} */,
  {32'hbe8bfcd2, 32'h3f1892a1} /* (26, 14, 20) {real, imag} */,
  {32'h3ec39bca, 32'h3f3a903e} /* (26, 14, 19) {real, imag} */,
  {32'h3f92d421, 32'hbff79839} /* (26, 14, 18) {real, imag} */,
  {32'hc012f959, 32'hbe1ca029} /* (26, 14, 17) {real, imag} */,
  {32'hbf168a00, 32'hbe8c3c4a} /* (26, 14, 16) {real, imag} */,
  {32'hbf8038a0, 32'h3e927024} /* (26, 14, 15) {real, imag} */,
  {32'hc0380554, 32'h3dc6889f} /* (26, 14, 14) {real, imag} */,
  {32'h3f3d53f5, 32'h3fd908a5} /* (26, 14, 13) {real, imag} */,
  {32'hbf3072df, 32'h3ff79f13} /* (26, 14, 12) {real, imag} */,
  {32'hbf751d56, 32'hbf874a55} /* (26, 14, 11) {real, imag} */,
  {32'h3f4184eb, 32'h3f589325} /* (26, 14, 10) {real, imag} */,
  {32'hc0418428, 32'h3e785146} /* (26, 14, 9) {real, imag} */,
  {32'h3e667988, 32'hbf221834} /* (26, 14, 8) {real, imag} */,
  {32'h3e823620, 32'hbf5e191a} /* (26, 14, 7) {real, imag} */,
  {32'hbfea2f11, 32'h3fd49f8d} /* (26, 14, 6) {real, imag} */,
  {32'hbd4e43fd, 32'hbedb85ca} /* (26, 14, 5) {real, imag} */,
  {32'hbfe038f8, 32'hbfcae717} /* (26, 14, 4) {real, imag} */,
  {32'h3fd6cb8b, 32'hc02c5662} /* (26, 14, 3) {real, imag} */,
  {32'hbef06cb3, 32'hbea1860f} /* (26, 14, 2) {real, imag} */,
  {32'hc016bc65, 32'h3f24580e} /* (26, 14, 1) {real, imag} */,
  {32'h3de8868e, 32'h3f411ca4} /* (26, 14, 0) {real, imag} */,
  {32'hbf3da694, 32'hbc9e55a3} /* (26, 13, 31) {real, imag} */,
  {32'h3f994a12, 32'hbfacb539} /* (26, 13, 30) {real, imag} */,
  {32'hbfb9439c, 32'hbdf3b881} /* (26, 13, 29) {real, imag} */,
  {32'hbe89f65c, 32'h3fbff52f} /* (26, 13, 28) {real, imag} */,
  {32'h3fbe167c, 32'h3f6d150b} /* (26, 13, 27) {real, imag} */,
  {32'hbfc31db9, 32'hbf368514} /* (26, 13, 26) {real, imag} */,
  {32'hbf68c4d4, 32'h3eeb61bc} /* (26, 13, 25) {real, imag} */,
  {32'h3f378d9b, 32'hbf694958} /* (26, 13, 24) {real, imag} */,
  {32'h40594f19, 32'h3f8b6966} /* (26, 13, 23) {real, imag} */,
  {32'h402233c9, 32'h3fa6798a} /* (26, 13, 22) {real, imag} */,
  {32'hbf315308, 32'hbfdc900b} /* (26, 13, 21) {real, imag} */,
  {32'hc0458014, 32'h3d191575} /* (26, 13, 20) {real, imag} */,
  {32'hbfad80f7, 32'h3f118369} /* (26, 13, 19) {real, imag} */,
  {32'hbf94ee72, 32'h4023de1e} /* (26, 13, 18) {real, imag} */,
  {32'hc007c12f, 32'h3f8b1e37} /* (26, 13, 17) {real, imag} */,
  {32'h3e52b36e, 32'hbe5718ef} /* (26, 13, 16) {real, imag} */,
  {32'h3f8cdc49, 32'hbf0499d8} /* (26, 13, 15) {real, imag} */,
  {32'hbe1c8b0d, 32'hbfdb2093} /* (26, 13, 14) {real, imag} */,
  {32'h3fbe0ebf, 32'h40150fe5} /* (26, 13, 13) {real, imag} */,
  {32'h3ea3cff3, 32'h40039d5c} /* (26, 13, 12) {real, imag} */,
  {32'h3e89e04f, 32'h3febc93a} /* (26, 13, 11) {real, imag} */,
  {32'hbefe5eb5, 32'hbfa3afcb} /* (26, 13, 10) {real, imag} */,
  {32'hbfd5eb4f, 32'hbe8def72} /* (26, 13, 9) {real, imag} */,
  {32'h4004a7c4, 32'h3f428274} /* (26, 13, 8) {real, imag} */,
  {32'hc05b2eab, 32'h3f03ac26} /* (26, 13, 7) {real, imag} */,
  {32'hbfbb4055, 32'hbf42ea02} /* (26, 13, 6) {real, imag} */,
  {32'hbe8e7f84, 32'h3e1091c4} /* (26, 13, 5) {real, imag} */,
  {32'hbf9438be, 32'h3fb000d8} /* (26, 13, 4) {real, imag} */,
  {32'hbf8cbee6, 32'hbf3f4fcd} /* (26, 13, 3) {real, imag} */,
  {32'h3ed1cfe3, 32'h3fe88c4f} /* (26, 13, 2) {real, imag} */,
  {32'hbf7c1efb, 32'hc03c92b5} /* (26, 13, 1) {real, imag} */,
  {32'hbec3cee4, 32'h3fb5a5bb} /* (26, 13, 0) {real, imag} */,
  {32'h3eeb8d7b, 32'h3f7df4f2} /* (26, 12, 31) {real, imag} */,
  {32'h3f9ce3b0, 32'hbe981c9e} /* (26, 12, 30) {real, imag} */,
  {32'hbfddfd54, 32'hbfc2ffdd} /* (26, 12, 29) {real, imag} */,
  {32'hbfdf0616, 32'hc001c05f} /* (26, 12, 28) {real, imag} */,
  {32'hbf82dd7b, 32'h4002f799} /* (26, 12, 27) {real, imag} */,
  {32'hc008aa14, 32'hbf91df3a} /* (26, 12, 26) {real, imag} */,
  {32'h3d825cce, 32'h3f8f5a4a} /* (26, 12, 25) {real, imag} */,
  {32'hc01877bf, 32'hbf3c385d} /* (26, 12, 24) {real, imag} */,
  {32'h3fb38ddb, 32'h3fc51eba} /* (26, 12, 23) {real, imag} */,
  {32'h3fb3be00, 32'h3f9b6703} /* (26, 12, 22) {real, imag} */,
  {32'h40154f6e, 32'hbfff1eeb} /* (26, 12, 21) {real, imag} */,
  {32'hbff79a8c, 32'h3fb28dda} /* (26, 12, 20) {real, imag} */,
  {32'h4020e3fb, 32'h3f1444f3} /* (26, 12, 19) {real, imag} */,
  {32'hbddb1dda, 32'hbf952fc6} /* (26, 12, 18) {real, imag} */,
  {32'h3f9da5e2, 32'hc0201a49} /* (26, 12, 17) {real, imag} */,
  {32'hbf45f626, 32'hc017fc8b} /* (26, 12, 16) {real, imag} */,
  {32'hbd506d93, 32'hbe961172} /* (26, 12, 15) {real, imag} */,
  {32'hbecaf370, 32'hc0477a9b} /* (26, 12, 14) {real, imag} */,
  {32'h3f51acfb, 32'h3f8a2f8c} /* (26, 12, 13) {real, imag} */,
  {32'h4022e10d, 32'hbeeb1bcb} /* (26, 12, 12) {real, imag} */,
  {32'hbfb53590, 32'h3fb03673} /* (26, 12, 11) {real, imag} */,
  {32'h3fe7de0c, 32'h40285933} /* (26, 12, 10) {real, imag} */,
  {32'hbfe52051, 32'hbfc61a3c} /* (26, 12, 9) {real, imag} */,
  {32'h3ffaffac, 32'h407b025b} /* (26, 12, 8) {real, imag} */,
  {32'h3d41d6ca, 32'hbf1fa7fc} /* (26, 12, 7) {real, imag} */,
  {32'h3f1fddd5, 32'h3e9b97d1} /* (26, 12, 6) {real, imag} */,
  {32'hbe261fbd, 32'hbfc81b52} /* (26, 12, 5) {real, imag} */,
  {32'hbead4053, 32'h3f7c74ac} /* (26, 12, 4) {real, imag} */,
  {32'hbe265477, 32'h4000b218} /* (26, 12, 3) {real, imag} */,
  {32'h4037584a, 32'hc00c50b3} /* (26, 12, 2) {real, imag} */,
  {32'hbff2083c, 32'hbf882801} /* (26, 12, 1) {real, imag} */,
  {32'h3f1eb140, 32'hbfdce5da} /* (26, 12, 0) {real, imag} */,
  {32'hc0504d15, 32'hbf699093} /* (26, 11, 31) {real, imag} */,
  {32'h405766be, 32'h3f76d3c1} /* (26, 11, 30) {real, imag} */,
  {32'h3febaf6b, 32'h3f45c435} /* (26, 11, 29) {real, imag} */,
  {32'hbf9b2463, 32'h40117b88} /* (26, 11, 28) {real, imag} */,
  {32'hc02a5ef7, 32'hbe259fa9} /* (26, 11, 27) {real, imag} */,
  {32'hbfa97466, 32'hbea0b213} /* (26, 11, 26) {real, imag} */,
  {32'hbfea71ca, 32'h401f788f} /* (26, 11, 25) {real, imag} */,
  {32'h3fd5816e, 32'hbeed123c} /* (26, 11, 24) {real, imag} */,
  {32'h3f260b2b, 32'hbfdc5d6d} /* (26, 11, 23) {real, imag} */,
  {32'h3ec40b2f, 32'h3f5a5371} /* (26, 11, 22) {real, imag} */,
  {32'hbfb03abc, 32'hbfb8c295} /* (26, 11, 21) {real, imag} */,
  {32'hc031df7a, 32'h40129383} /* (26, 11, 20) {real, imag} */,
  {32'h3e9bdb81, 32'h403db982} /* (26, 11, 19) {real, imag} */,
  {32'hbf837a57, 32'hbfea750e} /* (26, 11, 18) {real, imag} */,
  {32'h3f98d877, 32'hbf4348c0} /* (26, 11, 17) {real, imag} */,
  {32'hbf145e60, 32'h3fa853ee} /* (26, 11, 16) {real, imag} */,
  {32'hbf6a35d3, 32'hc0372cbe} /* (26, 11, 15) {real, imag} */,
  {32'h3f49e1b2, 32'hbdbfcedd} /* (26, 11, 14) {real, imag} */,
  {32'hbfe83507, 32'h404e0f68} /* (26, 11, 13) {real, imag} */,
  {32'hbef7b444, 32'h4005ad85} /* (26, 11, 12) {real, imag} */,
  {32'hbfc9cd18, 32'hbff3fa22} /* (26, 11, 11) {real, imag} */,
  {32'hbf648dc7, 32'hbf62ed24} /* (26, 11, 10) {real, imag} */,
  {32'h3fa5731c, 32'h4095ddce} /* (26, 11, 9) {real, imag} */,
  {32'h3f94a603, 32'h40157fcb} /* (26, 11, 8) {real, imag} */,
  {32'h3e114a99, 32'hbfbe15a4} /* (26, 11, 7) {real, imag} */,
  {32'hc0124191, 32'hbfaf9aaa} /* (26, 11, 6) {real, imag} */,
  {32'hbec700ce, 32'h3ecf952d} /* (26, 11, 5) {real, imag} */,
  {32'h3f46f33d, 32'h40469c0e} /* (26, 11, 4) {real, imag} */,
  {32'hc0542366, 32'hbf28de7a} /* (26, 11, 3) {real, imag} */,
  {32'hbf430dea, 32'h3f01dec6} /* (26, 11, 2) {real, imag} */,
  {32'h3fac1e4d, 32'hbfc3bcaf} /* (26, 11, 1) {real, imag} */,
  {32'h3fbc6fcb, 32'h3e9b7369} /* (26, 11, 0) {real, imag} */,
  {32'hbf0d93fd, 32'hbf98ab3e} /* (26, 10, 31) {real, imag} */,
  {32'hc001c3de, 32'hbf7d26af} /* (26, 10, 30) {real, imag} */,
  {32'h4060e267, 32'hbdf5a5e9} /* (26, 10, 29) {real, imag} */,
  {32'hbe830664, 32'hbf3c6f5f} /* (26, 10, 28) {real, imag} */,
  {32'hbf93bbce, 32'hc05b1249} /* (26, 10, 27) {real, imag} */,
  {32'hbeddbd5c, 32'h40886e28} /* (26, 10, 26) {real, imag} */,
  {32'hbfdde9d8, 32'hc000d3ac} /* (26, 10, 25) {real, imag} */,
  {32'h40a1f8cd, 32'h3ff049d1} /* (26, 10, 24) {real, imag} */,
  {32'h3fbdd49b, 32'hbeefce2e} /* (26, 10, 23) {real, imag} */,
  {32'h3f0355dd, 32'hc0540987} /* (26, 10, 22) {real, imag} */,
  {32'hbf54d6b7, 32'h3e12720f} /* (26, 10, 21) {real, imag} */,
  {32'h3fcd4c26, 32'h3e6a4486} /* (26, 10, 20) {real, imag} */,
  {32'hbfad5b9d, 32'h3edc2110} /* (26, 10, 19) {real, imag} */,
  {32'h3f3863dc, 32'h3f336661} /* (26, 10, 18) {real, imag} */,
  {32'hbd9654fe, 32'h407163ec} /* (26, 10, 17) {real, imag} */,
  {32'h4020a0ac, 32'hbf2f3994} /* (26, 10, 16) {real, imag} */,
  {32'hbe1ea961, 32'hbea09db2} /* (26, 10, 15) {real, imag} */,
  {32'h3f2341e0, 32'hbfe6a8ba} /* (26, 10, 14) {real, imag} */,
  {32'hbf9a949f, 32'h3e4876b5} /* (26, 10, 13) {real, imag} */,
  {32'h3f750440, 32'h3ea9bfd9} /* (26, 10, 12) {real, imag} */,
  {32'hbf88875d, 32'hbf4292f7} /* (26, 10, 11) {real, imag} */,
  {32'hbfd56ea7, 32'h3f956477} /* (26, 10, 10) {real, imag} */,
  {32'hbeda8626, 32'h3fb9d406} /* (26, 10, 9) {real, imag} */,
  {32'h400b0f64, 32'hc0739fb8} /* (26, 10, 8) {real, imag} */,
  {32'hbcf63948, 32'h3f754171} /* (26, 10, 7) {real, imag} */,
  {32'h40716def, 32'h3f4953f4} /* (26, 10, 6) {real, imag} */,
  {32'h3f4694b8, 32'h3dd5e9ca} /* (26, 10, 5) {real, imag} */,
  {32'hbf6943a7, 32'h404a5ae7} /* (26, 10, 4) {real, imag} */,
  {32'h40367e17, 32'hc008ba84} /* (26, 10, 3) {real, imag} */,
  {32'hbf4d1a99, 32'hbf7538be} /* (26, 10, 2) {real, imag} */,
  {32'h3badb1f8, 32'h3e8c3066} /* (26, 10, 1) {real, imag} */,
  {32'hc01f3402, 32'h3fad6705} /* (26, 10, 0) {real, imag} */,
  {32'h3ee28613, 32'hbf087f8c} /* (26, 9, 31) {real, imag} */,
  {32'hbe1915bc, 32'h4067b636} /* (26, 9, 30) {real, imag} */,
  {32'hbd937977, 32'hc01adf6c} /* (26, 9, 29) {real, imag} */,
  {32'hc0136ac7, 32'hbf8f1f33} /* (26, 9, 28) {real, imag} */,
  {32'h3fc753bf, 32'hc04d25db} /* (26, 9, 27) {real, imag} */,
  {32'h3fce6dd5, 32'h3f26e700} /* (26, 9, 26) {real, imag} */,
  {32'h3e756695, 32'hc003afb6} /* (26, 9, 25) {real, imag} */,
  {32'hc0000a3f, 32'hbedbf650} /* (26, 9, 24) {real, imag} */,
  {32'hbf12af5a, 32'h3fdea230} /* (26, 9, 23) {real, imag} */,
  {32'h3fbab614, 32'h40480109} /* (26, 9, 22) {real, imag} */,
  {32'h3f529885, 32'hc04050e4} /* (26, 9, 21) {real, imag} */,
  {32'h3feb4767, 32'h3fd7dfd5} /* (26, 9, 20) {real, imag} */,
  {32'hbf38dd39, 32'hbf552b4c} /* (26, 9, 19) {real, imag} */,
  {32'hbf9f7053, 32'h40608809} /* (26, 9, 18) {real, imag} */,
  {32'hbf8d9d1e, 32'h3f2702f6} /* (26, 9, 17) {real, imag} */,
  {32'hc02e4054, 32'h402143eb} /* (26, 9, 16) {real, imag} */,
  {32'hbfc50b5b, 32'h3f23a92a} /* (26, 9, 15) {real, imag} */,
  {32'h3fd7ce5b, 32'hbfbbecc9} /* (26, 9, 14) {real, imag} */,
  {32'hbe8cf9b4, 32'h3f8fda35} /* (26, 9, 13) {real, imag} */,
  {32'hbfd1e4a7, 32'h3f21a59a} /* (26, 9, 12) {real, imag} */,
  {32'h3f80c8b6, 32'hc028c41a} /* (26, 9, 11) {real, imag} */,
  {32'hbf7055cd, 32'hc049c947} /* (26, 9, 10) {real, imag} */,
  {32'h40803e4d, 32'hbf499bfb} /* (26, 9, 9) {real, imag} */,
  {32'hbf0962c6, 32'h3fbc6d64} /* (26, 9, 8) {real, imag} */,
  {32'h4027aea4, 32'h3e293302} /* (26, 9, 7) {real, imag} */,
  {32'h3e328e84, 32'hc03e0b6e} /* (26, 9, 6) {real, imag} */,
  {32'h3f2c97a3, 32'h3f44e224} /* (26, 9, 5) {real, imag} */,
  {32'h3f886811, 32'h3f9a6cf2} /* (26, 9, 4) {real, imag} */,
  {32'h400684b4, 32'h3f0ed66a} /* (26, 9, 3) {real, imag} */,
  {32'h3ff5dcb1, 32'h3f93d682} /* (26, 9, 2) {real, imag} */,
  {32'h3f239512, 32'h3f1431b0} /* (26, 9, 1) {real, imag} */,
  {32'h3ff85cd1, 32'h3fd4b9ea} /* (26, 9, 0) {real, imag} */,
  {32'hbf8869c0, 32'h3f071898} /* (26, 8, 31) {real, imag} */,
  {32'hc095a5b9, 32'hc0b53167} /* (26, 8, 30) {real, imag} */,
  {32'hbe864b22, 32'h404cd06a} /* (26, 8, 29) {real, imag} */,
  {32'h3f848552, 32'hc004789d} /* (26, 8, 28) {real, imag} */,
  {32'hbf1906b4, 32'hbe69efba} /* (26, 8, 27) {real, imag} */,
  {32'hc026e30e, 32'h406d2f8c} /* (26, 8, 26) {real, imag} */,
  {32'h3ed166e2, 32'hbde0e576} /* (26, 8, 25) {real, imag} */,
  {32'hc078ac17, 32'h3db88990} /* (26, 8, 24) {real, imag} */,
  {32'h3f23844b, 32'h3f993ecc} /* (26, 8, 23) {real, imag} */,
  {32'h3fe70ff9, 32'hbfe9ae72} /* (26, 8, 22) {real, imag} */,
  {32'hbffee716, 32'h404139a2} /* (26, 8, 21) {real, imag} */,
  {32'h400e415c, 32'h3f86c9c9} /* (26, 8, 20) {real, imag} */,
  {32'hbf00c181, 32'hbf975ffe} /* (26, 8, 19) {real, imag} */,
  {32'h3f261578, 32'h40392448} /* (26, 8, 18) {real, imag} */,
  {32'h3e99dfcd, 32'hbf66cbaa} /* (26, 8, 17) {real, imag} */,
  {32'hbf8a5fc4, 32'hbfe1f0bd} /* (26, 8, 16) {real, imag} */,
  {32'hbf958a85, 32'h3fe752da} /* (26, 8, 15) {real, imag} */,
  {32'h4022367a, 32'h3fccff81} /* (26, 8, 14) {real, imag} */,
  {32'hc01bf957, 32'hbff54035} /* (26, 8, 13) {real, imag} */,
  {32'hbf62ea5c, 32'h3fa8f3a8} /* (26, 8, 12) {real, imag} */,
  {32'hbfb83cc4, 32'h401a48e8} /* (26, 8, 11) {real, imag} */,
  {32'hbf574be2, 32'h4053d54a} /* (26, 8, 10) {real, imag} */,
  {32'h403fbe8c, 32'h3fcccaeb} /* (26, 8, 9) {real, imag} */,
  {32'h3f81c9c4, 32'hbfab381c} /* (26, 8, 8) {real, imag} */,
  {32'h408fa381, 32'hbf89addc} /* (26, 8, 7) {real, imag} */,
  {32'h3f1f4db1, 32'h3e955dc6} /* (26, 8, 6) {real, imag} */,
  {32'hbfc31a28, 32'hbed2055a} /* (26, 8, 5) {real, imag} */,
  {32'h401d8a31, 32'h3f6df5a4} /* (26, 8, 4) {real, imag} */,
  {32'hbdd25c3e, 32'h4034d3d1} /* (26, 8, 3) {real, imag} */,
  {32'h402373d0, 32'h40d1d23a} /* (26, 8, 2) {real, imag} */,
  {32'hc0096f50, 32'hbfc23a5a} /* (26, 8, 1) {real, imag} */,
  {32'h407f328e, 32'hbfaf2abb} /* (26, 8, 0) {real, imag} */,
  {32'h4027f683, 32'h407608ee} /* (26, 7, 31) {real, imag} */,
  {32'hbfc6efe9, 32'h3f1144a0} /* (26, 7, 30) {real, imag} */,
  {32'h3d275fd6, 32'h3fd15348} /* (26, 7, 29) {real, imag} */,
  {32'hc033060b, 32'h402a7e9c} /* (26, 7, 28) {real, imag} */,
  {32'h3e973b18, 32'hc0345d9e} /* (26, 7, 27) {real, imag} */,
  {32'hbfa2af1e, 32'h3ff0162f} /* (26, 7, 26) {real, imag} */,
  {32'h3f85363c, 32'hbf8b8b2a} /* (26, 7, 25) {real, imag} */,
  {32'hc07deed9, 32'h3f4e598a} /* (26, 7, 24) {real, imag} */,
  {32'h3efda3c1, 32'h3e0ea315} /* (26, 7, 23) {real, imag} */,
  {32'hbeaa2038, 32'hbfea8e85} /* (26, 7, 22) {real, imag} */,
  {32'h401ccabe, 32'h4046ed68} /* (26, 7, 21) {real, imag} */,
  {32'hbfe46db5, 32'hbd929421} /* (26, 7, 20) {real, imag} */,
  {32'hbee93d12, 32'h400980f9} /* (26, 7, 19) {real, imag} */,
  {32'hc00d2086, 32'hbfd42523} /* (26, 7, 18) {real, imag} */,
  {32'h3f5a7ac4, 32'hbfc038d6} /* (26, 7, 17) {real, imag} */,
  {32'hbfb0151c, 32'hbfb39029} /* (26, 7, 16) {real, imag} */,
  {32'hbea016c8, 32'h40478830} /* (26, 7, 15) {real, imag} */,
  {32'hbdb19a6f, 32'h40330e6d} /* (26, 7, 14) {real, imag} */,
  {32'hbf3dd29c, 32'h3e388f19} /* (26, 7, 13) {real, imag} */,
  {32'h3f5666d1, 32'h3d1b18f0} /* (26, 7, 12) {real, imag} */,
  {32'h3ff73552, 32'hbf7ad227} /* (26, 7, 11) {real, imag} */,
  {32'hbffd035f, 32'hbee137d8} /* (26, 7, 10) {real, imag} */,
  {32'hbf168e53, 32'hbf09e990} /* (26, 7, 9) {real, imag} */,
  {32'h3f798c15, 32'hc03b54ca} /* (26, 7, 8) {real, imag} */,
  {32'hbea862c4, 32'h401958cb} /* (26, 7, 7) {real, imag} */,
  {32'hbf8b2221, 32'h4041ba8d} /* (26, 7, 6) {real, imag} */,
  {32'h3f4486d6, 32'hbeeebb07} /* (26, 7, 5) {real, imag} */,
  {32'h3f52f834, 32'hbeb1e40b} /* (26, 7, 4) {real, imag} */,
  {32'h3e0871a2, 32'hc0bccca5} /* (26, 7, 3) {real, imag} */,
  {32'hbebe0d19, 32'hbf7480b4} /* (26, 7, 2) {real, imag} */,
  {32'h4045a726, 32'h40602031} /* (26, 7, 1) {real, imag} */,
  {32'hbfd8c48a, 32'h403cca96} /* (26, 7, 0) {real, imag} */,
  {32'h4012668f, 32'h3f9f6f37} /* (26, 6, 31) {real, imag} */,
  {32'hc053b6dd, 32'hbe8e9dc6} /* (26, 6, 30) {real, imag} */,
  {32'h40bf994b, 32'h3d90861b} /* (26, 6, 29) {real, imag} */,
  {32'h3fa0d772, 32'hc07bbac4} /* (26, 6, 28) {real, imag} */,
  {32'h401e87aa, 32'hbe95b78d} /* (26, 6, 27) {real, imag} */,
  {32'h4082fd32, 32'hc02d521c} /* (26, 6, 26) {real, imag} */,
  {32'hbfe90737, 32'h40a0847b} /* (26, 6, 25) {real, imag} */,
  {32'hbfbe5913, 32'h3f4227f8} /* (26, 6, 24) {real, imag} */,
  {32'h3da34456, 32'hbe282ce2} /* (26, 6, 23) {real, imag} */,
  {32'hbff9459b, 32'h3f3452e9} /* (26, 6, 22) {real, imag} */,
  {32'h3fe46e25, 32'hbf2d2557} /* (26, 6, 21) {real, imag} */,
  {32'h3f15ae96, 32'h3f5e6dc9} /* (26, 6, 20) {real, imag} */,
  {32'hc01b84ee, 32'h3fa0909b} /* (26, 6, 19) {real, imag} */,
  {32'h3e2db08c, 32'h3fb1ade7} /* (26, 6, 18) {real, imag} */,
  {32'hbf334d4c, 32'h3d1d3416} /* (26, 6, 17) {real, imag} */,
  {32'h3fb1222c, 32'h3cccc8db} /* (26, 6, 16) {real, imag} */,
  {32'hbec67627, 32'hbf89ad34} /* (26, 6, 15) {real, imag} */,
  {32'h3f38befd, 32'h3ece0efa} /* (26, 6, 14) {real, imag} */,
  {32'hbfe51150, 32'hc08681b4} /* (26, 6, 13) {real, imag} */,
  {32'h3f51c390, 32'h3f8dfd1e} /* (26, 6, 12) {real, imag} */,
  {32'hbe98ff5f, 32'h3f3f18db} /* (26, 6, 11) {real, imag} */,
  {32'hc025a35b, 32'hbe779edb} /* (26, 6, 10) {real, imag} */,
  {32'h401a09d1, 32'hc0184347} /* (26, 6, 9) {real, imag} */,
  {32'h3e9c08aa, 32'hc080c27a} /* (26, 6, 8) {real, imag} */,
  {32'h400c246d, 32'h3f83a9ef} /* (26, 6, 7) {real, imag} */,
  {32'h3f2ea376, 32'hbfa68235} /* (26, 6, 6) {real, imag} */,
  {32'hbf512d37, 32'h3e9a2e06} /* (26, 6, 5) {real, imag} */,
  {32'hbeae2ceb, 32'h407267fd} /* (26, 6, 4) {real, imag} */,
  {32'hbf74c9ad, 32'hc07d73ba} /* (26, 6, 3) {real, imag} */,
  {32'hbf0cd021, 32'hbf657d6a} /* (26, 6, 2) {real, imag} */,
  {32'h407fd40c, 32'h40638119} /* (26, 6, 1) {real, imag} */,
  {32'h3f7bb9c8, 32'hc0b5e67e} /* (26, 6, 0) {real, imag} */,
  {32'hc041f344, 32'h4014fcb7} /* (26, 5, 31) {real, imag} */,
  {32'h3f6e1b5a, 32'hbe5ab591} /* (26, 5, 30) {real, imag} */,
  {32'hbfb3ae66, 32'hbf843f04} /* (26, 5, 29) {real, imag} */,
  {32'hc00edfc0, 32'h3f6a1740} /* (26, 5, 28) {real, imag} */,
  {32'h3e79dd38, 32'h40a0714f} /* (26, 5, 27) {real, imag} */,
  {32'h3eb8c134, 32'hbe9735b3} /* (26, 5, 26) {real, imag} */,
  {32'h3fdf2eaa, 32'hbe48e60c} /* (26, 5, 25) {real, imag} */,
  {32'hbea036cc, 32'h4023123b} /* (26, 5, 24) {real, imag} */,
  {32'h3f0045d0, 32'h4015d09b} /* (26, 5, 23) {real, imag} */,
  {32'hc04b7dc0, 32'hbf736c29} /* (26, 5, 22) {real, imag} */,
  {32'h3fcc51cc, 32'hbf57b106} /* (26, 5, 21) {real, imag} */,
  {32'h40955986, 32'hbfd4b328} /* (26, 5, 20) {real, imag} */,
  {32'hbfbb0383, 32'h3f907eeb} /* (26, 5, 19) {real, imag} */,
  {32'h3e5d6c82, 32'hbf9cbac6} /* (26, 5, 18) {real, imag} */,
  {32'hbf2523d3, 32'hbf9742c8} /* (26, 5, 17) {real, imag} */,
  {32'hbf810d47, 32'h3fc71d3d} /* (26, 5, 16) {real, imag} */,
  {32'hbe1db2ab, 32'hbe72821c} /* (26, 5, 15) {real, imag} */,
  {32'h3f1dc045, 32'hbf93c006} /* (26, 5, 14) {real, imag} */,
  {32'h3fb9b661, 32'h407d0247} /* (26, 5, 13) {real, imag} */,
  {32'h3fb997d7, 32'h3f844677} /* (26, 5, 12) {real, imag} */,
  {32'hbdc91340, 32'h3ec19f91} /* (26, 5, 11) {real, imag} */,
  {32'h40389e5d, 32'hbfb2d19e} /* (26, 5, 10) {real, imag} */,
  {32'h3d7939d4, 32'hbe5e9dd1} /* (26, 5, 9) {real, imag} */,
  {32'h40401b54, 32'h40316028} /* (26, 5, 8) {real, imag} */,
  {32'hc0400107, 32'hbf7dd6bc} /* (26, 5, 7) {real, imag} */,
  {32'h3e8f34e1, 32'hbec368d2} /* (26, 5, 6) {real, imag} */,
  {32'hbfa23f54, 32'hbe0533d9} /* (26, 5, 5) {real, imag} */,
  {32'hc08443cd, 32'h3f4cd1c0} /* (26, 5, 4) {real, imag} */,
  {32'hbeb7180a, 32'hbffc4edb} /* (26, 5, 3) {real, imag} */,
  {32'h409d49e0, 32'h4022b966} /* (26, 5, 2) {real, imag} */,
  {32'hbf6ef52d, 32'hc0015d19} /* (26, 5, 1) {real, imag} */,
  {32'h3de67127, 32'h4079fc0a} /* (26, 5, 0) {real, imag} */,
  {32'hc07e77d3, 32'hbfd00d29} /* (26, 4, 31) {real, imag} */,
  {32'h40a1d87e, 32'hc07236a8} /* (26, 4, 30) {real, imag} */,
  {32'h408f1c6c, 32'hbfe20139} /* (26, 4, 29) {real, imag} */,
  {32'h4053777a, 32'hbffbf9e4} /* (26, 4, 28) {real, imag} */,
  {32'h3bda0664, 32'h40530912} /* (26, 4, 27) {real, imag} */,
  {32'hbfb30897, 32'h40b5c00a} /* (26, 4, 26) {real, imag} */,
  {32'h40b3868f, 32'h3f85b8f8} /* (26, 4, 25) {real, imag} */,
  {32'h4020486b, 32'hbed47f04} /* (26, 4, 24) {real, imag} */,
  {32'h3f535b1a, 32'hbfe70b42} /* (26, 4, 23) {real, imag} */,
  {32'h3f09c873, 32'hbffae799} /* (26, 4, 22) {real, imag} */,
  {32'hc02638d0, 32'hc0117072} /* (26, 4, 21) {real, imag} */,
  {32'h402ef3a7, 32'h40596042} /* (26, 4, 20) {real, imag} */,
  {32'hbfdc5b77, 32'h40914cb2} /* (26, 4, 19) {real, imag} */,
  {32'h3fd0a438, 32'h3ea60d62} /* (26, 4, 18) {real, imag} */,
  {32'h3fd02a02, 32'h3ea72367} /* (26, 4, 17) {real, imag} */,
  {32'hbf36a517, 32'h3f82e1f2} /* (26, 4, 16) {real, imag} */,
  {32'hbfd23211, 32'h4021431c} /* (26, 4, 15) {real, imag} */,
  {32'h3f066a41, 32'h3eb30d74} /* (26, 4, 14) {real, imag} */,
  {32'hc05b30cf, 32'hbface9bf} /* (26, 4, 13) {real, imag} */,
  {32'h3ffdc406, 32'h3f86ba46} /* (26, 4, 12) {real, imag} */,
  {32'hbeaa11a7, 32'hbfded89e} /* (26, 4, 11) {real, imag} */,
  {32'h3e40b5f3, 32'hbf4596f1} /* (26, 4, 10) {real, imag} */,
  {32'hbf044f67, 32'h3f83aff5} /* (26, 4, 9) {real, imag} */,
  {32'h40549c5e, 32'h3f40ce57} /* (26, 4, 8) {real, imag} */,
  {32'h401ed6ed, 32'hc014be2c} /* (26, 4, 7) {real, imag} */,
  {32'hc09fcf94, 32'hbf33f96e} /* (26, 4, 6) {real, imag} */,
  {32'h4077529e, 32'hc0265fbf} /* (26, 4, 5) {real, imag} */,
  {32'h3f626f31, 32'h4034ec67} /* (26, 4, 4) {real, imag} */,
  {32'h40d347eb, 32'h408541d7} /* (26, 4, 3) {real, imag} */,
  {32'hc0ba8a74, 32'hbf012ec4} /* (26, 4, 2) {real, imag} */,
  {32'hc06e67b9, 32'h40868ee7} /* (26, 4, 1) {real, imag} */,
  {32'h3f37aa4c, 32'hbf173cee} /* (26, 4, 0) {real, imag} */,
  {32'h401b7bc4, 32'hbeca723c} /* (26, 3, 31) {real, imag} */,
  {32'hc022b852, 32'hc0dfdcd3} /* (26, 3, 30) {real, imag} */,
  {32'h4001e697, 32'hc0afb0e1} /* (26, 3, 29) {real, imag} */,
  {32'hc03d4aca, 32'h3ec1944f} /* (26, 3, 28) {real, imag} */,
  {32'hc01b69dc, 32'h40a82bd9} /* (26, 3, 27) {real, imag} */,
  {32'h3f709778, 32'hbfd681c6} /* (26, 3, 26) {real, imag} */,
  {32'h3fb0290b, 32'h3fa1b565} /* (26, 3, 25) {real, imag} */,
  {32'h40a79437, 32'hbee8172e} /* (26, 3, 24) {real, imag} */,
  {32'h3f36b948, 32'h3fc0772a} /* (26, 3, 23) {real, imag} */,
  {32'hbfd2946c, 32'hbe812f16} /* (26, 3, 22) {real, imag} */,
  {32'h3fabc9e5, 32'h40828371} /* (26, 3, 21) {real, imag} */,
  {32'h403ce0e8, 32'hbf67c354} /* (26, 3, 20) {real, imag} */,
  {32'hbfb456be, 32'hbf78a949} /* (26, 3, 19) {real, imag} */,
  {32'hbffbf68b, 32'hc02901b6} /* (26, 3, 18) {real, imag} */,
  {32'h3f3bbe94, 32'hbf5b9b76} /* (26, 3, 17) {real, imag} */,
  {32'h3f6657b6, 32'h3f344b98} /* (26, 3, 16) {real, imag} */,
  {32'h3f9673f1, 32'h3f581255} /* (26, 3, 15) {real, imag} */,
  {32'h401bc0c1, 32'hbf2745d1} /* (26, 3, 14) {real, imag} */,
  {32'h4055d242, 32'hbfb6c20f} /* (26, 3, 13) {real, imag} */,
  {32'h3ea2291c, 32'hc02461bd} /* (26, 3, 12) {real, imag} */,
  {32'h4058d8a9, 32'h407c653c} /* (26, 3, 11) {real, imag} */,
  {32'hbf6208d2, 32'h3f9a1052} /* (26, 3, 10) {real, imag} */,
  {32'hc055f41c, 32'h40405bf8} /* (26, 3, 9) {real, imag} */,
  {32'hbf351a67, 32'hc014e206} /* (26, 3, 8) {real, imag} */,
  {32'hc03840cd, 32'hbc486142} /* (26, 3, 7) {real, imag} */,
  {32'h3ed96380, 32'hc0084fcc} /* (26, 3, 6) {real, imag} */,
  {32'hbf001827, 32'h3ff5124b} /* (26, 3, 5) {real, imag} */,
  {32'hc0434c4d, 32'hbf9afad8} /* (26, 3, 4) {real, imag} */,
  {32'h40b9a660, 32'hbf98d99d} /* (26, 3, 3) {real, imag} */,
  {32'h401e6c9b, 32'hc0aebf2b} /* (26, 3, 2) {real, imag} */,
  {32'hbf9454f0, 32'h40e51da8} /* (26, 3, 1) {real, imag} */,
  {32'h40e2155e, 32'h412fc090} /* (26, 3, 0) {real, imag} */,
  {32'hc0ba9cbf, 32'hc029c230} /* (26, 2, 31) {real, imag} */,
  {32'h40d651aa, 32'h4107dc6a} /* (26, 2, 30) {real, imag} */,
  {32'hc01db557, 32'hc0da2d9c} /* (26, 2, 29) {real, imag} */,
  {32'h3ffeab76, 32'h40c06cc7} /* (26, 2, 28) {real, imag} */,
  {32'hc0a33c7a, 32'hc0934697} /* (26, 2, 27) {real, imag} */,
  {32'h3f48b696, 32'h40808286} /* (26, 2, 26) {real, imag} */,
  {32'h3eb1aeed, 32'h3eb6fe7b} /* (26, 2, 25) {real, imag} */,
  {32'h3fd048f8, 32'hc0298a85} /* (26, 2, 24) {real, imag} */,
  {32'h3f6acf5c, 32'hbc28fcd2} /* (26, 2, 23) {real, imag} */,
  {32'hc0891cb5, 32'h3fe84ce9} /* (26, 2, 22) {real, imag} */,
  {32'h3f0ce1e2, 32'hbdd00cf7} /* (26, 2, 21) {real, imag} */,
  {32'h3ea4bb1a, 32'h4017cd78} /* (26, 2, 20) {real, imag} */,
  {32'hbe2f8d37, 32'hbf437bba} /* (26, 2, 19) {real, imag} */,
  {32'hbca002e4, 32'h3e5e7e03} /* (26, 2, 18) {real, imag} */,
  {32'hbfd83313, 32'hbf8000fa} /* (26, 2, 17) {real, imag} */,
  {32'hbf0d0276, 32'h3ed022df} /* (26, 2, 16) {real, imag} */,
  {32'hbf84de0b, 32'h3ed6a8a5} /* (26, 2, 15) {real, imag} */,
  {32'hbf62826c, 32'h3ebb04c4} /* (26, 2, 14) {real, imag} */,
  {32'h3ec40815, 32'h4017bce9} /* (26, 2, 13) {real, imag} */,
  {32'hc0878c23, 32'hc02d828f} /* (26, 2, 12) {real, imag} */,
  {32'h3c7a18c9, 32'hbfa4a40e} /* (26, 2, 11) {real, imag} */,
  {32'hc01a7233, 32'hbc690f17} /* (26, 2, 10) {real, imag} */,
  {32'hc052e9b1, 32'h3faf5b92} /* (26, 2, 9) {real, imag} */,
  {32'h3dfd3081, 32'hc018b9de} /* (26, 2, 8) {real, imag} */,
  {32'hbe9604e8, 32'hbedb0737} /* (26, 2, 7) {real, imag} */,
  {32'hbff8d806, 32'h3f4e5b6f} /* (26, 2, 6) {real, imag} */,
  {32'h3ee4e156, 32'h3f799317} /* (26, 2, 5) {real, imag} */,
  {32'hc02c1aaa, 32'hc066b20a} /* (26, 2, 4) {real, imag} */,
  {32'h40a89385, 32'h3fa2fea4} /* (26, 2, 3) {real, imag} */,
  {32'h40b15230, 32'hbf8b6a49} /* (26, 2, 2) {real, imag} */,
  {32'h410ac75d, 32'hbfd4ec1e} /* (26, 2, 1) {real, imag} */,
  {32'hc0738015, 32'h3fb7635f} /* (26, 2, 0) {real, imag} */,
  {32'hbee9b043, 32'h3fe851d9} /* (26, 1, 31) {real, imag} */,
  {32'h40f09af1, 32'hc0bbb4a9} /* (26, 1, 30) {real, imag} */,
  {32'h3f29b795, 32'h41053939} /* (26, 1, 29) {real, imag} */,
  {32'hc0acfb26, 32'hc0f6dc31} /* (26, 1, 28) {real, imag} */,
  {32'h3fb9ab28, 32'hc008ef1a} /* (26, 1, 27) {real, imag} */,
  {32'hc02cc300, 32'h40666ca5} /* (26, 1, 26) {real, imag} */,
  {32'hc0035216, 32'hc042491f} /* (26, 1, 25) {real, imag} */,
  {32'h3f61a052, 32'h3f97bf82} /* (26, 1, 24) {real, imag} */,
  {32'h405c55c0, 32'hbffc686a} /* (26, 1, 23) {real, imag} */,
  {32'hbfda0198, 32'hbf08c799} /* (26, 1, 22) {real, imag} */,
  {32'hc031eeac, 32'hbde4d6c1} /* (26, 1, 21) {real, imag} */,
  {32'h405e2c8c, 32'hc00d2ddd} /* (26, 1, 20) {real, imag} */,
  {32'hbf6273a7, 32'hbf5f23dd} /* (26, 1, 19) {real, imag} */,
  {32'h3f8ca5b0, 32'h3fabfd79} /* (26, 1, 18) {real, imag} */,
  {32'h3f06d585, 32'h3e0debbe} /* (26, 1, 17) {real, imag} */,
  {32'hbdf554ac, 32'hbe92891c} /* (26, 1, 16) {real, imag} */,
  {32'hbebb3906, 32'h40147820} /* (26, 1, 15) {real, imag} */,
  {32'h3e5f49ad, 32'hbe416d2a} /* (26, 1, 14) {real, imag} */,
  {32'h402ea663, 32'hc044d3a3} /* (26, 1, 13) {real, imag} */,
  {32'hbf01a688, 32'h4024e197} /* (26, 1, 12) {real, imag} */,
  {32'hbf85adaa, 32'hbfb20aa0} /* (26, 1, 11) {real, imag} */,
  {32'hc02424cf, 32'hbf75d9de} /* (26, 1, 10) {real, imag} */,
  {32'h40222462, 32'h3dc9cc69} /* (26, 1, 9) {real, imag} */,
  {32'hc02cbc29, 32'h400163d0} /* (26, 1, 8) {real, imag} */,
  {32'h404074f6, 32'hbfb1156b} /* (26, 1, 7) {real, imag} */,
  {32'hbf261d28, 32'h4041b257} /* (26, 1, 6) {real, imag} */,
  {32'hbeb8a664, 32'hbf6f2b14} /* (26, 1, 5) {real, imag} */,
  {32'hbf9058a9, 32'hc0bbe310} /* (26, 1, 4) {real, imag} */,
  {32'h41382502, 32'hbfd3efca} /* (26, 1, 3) {real, imag} */,
  {32'hbf913e86, 32'h4036d137} /* (26, 1, 2) {real, imag} */,
  {32'hc0890c3e, 32'h400c9d5f} /* (26, 1, 1) {real, imag} */,
  {32'hc112c05e, 32'h3ef71cae} /* (26, 1, 0) {real, imag} */,
  {32'h40737003, 32'hbfa344c0} /* (26, 0, 31) {real, imag} */,
  {32'h40bc2028, 32'hc0db7cb5} /* (26, 0, 30) {real, imag} */,
  {32'h3e7dbb0b, 32'hc007a621} /* (26, 0, 29) {real, imag} */,
  {32'hc02b48eb, 32'h4095414c} /* (26, 0, 28) {real, imag} */,
  {32'hbfc27fa9, 32'h406aae23} /* (26, 0, 27) {real, imag} */,
  {32'hbf0c8e4a, 32'hbfd787ce} /* (26, 0, 26) {real, imag} */,
  {32'h40a61a8b, 32'h4019199d} /* (26, 0, 25) {real, imag} */,
  {32'hbf968e29, 32'h3f50adcd} /* (26, 0, 24) {real, imag} */,
  {32'hbf7a539e, 32'h3fadfb1a} /* (26, 0, 23) {real, imag} */,
  {32'hbf990497, 32'h4028456c} /* (26, 0, 22) {real, imag} */,
  {32'h3f2e2b6b, 32'h4052b595} /* (26, 0, 21) {real, imag} */,
  {32'h3ee38372, 32'h3fe61ccd} /* (26, 0, 20) {real, imag} */,
  {32'hc05269f2, 32'h3ff7c591} /* (26, 0, 19) {real, imag} */,
  {32'h3fbb126b, 32'hc02da3b5} /* (26, 0, 18) {real, imag} */,
  {32'hbf111999, 32'h3f271b7e} /* (26, 0, 17) {real, imag} */,
  {32'hbef56a0b, 32'hc00732f1} /* (26, 0, 16) {real, imag} */,
  {32'hbff50780, 32'hbe8f0233} /* (26, 0, 15) {real, imag} */,
  {32'hbfdd25f5, 32'hbe6d4e17} /* (26, 0, 14) {real, imag} */,
  {32'h3f3c2d37, 32'hbfb4a9e9} /* (26, 0, 13) {real, imag} */,
  {32'h3f7d94d2, 32'hbeae23dd} /* (26, 0, 12) {real, imag} */,
  {32'hbf45ebd9, 32'h3f04edc0} /* (26, 0, 11) {real, imag} */,
  {32'h3fedc330, 32'hbfde1e51} /* (26, 0, 10) {real, imag} */,
  {32'hbfe42acf, 32'hbf66f86b} /* (26, 0, 9) {real, imag} */,
  {32'hbf7c3987, 32'h409b274a} /* (26, 0, 8) {real, imag} */,
  {32'h3fae9a81, 32'h3fc39489} /* (26, 0, 7) {real, imag} */,
  {32'h3e4b256f, 32'hbfe8122e} /* (26, 0, 6) {real, imag} */,
  {32'h4092bdb7, 32'hc10bbc7b} /* (26, 0, 5) {real, imag} */,
  {32'hbf97bb6a, 32'h4084127d} /* (26, 0, 4) {real, imag} */,
  {32'h3e1fd7e6, 32'hbd5d435f} /* (26, 0, 3) {real, imag} */,
  {32'hc0dc3da7, 32'h3f64887e} /* (26, 0, 2) {real, imag} */,
  {32'h3f381d16, 32'hc0c43062} /* (26, 0, 1) {real, imag} */,
  {32'h40fce6ce, 32'hc0e29fd0} /* (26, 0, 0) {real, imag} */,
  {32'h409763a3, 32'h407a1664} /* (25, 31, 31) {real, imag} */,
  {32'hc0490f6d, 32'hc0a2cb24} /* (25, 31, 30) {real, imag} */,
  {32'hbdd3430e, 32'h409a65ea} /* (25, 31, 29) {real, imag} */,
  {32'h3d3be098, 32'hbdcfd68d} /* (25, 31, 28) {real, imag} */,
  {32'hbf4d7b3e, 32'h3fa97efa} /* (25, 31, 27) {real, imag} */,
  {32'h40629c76, 32'h40d22625} /* (25, 31, 26) {real, imag} */,
  {32'h3d16874d, 32'hbfdd2beb} /* (25, 31, 25) {real, imag} */,
  {32'hbfa65773, 32'h3e97de3b} /* (25, 31, 24) {real, imag} */,
  {32'h3f008fc9, 32'h3da75a67} /* (25, 31, 23) {real, imag} */,
  {32'hc0556c23, 32'h3f9fa9ee} /* (25, 31, 22) {real, imag} */,
  {32'hbf836365, 32'h40369d50} /* (25, 31, 21) {real, imag} */,
  {32'h3d48f037, 32'hbfa65995} /* (25, 31, 20) {real, imag} */,
  {32'h3fbc0a26, 32'hbf0f296c} /* (25, 31, 19) {real, imag} */,
  {32'h3e16bb1f, 32'h3fd336e0} /* (25, 31, 18) {real, imag} */,
  {32'hbf279ac2, 32'hbf4069d9} /* (25, 31, 17) {real, imag} */,
  {32'h3f197904, 32'h3ee462f4} /* (25, 31, 16) {real, imag} */,
  {32'hbf02c5c8, 32'hbf9767f4} /* (25, 31, 15) {real, imag} */,
  {32'hc00bad2c, 32'hbf809ccf} /* (25, 31, 14) {real, imag} */,
  {32'h3f9db8d9, 32'h400c15a5} /* (25, 31, 13) {real, imag} */,
  {32'hbfc55d66, 32'hbfe21a43} /* (25, 31, 12) {real, imag} */,
  {32'hbff1cbbb, 32'h3fbc7764} /* (25, 31, 11) {real, imag} */,
  {32'hc08dfb6f, 32'hbfb1550d} /* (25, 31, 10) {real, imag} */,
  {32'h3fc57399, 32'h4091676b} /* (25, 31, 9) {real, imag} */,
  {32'h3f461ace, 32'h3fe8a5a4} /* (25, 31, 8) {real, imag} */,
  {32'h3fe24452, 32'hc09dbc5b} /* (25, 31, 7) {real, imag} */,
  {32'h3f886cd6, 32'hbf4faf88} /* (25, 31, 6) {real, imag} */,
  {32'h402b6528, 32'hc0c76abe} /* (25, 31, 5) {real, imag} */,
  {32'h40772e6c, 32'h3fa06ff3} /* (25, 31, 4) {real, imag} */,
  {32'h3ebcef90, 32'hc001a5cc} /* (25, 31, 3) {real, imag} */,
  {32'hc0c51e8f, 32'hc0931558} /* (25, 31, 2) {real, imag} */,
  {32'h3de7cae4, 32'h40f47d5d} /* (25, 31, 1) {real, imag} */,
  {32'h3f6fab2c, 32'hc06c72c2} /* (25, 31, 0) {real, imag} */,
  {32'hbf6b7468, 32'hbfe6bd0a} /* (25, 30, 31) {real, imag} */,
  {32'hc07895b2, 32'h402c0f95} /* (25, 30, 30) {real, imag} */,
  {32'h40778266, 32'h3e9af201} /* (25, 30, 29) {real, imag} */,
  {32'h3fbc3799, 32'h3f84f7a0} /* (25, 30, 28) {real, imag} */,
  {32'h4065cc30, 32'h3fc3022d} /* (25, 30, 27) {real, imag} */,
  {32'hbfd1690d, 32'hbfa3b5fd} /* (25, 30, 26) {real, imag} */,
  {32'h3f86c24e, 32'h3dd29f9b} /* (25, 30, 25) {real, imag} */,
  {32'h3fa0cec5, 32'hbd617b9b} /* (25, 30, 24) {real, imag} */,
  {32'h40708586, 32'hbe861fc6} /* (25, 30, 23) {real, imag} */,
  {32'hc05169ec, 32'h3d5e8957} /* (25, 30, 22) {real, imag} */,
  {32'hc091ad36, 32'h3ff4a0aa} /* (25, 30, 21) {real, imag} */,
  {32'h3fd49c5f, 32'hbf18b534} /* (25, 30, 20) {real, imag} */,
  {32'hbeb4fcfe, 32'hbef2b1a0} /* (25, 30, 19) {real, imag} */,
  {32'h3fbc6c46, 32'hbe93095b} /* (25, 30, 18) {real, imag} */,
  {32'hbd8fa4b4, 32'hbe5176d8} /* (25, 30, 17) {real, imag} */,
  {32'h3ea74fbb, 32'h3f848bc9} /* (25, 30, 16) {real, imag} */,
  {32'h3f3b34b3, 32'hc0413ea5} /* (25, 30, 15) {real, imag} */,
  {32'h3ea490c1, 32'h3fca6d9e} /* (25, 30, 14) {real, imag} */,
  {32'hbeb9d596, 32'hbf7ad8ee} /* (25, 30, 13) {real, imag} */,
  {32'h3fe4f444, 32'hbf3328db} /* (25, 30, 12) {real, imag} */,
  {32'hc03b03ee, 32'h3ef6e33f} /* (25, 30, 11) {real, imag} */,
  {32'hbfcf3ef3, 32'hbf63649c} /* (25, 30, 10) {real, imag} */,
  {32'h3fcd4468, 32'hbf169679} /* (25, 30, 9) {real, imag} */,
  {32'h3fadeef4, 32'h408c29e1} /* (25, 30, 8) {real, imag} */,
  {32'h3ea8ef7a, 32'hc041e13e} /* (25, 30, 7) {real, imag} */,
  {32'hbfa52dea, 32'hbf445802} /* (25, 30, 6) {real, imag} */,
  {32'hc02f02fd, 32'hbff2279f} /* (25, 30, 5) {real, imag} */,
  {32'h4075b2ad, 32'h40a43eca} /* (25, 30, 4) {real, imag} */,
  {32'hc0d9afc8, 32'h40addadc} /* (25, 30, 3) {real, imag} */,
  {32'hbfeedbdc, 32'h40bf490c} /* (25, 30, 2) {real, imag} */,
  {32'hc037f6c1, 32'hc03d50d4} /* (25, 30, 1) {real, imag} */,
  {32'hbf82554f, 32'hc03e8a55} /* (25, 30, 0) {real, imag} */,
  {32'h407002c3, 32'hbf5859f4} /* (25, 29, 31) {real, imag} */,
  {32'h3fc6b4df, 32'h3fd239b9} /* (25, 29, 30) {real, imag} */,
  {32'h40b7ea11, 32'hbe1bad15} /* (25, 29, 29) {real, imag} */,
  {32'h406b4b67, 32'h3e005b62} /* (25, 29, 28) {real, imag} */,
  {32'hc0145cc2, 32'h40813cc0} /* (25, 29, 27) {real, imag} */,
  {32'hc026ac0d, 32'hc020d137} /* (25, 29, 26) {real, imag} */,
  {32'hc0837067, 32'hbf11118c} /* (25, 29, 25) {real, imag} */,
  {32'h3ea498c6, 32'hbf879e63} /* (25, 29, 24) {real, imag} */,
  {32'h3ea813ed, 32'h405b232f} /* (25, 29, 23) {real, imag} */,
  {32'h3efb8eca, 32'h3fccc4de} /* (25, 29, 22) {real, imag} */,
  {32'h4018e8e9, 32'h3e904283} /* (25, 29, 21) {real, imag} */,
  {32'h3f7e4ee4, 32'h4027b10c} /* (25, 29, 20) {real, imag} */,
  {32'hbe249acf, 32'hbe93e64a} /* (25, 29, 19) {real, imag} */,
  {32'hc0897ba4, 32'h3fb37b14} /* (25, 29, 18) {real, imag} */,
  {32'h3f829fdf, 32'h3eaffe45} /* (25, 29, 17) {real, imag} */,
  {32'hbf285bad, 32'h3ee73729} /* (25, 29, 16) {real, imag} */,
  {32'hbf1a62a5, 32'h3f50d116} /* (25, 29, 15) {real, imag} */,
  {32'h3f6d3472, 32'h3f20433a} /* (25, 29, 14) {real, imag} */,
  {32'hbf273200, 32'hc04ed7f6} /* (25, 29, 13) {real, imag} */,
  {32'h404a8983, 32'h409cb89d} /* (25, 29, 12) {real, imag} */,
  {32'hbe82ad2b, 32'h3f82c020} /* (25, 29, 11) {real, imag} */,
  {32'hbf2bc28c, 32'hbfcfcb4e} /* (25, 29, 10) {real, imag} */,
  {32'h3fa3b94b, 32'hc0646ebd} /* (25, 29, 9) {real, imag} */,
  {32'h3fdd2b4b, 32'h3e99839d} /* (25, 29, 8) {real, imag} */,
  {32'h3fb89379, 32'h3f4ed297} /* (25, 29, 7) {real, imag} */,
  {32'h3fa99b2b, 32'h401b90fd} /* (25, 29, 6) {real, imag} */,
  {32'h3de8c478, 32'h3fec5eb9} /* (25, 29, 5) {real, imag} */,
  {32'hbef4b4e7, 32'h4024fce1} /* (25, 29, 4) {real, imag} */,
  {32'hbe020d8f, 32'hc0c90093} /* (25, 29, 3) {real, imag} */,
  {32'h3e56f5aa, 32'hc03f10aa} /* (25, 29, 2) {real, imag} */,
  {32'hc0c361d7, 32'h4097e66b} /* (25, 29, 1) {real, imag} */,
  {32'h40821060, 32'hbeeff27e} /* (25, 29, 0) {real, imag} */,
  {32'hbedc56f7, 32'hc01d25d2} /* (25, 28, 31) {real, imag} */,
  {32'h3fd81941, 32'h40e6085e} /* (25, 28, 30) {real, imag} */,
  {32'hc03ca09e, 32'hc04abd27} /* (25, 28, 29) {real, imag} */,
  {32'h40a9cd28, 32'h3b8eb776} /* (25, 28, 28) {real, imag} */,
  {32'h3f9b398a, 32'hbfa7aa30} /* (25, 28, 27) {real, imag} */,
  {32'h3f326465, 32'hc00cac98} /* (25, 28, 26) {real, imag} */,
  {32'hc0443ea8, 32'h3fad079a} /* (25, 28, 25) {real, imag} */,
  {32'h402b051e, 32'hc025c588} /* (25, 28, 24) {real, imag} */,
  {32'hbfdc52f5, 32'h4007ce17} /* (25, 28, 23) {real, imag} */,
  {32'h3eaa5e78, 32'h3f99d914} /* (25, 28, 22) {real, imag} */,
  {32'h3f95f93d, 32'hc0292bf4} /* (25, 28, 21) {real, imag} */,
  {32'h3fb39e82, 32'h3fec99e6} /* (25, 28, 20) {real, imag} */,
  {32'hc0803d18, 32'h3f7b7788} /* (25, 28, 19) {real, imag} */,
  {32'h3ef51379, 32'hc0121b86} /* (25, 28, 18) {real, imag} */,
  {32'h3eac0742, 32'h3df922db} /* (25, 28, 17) {real, imag} */,
  {32'h3ec07c23, 32'hbed6a5a2} /* (25, 28, 16) {real, imag} */,
  {32'hbe80cda6, 32'h3f8cabe5} /* (25, 28, 15) {real, imag} */,
  {32'hbf6efca5, 32'hc05997db} /* (25, 28, 14) {real, imag} */,
  {32'hbfa59aa2, 32'h3e2ac4c3} /* (25, 28, 13) {real, imag} */,
  {32'h3ef2b476, 32'hbe5baa05} /* (25, 28, 12) {real, imag} */,
  {32'hc06bd578, 32'h4002a3e3} /* (25, 28, 11) {real, imag} */,
  {32'hbf6d823d, 32'hc0694904} /* (25, 28, 10) {real, imag} */,
  {32'hbd7704c9, 32'hbc8c7efa} /* (25, 28, 9) {real, imag} */,
  {32'h40343ddd, 32'hc005b946} /* (25, 28, 8) {real, imag} */,
  {32'h3f6645d6, 32'hbff24a22} /* (25, 28, 7) {real, imag} */,
  {32'hbfcac594, 32'hc00457c7} /* (25, 28, 6) {real, imag} */,
  {32'h4071cd51, 32'h4041aad2} /* (25, 28, 5) {real, imag} */,
  {32'hc0162930, 32'hc05439b7} /* (25, 28, 4) {real, imag} */,
  {32'hbf6db6e9, 32'h40249f7e} /* (25, 28, 3) {real, imag} */,
  {32'h405dc3af, 32'h4091c81a} /* (25, 28, 2) {real, imag} */,
  {32'h3fdd7fbc, 32'h3ff9aba1} /* (25, 28, 1) {real, imag} */,
  {32'hbf1a5b02, 32'hc01fa95b} /* (25, 28, 0) {real, imag} */,
  {32'hbffb6a83, 32'h3f610af9} /* (25, 27, 31) {real, imag} */,
  {32'hc044a891, 32'hc04357c8} /* (25, 27, 30) {real, imag} */,
  {32'hbf84621c, 32'h403ea424} /* (25, 27, 29) {real, imag} */,
  {32'h3fb4996e, 32'hbff4ce17} /* (25, 27, 28) {real, imag} */,
  {32'hbf6426a4, 32'hbf9b8c82} /* (25, 27, 27) {real, imag} */,
  {32'hc019f548, 32'hbf1ed62b} /* (25, 27, 26) {real, imag} */,
  {32'h40227cc1, 32'h4040f060} /* (25, 27, 25) {real, imag} */,
  {32'h3f3ff1af, 32'hbfd83755} /* (25, 27, 24) {real, imag} */,
  {32'h3de9794a, 32'hc05276c1} /* (25, 27, 23) {real, imag} */,
  {32'hbf09a76b, 32'hc0a89c3b} /* (25, 27, 22) {real, imag} */,
  {32'hbd59ceb8, 32'h4025d394} /* (25, 27, 21) {real, imag} */,
  {32'h3f07ac39, 32'h3fc6ad2c} /* (25, 27, 20) {real, imag} */,
  {32'h3f8fd92f, 32'h3f8e8160} /* (25, 27, 19) {real, imag} */,
  {32'h3f924607, 32'hbec87350} /* (25, 27, 18) {real, imag} */,
  {32'h3fbb3296, 32'h3f5c0b5b} /* (25, 27, 17) {real, imag} */,
  {32'h3fae5f0b, 32'hbe2f4c76} /* (25, 27, 16) {real, imag} */,
  {32'h3e56715e, 32'hbf75a46c} /* (25, 27, 15) {real, imag} */,
  {32'h4073a847, 32'hbfb5c189} /* (25, 27, 14) {real, imag} */,
  {32'hc08aca65, 32'hbf242182} /* (25, 27, 13) {real, imag} */,
  {32'hbff78a89, 32'h3f298e58} /* (25, 27, 12) {real, imag} */,
  {32'hbffeec3a, 32'h3f7045b9} /* (25, 27, 11) {real, imag} */,
  {32'h3f2b8109, 32'hbeb64880} /* (25, 27, 10) {real, imag} */,
  {32'h404f4cc7, 32'hc0475a97} /* (25, 27, 9) {real, imag} */,
  {32'hbe52d29a, 32'h3fa995b2} /* (25, 27, 8) {real, imag} */,
  {32'h4019b29f, 32'hc099d42b} /* (25, 27, 7) {real, imag} */,
  {32'hc062a917, 32'hbf25012f} /* (25, 27, 6) {real, imag} */,
  {32'h409a441f, 32'h4036ef07} /* (25, 27, 5) {real, imag} */,
  {32'h3f6f6dcb, 32'h3fe73126} /* (25, 27, 4) {real, imag} */,
  {32'h3fa5982e, 32'hbee52088} /* (25, 27, 3) {real, imag} */,
  {32'hbe5254aa, 32'hc0e05c31} /* (25, 27, 2) {real, imag} */,
  {32'h3fc45461, 32'hbfad402b} /* (25, 27, 1) {real, imag} */,
  {32'h3f9f48c0, 32'h40cc51fe} /* (25, 27, 0) {real, imag} */,
  {32'h4084c039, 32'hbff2eb66} /* (25, 26, 31) {real, imag} */,
  {32'hbfaad2ba, 32'h4048da45} /* (25, 26, 30) {real, imag} */,
  {32'hbe87c8cb, 32'h3ee06e91} /* (25, 26, 29) {real, imag} */,
  {32'h3fd3a594, 32'hbebbef6b} /* (25, 26, 28) {real, imag} */,
  {32'hbfe2724e, 32'h3fa8b143} /* (25, 26, 27) {real, imag} */,
  {32'hbec408c3, 32'h3ec9fa3b} /* (25, 26, 26) {real, imag} */,
  {32'hbf1e9f13, 32'h4009e43e} /* (25, 26, 25) {real, imag} */,
  {32'hc017f1e5, 32'hc006826b} /* (25, 26, 24) {real, imag} */,
  {32'h3fa3cbcf, 32'h401deea7} /* (25, 26, 23) {real, imag} */,
  {32'h3f46d172, 32'h3f0f966d} /* (25, 26, 22) {real, imag} */,
  {32'hbc3bb38b, 32'hc03c6002} /* (25, 26, 21) {real, imag} */,
  {32'h3c4bb7a4, 32'h3f90ca8e} /* (25, 26, 20) {real, imag} */,
  {32'h3e826534, 32'hc0521c35} /* (25, 26, 19) {real, imag} */,
  {32'h3f59e21a, 32'h3ed42ee7} /* (25, 26, 18) {real, imag} */,
  {32'h3ee3b1dc, 32'hbeee8b53} /* (25, 26, 17) {real, imag} */,
  {32'h3e9bfd4a, 32'h3f0b6536} /* (25, 26, 16) {real, imag} */,
  {32'hbe5f9f43, 32'hbfc18d28} /* (25, 26, 15) {real, imag} */,
  {32'hbe96ecb4, 32'h3ef3f5b9} /* (25, 26, 14) {real, imag} */,
  {32'hbf8a010d, 32'h40082647} /* (25, 26, 13) {real, imag} */,
  {32'h3e526a36, 32'h3fb9fbc2} /* (25, 26, 12) {real, imag} */,
  {32'h4020a027, 32'hc03aea57} /* (25, 26, 11) {real, imag} */,
  {32'hc0599002, 32'hbfb4da83} /* (25, 26, 10) {real, imag} */,
  {32'h400ae0bd, 32'hbc996bfa} /* (25, 26, 9) {real, imag} */,
  {32'hbfad50d5, 32'hbf679588} /* (25, 26, 8) {real, imag} */,
  {32'h4039cbac, 32'h3f39b60f} /* (25, 26, 7) {real, imag} */,
  {32'hbfd35fe4, 32'hbcebeab9} /* (25, 26, 6) {real, imag} */,
  {32'hc011e565, 32'hc02e2e34} /* (25, 26, 5) {real, imag} */,
  {32'h3ed43ec5, 32'hbfcc866d} /* (25, 26, 4) {real, imag} */,
  {32'h3f128cc0, 32'hc04cefe0} /* (25, 26, 3) {real, imag} */,
  {32'h408897d5, 32'hbf079b69} /* (25, 26, 2) {real, imag} */,
  {32'hbfee4a2b, 32'h3ff72a9a} /* (25, 26, 1) {real, imag} */,
  {32'hbe9d8e07, 32'h3f51abcf} /* (25, 26, 0) {real, imag} */,
  {32'h40161171, 32'h3f8c6339} /* (25, 25, 31) {real, imag} */,
  {32'h3fa5c054, 32'hbfb9ba53} /* (25, 25, 30) {real, imag} */,
  {32'hc045c3d9, 32'hbf19e8b0} /* (25, 25, 29) {real, imag} */,
  {32'hbf8338f1, 32'h3f7a1b2a} /* (25, 25, 28) {real, imag} */,
  {32'h3ed9be5d, 32'hc04ddeec} /* (25, 25, 27) {real, imag} */,
  {32'h3e1e7efa, 32'hc00ace6b} /* (25, 25, 26) {real, imag} */,
  {32'h4002f005, 32'hbdb33e6c} /* (25, 25, 25) {real, imag} */,
  {32'h3f339e92, 32'h3fca0900} /* (25, 25, 24) {real, imag} */,
  {32'hbfea40ab, 32'h4038d59a} /* (25, 25, 23) {real, imag} */,
  {32'hbe5e53c8, 32'h3e84f3a0} /* (25, 25, 22) {real, imag} */,
  {32'hbd86ed63, 32'hbf663317} /* (25, 25, 21) {real, imag} */,
  {32'hbfa3057b, 32'hbee219a4} /* (25, 25, 20) {real, imag} */,
  {32'h3fe81977, 32'h3f7a188c} /* (25, 25, 19) {real, imag} */,
  {32'hbdbe2227, 32'h3f70ecb3} /* (25, 25, 18) {real, imag} */,
  {32'h3f9d25cd, 32'hbfad5feb} /* (25, 25, 17) {real, imag} */,
  {32'h3f3c6ba4, 32'hbc524cc6} /* (25, 25, 16) {real, imag} */,
  {32'h3f8c6f5a, 32'h3f272456} /* (25, 25, 15) {real, imag} */,
  {32'hbea046fb, 32'hc011ac94} /* (25, 25, 14) {real, imag} */,
  {32'hbf4a67cc, 32'h3efc7ebb} /* (25, 25, 13) {real, imag} */,
  {32'h4029d02a, 32'h3f7e8993} /* (25, 25, 12) {real, imag} */,
  {32'h3ffb70a2, 32'hc03fbff3} /* (25, 25, 11) {real, imag} */,
  {32'h4013f104, 32'h3fea99f2} /* (25, 25, 10) {real, imag} */,
  {32'h3ee65d6b, 32'hbfb83b8d} /* (25, 25, 9) {real, imag} */,
  {32'hbee59afd, 32'h3ed50136} /* (25, 25, 8) {real, imag} */,
  {32'h3e625e9b, 32'h4027a426} /* (25, 25, 7) {real, imag} */,
  {32'hc01489d0, 32'h3d51e11c} /* (25, 25, 6) {real, imag} */,
  {32'hbf86a372, 32'hbf1d2347} /* (25, 25, 5) {real, imag} */,
  {32'h3f2478a7, 32'hbf43b812} /* (25, 25, 4) {real, imag} */,
  {32'h402d93f1, 32'hc0431e13} /* (25, 25, 3) {real, imag} */,
  {32'h3fe4795c, 32'hc048b65d} /* (25, 25, 2) {real, imag} */,
  {32'h3f3b8faf, 32'h3f2438ef} /* (25, 25, 1) {real, imag} */,
  {32'hc00aba2c, 32'h3f95e35c} /* (25, 25, 0) {real, imag} */,
  {32'hc00f4bed, 32'h40338d18} /* (25, 24, 31) {real, imag} */,
  {32'hbf5a0c36, 32'h40107047} /* (25, 24, 30) {real, imag} */,
  {32'hbc8d55f1, 32'hbe373fd8} /* (25, 24, 29) {real, imag} */,
  {32'h4021c0b3, 32'hbfc21381} /* (25, 24, 28) {real, imag} */,
  {32'hbfd8eb8a, 32'hbf8baa9e} /* (25, 24, 27) {real, imag} */,
  {32'h3fb4ac91, 32'hbf3021ca} /* (25, 24, 26) {real, imag} */,
  {32'h407b37da, 32'hbf1dfd67} /* (25, 24, 25) {real, imag} */,
  {32'h3f1bfa81, 32'h3e716631} /* (25, 24, 24) {real, imag} */,
  {32'h405d6e0d, 32'hc0412bee} /* (25, 24, 23) {real, imag} */,
  {32'h3fc524e9, 32'h400db481} /* (25, 24, 22) {real, imag} */,
  {32'h40aed304, 32'hbf0589a7} /* (25, 24, 21) {real, imag} */,
  {32'hc06a6491, 32'hbe3a5ccf} /* (25, 24, 20) {real, imag} */,
  {32'hbe8fa90e, 32'h3f83435b} /* (25, 24, 19) {real, imag} */,
  {32'hbf0cb0ac, 32'hbfaaf334} /* (25, 24, 18) {real, imag} */,
  {32'hbf1808e9, 32'h40272339} /* (25, 24, 17) {real, imag} */,
  {32'hbdde132e, 32'h3fb14b83} /* (25, 24, 16) {real, imag} */,
  {32'hc02332ab, 32'hbed9cb7c} /* (25, 24, 15) {real, imag} */,
  {32'hbee35ee8, 32'h3f6daf19} /* (25, 24, 14) {real, imag} */,
  {32'h3fe7905f, 32'hbf066abb} /* (25, 24, 13) {real, imag} */,
  {32'h3efe382a, 32'h3f4cfe3d} /* (25, 24, 12) {real, imag} */,
  {32'hbf70c0dd, 32'hbe6dd0b4} /* (25, 24, 11) {real, imag} */,
  {32'hbfd30276, 32'h40265717} /* (25, 24, 10) {real, imag} */,
  {32'hc0826949, 32'h3f6a2e1e} /* (25, 24, 9) {real, imag} */,
  {32'hbfbb301d, 32'hbf4091b3} /* (25, 24, 8) {real, imag} */,
  {32'hc00fa17b, 32'h3ee9d406} /* (25, 24, 7) {real, imag} */,
  {32'h3f0ec09e, 32'h407d27c5} /* (25, 24, 6) {real, imag} */,
  {32'h3fd4c5f4, 32'hc0363099} /* (25, 24, 5) {real, imag} */,
  {32'hbf0e7b15, 32'hc0549edb} /* (25, 24, 4) {real, imag} */,
  {32'h4073d52c, 32'h3e950630} /* (25, 24, 3) {real, imag} */,
  {32'hbfaea303, 32'hbf54c91b} /* (25, 24, 2) {real, imag} */,
  {32'hbe843ca6, 32'hbf9430c8} /* (25, 24, 1) {real, imag} */,
  {32'h3f46e8bb, 32'hc07cfcb6} /* (25, 24, 0) {real, imag} */,
  {32'h3fb97970, 32'hbfad2e6c} /* (25, 23, 31) {real, imag} */,
  {32'h40b38d30, 32'hbeb84ee4} /* (25, 23, 30) {real, imag} */,
  {32'h3d70c82f, 32'hbf1af408} /* (25, 23, 29) {real, imag} */,
  {32'hbf8275d8, 32'hbf978c97} /* (25, 23, 28) {real, imag} */,
  {32'hbe131520, 32'h3ea153bc} /* (25, 23, 27) {real, imag} */,
  {32'hbfab900a, 32'h40666382} /* (25, 23, 26) {real, imag} */,
  {32'hc00fbd00, 32'hc0a88b3f} /* (25, 23, 25) {real, imag} */,
  {32'h3ff2d3d5, 32'hbfa065b0} /* (25, 23, 24) {real, imag} */,
  {32'hbf000d26, 32'h40797eb3} /* (25, 23, 23) {real, imag} */,
  {32'h40389a42, 32'hc067df92} /* (25, 23, 22) {real, imag} */,
  {32'hc0112c65, 32'h3f84dfe0} /* (25, 23, 21) {real, imag} */,
  {32'h3f9d821b, 32'hbee2f59f} /* (25, 23, 20) {real, imag} */,
  {32'h40125509, 32'h3f0745dc} /* (25, 23, 19) {real, imag} */,
  {32'h3f0b2845, 32'hbfa55e71} /* (25, 23, 18) {real, imag} */,
  {32'h3eea8939, 32'h3f8aefb8} /* (25, 23, 17) {real, imag} */,
  {32'h3ee8a782, 32'h3f9d10de} /* (25, 23, 16) {real, imag} */,
  {32'hbf79342f, 32'hbffa0c8f} /* (25, 23, 15) {real, imag} */,
  {32'h3f6b6e98, 32'h40008ace} /* (25, 23, 14) {real, imag} */,
  {32'h3fe9b021, 32'h3fe6bb79} /* (25, 23, 13) {real, imag} */,
  {32'hbf95889e, 32'hbecd7cef} /* (25, 23, 12) {real, imag} */,
  {32'hc050ea16, 32'hbf943498} /* (25, 23, 11) {real, imag} */,
  {32'h404a3bc5, 32'hc01a2dee} /* (25, 23, 10) {real, imag} */,
  {32'h3f96a4e1, 32'h3f0218e5} /* (25, 23, 9) {real, imag} */,
  {32'hbbb6b89a, 32'h3fee16b4} /* (25, 23, 8) {real, imag} */,
  {32'h4073acb9, 32'hbf40eaeb} /* (25, 23, 7) {real, imag} */,
  {32'hbfcd55b6, 32'hbeb63c82} /* (25, 23, 6) {real, imag} */,
  {32'hbf6d5ef7, 32'h3ffe01bd} /* (25, 23, 5) {real, imag} */,
  {32'h400e4a37, 32'h3e87f8ae} /* (25, 23, 4) {real, imag} */,
  {32'hbf42742c, 32'hbf9cf707} /* (25, 23, 3) {real, imag} */,
  {32'h3fb9d499, 32'hbeef80d6} /* (25, 23, 2) {real, imag} */,
  {32'h3f62a0be, 32'h3fd201fb} /* (25, 23, 1) {real, imag} */,
  {32'hbf826782, 32'hc0363344} /* (25, 23, 0) {real, imag} */,
  {32'h3f0895d2, 32'h3f9073a0} /* (25, 22, 31) {real, imag} */,
  {32'h40161005, 32'hc0298ee6} /* (25, 22, 30) {real, imag} */,
  {32'hbeafeff3, 32'h4048c269} /* (25, 22, 29) {real, imag} */,
  {32'hbffdf99e, 32'h3eed29a6} /* (25, 22, 28) {real, imag} */,
  {32'hbfb7276d, 32'hbfb7faf5} /* (25, 22, 27) {real, imag} */,
  {32'hbf9b6b54, 32'hbfeb90cb} /* (25, 22, 26) {real, imag} */,
  {32'h3faaeb37, 32'hbc8417fd} /* (25, 22, 25) {real, imag} */,
  {32'hbf3b0651, 32'hbfac6cde} /* (25, 22, 24) {real, imag} */,
  {32'hbe059e56, 32'h3f84e753} /* (25, 22, 23) {real, imag} */,
  {32'h3ef8e661, 32'h401fcd66} /* (25, 22, 22) {real, imag} */,
  {32'hbf0dd4fe, 32'hbe6e0e23} /* (25, 22, 21) {real, imag} */,
  {32'h403fc72d, 32'h3fad088f} /* (25, 22, 20) {real, imag} */,
  {32'hbea2357e, 32'hbfe469c2} /* (25, 22, 19) {real, imag} */,
  {32'hbec99b03, 32'h3fae5fc3} /* (25, 22, 18) {real, imag} */,
  {32'hbf9399d3, 32'hbf0e3783} /* (25, 22, 17) {real, imag} */,
  {32'hbe38ae3b, 32'h3e885104} /* (25, 22, 16) {real, imag} */,
  {32'hbd76a4aa, 32'h40230003} /* (25, 22, 15) {real, imag} */,
  {32'h3f01de98, 32'h3ebe48e9} /* (25, 22, 14) {real, imag} */,
  {32'hc0881e30, 32'hbf720a2c} /* (25, 22, 13) {real, imag} */,
  {32'hc0372de5, 32'hbf379900} /* (25, 22, 12) {real, imag} */,
  {32'hc03d7d5d, 32'hbffbb7aa} /* (25, 22, 11) {real, imag} */,
  {32'h4051141d, 32'h3fbab7e9} /* (25, 22, 10) {real, imag} */,
  {32'hbf4870b5, 32'h404b4cdb} /* (25, 22, 9) {real, imag} */,
  {32'h3fbfd717, 32'hc00fc79e} /* (25, 22, 8) {real, imag} */,
  {32'h3ff991d7, 32'h4035c019} /* (25, 22, 7) {real, imag} */,
  {32'h3f4f84ef, 32'hc0650fad} /* (25, 22, 6) {real, imag} */,
  {32'h3f2d56ff, 32'hbffee69e} /* (25, 22, 5) {real, imag} */,
  {32'hc049b161, 32'h3f3e1e78} /* (25, 22, 4) {real, imag} */,
  {32'hbfb1955a, 32'hc032c38a} /* (25, 22, 3) {real, imag} */,
  {32'hbfc3c00c, 32'h40438ccd} /* (25, 22, 2) {real, imag} */,
  {32'h3e643d74, 32'h3fb32e90} /* (25, 22, 1) {real, imag} */,
  {32'h3fbcf87a, 32'hbe90c6aa} /* (25, 22, 0) {real, imag} */,
  {32'hc06e8f33, 32'h401bb747} /* (25, 21, 31) {real, imag} */,
  {32'h404771ad, 32'h3fc87e5f} /* (25, 21, 30) {real, imag} */,
  {32'hbf8904f9, 32'hbfd10444} /* (25, 21, 29) {real, imag} */,
  {32'hbf96f087, 32'h3f1d441d} /* (25, 21, 28) {real, imag} */,
  {32'hbede4b0e, 32'h3f854960} /* (25, 21, 27) {real, imag} */,
  {32'hc0153e0d, 32'hc00e1857} /* (25, 21, 26) {real, imag} */,
  {32'h40804333, 32'hbf0aab69} /* (25, 21, 25) {real, imag} */,
  {32'h3f51b686, 32'h3ca25ebd} /* (25, 21, 24) {real, imag} */,
  {32'hc03560cc, 32'hbf95eda9} /* (25, 21, 23) {real, imag} */,
  {32'hc04e9b08, 32'h3f71ddfe} /* (25, 21, 22) {real, imag} */,
  {32'hbfeddba4, 32'h3f40d054} /* (25, 21, 21) {real, imag} */,
  {32'h3e72b425, 32'h3fbea9ff} /* (25, 21, 20) {real, imag} */,
  {32'h3fda1f6f, 32'h4092c1df} /* (25, 21, 19) {real, imag} */,
  {32'h4047c21d, 32'h3e1bacd1} /* (25, 21, 18) {real, imag} */,
  {32'hbf3ff85e, 32'hc01b032e} /* (25, 21, 17) {real, imag} */,
  {32'h3fe9da91, 32'h3fa9ce0d} /* (25, 21, 16) {real, imag} */,
  {32'hbdaf0f96, 32'h3e75faa1} /* (25, 21, 15) {real, imag} */,
  {32'hbf7810be, 32'h3fc574c9} /* (25, 21, 14) {real, imag} */,
  {32'hbfa964f7, 32'hc006b899} /* (25, 21, 13) {real, imag} */,
  {32'h3f090b59, 32'hc01a8b3c} /* (25, 21, 12) {real, imag} */,
  {32'h3f305e3b, 32'h3e71342c} /* (25, 21, 11) {real, imag} */,
  {32'h3f96caef, 32'h3ef26764} /* (25, 21, 10) {real, imag} */,
  {32'hbf90687e, 32'h4092aea5} /* (25, 21, 9) {real, imag} */,
  {32'hbedfb4bb, 32'h402db096} /* (25, 21, 8) {real, imag} */,
  {32'h3febd5a2, 32'h400c500f} /* (25, 21, 7) {real, imag} */,
  {32'hbe056a2a, 32'h3f993dd2} /* (25, 21, 6) {real, imag} */,
  {32'h405fa76b, 32'hc06b4251} /* (25, 21, 5) {real, imag} */,
  {32'hbe642d64, 32'hbf1aaecf} /* (25, 21, 4) {real, imag} */,
  {32'hc0263923, 32'hbfd3ba86} /* (25, 21, 3) {real, imag} */,
  {32'hbffc01d9, 32'h4022df3e} /* (25, 21, 2) {real, imag} */,
  {32'hbfd780e9, 32'hbe6199e8} /* (25, 21, 1) {real, imag} */,
  {32'hbf639671, 32'h3f961d0c} /* (25, 21, 0) {real, imag} */,
  {32'hbf104d9a, 32'hbfc46b2b} /* (25, 20, 31) {real, imag} */,
  {32'hbf5dcef1, 32'h3f1dbf4c} /* (25, 20, 30) {real, imag} */,
  {32'h3e81c4bd, 32'hbe86d6b1} /* (25, 20, 29) {real, imag} */,
  {32'hbf33493c, 32'h3ee0e89f} /* (25, 20, 28) {real, imag} */,
  {32'h403e47e8, 32'hbfea3efe} /* (25, 20, 27) {real, imag} */,
  {32'h3e45d243, 32'h3f0ccd11} /* (25, 20, 26) {real, imag} */,
  {32'hc00d64db, 32'h3f8df64f} /* (25, 20, 25) {real, imag} */,
  {32'h3eb7b0a3, 32'h4088fcb4} /* (25, 20, 24) {real, imag} */,
  {32'h40703106, 32'hc014e6b3} /* (25, 20, 23) {real, imag} */,
  {32'hbfe489be, 32'hbf8b01a2} /* (25, 20, 22) {real, imag} */,
  {32'hbda7b70e, 32'hbf778469} /* (25, 20, 21) {real, imag} */,
  {32'hbf40b06d, 32'hbfeb6d64} /* (25, 20, 20) {real, imag} */,
  {32'h3f74a211, 32'h3f934a72} /* (25, 20, 19) {real, imag} */,
  {32'hbff9f654, 32'h3fbb2b5f} /* (25, 20, 18) {real, imag} */,
  {32'h3efbb759, 32'h3fcb7b51} /* (25, 20, 17) {real, imag} */,
  {32'hbf303f5b, 32'h3f662205} /* (25, 20, 16) {real, imag} */,
  {32'hbfd942d3, 32'h40250f22} /* (25, 20, 15) {real, imag} */,
  {32'h3f77bcda, 32'h400bb020} /* (25, 20, 14) {real, imag} */,
  {32'h405feaac, 32'h3fe82c2f} /* (25, 20, 13) {real, imag} */,
  {32'h3eb5d95b, 32'h3f5789ce} /* (25, 20, 12) {real, imag} */,
  {32'h4036aa15, 32'hc0a4b64c} /* (25, 20, 11) {real, imag} */,
  {32'h3f88ee07, 32'hbf352065} /* (25, 20, 10) {real, imag} */,
  {32'h400f87c2, 32'hbd4a2d87} /* (25, 20, 9) {real, imag} */,
  {32'hbff75c93, 32'hbfd3f5b7} /* (25, 20, 8) {real, imag} */,
  {32'hbf865ab2, 32'h3fc95300} /* (25, 20, 7) {real, imag} */,
  {32'hbe3362e9, 32'h4096585f} /* (25, 20, 6) {real, imag} */,
  {32'hbf9fe78d, 32'hbf9f9927} /* (25, 20, 5) {real, imag} */,
  {32'hbd925de7, 32'h405a310b} /* (25, 20, 4) {real, imag} */,
  {32'hbf1aa9d7, 32'hc0195999} /* (25, 20, 3) {real, imag} */,
  {32'hbf0d2110, 32'h3f89cae3} /* (25, 20, 2) {real, imag} */,
  {32'h3e3779bd, 32'h3fdf4905} /* (25, 20, 1) {real, imag} */,
  {32'hbe62ab3b, 32'h3f517cde} /* (25, 20, 0) {real, imag} */,
  {32'h403430c5, 32'h3f19b11e} /* (25, 19, 31) {real, imag} */,
  {32'h3f8e9bed, 32'hbf091130} /* (25, 19, 30) {real, imag} */,
  {32'h3d1733f4, 32'h3ea2bcbe} /* (25, 19, 29) {real, imag} */,
  {32'hbef111bc, 32'hbfa630fa} /* (25, 19, 28) {real, imag} */,
  {32'h3f96fbb2, 32'h3d7d0153} /* (25, 19, 27) {real, imag} */,
  {32'hbf81af2e, 32'h409b8d57} /* (25, 19, 26) {real, imag} */,
  {32'hc009039b, 32'hbfc1b0ba} /* (25, 19, 25) {real, imag} */,
  {32'hbf4f9ff1, 32'h3dd300d6} /* (25, 19, 24) {real, imag} */,
  {32'h3f06957c, 32'hc02c416f} /* (25, 19, 23) {real, imag} */,
  {32'h3f9e8f4d, 32'hbfa57906} /* (25, 19, 22) {real, imag} */,
  {32'h40171035, 32'hbf10280a} /* (25, 19, 21) {real, imag} */,
  {32'h3f4e893f, 32'hbf7a9da4} /* (25, 19, 20) {real, imag} */,
  {32'h3fc91cc4, 32'h3ffbd3ac} /* (25, 19, 19) {real, imag} */,
  {32'hbfea4233, 32'h4048145b} /* (25, 19, 18) {real, imag} */,
  {32'h3de9fa41, 32'hc06c9397} /* (25, 19, 17) {real, imag} */,
  {32'h402fc34c, 32'hbf176334} /* (25, 19, 16) {real, imag} */,
  {32'hbf5ba566, 32'hbdf619a6} /* (25, 19, 15) {real, imag} */,
  {32'hbe9f4233, 32'hc0584bee} /* (25, 19, 14) {real, imag} */,
  {32'hbe5302fb, 32'h3ff0f51c} /* (25, 19, 13) {real, imag} */,
  {32'hbf98f727, 32'hc054ac24} /* (25, 19, 12) {real, imag} */,
  {32'h3e9ac23b, 32'h4025ae06} /* (25, 19, 11) {real, imag} */,
  {32'h3f27bb7e, 32'hbfd127f5} /* (25, 19, 10) {real, imag} */,
  {32'h3d183abb, 32'hbf831c5f} /* (25, 19, 9) {real, imag} */,
  {32'h402af66a, 32'h3dc856f9} /* (25, 19, 8) {real, imag} */,
  {32'hbf0c2a30, 32'hbe61a092} /* (25, 19, 7) {real, imag} */,
  {32'hbfbbb70e, 32'h3f83fdbc} /* (25, 19, 6) {real, imag} */,
  {32'h4018056d, 32'hbee5da2c} /* (25, 19, 5) {real, imag} */,
  {32'hbfea11f1, 32'h3f8b20d2} /* (25, 19, 4) {real, imag} */,
  {32'hc029f1be, 32'h40166653} /* (25, 19, 3) {real, imag} */,
  {32'h3f888216, 32'hbf3f463c} /* (25, 19, 2) {real, imag} */,
  {32'hbe3a8b13, 32'hbed217f5} /* (25, 19, 1) {real, imag} */,
  {32'hbfd2c82e, 32'h4013469e} /* (25, 19, 0) {real, imag} */,
  {32'hc01a0610, 32'hbf63e6c0} /* (25, 18, 31) {real, imag} */,
  {32'hbf224c3f, 32'hbfe80e65} /* (25, 18, 30) {real, imag} */,
  {32'h3f6db535, 32'hbe3849b4} /* (25, 18, 29) {real, imag} */,
  {32'hbe8d9d81, 32'hbf6768d9} /* (25, 18, 28) {real, imag} */,
  {32'h3e4ec77c, 32'hbea98952} /* (25, 18, 27) {real, imag} */,
  {32'h4059f775, 32'h3fb8a1a4} /* (25, 18, 26) {real, imag} */,
  {32'h4033d0e1, 32'h3f28f05e} /* (25, 18, 25) {real, imag} */,
  {32'hbf9cc512, 32'h3ecf681d} /* (25, 18, 24) {real, imag} */,
  {32'hbf257f75, 32'h3fa4c3cb} /* (25, 18, 23) {real, imag} */,
  {32'h3fba3072, 32'h3fc5c3c0} /* (25, 18, 22) {real, imag} */,
  {32'h3f2d7ac7, 32'h3f441b1b} /* (25, 18, 21) {real, imag} */,
  {32'h400f3d49, 32'hbf699d75} /* (25, 18, 20) {real, imag} */,
  {32'hbfaafe91, 32'hbf9ade1a} /* (25, 18, 19) {real, imag} */,
  {32'hbf118ee8, 32'hbf620893} /* (25, 18, 18) {real, imag} */,
  {32'hbe5d5e3f, 32'h3faf99b5} /* (25, 18, 17) {real, imag} */,
  {32'h3f2650a9, 32'hbe9c9530} /* (25, 18, 16) {real, imag} */,
  {32'h4003bcb6, 32'h3d02ae1d} /* (25, 18, 15) {real, imag} */,
  {32'h3ff43218, 32'hbf46f779} /* (25, 18, 14) {real, imag} */,
  {32'h3f31a221, 32'h3effa280} /* (25, 18, 13) {real, imag} */,
  {32'h3eee4c49, 32'h3fb0bd40} /* (25, 18, 12) {real, imag} */,
  {32'hbf864bf2, 32'hbfed7c89} /* (25, 18, 11) {real, imag} */,
  {32'hbea47d0a, 32'h3fcc4da8} /* (25, 18, 10) {real, imag} */,
  {32'hbed2744f, 32'hbf0fb9e0} /* (25, 18, 9) {real, imag} */,
  {32'hbed67745, 32'hbfcda9a3} /* (25, 18, 8) {real, imag} */,
  {32'h3fd501c7, 32'h3fdcf48f} /* (25, 18, 7) {real, imag} */,
  {32'hc03d7015, 32'hbfa98cbe} /* (25, 18, 6) {real, imag} */,
  {32'h3ffe556b, 32'h407b378a} /* (25, 18, 5) {real, imag} */,
  {32'hbf23ce66, 32'h3fe68395} /* (25, 18, 4) {real, imag} */,
  {32'h3fcce273, 32'hbf888e98} /* (25, 18, 3) {real, imag} */,
  {32'h3ed1c043, 32'hbf67891c} /* (25, 18, 2) {real, imag} */,
  {32'hbe8ed0ef, 32'h3e15a1a1} /* (25, 18, 1) {real, imag} */,
  {32'hbf667ac2, 32'hbd992f4b} /* (25, 18, 0) {real, imag} */,
  {32'h3e831aa6, 32'h4029a2db} /* (25, 17, 31) {real, imag} */,
  {32'h3f0ff1a4, 32'h3f978770} /* (25, 17, 30) {real, imag} */,
  {32'h3f435af4, 32'h3eb7508b} /* (25, 17, 29) {real, imag} */,
  {32'h3efb557a, 32'h40081e1e} /* (25, 17, 28) {real, imag} */,
  {32'h3e876d37, 32'hbff9ec34} /* (25, 17, 27) {real, imag} */,
  {32'hbdbce961, 32'hbf3368e2} /* (25, 17, 26) {real, imag} */,
  {32'h4007dd80, 32'hc00b0c3d} /* (25, 17, 25) {real, imag} */,
  {32'hbd61144c, 32'h4009138e} /* (25, 17, 24) {real, imag} */,
  {32'h3fab7c65, 32'hbfff3ccf} /* (25, 17, 23) {real, imag} */,
  {32'hc01c61a6, 32'h3f42e323} /* (25, 17, 22) {real, imag} */,
  {32'hbe9ddd8b, 32'hbfb22cff} /* (25, 17, 21) {real, imag} */,
  {32'hbf8439b6, 32'h3f13e63a} /* (25, 17, 20) {real, imag} */,
  {32'h3e8c63df, 32'hbf98278b} /* (25, 17, 19) {real, imag} */,
  {32'hbfe277dd, 32'h3bede588} /* (25, 17, 18) {real, imag} */,
  {32'h3eec6bae, 32'h3f028615} /* (25, 17, 17) {real, imag} */,
  {32'hbda9cc77, 32'hbea4554b} /* (25, 17, 16) {real, imag} */,
  {32'h3f91f03c, 32'h3eba9a7c} /* (25, 17, 15) {real, imag} */,
  {32'h3fc39922, 32'hbf1ec5f8} /* (25, 17, 14) {real, imag} */,
  {32'h3f2e1f8d, 32'hbd783c9a} /* (25, 17, 13) {real, imag} */,
  {32'hbf26a59a, 32'hbf19f8ad} /* (25, 17, 12) {real, imag} */,
  {32'h40153ee6, 32'h3f9964f3} /* (25, 17, 11) {real, imag} */,
  {32'h3e86bc5f, 32'hc016d28b} /* (25, 17, 10) {real, imag} */,
  {32'h3f8d8c16, 32'h3fa18e99} /* (25, 17, 9) {real, imag} */,
  {32'hbf99b70b, 32'hbfb508f1} /* (25, 17, 8) {real, imag} */,
  {32'h405eacc1, 32'hbf20879c} /* (25, 17, 7) {real, imag} */,
  {32'hbd3d5b74, 32'h3fc36fea} /* (25, 17, 6) {real, imag} */,
  {32'h3b640088, 32'hbfca3336} /* (25, 17, 5) {real, imag} */,
  {32'hbe414179, 32'hbff4910a} /* (25, 17, 4) {real, imag} */,
  {32'hbe862136, 32'hbf034495} /* (25, 17, 3) {real, imag} */,
  {32'hbfb2f9da, 32'h3f27b1a8} /* (25, 17, 2) {real, imag} */,
  {32'h3f7b2db4, 32'h3f5d1e9d} /* (25, 17, 1) {real, imag} */,
  {32'hc0268683, 32'h3f329d11} /* (25, 17, 0) {real, imag} */,
  {32'hbff80ce5, 32'h3f8a7217} /* (25, 16, 31) {real, imag} */,
  {32'hbfd0a00f, 32'h3d80fa73} /* (25, 16, 30) {real, imag} */,
  {32'h3e81a4d1, 32'h3f043e83} /* (25, 16, 29) {real, imag} */,
  {32'hbe2afca9, 32'hbf3c9573} /* (25, 16, 28) {real, imag} */,
  {32'h3f23ccd1, 32'hbf53eb2c} /* (25, 16, 27) {real, imag} */,
  {32'h3ede3b84, 32'hbf1018ed} /* (25, 16, 26) {real, imag} */,
  {32'hc0122a6c, 32'hbbe52054} /* (25, 16, 25) {real, imag} */,
  {32'h3e456aa9, 32'hbfc232c7} /* (25, 16, 24) {real, imag} */,
  {32'h3e25f9b4, 32'hc0128930} /* (25, 16, 23) {real, imag} */,
  {32'hbf848481, 32'h401523b5} /* (25, 16, 22) {real, imag} */,
  {32'hbf2764eb, 32'hc00c599c} /* (25, 16, 21) {real, imag} */,
  {32'h3e8a2cb0, 32'hbe6b4a78} /* (25, 16, 20) {real, imag} */,
  {32'h3d9273be, 32'h3fc7d5d3} /* (25, 16, 19) {real, imag} */,
  {32'hbf006ce2, 32'h3f5eb722} /* (25, 16, 18) {real, imag} */,
  {32'h3f05ec40, 32'h3e3497fe} /* (25, 16, 17) {real, imag} */,
  {32'hbe9f30cd, 32'h3f4e425a} /* (25, 16, 16) {real, imag} */,
  {32'hbfd953f7, 32'hbea42a8c} /* (25, 16, 15) {real, imag} */,
  {32'hbf8f029d, 32'h3fa76cac} /* (25, 16, 14) {real, imag} */,
  {32'h3f9a0680, 32'h400e57ed} /* (25, 16, 13) {real, imag} */,
  {32'hbfc624e3, 32'h3f85be44} /* (25, 16, 12) {real, imag} */,
  {32'h3f6feefb, 32'hbf910997} /* (25, 16, 11) {real, imag} */,
  {32'h3f231a3a, 32'hbec9683c} /* (25, 16, 10) {real, imag} */,
  {32'hbe9b7a05, 32'h3f193395} /* (25, 16, 9) {real, imag} */,
  {32'h3f9f1295, 32'hbe5f0f1e} /* (25, 16, 8) {real, imag} */,
  {32'h3f23bcfd, 32'h3f522bf7} /* (25, 16, 7) {real, imag} */,
  {32'hbfecb8ed, 32'h3f8d8dfd} /* (25, 16, 6) {real, imag} */,
  {32'hbf2035cd, 32'h3d1b7da2} /* (25, 16, 5) {real, imag} */,
  {32'h401ec460, 32'hbcc53534} /* (25, 16, 4) {real, imag} */,
  {32'h3fbe6281, 32'h3f7fbcb4} /* (25, 16, 3) {real, imag} */,
  {32'hbfaf0435, 32'h3f9f4fc2} /* (25, 16, 2) {real, imag} */,
  {32'h3f97c8bd, 32'hbf6fb3b0} /* (25, 16, 1) {real, imag} */,
  {32'h3eb7f7ac, 32'hbcf99927} /* (25, 16, 0) {real, imag} */,
  {32'hb9c1e304, 32'hbf7a7696} /* (25, 15, 31) {real, imag} */,
  {32'h3f2284a5, 32'h401c1511} /* (25, 15, 30) {real, imag} */,
  {32'h3f3f6200, 32'h3f0755a2} /* (25, 15, 29) {real, imag} */,
  {32'hbf56352f, 32'h3e9ea328} /* (25, 15, 28) {real, imag} */,
  {32'hbf694bbb, 32'hbe01bb0e} /* (25, 15, 27) {real, imag} */,
  {32'hc01a8d6a, 32'hbffe4c24} /* (25, 15, 26) {real, imag} */,
  {32'hbeae7891, 32'h3f10c45f} /* (25, 15, 25) {real, imag} */,
  {32'hbed7cbd3, 32'hbf74d578} /* (25, 15, 24) {real, imag} */,
  {32'hbf34f635, 32'hc00ac1a1} /* (25, 15, 23) {real, imag} */,
  {32'h3e2d7dc7, 32'hbf13ad2f} /* (25, 15, 22) {real, imag} */,
  {32'h3e811573, 32'h3fa8a98a} /* (25, 15, 21) {real, imag} */,
  {32'hbf5c21bf, 32'h3f05d98e} /* (25, 15, 20) {real, imag} */,
  {32'h405706dc, 32'h3ff1c3bc} /* (25, 15, 19) {real, imag} */,
  {32'h3f911546, 32'hc0347030} /* (25, 15, 18) {real, imag} */,
  {32'h3fba0dcf, 32'hc001a687} /* (25, 15, 17) {real, imag} */,
  {32'h3fb9237f, 32'h3ed8a814} /* (25, 15, 16) {real, imag} */,
  {32'hbf166896, 32'hbf6629a9} /* (25, 15, 15) {real, imag} */,
  {32'h3fb42991, 32'hbd7a5fba} /* (25, 15, 14) {real, imag} */,
  {32'hbfb8ff5a, 32'hbff356bb} /* (25, 15, 13) {real, imag} */,
  {32'h3f364cd1, 32'hbf0bb3ee} /* (25, 15, 12) {real, imag} */,
  {32'hc05b5b37, 32'h3c916eba} /* (25, 15, 11) {real, imag} */,
  {32'hbf59370e, 32'h3f988d09} /* (25, 15, 10) {real, imag} */,
  {32'hbef9e0a7, 32'h3f06be46} /* (25, 15, 9) {real, imag} */,
  {32'h3f81070c, 32'h400e346b} /* (25, 15, 8) {real, imag} */,
  {32'h3ea3e728, 32'h3fbb78c5} /* (25, 15, 7) {real, imag} */,
  {32'h3ffaa34f, 32'hbfd5a930} /* (25, 15, 6) {real, imag} */,
  {32'h3e94c45a, 32'hbe02a6b6} /* (25, 15, 5) {real, imag} */,
  {32'h3ea37ec4, 32'hbf3c7c3e} /* (25, 15, 4) {real, imag} */,
  {32'hbf3aa749, 32'hbebaeb17} /* (25, 15, 3) {real, imag} */,
  {32'h3e360d5f, 32'h3e2da011} /* (25, 15, 2) {real, imag} */,
  {32'h3ef15289, 32'h3f486477} /* (25, 15, 1) {real, imag} */,
  {32'hc03876ba, 32'hbf497afe} /* (25, 15, 0) {real, imag} */,
  {32'hbf662bb9, 32'hbef0c974} /* (25, 14, 31) {real, imag} */,
  {32'h3eed62fd, 32'hbfaa0f87} /* (25, 14, 30) {real, imag} */,
  {32'hc0223d72, 32'h3ea20400} /* (25, 14, 29) {real, imag} */,
  {32'hbffb3af8, 32'h3fa869c8} /* (25, 14, 28) {real, imag} */,
  {32'hbe329080, 32'hbe6f3313} /* (25, 14, 27) {real, imag} */,
  {32'hbf877631, 32'h3fd23621} /* (25, 14, 26) {real, imag} */,
  {32'h3e5f59b1, 32'hc0564956} /* (25, 14, 25) {real, imag} */,
  {32'h3fdfb0d2, 32'hc009300b} /* (25, 14, 24) {real, imag} */,
  {32'h401e250c, 32'h3f0f00a3} /* (25, 14, 23) {real, imag} */,
  {32'h3fa9b172, 32'hbf9af729} /* (25, 14, 22) {real, imag} */,
  {32'h3fd96b3f, 32'h3ef7b129} /* (25, 14, 21) {real, imag} */,
  {32'h3fdf6a80, 32'hbf90d508} /* (25, 14, 20) {real, imag} */,
  {32'h3ffe6a6d, 32'h3edc09d4} /* (25, 14, 19) {real, imag} */,
  {32'h40796360, 32'hbf021318} /* (25, 14, 18) {real, imag} */,
  {32'hc003a7f0, 32'h3ee89d27} /* (25, 14, 17) {real, imag} */,
  {32'hbf8a56e9, 32'hbf723e58} /* (25, 14, 16) {real, imag} */,
  {32'hbe97cc0b, 32'hbfa05456} /* (25, 14, 15) {real, imag} */,
  {32'h3e2d2737, 32'hbe899ac5} /* (25, 14, 14) {real, imag} */,
  {32'h3fbbf043, 32'h3fa3010a} /* (25, 14, 13) {real, imag} */,
  {32'h3e9906f7, 32'h3f06037e} /* (25, 14, 12) {real, imag} */,
  {32'h3f622db0, 32'hbf5c267d} /* (25, 14, 11) {real, imag} */,
  {32'hbd13bf43, 32'h4085d41a} /* (25, 14, 10) {real, imag} */,
  {32'hbf75fbf6, 32'hbf8b220b} /* (25, 14, 9) {real, imag} */,
  {32'hbea58867, 32'hc01f9997} /* (25, 14, 8) {real, imag} */,
  {32'h3f01ae9a, 32'h3c209c8f} /* (25, 14, 7) {real, imag} */,
  {32'hc0173f50, 32'h3e347af2} /* (25, 14, 6) {real, imag} */,
  {32'hc04ea44b, 32'hc06b25d1} /* (25, 14, 5) {real, imag} */,
  {32'h3fa95a1e, 32'hbf9c3a2d} /* (25, 14, 4) {real, imag} */,
  {32'h3f4d6d30, 32'hbfbb7bef} /* (25, 14, 3) {real, imag} */,
  {32'hc01af198, 32'h3edca988} /* (25, 14, 2) {real, imag} */,
  {32'hbf9afbf9, 32'hbfaa0d60} /* (25, 14, 1) {real, imag} */,
  {32'h3fe5e6c2, 32'hbf3787a5} /* (25, 14, 0) {real, imag} */,
  {32'h3fa25e28, 32'h3e548924} /* (25, 13, 31) {real, imag} */,
  {32'h3f6fb035, 32'h4043ed04} /* (25, 13, 30) {real, imag} */,
  {32'hbf91308d, 32'hbfdeddd4} /* (25, 13, 29) {real, imag} */,
  {32'hbe57abb1, 32'hbf15eec7} /* (25, 13, 28) {real, imag} */,
  {32'hbf987d1b, 32'h3f0af0f9} /* (25, 13, 27) {real, imag} */,
  {32'h3f1673e2, 32'hc0164f26} /* (25, 13, 26) {real, imag} */,
  {32'h3f024e7a, 32'hbf069717} /* (25, 13, 25) {real, imag} */,
  {32'hbf79b1de, 32'h3f20ed1e} /* (25, 13, 24) {real, imag} */,
  {32'h3e8e7e07, 32'h3ef00bc2} /* (25, 13, 23) {real, imag} */,
  {32'h3f1f4344, 32'hbf297030} /* (25, 13, 22) {real, imag} */,
  {32'h3ff8721b, 32'hc009e436} /* (25, 13, 21) {real, imag} */,
  {32'h40cb9fbc, 32'hbe2103d7} /* (25, 13, 20) {real, imag} */,
  {32'hbed08cc3, 32'hc00323ee} /* (25, 13, 19) {real, imag} */,
  {32'h3e332537, 32'hbe59d887} /* (25, 13, 18) {real, imag} */,
  {32'hbe077a2e, 32'h400b8c51} /* (25, 13, 17) {real, imag} */,
  {32'h3f4baf5c, 32'h400e00e1} /* (25, 13, 16) {real, imag} */,
  {32'hbfbe03d8, 32'hbfc0088e} /* (25, 13, 15) {real, imag} */,
  {32'hbfd36005, 32'hbe01f51b} /* (25, 13, 14) {real, imag} */,
  {32'hbeeba876, 32'hbe631e52} /* (25, 13, 13) {real, imag} */,
  {32'hbed4ee49, 32'h3fd6137e} /* (25, 13, 12) {real, imag} */,
  {32'hbf857d93, 32'h3f11d507} /* (25, 13, 11) {real, imag} */,
  {32'h402deb20, 32'hbfee7d63} /* (25, 13, 10) {real, imag} */,
  {32'h3fc5c3db, 32'hbfa13dcd} /* (25, 13, 9) {real, imag} */,
  {32'hbe017fd9, 32'h3ead39ea} /* (25, 13, 8) {real, imag} */,
  {32'hc027e3f3, 32'hc0b1d856} /* (25, 13, 7) {real, imag} */,
  {32'hbf47a981, 32'h3f3924bb} /* (25, 13, 6) {real, imag} */,
  {32'hbf0ddcfe, 32'h3f1f3417} /* (25, 13, 5) {real, imag} */,
  {32'hbf23a618, 32'hbfeb17d8} /* (25, 13, 4) {real, imag} */,
  {32'hbf89aabf, 32'hbfd6ba76} /* (25, 13, 3) {real, imag} */,
  {32'h4084294f, 32'h3f840c9c} /* (25, 13, 2) {real, imag} */,
  {32'h3f262e97, 32'h3ff0d895} /* (25, 13, 1) {real, imag} */,
  {32'h3eb5398c, 32'h3ede21fe} /* (25, 13, 0) {real, imag} */,
  {32'hbf3af07c, 32'h3fe26905} /* (25, 12, 31) {real, imag} */,
  {32'h402821b8, 32'hbf40d907} /* (25, 12, 30) {real, imag} */,
  {32'hbf9ca249, 32'h3e55988b} /* (25, 12, 29) {real, imag} */,
  {32'h3e60f4be, 32'h402b78ad} /* (25, 12, 28) {real, imag} */,
  {32'h3ebcd6c9, 32'h3f2e195c} /* (25, 12, 27) {real, imag} */,
  {32'hc0432499, 32'h3e6e4534} /* (25, 12, 26) {real, imag} */,
  {32'h3fafc5ef, 32'hc04f6365} /* (25, 12, 25) {real, imag} */,
  {32'hc029b92c, 32'h3f28da70} /* (25, 12, 24) {real, imag} */,
  {32'hc049f94c, 32'hc0264cf7} /* (25, 12, 23) {real, imag} */,
  {32'hbeb7b1a4, 32'hbfb7fc28} /* (25, 12, 22) {real, imag} */,
  {32'hc0045569, 32'hbfbdaed7} /* (25, 12, 21) {real, imag} */,
  {32'hbfd5d06b, 32'h40a5364b} /* (25, 12, 20) {real, imag} */,
  {32'hbfd707d0, 32'h3fb3238f} /* (25, 12, 19) {real, imag} */,
  {32'hbf047930, 32'hbf7a7ef3} /* (25, 12, 18) {real, imag} */,
  {32'hbe7ef06e, 32'h3f888aba} /* (25, 12, 17) {real, imag} */,
  {32'h3fafa264, 32'hbe42cc09} /* (25, 12, 16) {real, imag} */,
  {32'hbfc0d69a, 32'h3fdf0c0f} /* (25, 12, 15) {real, imag} */,
  {32'hbeb0c5af, 32'hc0472c74} /* (25, 12, 14) {real, imag} */,
  {32'h3f0e0ad4, 32'h3e5fb4e4} /* (25, 12, 13) {real, imag} */,
  {32'hc080d573, 32'hc0021192} /* (25, 12, 12) {real, imag} */,
  {32'h3fb0f92a, 32'hbd6d9197} /* (25, 12, 11) {real, imag} */,
  {32'h3fa7722d, 32'hc0768dae} /* (25, 12, 10) {real, imag} */,
  {32'h3e856b01, 32'h3e8e0ddb} /* (25, 12, 9) {real, imag} */,
  {32'h3f513613, 32'hc08b0214} /* (25, 12, 8) {real, imag} */,
  {32'hbed2e008, 32'h3f722a60} /* (25, 12, 7) {real, imag} */,
  {32'hbfc02ce2, 32'hbf9e4b8d} /* (25, 12, 6) {real, imag} */,
  {32'h3fc0ad6b, 32'hbe2f8e16} /* (25, 12, 5) {real, imag} */,
  {32'h3e11cbfa, 32'h401aacff} /* (25, 12, 4) {real, imag} */,
  {32'h3fbb9325, 32'hbf8d93bd} /* (25, 12, 3) {real, imag} */,
  {32'hbebcfc20, 32'hbf38bb78} /* (25, 12, 2) {real, imag} */,
  {32'h3d918fd0, 32'h3e9ab044} /* (25, 12, 1) {real, imag} */,
  {32'h3f97e552, 32'hbf9d3c56} /* (25, 12, 0) {real, imag} */,
  {32'hbf59bd6f, 32'h3f1d2d3e} /* (25, 11, 31) {real, imag} */,
  {32'h3f9f0110, 32'h3ee4b66a} /* (25, 11, 30) {real, imag} */,
  {32'hc0218a65, 32'h3e2eb095} /* (25, 11, 29) {real, imag} */,
  {32'h400273bf, 32'hbec692c8} /* (25, 11, 28) {real, imag} */,
  {32'hbe5933c7, 32'h3fc135a4} /* (25, 11, 27) {real, imag} */,
  {32'h4009b8de, 32'h3fb596d2} /* (25, 11, 26) {real, imag} */,
  {32'h40358be4, 32'hbea2bc6d} /* (25, 11, 25) {real, imag} */,
  {32'hbff34f11, 32'h3f5c461d} /* (25, 11, 24) {real, imag} */,
  {32'h40639b7c, 32'hbec594da} /* (25, 11, 23) {real, imag} */,
  {32'h3f058c0d, 32'h3fd52d6c} /* (25, 11, 22) {real, imag} */,
  {32'hc00d2dfd, 32'h3f808387} /* (25, 11, 21) {real, imag} */,
  {32'hc01c233e, 32'hc00012ac} /* (25, 11, 20) {real, imag} */,
  {32'hbfaea4ab, 32'h3f3e32d2} /* (25, 11, 19) {real, imag} */,
  {32'hc0225058, 32'h40450dc8} /* (25, 11, 18) {real, imag} */,
  {32'hbec2fdc3, 32'hc0581fc3} /* (25, 11, 17) {real, imag} */,
  {32'hbf61a597, 32'h3fde0e2f} /* (25, 11, 16) {real, imag} */,
  {32'hc00af3fb, 32'h3ef9b51d} /* (25, 11, 15) {real, imag} */,
  {32'h3fccb2be, 32'hbf0d5a92} /* (25, 11, 14) {real, imag} */,
  {32'h4003ce88, 32'h3f97f2d0} /* (25, 11, 13) {real, imag} */,
  {32'hbfa23a02, 32'h401f0ac7} /* (25, 11, 12) {real, imag} */,
  {32'h4061c0fd, 32'hbf15e517} /* (25, 11, 11) {real, imag} */,
  {32'h3ea7a224, 32'hc0145936} /* (25, 11, 10) {real, imag} */,
  {32'h3fb09922, 32'h407dff7a} /* (25, 11, 9) {real, imag} */,
  {32'hc0149d5f, 32'hbf9dfb61} /* (25, 11, 8) {real, imag} */,
  {32'hbf437ee5, 32'hc0011797} /* (25, 11, 7) {real, imag} */,
  {32'h3fa46ec4, 32'h3ebd6389} /* (25, 11, 6) {real, imag} */,
  {32'hc076fc7d, 32'h3dcfe68e} /* (25, 11, 5) {real, imag} */,
  {32'h3f544c06, 32'hc00f0dc8} /* (25, 11, 4) {real, imag} */,
  {32'hbf3a7f20, 32'h3ff302e4} /* (25, 11, 3) {real, imag} */,
  {32'hbfaa6f32, 32'h3d404f0d} /* (25, 11, 2) {real, imag} */,
  {32'h403bf995, 32'h40281c4f} /* (25, 11, 1) {real, imag} */,
  {32'hbe36d0c6, 32'h3ef2d20c} /* (25, 11, 0) {real, imag} */,
  {32'h3dc81d00, 32'hbf35d16f} /* (25, 10, 31) {real, imag} */,
  {32'h3e11cd5f, 32'hc0aca365} /* (25, 10, 30) {real, imag} */,
  {32'hbf113990, 32'hbfa03c48} /* (25, 10, 29) {real, imag} */,
  {32'h3f9f7f62, 32'hc057c049} /* (25, 10, 28) {real, imag} */,
  {32'hbe0a7780, 32'h3f7455dc} /* (25, 10, 27) {real, imag} */,
  {32'h4007e108, 32'h3fcb18ba} /* (25, 10, 26) {real, imag} */,
  {32'h3cb2c4fe, 32'h405e8a9f} /* (25, 10, 25) {real, imag} */,
  {32'h3e030052, 32'h3f6cd4f3} /* (25, 10, 24) {real, imag} */,
  {32'h4060c6d7, 32'h408542cf} /* (25, 10, 23) {real, imag} */,
  {32'hc0807991, 32'hbfc441f8} /* (25, 10, 22) {real, imag} */,
  {32'hbf00dece, 32'h3e819277} /* (25, 10, 21) {real, imag} */,
  {32'h3fde7928, 32'hbca010c6} /* (25, 10, 20) {real, imag} */,
  {32'hbf593cf1, 32'hc01a08f9} /* (25, 10, 19) {real, imag} */,
  {32'hc006521a, 32'hbefad008} /* (25, 10, 18) {real, imag} */,
  {32'h3f155a2c, 32'hbf831a1a} /* (25, 10, 17) {real, imag} */,
  {32'h3f9a75a0, 32'hc02c1d35} /* (25, 10, 16) {real, imag} */,
  {32'hbf824fef, 32'hbf106367} /* (25, 10, 15) {real, imag} */,
  {32'h3edafee1, 32'hbfb00ecf} /* (25, 10, 14) {real, imag} */,
  {32'hbfff7609, 32'h40450184} /* (25, 10, 13) {real, imag} */,
  {32'h3fb118f6, 32'hc03cf0f3} /* (25, 10, 12) {real, imag} */,
  {32'h3f82231e, 32'h402675fe} /* (25, 10, 11) {real, imag} */,
  {32'hbf9e1d1d, 32'hbf573d1b} /* (25, 10, 10) {real, imag} */,
  {32'hbf4e0c87, 32'hc0535a25} /* (25, 10, 9) {real, imag} */,
  {32'h3e362b96, 32'h4009c2b4} /* (25, 10, 8) {real, imag} */,
  {32'hbdc5c2b8, 32'h3e91df38} /* (25, 10, 7) {real, imag} */,
  {32'hc02ca6ba, 32'h400b549e} /* (25, 10, 6) {real, imag} */,
  {32'hc00b7bc3, 32'hbf57fc91} /* (25, 10, 5) {real, imag} */,
  {32'h402bf9e0, 32'hc0055c6d} /* (25, 10, 4) {real, imag} */,
  {32'hc04029f9, 32'hc030f40a} /* (25, 10, 3) {real, imag} */,
  {32'h3fd37b96, 32'h4071d9d8} /* (25, 10, 2) {real, imag} */,
  {32'h3fdb5fb2, 32'h402480b0} /* (25, 10, 1) {real, imag} */,
  {32'h3e90b0cc, 32'h3fa4d4e3} /* (25, 10, 0) {real, imag} */,
  {32'h402287bb, 32'hc04295c9} /* (25, 9, 31) {real, imag} */,
  {32'h3fba631f, 32'hbf1b2d85} /* (25, 9, 30) {real, imag} */,
  {32'hbecb3d53, 32'h3dcf21d9} /* (25, 9, 29) {real, imag} */,
  {32'hbf544b44, 32'h3dbcc4d1} /* (25, 9, 28) {real, imag} */,
  {32'h3faa5e2b, 32'hbf0c2a22} /* (25, 9, 27) {real, imag} */,
  {32'hbeb620a8, 32'hbf759de7} /* (25, 9, 26) {real, imag} */,
  {32'hbe939064, 32'h40787d39} /* (25, 9, 25) {real, imag} */,
  {32'h401144d9, 32'hbe01e74e} /* (25, 9, 24) {real, imag} */,
  {32'h3f011a70, 32'hbea82b33} /* (25, 9, 23) {real, imag} */,
  {32'hbf3f3152, 32'hbf999b27} /* (25, 9, 22) {real, imag} */,
  {32'h3f2a71ff, 32'hbfa2a80d} /* (25, 9, 21) {real, imag} */,
  {32'hbefcafe0, 32'hbea4da65} /* (25, 9, 20) {real, imag} */,
  {32'hc09258fc, 32'hbdb4b317} /* (25, 9, 19) {real, imag} */,
  {32'hbf89432d, 32'h3f82aa9f} /* (25, 9, 18) {real, imag} */,
  {32'h3e0b1c4a, 32'h3ea24a9d} /* (25, 9, 17) {real, imag} */,
  {32'h3f60a407, 32'h3e406be1} /* (25, 9, 16) {real, imag} */,
  {32'h3f870cc0, 32'hc017a7a2} /* (25, 9, 15) {real, imag} */,
  {32'h3ecb6a11, 32'hc0380633} /* (25, 9, 14) {real, imag} */,
  {32'h4049b386, 32'h3f6555aa} /* (25, 9, 13) {real, imag} */,
  {32'hbfcb1f91, 32'h3f2404b4} /* (25, 9, 12) {real, imag} */,
  {32'hbe8ac951, 32'hbf94fa15} /* (25, 9, 11) {real, imag} */,
  {32'h40915297, 32'h3fb5f3a4} /* (25, 9, 10) {real, imag} */,
  {32'hc0891b86, 32'hc012b38e} /* (25, 9, 9) {real, imag} */,
  {32'h3fa1c425, 32'h3f953a26} /* (25, 9, 8) {real, imag} */,
  {32'h3de2bb33, 32'h3fa4cd42} /* (25, 9, 7) {real, imag} */,
  {32'hbfc737e8, 32'h405da5f9} /* (25, 9, 6) {real, imag} */,
  {32'hc02a38ee, 32'hbfb18aa0} /* (25, 9, 5) {real, imag} */,
  {32'h4040df5b, 32'hc0005af6} /* (25, 9, 4) {real, imag} */,
  {32'h3d6e8eb2, 32'h408a21fe} /* (25, 9, 3) {real, imag} */,
  {32'h405087c9, 32'h3fdd0dd7} /* (25, 9, 2) {real, imag} */,
  {32'hc0137502, 32'hc038c94a} /* (25, 9, 1) {real, imag} */,
  {32'hbf1da61d, 32'h3f37c8c9} /* (25, 9, 0) {real, imag} */,
  {32'hbf8ee309, 32'hbfdf9817} /* (25, 8, 31) {real, imag} */,
  {32'hc01d2db7, 32'hbeab2c8b} /* (25, 8, 30) {real, imag} */,
  {32'h4039f3c6, 32'h3f910dc0} /* (25, 8, 29) {real, imag} */,
  {32'hbffec264, 32'hc00e16f1} /* (25, 8, 28) {real, imag} */,
  {32'hc008191a, 32'hbedab1e6} /* (25, 8, 27) {real, imag} */,
  {32'hbf8aaa69, 32'hbffe393d} /* (25, 8, 26) {real, imag} */,
  {32'h4088d6b5, 32'h4013b311} /* (25, 8, 25) {real, imag} */,
  {32'hbfcd447b, 32'h3f964edf} /* (25, 8, 24) {real, imag} */,
  {32'hc05d8ea6, 32'h3f86c429} /* (25, 8, 23) {real, imag} */,
  {32'hc074ad83, 32'h4087adbf} /* (25, 8, 22) {real, imag} */,
  {32'h3eb2194c, 32'h3fdacd19} /* (25, 8, 21) {real, imag} */,
  {32'hbf874c59, 32'hc0893d08} /* (25, 8, 20) {real, imag} */,
  {32'h3fe03012, 32'h3fc2d7de} /* (25, 8, 19) {real, imag} */,
  {32'h3d8cb9f9, 32'hbd2d2ccd} /* (25, 8, 18) {real, imag} */,
  {32'h3f8a4fd2, 32'hc01349e4} /* (25, 8, 17) {real, imag} */,
  {32'h3e5b46d3, 32'hbe95b079} /* (25, 8, 16) {real, imag} */,
  {32'hbf2b55b9, 32'hbe5fa53c} /* (25, 8, 15) {real, imag} */,
  {32'hbd99ec20, 32'h40668c58} /* (25, 8, 14) {real, imag} */,
  {32'h3f43aa5e, 32'hbecc9e77} /* (25, 8, 13) {real, imag} */,
  {32'h3f2ad0c8, 32'hc02927cb} /* (25, 8, 12) {real, imag} */,
  {32'h3d904e1b, 32'hbefc1d03} /* (25, 8, 11) {real, imag} */,
  {32'hc0098752, 32'hbfc6d864} /* (25, 8, 10) {real, imag} */,
  {32'h3ebab182, 32'h3d1debbb} /* (25, 8, 9) {real, imag} */,
  {32'hbefd97f8, 32'h3f874c03} /* (25, 8, 8) {real, imag} */,
  {32'h4101ce9f, 32'h3eae6215} /* (25, 8, 7) {real, imag} */,
  {32'h4014f1c4, 32'h3faab159} /* (25, 8, 6) {real, imag} */,
  {32'h4064e831, 32'hc02c0855} /* (25, 8, 5) {real, imag} */,
  {32'h400ce7f1, 32'h3e5d07bf} /* (25, 8, 4) {real, imag} */,
  {32'h3f3e9cc2, 32'hc03b5d72} /* (25, 8, 3) {real, imag} */,
  {32'h3d23f5aa, 32'hc00ba12e} /* (25, 8, 2) {real, imag} */,
  {32'hc037661b, 32'h3fd27834} /* (25, 8, 1) {real, imag} */,
  {32'h3e912429, 32'h40801be2} /* (25, 8, 0) {real, imag} */,
  {32'hc034d32b, 32'hbdfc8988} /* (25, 7, 31) {real, imag} */,
  {32'hbfd850c5, 32'hbfe7a685} /* (25, 7, 30) {real, imag} */,
  {32'hbeffbd60, 32'hbf8e316f} /* (25, 7, 29) {real, imag} */,
  {32'h4042cb8a, 32'hc09023b1} /* (25, 7, 28) {real, imag} */,
  {32'hc0481e53, 32'h3e107608} /* (25, 7, 27) {real, imag} */,
  {32'h403ebdac, 32'hc04c3564} /* (25, 7, 26) {real, imag} */,
  {32'hbf1b2a95, 32'hc00524f1} /* (25, 7, 25) {real, imag} */,
  {32'hbf483117, 32'h3fc0fcfa} /* (25, 7, 24) {real, imag} */,
  {32'h3f373123, 32'hbf76bd35} /* (25, 7, 23) {real, imag} */,
  {32'h402fe286, 32'hc03907de} /* (25, 7, 22) {real, imag} */,
  {32'hc00bc072, 32'h3f875cc3} /* (25, 7, 21) {real, imag} */,
  {32'h40339067, 32'hc034c106} /* (25, 7, 20) {real, imag} */,
  {32'h3f95c039, 32'h402b94c7} /* (25, 7, 19) {real, imag} */,
  {32'h3f1fddbb, 32'hbd14a311} /* (25, 7, 18) {real, imag} */,
  {32'h40283944, 32'hbf002186} /* (25, 7, 17) {real, imag} */,
  {32'h401057f3, 32'hbf657e48} /* (25, 7, 16) {real, imag} */,
  {32'hbf2c2040, 32'hc012e86c} /* (25, 7, 15) {real, imag} */,
  {32'h3eef9cba, 32'h403262bb} /* (25, 7, 14) {real, imag} */,
  {32'hc063d9ab, 32'h3fb9a933} /* (25, 7, 13) {real, imag} */,
  {32'hbfc893b9, 32'h3fa784a3} /* (25, 7, 12) {real, imag} */,
  {32'h3d6a1faa, 32'hbe2e1fc0} /* (25, 7, 11) {real, imag} */,
  {32'hc010031c, 32'h3f259c04} /* (25, 7, 10) {real, imag} */,
  {32'h3f72c04d, 32'h4005451b} /* (25, 7, 9) {real, imag} */,
  {32'hbfc8bb9f, 32'hbfef260c} /* (25, 7, 8) {real, imag} */,
  {32'hbff8c758, 32'h3e5fc453} /* (25, 7, 7) {real, imag} */,
  {32'h3fee95e3, 32'h3fa2f374} /* (25, 7, 6) {real, imag} */,
  {32'h3d34f8aa, 32'hc00ee6c1} /* (25, 7, 5) {real, imag} */,
  {32'hc06a25e8, 32'h404e9404} /* (25, 7, 4) {real, imag} */,
  {32'h3fc44635, 32'hbfa664e7} /* (25, 7, 3) {real, imag} */,
  {32'hbfb15e50, 32'hbf8d2d8a} /* (25, 7, 2) {real, imag} */,
  {32'h4066b529, 32'hbfca23e8} /* (25, 7, 1) {real, imag} */,
  {32'h4000264f, 32'h3f599dbf} /* (25, 7, 0) {real, imag} */,
  {32'hbf35bb0e, 32'hbf19fd84} /* (25, 6, 31) {real, imag} */,
  {32'h3de6eea5, 32'hbe7d0efb} /* (25, 6, 30) {real, imag} */,
  {32'hc016845a, 32'hbfa59e29} /* (25, 6, 29) {real, imag} */,
  {32'hbf88f9e8, 32'h40870178} /* (25, 6, 28) {real, imag} */,
  {32'h401cdd73, 32'h3d2e1018} /* (25, 6, 27) {real, imag} */,
  {32'h3f8c5624, 32'hbfd1fee0} /* (25, 6, 26) {real, imag} */,
  {32'hc07046e4, 32'hbf4fc5d4} /* (25, 6, 25) {real, imag} */,
  {32'h3e728368, 32'hbfc47650} /* (25, 6, 24) {real, imag} */,
  {32'hc04525c2, 32'h3d9e1569} /* (25, 6, 23) {real, imag} */,
  {32'hbd0d4d99, 32'hbf9460b5} /* (25, 6, 22) {real, imag} */,
  {32'hbf44a57f, 32'hc0055130} /* (25, 6, 21) {real, imag} */,
  {32'hbf488a66, 32'h40376fd6} /* (25, 6, 20) {real, imag} */,
  {32'h40898a11, 32'h3fba6daf} /* (25, 6, 19) {real, imag} */,
  {32'h4010e53d, 32'hbf9073d9} /* (25, 6, 18) {real, imag} */,
  {32'hbf036fdb, 32'hbf135e27} /* (25, 6, 17) {real, imag} */,
  {32'hbf926d46, 32'h3fb97530} /* (25, 6, 16) {real, imag} */,
  {32'h3e900ffe, 32'hbf3f5571} /* (25, 6, 15) {real, imag} */,
  {32'hbfd10fc3, 32'hc018bfda} /* (25, 6, 14) {real, imag} */,
  {32'hbff40732, 32'h3d9a4371} /* (25, 6, 13) {real, imag} */,
  {32'h40701070, 32'h3fb220d4} /* (25, 6, 12) {real, imag} */,
  {32'hbe9c5afb, 32'h405a0f47} /* (25, 6, 11) {real, imag} */,
  {32'hc03c049b, 32'h404e663f} /* (25, 6, 10) {real, imag} */,
  {32'h3e4941a2, 32'hbfbd7ecf} /* (25, 6, 9) {real, imag} */,
  {32'hbf9e549c, 32'hbc050659} /* (25, 6, 8) {real, imag} */,
  {32'h40205d4a, 32'h3fad8b31} /* (25, 6, 7) {real, imag} */,
  {32'hc016d649, 32'h40013895} /* (25, 6, 6) {real, imag} */,
  {32'hc002e719, 32'h402cfe3e} /* (25, 6, 5) {real, imag} */,
  {32'hc04919a3, 32'h3ebb88a5} /* (25, 6, 4) {real, imag} */,
  {32'h3f80a608, 32'hbfbba8cd} /* (25, 6, 3) {real, imag} */,
  {32'hbe8e1bbc, 32'h3f60c3ee} /* (25, 6, 2) {real, imag} */,
  {32'hc03b792f, 32'hc05c08c3} /* (25, 6, 1) {real, imag} */,
  {32'hbceb9042, 32'hbee33e1a} /* (25, 6, 0) {real, imag} */,
  {32'hc0720a53, 32'h40485b11} /* (25, 5, 31) {real, imag} */,
  {32'hc07db18d, 32'h40185c1a} /* (25, 5, 30) {real, imag} */,
  {32'hbec1525b, 32'hc02517d8} /* (25, 5, 29) {real, imag} */,
  {32'hc029aee3, 32'hc0ab7e79} /* (25, 5, 28) {real, imag} */,
  {32'hc0199c66, 32'hbed1dfe8} /* (25, 5, 27) {real, imag} */,
  {32'h40855bfa, 32'h40ab1488} /* (25, 5, 26) {real, imag} */,
  {32'h3f238a05, 32'hbfe369b1} /* (25, 5, 25) {real, imag} */,
  {32'hbe31e65e, 32'hc03fef90} /* (25, 5, 24) {real, imag} */,
  {32'h40394646, 32'h3f6d576d} /* (25, 5, 23) {real, imag} */,
  {32'hc038eecb, 32'hc0162d06} /* (25, 5, 22) {real, imag} */,
  {32'h3fe5848d, 32'h3f7fa0f7} /* (25, 5, 21) {real, imag} */,
  {32'hbfced8dd, 32'hc008dbf8} /* (25, 5, 20) {real, imag} */,
  {32'hbfcbb8da, 32'h3f7f6ae8} /* (25, 5, 19) {real, imag} */,
  {32'h3d59f182, 32'h3e31fd63} /* (25, 5, 18) {real, imag} */,
  {32'h3f185986, 32'h3e524a8e} /* (25, 5, 17) {real, imag} */,
  {32'hbf27abc3, 32'h3f286e1e} /* (25, 5, 16) {real, imag} */,
  {32'hbe556e1c, 32'h3dfca2b6} /* (25, 5, 15) {real, imag} */,
  {32'h403f747b, 32'h3ed3fa3c} /* (25, 5, 14) {real, imag} */,
  {32'h3f1f9a8c, 32'h3f4936ad} /* (25, 5, 13) {real, imag} */,
  {32'hbfc147c5, 32'hbf9febb3} /* (25, 5, 12) {real, imag} */,
  {32'hbfe46ccb, 32'h3fa8b3fd} /* (25, 5, 11) {real, imag} */,
  {32'h3c6a9c97, 32'h3f0fa9e5} /* (25, 5, 10) {real, imag} */,
  {32'h3fc29a73, 32'hc0ae67fa} /* (25, 5, 9) {real, imag} */,
  {32'hbfd8510b, 32'hbea1a95c} /* (25, 5, 8) {real, imag} */,
  {32'h3ef0185d, 32'hbfeac28a} /* (25, 5, 7) {real, imag} */,
  {32'h3e79655b, 32'h3f2564c2} /* (25, 5, 6) {real, imag} */,
  {32'h3eac8b80, 32'hc0113fe1} /* (25, 5, 5) {real, imag} */,
  {32'hbe8ea19f, 32'h40b92a0d} /* (25, 5, 4) {real, imag} */,
  {32'h3faceb19, 32'h4027a32c} /* (25, 5, 3) {real, imag} */,
  {32'h3f713ea1, 32'hbff0373c} /* (25, 5, 2) {real, imag} */,
  {32'hc03fbc73, 32'hc056ff46} /* (25, 5, 1) {real, imag} */,
  {32'h407281a3, 32'hc0756d0d} /* (25, 5, 0) {real, imag} */,
  {32'hbf8afdc5, 32'h3fa31a5b} /* (25, 4, 31) {real, imag} */,
  {32'h3c42d5f9, 32'h4004103e} /* (25, 4, 30) {real, imag} */,
  {32'h3f4886bc, 32'hbfc2225a} /* (25, 4, 29) {real, imag} */,
  {32'h4008dd6b, 32'h3e696de1} /* (25, 4, 28) {real, imag} */,
  {32'hbfcac4a3, 32'hc0004c77} /* (25, 4, 27) {real, imag} */,
  {32'hbfa38abb, 32'h40ad94f4} /* (25, 4, 26) {real, imag} */,
  {32'hbeab315d, 32'h3ec52236} /* (25, 4, 25) {real, imag} */,
  {32'hbfb40e98, 32'h3f40f46b} /* (25, 4, 24) {real, imag} */,
  {32'h3fcc925e, 32'h40116460} /* (25, 4, 23) {real, imag} */,
  {32'h3f669aae, 32'hc005facc} /* (25, 4, 22) {real, imag} */,
  {32'h402e0489, 32'h4025f0c6} /* (25, 4, 21) {real, imag} */,
  {32'hbe9f457f, 32'hbf4418b5} /* (25, 4, 20) {real, imag} */,
  {32'h3e79e616, 32'hc0266743} /* (25, 4, 19) {real, imag} */,
  {32'hbf1f3712, 32'hbf0709ff} /* (25, 4, 18) {real, imag} */,
  {32'hbeb2a973, 32'hbde4afa5} /* (25, 4, 17) {real, imag} */,
  {32'hbf8c2c54, 32'hbff2406c} /* (25, 4, 16) {real, imag} */,
  {32'h3f228e00, 32'hbf749824} /* (25, 4, 15) {real, imag} */,
  {32'hbf6e8591, 32'h3f8477dd} /* (25, 4, 14) {real, imag} */,
  {32'h3fadfc82, 32'h3fbec6c0} /* (25, 4, 13) {real, imag} */,
  {32'hbfea598b, 32'hbf554d1e} /* (25, 4, 12) {real, imag} */,
  {32'hc02bae47, 32'hbf5ac2b1} /* (25, 4, 11) {real, imag} */,
  {32'h4078b98c, 32'h3f1b4cf3} /* (25, 4, 10) {real, imag} */,
  {32'h401c334e, 32'h3e951e92} /* (25, 4, 9) {real, imag} */,
  {32'hc02c053c, 32'hc04ec698} /* (25, 4, 8) {real, imag} */,
  {32'h3f3606ab, 32'hc010762f} /* (25, 4, 7) {real, imag} */,
  {32'hbd1c1a5d, 32'hc062e029} /* (25, 4, 6) {real, imag} */,
  {32'hc054cccf, 32'h3e8f006e} /* (25, 4, 5) {real, imag} */,
  {32'h4097ffdf, 32'h3e25ad08} /* (25, 4, 4) {real, imag} */,
  {32'h3f3947e7, 32'h40660463} /* (25, 4, 3) {real, imag} */,
  {32'hbf8d3102, 32'hbfd7acfb} /* (25, 4, 2) {real, imag} */,
  {32'hbf800a15, 32'hc0347513} /* (25, 4, 1) {real, imag} */,
  {32'h3f5ff2dc, 32'h40994c7c} /* (25, 4, 0) {real, imag} */,
  {32'hbfbcb86f, 32'hbf92d748} /* (25, 3, 31) {real, imag} */,
  {32'h3f67d955, 32'h3fb6ea18} /* (25, 3, 30) {real, imag} */,
  {32'h3f7ea417, 32'hbb94497a} /* (25, 3, 29) {real, imag} */,
  {32'hc017ebe2, 32'h3fa3bcbe} /* (25, 3, 28) {real, imag} */,
  {32'hbf7959e5, 32'hc0bf3dfb} /* (25, 3, 27) {real, imag} */,
  {32'hc028d608, 32'h3e6d5bf1} /* (25, 3, 26) {real, imag} */,
  {32'h400080b8, 32'hc05ec89a} /* (25, 3, 25) {real, imag} */,
  {32'h3faa5918, 32'hbf84dc9a} /* (25, 3, 24) {real, imag} */,
  {32'hbff0c34a, 32'h40216c6e} /* (25, 3, 23) {real, imag} */,
  {32'hbe8b299f, 32'hbfb13bb7} /* (25, 3, 22) {real, imag} */,
  {32'hbfa70fd9, 32'hc019cbf9} /* (25, 3, 21) {real, imag} */,
  {32'hbeba95ab, 32'hc0251d64} /* (25, 3, 20) {real, imag} */,
  {32'hbeb18947, 32'hbfae9cf4} /* (25, 3, 19) {real, imag} */,
  {32'hbd833d21, 32'h40372b1d} /* (25, 3, 18) {real, imag} */,
  {32'hbf9f0acb, 32'hbf98f736} /* (25, 3, 17) {real, imag} */,
  {32'h3fae9413, 32'hbf1b55bf} /* (25, 3, 16) {real, imag} */,
  {32'h3f186b3a, 32'hbdd57f25} /* (25, 3, 15) {real, imag} */,
  {32'hbf607120, 32'h3fb19713} /* (25, 3, 14) {real, imag} */,
  {32'hbe061ac6, 32'hbfc94652} /* (25, 3, 13) {real, imag} */,
  {32'hbf0febdd, 32'hbbe703ab} /* (25, 3, 12) {real, imag} */,
  {32'h3e115a20, 32'h3f17388b} /* (25, 3, 11) {real, imag} */,
  {32'hbfed66db, 32'h406b0d21} /* (25, 3, 10) {real, imag} */,
  {32'h3fc49393, 32'hbf49c880} /* (25, 3, 9) {real, imag} */,
  {32'h3f1ab382, 32'hbc3427f9} /* (25, 3, 8) {real, imag} */,
  {32'hc04dd678, 32'hbf32882b} /* (25, 3, 7) {real, imag} */,
  {32'h3ee35f1a, 32'hc094bdc4} /* (25, 3, 6) {real, imag} */,
  {32'h40a3f6f6, 32'h3f43d54f} /* (25, 3, 5) {real, imag} */,
  {32'hc007f4f2, 32'h3f94fcc1} /* (25, 3, 4) {real, imag} */,
  {32'hc02a712f, 32'h3f6b5194} /* (25, 3, 3) {real, imag} */,
  {32'hc0a0f453, 32'h3ee710bf} /* (25, 3, 2) {real, imag} */,
  {32'h3f0fd115, 32'hbfdf7a81} /* (25, 3, 1) {real, imag} */,
  {32'hc0b21258, 32'hc01a3c4c} /* (25, 3, 0) {real, imag} */,
  {32'h408aa45f, 32'hc098329c} /* (25, 2, 31) {real, imag} */,
  {32'h3f0b72f8, 32'hc0b2023a} /* (25, 2, 30) {real, imag} */,
  {32'h405bfcb1, 32'h40215fcf} /* (25, 2, 29) {real, imag} */,
  {32'hc051e869, 32'h40976d45} /* (25, 2, 28) {real, imag} */,
  {32'h3ee0dc9a, 32'h3f15179d} /* (25, 2, 27) {real, imag} */,
  {32'hc0c1711c, 32'hbde3b5aa} /* (25, 2, 26) {real, imag} */,
  {32'hc0006a83, 32'hbfbe6090} /* (25, 2, 25) {real, imag} */,
  {32'h3f922a96, 32'h3f40fd02} /* (25, 2, 24) {real, imag} */,
  {32'h3f9e8aba, 32'hbec566c7} /* (25, 2, 23) {real, imag} */,
  {32'h403ca5ae, 32'h401f28a5} /* (25, 2, 22) {real, imag} */,
  {32'h3dc28706, 32'hbf15f0b1} /* (25, 2, 21) {real, imag} */,
  {32'hbede4394, 32'h3ec6b798} /* (25, 2, 20) {real, imag} */,
  {32'hbea63fe0, 32'h3d6c7ca7} /* (25, 2, 19) {real, imag} */,
  {32'h405541c9, 32'hbedccee1} /* (25, 2, 18) {real, imag} */,
  {32'h3f94a303, 32'hbfd30bae} /* (25, 2, 17) {real, imag} */,
  {32'h3f8129b8, 32'hbf1ee425} /* (25, 2, 16) {real, imag} */,
  {32'h3fc03d62, 32'h3fbdf331} /* (25, 2, 15) {real, imag} */,
  {32'hbee92878, 32'hbe5ba02e} /* (25, 2, 14) {real, imag} */,
  {32'hbf33e7dd, 32'hbf8a925b} /* (25, 2, 13) {real, imag} */,
  {32'hbf633759, 32'hc076ccbb} /* (25, 2, 12) {real, imag} */,
  {32'hbf73e0de, 32'hbff8a3b5} /* (25, 2, 11) {real, imag} */,
  {32'hc0219a48, 32'hc0589fe4} /* (25, 2, 10) {real, imag} */,
  {32'hbfd79df7, 32'h4037d647} /* (25, 2, 9) {real, imag} */,
  {32'h401ad3e7, 32'h3fbc43bf} /* (25, 2, 8) {real, imag} */,
  {32'hc08f712b, 32'h4034d699} /* (25, 2, 7) {real, imag} */,
  {32'h40700ad4, 32'hbea14461} /* (25, 2, 6) {real, imag} */,
  {32'h3fe0f596, 32'hbf2c02c5} /* (25, 2, 5) {real, imag} */,
  {32'hbf8fbde9, 32'h4016e88b} /* (25, 2, 4) {real, imag} */,
  {32'h3f86a6ec, 32'h40879d66} /* (25, 2, 3) {real, imag} */,
  {32'hbf813f21, 32'h3eba3ebf} /* (25, 2, 2) {real, imag} */,
  {32'hbfe79119, 32'hbf92dbe8} /* (25, 2, 1) {real, imag} */,
  {32'hc04bdd0b, 32'hc1062499} /* (25, 2, 0) {real, imag} */,
  {32'hbfe2bdb8, 32'hc027109d} /* (25, 1, 31) {real, imag} */,
  {32'h3f8cfb77, 32'hc0bf5f84} /* (25, 1, 30) {real, imag} */,
  {32'hbbec520d, 32'h40171c6d} /* (25, 1, 29) {real, imag} */,
  {32'hc0a68f88, 32'h40970734} /* (25, 1, 28) {real, imag} */,
  {32'hc05213bc, 32'hbf496679} /* (25, 1, 27) {real, imag} */,
  {32'h3fb68ae1, 32'hc02372a8} /* (25, 1, 26) {real, imag} */,
  {32'hc0258f50, 32'h3ea5b3f2} /* (25, 1, 25) {real, imag} */,
  {32'hbf18776f, 32'hbf871c2f} /* (25, 1, 24) {real, imag} */,
  {32'h3e84f333, 32'hbfb37ced} /* (25, 1, 23) {real, imag} */,
  {32'hc01999c7, 32'h3f2e109f} /* (25, 1, 22) {real, imag} */,
  {32'hbfc110d1, 32'hbffc17f1} /* (25, 1, 21) {real, imag} */,
  {32'hbf8d3655, 32'hbee6f24d} /* (25, 1, 20) {real, imag} */,
  {32'h3f8d5a4c, 32'hbf886406} /* (25, 1, 19) {real, imag} */,
  {32'h3ff1fde2, 32'hbfb045b2} /* (25, 1, 18) {real, imag} */,
  {32'h3f27a5ea, 32'hbe22938b} /* (25, 1, 17) {real, imag} */,
  {32'h3f262fb5, 32'h3e364841} /* (25, 1, 16) {real, imag} */,
  {32'h3f382851, 32'h3f56d160} /* (25, 1, 15) {real, imag} */,
  {32'h3fa10d92, 32'h3ef20f97} /* (25, 1, 14) {real, imag} */,
  {32'h3fc2d836, 32'h3fa1c604} /* (25, 1, 13) {real, imag} */,
  {32'h3ecb01ee, 32'hbff0cb9c} /* (25, 1, 12) {real, imag} */,
  {32'h3f61b173, 32'hbf376f89} /* (25, 1, 11) {real, imag} */,
  {32'h401dff51, 32'h3ec4ed4d} /* (25, 1, 10) {real, imag} */,
  {32'hc0a4dc9a, 32'h3e8ed65a} /* (25, 1, 9) {real, imag} */,
  {32'h40369024, 32'h3f8e8671} /* (25, 1, 8) {real, imag} */,
  {32'hbecff1c8, 32'hbe991447} /* (25, 1, 7) {real, imag} */,
  {32'hbf0d4940, 32'hc085246d} /* (25, 1, 6) {real, imag} */,
  {32'h400d777a, 32'hc070cacc} /* (25, 1, 5) {real, imag} */,
  {32'h3f1acaa7, 32'h40a3e10e} /* (25, 1, 4) {real, imag} */,
  {32'hc10aee11, 32'h3fa2da0b} /* (25, 1, 3) {real, imag} */,
  {32'h409be686, 32'hc04c82c3} /* (25, 1, 2) {real, imag} */,
  {32'h4068e8f7, 32'h40cb8ad7} /* (25, 1, 1) {real, imag} */,
  {32'hc06de830, 32'h40592fd6} /* (25, 1, 0) {real, imag} */,
  {32'h40215e4a, 32'hbfd92793} /* (25, 0, 31) {real, imag} */,
  {32'hbfc9992d, 32'h40af316a} /* (25, 0, 30) {real, imag} */,
  {32'h404db148, 32'hbfceeaa4} /* (25, 0, 29) {real, imag} */,
  {32'h4098350f, 32'hc081118b} /* (25, 0, 28) {real, imag} */,
  {32'hc067b81c, 32'h3e9d8e39} /* (25, 0, 27) {real, imag} */,
  {32'h40584196, 32'h3f2a0ad3} /* (25, 0, 26) {real, imag} */,
  {32'hbf532a8e, 32'h4023aabd} /* (25, 0, 25) {real, imag} */,
  {32'h4000e5e6, 32'h3f895439} /* (25, 0, 24) {real, imag} */,
  {32'hbea07ab2, 32'hc01a5b47} /* (25, 0, 23) {real, imag} */,
  {32'hbe2481f8, 32'h3fb968d7} /* (25, 0, 22) {real, imag} */,
  {32'hc02726a4, 32'h3fc4fcdd} /* (25, 0, 21) {real, imag} */,
  {32'h3e917c57, 32'h40879cbb} /* (25, 0, 20) {real, imag} */,
  {32'hbfce0a37, 32'hc03c9796} /* (25, 0, 19) {real, imag} */,
  {32'h3f7306fc, 32'h3f16bda2} /* (25, 0, 18) {real, imag} */,
  {32'hbf6faf1f, 32'h3fc2275f} /* (25, 0, 17) {real, imag} */,
  {32'hbf89737c, 32'h3f9c7286} /* (25, 0, 16) {real, imag} */,
  {32'hbfea1094, 32'hc04d2377} /* (25, 0, 15) {real, imag} */,
  {32'hbeca1760, 32'h3e79220f} /* (25, 0, 14) {real, imag} */,
  {32'h3fddd953, 32'hbdf4e206} /* (25, 0, 13) {real, imag} */,
  {32'h3fc8cd3d, 32'hbf867565} /* (25, 0, 12) {real, imag} */,
  {32'h3f95c853, 32'h3fa24fd5} /* (25, 0, 11) {real, imag} */,
  {32'hc06963cd, 32'h3c837845} /* (25, 0, 10) {real, imag} */,
  {32'hbfa9afed, 32'h3f07a34a} /* (25, 0, 9) {real, imag} */,
  {32'h3fc5f2c2, 32'hc02e0a14} /* (25, 0, 8) {real, imag} */,
  {32'h3f1aaa81, 32'h3bef4a07} /* (25, 0, 7) {real, imag} */,
  {32'h408d96a7, 32'h3fcba01b} /* (25, 0, 6) {real, imag} */,
  {32'hbf689f13, 32'hc0694b1d} /* (25, 0, 5) {real, imag} */,
  {32'hbfe22fa1, 32'hc0b5d2c9} /* (25, 0, 4) {real, imag} */,
  {32'hbfbe7592, 32'hbfc9b686} /* (25, 0, 3) {real, imag} */,
  {32'hbf386261, 32'hbf9f3684} /* (25, 0, 2) {real, imag} */,
  {32'hbc38e6f5, 32'hc0596853} /* (25, 0, 1) {real, imag} */,
  {32'hbe9f7d7b, 32'h40c1131b} /* (25, 0, 0) {real, imag} */,
  {32'hc1d113d0, 32'hc0be6938} /* (24, 31, 31) {real, imag} */,
  {32'h418f193a, 32'h401920a2} /* (24, 31, 30) {real, imag} */,
  {32'h3fd1614c, 32'hbfe58171} /* (24, 31, 29) {real, imag} */,
  {32'h3f9a7777, 32'h40bc6560} /* (24, 31, 28) {real, imag} */,
  {32'h40ebcf1f, 32'h3f368d25} /* (24, 31, 27) {real, imag} */,
  {32'h3fe642a9, 32'hbfc18be2} /* (24, 31, 26) {real, imag} */,
  {32'hc0c442bb, 32'h3f6b9e72} /* (24, 31, 25) {real, imag} */,
  {32'h40a13655, 32'hbefe2e55} /* (24, 31, 24) {real, imag} */,
  {32'h3d52b90d, 32'h402c88d2} /* (24, 31, 23) {real, imag} */,
  {32'hbce7a44c, 32'hc022094d} /* (24, 31, 22) {real, imag} */,
  {32'h3f1c52cb, 32'hbf933ad1} /* (24, 31, 21) {real, imag} */,
  {32'hc015236b, 32'h40919868} /* (24, 31, 20) {real, imag} */,
  {32'hbfacb9cb, 32'hbe984056} /* (24, 31, 19) {real, imag} */,
  {32'h3f6625c5, 32'hbf701cff} /* (24, 31, 18) {real, imag} */,
  {32'h3e1ceff0, 32'hbf54ef32} /* (24, 31, 17) {real, imag} */,
  {32'h3e999674, 32'hbddee17a} /* (24, 31, 16) {real, imag} */,
  {32'h3eeb19c7, 32'hbedeb623} /* (24, 31, 15) {real, imag} */,
  {32'h3ff8cb82, 32'h3f6fe752} /* (24, 31, 14) {real, imag} */,
  {32'hc041e14e, 32'hbe97b355} /* (24, 31, 13) {real, imag} */,
  {32'hc022e245, 32'h401d890c} /* (24, 31, 12) {real, imag} */,
  {32'hbf9f6ecc, 32'h40ae318e} /* (24, 31, 11) {real, imag} */,
  {32'hc016eb8d, 32'hbf21b606} /* (24, 31, 10) {real, imag} */,
  {32'hbddf95a5, 32'hc011f28f} /* (24, 31, 9) {real, imag} */,
  {32'hbf834267, 32'h409c8e4e} /* (24, 31, 8) {real, imag} */,
  {32'hc0acfdba, 32'hbec1145b} /* (24, 31, 7) {real, imag} */,
  {32'hc003e4b5, 32'hc007aa44} /* (24, 31, 6) {real, imag} */,
  {32'h4067a85b, 32'h408d3bcd} /* (24, 31, 5) {real, imag} */,
  {32'hc0020e1d, 32'h3fe73d4c} /* (24, 31, 4) {real, imag} */,
  {32'h3e833c93, 32'hbff07022} /* (24, 31, 3) {real, imag} */,
  {32'hbf850bac, 32'h40eaa787} /* (24, 31, 2) {real, imag} */,
  {32'hc147f7b4, 32'hc18d40ad} /* (24, 31, 1) {real, imag} */,
  {32'hc11b6bdf, 32'hc14197be} /* (24, 31, 0) {real, imag} */,
  {32'h41377b40, 32'h413ddd4c} /* (24, 30, 31) {real, imag} */,
  {32'hc02e38c4, 32'hc0a92edc} /* (24, 30, 30) {real, imag} */,
  {32'h3f0c0ff0, 32'h3ff0ba2f} /* (24, 30, 29) {real, imag} */,
  {32'h40b5338d, 32'h40aec42f} /* (24, 30, 28) {real, imag} */,
  {32'hc0b39358, 32'h3ff2ffb4} /* (24, 30, 27) {real, imag} */,
  {32'h402fbc48, 32'hbef82051} /* (24, 30, 26) {real, imag} */,
  {32'h3f6c0b40, 32'h3ec4c56e} /* (24, 30, 25) {real, imag} */,
  {32'hc0a93501, 32'hbfa62ed5} /* (24, 30, 24) {real, imag} */,
  {32'hc01b0b8e, 32'hbeaf3b58} /* (24, 30, 23) {real, imag} */,
  {32'hbf6c0ee3, 32'h3f49f4d7} /* (24, 30, 22) {real, imag} */,
  {32'hc07d8d66, 32'h40608f29} /* (24, 30, 21) {real, imag} */,
  {32'hbfa7470d, 32'h3e7aef39} /* (24, 30, 20) {real, imag} */,
  {32'hbe771607, 32'h3fe483ef} /* (24, 30, 19) {real, imag} */,
  {32'hc01e1211, 32'hbf8f2e45} /* (24, 30, 18) {real, imag} */,
  {32'hbaab9847, 32'hc01d3488} /* (24, 30, 17) {real, imag} */,
  {32'hbf90ac27, 32'hbddc047a} /* (24, 30, 16) {real, imag} */,
  {32'hc01d141e, 32'hbf35fcd9} /* (24, 30, 15) {real, imag} */,
  {32'hbee81c9d, 32'hbea420e6} /* (24, 30, 14) {real, imag} */,
  {32'hbfb43e18, 32'h3f1bbd2e} /* (24, 30, 13) {real, imag} */,
  {32'h3f6fcc0b, 32'h3fbdce65} /* (24, 30, 12) {real, imag} */,
  {32'h3df24f8b, 32'hbf127d44} /* (24, 30, 11) {real, imag} */,
  {32'h3f9a1990, 32'h3e2bdbf7} /* (24, 30, 10) {real, imag} */,
  {32'h3f143e2d, 32'hbf8e8829} /* (24, 30, 9) {real, imag} */,
  {32'h3c56737c, 32'hc099a259} /* (24, 30, 8) {real, imag} */,
  {32'h3faf3379, 32'h3f8c70e9} /* (24, 30, 7) {real, imag} */,
  {32'hbf8dbe7e, 32'hbffead18} /* (24, 30, 6) {real, imag} */,
  {32'hbf22d783, 32'h3ee1a093} /* (24, 30, 5) {real, imag} */,
  {32'hbf9b82ce, 32'h3fa5a21c} /* (24, 30, 4) {real, imag} */,
  {32'hbfc37788, 32'h404da494} /* (24, 30, 3) {real, imag} */,
  {32'hc1221985, 32'hc1418729} /* (24, 30, 2) {real, imag} */,
  {32'h418a52a7, 32'h413f6e8b} /* (24, 30, 1) {real, imag} */,
  {32'h413aa1d1, 32'h40edd0d4} /* (24, 30, 0) {real, imag} */,
  {32'hc0b46bec, 32'hbf7af1c3} /* (24, 29, 31) {real, imag} */,
  {32'h40b25e52, 32'hbf605d75} /* (24, 29, 30) {real, imag} */,
  {32'h3fb264fd, 32'h3f0dd07a} /* (24, 29, 29) {real, imag} */,
  {32'h40049929, 32'h3fcbbfed} /* (24, 29, 28) {real, imag} */,
  {32'h3fa69ad1, 32'hbf5b36ff} /* (24, 29, 27) {real, imag} */,
  {32'hc00da0b2, 32'hbfcfc726} /* (24, 29, 26) {real, imag} */,
  {32'hbebf2ac9, 32'h406364d2} /* (24, 29, 25) {real, imag} */,
  {32'h3fe109ae, 32'hc058b63d} /* (24, 29, 24) {real, imag} */,
  {32'hc08634e1, 32'hc079383e} /* (24, 29, 23) {real, imag} */,
  {32'h3ff59577, 32'h401d2d40} /* (24, 29, 22) {real, imag} */,
  {32'h40020bad, 32'h3fac8376} /* (24, 29, 21) {real, imag} */,
  {32'h3fdc1dff, 32'h3fcaa280} /* (24, 29, 20) {real, imag} */,
  {32'hbff7bfd9, 32'h3fa54964} /* (24, 29, 19) {real, imag} */,
  {32'hbfb8bb56, 32'h3ee15383} /* (24, 29, 18) {real, imag} */,
  {32'hbf00ce95, 32'h3ffaa248} /* (24, 29, 17) {real, imag} */,
  {32'h3f1747c6, 32'hc01254a4} /* (24, 29, 16) {real, imag} */,
  {32'hc024318f, 32'h3f1bb01f} /* (24, 29, 15) {real, imag} */,
  {32'h3dbf5c17, 32'hc02f4425} /* (24, 29, 14) {real, imag} */,
  {32'hc042e15e, 32'h40058722} /* (24, 29, 13) {real, imag} */,
  {32'h402a8bb7, 32'h3fb9e4d5} /* (24, 29, 12) {real, imag} */,
  {32'h3fef972a, 32'hbfdf9f27} /* (24, 29, 11) {real, imag} */,
  {32'h4072adae, 32'hbf8b2986} /* (24, 29, 10) {real, imag} */,
  {32'hbe1374f0, 32'hbeadd8af} /* (24, 29, 9) {real, imag} */,
  {32'hbfa6af4d, 32'h4088221b} /* (24, 29, 8) {real, imag} */,
  {32'hbf9af070, 32'hbfe3bc93} /* (24, 29, 7) {real, imag} */,
  {32'hbfba1e2b, 32'hc02f3d3b} /* (24, 29, 6) {real, imag} */,
  {32'hbf8bbac1, 32'h3f63164f} /* (24, 29, 5) {real, imag} */,
  {32'hc0887583, 32'hbfd9c269} /* (24, 29, 4) {real, imag} */,
  {32'h4095af02, 32'h3e5d8c1c} /* (24, 29, 3) {real, imag} */,
  {32'h40068ba2, 32'hc0110168} /* (24, 29, 2) {real, imag} */,
  {32'hc01df710, 32'h40bc59ec} /* (24, 29, 1) {real, imag} */,
  {32'hc0198b69, 32'h401042fc} /* (24, 29, 0) {real, imag} */,
  {32'hc0f7e71a, 32'hc05d9d64} /* (24, 28, 31) {real, imag} */,
  {32'h40ea6c66, 32'h4014fc6d} /* (24, 28, 30) {real, imag} */,
  {32'h3f886eda, 32'hc000c538} /* (24, 28, 29) {real, imag} */,
  {32'hc00dec04, 32'h40d61f2f} /* (24, 28, 28) {real, imag} */,
  {32'h3fc9b4ff, 32'hbdf3a32a} /* (24, 28, 27) {real, imag} */,
  {32'h40055f4c, 32'h406b31fe} /* (24, 28, 26) {real, imag} */,
  {32'hc0be84d6, 32'hbf4ea635} /* (24, 28, 25) {real, imag} */,
  {32'h405460ce, 32'h40a9d0f5} /* (24, 28, 24) {real, imag} */,
  {32'hc031b069, 32'hbfe7d719} /* (24, 28, 23) {real, imag} */,
  {32'h3e99094b, 32'h4047c216} /* (24, 28, 22) {real, imag} */,
  {32'hbf84e837, 32'h401ca4f9} /* (24, 28, 21) {real, imag} */,
  {32'h3e646fca, 32'hc0100856} /* (24, 28, 20) {real, imag} */,
  {32'hc056d4e4, 32'hc0303edd} /* (24, 28, 19) {real, imag} */,
  {32'hbfc1ce73, 32'hbfb4da9a} /* (24, 28, 18) {real, imag} */,
  {32'hbe126820, 32'h3f86c7a1} /* (24, 28, 17) {real, imag} */,
  {32'h400174bc, 32'h3f405fd3} /* (24, 28, 16) {real, imag} */,
  {32'hbf55d955, 32'hbfde7175} /* (24, 28, 15) {real, imag} */,
  {32'h40391619, 32'hbfbfa436} /* (24, 28, 14) {real, imag} */,
  {32'h3fba181c, 32'h3e398389} /* (24, 28, 13) {real, imag} */,
  {32'hbf6ed86f, 32'hbdd7df8f} /* (24, 28, 12) {real, imag} */,
  {32'h401d7724, 32'hbf4c83c5} /* (24, 28, 11) {real, imag} */,
  {32'h3ecd79bc, 32'h3ec7357f} /* (24, 28, 10) {real, imag} */,
  {32'hbfdf6616, 32'h3f6fcaa0} /* (24, 28, 9) {real, imag} */,
  {32'h3ff4c602, 32'h3e58d007} /* (24, 28, 8) {real, imag} */,
  {32'h405248c1, 32'h3faeaab9} /* (24, 28, 7) {real, imag} */,
  {32'hbfd18b62, 32'h404100e9} /* (24, 28, 6) {real, imag} */,
  {32'h3f40ff95, 32'h3dcf327b} /* (24, 28, 5) {real, imag} */,
  {32'hbf35cf2f, 32'hbf8a6164} /* (24, 28, 4) {real, imag} */,
  {32'h401048ff, 32'h3fe150fd} /* (24, 28, 3) {real, imag} */,
  {32'h40e66195, 32'h3f059971} /* (24, 28, 2) {real, imag} */,
  {32'hc0599ce1, 32'h40542d74} /* (24, 28, 1) {real, imag} */,
  {32'hbf5022cf, 32'h3f2af00b} /* (24, 28, 0) {real, imag} */,
  {32'h40390c61, 32'hbfbdb0b6} /* (24, 27, 31) {real, imag} */,
  {32'hc0251a4d, 32'h401855a3} /* (24, 27, 30) {real, imag} */,
  {32'h4003d02c, 32'h4001146e} /* (24, 27, 29) {real, imag} */,
  {32'h40180b63, 32'hc096e41a} /* (24, 27, 28) {real, imag} */,
  {32'h40688344, 32'hc03170d8} /* (24, 27, 27) {real, imag} */,
  {32'hbfe5e3a3, 32'hbc773557} /* (24, 27, 26) {real, imag} */,
  {32'h3ea9ec2d, 32'hbfc13ea6} /* (24, 27, 25) {real, imag} */,
  {32'hbf99c8a3, 32'hbed6a4c7} /* (24, 27, 24) {real, imag} */,
  {32'hbfd8b6d2, 32'hbe0716dc} /* (24, 27, 23) {real, imag} */,
  {32'h3f199ad3, 32'h3f8689f5} /* (24, 27, 22) {real, imag} */,
  {32'h4064c769, 32'h4003069f} /* (24, 27, 21) {real, imag} */,
  {32'h3f8b74d5, 32'hbecc6a14} /* (24, 27, 20) {real, imag} */,
  {32'hbfd570e3, 32'h40363173} /* (24, 27, 19) {real, imag} */,
  {32'hbf637af7, 32'h403d72bb} /* (24, 27, 18) {real, imag} */,
  {32'h402605b5, 32'hbf87fd7b} /* (24, 27, 17) {real, imag} */,
  {32'h3f0d7b46, 32'hbf670f26} /* (24, 27, 16) {real, imag} */,
  {32'hbf21cec5, 32'h3e019198} /* (24, 27, 15) {real, imag} */,
  {32'h3f6ad938, 32'hbf7afd89} /* (24, 27, 14) {real, imag} */,
  {32'hbf780e73, 32'hbfb3a2ec} /* (24, 27, 13) {real, imag} */,
  {32'hbf6c2a76, 32'hbf5b8c7c} /* (24, 27, 12) {real, imag} */,
  {32'hbfb0e1b9, 32'h3e9ae9c1} /* (24, 27, 11) {real, imag} */,
  {32'hbe9b35c2, 32'hc055a960} /* (24, 27, 10) {real, imag} */,
  {32'h3f8e29e2, 32'h3da6cb58} /* (24, 27, 9) {real, imag} */,
  {32'h3fc575cb, 32'h3f85edd3} /* (24, 27, 8) {real, imag} */,
  {32'h3ffcb912, 32'h3fd13dd8} /* (24, 27, 7) {real, imag} */,
  {32'h3fc40b46, 32'h3e1500c6} /* (24, 27, 6) {real, imag} */,
  {32'h3fb62130, 32'hc00ffbf7} /* (24, 27, 5) {real, imag} */,
  {32'h4060b3c4, 32'hbe5f37c8} /* (24, 27, 4) {real, imag} */,
  {32'h3f611447, 32'h3f083ae3} /* (24, 27, 3) {real, imag} */,
  {32'hc05de3e6, 32'hc01d8cb4} /* (24, 27, 2) {real, imag} */,
  {32'h4089e028, 32'h40d60d12} /* (24, 27, 1) {real, imag} */,
  {32'h40c93c1a, 32'h403a652f} /* (24, 27, 0) {real, imag} */,
  {32'h4028e993, 32'hbf19d209} /* (24, 26, 31) {real, imag} */,
  {32'h3f5a0750, 32'h3f28abfc} /* (24, 26, 30) {real, imag} */,
  {32'hbfe48670, 32'hc051c608} /* (24, 26, 29) {real, imag} */,
  {32'h3e030747, 32'h3f06cc79} /* (24, 26, 28) {real, imag} */,
  {32'h3fd066b7, 32'h3fbec40c} /* (24, 26, 27) {real, imag} */,
  {32'hc0031099, 32'h3f636265} /* (24, 26, 26) {real, imag} */,
  {32'hc028b9c0, 32'hbfec431f} /* (24, 26, 25) {real, imag} */,
  {32'hc01e96ba, 32'h4080184e} /* (24, 26, 24) {real, imag} */,
  {32'h3eb924fc, 32'h4090728a} /* (24, 26, 23) {real, imag} */,
  {32'hbfda4d8a, 32'hbf2091ad} /* (24, 26, 22) {real, imag} */,
  {32'h3eaf4fcc, 32'hbff74801} /* (24, 26, 21) {real, imag} */,
  {32'h400c38e3, 32'h3fc23ddb} /* (24, 26, 20) {real, imag} */,
  {32'hbf39bef4, 32'h3fe26b52} /* (24, 26, 19) {real, imag} */,
  {32'h3e8a8adf, 32'hbe207cc2} /* (24, 26, 18) {real, imag} */,
  {32'h3f1ceaa0, 32'h3e59d933} /* (24, 26, 17) {real, imag} */,
  {32'hbf8bf209, 32'h3f600c2c} /* (24, 26, 16) {real, imag} */,
  {32'h40838c00, 32'hbfcd5331} /* (24, 26, 15) {real, imag} */,
  {32'h3ea1071b, 32'h401320f9} /* (24, 26, 14) {real, imag} */,
  {32'hbf8b275e, 32'h3f848dc0} /* (24, 26, 13) {real, imag} */,
  {32'h3ecc39ae, 32'h401f4638} /* (24, 26, 12) {real, imag} */,
  {32'hbf3a63c9, 32'h3e3e7e0d} /* (24, 26, 11) {real, imag} */,
  {32'h3f85f1fd, 32'hbf8f79a5} /* (24, 26, 10) {real, imag} */,
  {32'h3f7e48e3, 32'hbf8fa671} /* (24, 26, 9) {real, imag} */,
  {32'h3ef4b6bf, 32'h3fa79f68} /* (24, 26, 8) {real, imag} */,
  {32'h407da905, 32'hbfb59158} /* (24, 26, 7) {real, imag} */,
  {32'hbf9dc94b, 32'h40418e2f} /* (24, 26, 6) {real, imag} */,
  {32'hc00a90d8, 32'hc00602fb} /* (24, 26, 5) {real, imag} */,
  {32'hc00fcf0a, 32'hbfeb0660} /* (24, 26, 4) {real, imag} */,
  {32'h406bef34, 32'h40560aee} /* (24, 26, 3) {real, imag} */,
  {32'h4046c2f7, 32'hc01fb7c4} /* (24, 26, 2) {real, imag} */,
  {32'h409baee7, 32'h3fb92203} /* (24, 26, 1) {real, imag} */,
  {32'hbedd3871, 32'h40342f26} /* (24, 26, 0) {real, imag} */,
  {32'h3fd9924a, 32'h40c3f90b} /* (24, 25, 31) {real, imag} */,
  {32'h3c9da54a, 32'h3e5f8a8e} /* (24, 25, 30) {real, imag} */,
  {32'hc06b862a, 32'hc0494699} /* (24, 25, 29) {real, imag} */,
  {32'hbf7e4d55, 32'hc0175b97} /* (24, 25, 28) {real, imag} */,
  {32'h40305f2a, 32'hc01bd4bc} /* (24, 25, 27) {real, imag} */,
  {32'hc012f825, 32'hbf1a6dd4} /* (24, 25, 26) {real, imag} */,
  {32'hbfe24565, 32'hc0002fdb} /* (24, 25, 25) {real, imag} */,
  {32'h3ee9c432, 32'hc098dc93} /* (24, 25, 24) {real, imag} */,
  {32'h3f94e675, 32'h3fece42f} /* (24, 25, 23) {real, imag} */,
  {32'h3e24b456, 32'hbede9741} /* (24, 25, 22) {real, imag} */,
  {32'h406a044b, 32'h3f0ab662} /* (24, 25, 21) {real, imag} */,
  {32'hbef44718, 32'hbf0d3e21} /* (24, 25, 20) {real, imag} */,
  {32'hc028cf20, 32'h3fc2ca47} /* (24, 25, 19) {real, imag} */,
  {32'h4026762f, 32'hbfd0a03e} /* (24, 25, 18) {real, imag} */,
  {32'hbe7c1b7a, 32'h3f0a7546} /* (24, 25, 17) {real, imag} */,
  {32'h3ef3e08c, 32'hbee22356} /* (24, 25, 16) {real, imag} */,
  {32'h3f5c9f8a, 32'hbfe8ea08} /* (24, 25, 15) {real, imag} */,
  {32'h3e3bb36c, 32'h4011e208} /* (24, 25, 14) {real, imag} */,
  {32'h3e767820, 32'hbc1075ba} /* (24, 25, 13) {real, imag} */,
  {32'h3f230410, 32'h3d8a31d7} /* (24, 25, 12) {real, imag} */,
  {32'hc02e0cc5, 32'hc00e3eab} /* (24, 25, 11) {real, imag} */,
  {32'h403438ba, 32'h3f4103ac} /* (24, 25, 10) {real, imag} */,
  {32'hbefe283b, 32'h3ea5941b} /* (24, 25, 9) {real, imag} */,
  {32'hbf8cfd78, 32'h3f6059fb} /* (24, 25, 8) {real, imag} */,
  {32'h3d846d97, 32'hc03ee135} /* (24, 25, 7) {real, imag} */,
  {32'h3fa70676, 32'h4008755e} /* (24, 25, 6) {real, imag} */,
  {32'hbfbd0f5e, 32'h3e3798d6} /* (24, 25, 5) {real, imag} */,
  {32'h3f7a5c7d, 32'hbf06a091} /* (24, 25, 4) {real, imag} */,
  {32'hc0353e6f, 32'h3f1ec191} /* (24, 25, 3) {real, imag} */,
  {32'hbe7c8d28, 32'h3f535da0} /* (24, 25, 2) {real, imag} */,
  {32'hc088c08e, 32'h3fe29bb3} /* (24, 25, 1) {real, imag} */,
  {32'h3fe73424, 32'hc056de71} /* (24, 25, 0) {real, imag} */,
  {32'h3f85c819, 32'hbfb5249b} /* (24, 24, 31) {real, imag} */,
  {32'hc104f28e, 32'hbe99b8d7} /* (24, 24, 30) {real, imag} */,
  {32'hbe938e34, 32'h3fd86c34} /* (24, 24, 29) {real, imag} */,
  {32'h40470fbc, 32'h40c8ecb4} /* (24, 24, 28) {real, imag} */,
  {32'h3fb7b7e7, 32'h3fbf33a7} /* (24, 24, 27) {real, imag} */,
  {32'h3ff5f6dc, 32'h3fd1af33} /* (24, 24, 26) {real, imag} */,
  {32'hc019521d, 32'hbf1dbd44} /* (24, 24, 25) {real, imag} */,
  {32'hbf95d52e, 32'h403cb7f7} /* (24, 24, 24) {real, imag} */,
  {32'h4096c2de, 32'h40413db1} /* (24, 24, 23) {real, imag} */,
  {32'h404c6632, 32'hc0488414} /* (24, 24, 22) {real, imag} */,
  {32'hc0851310, 32'h3e5401e1} /* (24, 24, 21) {real, imag} */,
  {32'h3edc8de6, 32'hbe98d82a} /* (24, 24, 20) {real, imag} */,
  {32'hbfb09404, 32'h3ef93d4f} /* (24, 24, 19) {real, imag} */,
  {32'hc054f896, 32'hc09bdf91} /* (24, 24, 18) {real, imag} */,
  {32'h4007035b, 32'h3e56f76f} /* (24, 24, 17) {real, imag} */,
  {32'h3fc1f54f, 32'h40591702} /* (24, 24, 16) {real, imag} */,
  {32'hbf74f8b0, 32'hbdf19db2} /* (24, 24, 15) {real, imag} */,
  {32'h3f6898c1, 32'hbe7ef864} /* (24, 24, 14) {real, imag} */,
  {32'hbf0f65b7, 32'h3f93cf7d} /* (24, 24, 13) {real, imag} */,
  {32'hbf91281c, 32'hbf36759f} /* (24, 24, 12) {real, imag} */,
  {32'h40152001, 32'hc01e7f87} /* (24, 24, 11) {real, imag} */,
  {32'hbeb8e6b4, 32'hc083b0d7} /* (24, 24, 10) {real, imag} */,
  {32'hbf69a182, 32'h404af914} /* (24, 24, 9) {real, imag} */,
  {32'hbff905b6, 32'h3fc3e516} /* (24, 24, 8) {real, imag} */,
  {32'h3c33ea20, 32'h40878c8a} /* (24, 24, 7) {real, imag} */,
  {32'hbf88056b, 32'h4021cc99} /* (24, 24, 6) {real, imag} */,
  {32'hbf7b0e35, 32'h3f3e0ef2} /* (24, 24, 5) {real, imag} */,
  {32'h407bfe82, 32'h40698e16} /* (24, 24, 4) {real, imag} */,
  {32'h4004d7cd, 32'h405c72f6} /* (24, 24, 3) {real, imag} */,
  {32'h3f9cdc34, 32'hbff71051} /* (24, 24, 2) {real, imag} */,
  {32'h404b198c, 32'h3f809cb8} /* (24, 24, 1) {real, imag} */,
  {32'h40188965, 32'hbf138815} /* (24, 24, 0) {real, imag} */,
  {32'hbfcc3d0d, 32'h3e43d6fd} /* (24, 23, 31) {real, imag} */,
  {32'hbea9044d, 32'hbecf1229} /* (24, 23, 30) {real, imag} */,
  {32'h4037cdea, 32'h40770a34} /* (24, 23, 29) {real, imag} */,
  {32'hbfec9c74, 32'hc02eb491} /* (24, 23, 28) {real, imag} */,
  {32'hbf4d4aa1, 32'h3f581fe6} /* (24, 23, 27) {real, imag} */,
  {32'hbfaf2bae, 32'hbf0ec0dd} /* (24, 23, 26) {real, imag} */,
  {32'hbe74859b, 32'hbe7b85e4} /* (24, 23, 25) {real, imag} */,
  {32'h3f8d6d1c, 32'h3f902b58} /* (24, 23, 24) {real, imag} */,
  {32'hc03647c2, 32'hc0035c71} /* (24, 23, 23) {real, imag} */,
  {32'h3f38e9f0, 32'hc007db34} /* (24, 23, 22) {real, imag} */,
  {32'hbef074b9, 32'h3fa96358} /* (24, 23, 21) {real, imag} */,
  {32'h405b83d4, 32'hc004e773} /* (24, 23, 20) {real, imag} */,
  {32'h406968f3, 32'h3e80bc31} /* (24, 23, 19) {real, imag} */,
  {32'h3cc57f88, 32'h3f1c45b5} /* (24, 23, 18) {real, imag} */,
  {32'h4001d217, 32'hc0120f4c} /* (24, 23, 17) {real, imag} */,
  {32'hbee85efe, 32'h3f96275f} /* (24, 23, 16) {real, imag} */,
  {32'h40203f65, 32'hbed30c46} /* (24, 23, 15) {real, imag} */,
  {32'hc01325e6, 32'h3e1101b1} /* (24, 23, 14) {real, imag} */,
  {32'h402d009f, 32'hc089d166} /* (24, 23, 13) {real, imag} */,
  {32'h3f805f73, 32'hbf221fa6} /* (24, 23, 12) {real, imag} */,
  {32'hbfd96a34, 32'h3f7906a8} /* (24, 23, 11) {real, imag} */,
  {32'h3ecbeb5f, 32'hbf00c43a} /* (24, 23, 10) {real, imag} */,
  {32'h3faf1104, 32'h402ffeb1} /* (24, 23, 9) {real, imag} */,
  {32'hbec50a7f, 32'hbfd55e15} /* (24, 23, 8) {real, imag} */,
  {32'h3f38c7fd, 32'h3e80da89} /* (24, 23, 7) {real, imag} */,
  {32'h3f54bdea, 32'hc0274056} /* (24, 23, 6) {real, imag} */,
  {32'h3f73e45c, 32'hbfbfad9a} /* (24, 23, 5) {real, imag} */,
  {32'hc03a9209, 32'h3fc5c806} /* (24, 23, 4) {real, imag} */,
  {32'h3f3c7f96, 32'h3fb0f10c} /* (24, 23, 3) {real, imag} */,
  {32'hbee6c34a, 32'h405dfc54} /* (24, 23, 2) {real, imag} */,
  {32'hc0241804, 32'h400c1be6} /* (24, 23, 1) {real, imag} */,
  {32'hc0211aa3, 32'h3fba1744} /* (24, 23, 0) {real, imag} */,
  {32'hbf7ea675, 32'hbfe17ac8} /* (24, 22, 31) {real, imag} */,
  {32'h40569bd2, 32'h3c8b304b} /* (24, 22, 30) {real, imag} */,
  {32'hc02ddce5, 32'h3f0452bc} /* (24, 22, 29) {real, imag} */,
  {32'hbebd856d, 32'h3e516c04} /* (24, 22, 28) {real, imag} */,
  {32'h3f3c6ea9, 32'hbe665376} /* (24, 22, 27) {real, imag} */,
  {32'hbfd478cf, 32'h400a4e20} /* (24, 22, 26) {real, imag} */,
  {32'hbd6ec555, 32'h4001ad57} /* (24, 22, 25) {real, imag} */,
  {32'hbff504e1, 32'hbf4c9af9} /* (24, 22, 24) {real, imag} */,
  {32'h3fb82a01, 32'hbe6d2a88} /* (24, 22, 23) {real, imag} */,
  {32'h40471e73, 32'h3fbe68c4} /* (24, 22, 22) {real, imag} */,
  {32'h3f9d53f7, 32'h3e5eecc6} /* (24, 22, 21) {real, imag} */,
  {32'hbfcb4f09, 32'hbe2b2019} /* (24, 22, 20) {real, imag} */,
  {32'h3e18f290, 32'hc030f6c3} /* (24, 22, 19) {real, imag} */,
  {32'hbfee1522, 32'hbeb07a62} /* (24, 22, 18) {real, imag} */,
  {32'h3fdb4698, 32'h3f83f81b} /* (24, 22, 17) {real, imag} */,
  {32'hbe88c5f6, 32'h3eb8f584} /* (24, 22, 16) {real, imag} */,
  {32'h3f5c84ac, 32'h3f8c31b5} /* (24, 22, 15) {real, imag} */,
  {32'h3e18f5e8, 32'h3f621759} /* (24, 22, 14) {real, imag} */,
  {32'h40112eec, 32'hc0080bdf} /* (24, 22, 13) {real, imag} */,
  {32'hbf11c69f, 32'hbedc50a1} /* (24, 22, 12) {real, imag} */,
  {32'h3feb0f79, 32'h3eb83c2c} /* (24, 22, 11) {real, imag} */,
  {32'h3eb1e8a1, 32'h3efa7d30} /* (24, 22, 10) {real, imag} */,
  {32'hc00eb0d6, 32'h3fa1e476} /* (24, 22, 9) {real, imag} */,
  {32'h3f81e806, 32'h3ecb87f8} /* (24, 22, 8) {real, imag} */,
  {32'hbd43f480, 32'h3e6ddeac} /* (24, 22, 7) {real, imag} */,
  {32'hbe7e8173, 32'hbd845900} /* (24, 22, 6) {real, imag} */,
  {32'h3e6fa912, 32'h3fbe09a6} /* (24, 22, 5) {real, imag} */,
  {32'hbf9a1a75, 32'hbfa06d93} /* (24, 22, 4) {real, imag} */,
  {32'h3eb63b1c, 32'hbe976334} /* (24, 22, 3) {real, imag} */,
  {32'h3e8d880e, 32'hc0009b07} /* (24, 22, 2) {real, imag} */,
  {32'hc03c600d, 32'h4060dbfe} /* (24, 22, 1) {real, imag} */,
  {32'hbfff24c2, 32'hbda9eb87} /* (24, 22, 0) {real, imag} */,
  {32'h3f5cb411, 32'hbf83c0ce} /* (24, 21, 31) {real, imag} */,
  {32'hc00b5e67, 32'h4058a06a} /* (24, 21, 30) {real, imag} */,
  {32'h3fa3b437, 32'h4017a7df} /* (24, 21, 29) {real, imag} */,
  {32'h3ff379f0, 32'h3fd9a15f} /* (24, 21, 28) {real, imag} */,
  {32'hbff1328a, 32'hbf31ad7c} /* (24, 21, 27) {real, imag} */,
  {32'h40087ea4, 32'h3f1e08d0} /* (24, 21, 26) {real, imag} */,
  {32'hc035fe4b, 32'hbfc103f5} /* (24, 21, 25) {real, imag} */,
  {32'hc00def69, 32'h40076489} /* (24, 21, 24) {real, imag} */,
  {32'h3fe8b6ae, 32'h3fbf5b15} /* (24, 21, 23) {real, imag} */,
  {32'hc075588e, 32'hc02c501a} /* (24, 21, 22) {real, imag} */,
  {32'hbf47cc31, 32'hc03cfb26} /* (24, 21, 21) {real, imag} */,
  {32'hc003b553, 32'h3deabc32} /* (24, 21, 20) {real, imag} */,
  {32'hc042e537, 32'h3fdb83ad} /* (24, 21, 19) {real, imag} */,
  {32'h3f4ab007, 32'h405dfcd7} /* (24, 21, 18) {real, imag} */,
  {32'h3e1f8326, 32'hbfd2f1d3} /* (24, 21, 17) {real, imag} */,
  {32'h3ee55716, 32'hbf1f29c2} /* (24, 21, 16) {real, imag} */,
  {32'hbfdc94a0, 32'hbe8e9272} /* (24, 21, 15) {real, imag} */,
  {32'hbf327cd9, 32'hbf6783a1} /* (24, 21, 14) {real, imag} */,
  {32'h3f8000ee, 32'h3f5c03b0} /* (24, 21, 13) {real, imag} */,
  {32'h3ee16d17, 32'hc016954b} /* (24, 21, 12) {real, imag} */,
  {32'hbea0a4c1, 32'hbfc08e29} /* (24, 21, 11) {real, imag} */,
  {32'h3fe7b713, 32'hbf88c911} /* (24, 21, 10) {real, imag} */,
  {32'hbec8b6fc, 32'h3fb18ca4} /* (24, 21, 9) {real, imag} */,
  {32'h3e3dc0c0, 32'hc000d850} /* (24, 21, 8) {real, imag} */,
  {32'hbfcf4e0f, 32'h3fb12de0} /* (24, 21, 7) {real, imag} */,
  {32'h40037cce, 32'hbf624ae9} /* (24, 21, 6) {real, imag} */,
  {32'hbf4f0823, 32'h4042a404} /* (24, 21, 5) {real, imag} */,
  {32'h3f4fb4c9, 32'h404daed6} /* (24, 21, 4) {real, imag} */,
  {32'h3c9724ff, 32'hbf784581} /* (24, 21, 3) {real, imag} */,
  {32'h3f62f4be, 32'hbf3da8cd} /* (24, 21, 2) {real, imag} */,
  {32'h4080be94, 32'hbfea3cdb} /* (24, 21, 1) {real, imag} */,
  {32'h3fd70bc2, 32'hc042add0} /* (24, 21, 0) {real, imag} */,
  {32'hbf8279a2, 32'h3eaf209f} /* (24, 20, 31) {real, imag} */,
  {32'hbf2f7179, 32'h3e8cb1bb} /* (24, 20, 30) {real, imag} */,
  {32'h3d1b83ec, 32'h3fe1db5f} /* (24, 20, 29) {real, imag} */,
  {32'hbf8a61ca, 32'hbfd2c996} /* (24, 20, 28) {real, imag} */,
  {32'h3fd9e973, 32'h401a2e21} /* (24, 20, 27) {real, imag} */,
  {32'h3eec1e8d, 32'h3fa1b2f6} /* (24, 20, 26) {real, imag} */,
  {32'h4043421f, 32'hc0651ca0} /* (24, 20, 25) {real, imag} */,
  {32'h3eec266d, 32'hc0a44370} /* (24, 20, 24) {real, imag} */,
  {32'h3f2cb7b4, 32'h3f7a85ea} /* (24, 20, 23) {real, imag} */,
  {32'hc0560cc0, 32'hbe1c9cc4} /* (24, 20, 22) {real, imag} */,
  {32'hbea596c7, 32'hbfd2e50b} /* (24, 20, 21) {real, imag} */,
  {32'h3f258ca5, 32'hbe09da80} /* (24, 20, 20) {real, imag} */,
  {32'hbf933751, 32'h400c1ce2} /* (24, 20, 19) {real, imag} */,
  {32'hbfd4c1f0, 32'h3ed90c38} /* (24, 20, 18) {real, imag} */,
  {32'h3dc82db8, 32'h40a2e797} /* (24, 20, 17) {real, imag} */,
  {32'h3fb0a15f, 32'hbfe711ae} /* (24, 20, 16) {real, imag} */,
  {32'h3fca8a87, 32'hbf16cbd8} /* (24, 20, 15) {real, imag} */,
  {32'hc040078a, 32'h3fdb666e} /* (24, 20, 14) {real, imag} */,
  {32'h4033c770, 32'h3f1ebb7c} /* (24, 20, 13) {real, imag} */,
  {32'hbf10a5fd, 32'h3fbd4745} /* (24, 20, 12) {real, imag} */,
  {32'hbff84502, 32'h403bcfa5} /* (24, 20, 11) {real, imag} */,
  {32'h3fb75646, 32'h4015f6c3} /* (24, 20, 10) {real, imag} */,
  {32'hbfae74c2, 32'h3f11b9bd} /* (24, 20, 9) {real, imag} */,
  {32'h40264257, 32'h3f617911} /* (24, 20, 8) {real, imag} */,
  {32'hbcc77cc1, 32'h3f5652d2} /* (24, 20, 7) {real, imag} */,
  {32'hbffc0c83, 32'hbfb89fb5} /* (24, 20, 6) {real, imag} */,
  {32'h3ed305a9, 32'h3ff9858d} /* (24, 20, 5) {real, imag} */,
  {32'hbe2f4b26, 32'h4071953a} /* (24, 20, 4) {real, imag} */,
  {32'hc02a5087, 32'hbfb7fc9f} /* (24, 20, 3) {real, imag} */,
  {32'hbaa96760, 32'h402948ee} /* (24, 20, 2) {real, imag} */,
  {32'hbf32d11e, 32'hc009c357} /* (24, 20, 1) {real, imag} */,
  {32'hbe8838ef, 32'hbf9c0eb9} /* (24, 20, 0) {real, imag} */,
  {32'hbf598cc5, 32'hbff77817} /* (24, 19, 31) {real, imag} */,
  {32'h3dd688f5, 32'h3fb71920} /* (24, 19, 30) {real, imag} */,
  {32'hbfb44685, 32'hbf4864f6} /* (24, 19, 29) {real, imag} */,
  {32'hbe91bfb9, 32'h40380493} /* (24, 19, 28) {real, imag} */,
  {32'h3f2b4e12, 32'hc021e3ff} /* (24, 19, 27) {real, imag} */,
  {32'h3f8574d5, 32'hbffb8d32} /* (24, 19, 26) {real, imag} */,
  {32'h3eec2a32, 32'h3f7f0f4e} /* (24, 19, 25) {real, imag} */,
  {32'h40466d06, 32'h3f693eb9} /* (24, 19, 24) {real, imag} */,
  {32'h4038bf6f, 32'hbf230238} /* (24, 19, 23) {real, imag} */,
  {32'h3fb24392, 32'h3ee0f0f5} /* (24, 19, 22) {real, imag} */,
  {32'hc086dca5, 32'h40486a71} /* (24, 19, 21) {real, imag} */,
  {32'h400ca397, 32'h3dd42c51} /* (24, 19, 20) {real, imag} */,
  {32'h3e1b9b53, 32'h3e85417f} /* (24, 19, 19) {real, imag} */,
  {32'h3da240d4, 32'h3fe358a1} /* (24, 19, 18) {real, imag} */,
  {32'h3ee943b8, 32'h3fd9abad} /* (24, 19, 17) {real, imag} */,
  {32'hc006c524, 32'hbf99e4fd} /* (24, 19, 16) {real, imag} */,
  {32'h3feb3afb, 32'hbeb0a0bf} /* (24, 19, 15) {real, imag} */,
  {32'h403a55ce, 32'h3ee98418} /* (24, 19, 14) {real, imag} */,
  {32'hbf892560, 32'hc024b617} /* (24, 19, 13) {real, imag} */,
  {32'h3fa59d32, 32'h3fee73a6} /* (24, 19, 12) {real, imag} */,
  {32'h3f83e7cc, 32'h40455803} /* (24, 19, 11) {real, imag} */,
  {32'hbf1d9da0, 32'h3ff8fb68} /* (24, 19, 10) {real, imag} */,
  {32'hc02214af, 32'hc053571b} /* (24, 19, 9) {real, imag} */,
  {32'hc00e6082, 32'hbec9f320} /* (24, 19, 8) {real, imag} */,
  {32'hbf611c71, 32'hc013fe53} /* (24, 19, 7) {real, imag} */,
  {32'h3c965504, 32'hbfa771f4} /* (24, 19, 6) {real, imag} */,
  {32'h3f957b21, 32'hbdeb74c8} /* (24, 19, 5) {real, imag} */,
  {32'h3fbd4122, 32'hbf900a0f} /* (24, 19, 4) {real, imag} */,
  {32'h3fda295c, 32'hbfc9978b} /* (24, 19, 3) {real, imag} */,
  {32'hbf2b1a5c, 32'h40148d6c} /* (24, 19, 2) {real, imag} */,
  {32'hbfcf5194, 32'hc00ee17d} /* (24, 19, 1) {real, imag} */,
  {32'h3db2e204, 32'h401a6733} /* (24, 19, 0) {real, imag} */,
  {32'h3ff19c16, 32'hbfc3bf13} /* (24, 18, 31) {real, imag} */,
  {32'hbf01ca49, 32'h3de4bba7} /* (24, 18, 30) {real, imag} */,
  {32'hbe6fb784, 32'hbf12b5e2} /* (24, 18, 29) {real, imag} */,
  {32'h3fed9598, 32'hbf60e696} /* (24, 18, 28) {real, imag} */,
  {32'hbdeca958, 32'hbf270547} /* (24, 18, 27) {real, imag} */,
  {32'hbea82c46, 32'h4026e974} /* (24, 18, 26) {real, imag} */,
  {32'h3f93c49d, 32'h3fb6d59b} /* (24, 18, 25) {real, imag} */,
  {32'hbfe0f7b6, 32'h403103f4} /* (24, 18, 24) {real, imag} */,
  {32'hbf55a814, 32'h401d97c8} /* (24, 18, 23) {real, imag} */,
  {32'h3f8919e9, 32'hbf88f9dc} /* (24, 18, 22) {real, imag} */,
  {32'h3de19c10, 32'hc0286923} /* (24, 18, 21) {real, imag} */,
  {32'h3ea73a72, 32'hbf5e9090} /* (24, 18, 20) {real, imag} */,
  {32'h3f34121c, 32'h3ebde759} /* (24, 18, 19) {real, imag} */,
  {32'h3f935f9a, 32'hc00a4831} /* (24, 18, 18) {real, imag} */,
  {32'hbf93a371, 32'h3fb73181} /* (24, 18, 17) {real, imag} */,
  {32'hbf896824, 32'h401c6b14} /* (24, 18, 16) {real, imag} */,
  {32'hbfee118a, 32'hc010dc14} /* (24, 18, 15) {real, imag} */,
  {32'h3fbf7987, 32'h40583443} /* (24, 18, 14) {real, imag} */,
  {32'hbdf6ad57, 32'h3f21d080} /* (24, 18, 13) {real, imag} */,
  {32'hbfdef551, 32'hc01984e9} /* (24, 18, 12) {real, imag} */,
  {32'h3f8c9ebc, 32'hbfe32244} /* (24, 18, 11) {real, imag} */,
  {32'hc00d5af1, 32'h3fa439fb} /* (24, 18, 10) {real, imag} */,
  {32'h4000d282, 32'hbf53c2bf} /* (24, 18, 9) {real, imag} */,
  {32'h3f36e1bd, 32'hbf999b05} /* (24, 18, 8) {real, imag} */,
  {32'h3fa3442c, 32'hc020a9bf} /* (24, 18, 7) {real, imag} */,
  {32'hc0140df4, 32'hbfa32959} /* (24, 18, 6) {real, imag} */,
  {32'h4016931a, 32'h3f0704ad} /* (24, 18, 5) {real, imag} */,
  {32'hbf63122f, 32'h40672904} /* (24, 18, 4) {real, imag} */,
  {32'hbed1e355, 32'h4019ffbc} /* (24, 18, 3) {real, imag} */,
  {32'hbfbd2913, 32'hbf91895e} /* (24, 18, 2) {real, imag} */,
  {32'h3da699ab, 32'hbfb26a04} /* (24, 18, 1) {real, imag} */,
  {32'h3fa0b741, 32'hbf551362} /* (24, 18, 0) {real, imag} */,
  {32'hbe50f42d, 32'hbf10f437} /* (24, 17, 31) {real, imag} */,
  {32'h3e5b047e, 32'hbff24546} /* (24, 17, 30) {real, imag} */,
  {32'hbededf1d, 32'h3fec210f} /* (24, 17, 29) {real, imag} */,
  {32'hbf757321, 32'hbfe4c3ad} /* (24, 17, 28) {real, imag} */,
  {32'hbfab280b, 32'hbef96d96} /* (24, 17, 27) {real, imag} */,
  {32'h3f88a362, 32'hbf83623b} /* (24, 17, 26) {real, imag} */,
  {32'hbe9237ce, 32'h3e98325a} /* (24, 17, 25) {real, imag} */,
  {32'hbfa17cdd, 32'hbeb2660d} /* (24, 17, 24) {real, imag} */,
  {32'hbf0926fd, 32'h3f2fe7a2} /* (24, 17, 23) {real, imag} */,
  {32'hbe976e30, 32'h3f38e918} /* (24, 17, 22) {real, imag} */,
  {32'h3e9ff539, 32'hbe9701cf} /* (24, 17, 21) {real, imag} */,
  {32'hc025592f, 32'h403b1793} /* (24, 17, 20) {real, imag} */,
  {32'h3f0b315b, 32'hbf41bc62} /* (24, 17, 19) {real, imag} */,
  {32'hbe238a01, 32'h3f76c4a4} /* (24, 17, 18) {real, imag} */,
  {32'hbeaeb6f9, 32'hbf9b24be} /* (24, 17, 17) {real, imag} */,
  {32'hbf60caad, 32'hbea84d54} /* (24, 17, 16) {real, imag} */,
  {32'hbf8f85e9, 32'hbe901f1e} /* (24, 17, 15) {real, imag} */,
  {32'hbe9cfcac, 32'hbf186fbe} /* (24, 17, 14) {real, imag} */,
  {32'hbf3b4e9d, 32'hbe33f57e} /* (24, 17, 13) {real, imag} */,
  {32'h3edcf558, 32'hbe30d9e3} /* (24, 17, 12) {real, imag} */,
  {32'hbeb2cb8b, 32'h3f35b875} /* (24, 17, 11) {real, imag} */,
  {32'hc00ac5b9, 32'h3fbd086b} /* (24, 17, 10) {real, imag} */,
  {32'h3e4927cc, 32'h3fee40f5} /* (24, 17, 9) {real, imag} */,
  {32'h3f0f4fbb, 32'h3f82ef82} /* (24, 17, 8) {real, imag} */,
  {32'hbfb9be52, 32'h3ffb5cf6} /* (24, 17, 7) {real, imag} */,
  {32'hbd889e3c, 32'hbf83c8d8} /* (24, 17, 6) {real, imag} */,
  {32'hbfaa386f, 32'h3f6ddac7} /* (24, 17, 5) {real, imag} */,
  {32'h3f472c16, 32'hbf8701f6} /* (24, 17, 4) {real, imag} */,
  {32'h3f81c89f, 32'h3d96fcbe} /* (24, 17, 3) {real, imag} */,
  {32'h3f026bc5, 32'hc00dae17} /* (24, 17, 2) {real, imag} */,
  {32'h3d2f5f64, 32'h4007f9fe} /* (24, 17, 1) {real, imag} */,
  {32'h3f377a23, 32'h401368ce} /* (24, 17, 0) {real, imag} */,
  {32'hbf135e8e, 32'hbe879e5d} /* (24, 16, 31) {real, imag} */,
  {32'h3f590cbe, 32'h3f2da9f4} /* (24, 16, 30) {real, imag} */,
  {32'h3ffe6504, 32'hbfdaf5af} /* (24, 16, 29) {real, imag} */,
  {32'h3fb39b8a, 32'hbfe0a979} /* (24, 16, 28) {real, imag} */,
  {32'h3ff44b76, 32'hbf2bf986} /* (24, 16, 27) {real, imag} */,
  {32'hbfd80e8f, 32'hc0037466} /* (24, 16, 26) {real, imag} */,
  {32'h3f427337, 32'hbf0a2343} /* (24, 16, 25) {real, imag} */,
  {32'h4024ecaf, 32'hbf73de37} /* (24, 16, 24) {real, imag} */,
  {32'hbde897ef, 32'h3f478540} /* (24, 16, 23) {real, imag} */,
  {32'hc00b9683, 32'hbea78e3b} /* (24, 16, 22) {real, imag} */,
  {32'hbf325ef7, 32'h3e5dcca1} /* (24, 16, 21) {real, imag} */,
  {32'h3e8581ee, 32'hbf8b4698} /* (24, 16, 20) {real, imag} */,
  {32'h3f6d9bb8, 32'hbf3a79cc} /* (24, 16, 19) {real, imag} */,
  {32'hbe97d747, 32'h3ee90fd4} /* (24, 16, 18) {real, imag} */,
  {32'hbd7e0484, 32'h3f0fb677} /* (24, 16, 17) {real, imag} */,
  {32'h3fef6f04, 32'hbf1e8ccb} /* (24, 16, 16) {real, imag} */,
  {32'h3f8ccddb, 32'hbe81a58a} /* (24, 16, 15) {real, imag} */,
  {32'hc0570d8f, 32'hbf1731d6} /* (24, 16, 14) {real, imag} */,
  {32'hbe11f38b, 32'hbf92f9ef} /* (24, 16, 13) {real, imag} */,
  {32'h3ef5c081, 32'h3fee26d6} /* (24, 16, 12) {real, imag} */,
  {32'hbf49d3e4, 32'hbfe4bfa1} /* (24, 16, 11) {real, imag} */,
  {32'hbf1eb2c9, 32'hbe687bd3} /* (24, 16, 10) {real, imag} */,
  {32'hbeed07e9, 32'hbf521e43} /* (24, 16, 9) {real, imag} */,
  {32'hbf481f85, 32'h3fc3862b} /* (24, 16, 8) {real, imag} */,
  {32'h3f907e5b, 32'hc001ef69} /* (24, 16, 7) {real, imag} */,
  {32'h3feab74a, 32'h3e1741be} /* (24, 16, 6) {real, imag} */,
  {32'hbfa8712e, 32'h3fce6892} /* (24, 16, 5) {real, imag} */,
  {32'hbfc80ee1, 32'hbdd2eb79} /* (24, 16, 4) {real, imag} */,
  {32'hbfd57071, 32'hbf6a4c3a} /* (24, 16, 3) {real, imag} */,
  {32'hbf90574e, 32'h3f432cb1} /* (24, 16, 2) {real, imag} */,
  {32'hc02c2d4d, 32'h3efcfc6c} /* (24, 16, 1) {real, imag} */,
  {32'hbef8eea7, 32'h40419af0} /* (24, 16, 0) {real, imag} */,
  {32'h4023c02f, 32'hbe70a683} /* (24, 15, 31) {real, imag} */,
  {32'hbf529a57, 32'h3e3f18e5} /* (24, 15, 30) {real, imag} */,
  {32'hc01a4a70, 32'h3f8346cc} /* (24, 15, 29) {real, imag} */,
  {32'hbf063c42, 32'hc00c34ca} /* (24, 15, 28) {real, imag} */,
  {32'h3ffee69b, 32'h3f5e1a92} /* (24, 15, 27) {real, imag} */,
  {32'h3f28b4a5, 32'hbf9585e3} /* (24, 15, 26) {real, imag} */,
  {32'h3feb77e2, 32'h3edfdc00} /* (24, 15, 25) {real, imag} */,
  {32'hbf78c41a, 32'h401c9a65} /* (24, 15, 24) {real, imag} */,
  {32'h3d8f889c, 32'h3d4991ca} /* (24, 15, 23) {real, imag} */,
  {32'h3f8a7921, 32'hc023fd86} /* (24, 15, 22) {real, imag} */,
  {32'hbfe7d3ac, 32'hbf917420} /* (24, 15, 21) {real, imag} */,
  {32'h3f647ed1, 32'h3f86fb99} /* (24, 15, 20) {real, imag} */,
  {32'h3faca6e5, 32'h3f30e0be} /* (24, 15, 19) {real, imag} */,
  {32'h3d471995, 32'hbd8ac1e0} /* (24, 15, 18) {real, imag} */,
  {32'hbcf0d3c7, 32'h40173e85} /* (24, 15, 17) {real, imag} */,
  {32'hbf0175fb, 32'h3f326f2b} /* (24, 15, 16) {real, imag} */,
  {32'h3c8beecf, 32'h3eda28b1} /* (24, 15, 15) {real, imag} */,
  {32'h3f5c431d, 32'hbf600ad3} /* (24, 15, 14) {real, imag} */,
  {32'h3eb9f539, 32'h3ff75057} /* (24, 15, 13) {real, imag} */,
  {32'hc02ce79d, 32'h3f2580c6} /* (24, 15, 12) {real, imag} */,
  {32'hbe38f35c, 32'hbf9574b5} /* (24, 15, 11) {real, imag} */,
  {32'h3f534955, 32'hc007747d} /* (24, 15, 10) {real, imag} */,
  {32'hbf1a2376, 32'hc05b1945} /* (24, 15, 9) {real, imag} */,
  {32'h3e9c70f9, 32'hc0445380} /* (24, 15, 8) {real, imag} */,
  {32'hbeae338f, 32'h3f8332cd} /* (24, 15, 7) {real, imag} */,
  {32'hbfacadb5, 32'hc04d72dd} /* (24, 15, 6) {real, imag} */,
  {32'h3ec88569, 32'hc02c9471} /* (24, 15, 5) {real, imag} */,
  {32'h3def66cb, 32'hbe2e1468} /* (24, 15, 4) {real, imag} */,
  {32'h3ed68f38, 32'h3f0635e6} /* (24, 15, 3) {real, imag} */,
  {32'hbeadfdf7, 32'h3ee20324} /* (24, 15, 2) {real, imag} */,
  {32'hbf6f6293, 32'h3f312106} /* (24, 15, 1) {real, imag} */,
  {32'hbe5e263f, 32'hbf16b252} /* (24, 15, 0) {real, imag} */,
  {32'hbf5463b9, 32'h4018ed72} /* (24, 14, 31) {real, imag} */,
  {32'h3f08f130, 32'h3e6b9745} /* (24, 14, 30) {real, imag} */,
  {32'hbf88a7e1, 32'h3ed91430} /* (24, 14, 29) {real, imag} */,
  {32'h401b619b, 32'hbf25bdbb} /* (24, 14, 28) {real, imag} */,
  {32'hbf780b09, 32'h3f5115f6} /* (24, 14, 27) {real, imag} */,
  {32'hc05124dd, 32'h3dc4d747} /* (24, 14, 26) {real, imag} */,
  {32'h3f47bdf4, 32'hbfd0de85} /* (24, 14, 25) {real, imag} */,
  {32'h40345720, 32'hbedaabe2} /* (24, 14, 24) {real, imag} */,
  {32'h408d8f22, 32'hbf079c3a} /* (24, 14, 23) {real, imag} */,
  {32'hbd10f733, 32'h3d7c138c} /* (24, 14, 22) {real, imag} */,
  {32'hbfa0d742, 32'h4050c68b} /* (24, 14, 21) {real, imag} */,
  {32'h3fbb869f, 32'hbfb3c908} /* (24, 14, 20) {real, imag} */,
  {32'hbf22f030, 32'hbf6033b6} /* (24, 14, 19) {real, imag} */,
  {32'hbefe3a91, 32'h400e0952} /* (24, 14, 18) {real, imag} */,
  {32'hbfc83d62, 32'hbf5364c2} /* (24, 14, 17) {real, imag} */,
  {32'h3fe51e1c, 32'h3f868985} /* (24, 14, 16) {real, imag} */,
  {32'h3e480091, 32'hbe2f722e} /* (24, 14, 15) {real, imag} */,
  {32'h3f0b2336, 32'h3d7afafe} /* (24, 14, 14) {real, imag} */,
  {32'hbe650d08, 32'h3f94f8b2} /* (24, 14, 13) {real, imag} */,
  {32'h40211068, 32'h40623e3f} /* (24, 14, 12) {real, imag} */,
  {32'h3f952608, 32'h4022c02a} /* (24, 14, 11) {real, imag} */,
  {32'hbfe828e3, 32'hbfa9efa3} /* (24, 14, 10) {real, imag} */,
  {32'h3fd72362, 32'h403deebd} /* (24, 14, 9) {real, imag} */,
  {32'h3fe262fa, 32'h3ca09f9c} /* (24, 14, 8) {real, imag} */,
  {32'h3f9eae69, 32'hc02ad165} /* (24, 14, 7) {real, imag} */,
  {32'hbfbc7eed, 32'h3e47e577} /* (24, 14, 6) {real, imag} */,
  {32'hbf20000d, 32'h3f452e64} /* (24, 14, 5) {real, imag} */,
  {32'h3e66eb59, 32'hbf901c7b} /* (24, 14, 4) {real, imag} */,
  {32'hbf227761, 32'hc06692f3} /* (24, 14, 3) {real, imag} */,
  {32'h3f5ab9e2, 32'hbfbf31e9} /* (24, 14, 2) {real, imag} */,
  {32'hbf89e306, 32'hbf187d8e} /* (24, 14, 1) {real, imag} */,
  {32'hc0103ba8, 32'h3f0a4c4a} /* (24, 14, 0) {real, imag} */,
  {32'hbfa96b44, 32'h401277f6} /* (24, 13, 31) {real, imag} */,
  {32'h3fd08426, 32'h3ffb5ae6} /* (24, 13, 30) {real, imag} */,
  {32'h3ec8715b, 32'h3f6e1f72} /* (24, 13, 29) {real, imag} */,
  {32'h3eb65c48, 32'hbfde7a5f} /* (24, 13, 28) {real, imag} */,
  {32'h403a221c, 32'h3ed2c3a1} /* (24, 13, 27) {real, imag} */,
  {32'h3f897517, 32'h403a39bb} /* (24, 13, 26) {real, imag} */,
  {32'hbe2b1aed, 32'hbfc4a587} /* (24, 13, 25) {real, imag} */,
  {32'hbf6ed8cd, 32'h402ada54} /* (24, 13, 24) {real, imag} */,
  {32'hbf41fccd, 32'hbf430f7e} /* (24, 13, 23) {real, imag} */,
  {32'hbff6e22a, 32'hbf3696b6} /* (24, 13, 22) {real, imag} */,
  {32'hc001f16e, 32'h3e455383} /* (24, 13, 21) {real, imag} */,
  {32'hc0433a64, 32'h3eae040d} /* (24, 13, 20) {real, imag} */,
  {32'h4080f25c, 32'hbfc59d19} /* (24, 13, 19) {real, imag} */,
  {32'hbfab34a0, 32'h3fe29321} /* (24, 13, 18) {real, imag} */,
  {32'h3cca1103, 32'hbf408a04} /* (24, 13, 17) {real, imag} */,
  {32'h3f37fa64, 32'hbf58ec4c} /* (24, 13, 16) {real, imag} */,
  {32'hbd32a24b, 32'hbfc2716a} /* (24, 13, 15) {real, imag} */,
  {32'hbf9a700d, 32'hbf778e12} /* (24, 13, 14) {real, imag} */,
  {32'h3f82b0b5, 32'h403d6369} /* (24, 13, 13) {real, imag} */,
  {32'h404d6c90, 32'hc06ad6d0} /* (24, 13, 12) {real, imag} */,
  {32'h4089be61, 32'hbebdccfb} /* (24, 13, 11) {real, imag} */,
  {32'h3e87697f, 32'hbf820af6} /* (24, 13, 10) {real, imag} */,
  {32'h3ed3e0db, 32'h3f84d3da} /* (24, 13, 9) {real, imag} */,
  {32'h40250c4b, 32'h3f0757e6} /* (24, 13, 8) {real, imag} */,
  {32'h3ff0d3c9, 32'hbfd6337c} /* (24, 13, 7) {real, imag} */,
  {32'hbff1788c, 32'hbebe577c} /* (24, 13, 6) {real, imag} */,
  {32'hbeb0e229, 32'hbe9b98c2} /* (24, 13, 5) {real, imag} */,
  {32'h40050c77, 32'hbf70cb85} /* (24, 13, 4) {real, imag} */,
  {32'h3f4cb597, 32'h3fb9b6fd} /* (24, 13, 3) {real, imag} */,
  {32'h3fa609fe, 32'hbc64e742} /* (24, 13, 2) {real, imag} */,
  {32'hbfba2814, 32'hc0435130} /* (24, 13, 1) {real, imag} */,
  {32'h3ff45703, 32'h3f2e1fe3} /* (24, 13, 0) {real, imag} */,
  {32'h3d33cf7c, 32'h3e419997} /* (24, 12, 31) {real, imag} */,
  {32'hbfad98d1, 32'hbf2866dc} /* (24, 12, 30) {real, imag} */,
  {32'hbfb52bce, 32'hc01b8ac4} /* (24, 12, 29) {real, imag} */,
  {32'hbfac1d89, 32'h402c4c16} /* (24, 12, 28) {real, imag} */,
  {32'hbfbd3e19, 32'h3ffa5eaa} /* (24, 12, 27) {real, imag} */,
  {32'hbf99724c, 32'hc03071b7} /* (24, 12, 26) {real, imag} */,
  {32'h3f739fdd, 32'h3f9f7a04} /* (24, 12, 25) {real, imag} */,
  {32'h3f93fc41, 32'h4067f84d} /* (24, 12, 24) {real, imag} */,
  {32'hbd50bb57, 32'h4003373d} /* (24, 12, 23) {real, imag} */,
  {32'hbf58bffe, 32'h3f374fbb} /* (24, 12, 22) {real, imag} */,
  {32'hbffd7ebe, 32'h401810e2} /* (24, 12, 21) {real, imag} */,
  {32'h3f89b713, 32'h3e5ddbe9} /* (24, 12, 20) {real, imag} */,
  {32'h3f0e1eb9, 32'h3fda5d67} /* (24, 12, 19) {real, imag} */,
  {32'h3f222865, 32'h402e2794} /* (24, 12, 18) {real, imag} */,
  {32'h3dcb4322, 32'hc021d0a0} /* (24, 12, 17) {real, imag} */,
  {32'hc004c911, 32'hbf86495a} /* (24, 12, 16) {real, imag} */,
  {32'hbfbb4735, 32'hbfe15654} /* (24, 12, 15) {real, imag} */,
  {32'h4056f8da, 32'h3f1ad316} /* (24, 12, 14) {real, imag} */,
  {32'h3fd17f4c, 32'h3fa063a1} /* (24, 12, 13) {real, imag} */,
  {32'hbf3234c1, 32'hbf8772e6} /* (24, 12, 12) {real, imag} */,
  {32'hbed32ae7, 32'hbfc6f9a0} /* (24, 12, 11) {real, imag} */,
  {32'h40827bd9, 32'hc003ae30} /* (24, 12, 10) {real, imag} */,
  {32'h3f8702c4, 32'h3f977b6e} /* (24, 12, 9) {real, imag} */,
  {32'h3f77a21f, 32'h3f5b80e4} /* (24, 12, 8) {real, imag} */,
  {32'hbeebc58a, 32'hc05f9c22} /* (24, 12, 7) {real, imag} */,
  {32'h3fa2c609, 32'h3f2e1460} /* (24, 12, 6) {real, imag} */,
  {32'hbfc0aab0, 32'hbf7d943f} /* (24, 12, 5) {real, imag} */,
  {32'hbfd5aee4, 32'h3fbcd579} /* (24, 12, 4) {real, imag} */,
  {32'hbebb454e, 32'hbfce4a4f} /* (24, 12, 3) {real, imag} */,
  {32'h3f8d1b81, 32'h4000edd7} /* (24, 12, 2) {real, imag} */,
  {32'h3ff92039, 32'h3fb7902f} /* (24, 12, 1) {real, imag} */,
  {32'hbf95c6ad, 32'h402d3695} /* (24, 12, 0) {real, imag} */,
  {32'h3fc1c473, 32'h40050130} /* (24, 11, 31) {real, imag} */,
  {32'h3e106350, 32'hbfafc8a9} /* (24, 11, 30) {real, imag} */,
  {32'hbf932217, 32'h3e902fea} /* (24, 11, 29) {real, imag} */,
  {32'h3d8ba7d5, 32'h40115e6f} /* (24, 11, 28) {real, imag} */,
  {32'h3f4c258f, 32'h3d2984e0} /* (24, 11, 27) {real, imag} */,
  {32'hbe860f04, 32'hc03728ef} /* (24, 11, 26) {real, imag} */,
  {32'hc00b7f64, 32'h3f2b26f5} /* (24, 11, 25) {real, imag} */,
  {32'hbfb490d2, 32'h3fb9d34e} /* (24, 11, 24) {real, imag} */,
  {32'h4015742b, 32'h3eb09856} /* (24, 11, 23) {real, imag} */,
  {32'h3f8c5bed, 32'h3dacfb0e} /* (24, 11, 22) {real, imag} */,
  {32'h4015f1fd, 32'hc094cdb4} /* (24, 11, 21) {real, imag} */,
  {32'hbf9eed0e, 32'hbdf7da54} /* (24, 11, 20) {real, imag} */,
  {32'hbf8758de, 32'h3ff9920a} /* (24, 11, 19) {real, imag} */,
  {32'h3e9dc48c, 32'hbe503df9} /* (24, 11, 18) {real, imag} */,
  {32'hbeab4d8d, 32'hbeb52eec} /* (24, 11, 17) {real, imag} */,
  {32'h3fca3ce5, 32'h3e40fc02} /* (24, 11, 16) {real, imag} */,
  {32'h3f5b5e5f, 32'hbf5d0ea7} /* (24, 11, 15) {real, imag} */,
  {32'h3e766cd6, 32'hbc052ff8} /* (24, 11, 14) {real, imag} */,
  {32'h3f3c6f9f, 32'hbea7ae1b} /* (24, 11, 13) {real, imag} */,
  {32'hc05c4bcc, 32'hbfcc9d13} /* (24, 11, 12) {real, imag} */,
  {32'h3fde813e, 32'hbe1c825b} /* (24, 11, 11) {real, imag} */,
  {32'hbf841672, 32'h4007947a} /* (24, 11, 10) {real, imag} */,
  {32'h3dd42154, 32'hbf772725} /* (24, 11, 9) {real, imag} */,
  {32'hbe2bee7b, 32'h3f60bcda} /* (24, 11, 8) {real, imag} */,
  {32'h3fc32768, 32'h3fe59f91} /* (24, 11, 7) {real, imag} */,
  {32'hbeb0587a, 32'hbf0071c6} /* (24, 11, 6) {real, imag} */,
  {32'hbfb6c5e9, 32'h3f99a7bb} /* (24, 11, 5) {real, imag} */,
  {32'hc07c68f4, 32'hc0917a49} /* (24, 11, 4) {real, imag} */,
  {32'h401f9023, 32'hbe1b9154} /* (24, 11, 3) {real, imag} */,
  {32'h3fcd0a29, 32'hbf866868} /* (24, 11, 2) {real, imag} */,
  {32'hbfd6e4cb, 32'h3fbc76c3} /* (24, 11, 1) {real, imag} */,
  {32'hbefd7ec7, 32'h3e0ac460} /* (24, 11, 0) {real, imag} */,
  {32'h409af695, 32'hbf9e5eec} /* (24, 10, 31) {real, imag} */,
  {32'hbfdaa122, 32'h408898f0} /* (24, 10, 30) {real, imag} */,
  {32'hc01dd2ec, 32'h3f81ed4a} /* (24, 10, 29) {real, imag} */,
  {32'h4027b998, 32'hc0146060} /* (24, 10, 28) {real, imag} */,
  {32'hbf955c89, 32'h408ee877} /* (24, 10, 27) {real, imag} */,
  {32'hc007f512, 32'h3f6f47fb} /* (24, 10, 26) {real, imag} */,
  {32'hbff32d59, 32'hbf93188e} /* (24, 10, 25) {real, imag} */,
  {32'h40064767, 32'hbe4dea37} /* (24, 10, 24) {real, imag} */,
  {32'h3fb0aac4, 32'hbfd1ecf9} /* (24, 10, 23) {real, imag} */,
  {32'hc02f8c10, 32'h4074f6af} /* (24, 10, 22) {real, imag} */,
  {32'h400fb16e, 32'h3d60911a} /* (24, 10, 21) {real, imag} */,
  {32'h4035c8e2, 32'hbdb4806d} /* (24, 10, 20) {real, imag} */,
  {32'hbe75eed1, 32'hbe16a5f6} /* (24, 10, 19) {real, imag} */,
  {32'hbf7faed8, 32'h3f29a535} /* (24, 10, 18) {real, imag} */,
  {32'h3e0f8fa6, 32'h3fde75e3} /* (24, 10, 17) {real, imag} */,
  {32'hbfd5e880, 32'h40244b7b} /* (24, 10, 16) {real, imag} */,
  {32'h3f82dd5c, 32'h4032626f} /* (24, 10, 15) {real, imag} */,
  {32'hc002e8c3, 32'hbea7725d} /* (24, 10, 14) {real, imag} */,
  {32'h3f5a3b46, 32'hbf81bacf} /* (24, 10, 13) {real, imag} */,
  {32'h3fd4ee42, 32'hc04889c5} /* (24, 10, 12) {real, imag} */,
  {32'hbd222105, 32'h3f2fe9d7} /* (24, 10, 11) {real, imag} */,
  {32'h3fb82880, 32'hbff49547} /* (24, 10, 10) {real, imag} */,
  {32'h3f9362a8, 32'h3f54be83} /* (24, 10, 9) {real, imag} */,
  {32'hbf96b30c, 32'h3eddb02c} /* (24, 10, 8) {real, imag} */,
  {32'hbf8edb33, 32'h3fe3598c} /* (24, 10, 7) {real, imag} */,
  {32'hbf86a598, 32'h3f696ae2} /* (24, 10, 6) {real, imag} */,
  {32'hbe52f120, 32'hc0aca82a} /* (24, 10, 5) {real, imag} */,
  {32'h405c4543, 32'hbf3f6e94} /* (24, 10, 4) {real, imag} */,
  {32'h3fd1e116, 32'hbe9eb1df} /* (24, 10, 3) {real, imag} */,
  {32'h3ffd5a5f, 32'hbe4c7b92} /* (24, 10, 2) {real, imag} */,
  {32'hbf970ef7, 32'h3f5adeac} /* (24, 10, 1) {real, imag} */,
  {32'hc00b6118, 32'hc0501a1b} /* (24, 10, 0) {real, imag} */,
  {32'h3cde947c, 32'h3fc5d969} /* (24, 9, 31) {real, imag} */,
  {32'h3f8c9b05, 32'hc08583e8} /* (24, 9, 30) {real, imag} */,
  {32'hbf8fb1a9, 32'hc0034005} /* (24, 9, 29) {real, imag} */,
  {32'h3e88bc2b, 32'hc00dd446} /* (24, 9, 28) {real, imag} */,
  {32'hc009bc3f, 32'h4008f0be} /* (24, 9, 27) {real, imag} */,
  {32'hbf61fc77, 32'h3f65b504} /* (24, 9, 26) {real, imag} */,
  {32'h3f15a46d, 32'hc01faf55} /* (24, 9, 25) {real, imag} */,
  {32'hbfe6b0cb, 32'h3fe258cf} /* (24, 9, 24) {real, imag} */,
  {32'hc00f0240, 32'h3f8c0798} /* (24, 9, 23) {real, imag} */,
  {32'hbed9f97e, 32'hbf961a0c} /* (24, 9, 22) {real, imag} */,
  {32'h3f528af8, 32'hc02b985a} /* (24, 9, 21) {real, imag} */,
  {32'h402ed0b9, 32'hbff7a508} /* (24, 9, 20) {real, imag} */,
  {32'hc0167e9c, 32'hbfa08064} /* (24, 9, 19) {real, imag} */,
  {32'hc0303eb8, 32'h40d50226} /* (24, 9, 18) {real, imag} */,
  {32'hbea4cb1e, 32'hc0698207} /* (24, 9, 17) {real, imag} */,
  {32'hbfc8d6dd, 32'hbe990e8f} /* (24, 9, 16) {real, imag} */,
  {32'hbe1a4712, 32'hbfae2abf} /* (24, 9, 15) {real, imag} */,
  {32'h40264227, 32'hbf12b357} /* (24, 9, 14) {real, imag} */,
  {32'hc0bd2bc7, 32'hbfafbfb6} /* (24, 9, 13) {real, imag} */,
  {32'h3f5d0d42, 32'hc01a702a} /* (24, 9, 12) {real, imag} */,
  {32'h3ef46629, 32'hc0585d9b} /* (24, 9, 11) {real, imag} */,
  {32'hbf8a6c01, 32'hbfa31f54} /* (24, 9, 10) {real, imag} */,
  {32'h3ef6a47b, 32'h4006a36e} /* (24, 9, 9) {real, imag} */,
  {32'hbf1421fe, 32'h3f09bdf4} /* (24, 9, 8) {real, imag} */,
  {32'h3febd5ce, 32'h3faac166} /* (24, 9, 7) {real, imag} */,
  {32'h3f54a110, 32'h3f23aa15} /* (24, 9, 6) {real, imag} */,
  {32'h3e4e190b, 32'h3f236e39} /* (24, 9, 5) {real, imag} */,
  {32'h40012b8e, 32'hbe4c1eeb} /* (24, 9, 4) {real, imag} */,
  {32'h3f0b3487, 32'hc0148b21} /* (24, 9, 3) {real, imag} */,
  {32'hbf855394, 32'h405b7306} /* (24, 9, 2) {real, imag} */,
  {32'hbf8fec25, 32'h406e37af} /* (24, 9, 1) {real, imag} */,
  {32'hbe84d13e, 32'hc0845dcb} /* (24, 9, 0) {real, imag} */,
  {32'h3db0e881, 32'h40d8e539} /* (24, 8, 31) {real, imag} */,
  {32'hc0856f3e, 32'hc0c2d127} /* (24, 8, 30) {real, imag} */,
  {32'h403d89a0, 32'h4062c656} /* (24, 8, 29) {real, imag} */,
  {32'h3ff2d67a, 32'hc0a08055} /* (24, 8, 28) {real, imag} */,
  {32'hbfd50256, 32'hbfd0bb3d} /* (24, 8, 27) {real, imag} */,
  {32'h3ff6da26, 32'hbe454a84} /* (24, 8, 26) {real, imag} */,
  {32'hc04cc6ef, 32'h3f211cda} /* (24, 8, 25) {real, imag} */,
  {32'hc09ac38c, 32'h3deec6fa} /* (24, 8, 24) {real, imag} */,
  {32'h3f50a3d8, 32'hbcb43b3b} /* (24, 8, 23) {real, imag} */,
  {32'hbfb82030, 32'h3f8297f7} /* (24, 8, 22) {real, imag} */,
  {32'hbecbe5fa, 32'h3ec6fbe8} /* (24, 8, 21) {real, imag} */,
  {32'h3fdf954e, 32'hbf601ba9} /* (24, 8, 20) {real, imag} */,
  {32'hbf897d97, 32'hbfc87b9b} /* (24, 8, 19) {real, imag} */,
  {32'h3f853d01, 32'h3ebbe18d} /* (24, 8, 18) {real, imag} */,
  {32'h3f935d0c, 32'h3e554049} /* (24, 8, 17) {real, imag} */,
  {32'hbd018bf5, 32'hbfc9bac7} /* (24, 8, 16) {real, imag} */,
  {32'hbed00231, 32'h3fd488b5} /* (24, 8, 15) {real, imag} */,
  {32'h3f896f09, 32'h3ff87b18} /* (24, 8, 14) {real, imag} */,
  {32'h400d6860, 32'h403ea852} /* (24, 8, 13) {real, imag} */,
  {32'h3f309b1a, 32'h3f8f63cf} /* (24, 8, 12) {real, imag} */,
  {32'h3f20a758, 32'h3fd77344} /* (24, 8, 11) {real, imag} */,
  {32'h3f852361, 32'hbf916a17} /* (24, 8, 10) {real, imag} */,
  {32'hbfb29a42, 32'h40403ea2} /* (24, 8, 9) {real, imag} */,
  {32'h3ff216df, 32'h3f2693ce} /* (24, 8, 8) {real, imag} */,
  {32'hc08d0146, 32'h3e9cb98a} /* (24, 8, 7) {real, imag} */,
  {32'h3e8bc5c5, 32'hc0006fe4} /* (24, 8, 6) {real, imag} */,
  {32'h3e70b571, 32'hc064645d} /* (24, 8, 5) {real, imag} */,
  {32'h3ff6a202, 32'hbf4cfafe} /* (24, 8, 4) {real, imag} */,
  {32'hc07f9759, 32'h3fd5ea30} /* (24, 8, 3) {real, imag} */,
  {32'hbec2af62, 32'hc038e26c} /* (24, 8, 2) {real, imag} */,
  {32'h4022beb3, 32'h40c9f02f} /* (24, 8, 1) {real, imag} */,
  {32'h402dc63a, 32'h3f963580} /* (24, 8, 0) {real, imag} */,
  {32'hbfe83aac, 32'h3f593256} /* (24, 7, 31) {real, imag} */,
  {32'h3fecccdb, 32'h40907925} /* (24, 7, 30) {real, imag} */,
  {32'h401687b1, 32'hbfb48a0f} /* (24, 7, 29) {real, imag} */,
  {32'hc00eb141, 32'hc03628da} /* (24, 7, 28) {real, imag} */,
  {32'hbeedda40, 32'hc06f5cbc} /* (24, 7, 27) {real, imag} */,
  {32'h3f6a943f, 32'hc0712c61} /* (24, 7, 26) {real, imag} */,
  {32'h403c31fe, 32'h404634a8} /* (24, 7, 25) {real, imag} */,
  {32'h40622b4c, 32'h3fae6536} /* (24, 7, 24) {real, imag} */,
  {32'h402ec423, 32'hbfa59977} /* (24, 7, 23) {real, imag} */,
  {32'hbf304d03, 32'hc055df68} /* (24, 7, 22) {real, imag} */,
  {32'hbf97e8b1, 32'hbf3152cb} /* (24, 7, 21) {real, imag} */,
  {32'hc00f1c4c, 32'h407550b5} /* (24, 7, 20) {real, imag} */,
  {32'h3f835075, 32'hbec7acc7} /* (24, 7, 19) {real, imag} */,
  {32'hbf03d28f, 32'h3ede2452} /* (24, 7, 18) {real, imag} */,
  {32'hbf8d970d, 32'h3f53d23b} /* (24, 7, 17) {real, imag} */,
  {32'h3d667af6, 32'hbff1743a} /* (24, 7, 16) {real, imag} */,
  {32'hbf02f168, 32'hbefbabf3} /* (24, 7, 15) {real, imag} */,
  {32'h40117946, 32'hbfca6058} /* (24, 7, 14) {real, imag} */,
  {32'hbf921a0e, 32'hc0115ae8} /* (24, 7, 13) {real, imag} */,
  {32'hbefd470c, 32'h3f7a4b57} /* (24, 7, 12) {real, imag} */,
  {32'h3f1ee1a5, 32'hbfbf5105} /* (24, 7, 11) {real, imag} */,
  {32'h403c563c, 32'hbff1fa6b} /* (24, 7, 10) {real, imag} */,
  {32'hbfaa8660, 32'h3ebda981} /* (24, 7, 9) {real, imag} */,
  {32'hbf7d8090, 32'h3fe8ec30} /* (24, 7, 8) {real, imag} */,
  {32'h3f9b9b50, 32'hbe7678bd} /* (24, 7, 7) {real, imag} */,
  {32'hc088387d, 32'hbffbec55} /* (24, 7, 6) {real, imag} */,
  {32'h3fe00cd7, 32'h4076fb7d} /* (24, 7, 5) {real, imag} */,
  {32'h3f3f6969, 32'h3f55a413} /* (24, 7, 4) {real, imag} */,
  {32'hc07ff1bb, 32'h3e9cbd5f} /* (24, 7, 3) {real, imag} */,
  {32'hbf65e14e, 32'hbf590af0} /* (24, 7, 2) {real, imag} */,
  {32'h3fc944ed, 32'h3da8c5b1} /* (24, 7, 1) {real, imag} */,
  {32'hbfe1bc8d, 32'hc093c6b7} /* (24, 7, 0) {real, imag} */,
  {32'hc076475d, 32'hbfaac55a} /* (24, 6, 31) {real, imag} */,
  {32'hbcdba04a, 32'h40a10d38} /* (24, 6, 30) {real, imag} */,
  {32'h4002383b, 32'hbf8a7e1d} /* (24, 6, 29) {real, imag} */,
  {32'h406c1d8e, 32'h409b4062} /* (24, 6, 28) {real, imag} */,
  {32'h408c3e11, 32'h3f986466} /* (24, 6, 27) {real, imag} */,
  {32'hc04abc21, 32'h3f6403bc} /* (24, 6, 26) {real, imag} */,
  {32'hbf5d393c, 32'h404a1e7d} /* (24, 6, 25) {real, imag} */,
  {32'hc02b0991, 32'hbfe19dda} /* (24, 6, 24) {real, imag} */,
  {32'hbfcec06a, 32'hbf93432f} /* (24, 6, 23) {real, imag} */,
  {32'hbf5cf2d6, 32'hc0245e9d} /* (24, 6, 22) {real, imag} */,
  {32'h3f46178b, 32'hbf7ad896} /* (24, 6, 21) {real, imag} */,
  {32'hbf047bc4, 32'hc0015670} /* (24, 6, 20) {real, imag} */,
  {32'h4083f2bd, 32'h404581ef} /* (24, 6, 19) {real, imag} */,
  {32'hc021c5c7, 32'hbfc00ce7} /* (24, 6, 18) {real, imag} */,
  {32'h3f60e330, 32'h3ecd52c1} /* (24, 6, 17) {real, imag} */,
  {32'hbe390bc5, 32'hbeb1752a} /* (24, 6, 16) {real, imag} */,
  {32'h3f45e901, 32'hbfe6adc9} /* (24, 6, 15) {real, imag} */,
  {32'h3f939c85, 32'hbd33ce51} /* (24, 6, 14) {real, imag} */,
  {32'h3fece129, 32'hbe346570} /* (24, 6, 13) {real, imag} */,
  {32'h3f89f65b, 32'h3f9c2a54} /* (24, 6, 12) {real, imag} */,
  {32'hc08be198, 32'h3fab74bc} /* (24, 6, 11) {real, imag} */,
  {32'hc0203493, 32'h404d0d31} /* (24, 6, 10) {real, imag} */,
  {32'h3e7372f4, 32'h3f4964f9} /* (24, 6, 9) {real, imag} */,
  {32'hbf63154e, 32'h3dffbaf6} /* (24, 6, 8) {real, imag} */,
  {32'hbd449725, 32'h407d8057} /* (24, 6, 7) {real, imag} */,
  {32'h3f897e95, 32'hbfd39486} /* (24, 6, 6) {real, imag} */,
  {32'h3ea36240, 32'hc086f02b} /* (24, 6, 5) {real, imag} */,
  {32'h4019a69b, 32'h3f3147fd} /* (24, 6, 4) {real, imag} */,
  {32'h403abadd, 32'hbf8695c7} /* (24, 6, 3) {real, imag} */,
  {32'h3f5886f8, 32'h3edfa4fd} /* (24, 6, 2) {real, imag} */,
  {32'h3f39593f, 32'hc04780cd} /* (24, 6, 1) {real, imag} */,
  {32'hc02525c3, 32'hbea5dace} /* (24, 6, 0) {real, imag} */,
  {32'h4006fdba, 32'h40534277} /* (24, 5, 31) {real, imag} */,
  {32'hbff5c55a, 32'hc04f2798} /* (24, 5, 30) {real, imag} */,
  {32'h3f505465, 32'h3ec1bb26} /* (24, 5, 29) {real, imag} */,
  {32'h3ff07814, 32'hbee0116d} /* (24, 5, 28) {real, imag} */,
  {32'hc0287bfe, 32'h3fa2f215} /* (24, 5, 27) {real, imag} */,
  {32'hbf95c49b, 32'h3f96c37e} /* (24, 5, 26) {real, imag} */,
  {32'h4021b97e, 32'h3f83ad38} /* (24, 5, 25) {real, imag} */,
  {32'hbf9ea7a0, 32'hbf8aac5f} /* (24, 5, 24) {real, imag} */,
  {32'h3f1c34c9, 32'hbdc1d931} /* (24, 5, 23) {real, imag} */,
  {32'hbd595f00, 32'hbe65444e} /* (24, 5, 22) {real, imag} */,
  {32'h3f1e0b19, 32'h402db0c7} /* (24, 5, 21) {real, imag} */,
  {32'hbfc28a58, 32'h3f0ee336} /* (24, 5, 20) {real, imag} */,
  {32'hbeb22f7a, 32'hbf348d97} /* (24, 5, 19) {real, imag} */,
  {32'hbfb7beac, 32'h3fcadea2} /* (24, 5, 18) {real, imag} */,
  {32'hbf13e13b, 32'hbf47d754} /* (24, 5, 17) {real, imag} */,
  {32'h3fdb15c3, 32'h406f5f64} /* (24, 5, 16) {real, imag} */,
  {32'hbf0f88a0, 32'hbfff02f3} /* (24, 5, 15) {real, imag} */,
  {32'hbfaa2d50, 32'h3fc4cfb2} /* (24, 5, 14) {real, imag} */,
  {32'hc0977cd8, 32'hbecf434f} /* (24, 5, 13) {real, imag} */,
  {32'h404c7ec2, 32'h3ec7c731} /* (24, 5, 12) {real, imag} */,
  {32'h3fa5441f, 32'hbeee09e5} /* (24, 5, 11) {real, imag} */,
  {32'hbf20c1d9, 32'hbc7a2994} /* (24, 5, 10) {real, imag} */,
  {32'h3f37444a, 32'h3f556545} /* (24, 5, 9) {real, imag} */,
  {32'h4032c488, 32'hc001635a} /* (24, 5, 8) {real, imag} */,
  {32'hc03df135, 32'h3fbe2a06} /* (24, 5, 7) {real, imag} */,
  {32'h3f6e7bdb, 32'h3e4937ee} /* (24, 5, 6) {real, imag} */,
  {32'h3f9fd05c, 32'h3df9f9d8} /* (24, 5, 5) {real, imag} */,
  {32'h4040f972, 32'hc06c2ede} /* (24, 5, 4) {real, imag} */,
  {32'h3e3cd7b7, 32'h3ca2fab1} /* (24, 5, 3) {real, imag} */,
  {32'h3f936aeb, 32'hc05a7ffa} /* (24, 5, 2) {real, imag} */,
  {32'hbfe92936, 32'h3f763e7c} /* (24, 5, 1) {real, imag} */,
  {32'h3f5fd3f5, 32'h40296de4} /* (24, 5, 0) {real, imag} */,
  {32'hbdc8299f, 32'hc02be5ae} /* (24, 4, 31) {real, imag} */,
  {32'h3fa71b21, 32'h40ca7a8e} /* (24, 4, 30) {real, imag} */,
  {32'h3fac6465, 32'hc0a7c524} /* (24, 4, 29) {real, imag} */,
  {32'hbffa6fef, 32'hbd93ebfb} /* (24, 4, 28) {real, imag} */,
  {32'h3eb1cf76, 32'hc0d8b883} /* (24, 4, 27) {real, imag} */,
  {32'h3f88c44f, 32'h3f1395d3} /* (24, 4, 26) {real, imag} */,
  {32'h3fad5868, 32'h3de11b4e} /* (24, 4, 25) {real, imag} */,
  {32'h401bf96d, 32'hbf89a9db} /* (24, 4, 24) {real, imag} */,
  {32'h3f94da11, 32'hbf70f248} /* (24, 4, 23) {real, imag} */,
  {32'h3ec827b4, 32'hc007e35f} /* (24, 4, 22) {real, imag} */,
  {32'hbf52552a, 32'hbf19328c} /* (24, 4, 21) {real, imag} */,
  {32'hbf1ada8e, 32'h3fa8e3fb} /* (24, 4, 20) {real, imag} */,
  {32'h3f3cc48b, 32'hbf7bda8a} /* (24, 4, 19) {real, imag} */,
  {32'hbfc913db, 32'h40040dfc} /* (24, 4, 18) {real, imag} */,
  {32'hbf2e9fe5, 32'h3fd5aa5a} /* (24, 4, 17) {real, imag} */,
  {32'h3e917385, 32'hbf458cb4} /* (24, 4, 16) {real, imag} */,
  {32'h3ed9593c, 32'h3f0483d6} /* (24, 4, 15) {real, imag} */,
  {32'hbe534efd, 32'h4024f027} /* (24, 4, 14) {real, imag} */,
  {32'h3f9f49c8, 32'hbfd8b267} /* (24, 4, 13) {real, imag} */,
  {32'hbf863f88, 32'hbf9d01c7} /* (24, 4, 12) {real, imag} */,
  {32'hc06b04b5, 32'h408aec72} /* (24, 4, 11) {real, imag} */,
  {32'h3fd24613, 32'h3f125cb5} /* (24, 4, 10) {real, imag} */,
  {32'hc0a1fa89, 32'h3fff493b} /* (24, 4, 9) {real, imag} */,
  {32'h3eb959ad, 32'h3e54f482} /* (24, 4, 8) {real, imag} */,
  {32'h3f492778, 32'hc0a98ea8} /* (24, 4, 7) {real, imag} */,
  {32'h3f0b96f1, 32'hbf0c9868} /* (24, 4, 6) {real, imag} */,
  {32'h3fa91cf5, 32'h3e969e2d} /* (24, 4, 5) {real, imag} */,
  {32'h405c0091, 32'hc08a42c9} /* (24, 4, 4) {real, imag} */,
  {32'hbf963530, 32'hc0a48062} /* (24, 4, 3) {real, imag} */,
  {32'hc015f9c4, 32'h40cc05c6} /* (24, 4, 2) {real, imag} */,
  {32'hbffbbe2b, 32'hc0fd4999} /* (24, 4, 1) {real, imag} */,
  {32'hbe22dbef, 32'hbf7523e4} /* (24, 4, 0) {real, imag} */,
  {32'h40a71ba9, 32'hbf3618d6} /* (24, 3, 31) {real, imag} */,
  {32'hc00b38b9, 32'hbffc2f8c} /* (24, 3, 30) {real, imag} */,
  {32'hc04080a8, 32'h40e52a61} /* (24, 3, 29) {real, imag} */,
  {32'h3fbc2c84, 32'hc0d97ae1} /* (24, 3, 28) {real, imag} */,
  {32'h4027ca12, 32'hbd252fcd} /* (24, 3, 27) {real, imag} */,
  {32'h4079c33d, 32'hc03ed1e7} /* (24, 3, 26) {real, imag} */,
  {32'hbfe6131c, 32'h3f5d336f} /* (24, 3, 25) {real, imag} */,
  {32'hbfe76184, 32'h40534954} /* (24, 3, 24) {real, imag} */,
  {32'h3f71f7fc, 32'h4023b259} /* (24, 3, 23) {real, imag} */,
  {32'h405fc0b6, 32'h3d8d4602} /* (24, 3, 22) {real, imag} */,
  {32'hc0391be9, 32'hc00bbea3} /* (24, 3, 21) {real, imag} */,
  {32'hbe4d225d, 32'h3ffa59c6} /* (24, 3, 20) {real, imag} */,
  {32'hbfd11528, 32'hbf38adf6} /* (24, 3, 19) {real, imag} */,
  {32'hc03943a1, 32'hc0053c07} /* (24, 3, 18) {real, imag} */,
  {32'h3e08aa62, 32'h3fa10f13} /* (24, 3, 17) {real, imag} */,
  {32'hbf6b8482, 32'h3f22fe9a} /* (24, 3, 16) {real, imag} */,
  {32'h3fa0c5ea, 32'h402d8c78} /* (24, 3, 15) {real, imag} */,
  {32'h3e8ed735, 32'hc0375bfc} /* (24, 3, 14) {real, imag} */,
  {32'hc02e29b4, 32'h3fb82e6a} /* (24, 3, 13) {real, imag} */,
  {32'hc0083636, 32'h404d6ff2} /* (24, 3, 12) {real, imag} */,
  {32'hbf131d2c, 32'hbf5f2302} /* (24, 3, 11) {real, imag} */,
  {32'h3ed63b64, 32'hbf260a6f} /* (24, 3, 10) {real, imag} */,
  {32'h3ef48cd2, 32'hbd93712c} /* (24, 3, 9) {real, imag} */,
  {32'h3fe5b1a9, 32'h3e073605} /* (24, 3, 8) {real, imag} */,
  {32'hc000cfd4, 32'hbe84f345} /* (24, 3, 7) {real, imag} */,
  {32'hbffd03ab, 32'h3e830eb3} /* (24, 3, 6) {real, imag} */,
  {32'h3f0b88a5, 32'hc0286c7b} /* (24, 3, 5) {real, imag} */,
  {32'h4016551b, 32'h40162b3a} /* (24, 3, 4) {real, imag} */,
  {32'h4079923f, 32'h406f860d} /* (24, 3, 3) {real, imag} */,
  {32'hc018f632, 32'h3fcf4d99} /* (24, 3, 2) {real, imag} */,
  {32'hbfaac526, 32'hc027b645} /* (24, 3, 1) {real, imag} */,
  {32'h401b26a6, 32'hbf8d57a3} /* (24, 3, 0) {real, imag} */,
  {32'h411fc6b6, 32'h418ec8ab} /* (24, 2, 31) {real, imag} */,
  {32'hc11771e0, 32'hc052697c} /* (24, 2, 30) {real, imag} */,
  {32'h404192d0, 32'h3fe30827} /* (24, 2, 29) {real, imag} */,
  {32'h3fe0ca6b, 32'hbfee1a85} /* (24, 2, 28) {real, imag} */,
  {32'hc0cadcfa, 32'hbf560c02} /* (24, 2, 27) {real, imag} */,
  {32'h403be27b, 32'h4094c0e4} /* (24, 2, 26) {real, imag} */,
  {32'h3f3991d9, 32'h3e6eb536} /* (24, 2, 25) {real, imag} */,
  {32'hc0e5cc89, 32'hbf8b7909} /* (24, 2, 24) {real, imag} */,
  {32'hbfa4da82, 32'h3f8d4278} /* (24, 2, 23) {real, imag} */,
  {32'h3f977384, 32'hbfa257db} /* (24, 2, 22) {real, imag} */,
  {32'h3f80d480, 32'h3f7d7657} /* (24, 2, 21) {real, imag} */,
  {32'hbf4b64ec, 32'hc086130c} /* (24, 2, 20) {real, imag} */,
  {32'h402549c6, 32'hbfe737f8} /* (24, 2, 19) {real, imag} */,
  {32'h3f597afe, 32'hbfdd4f33} /* (24, 2, 18) {real, imag} */,
  {32'hbec70f61, 32'hbca71186} /* (24, 2, 17) {real, imag} */,
  {32'h3f5a4ab6, 32'h3f90c299} /* (24, 2, 16) {real, imag} */,
  {32'hbf2dc6a5, 32'hbe99ca75} /* (24, 2, 15) {real, imag} */,
  {32'hbea0f244, 32'h3eb811ff} /* (24, 2, 14) {real, imag} */,
  {32'h3f1a376c, 32'h3d506f5f} /* (24, 2, 13) {real, imag} */,
  {32'h402c2b10, 32'h402f0620} /* (24, 2, 12) {real, imag} */,
  {32'h3f8b0811, 32'hbeecbb8c} /* (24, 2, 11) {real, imag} */,
  {32'hbfd7ba62, 32'hbf06cfc8} /* (24, 2, 10) {real, imag} */,
  {32'hbdac4e0e, 32'h3f832ec8} /* (24, 2, 9) {real, imag} */,
  {32'hbf015189, 32'hc0883606} /* (24, 2, 8) {real, imag} */,
  {32'hbfb69288, 32'hc02da91c} /* (24, 2, 7) {real, imag} */,
  {32'h3e4d7df5, 32'hbf186f2a} /* (24, 2, 6) {real, imag} */,
  {32'h40183e01, 32'hc0e08e3a} /* (24, 2, 5) {real, imag} */,
  {32'h4086965f, 32'h3ff0e715} /* (24, 2, 4) {real, imag} */,
  {32'h407bf02d, 32'hbfaf7adc} /* (24, 2, 3) {real, imag} */,
  {32'hc136d204, 32'hc1632eec} /* (24, 2, 2) {real, imag} */,
  {32'h413ad087, 32'h3f9e23e5} /* (24, 2, 1) {real, imag} */,
  {32'h4093fb62, 32'h412332ec} /* (24, 2, 0) {real, imag} */,
  {32'hc127fe79, 32'hc130aa59} /* (24, 1, 31) {real, imag} */,
  {32'h40fa8ebe, 32'h40b3c9b3} /* (24, 1, 30) {real, imag} */,
  {32'h3f5fb74e, 32'h3f53c37e} /* (24, 1, 29) {real, imag} */,
  {32'h3fb3eba7, 32'hc0750f12} /* (24, 1, 28) {real, imag} */,
  {32'h4020d0b0, 32'h40d14ab4} /* (24, 1, 27) {real, imag} */,
  {32'hc012d13f, 32'h3f29efec} /* (24, 1, 26) {real, imag} */,
  {32'h4042a95d, 32'hbf0a3d47} /* (24, 1, 25) {real, imag} */,
  {32'h3f1ac76e, 32'hbfd8a2a9} /* (24, 1, 24) {real, imag} */,
  {32'h3f3cb06d, 32'h4087c4d2} /* (24, 1, 23) {real, imag} */,
  {32'hbe7f9e17, 32'hbdbb3276} /* (24, 1, 22) {real, imag} */,
  {32'hbf8aa415, 32'hbfb737a3} /* (24, 1, 21) {real, imag} */,
  {32'h3e945379, 32'hbfa1aab1} /* (24, 1, 20) {real, imag} */,
  {32'h3e14c8ed, 32'h3fd4ac8c} /* (24, 1, 19) {real, imag} */,
  {32'h3f7d2d34, 32'hc07dab9e} /* (24, 1, 18) {real, imag} */,
  {32'hbf5f97ad, 32'h3f733048} /* (24, 1, 17) {real, imag} */,
  {32'hbf927fe3, 32'hbf96aff4} /* (24, 1, 16) {real, imag} */,
  {32'h409cca41, 32'h3dba117c} /* (24, 1, 15) {real, imag} */,
  {32'hbf7e1054, 32'hbc924251} /* (24, 1, 14) {real, imag} */,
  {32'hbe5599f4, 32'hbfaff77f} /* (24, 1, 13) {real, imag} */,
  {32'hc01fc3b8, 32'h3e750a29} /* (24, 1, 12) {real, imag} */,
  {32'h3e8b4a9d, 32'h407772c6} /* (24, 1, 11) {real, imag} */,
  {32'h405be2bd, 32'hc02bd702} /* (24, 1, 10) {real, imag} */,
  {32'hc05525c1, 32'h3f89d94f} /* (24, 1, 9) {real, imag} */,
  {32'hc054765d, 32'h408f18a2} /* (24, 1, 8) {real, imag} */,
  {32'hbfa9ab52, 32'hbe77cb01} /* (24, 1, 7) {real, imag} */,
  {32'hbee83711, 32'hbe61a2ea} /* (24, 1, 6) {real, imag} */,
  {32'h3f68f5d2, 32'h40971572} /* (24, 1, 5) {real, imag} */,
  {32'h4057a30f, 32'h402a42f5} /* (24, 1, 4) {real, imag} */,
  {32'hbe699550, 32'hbf353691} /* (24, 1, 3) {real, imag} */,
  {32'hc0017c6b, 32'h4191019a} /* (24, 1, 2) {real, imag} */,
  {32'hc0b68caa, 32'hc1dcba48} /* (24, 1, 1) {real, imag} */,
  {32'hc10d65e9, 32'hc186824f} /* (24, 1, 0) {real, imag} */,
  {32'hc14d4dab, 32'hc05f092b} /* (24, 0, 31) {real, imag} */,
  {32'h40961550, 32'hc083fece} /* (24, 0, 30) {real, imag} */,
  {32'h3f8078cd, 32'h4096e363} /* (24, 0, 29) {real, imag} */,
  {32'hbec4f62b, 32'hbf992d77} /* (24, 0, 28) {real, imag} */,
  {32'h4085d9f2, 32'h401066ce} /* (24, 0, 27) {real, imag} */,
  {32'h4062294a, 32'hc0494b4b} /* (24, 0, 26) {real, imag} */,
  {32'hc09c5354, 32'hc0494d7f} /* (24, 0, 25) {real, imag} */,
  {32'h4023b349, 32'h4014b47f} /* (24, 0, 24) {real, imag} */,
  {32'h3fb4db4a, 32'hbfc200f0} /* (24, 0, 23) {real, imag} */,
  {32'hc081e7ed, 32'h40737537} /* (24, 0, 22) {real, imag} */,
  {32'h3fe6fb1d, 32'h3f5a5215} /* (24, 0, 21) {real, imag} */,
  {32'hbf86e8e7, 32'hbf970e3b} /* (24, 0, 20) {real, imag} */,
  {32'hbf9b72e1, 32'h3fe4c5ee} /* (24, 0, 19) {real, imag} */,
  {32'h4065b005, 32'hc067e2b1} /* (24, 0, 18) {real, imag} */,
  {32'hc01750a2, 32'hc025af6f} /* (24, 0, 17) {real, imag} */,
  {32'hbf823d68, 32'hbe9eb703} /* (24, 0, 16) {real, imag} */,
  {32'hbf84a399, 32'hbe91a3a3} /* (24, 0, 15) {real, imag} */,
  {32'hbf207fda, 32'hbf1d2b1d} /* (24, 0, 14) {real, imag} */,
  {32'h3e1abb31, 32'h3ff820b6} /* (24, 0, 13) {real, imag} */,
  {32'hbfb4a37b, 32'h3deb692b} /* (24, 0, 12) {real, imag} */,
  {32'hc031ebdd, 32'h3f3becd8} /* (24, 0, 11) {real, imag} */,
  {32'hbeb77af3, 32'h3f189f6c} /* (24, 0, 10) {real, imag} */,
  {32'h3fa571d1, 32'hbf91f7f5} /* (24, 0, 9) {real, imag} */,
  {32'hc086ec75, 32'h3f329e91} /* (24, 0, 8) {real, imag} */,
  {32'h40514d9d, 32'hc025df23} /* (24, 0, 7) {real, imag} */,
  {32'hbfc65bff, 32'h402e2307} /* (24, 0, 6) {real, imag} */,
  {32'hbe7c4009, 32'h40887065} /* (24, 0, 5) {real, imag} */,
  {32'hc0832be1, 32'h3f28d8af} /* (24, 0, 4) {real, imag} */,
  {32'h40251ca1, 32'hbff25aa9} /* (24, 0, 3) {real, imag} */,
  {32'hbfa65c3b, 32'h404fd79b} /* (24, 0, 2) {real, imag} */,
  {32'hc0d6af11, 32'hc16fcae3} /* (24, 0, 1) {real, imag} */,
  {32'hc0a7ed62, 32'hc0ee2d8e} /* (24, 0, 0) {real, imag} */,
  {32'hc0b610c6, 32'h3ed07cdb} /* (23, 31, 31) {real, imag} */,
  {32'h40ab1cac, 32'h4078dc3d} /* (23, 31, 30) {real, imag} */,
  {32'h3ed4e7bd, 32'h410f0324} /* (23, 31, 29) {real, imag} */,
  {32'hbf1c9d85, 32'hc017bdc4} /* (23, 31, 28) {real, imag} */,
  {32'h402a5695, 32'h3efb70a5} /* (23, 31, 27) {real, imag} */,
  {32'h3fd5afbc, 32'h3fc8f943} /* (23, 31, 26) {real, imag} */,
  {32'h3ff9993d, 32'hbfd39f1b} /* (23, 31, 25) {real, imag} */,
  {32'hc03fd469, 32'hc0be2e36} /* (23, 31, 24) {real, imag} */,
  {32'h3fae36fe, 32'hc03b26a2} /* (23, 31, 23) {real, imag} */,
  {32'hbfca08bf, 32'hbfe70597} /* (23, 31, 22) {real, imag} */,
  {32'hbfbcb05e, 32'h3cfb0928} /* (23, 31, 21) {real, imag} */,
  {32'hbf999226, 32'hbeeb1789} /* (23, 31, 20) {real, imag} */,
  {32'hbebbb032, 32'h403796ca} /* (23, 31, 19) {real, imag} */,
  {32'hbfbeeee5, 32'h3f3a040e} /* (23, 31, 18) {real, imag} */,
  {32'h3f2d60eb, 32'h3db55d04} /* (23, 31, 17) {real, imag} */,
  {32'h3f2cd194, 32'h3febdbbf} /* (23, 31, 16) {real, imag} */,
  {32'h3f2339fb, 32'hbfae282e} /* (23, 31, 15) {real, imag} */,
  {32'h3f63549e, 32'h3f683da2} /* (23, 31, 14) {real, imag} */,
  {32'h3fc952e5, 32'h3fdfeb82} /* (23, 31, 13) {real, imag} */,
  {32'hc0491cbc, 32'h3f334756} /* (23, 31, 12) {real, imag} */,
  {32'h3fe0c154, 32'hbf082c7c} /* (23, 31, 11) {real, imag} */,
  {32'h401a184a, 32'h3fac0cde} /* (23, 31, 10) {real, imag} */,
  {32'h3ea061f3, 32'h3fbeebf1} /* (23, 31, 9) {real, imag} */,
  {32'h3f3b8934, 32'h3fa29869} /* (23, 31, 8) {real, imag} */,
  {32'hc02c0a97, 32'hbf99fb0c} /* (23, 31, 7) {real, imag} */,
  {32'hc0812aa1, 32'hc03a4fc4} /* (23, 31, 6) {real, imag} */,
  {32'h3f6715bf, 32'hbfc85114} /* (23, 31, 5) {real, imag} */,
  {32'hbc9e394e, 32'hbfb4ca3b} /* (23, 31, 4) {real, imag} */,
  {32'h3e3f5e91, 32'h3da627d4} /* (23, 31, 3) {real, imag} */,
  {32'h4022aa49, 32'h405c953f} /* (23, 31, 2) {real, imag} */,
  {32'hbf94afa2, 32'hc0891c5a} /* (23, 31, 1) {real, imag} */,
  {32'hc0a72a0d, 32'h4017e4c4} /* (23, 31, 0) {real, imag} */,
  {32'h406c017c, 32'h40820344} /* (23, 30, 31) {real, imag} */,
  {32'h3fe1a416, 32'hc0ee9c4a} /* (23, 30, 30) {real, imag} */,
  {32'hc00e4f6d, 32'hc071f8f4} /* (23, 30, 29) {real, imag} */,
  {32'h3ff2b67b, 32'h408f2e1b} /* (23, 30, 28) {real, imag} */,
  {32'hc02b3f91, 32'h3f8f3f1f} /* (23, 30, 27) {real, imag} */,
  {32'h40226ac5, 32'hbf9ff0c2} /* (23, 30, 26) {real, imag} */,
  {32'h408789f5, 32'h3f6d32a2} /* (23, 30, 25) {real, imag} */,
  {32'hc05ada4d, 32'hbf8eeda7} /* (23, 30, 24) {real, imag} */,
  {32'hbda36622, 32'h3fc1b402} /* (23, 30, 23) {real, imag} */,
  {32'h402b98b8, 32'hc01af434} /* (23, 30, 22) {real, imag} */,
  {32'hc04393b3, 32'h3fbce410} /* (23, 30, 21) {real, imag} */,
  {32'h3f94f51a, 32'h3f10310a} /* (23, 30, 20) {real, imag} */,
  {32'hbf581265, 32'h3f90145d} /* (23, 30, 19) {real, imag} */,
  {32'h401d89c3, 32'h3f065fde} /* (23, 30, 18) {real, imag} */,
  {32'h403496e8, 32'hc0148395} /* (23, 30, 17) {real, imag} */,
  {32'h3fa7fd29, 32'h3e8b7be0} /* (23, 30, 16) {real, imag} */,
  {32'hbf0cad44, 32'hbe9ed13d} /* (23, 30, 15) {real, imag} */,
  {32'h3f9da7fa, 32'hc029cd58} /* (23, 30, 14) {real, imag} */,
  {32'hc04e2125, 32'hbfb61fc7} /* (23, 30, 13) {real, imag} */,
  {32'h3eae206b, 32'h40182c87} /* (23, 30, 12) {real, imag} */,
  {32'h3fdbb9c1, 32'hbf524e41} /* (23, 30, 11) {real, imag} */,
  {32'h405d11a7, 32'hbfa82d3f} /* (23, 30, 10) {real, imag} */,
  {32'hbf7f47e2, 32'h3f6c0d50} /* (23, 30, 9) {real, imag} */,
  {32'hbfa14203, 32'h3f30b40a} /* (23, 30, 8) {real, imag} */,
  {32'h3f2c78b1, 32'hc009e451} /* (23, 30, 7) {real, imag} */,
  {32'h3fbe06ef, 32'hc0424e9b} /* (23, 30, 6) {real, imag} */,
  {32'h3d92a698, 32'hbf83ffb5} /* (23, 30, 5) {real, imag} */,
  {32'hc03396bf, 32'h40850785} /* (23, 30, 4) {real, imag} */,
  {32'hc0a5d16b, 32'hbb7376c4} /* (23, 30, 3) {real, imag} */,
  {32'hbfb882e9, 32'hc0be8d4b} /* (23, 30, 2) {real, imag} */,
  {32'h3f93fb79, 32'h405db407} /* (23, 30, 1) {real, imag} */,
  {32'h3f53835d, 32'h40840c4a} /* (23, 30, 0) {real, imag} */,
  {32'hbe8bf30d, 32'h3fb4151d} /* (23, 29, 31) {real, imag} */,
  {32'hc053c5ba, 32'h40bd31c7} /* (23, 29, 30) {real, imag} */,
  {32'h404a9674, 32'h3f853b92} /* (23, 29, 29) {real, imag} */,
  {32'hbed41e36, 32'hc0581431} /* (23, 29, 28) {real, imag} */,
  {32'h40334283, 32'hbea5eeda} /* (23, 29, 27) {real, imag} */,
  {32'h40196575, 32'h4088867a} /* (23, 29, 26) {real, imag} */,
  {32'hc005189a, 32'hbff818b5} /* (23, 29, 25) {real, imag} */,
  {32'h3ffc95c5, 32'hbf08baad} /* (23, 29, 24) {real, imag} */,
  {32'hbf361f91, 32'h3d75c4b8} /* (23, 29, 23) {real, imag} */,
  {32'hbe3e2f17, 32'hbe986382} /* (23, 29, 22) {real, imag} */,
  {32'hbf3b7e87, 32'hc0670d4c} /* (23, 29, 21) {real, imag} */,
  {32'h3ff64458, 32'h3fa251ae} /* (23, 29, 20) {real, imag} */,
  {32'h3f191754, 32'h40a7dea3} /* (23, 29, 19) {real, imag} */,
  {32'hc033db19, 32'hbf7a9d28} /* (23, 29, 18) {real, imag} */,
  {32'hbf33b5b9, 32'hc00846ad} /* (23, 29, 17) {real, imag} */,
  {32'hbea4cca3, 32'hbf44a1b1} /* (23, 29, 16) {real, imag} */,
  {32'h400a3db8, 32'h3f0e127a} /* (23, 29, 15) {real, imag} */,
  {32'hc01c6b5a, 32'hbe2bd09e} /* (23, 29, 14) {real, imag} */,
  {32'h4022bbf5, 32'h3e5c62a2} /* (23, 29, 13) {real, imag} */,
  {32'h3e2141a4, 32'hbfa4d060} /* (23, 29, 12) {real, imag} */,
  {32'h3f0bf89d, 32'h3f926f3a} /* (23, 29, 11) {real, imag} */,
  {32'hc03c504f, 32'hbdb1a6bb} /* (23, 29, 10) {real, imag} */,
  {32'hbfaaa029, 32'h407008b7} /* (23, 29, 9) {real, imag} */,
  {32'hbbe86860, 32'hbf0e52b9} /* (23, 29, 8) {real, imag} */,
  {32'h3fd6c827, 32'hbff7427a} /* (23, 29, 7) {real, imag} */,
  {32'h3f881e1f, 32'h40236057} /* (23, 29, 6) {real, imag} */,
  {32'h3f5302ff, 32'hbf8134fb} /* (23, 29, 5) {real, imag} */,
  {32'hbdac85c4, 32'hbf7f6ce6} /* (23, 29, 4) {real, imag} */,
  {32'h406d8087, 32'hbefe7171} /* (23, 29, 3) {real, imag} */,
  {32'hbea7d01e, 32'hbf9979e6} /* (23, 29, 2) {real, imag} */,
  {32'hbdea6b3b, 32'hbe225eab} /* (23, 29, 1) {real, imag} */,
  {32'h4045de60, 32'h3eef567a} /* (23, 29, 0) {real, imag} */,
  {32'hbe443d65, 32'hbfb28a2a} /* (23, 28, 31) {real, imag} */,
  {32'hbd6f8a91, 32'hbf654a3d} /* (23, 28, 30) {real, imag} */,
  {32'h4083391c, 32'hbe5633e7} /* (23, 28, 29) {real, imag} */,
  {32'hbf747114, 32'hbf8a411f} /* (23, 28, 28) {real, imag} */,
  {32'hbf82a5df, 32'h3f3a1b57} /* (23, 28, 27) {real, imag} */,
  {32'hc0784cf0, 32'hc01fade9} /* (23, 28, 26) {real, imag} */,
  {32'h3f59c70c, 32'h3fccdbdc} /* (23, 28, 25) {real, imag} */,
  {32'hbf998bae, 32'h3f920c4f} /* (23, 28, 24) {real, imag} */,
  {32'h3fda0671, 32'hc0292900} /* (23, 28, 23) {real, imag} */,
  {32'h3fad266e, 32'h4005ebd4} /* (23, 28, 22) {real, imag} */,
  {32'h408531b1, 32'h3fbb0f39} /* (23, 28, 21) {real, imag} */,
  {32'hbef2e2dd, 32'h3febfb49} /* (23, 28, 20) {real, imag} */,
  {32'h3fba47ef, 32'hbfc6594d} /* (23, 28, 19) {real, imag} */,
  {32'h3f492bfb, 32'h3f7e170f} /* (23, 28, 18) {real, imag} */,
  {32'hc01a2f13, 32'hbf91cf40} /* (23, 28, 17) {real, imag} */,
  {32'hbf09c9f0, 32'hbf443f13} /* (23, 28, 16) {real, imag} */,
  {32'hbfce91d2, 32'hbf351988} /* (23, 28, 15) {real, imag} */,
  {32'h3f9c1a1b, 32'hbf8f23d5} /* (23, 28, 14) {real, imag} */,
  {32'h3d95979c, 32'hc021d9e9} /* (23, 28, 13) {real, imag} */,
  {32'h3f21fea5, 32'hc014fb1d} /* (23, 28, 12) {real, imag} */,
  {32'h3f363454, 32'h3fe2c579} /* (23, 28, 11) {real, imag} */,
  {32'hc0600d20, 32'h400f678d} /* (23, 28, 10) {real, imag} */,
  {32'hbff022d4, 32'h3fc33b4a} /* (23, 28, 9) {real, imag} */,
  {32'hc014912e, 32'hbfcf76cc} /* (23, 28, 8) {real, imag} */,
  {32'h40b9470c, 32'hbf8e863e} /* (23, 28, 7) {real, imag} */,
  {32'h3f513d3a, 32'hc02c195a} /* (23, 28, 6) {real, imag} */,
  {32'hc072ed4d, 32'hc099880e} /* (23, 28, 5) {real, imag} */,
  {32'h40007c0c, 32'h3ef1241d} /* (23, 28, 4) {real, imag} */,
  {32'h3f23121f, 32'hc08ab943} /* (23, 28, 3) {real, imag} */,
  {32'h3fd7c9d6, 32'h3feec363} /* (23, 28, 2) {real, imag} */,
  {32'h3ff0ade2, 32'hbf894f97} /* (23, 28, 1) {real, imag} */,
  {32'h3e3e2208, 32'hbf032feb} /* (23, 28, 0) {real, imag} */,
  {32'h3fddb791, 32'h3f3754df} /* (23, 27, 31) {real, imag} */,
  {32'h3fb3450d, 32'h401838b8} /* (23, 27, 30) {real, imag} */,
  {32'hc04ab467, 32'h3ec9c2c0} /* (23, 27, 29) {real, imag} */,
  {32'hbfc096d6, 32'hc01b6a1b} /* (23, 27, 28) {real, imag} */,
  {32'h4014c1e1, 32'h3ddab100} /* (23, 27, 27) {real, imag} */,
  {32'hc06c66a5, 32'h3e7aac49} /* (23, 27, 26) {real, imag} */,
  {32'h403e23d5, 32'h3e47d633} /* (23, 27, 25) {real, imag} */,
  {32'h3e2dbcb3, 32'h3f6d4a2b} /* (23, 27, 24) {real, imag} */,
  {32'h403293e9, 32'h4008045d} /* (23, 27, 23) {real, imag} */,
  {32'hbe8b0948, 32'hbea871da} /* (23, 27, 22) {real, imag} */,
  {32'hc0283eec, 32'h40b13eea} /* (23, 27, 21) {real, imag} */,
  {32'h3fd949df, 32'hbf4478ea} /* (23, 27, 20) {real, imag} */,
  {32'h40102ddb, 32'h3f993dde} /* (23, 27, 19) {real, imag} */,
  {32'hbea96874, 32'hbf51a117} /* (23, 27, 18) {real, imag} */,
  {32'h3fb8b85d, 32'h40550381} /* (23, 27, 17) {real, imag} */,
  {32'hbeac56ea, 32'h3ea25177} /* (23, 27, 16) {real, imag} */,
  {32'h3f1c9598, 32'h3f3427d8} /* (23, 27, 15) {real, imag} */,
  {32'h4002498d, 32'h3e8e77f6} /* (23, 27, 14) {real, imag} */,
  {32'h40a0aef1, 32'h40165597} /* (23, 27, 13) {real, imag} */,
  {32'hbce4a788, 32'hbfe2e1ac} /* (23, 27, 12) {real, imag} */,
  {32'hbfdb40b8, 32'hbf37eb17} /* (23, 27, 11) {real, imag} */,
  {32'h3fe82b0c, 32'h3e09f7dd} /* (23, 27, 10) {real, imag} */,
  {32'hbfc3ffad, 32'h403bff91} /* (23, 27, 9) {real, imag} */,
  {32'hbfcd482e, 32'h40a0859f} /* (23, 27, 8) {real, imag} */,
  {32'h3e129b63, 32'hc00106e8} /* (23, 27, 7) {real, imag} */,
  {32'h3fbf5924, 32'h3e61f20b} /* (23, 27, 6) {real, imag} */,
  {32'h3ed14f0b, 32'hc006b1ed} /* (23, 27, 5) {real, imag} */,
  {32'h3ff02108, 32'h3fba0b79} /* (23, 27, 4) {real, imag} */,
  {32'hc012c316, 32'h405094f8} /* (23, 27, 3) {real, imag} */,
  {32'hc04bac71, 32'hc00075f2} /* (23, 27, 2) {real, imag} */,
  {32'hbe6f2eba, 32'h4002c889} /* (23, 27, 1) {real, imag} */,
  {32'h4029aef4, 32'h403d7f3b} /* (23, 27, 0) {real, imag} */,
  {32'h403c063b, 32'h3f669e22} /* (23, 26, 31) {real, imag} */,
  {32'h3f9989d2, 32'hc0a0dfbe} /* (23, 26, 30) {real, imag} */,
  {32'h3f36c393, 32'hbeaddc1d} /* (23, 26, 29) {real, imag} */,
  {32'hc01d2098, 32'h403cd6fc} /* (23, 26, 28) {real, imag} */,
  {32'hc023d39b, 32'hbf19a6e6} /* (23, 26, 27) {real, imag} */,
  {32'hbfb9fccc, 32'h4022f7a1} /* (23, 26, 26) {real, imag} */,
  {32'h3fd834b4, 32'h3fb39f1a} /* (23, 26, 25) {real, imag} */,
  {32'h40021d0f, 32'h3f8d7ee4} /* (23, 26, 24) {real, imag} */,
  {32'h3f3896c3, 32'hbee328ca} /* (23, 26, 23) {real, imag} */,
  {32'h3fba306f, 32'h3f188372} /* (23, 26, 22) {real, imag} */,
  {32'hbf3ca313, 32'h4071c129} /* (23, 26, 21) {real, imag} */,
  {32'h407ee619, 32'hbe70f368} /* (23, 26, 20) {real, imag} */,
  {32'h3fd32a1f, 32'h3f895a10} /* (23, 26, 19) {real, imag} */,
  {32'hbfc108f7, 32'hc00be29f} /* (23, 26, 18) {real, imag} */,
  {32'h3f1a7ebd, 32'hbf7fa184} /* (23, 26, 17) {real, imag} */,
  {32'h3fd39da0, 32'h3f50e2be} /* (23, 26, 16) {real, imag} */,
  {32'hbda15e16, 32'h3edb142b} /* (23, 26, 15) {real, imag} */,
  {32'hc00425e6, 32'hc0037391} /* (23, 26, 14) {real, imag} */,
  {32'h3eb91dcd, 32'hbf1e5d0b} /* (23, 26, 13) {real, imag} */,
  {32'hbfd34540, 32'hc03fb550} /* (23, 26, 12) {real, imag} */,
  {32'h3ed1990d, 32'h3f04e1c5} /* (23, 26, 11) {real, imag} */,
  {32'h3ec369d7, 32'h3d802423} /* (23, 26, 10) {real, imag} */,
  {32'h4072ffd5, 32'hbf8a8c5d} /* (23, 26, 9) {real, imag} */,
  {32'h3f96f40d, 32'hbf4b4d0e} /* (23, 26, 8) {real, imag} */,
  {32'h3f2db2ff, 32'h3ee63088} /* (23, 26, 7) {real, imag} */,
  {32'h3fe628f7, 32'hc0a179ce} /* (23, 26, 6) {real, imag} */,
  {32'h3ecef923, 32'h3f41e415} /* (23, 26, 5) {real, imag} */,
  {32'hbfbd5c16, 32'h3fb51d7e} /* (23, 26, 4) {real, imag} */,
  {32'h3e9dd5a8, 32'hbeddd2a6} /* (23, 26, 3) {real, imag} */,
  {32'h402f741c, 32'hc004b847} /* (23, 26, 2) {real, imag} */,
  {32'h403ca14f, 32'h3f569625} /* (23, 26, 1) {real, imag} */,
  {32'hc076aa4f, 32'hbec47798} /* (23, 26, 0) {real, imag} */,
  {32'hbf625f1d, 32'h408ace93} /* (23, 25, 31) {real, imag} */,
  {32'hc056a3a7, 32'h3f45057f} /* (23, 25, 30) {real, imag} */,
  {32'hbf8afb51, 32'hc0186e39} /* (23, 25, 29) {real, imag} */,
  {32'hc02fe68e, 32'hbeaf2795} /* (23, 25, 28) {real, imag} */,
  {32'h3e7a5752, 32'h3fb1cadf} /* (23, 25, 27) {real, imag} */,
  {32'h3f556517, 32'hbf33b8fa} /* (23, 25, 26) {real, imag} */,
  {32'hbfe6374c, 32'hbf7db322} /* (23, 25, 25) {real, imag} */,
  {32'hbfe6e0cc, 32'h40991d2c} /* (23, 25, 24) {real, imag} */,
  {32'hc003262e, 32'hbf81e0e7} /* (23, 25, 23) {real, imag} */,
  {32'hbfed6608, 32'h3fb94a08} /* (23, 25, 22) {real, imag} */,
  {32'h3f9d9882, 32'hbf2f6a5d} /* (23, 25, 21) {real, imag} */,
  {32'hc00bce92, 32'hc02f9a16} /* (23, 25, 20) {real, imag} */,
  {32'hbf1e3a27, 32'hc0a4a81d} /* (23, 25, 19) {real, imag} */,
  {32'h3f7001ec, 32'hbf718d8e} /* (23, 25, 18) {real, imag} */,
  {32'hbfdb9301, 32'hbf12c45c} /* (23, 25, 17) {real, imag} */,
  {32'hbfc5a2ef, 32'hbef36fae} /* (23, 25, 16) {real, imag} */,
  {32'hbfb15951, 32'hbf280180} /* (23, 25, 15) {real, imag} */,
  {32'h3fd8ae0d, 32'h3fd4ef6c} /* (23, 25, 14) {real, imag} */,
  {32'hbfcca234, 32'hc017d3fc} /* (23, 25, 13) {real, imag} */,
  {32'h402a3d88, 32'h4089d349} /* (23, 25, 12) {real, imag} */,
  {32'hbea8fa71, 32'h3f76212e} /* (23, 25, 11) {real, imag} */,
  {32'hbf8c040f, 32'hbe3961a9} /* (23, 25, 10) {real, imag} */,
  {32'h40022acd, 32'h3f34b0f9} /* (23, 25, 9) {real, imag} */,
  {32'hc0dd9195, 32'hbc93c59e} /* (23, 25, 8) {real, imag} */,
  {32'hbf63a57c, 32'h3ecbf20c} /* (23, 25, 7) {real, imag} */,
  {32'hbee46497, 32'h407dfc36} /* (23, 25, 6) {real, imag} */,
  {32'h3f376268, 32'h402a42fd} /* (23, 25, 5) {real, imag} */,
  {32'h409df532, 32'hbee83376} /* (23, 25, 4) {real, imag} */,
  {32'hc009f2f7, 32'h3fba51ff} /* (23, 25, 3) {real, imag} */,
  {32'h4005c648, 32'hc04d1323} /* (23, 25, 2) {real, imag} */,
  {32'hbf3df1dc, 32'hbe87bf23} /* (23, 25, 1) {real, imag} */,
  {32'hc0225ccb, 32'hc00c7df1} /* (23, 25, 0) {real, imag} */,
  {32'h4058c030, 32'h3f97c090} /* (23, 24, 31) {real, imag} */,
  {32'h3e0d8906, 32'hbea2361d} /* (23, 24, 30) {real, imag} */,
  {32'h3f550148, 32'h3fe3c3f3} /* (23, 24, 29) {real, imag} */,
  {32'h3fa90101, 32'hc07ce36d} /* (23, 24, 28) {real, imag} */,
  {32'hc0984ad0, 32'hbfc0987c} /* (23, 24, 27) {real, imag} */,
  {32'hbfe8e60d, 32'hbef38d90} /* (23, 24, 26) {real, imag} */,
  {32'hbf6668d7, 32'h3f9ca17b} /* (23, 24, 25) {real, imag} */,
  {32'hbf4f03b3, 32'hbfb9c8d7} /* (23, 24, 24) {real, imag} */,
  {32'hbece7c44, 32'h408b5067} /* (23, 24, 23) {real, imag} */,
  {32'h3ed5e31a, 32'h40731855} /* (23, 24, 22) {real, imag} */,
  {32'h3fcfd71f, 32'hbf844d17} /* (23, 24, 21) {real, imag} */,
  {32'hbfa94c56, 32'hc0097a58} /* (23, 24, 20) {real, imag} */,
  {32'hbfef0b3d, 32'hbe05fc50} /* (23, 24, 19) {real, imag} */,
  {32'h40192b43, 32'hbe87386a} /* (23, 24, 18) {real, imag} */,
  {32'hbf7e410d, 32'h400661c5} /* (23, 24, 17) {real, imag} */,
  {32'hbf745773, 32'h3fd1e5e2} /* (23, 24, 16) {real, imag} */,
  {32'hc037dbc4, 32'hbe9aa30e} /* (23, 24, 15) {real, imag} */,
  {32'h3e93df68, 32'h3f4b01fc} /* (23, 24, 14) {real, imag} */,
  {32'hbdaf4aaf, 32'hc0549abb} /* (23, 24, 13) {real, imag} */,
  {32'hbeb0af6e, 32'hbf060d19} /* (23, 24, 12) {real, imag} */,
  {32'hc02dff8a, 32'hbfb8c80d} /* (23, 24, 11) {real, imag} */,
  {32'h3f804f97, 32'h3f8ff5c4} /* (23, 24, 10) {real, imag} */,
  {32'h3d4dd413, 32'hbd636c87} /* (23, 24, 9) {real, imag} */,
  {32'hbf910e8a, 32'h40033889} /* (23, 24, 8) {real, imag} */,
  {32'hbea6aa0b, 32'h3e67cb85} /* (23, 24, 7) {real, imag} */,
  {32'h40b0e5f6, 32'h3f2bf2e6} /* (23, 24, 6) {real, imag} */,
  {32'h3eb6036f, 32'h3f3087dd} /* (23, 24, 5) {real, imag} */,
  {32'hbf1cb02e, 32'h40050079} /* (23, 24, 4) {real, imag} */,
  {32'h3f36a20e, 32'hbfc9acf7} /* (23, 24, 3) {real, imag} */,
  {32'hbff96900, 32'hbfc8e5be} /* (23, 24, 2) {real, imag} */,
  {32'hc07b5bd9, 32'h3fb9f17b} /* (23, 24, 1) {real, imag} */,
  {32'h40d79b1a, 32'h3f198ed6} /* (23, 24, 0) {real, imag} */,
  {32'hbfcb7f9c, 32'h3fb97542} /* (23, 23, 31) {real, imag} */,
  {32'h3fe67506, 32'hbfb106da} /* (23, 23, 30) {real, imag} */,
  {32'h3fbe2006, 32'hbd8736b3} /* (23, 23, 29) {real, imag} */,
  {32'h3f4b679d, 32'h40254adf} /* (23, 23, 28) {real, imag} */,
  {32'h4009c474, 32'hbdf85654} /* (23, 23, 27) {real, imag} */,
  {32'h3f3d8c92, 32'h400ecceb} /* (23, 23, 26) {real, imag} */,
  {32'hc05cd6c3, 32'h3fc3f7eb} /* (23, 23, 25) {real, imag} */,
  {32'hc019e2bc, 32'h3fa82735} /* (23, 23, 24) {real, imag} */,
  {32'hc00264eb, 32'h3fe4575b} /* (23, 23, 23) {real, imag} */,
  {32'h3ff8e9b5, 32'hc06cee5d} /* (23, 23, 22) {real, imag} */,
  {32'hc00dda31, 32'hbfda676c} /* (23, 23, 21) {real, imag} */,
  {32'hc0229e00, 32'h406ddd51} /* (23, 23, 20) {real, imag} */,
  {32'hbed9019c, 32'hbea0ee6f} /* (23, 23, 19) {real, imag} */,
  {32'hbf8471f5, 32'hbfecf7d0} /* (23, 23, 18) {real, imag} */,
  {32'hbef9ae05, 32'h3f1aded0} /* (23, 23, 17) {real, imag} */,
  {32'h3e0e76dc, 32'h3ff7a879} /* (23, 23, 16) {real, imag} */,
  {32'hbf39f8f1, 32'h3fcefdfd} /* (23, 23, 15) {real, imag} */,
  {32'h3bc98101, 32'hbe5a2630} /* (23, 23, 14) {real, imag} */,
  {32'h402c9d8a, 32'h40339f9d} /* (23, 23, 13) {real, imag} */,
  {32'h3fe827ef, 32'hbfdfdbd4} /* (23, 23, 12) {real, imag} */,
  {32'h400284d4, 32'h3f2c123c} /* (23, 23, 11) {real, imag} */,
  {32'h3e0ce500, 32'h4088bf68} /* (23, 23, 10) {real, imag} */,
  {32'hbe0c3a69, 32'hbe5bdd8b} /* (23, 23, 9) {real, imag} */,
  {32'h3ddfaf54, 32'hbe6f1be3} /* (23, 23, 8) {real, imag} */,
  {32'hc02f73ac, 32'hc005a414} /* (23, 23, 7) {real, imag} */,
  {32'hc03b030c, 32'h401181c5} /* (23, 23, 6) {real, imag} */,
  {32'hbf5a2846, 32'h3eea76a3} /* (23, 23, 5) {real, imag} */,
  {32'h3fce36f8, 32'hbfbcb4e5} /* (23, 23, 4) {real, imag} */,
  {32'h3f327902, 32'hbf06937a} /* (23, 23, 3) {real, imag} */,
  {32'h401988ff, 32'h3febee37} /* (23, 23, 2) {real, imag} */,
  {32'hc022111f, 32'hbfd6d9a6} /* (23, 23, 1) {real, imag} */,
  {32'hbfb6e826, 32'hc065a94e} /* (23, 23, 0) {real, imag} */,
  {32'hbeff9441, 32'h3cab2acb} /* (23, 22, 31) {real, imag} */,
  {32'h409cbffb, 32'hbeab053d} /* (23, 22, 30) {real, imag} */,
  {32'hc028c3a6, 32'hc0372761} /* (23, 22, 29) {real, imag} */,
  {32'h3cda1e06, 32'hbf90d47f} /* (23, 22, 28) {real, imag} */,
  {32'h3f3fc053, 32'hbfaef594} /* (23, 22, 27) {real, imag} */,
  {32'hbe6f66f4, 32'h3f5b8c4a} /* (23, 22, 26) {real, imag} */,
  {32'hbff9ce8c, 32'h3f50f466} /* (23, 22, 25) {real, imag} */,
  {32'h3f4ae95b, 32'h3facb308} /* (23, 22, 24) {real, imag} */,
  {32'h3f6dbd98, 32'hbf82a51e} /* (23, 22, 23) {real, imag} */,
  {32'hbee21476, 32'h3ffd04ae} /* (23, 22, 22) {real, imag} */,
  {32'h402ca666, 32'hbd85e7fb} /* (23, 22, 21) {real, imag} */,
  {32'h3fbc4052, 32'h3fbc6e45} /* (23, 22, 20) {real, imag} */,
  {32'hbee0a02b, 32'h3fbbbd7c} /* (23, 22, 19) {real, imag} */,
  {32'hbea6b2ea, 32'h403552e2} /* (23, 22, 18) {real, imag} */,
  {32'hc002f9bb, 32'h40068384} /* (23, 22, 17) {real, imag} */,
  {32'h3fc05df6, 32'hc0211ae2} /* (23, 22, 16) {real, imag} */,
  {32'h3fc6e694, 32'h3f203fea} /* (23, 22, 15) {real, imag} */,
  {32'h3f9d2c70, 32'h403753e7} /* (23, 22, 14) {real, imag} */,
  {32'hc08a4673, 32'h40097116} /* (23, 22, 13) {real, imag} */,
  {32'hbe81cfcb, 32'h408ee777} /* (23, 22, 12) {real, imag} */,
  {32'h4023837e, 32'hbeb47964} /* (23, 22, 11) {real, imag} */,
  {32'hbf629766, 32'hbfd02024} /* (23, 22, 10) {real, imag} */,
  {32'h402b5225, 32'hc010a382} /* (23, 22, 9) {real, imag} */,
  {32'hbf5cdaae, 32'hc01619c8} /* (23, 22, 8) {real, imag} */,
  {32'h40098d08, 32'hba9aecbf} /* (23, 22, 7) {real, imag} */,
  {32'h3fa69518, 32'hc01e8f20} /* (23, 22, 6) {real, imag} */,
  {32'h40511454, 32'h3fcbe563} /* (23, 22, 5) {real, imag} */,
  {32'h3e38411e, 32'hbf13cea0} /* (23, 22, 4) {real, imag} */,
  {32'h3eceae8f, 32'h3f89dc8b} /* (23, 22, 3) {real, imag} */,
  {32'hc0284e2c, 32'h3f2622fa} /* (23, 22, 2) {real, imag} */,
  {32'h3f79a495, 32'h3fa0fe17} /* (23, 22, 1) {real, imag} */,
  {32'hbfae5fff, 32'hbf7779ee} /* (23, 22, 0) {real, imag} */,
  {32'h4020f36d, 32'hbf1e9735} /* (23, 21, 31) {real, imag} */,
  {32'hbe6d371b, 32'hbfc73765} /* (23, 21, 30) {real, imag} */,
  {32'hbff20695, 32'hc080ddd9} /* (23, 21, 29) {real, imag} */,
  {32'h3fce272b, 32'h3fa4a288} /* (23, 21, 28) {real, imag} */,
  {32'h40436bc9, 32'hc0652a47} /* (23, 21, 27) {real, imag} */,
  {32'h3f7beeaa, 32'hc01129d5} /* (23, 21, 26) {real, imag} */,
  {32'h40175d68, 32'hbfdadbae} /* (23, 21, 25) {real, imag} */,
  {32'h40063b05, 32'hbfd48214} /* (23, 21, 24) {real, imag} */,
  {32'h405c94b1, 32'h3e1478a1} /* (23, 21, 23) {real, imag} */,
  {32'h3fe16bfc, 32'hc0812dca} /* (23, 21, 22) {real, imag} */,
  {32'hc02ea8b1, 32'h3e5fc7da} /* (23, 21, 21) {real, imag} */,
  {32'h3fbad6dc, 32'hbfa1eaf9} /* (23, 21, 20) {real, imag} */,
  {32'h3e6412cd, 32'hbfec2fdb} /* (23, 21, 19) {real, imag} */,
  {32'h3fe73e75, 32'hbf293f4d} /* (23, 21, 18) {real, imag} */,
  {32'hbfe3a2be, 32'hbfbd23aa} /* (23, 21, 17) {real, imag} */,
  {32'hbe9d34e6, 32'h3f8e0200} /* (23, 21, 16) {real, imag} */,
  {32'h3fa536c5, 32'h402775c0} /* (23, 21, 15) {real, imag} */,
  {32'hbe72262c, 32'hbfefe00b} /* (23, 21, 14) {real, imag} */,
  {32'h3ffada80, 32'h3f87f42a} /* (23, 21, 13) {real, imag} */,
  {32'h3f906ecc, 32'h400a6f88} /* (23, 21, 12) {real, imag} */,
  {32'hc03faa41, 32'h4042deae} /* (23, 21, 11) {real, imag} */,
  {32'hbda72796, 32'hbfee1654} /* (23, 21, 10) {real, imag} */,
  {32'hc08272bb, 32'h3ef36b3c} /* (23, 21, 9) {real, imag} */,
  {32'h405e1900, 32'h3e7874ee} /* (23, 21, 8) {real, imag} */,
  {32'h40854ae2, 32'hc01599a9} /* (23, 21, 7) {real, imag} */,
  {32'h3fa9c588, 32'hc0104b74} /* (23, 21, 6) {real, imag} */,
  {32'hc082594b, 32'hbfa77802} /* (23, 21, 5) {real, imag} */,
  {32'hbfc40310, 32'h3eeb4664} /* (23, 21, 4) {real, imag} */,
  {32'hc026f07a, 32'h3f66638d} /* (23, 21, 3) {real, imag} */,
  {32'hbe96f736, 32'h400be92c} /* (23, 21, 2) {real, imag} */,
  {32'hbf320b7f, 32'h3f4afcc1} /* (23, 21, 1) {real, imag} */,
  {32'hc029d401, 32'hbf886829} /* (23, 21, 0) {real, imag} */,
  {32'h4017e819, 32'h3fbc6fae} /* (23, 20, 31) {real, imag} */,
  {32'h401145ff, 32'hbf024809} /* (23, 20, 30) {real, imag} */,
  {32'hbfbcf93e, 32'hbd2d99ee} /* (23, 20, 29) {real, imag} */,
  {32'h3f19756f, 32'hbeb8ad75} /* (23, 20, 28) {real, imag} */,
  {32'h3fa04d8f, 32'h3ff1573b} /* (23, 20, 27) {real, imag} */,
  {32'h3f3f1d99, 32'hbf656beb} /* (23, 20, 26) {real, imag} */,
  {32'h3fe38429, 32'hbebbb3bf} /* (23, 20, 25) {real, imag} */,
  {32'hbd6b0d36, 32'hc009f749} /* (23, 20, 24) {real, imag} */,
  {32'h3c27b10d, 32'h40226588} /* (23, 20, 23) {real, imag} */,
  {32'hbf79577f, 32'hbff68c1e} /* (23, 20, 22) {real, imag} */,
  {32'h3fe2fa5f, 32'h3f66522c} /* (23, 20, 21) {real, imag} */,
  {32'h3fa5325f, 32'h3e1b4b1f} /* (23, 20, 20) {real, imag} */,
  {32'h3ff4eceb, 32'hbfe84b38} /* (23, 20, 19) {real, imag} */,
  {32'h3f0a0db5, 32'h3f7bd7ab} /* (23, 20, 18) {real, imag} */,
  {32'hbeabe509, 32'h3f6b7d0d} /* (23, 20, 17) {real, imag} */,
  {32'hc019fb8b, 32'h3f5aaa89} /* (23, 20, 16) {real, imag} */,
  {32'h4022c8f8, 32'hbf34fc0b} /* (23, 20, 15) {real, imag} */,
  {32'h406b1ad3, 32'hbef1a48a} /* (23, 20, 14) {real, imag} */,
  {32'h400f5ef9, 32'h3f0047e6} /* (23, 20, 13) {real, imag} */,
  {32'h3eb82e41, 32'hbdbab44f} /* (23, 20, 12) {real, imag} */,
  {32'h3fe6190d, 32'hc08970c6} /* (23, 20, 11) {real, imag} */,
  {32'hbfc13925, 32'h3faa2699} /* (23, 20, 10) {real, imag} */,
  {32'hbf9d983e, 32'hc050a318} /* (23, 20, 9) {real, imag} */,
  {32'h3fd551d4, 32'hbfb19888} /* (23, 20, 8) {real, imag} */,
  {32'hbf2d23b1, 32'h3ffd2219} /* (23, 20, 7) {real, imag} */,
  {32'hc04741f7, 32'hc030b850} /* (23, 20, 6) {real, imag} */,
  {32'hbf604ae0, 32'h40102067} /* (23, 20, 5) {real, imag} */,
  {32'hbe6e5ac1, 32'hbfe48789} /* (23, 20, 4) {real, imag} */,
  {32'hc01edcfa, 32'hbeb3473e} /* (23, 20, 3) {real, imag} */,
  {32'hbf2e980a, 32'hbed33c99} /* (23, 20, 2) {real, imag} */,
  {32'h3fecb699, 32'hc0280949} /* (23, 20, 1) {real, imag} */,
  {32'hbfc99c3d, 32'hbf0acaaf} /* (23, 20, 0) {real, imag} */,
  {32'hc023ccc4, 32'h3f4a415c} /* (23, 19, 31) {real, imag} */,
  {32'hbf5b566c, 32'h3fcfa0ce} /* (23, 19, 30) {real, imag} */,
  {32'hbf31c132, 32'h40240681} /* (23, 19, 29) {real, imag} */,
  {32'h40587ba0, 32'hbf59d3fc} /* (23, 19, 28) {real, imag} */,
  {32'hc05657e9, 32'hbfbe896f} /* (23, 19, 27) {real, imag} */,
  {32'h3d742bc8, 32'hbf93f0b4} /* (23, 19, 26) {real, imag} */,
  {32'hbd0e830a, 32'h3d149e4e} /* (23, 19, 25) {real, imag} */,
  {32'hbfda96f6, 32'h3f84e225} /* (23, 19, 24) {real, imag} */,
  {32'hc033a6be, 32'hc003ad44} /* (23, 19, 23) {real, imag} */,
  {32'hc0257d2d, 32'hbfd948df} /* (23, 19, 22) {real, imag} */,
  {32'h407b2778, 32'h3fe09245} /* (23, 19, 21) {real, imag} */,
  {32'hbec284bc, 32'hc04f7c50} /* (23, 19, 20) {real, imag} */,
  {32'h3f9365a1, 32'hbff651fd} /* (23, 19, 19) {real, imag} */,
  {32'h3e1beadf, 32'hbf254493} /* (23, 19, 18) {real, imag} */,
  {32'hbf780e0f, 32'h3ef8c572} /* (23, 19, 17) {real, imag} */,
  {32'hbe3d89c6, 32'hbde0ea18} /* (23, 19, 16) {real, imag} */,
  {32'h3faaa389, 32'hbfb35754} /* (23, 19, 15) {real, imag} */,
  {32'h3ed59c9b, 32'h3e175254} /* (23, 19, 14) {real, imag} */,
  {32'h3f1e4111, 32'hc0609a50} /* (23, 19, 13) {real, imag} */,
  {32'hbe543ce2, 32'h40296ab6} /* (23, 19, 12) {real, imag} */,
  {32'h3e8c453d, 32'hbf29fe08} /* (23, 19, 11) {real, imag} */,
  {32'h3fa3129c, 32'h3fc945ac} /* (23, 19, 10) {real, imag} */,
  {32'h3ef3d317, 32'h3f960a41} /* (23, 19, 9) {real, imag} */,
  {32'h3f8a1812, 32'h4042a340} /* (23, 19, 8) {real, imag} */,
  {32'h3efe313e, 32'hbf295541} /* (23, 19, 7) {real, imag} */,
  {32'hbfd6ac68, 32'h3f72be00} /* (23, 19, 6) {real, imag} */,
  {32'h3ef800ec, 32'h3f4a9435} /* (23, 19, 5) {real, imag} */,
  {32'h3f177e7a, 32'h404d31bb} /* (23, 19, 4) {real, imag} */,
  {32'h3e165320, 32'hbfc80033} /* (23, 19, 3) {real, imag} */,
  {32'h400e6d33, 32'h3ea534e0} /* (23, 19, 2) {real, imag} */,
  {32'hbede8263, 32'h3fc6f924} /* (23, 19, 1) {real, imag} */,
  {32'hbe37d244, 32'h3efd3603} /* (23, 19, 0) {real, imag} */,
  {32'hbf82d915, 32'hbfeec0ae} /* (23, 18, 31) {real, imag} */,
  {32'hbfbc4d46, 32'hbdcb897b} /* (23, 18, 30) {real, imag} */,
  {32'h3f15e2fb, 32'hbfe0098b} /* (23, 18, 29) {real, imag} */,
  {32'h4034a3e6, 32'hc05475cc} /* (23, 18, 28) {real, imag} */,
  {32'h3f942711, 32'hbe9e4618} /* (23, 18, 27) {real, imag} */,
  {32'h3dda5bb8, 32'hbe38beae} /* (23, 18, 26) {real, imag} */,
  {32'hc094ad49, 32'h3f9d8b69} /* (23, 18, 25) {real, imag} */,
  {32'h3fd76763, 32'h3ff32086} /* (23, 18, 24) {real, imag} */,
  {32'hbfc97631, 32'hbf9a1d9a} /* (23, 18, 23) {real, imag} */,
  {32'hbf03f4e7, 32'hc03a84e0} /* (23, 18, 22) {real, imag} */,
  {32'h3f972402, 32'hbfb86e1a} /* (23, 18, 21) {real, imag} */,
  {32'hbf518f8e, 32'h3d92d2bb} /* (23, 18, 20) {real, imag} */,
  {32'h3c93484b, 32'hbee580ee} /* (23, 18, 19) {real, imag} */,
  {32'hbf2b9b10, 32'h3f578d83} /* (23, 18, 18) {real, imag} */,
  {32'hbf136f93, 32'h3d97011a} /* (23, 18, 17) {real, imag} */,
  {32'hbf1f3fcf, 32'hbf06afcf} /* (23, 18, 16) {real, imag} */,
  {32'h3ef34559, 32'h3fe6f128} /* (23, 18, 15) {real, imag} */,
  {32'hbc007ed6, 32'hbec4ae78} /* (23, 18, 14) {real, imag} */,
  {32'hbfce3d25, 32'h400a1228} /* (23, 18, 13) {real, imag} */,
  {32'hbf64e02a, 32'hbfbfef1e} /* (23, 18, 12) {real, imag} */,
  {32'hbfa6d6da, 32'h3fce79da} /* (23, 18, 11) {real, imag} */,
  {32'h3e8ebf59, 32'h3fe287ad} /* (23, 18, 10) {real, imag} */,
  {32'h3d99cb12, 32'h3fe8f128} /* (23, 18, 9) {real, imag} */,
  {32'hbf650c94, 32'h3de37e46} /* (23, 18, 8) {real, imag} */,
  {32'hc01c6af1, 32'h3fa4cff8} /* (23, 18, 7) {real, imag} */,
  {32'hbfa3646a, 32'h3ee8d012} /* (23, 18, 6) {real, imag} */,
  {32'hbd1603d0, 32'h4013fe01} /* (23, 18, 5) {real, imag} */,
  {32'h3fb6bef6, 32'hc064f356} /* (23, 18, 4) {real, imag} */,
  {32'hc012a127, 32'hbeadb345} /* (23, 18, 3) {real, imag} */,
  {32'hc011a5e8, 32'h3f245269} /* (23, 18, 2) {real, imag} */,
  {32'h3f741555, 32'hbf0be4ff} /* (23, 18, 1) {real, imag} */,
  {32'hbeea9cf2, 32'hc004fed9} /* (23, 18, 0) {real, imag} */,
  {32'hbfe283d9, 32'hbfc875c0} /* (23, 17, 31) {real, imag} */,
  {32'hbd89ec92, 32'hbf8f5892} /* (23, 17, 30) {real, imag} */,
  {32'h3e8dd83a, 32'h3f12e251} /* (23, 17, 29) {real, imag} */,
  {32'hbfe4bef2, 32'h3dd12ada} /* (23, 17, 28) {real, imag} */,
  {32'hbf7fb184, 32'h3ede322b} /* (23, 17, 27) {real, imag} */,
  {32'hc0060ed0, 32'hbf350f69} /* (23, 17, 26) {real, imag} */,
  {32'h3f26afb9, 32'h3f823536} /* (23, 17, 25) {real, imag} */,
  {32'h402337ff, 32'h3edf8d05} /* (23, 17, 24) {real, imag} */,
  {32'hbeef2bc2, 32'h3f1d48c7} /* (23, 17, 23) {real, imag} */,
  {32'h3fd34d31, 32'hc016a1d8} /* (23, 17, 22) {real, imag} */,
  {32'hbffdbccf, 32'hbf812175} /* (23, 17, 21) {real, imag} */,
  {32'hbf99db31, 32'h3fc0fc84} /* (23, 17, 20) {real, imag} */,
  {32'h403347ec, 32'h3ef96fa0} /* (23, 17, 19) {real, imag} */,
  {32'h3ff6e5fc, 32'h3fe29496} /* (23, 17, 18) {real, imag} */,
  {32'h4037670e, 32'hbf9a7dd8} /* (23, 17, 17) {real, imag} */,
  {32'hbf34e185, 32'h3f58dbee} /* (23, 17, 16) {real, imag} */,
  {32'h3f448e39, 32'h3efc8c3e} /* (23, 17, 15) {real, imag} */,
  {32'h3e720c25, 32'hbed06f19} /* (23, 17, 14) {real, imag} */,
  {32'h3fb841ed, 32'hc0081b81} /* (23, 17, 13) {real, imag} */,
  {32'hbee06e9d, 32'h3fe197c5} /* (23, 17, 12) {real, imag} */,
  {32'hbe727dd1, 32'hbf9afdb2} /* (23, 17, 11) {real, imag} */,
  {32'hc0127789, 32'h3f899f10} /* (23, 17, 10) {real, imag} */,
  {32'hbf6a77d2, 32'h3eef68d5} /* (23, 17, 9) {real, imag} */,
  {32'hbf5f69fa, 32'h3f380d28} /* (23, 17, 8) {real, imag} */,
  {32'hbfd99d06, 32'h3f86d7d7} /* (23, 17, 7) {real, imag} */,
  {32'h3f0e0cf8, 32'hbe77aa3e} /* (23, 17, 6) {real, imag} */,
  {32'h3f1cd9c8, 32'hc00f7abc} /* (23, 17, 5) {real, imag} */,
  {32'hbf85d4e2, 32'h3f633958} /* (23, 17, 4) {real, imag} */,
  {32'h3fe81a1d, 32'hbff2e3a1} /* (23, 17, 3) {real, imag} */,
  {32'h3e8353dc, 32'hbf8b1737} /* (23, 17, 2) {real, imag} */,
  {32'hbea9dc68, 32'h3ce411b3} /* (23, 17, 1) {real, imag} */,
  {32'h3f4fd711, 32'h3f0eb377} /* (23, 17, 0) {real, imag} */,
  {32'h3f9baa43, 32'hbfae4b03} /* (23, 16, 31) {real, imag} */,
  {32'hbf0747ed, 32'h3e050f39} /* (23, 16, 30) {real, imag} */,
  {32'hbf145187, 32'hbf12e541} /* (23, 16, 29) {real, imag} */,
  {32'h3f20ecd3, 32'h3fed8738} /* (23, 16, 28) {real, imag} */,
  {32'h3ff6c504, 32'h3fa62a73} /* (23, 16, 27) {real, imag} */,
  {32'h3e1347be, 32'hbfe69eca} /* (23, 16, 26) {real, imag} */,
  {32'h3f61a49f, 32'hbfbadf7b} /* (23, 16, 25) {real, imag} */,
  {32'h3f333cf4, 32'hbfe189e1} /* (23, 16, 24) {real, imag} */,
  {32'h3d17ecfb, 32'h3f650485} /* (23, 16, 23) {real, imag} */,
  {32'h3ebe0ca1, 32'hbf26beae} /* (23, 16, 22) {real, imag} */,
  {32'h3f049f35, 32'hc00f124e} /* (23, 16, 21) {real, imag} */,
  {32'hbf91d25c, 32'h3fd003be} /* (23, 16, 20) {real, imag} */,
  {32'hc023e0af, 32'h3f91a5a2} /* (23, 16, 19) {real, imag} */,
  {32'hbff91166, 32'h3eb0384f} /* (23, 16, 18) {real, imag} */,
  {32'h3fbb722c, 32'h3f288735} /* (23, 16, 17) {real, imag} */,
  {32'hbf4a02a2, 32'h400f3871} /* (23, 16, 16) {real, imag} */,
  {32'hbfc15ce8, 32'h3ffa315a} /* (23, 16, 15) {real, imag} */,
  {32'h3ee035d6, 32'h3e4e0af1} /* (23, 16, 14) {real, imag} */,
  {32'h3f9f6a95, 32'h3e2a7b91} /* (23, 16, 13) {real, imag} */,
  {32'hbfc307e4, 32'hc0663ee8} /* (23, 16, 12) {real, imag} */,
  {32'hbe39e4f3, 32'h3fbdf706} /* (23, 16, 11) {real, imag} */,
  {32'h3ed390b1, 32'hbfc008ed} /* (23, 16, 10) {real, imag} */,
  {32'h3f897879, 32'hbf8360ee} /* (23, 16, 9) {real, imag} */,
  {32'hbf48aa8c, 32'h3f3bc06f} /* (23, 16, 8) {real, imag} */,
  {32'hbe83bd65, 32'h3f3843c9} /* (23, 16, 7) {real, imag} */,
  {32'h3f87abd4, 32'hbf83d20a} /* (23, 16, 6) {real, imag} */,
  {32'h3e897f5d, 32'hbecf734f} /* (23, 16, 5) {real, imag} */,
  {32'h3e936e1d, 32'hbf96bc94} /* (23, 16, 4) {real, imag} */,
  {32'h3f131eca, 32'h3f533f3e} /* (23, 16, 3) {real, imag} */,
  {32'h3f4fb198, 32'h3e82b21e} /* (23, 16, 2) {real, imag} */,
  {32'hbefd2ba3, 32'hbf2bd271} /* (23, 16, 1) {real, imag} */,
  {32'h3f2c2349, 32'h40003d48} /* (23, 16, 0) {real, imag} */,
  {32'h3f933411, 32'h3f35f179} /* (23, 15, 31) {real, imag} */,
  {32'hbb7b9626, 32'h3fe9c1c9} /* (23, 15, 30) {real, imag} */,
  {32'hbe83da49, 32'hbf677a2a} /* (23, 15, 29) {real, imag} */,
  {32'h3fc2bc36, 32'h3f9c5e63} /* (23, 15, 28) {real, imag} */,
  {32'hbed00341, 32'h3e08ccb8} /* (23, 15, 27) {real, imag} */,
  {32'hbf90f2d4, 32'h401dd175} /* (23, 15, 26) {real, imag} */,
  {32'hbf106048, 32'hbf844713} /* (23, 15, 25) {real, imag} */,
  {32'hbe853cba, 32'hbf8e1c7a} /* (23, 15, 24) {real, imag} */,
  {32'h402d5388, 32'hbf014b09} /* (23, 15, 23) {real, imag} */,
  {32'h3ee53a32, 32'hbfdc70e7} /* (23, 15, 22) {real, imag} */,
  {32'hbfa241dd, 32'h406ba6ea} /* (23, 15, 21) {real, imag} */,
  {32'h3f66f9a3, 32'hc00ad2e1} /* (23, 15, 20) {real, imag} */,
  {32'hbe458612, 32'h3ff312ae} /* (23, 15, 19) {real, imag} */,
  {32'hbec6ee28, 32'h3f3379fb} /* (23, 15, 18) {real, imag} */,
  {32'hbf67ea5f, 32'hbf0bb671} /* (23, 15, 17) {real, imag} */,
  {32'hbfefcebf, 32'hbdc4afe3} /* (23, 15, 16) {real, imag} */,
  {32'hbfa152d3, 32'h3ff477ba} /* (23, 15, 15) {real, imag} */,
  {32'h3e936cb1, 32'hbf81db40} /* (23, 15, 14) {real, imag} */,
  {32'h3fa77384, 32'hbf71f340} /* (23, 15, 13) {real, imag} */,
  {32'h3f831d43, 32'hbf8d19e9} /* (23, 15, 12) {real, imag} */,
  {32'hbf875c67, 32'hbda1e611} /* (23, 15, 11) {real, imag} */,
  {32'h3f2b557c, 32'hbee73a98} /* (23, 15, 10) {real, imag} */,
  {32'h40192aa4, 32'hbf812629} /* (23, 15, 9) {real, imag} */,
  {32'h408fb545, 32'hbfee17ad} /* (23, 15, 8) {real, imag} */,
  {32'h3dcefd24, 32'hbf81fb34} /* (23, 15, 7) {real, imag} */,
  {32'hbfef754c, 32'h3fef14f8} /* (23, 15, 6) {real, imag} */,
  {32'h3eeeb2e6, 32'hc0199b7d} /* (23, 15, 5) {real, imag} */,
  {32'hbfd8d04c, 32'h3e0d5d9a} /* (23, 15, 4) {real, imag} */,
  {32'h3f9d04c0, 32'hbf2e8a4b} /* (23, 15, 3) {real, imag} */,
  {32'h3e4bcf0f, 32'h40052852} /* (23, 15, 2) {real, imag} */,
  {32'hbf82982b, 32'hbf94f5c4} /* (23, 15, 1) {real, imag} */,
  {32'h3ff80c0c, 32'h3e38f19e} /* (23, 15, 0) {real, imag} */,
  {32'hbf01e355, 32'hbf5aaeb5} /* (23, 14, 31) {real, imag} */,
  {32'hbf8b290b, 32'h3fd752bd} /* (23, 14, 30) {real, imag} */,
  {32'h3fbc3c51, 32'hbfa3a288} /* (23, 14, 29) {real, imag} */,
  {32'hbf9817fe, 32'hbf99e51b} /* (23, 14, 28) {real, imag} */,
  {32'h3fa0e388, 32'hc042c7fa} /* (23, 14, 27) {real, imag} */,
  {32'h3fc2e92a, 32'hbf241456} /* (23, 14, 26) {real, imag} */,
  {32'hc00d55ee, 32'hbdf1184d} /* (23, 14, 25) {real, imag} */,
  {32'hc037dded, 32'h40107b4e} /* (23, 14, 24) {real, imag} */,
  {32'hbf20ab09, 32'h3fe0f14c} /* (23, 14, 23) {real, imag} */,
  {32'h3fdaaeca, 32'h3fa3ab88} /* (23, 14, 22) {real, imag} */,
  {32'hbdf01ea6, 32'h3fe0ec05} /* (23, 14, 21) {real, imag} */,
  {32'h3fdc6f6c, 32'hbe74bb0d} /* (23, 14, 20) {real, imag} */,
  {32'h3f94a5bb, 32'h3fd103f5} /* (23, 14, 19) {real, imag} */,
  {32'h3f7c2137, 32'hbf8a409f} /* (23, 14, 18) {real, imag} */,
  {32'h3f52fbda, 32'h3fb913d5} /* (23, 14, 17) {real, imag} */,
  {32'hbf112645, 32'h3f5982c2} /* (23, 14, 16) {real, imag} */,
  {32'hbfd805fa, 32'hbf7535be} /* (23, 14, 15) {real, imag} */,
  {32'h3fa39bd7, 32'h3e85394b} /* (23, 14, 14) {real, imag} */,
  {32'hbf3ac754, 32'h3f6ae710} /* (23, 14, 13) {real, imag} */,
  {32'h401c4953, 32'hc091bef0} /* (23, 14, 12) {real, imag} */,
  {32'h3cfcac86, 32'h4018e331} /* (23, 14, 11) {real, imag} */,
  {32'h402e474a, 32'hbf4517de} /* (23, 14, 10) {real, imag} */,
  {32'h3ee6e345, 32'h3e18691d} /* (23, 14, 9) {real, imag} */,
  {32'hbe29b724, 32'hbee9d7ce} /* (23, 14, 8) {real, imag} */,
  {32'h3f3d0be8, 32'hbf50db64} /* (23, 14, 7) {real, imag} */,
  {32'h3eff622e, 32'h3f8b55ed} /* (23, 14, 6) {real, imag} */,
  {32'hbff0cf1b, 32'h3e4709bd} /* (23, 14, 5) {real, imag} */,
  {32'hbf7853aa, 32'h3fad3737} /* (23, 14, 4) {real, imag} */,
  {32'hbe81080f, 32'hbf6613e6} /* (23, 14, 3) {real, imag} */,
  {32'h3f8b08eb, 32'h400f0ab3} /* (23, 14, 2) {real, imag} */,
  {32'h3ef629c7, 32'hbfcced10} /* (23, 14, 1) {real, imag} */,
  {32'h3e965097, 32'h3f293d1e} /* (23, 14, 0) {real, imag} */,
  {32'h3f1135f0, 32'h3ff3f4ca} /* (23, 13, 31) {real, imag} */,
  {32'hbe847887, 32'h3f658aa3} /* (23, 13, 30) {real, imag} */,
  {32'h3f770754, 32'hbff55952} /* (23, 13, 29) {real, imag} */,
  {32'hbfa2ea40, 32'h4062c51a} /* (23, 13, 28) {real, imag} */,
  {32'hbef31227, 32'hbfc6c667} /* (23, 13, 27) {real, imag} */,
  {32'hbffc42e8, 32'h3e8a6e4d} /* (23, 13, 26) {real, imag} */,
  {32'hbebd1eb5, 32'hbdffdf45} /* (23, 13, 25) {real, imag} */,
  {32'hbe495688, 32'h3f342a06} /* (23, 13, 24) {real, imag} */,
  {32'h3f5d6560, 32'h3f10ce59} /* (23, 13, 23) {real, imag} */,
  {32'hc06a8826, 32'hbe95dff8} /* (23, 13, 22) {real, imag} */,
  {32'hbf4dc1ee, 32'h404839fd} /* (23, 13, 21) {real, imag} */,
  {32'hbf37adef, 32'hbf2c45e3} /* (23, 13, 20) {real, imag} */,
  {32'h401201de, 32'hbe01d939} /* (23, 13, 19) {real, imag} */,
  {32'h3f7350ee, 32'hbfdc2476} /* (23, 13, 18) {real, imag} */,
  {32'h3f9cd22c, 32'hc0541a71} /* (23, 13, 17) {real, imag} */,
  {32'h3e069dbe, 32'h3e8dd6f8} /* (23, 13, 16) {real, imag} */,
  {32'hc001794c, 32'h3fe2599e} /* (23, 13, 15) {real, imag} */,
  {32'h3ff1c125, 32'h3f8a7348} /* (23, 13, 14) {real, imag} */,
  {32'h3f9da7a6, 32'h40053a7f} /* (23, 13, 13) {real, imag} */,
  {32'h3fd1425c, 32'h40486079} /* (23, 13, 12) {real, imag} */,
  {32'hc0226f8d, 32'hbec361e5} /* (23, 13, 11) {real, imag} */,
  {32'hc0085bfa, 32'hbeccc82d} /* (23, 13, 10) {real, imag} */,
  {32'hbf150990, 32'h3f8eba21} /* (23, 13, 9) {real, imag} */,
  {32'h4049783f, 32'hbfc8bc3c} /* (23, 13, 8) {real, imag} */,
  {32'h3fc0f1fd, 32'hbf3ae3da} /* (23, 13, 7) {real, imag} */,
  {32'hbd8a024c, 32'hbf35734a} /* (23, 13, 6) {real, imag} */,
  {32'h3f770f94, 32'hc0179f45} /* (23, 13, 5) {real, imag} */,
  {32'hc001f283, 32'hbed7e745} /* (23, 13, 4) {real, imag} */,
  {32'h3f634d83, 32'h3f871686} /* (23, 13, 3) {real, imag} */,
  {32'hbf60613b, 32'hbe8714a0} /* (23, 13, 2) {real, imag} */,
  {32'hbc5d6502, 32'h3f104937} /* (23, 13, 1) {real, imag} */,
  {32'hc01293d0, 32'h408bfbc8} /* (23, 13, 0) {real, imag} */,
  {32'h3eb53e03, 32'h3fdb28fc} /* (23, 12, 31) {real, imag} */,
  {32'hbfcf89f2, 32'h3f62c604} /* (23, 12, 30) {real, imag} */,
  {32'hc00d3275, 32'h4014762b} /* (23, 12, 29) {real, imag} */,
  {32'h3f70f6f9, 32'hbf9e492c} /* (23, 12, 28) {real, imag} */,
  {32'h3ec15963, 32'hbd831297} /* (23, 12, 27) {real, imag} */,
  {32'h3fad766c, 32'h402c1507} /* (23, 12, 26) {real, imag} */,
  {32'hbfd736b5, 32'h3f2f0edd} /* (23, 12, 25) {real, imag} */,
  {32'h3ffd944f, 32'h3fa33b5c} /* (23, 12, 24) {real, imag} */,
  {32'hc005c47b, 32'h3fbfb2e8} /* (23, 12, 23) {real, imag} */,
  {32'h3ff6e304, 32'h3fba437b} /* (23, 12, 22) {real, imag} */,
  {32'hc02e219a, 32'hc043f163} /* (23, 12, 21) {real, imag} */,
  {32'hbf1f698b, 32'hbfb6c1b5} /* (23, 12, 20) {real, imag} */,
  {32'h3fe50a2b, 32'hbea716ba} /* (23, 12, 19) {real, imag} */,
  {32'hbf345e53, 32'hc0154866} /* (23, 12, 18) {real, imag} */,
  {32'hbf486a46, 32'hbf3efdff} /* (23, 12, 17) {real, imag} */,
  {32'hbed6c996, 32'hbf9e0d4d} /* (23, 12, 16) {real, imag} */,
  {32'h3f134d5c, 32'hbf43d92b} /* (23, 12, 15) {real, imag} */,
  {32'h3f8bcc7d, 32'h3ffc23e2} /* (23, 12, 14) {real, imag} */,
  {32'h3f6047ea, 32'hc0474382} /* (23, 12, 13) {real, imag} */,
  {32'h3fe533ea, 32'h40a84dfd} /* (23, 12, 12) {real, imag} */,
  {32'hbff39a91, 32'h3c98e734} /* (23, 12, 11) {real, imag} */,
  {32'hbf3b770d, 32'hbf3f78f0} /* (23, 12, 10) {real, imag} */,
  {32'hc0862b8b, 32'hbed3e5ae} /* (23, 12, 9) {real, imag} */,
  {32'hbfef1bee, 32'h3e46e92e} /* (23, 12, 8) {real, imag} */,
  {32'h3f276018, 32'hc0802e2a} /* (23, 12, 7) {real, imag} */,
  {32'h3ebb17a8, 32'h3ed15870} /* (23, 12, 6) {real, imag} */,
  {32'hc0081d20, 32'h3e909158} /* (23, 12, 5) {real, imag} */,
  {32'h3f9727c1, 32'hbf7f8688} /* (23, 12, 4) {real, imag} */,
  {32'h3fb802c1, 32'h3f5f5761} /* (23, 12, 3) {real, imag} */,
  {32'h3fba32ae, 32'hbf46b4c0} /* (23, 12, 2) {real, imag} */,
  {32'h3f21df2b, 32'hbeb6a106} /* (23, 12, 1) {real, imag} */,
  {32'h3fb3e015, 32'hbe73b4d7} /* (23, 12, 0) {real, imag} */,
  {32'h3f056e42, 32'h3ebc14bd} /* (23, 11, 31) {real, imag} */,
  {32'h3f922314, 32'hbfcc5df7} /* (23, 11, 30) {real, imag} */,
  {32'hbdb7f06d, 32'h3f0dc19f} /* (23, 11, 29) {real, imag} */,
  {32'hc02c7a66, 32'h4001918a} /* (23, 11, 28) {real, imag} */,
  {32'h405d7357, 32'hbeef0dd5} /* (23, 11, 27) {real, imag} */,
  {32'h3f054095, 32'h4057c841} /* (23, 11, 26) {real, imag} */,
  {32'h3f1fb6e4, 32'h3f7b9aa6} /* (23, 11, 25) {real, imag} */,
  {32'h3eeb6b80, 32'hbfc6f8a8} /* (23, 11, 24) {real, imag} */,
  {32'hc0929feb, 32'hbe85deec} /* (23, 11, 23) {real, imag} */,
  {32'hbf86dd36, 32'hbffc5d92} /* (23, 11, 22) {real, imag} */,
  {32'h40123b9e, 32'hbfd244bf} /* (23, 11, 21) {real, imag} */,
  {32'h3fe65ba9, 32'hbf6d6edc} /* (23, 11, 20) {real, imag} */,
  {32'hbf1a87e2, 32'hbe217027} /* (23, 11, 19) {real, imag} */,
  {32'hbf6f4f54, 32'h3e50d0e5} /* (23, 11, 18) {real, imag} */,
  {32'h3cb48e7b, 32'h3f4a7ee3} /* (23, 11, 17) {real, imag} */,
  {32'h3cf91bcf, 32'h3eea490b} /* (23, 11, 16) {real, imag} */,
  {32'h3f4de953, 32'hbfa953b5} /* (23, 11, 15) {real, imag} */,
  {32'h4060fdfe, 32'h3f7af6bf} /* (23, 11, 14) {real, imag} */,
  {32'hbf75b414, 32'hc039e9a6} /* (23, 11, 13) {real, imag} */,
  {32'hbfcc4ba3, 32'hbf0f1d18} /* (23, 11, 12) {real, imag} */,
  {32'hbf8aa64e, 32'hbf3ccea3} /* (23, 11, 11) {real, imag} */,
  {32'hbd507cf4, 32'hbfce7ebb} /* (23, 11, 10) {real, imag} */,
  {32'hbf06c4af, 32'h3edfd13b} /* (23, 11, 9) {real, imag} */,
  {32'h3c9b4b9a, 32'hbf8e54c1} /* (23, 11, 8) {real, imag} */,
  {32'h404167fa, 32'hbf9fd417} /* (23, 11, 7) {real, imag} */,
  {32'h4085a8d5, 32'h401e89a9} /* (23, 11, 6) {real, imag} */,
  {32'hbf47814f, 32'hc003c81d} /* (23, 11, 5) {real, imag} */,
  {32'hbf47b9d8, 32'h403567a6} /* (23, 11, 4) {real, imag} */,
  {32'hbf288060, 32'hc0156c57} /* (23, 11, 3) {real, imag} */,
  {32'h3f982105, 32'h40139c1b} /* (23, 11, 2) {real, imag} */,
  {32'hbfb7d2c6, 32'hbf61331a} /* (23, 11, 1) {real, imag} */,
  {32'h3f8249bb, 32'hbfaf3e72} /* (23, 11, 0) {real, imag} */,
  {32'h3fd115e8, 32'h3fca4872} /* (23, 10, 31) {real, imag} */,
  {32'h3e864133, 32'hbe8eacca} /* (23, 10, 30) {real, imag} */,
  {32'h3ffb056d, 32'h3d508c0e} /* (23, 10, 29) {real, imag} */,
  {32'h3f021bcb, 32'h40886396} /* (23, 10, 28) {real, imag} */,
  {32'h3e2db7ad, 32'hbfa151f6} /* (23, 10, 27) {real, imag} */,
  {32'h3f513ac4, 32'hc051335a} /* (23, 10, 26) {real, imag} */,
  {32'h3f917b22, 32'h3ea27a04} /* (23, 10, 25) {real, imag} */,
  {32'hbf7ea01c, 32'h3ec1c92f} /* (23, 10, 24) {real, imag} */,
  {32'h3f181b4b, 32'hc025618a} /* (23, 10, 23) {real, imag} */,
  {32'h3eff2056, 32'h400bdfe1} /* (23, 10, 22) {real, imag} */,
  {32'h40295632, 32'hbfec0842} /* (23, 10, 21) {real, imag} */,
  {32'h3fe71f2f, 32'h3fa9801f} /* (23, 10, 20) {real, imag} */,
  {32'hbf8f1d62, 32'h4085cb11} /* (23, 10, 19) {real, imag} */,
  {32'h3db96266, 32'h3f9485e6} /* (23, 10, 18) {real, imag} */,
  {32'hbf0d57ab, 32'hbf07832b} /* (23, 10, 17) {real, imag} */,
  {32'h3c477ec5, 32'hc004ce44} /* (23, 10, 16) {real, imag} */,
  {32'h3ca755d4, 32'h3c2800b5} /* (23, 10, 15) {real, imag} */,
  {32'hbf798d14, 32'hbec39c5c} /* (23, 10, 14) {real, imag} */,
  {32'hbe7adc2d, 32'h401870e0} /* (23, 10, 13) {real, imag} */,
  {32'h4078ad70, 32'h3ffa8b84} /* (23, 10, 12) {real, imag} */,
  {32'hbf8e7b29, 32'h3e04e27b} /* (23, 10, 11) {real, imag} */,
  {32'h3f68c817, 32'h3f5f94a3} /* (23, 10, 10) {real, imag} */,
  {32'h3f3cd5f9, 32'h400120f6} /* (23, 10, 9) {real, imag} */,
  {32'hc0022602, 32'hbfc0e573} /* (23, 10, 8) {real, imag} */,
  {32'hc08a9ffe, 32'hbffc41a8} /* (23, 10, 7) {real, imag} */,
  {32'h401d3484, 32'h3e06a0d9} /* (23, 10, 6) {real, imag} */,
  {32'h3f0fed89, 32'hbfba361f} /* (23, 10, 5) {real, imag} */,
  {32'h3e8e1b11, 32'hc02c7ebc} /* (23, 10, 4) {real, imag} */,
  {32'hbfa03846, 32'hbf3dd51a} /* (23, 10, 3) {real, imag} */,
  {32'hbe8de840, 32'h408188e9} /* (23, 10, 2) {real, imag} */,
  {32'hbfdeccc6, 32'hc038f664} /* (23, 10, 1) {real, imag} */,
  {32'h3f3049e5, 32'hbe1f653b} /* (23, 10, 0) {real, imag} */,
  {32'h3f4cea85, 32'hc0262cfa} /* (23, 9, 31) {real, imag} */,
  {32'hbf42dd17, 32'h3f00dd19} /* (23, 9, 30) {real, imag} */,
  {32'h3eab0d76, 32'h3f73ccd0} /* (23, 9, 29) {real, imag} */,
  {32'hbfb22c5c, 32'hc089fff7} /* (23, 9, 28) {real, imag} */,
  {32'h3ff9a90c, 32'hbfa7a63a} /* (23, 9, 27) {real, imag} */,
  {32'h40058b56, 32'hbf3bcbb7} /* (23, 9, 26) {real, imag} */,
  {32'h3e1b6633, 32'h3f736339} /* (23, 9, 25) {real, imag} */,
  {32'h40c6b775, 32'h3f490c65} /* (23, 9, 24) {real, imag} */,
  {32'hc0145a95, 32'hbee591cc} /* (23, 9, 23) {real, imag} */,
  {32'hbfeb0828, 32'hbff9a610} /* (23, 9, 22) {real, imag} */,
  {32'hbfbb8e34, 32'hbf8b1ffb} /* (23, 9, 21) {real, imag} */,
  {32'hbffc20e7, 32'hbe80ae7c} /* (23, 9, 20) {real, imag} */,
  {32'h40135703, 32'h3f99433a} /* (23, 9, 19) {real, imag} */,
  {32'hbfb921ce, 32'hbef22b73} /* (23, 9, 18) {real, imag} */,
  {32'hbf5e7444, 32'h3f1a9683} /* (23, 9, 17) {real, imag} */,
  {32'h3ee325a7, 32'hbeb4b580} /* (23, 9, 16) {real, imag} */,
  {32'h4004fea7, 32'h3eba27b7} /* (23, 9, 15) {real, imag} */,
  {32'hbfb2f7ec, 32'hbef99571} /* (23, 9, 14) {real, imag} */,
  {32'hc00fc5a7, 32'hbf95cb6f} /* (23, 9, 13) {real, imag} */,
  {32'h3fc52a9f, 32'h3fe047e4} /* (23, 9, 12) {real, imag} */,
  {32'hc0149c67, 32'hbf61386c} /* (23, 9, 11) {real, imag} */,
  {32'hbf8d7c44, 32'h3f93dc16} /* (23, 9, 10) {real, imag} */,
  {32'hbfb905eb, 32'hbde0cb43} /* (23, 9, 9) {real, imag} */,
  {32'hbf42aa57, 32'h3f2d7bd5} /* (23, 9, 8) {real, imag} */,
  {32'hbffbe287, 32'hbfb7d9cc} /* (23, 9, 7) {real, imag} */,
  {32'h3f8874ee, 32'hc021311a} /* (23, 9, 6) {real, imag} */,
  {32'hbf9f90e4, 32'h3cdecbab} /* (23, 9, 5) {real, imag} */,
  {32'h3f987b94, 32'hbf8a100d} /* (23, 9, 4) {real, imag} */,
  {32'hbe89b1f7, 32'h3f74f951} /* (23, 9, 3) {real, imag} */,
  {32'h3f8096cb, 32'h3eee0c02} /* (23, 9, 2) {real, imag} */,
  {32'hc041209f, 32'h409ff4f2} /* (23, 9, 1) {real, imag} */,
  {32'h3f1eb59a, 32'hbef9f15d} /* (23, 9, 0) {real, imag} */,
  {32'h3f5aea9f, 32'h3ed4987a} /* (23, 8, 31) {real, imag} */,
  {32'hbeea31c8, 32'hc01c2275} /* (23, 8, 30) {real, imag} */,
  {32'hbf0b37d3, 32'h3f30f12f} /* (23, 8, 29) {real, imag} */,
  {32'h405d6cd9, 32'h3f55921d} /* (23, 8, 28) {real, imag} */,
  {32'h3ec28791, 32'hc04089b7} /* (23, 8, 27) {real, imag} */,
  {32'hbe9cd8b4, 32'hbe7cd07b} /* (23, 8, 26) {real, imag} */,
  {32'hbe9e522a, 32'hbf91292e} /* (23, 8, 25) {real, imag} */,
  {32'hbfcdc65f, 32'hc01712b5} /* (23, 8, 24) {real, imag} */,
  {32'h3fab9d3e, 32'hbfd96774} /* (23, 8, 23) {real, imag} */,
  {32'h40437c57, 32'h3ec45884} /* (23, 8, 22) {real, imag} */,
  {32'hbd3efb09, 32'h4062cbbe} /* (23, 8, 21) {real, imag} */,
  {32'hbd220ae9, 32'h40574af5} /* (23, 8, 20) {real, imag} */,
  {32'h3fe0590e, 32'hc082850f} /* (23, 8, 19) {real, imag} */,
  {32'h3fd88c23, 32'hbf6bb7b5} /* (23, 8, 18) {real, imag} */,
  {32'hbf42a106, 32'h401b22cc} /* (23, 8, 17) {real, imag} */,
  {32'hbf1b962a, 32'hc016872c} /* (23, 8, 16) {real, imag} */,
  {32'hbf295758, 32'h3ca484f6} /* (23, 8, 15) {real, imag} */,
  {32'h4048f626, 32'h3f05f913} /* (23, 8, 14) {real, imag} */,
  {32'h3f8b7dfb, 32'hbf948bee} /* (23, 8, 13) {real, imag} */,
  {32'hbe5bb8cd, 32'hc03d69b2} /* (23, 8, 12) {real, imag} */,
  {32'h3e1c3da9, 32'h3f1fa28c} /* (23, 8, 11) {real, imag} */,
  {32'h3ed70fd4, 32'h401856b6} /* (23, 8, 10) {real, imag} */,
  {32'hbf85efbb, 32'h3f49239d} /* (23, 8, 9) {real, imag} */,
  {32'h40367a95, 32'h3f1f855b} /* (23, 8, 8) {real, imag} */,
  {32'hbfd68c5a, 32'hc019493f} /* (23, 8, 7) {real, imag} */,
  {32'hbfea674e, 32'h3ffceb00} /* (23, 8, 6) {real, imag} */,
  {32'h3fd11c06, 32'h4076648b} /* (23, 8, 5) {real, imag} */,
  {32'hbf84fdaa, 32'hbfe8a16f} /* (23, 8, 4) {real, imag} */,
  {32'hbf7f2d6f, 32'h3f9094ee} /* (23, 8, 3) {real, imag} */,
  {32'hbfe24b2f, 32'hbfac7aef} /* (23, 8, 2) {real, imag} */,
  {32'h3dd85674, 32'hc029c27e} /* (23, 8, 1) {real, imag} */,
  {32'hbf7a4474, 32'h4040d217} /* (23, 8, 0) {real, imag} */,
  {32'h3fb713a0, 32'hc0a1ee17} /* (23, 7, 31) {real, imag} */,
  {32'h3f0877c1, 32'h3fb91dd1} /* (23, 7, 30) {real, imag} */,
  {32'h3fd8e17f, 32'h3fe8727b} /* (23, 7, 29) {real, imag} */,
  {32'h3f9e123a, 32'h3f923749} /* (23, 7, 28) {real, imag} */,
  {32'h40908d43, 32'h40c27e3e} /* (23, 7, 27) {real, imag} */,
  {32'hc03d0d7f, 32'hbe1b07a4} /* (23, 7, 26) {real, imag} */,
  {32'h3f528d4f, 32'hbfc15caa} /* (23, 7, 25) {real, imag} */,
  {32'h400853da, 32'hbff04667} /* (23, 7, 24) {real, imag} */,
  {32'hbfe84857, 32'hbfd512fc} /* (23, 7, 23) {real, imag} */,
  {32'hc05aca0d, 32'hc00f3a38} /* (23, 7, 22) {real, imag} */,
  {32'hbff649d3, 32'h3edd740f} /* (23, 7, 21) {real, imag} */,
  {32'hbf5205ad, 32'h3f27ec5b} /* (23, 7, 20) {real, imag} */,
  {32'h3ec82e1b, 32'h3fca3be6} /* (23, 7, 19) {real, imag} */,
  {32'h3efae09f, 32'h3fb4ea30} /* (23, 7, 18) {real, imag} */,
  {32'hbf874103, 32'hbebafe79} /* (23, 7, 17) {real, imag} */,
  {32'h3f707ebb, 32'h3face86e} /* (23, 7, 16) {real, imag} */,
  {32'h4006f098, 32'hbfc29936} /* (23, 7, 15) {real, imag} */,
  {32'h3fd79863, 32'hbf22c321} /* (23, 7, 14) {real, imag} */,
  {32'hbfc67561, 32'h403834b8} /* (23, 7, 13) {real, imag} */,
  {32'hbc8f7591, 32'hbdecb28e} /* (23, 7, 12) {real, imag} */,
  {32'hc0188327, 32'h402ad367} /* (23, 7, 11) {real, imag} */,
  {32'hc02bcd7e, 32'hc049a94a} /* (23, 7, 10) {real, imag} */,
  {32'hc001eeb9, 32'hbeadd4fd} /* (23, 7, 9) {real, imag} */,
  {32'h3fe3a70e, 32'h3f4a54fd} /* (23, 7, 8) {real, imag} */,
  {32'hbf662aa7, 32'hbf24eb19} /* (23, 7, 7) {real, imag} */,
  {32'hc041fd3a, 32'hbfa65901} /* (23, 7, 6) {real, imag} */,
  {32'hbfaf3161, 32'hc035d11a} /* (23, 7, 5) {real, imag} */,
  {32'h3f742777, 32'hbf87ed14} /* (23, 7, 4) {real, imag} */,
  {32'hbd97f52c, 32'hbe541a1f} /* (23, 7, 3) {real, imag} */,
  {32'h3e6e2442, 32'h40589349} /* (23, 7, 2) {real, imag} */,
  {32'h3fed628e, 32'h3f9bba7c} /* (23, 7, 1) {real, imag} */,
  {32'h3f6e7c90, 32'h3f16876e} /* (23, 7, 0) {real, imag} */,
  {32'h403f89fc, 32'hbf29586e} /* (23, 6, 31) {real, imag} */,
  {32'hbf834d4a, 32'hbea9387b} /* (23, 6, 30) {real, imag} */,
  {32'hc0463b53, 32'h3ea7aff5} /* (23, 6, 29) {real, imag} */,
  {32'h3fffae94, 32'hc042ea0d} /* (23, 6, 28) {real, imag} */,
  {32'hc06a8daa, 32'hbf1cbdf5} /* (23, 6, 27) {real, imag} */,
  {32'hc00de6a8, 32'hc0131a71} /* (23, 6, 26) {real, imag} */,
  {32'h3f100527, 32'hc0105218} /* (23, 6, 25) {real, imag} */,
  {32'hbf16c3fa, 32'h4032b249} /* (23, 6, 24) {real, imag} */,
  {32'h3fb77d9a, 32'hbc5744c2} /* (23, 6, 23) {real, imag} */,
  {32'hc06d250d, 32'h40a3f5cb} /* (23, 6, 22) {real, imag} */,
  {32'h3f3f7223, 32'hc00d4ab6} /* (23, 6, 21) {real, imag} */,
  {32'h3fbaceb2, 32'hbf9ddd93} /* (23, 6, 20) {real, imag} */,
  {32'hbf0e2e2d, 32'hbe5ac6fa} /* (23, 6, 19) {real, imag} */,
  {32'hbeb1b596, 32'h3f5c1aaa} /* (23, 6, 18) {real, imag} */,
  {32'h40819090, 32'h3fdd5e2b} /* (23, 6, 17) {real, imag} */,
  {32'hbf92ae04, 32'h3fd1604a} /* (23, 6, 16) {real, imag} */,
  {32'hbfe40a5c, 32'hbe51ebab} /* (23, 6, 15) {real, imag} */,
  {32'hc02de3dd, 32'h40105eb9} /* (23, 6, 14) {real, imag} */,
  {32'hbf48a343, 32'h3f583406} /* (23, 6, 13) {real, imag} */,
  {32'hbfda9ead, 32'h4044332f} /* (23, 6, 12) {real, imag} */,
  {32'h3e97a5bf, 32'hc081cc98} /* (23, 6, 11) {real, imag} */,
  {32'hbdf9e090, 32'h400dadb4} /* (23, 6, 10) {real, imag} */,
  {32'h402e7d63, 32'hbff530fd} /* (23, 6, 9) {real, imag} */,
  {32'hbece8a1b, 32'hbfba09f3} /* (23, 6, 8) {real, imag} */,
  {32'h3f9ca35a, 32'h3d0752c0} /* (23, 6, 7) {real, imag} */,
  {32'h3f08b514, 32'h3f919d0d} /* (23, 6, 6) {real, imag} */,
  {32'hbfb7a40d, 32'hbf28a956} /* (23, 6, 5) {real, imag} */,
  {32'h401a6caa, 32'hbe4f9e07} /* (23, 6, 4) {real, imag} */,
  {32'h400d0a80, 32'h40d78fc9} /* (23, 6, 3) {real, imag} */,
  {32'h3fee28c9, 32'h3f557e14} /* (23, 6, 2) {real, imag} */,
  {32'hc02a1e1a, 32'h403d1472} /* (23, 6, 1) {real, imag} */,
  {32'hc0098b8a, 32'h3ebb9601} /* (23, 6, 0) {real, imag} */,
  {32'hbf9de27b, 32'h3fc31c7a} /* (23, 5, 31) {real, imag} */,
  {32'h3ffa48b2, 32'hc0035df3} /* (23, 5, 30) {real, imag} */,
  {32'hc048f778, 32'hbfc94b3c} /* (23, 5, 29) {real, imag} */,
  {32'hbec02ca0, 32'h3f4dc756} /* (23, 5, 28) {real, imag} */,
  {32'h3cd5fa22, 32'hc01bbe9c} /* (23, 5, 27) {real, imag} */,
  {32'hbfc12cd1, 32'hc0442ec8} /* (23, 5, 26) {real, imag} */,
  {32'h4014d275, 32'hbe31bc41} /* (23, 5, 25) {real, imag} */,
  {32'h4053f79e, 32'hc03ffdea} /* (23, 5, 24) {real, imag} */,
  {32'h4035f7bb, 32'hc0540a45} /* (23, 5, 23) {real, imag} */,
  {32'h3fd5d054, 32'h407bde98} /* (23, 5, 22) {real, imag} */,
  {32'hbff186a7, 32'h3f0e3c3b} /* (23, 5, 21) {real, imag} */,
  {32'h3f8f2c34, 32'h3edcf1bb} /* (23, 5, 20) {real, imag} */,
  {32'hbf1195b1, 32'h3f98c398} /* (23, 5, 19) {real, imag} */,
  {32'hbff3e4c3, 32'h40130e1d} /* (23, 5, 18) {real, imag} */,
  {32'hbd938016, 32'hbe36bf1d} /* (23, 5, 17) {real, imag} */,
  {32'hbfa470bf, 32'hbf9b8a6f} /* (23, 5, 16) {real, imag} */,
  {32'h3f8410d5, 32'h3fd8356c} /* (23, 5, 15) {real, imag} */,
  {32'h3e18e900, 32'h3f70cfa7} /* (23, 5, 14) {real, imag} */,
  {32'h3dcbfa2b, 32'hbf82425d} /* (23, 5, 13) {real, imag} */,
  {32'hc07eacf1, 32'h3d8144e1} /* (23, 5, 12) {real, imag} */,
  {32'h3e9905ed, 32'hc01b70c5} /* (23, 5, 11) {real, imag} */,
  {32'h3d6dd515, 32'hc0879e88} /* (23, 5, 10) {real, imag} */,
  {32'hbfbbcb26, 32'hc0747a1f} /* (23, 5, 9) {real, imag} */,
  {32'hbf73bd75, 32'h4030d6dd} /* (23, 5, 8) {real, imag} */,
  {32'h400dce51, 32'h4083d6fc} /* (23, 5, 7) {real, imag} */,
  {32'hc00d0095, 32'hc04e5e9a} /* (23, 5, 6) {real, imag} */,
  {32'h3f911d87, 32'hbe87af9a} /* (23, 5, 5) {real, imag} */,
  {32'h3f2f2128, 32'h3fd9c576} /* (23, 5, 4) {real, imag} */,
  {32'h4028f603, 32'h3f87f3bc} /* (23, 5, 3) {real, imag} */,
  {32'hc0134480, 32'hbff8d91e} /* (23, 5, 2) {real, imag} */,
  {32'h4014e92a, 32'h4083a0a6} /* (23, 5, 1) {real, imag} */,
  {32'h3f676323, 32'hbfaf8a11} /* (23, 5, 0) {real, imag} */,
  {32'h3ff9d852, 32'hc05b0d7a} /* (23, 4, 31) {real, imag} */,
  {32'hbfd64f74, 32'h404acf98} /* (23, 4, 30) {real, imag} */,
  {32'hc00fbf40, 32'hc0152154} /* (23, 4, 29) {real, imag} */,
  {32'hbfac0f31, 32'hbeb87404} /* (23, 4, 28) {real, imag} */,
  {32'hbf9cbc63, 32'h3ffc5bbb} /* (23, 4, 27) {real, imag} */,
  {32'h3fb1680f, 32'hbf6e504b} /* (23, 4, 26) {real, imag} */,
  {32'h3f5e2984, 32'h3fbf2f29} /* (23, 4, 25) {real, imag} */,
  {32'hc0c66462, 32'h3fe44d79} /* (23, 4, 24) {real, imag} */,
  {32'hbfe34b7d, 32'hbf4054e2} /* (23, 4, 23) {real, imag} */,
  {32'hbf8c48f6, 32'h3fe888de} /* (23, 4, 22) {real, imag} */,
  {32'hbf683337, 32'hbf9d763e} /* (23, 4, 21) {real, imag} */,
  {32'hbeb72828, 32'h3f0a0cbf} /* (23, 4, 20) {real, imag} */,
  {32'hbfb8d9d0, 32'h3fdce455} /* (23, 4, 19) {real, imag} */,
  {32'h3fe4e549, 32'hc0512365} /* (23, 4, 18) {real, imag} */,
  {32'h3ea556e7, 32'h3fbbf704} /* (23, 4, 17) {real, imag} */,
  {32'h3fb58293, 32'hbfc95495} /* (23, 4, 16) {real, imag} */,
  {32'hbfa3929b, 32'h3e513591} /* (23, 4, 15) {real, imag} */,
  {32'hbf773e55, 32'hc0090f2e} /* (23, 4, 14) {real, imag} */,
  {32'hbfde4275, 32'hbff40104} /* (23, 4, 13) {real, imag} */,
  {32'h404b34b5, 32'hc0185780} /* (23, 4, 12) {real, imag} */,
  {32'h3e08f994, 32'h3fb637be} /* (23, 4, 11) {real, imag} */,
  {32'h3fef7dc5, 32'hbee6c5dd} /* (23, 4, 10) {real, imag} */,
  {32'h3fd440ce, 32'hbfd15940} /* (23, 4, 9) {real, imag} */,
  {32'h405b6b6c, 32'h40012418} /* (23, 4, 8) {real, imag} */,
  {32'hbf46b170, 32'h3ffc6676} /* (23, 4, 7) {real, imag} */,
  {32'h4042c4d5, 32'h4060c04e} /* (23, 4, 6) {real, imag} */,
  {32'h4020bb48, 32'h401d47e5} /* (23, 4, 5) {real, imag} */,
  {32'h400956fc, 32'h3e624fd6} /* (23, 4, 4) {real, imag} */,
  {32'hbf05f2ae, 32'hc01c08ec} /* (23, 4, 3) {real, imag} */,
  {32'hbfd258e9, 32'hbf8d221d} /* (23, 4, 2) {real, imag} */,
  {32'h3f9efcdf, 32'h3fe404c9} /* (23, 4, 1) {real, imag} */,
  {32'h3f7446d4, 32'h405a4495} /* (23, 4, 0) {real, imag} */,
  {32'hbce755bc, 32'h4094a05e} /* (23, 3, 31) {real, imag} */,
  {32'hc09f517d, 32'h40453953} /* (23, 3, 30) {real, imag} */,
  {32'hbe0b221e, 32'hbf727172} /* (23, 3, 29) {real, imag} */,
  {32'hc030707e, 32'hbf73d795} /* (23, 3, 28) {real, imag} */,
  {32'h404344ef, 32'hc0167f9a} /* (23, 3, 27) {real, imag} */,
  {32'h3eda0eaf, 32'hbfcc3e98} /* (23, 3, 26) {real, imag} */,
  {32'hbf46b213, 32'hbf817bbd} /* (23, 3, 25) {real, imag} */,
  {32'h400bf5e6, 32'h40194128} /* (23, 3, 24) {real, imag} */,
  {32'hbf24d7d3, 32'h3f85b729} /* (23, 3, 23) {real, imag} */,
  {32'h4058a784, 32'hbf254ad2} /* (23, 3, 22) {real, imag} */,
  {32'hbf89d165, 32'hbe3b2e3c} /* (23, 3, 21) {real, imag} */,
  {32'h3fcdc884, 32'h4007cfd5} /* (23, 3, 20) {real, imag} */,
  {32'h3f28be6b, 32'hc018d869} /* (23, 3, 19) {real, imag} */,
  {32'h3f8274b4, 32'hbef21d7b} /* (23, 3, 18) {real, imag} */,
  {32'hc0077093, 32'h3f8889e3} /* (23, 3, 17) {real, imag} */,
  {32'hbf1d80fc, 32'h3e65b04e} /* (23, 3, 16) {real, imag} */,
  {32'hbec1a5c6, 32'hbf3ddf20} /* (23, 3, 15) {real, imag} */,
  {32'h3f309dfa, 32'hbfa4ffff} /* (23, 3, 14) {real, imag} */,
  {32'hbfbc172f, 32'h3fb2a52c} /* (23, 3, 13) {real, imag} */,
  {32'hc0078891, 32'h407b7b3d} /* (23, 3, 12) {real, imag} */,
  {32'hbfee4223, 32'hc01d67cf} /* (23, 3, 11) {real, imag} */,
  {32'h4008887d, 32'h3fe2fdb6} /* (23, 3, 10) {real, imag} */,
  {32'h3f97ff0b, 32'hbfbce95a} /* (23, 3, 9) {real, imag} */,
  {32'hbc6f985d, 32'hc0136166} /* (23, 3, 8) {real, imag} */,
  {32'h3fa62fdd, 32'hbf852626} /* (23, 3, 7) {real, imag} */,
  {32'hbf7f1795, 32'hbf84befc} /* (23, 3, 6) {real, imag} */,
  {32'h3f96a2ce, 32'hc02493ed} /* (23, 3, 5) {real, imag} */,
  {32'h3de40bdd, 32'hbfcbf35c} /* (23, 3, 4) {real, imag} */,
  {32'h403ccb35, 32'hc0249750} /* (23, 3, 3) {real, imag} */,
  {32'hc09e6758, 32'h409d48f0} /* (23, 3, 2) {real, imag} */,
  {32'hbec1e0fc, 32'hc05dfdc6} /* (23, 3, 1) {real, imag} */,
  {32'hbdb38734, 32'hc0193730} /* (23, 3, 0) {real, imag} */,
  {32'h408f90bc, 32'h402b0af6} /* (23, 2, 31) {real, imag} */,
  {32'hc06140ec, 32'hc04f6867} /* (23, 2, 30) {real, imag} */,
  {32'hc09df5cb, 32'hc00d7d4f} /* (23, 2, 29) {real, imag} */,
  {32'h403edb13, 32'hbce35992} /* (23, 2, 28) {real, imag} */,
  {32'hbee34bb2, 32'h3fd7287d} /* (23, 2, 27) {real, imag} */,
  {32'hc097bbd2, 32'hc00ea312} /* (23, 2, 26) {real, imag} */,
  {32'h3e94fbfb, 32'h407d0d32} /* (23, 2, 25) {real, imag} */,
  {32'hbfdaa068, 32'h401bf77f} /* (23, 2, 24) {real, imag} */,
  {32'h3f0c1eb8, 32'hbfb22a83} /* (23, 2, 23) {real, imag} */,
  {32'h3fc2cf91, 32'h40425139} /* (23, 2, 22) {real, imag} */,
  {32'hbf1bad4e, 32'hc0845108} /* (23, 2, 21) {real, imag} */,
  {32'hbe3487a6, 32'hc02bae58} /* (23, 2, 20) {real, imag} */,
  {32'h4015b910, 32'hbe3cba08} /* (23, 2, 19) {real, imag} */,
  {32'hbef59f1d, 32'h4018d31e} /* (23, 2, 18) {real, imag} */,
  {32'h3e6e4797, 32'h3fc307e8} /* (23, 2, 17) {real, imag} */,
  {32'hbf5fb73e, 32'h3e3162d7} /* (23, 2, 16) {real, imag} */,
  {32'h3f654553, 32'hbf0d3a26} /* (23, 2, 15) {real, imag} */,
  {32'hbf2b0188, 32'h3f22503b} /* (23, 2, 14) {real, imag} */,
  {32'hbfe4052e, 32'h400a3a2b} /* (23, 2, 13) {real, imag} */,
  {32'h3e487ff3, 32'hbfed3350} /* (23, 2, 12) {real, imag} */,
  {32'h3f434c88, 32'hc03e2f77} /* (23, 2, 11) {real, imag} */,
  {32'hbfedcadc, 32'hc0001d24} /* (23, 2, 10) {real, imag} */,
  {32'h3fd2fb1f, 32'hbfaa02f2} /* (23, 2, 9) {real, imag} */,
  {32'h3fbef27b, 32'hc09bd6bb} /* (23, 2, 8) {real, imag} */,
  {32'h402c6be5, 32'h3f931256} /* (23, 2, 7) {real, imag} */,
  {32'hbf58da36, 32'h3fa7ab98} /* (23, 2, 6) {real, imag} */,
  {32'hbe2fd68f, 32'h404735e4} /* (23, 2, 5) {real, imag} */,
  {32'hbff79f84, 32'h3fe1747a} /* (23, 2, 4) {real, imag} */,
  {32'h3fa5be0e, 32'h405bbdbd} /* (23, 2, 3) {real, imag} */,
  {32'hbfee7678, 32'hc0bc1e31} /* (23, 2, 2) {real, imag} */,
  {32'h408ad91b, 32'hc0197944} /* (23, 2, 1) {real, imag} */,
  {32'hbdd16f89, 32'h4013ae42} /* (23, 2, 0) {real, imag} */,
  {32'hc02ed7e0, 32'hc0750b3d} /* (23, 1, 31) {real, imag} */,
  {32'hbee0795d, 32'hbf853feb} /* (23, 1, 30) {real, imag} */,
  {32'h402ca188, 32'hc019ac45} /* (23, 1, 29) {real, imag} */,
  {32'hbfde0a13, 32'hbfbca16b} /* (23, 1, 28) {real, imag} */,
  {32'h3fa9ecda, 32'h3fcadf11} /* (23, 1, 27) {real, imag} */,
  {32'h3f08902e, 32'h3dbeb6aa} /* (23, 1, 26) {real, imag} */,
  {32'h3fc8e050, 32'hbfe14e42} /* (23, 1, 25) {real, imag} */,
  {32'hbf9d6ecb, 32'h3faeb2e4} /* (23, 1, 24) {real, imag} */,
  {32'h3f81418c, 32'h3fff66be} /* (23, 1, 23) {real, imag} */,
  {32'h3f1bbd10, 32'hbe770cb3} /* (23, 1, 22) {real, imag} */,
  {32'h405c0c4a, 32'hbf86dbe6} /* (23, 1, 21) {real, imag} */,
  {32'h401ef282, 32'hbeac95e9} /* (23, 1, 20) {real, imag} */,
  {32'hbfd90c67, 32'h3fbf1f68} /* (23, 1, 19) {real, imag} */,
  {32'h3fa4b829, 32'h3f7a87c1} /* (23, 1, 18) {real, imag} */,
  {32'h3ff247b3, 32'h400469b1} /* (23, 1, 17) {real, imag} */,
  {32'h40072a6f, 32'hbfb77283} /* (23, 1, 16) {real, imag} */,
  {32'hbcba9dde, 32'h3ef7415e} /* (23, 1, 15) {real, imag} */,
  {32'hc02cc534, 32'h3fdb6b0c} /* (23, 1, 14) {real, imag} */,
  {32'hbf590bab, 32'hbf2b8d53} /* (23, 1, 13) {real, imag} */,
  {32'h3f28e0d2, 32'h4000a2bd} /* (23, 1, 12) {real, imag} */,
  {32'h4015d8fd, 32'h4006ea8c} /* (23, 1, 11) {real, imag} */,
  {32'hbf6ac2d7, 32'hbfed6f8f} /* (23, 1, 10) {real, imag} */,
  {32'hbf2dfccb, 32'hc0599e8a} /* (23, 1, 9) {real, imag} */,
  {32'hbf955d41, 32'h40774128} /* (23, 1, 8) {real, imag} */,
  {32'h400728c1, 32'h3f5392f9} /* (23, 1, 7) {real, imag} */,
  {32'hbf9d96ac, 32'hbf208883} /* (23, 1, 6) {real, imag} */,
  {32'h3fd653dd, 32'hbf267a08} /* (23, 1, 5) {real, imag} */,
  {32'hbf3046d0, 32'hc02de475} /* (23, 1, 4) {real, imag} */,
  {32'hbfbc6c65, 32'hbea5f303} /* (23, 1, 3) {real, imag} */,
  {32'hbf4e8aea, 32'h408cc193} /* (23, 1, 2) {real, imag} */,
  {32'hc0531de6, 32'hc0d21818} /* (23, 1, 1) {real, imag} */,
  {32'hc093381e, 32'hc099176f} /* (23, 1, 0) {real, imag} */,
  {32'hc09a5d46, 32'h4015fe48} /* (23, 0, 31) {real, imag} */,
  {32'hc0021e29, 32'h3f03f796} /* (23, 0, 30) {real, imag} */,
  {32'h40afc7ae, 32'h3f06c377} /* (23, 0, 29) {real, imag} */,
  {32'hc02c8495, 32'hc0153e38} /* (23, 0, 28) {real, imag} */,
  {32'h401bd1ef, 32'h3fcb4204} /* (23, 0, 27) {real, imag} */,
  {32'hbf1b0960, 32'h402e1c5c} /* (23, 0, 26) {real, imag} */,
  {32'hbfe691ea, 32'hc00263d2} /* (23, 0, 25) {real, imag} */,
  {32'h40654fa5, 32'hc0be5f0e} /* (23, 0, 24) {real, imag} */,
  {32'h3fae1b9e, 32'h3e91d2c3} /* (23, 0, 23) {real, imag} */,
  {32'hbfc46b08, 32'hc007097f} /* (23, 0, 22) {real, imag} */,
  {32'hbf54bb1b, 32'h401e43ac} /* (23, 0, 21) {real, imag} */,
  {32'h3ec04596, 32'hbf8b6c48} /* (23, 0, 20) {real, imag} */,
  {32'hbffb400d, 32'hbf303189} /* (23, 0, 19) {real, imag} */,
  {32'h3fae65eb, 32'hbfef1c08} /* (23, 0, 18) {real, imag} */,
  {32'hbe852b95, 32'h3f3727cc} /* (23, 0, 17) {real, imag} */,
  {32'h3ef93f34, 32'h3fc5475c} /* (23, 0, 16) {real, imag} */,
  {32'hbf131872, 32'hbf10de1b} /* (23, 0, 15) {real, imag} */,
  {32'hbfb2dcd6, 32'h3f84ccad} /* (23, 0, 14) {real, imag} */,
  {32'h40262e93, 32'h3f25c551} /* (23, 0, 13) {real, imag} */,
  {32'h3e2b9282, 32'h3d2f7457} /* (23, 0, 12) {real, imag} */,
  {32'hbf8fa1fc, 32'hbe2b4619} /* (23, 0, 11) {real, imag} */,
  {32'h409895ca, 32'h3f66736f} /* (23, 0, 10) {real, imag} */,
  {32'h3f751e28, 32'h403b4a7d} /* (23, 0, 9) {real, imag} */,
  {32'hc0503152, 32'h4068e117} /* (23, 0, 8) {real, imag} */,
  {32'h3f1efe38, 32'hbfa86126} /* (23, 0, 7) {real, imag} */,
  {32'hc02adc2c, 32'hbf1dc253} /* (23, 0, 6) {real, imag} */,
  {32'h3fede971, 32'h3e9e9138} /* (23, 0, 5) {real, imag} */,
  {32'h3fee085d, 32'hbeb5ab91} /* (23, 0, 4) {real, imag} */,
  {32'hc032302b, 32'hbf1e4a15} /* (23, 0, 3) {real, imag} */,
  {32'h3f8ecfa0, 32'h3f6f1d6f} /* (23, 0, 2) {real, imag} */,
  {32'hc00ee180, 32'hc0837ce9} /* (23, 0, 1) {real, imag} */,
  {32'hbf3cbe3f, 32'hc0daa393} /* (23, 0, 0) {real, imag} */,
  {32'hc0c6f1ad, 32'h3ffb317d} /* (22, 31, 31) {real, imag} */,
  {32'h3f99d0bf, 32'h4017ac5f} /* (22, 31, 30) {real, imag} */,
  {32'h3fff5fcc, 32'hc03ae37e} /* (22, 31, 29) {real, imag} */,
  {32'hbfa75200, 32'hbfab561f} /* (22, 31, 28) {real, imag} */,
  {32'h3ed04664, 32'h3f3cd501} /* (22, 31, 27) {real, imag} */,
  {32'h3fa9356a, 32'hbfdc50e6} /* (22, 31, 26) {real, imag} */,
  {32'h3fad3868, 32'hbf623d4c} /* (22, 31, 25) {real, imag} */,
  {32'hbfdaf627, 32'hbe34f5df} /* (22, 31, 24) {real, imag} */,
  {32'h40091df0, 32'hbf7fc3a1} /* (22, 31, 23) {real, imag} */,
  {32'h3d4f296c, 32'hbec3919a} /* (22, 31, 22) {real, imag} */,
  {32'h3fe457d7, 32'hc04cb76c} /* (22, 31, 21) {real, imag} */,
  {32'hbfa944f9, 32'hbe475b76} /* (22, 31, 20) {real, imag} */,
  {32'hbf473146, 32'hbc998392} /* (22, 31, 19) {real, imag} */,
  {32'h3ec112da, 32'hc06d9826} /* (22, 31, 18) {real, imag} */,
  {32'h3d2b31ae, 32'h400e2cb3} /* (22, 31, 17) {real, imag} */,
  {32'hbfcedf37, 32'hbfeeaf51} /* (22, 31, 16) {real, imag} */,
  {32'hc0026a9a, 32'h3e6843ca} /* (22, 31, 15) {real, imag} */,
  {32'hbe35c250, 32'h3ed4c88d} /* (22, 31, 14) {real, imag} */,
  {32'h3fa80ee0, 32'h3ddbf6c1} /* (22, 31, 13) {real, imag} */,
  {32'h3f99424a, 32'hbfb00233} /* (22, 31, 12) {real, imag} */,
  {32'h40493d46, 32'h3f2361d2} /* (22, 31, 11) {real, imag} */,
  {32'hc033cd48, 32'hbfb0319b} /* (22, 31, 10) {real, imag} */,
  {32'hbe99f76b, 32'hbfd98705} /* (22, 31, 9) {real, imag} */,
  {32'h3e194e06, 32'h3ebb746a} /* (22, 31, 8) {real, imag} */,
  {32'h3f063af6, 32'h3f53f031} /* (22, 31, 7) {real, imag} */,
  {32'h4084dd57, 32'hc07c1fac} /* (22, 31, 6) {real, imag} */,
  {32'h405855a2, 32'h3ffbda73} /* (22, 31, 5) {real, imag} */,
  {32'hbf889eab, 32'hc093c751} /* (22, 31, 4) {real, imag} */,
  {32'h3f817d9d, 32'h3ff3b824} /* (22, 31, 3) {real, imag} */,
  {32'h403e6834, 32'hbf39062d} /* (22, 31, 2) {real, imag} */,
  {32'hc0802796, 32'hc013f0bd} /* (22, 31, 1) {real, imag} */,
  {32'hc0112cf1, 32'hbfdbcdff} /* (22, 31, 0) {real, imag} */,
  {32'h4034da8f, 32'h3e3ca191} /* (22, 30, 31) {real, imag} */,
  {32'hc079d3ab, 32'h3d817b95} /* (22, 30, 30) {real, imag} */,
  {32'hbfcd3a82, 32'hbffbbccf} /* (22, 30, 29) {real, imag} */,
  {32'h3dd03329, 32'h403bac2a} /* (22, 30, 28) {real, imag} */,
  {32'hc029807c, 32'hbed96395} /* (22, 30, 27) {real, imag} */,
  {32'h400e869e, 32'h3f066719} /* (22, 30, 26) {real, imag} */,
  {32'h402587cd, 32'h3fda8676} /* (22, 30, 25) {real, imag} */,
  {32'hbfff0db0, 32'hc04a85f1} /* (22, 30, 24) {real, imag} */,
  {32'hbfc59f61, 32'h3f990dad} /* (22, 30, 23) {real, imag} */,
  {32'h3f80f979, 32'hbf612bbd} /* (22, 30, 22) {real, imag} */,
  {32'h4009742f, 32'h402b42d1} /* (22, 30, 21) {real, imag} */,
  {32'hbf676d5a, 32'h3f0290b1} /* (22, 30, 20) {real, imag} */,
  {32'hbf1b01d4, 32'hc063094b} /* (22, 30, 19) {real, imag} */,
  {32'hc048d2a2, 32'hbfae1f35} /* (22, 30, 18) {real, imag} */,
  {32'h403c0e32, 32'h400d6e43} /* (22, 30, 17) {real, imag} */,
  {32'h3ff26f0b, 32'h3e350b2b} /* (22, 30, 16) {real, imag} */,
  {32'hc043fcb6, 32'h3e8cc3f2} /* (22, 30, 15) {real, imag} */,
  {32'h3fc34ac9, 32'h3f9be0c6} /* (22, 30, 14) {real, imag} */,
  {32'hc01ad820, 32'hc014a858} /* (22, 30, 13) {real, imag} */,
  {32'hbffff781, 32'hbf923027} /* (22, 30, 12) {real, imag} */,
  {32'hbd443505, 32'h3f03fc25} /* (22, 30, 11) {real, imag} */,
  {32'h40827059, 32'hc01bf96a} /* (22, 30, 10) {real, imag} */,
  {32'hc00242f5, 32'h3f213c4a} /* (22, 30, 9) {real, imag} */,
  {32'h40ba3aa8, 32'h400e4500} /* (22, 30, 8) {real, imag} */,
  {32'hbe6144e5, 32'h3e8d28a0} /* (22, 30, 7) {real, imag} */,
  {32'hbf2994bc, 32'h3fe0ad3e} /* (22, 30, 6) {real, imag} */,
  {32'hbf73ae5d, 32'hbca28444} /* (22, 30, 5) {real, imag} */,
  {32'h40071ddf, 32'h3ffafc0c} /* (22, 30, 4) {real, imag} */,
  {32'hc01f9bef, 32'h4058b26c} /* (22, 30, 3) {real, imag} */,
  {32'hc0b49156, 32'h3ea2a22d} /* (22, 30, 2) {real, imag} */,
  {32'h40915925, 32'hbef604b4} /* (22, 30, 1) {real, imag} */,
  {32'h3fc99a19, 32'h3eef91fa} /* (22, 30, 0) {real, imag} */,
  {32'h3f0f3155, 32'hc00b471e} /* (22, 29, 31) {real, imag} */,
  {32'h40738009, 32'hc00f20eb} /* (22, 29, 30) {real, imag} */,
  {32'hbfa96f00, 32'h402d30c0} /* (22, 29, 29) {real, imag} */,
  {32'h3f8645c3, 32'h3fcf8dbf} /* (22, 29, 28) {real, imag} */,
  {32'h3ee42af1, 32'hbbaa31c3} /* (22, 29, 27) {real, imag} */,
  {32'h3e9ddc3a, 32'h3fe5dbbc} /* (22, 29, 26) {real, imag} */,
  {32'hbe342cd2, 32'h3f2859d1} /* (22, 29, 25) {real, imag} */,
  {32'h3f851839, 32'h3fced198} /* (22, 29, 24) {real, imag} */,
  {32'hbf6c1703, 32'h3ff9498d} /* (22, 29, 23) {real, imag} */,
  {32'hbfbcba60, 32'hbf1bf204} /* (22, 29, 22) {real, imag} */,
  {32'h3f922476, 32'h40275a31} /* (22, 29, 21) {real, imag} */,
  {32'h3ee79ed2, 32'h3f44b069} /* (22, 29, 20) {real, imag} */,
  {32'hbf9e48dc, 32'h3f97340c} /* (22, 29, 19) {real, imag} */,
  {32'hbe787dfe, 32'hbf11ca2b} /* (22, 29, 18) {real, imag} */,
  {32'h3e2ba2b6, 32'h3f37f8da} /* (22, 29, 17) {real, imag} */,
  {32'hbe8ee991, 32'h3f818b18} /* (22, 29, 16) {real, imag} */,
  {32'hbf051afc, 32'hbe179a26} /* (22, 29, 15) {real, imag} */,
  {32'h3f35904d, 32'hc017409f} /* (22, 29, 14) {real, imag} */,
  {32'h3f9d58a3, 32'hc032c67e} /* (22, 29, 13) {real, imag} */,
  {32'hc05324ba, 32'hbf42dfed} /* (22, 29, 12) {real, imag} */,
  {32'h3f05b7de, 32'hbe1b4bab} /* (22, 29, 11) {real, imag} */,
  {32'hbfc7a916, 32'h3f04d7d8} /* (22, 29, 10) {real, imag} */,
  {32'hbf9aa05f, 32'hc034a5cc} /* (22, 29, 9) {real, imag} */,
  {32'h40238516, 32'hc07c3593} /* (22, 29, 8) {real, imag} */,
  {32'h3f3ad48a, 32'h3e486953} /* (22, 29, 7) {real, imag} */,
  {32'hbfce0fb8, 32'hc02d170c} /* (22, 29, 6) {real, imag} */,
  {32'h4028e837, 32'h40117534} /* (22, 29, 5) {real, imag} */,
  {32'h3dc65705, 32'hbfb14634} /* (22, 29, 4) {real, imag} */,
  {32'h3f1a79ca, 32'h40406fc1} /* (22, 29, 3) {real, imag} */,
  {32'h40af9652, 32'h3c97124a} /* (22, 29, 2) {real, imag} */,
  {32'h40000009, 32'hc00e55aa} /* (22, 29, 1) {real, imag} */,
  {32'hbf6fde3f, 32'h3eb2a3d7} /* (22, 29, 0) {real, imag} */,
  {32'hbf8ed19a, 32'h409b5e6f} /* (22, 28, 31) {real, imag} */,
  {32'h40469f43, 32'hbfd7642a} /* (22, 28, 30) {real, imag} */,
  {32'hc029b529, 32'hc02fd856} /* (22, 28, 29) {real, imag} */,
  {32'hbd80e380, 32'h402672cf} /* (22, 28, 28) {real, imag} */,
  {32'hbed0378e, 32'h3fd756d7} /* (22, 28, 27) {real, imag} */,
  {32'hbfcd4867, 32'hbe85733f} /* (22, 28, 26) {real, imag} */,
  {32'hc08624e3, 32'h3ffffa36} /* (22, 28, 25) {real, imag} */,
  {32'hbf8faacf, 32'h3f95eae2} /* (22, 28, 24) {real, imag} */,
  {32'hbe5f1607, 32'h404aa0cb} /* (22, 28, 23) {real, imag} */,
  {32'h3f60b1b0, 32'hbf9f26b7} /* (22, 28, 22) {real, imag} */,
  {32'hc0040c3e, 32'hbedccd16} /* (22, 28, 21) {real, imag} */,
  {32'hbeb8f922, 32'hbfc5db16} /* (22, 28, 20) {real, imag} */,
  {32'h3f9f9aa4, 32'h3e66976f} /* (22, 28, 19) {real, imag} */,
  {32'h3dc9a35f, 32'hc022921d} /* (22, 28, 18) {real, imag} */,
  {32'hc019dd9c, 32'hbf4d921f} /* (22, 28, 17) {real, imag} */,
  {32'h3e39cf40, 32'h3ea3f13c} /* (22, 28, 16) {real, imag} */,
  {32'h3e960f90, 32'h3e5c2d37} /* (22, 28, 15) {real, imag} */,
  {32'h3f884887, 32'hc01b23f1} /* (22, 28, 14) {real, imag} */,
  {32'h3f3ddda8, 32'h40ae73b3} /* (22, 28, 13) {real, imag} */,
  {32'hbf83f56f, 32'hc00098c5} /* (22, 28, 12) {real, imag} */,
  {32'hbe1b9f31, 32'h3f37245d} /* (22, 28, 11) {real, imag} */,
  {32'hbfdb7c71, 32'h407163c1} /* (22, 28, 10) {real, imag} */,
  {32'hbff391fb, 32'h401f3d1e} /* (22, 28, 9) {real, imag} */,
  {32'hbf2f34a2, 32'h4093e56a} /* (22, 28, 8) {real, imag} */,
  {32'h3faaa25c, 32'hbf5ecd1e} /* (22, 28, 7) {real, imag} */,
  {32'hbfdbff57, 32'hc001ca60} /* (22, 28, 6) {real, imag} */,
  {32'h3f750961, 32'hbfafb6f3} /* (22, 28, 5) {real, imag} */,
  {32'h408e6ce8, 32'hbf34f7fb} /* (22, 28, 4) {real, imag} */,
  {32'hc05b4105, 32'hc059fd8b} /* (22, 28, 3) {real, imag} */,
  {32'h405bb3d5, 32'h3dd7b80f} /* (22, 28, 2) {real, imag} */,
  {32'h3eeaa31d, 32'h3e416681} /* (22, 28, 1) {real, imag} */,
  {32'hc0538784, 32'h3f73d7e0} /* (22, 28, 0) {real, imag} */,
  {32'h400aa003, 32'hc05a5646} /* (22, 27, 31) {real, imag} */,
  {32'h3de1832d, 32'h3f94d869} /* (22, 27, 30) {real, imag} */,
  {32'h3f34cee9, 32'h3f5e10f0} /* (22, 27, 29) {real, imag} */,
  {32'h3fdd0b8d, 32'h3fd65f7b} /* (22, 27, 28) {real, imag} */,
  {32'hc034f1d3, 32'hbfe9f1c2} /* (22, 27, 27) {real, imag} */,
  {32'hbffac1ce, 32'hc025ab2e} /* (22, 27, 26) {real, imag} */,
  {32'h4074b05b, 32'hbe702a62} /* (22, 27, 25) {real, imag} */,
  {32'hbe82b86d, 32'h3fc80b81} /* (22, 27, 24) {real, imag} */,
  {32'h3fbb4cba, 32'h3d6183bd} /* (22, 27, 23) {real, imag} */,
  {32'hbfce1b3f, 32'h40153e95} /* (22, 27, 22) {real, imag} */,
  {32'hbf512710, 32'hc0277dfd} /* (22, 27, 21) {real, imag} */,
  {32'h3f6551d8, 32'hbd42f0d0} /* (22, 27, 20) {real, imag} */,
  {32'hc00796da, 32'h400f4e61} /* (22, 27, 19) {real, imag} */,
  {32'h40270950, 32'h3faa3e2e} /* (22, 27, 18) {real, imag} */,
  {32'hbfc67d3d, 32'hbf7aec49} /* (22, 27, 17) {real, imag} */,
  {32'hbf93a3ee, 32'h3e8a5f2c} /* (22, 27, 16) {real, imag} */,
  {32'h3fedaaa1, 32'h3e77a1f4} /* (22, 27, 15) {real, imag} */,
  {32'hbef69b1d, 32'h3fd78ca4} /* (22, 27, 14) {real, imag} */,
  {32'hbef6121f, 32'h3fcaaa27} /* (22, 27, 13) {real, imag} */,
  {32'hbc29e98c, 32'hbf9c3510} /* (22, 27, 12) {real, imag} */,
  {32'h3fa86a19, 32'h3f7b5156} /* (22, 27, 11) {real, imag} */,
  {32'hbfc9d177, 32'hc0acab65} /* (22, 27, 10) {real, imag} */,
  {32'h3bbd4e62, 32'hbfba76d5} /* (22, 27, 9) {real, imag} */,
  {32'hbfca9484, 32'h3fc37305} /* (22, 27, 8) {real, imag} */,
  {32'hbdadd4d1, 32'h3f074483} /* (22, 27, 7) {real, imag} */,
  {32'h3ffba6f1, 32'hc017c68b} /* (22, 27, 6) {real, imag} */,
  {32'hc0335a35, 32'h3f157e4c} /* (22, 27, 5) {real, imag} */,
  {32'hbf21496b, 32'h3f9af39e} /* (22, 27, 4) {real, imag} */,
  {32'h3ffb724c, 32'hbd1f73dd} /* (22, 27, 3) {real, imag} */,
  {32'hbf29d46e, 32'hc012d480} /* (22, 27, 2) {real, imag} */,
  {32'hc003262f, 32'h40a801b3} /* (22, 27, 1) {real, imag} */,
  {32'h40168054, 32'h404c39a3} /* (22, 27, 0) {real, imag} */,
  {32'h3f4d6435, 32'hc0537bfa} /* (22, 26, 31) {real, imag} */,
  {32'hc06ff9db, 32'h3fc66f5f} /* (22, 26, 30) {real, imag} */,
  {32'h4002e242, 32'hbfa3869b} /* (22, 26, 29) {real, imag} */,
  {32'h3dd39a64, 32'hbf4cc599} /* (22, 26, 28) {real, imag} */,
  {32'hbf8d310e, 32'h3f9b9fec} /* (22, 26, 27) {real, imag} */,
  {32'h3eb3fba7, 32'hbfe28c2f} /* (22, 26, 26) {real, imag} */,
  {32'h3f845d82, 32'h403b74a2} /* (22, 26, 25) {real, imag} */,
  {32'h408aa356, 32'hbfd67756} /* (22, 26, 24) {real, imag} */,
  {32'hbfbd2a2d, 32'hbdd2fa33} /* (22, 26, 23) {real, imag} */,
  {32'hc0674205, 32'h3ff88a96} /* (22, 26, 22) {real, imag} */,
  {32'hbd4f4668, 32'hc06f1b51} /* (22, 26, 21) {real, imag} */,
  {32'hbe2c5411, 32'hbfe0b90b} /* (22, 26, 20) {real, imag} */,
  {32'h3f3f5d85, 32'h4014e0af} /* (22, 26, 19) {real, imag} */,
  {32'h3e1710c9, 32'hbfddae66} /* (22, 26, 18) {real, imag} */,
  {32'hc01d659a, 32'hc00713ee} /* (22, 26, 17) {real, imag} */,
  {32'hbfb81417, 32'hbe91219d} /* (22, 26, 16) {real, imag} */,
  {32'hbf565831, 32'hbf068e6d} /* (22, 26, 15) {real, imag} */,
  {32'h3d24f8b4, 32'h404c4ad0} /* (22, 26, 14) {real, imag} */,
  {32'hbe178999, 32'hc005569d} /* (22, 26, 13) {real, imag} */,
  {32'h3ff485bd, 32'h3dd5fe71} /* (22, 26, 12) {real, imag} */,
  {32'hbdc4499d, 32'h3f021626} /* (22, 26, 11) {real, imag} */,
  {32'hbf6269f7, 32'hc095a3ca} /* (22, 26, 10) {real, imag} */,
  {32'h40402f5c, 32'h401a24c5} /* (22, 26, 9) {real, imag} */,
  {32'h3ea67c83, 32'hbf6df1ce} /* (22, 26, 8) {real, imag} */,
  {32'h3e7a7bc1, 32'h3f0690ac} /* (22, 26, 7) {real, imag} */,
  {32'hbe20dfb3, 32'h3ee16a7b} /* (22, 26, 6) {real, imag} */,
  {32'hbeb9180f, 32'h40476c33} /* (22, 26, 5) {real, imag} */,
  {32'h405845be, 32'hbe13b4c9} /* (22, 26, 4) {real, imag} */,
  {32'hc091fbb4, 32'h3d1ba9bc} /* (22, 26, 3) {real, imag} */,
  {32'h3e1a7411, 32'hbfa01c07} /* (22, 26, 2) {real, imag} */,
  {32'h3fd36b9b, 32'h3fa1ea66} /* (22, 26, 1) {real, imag} */,
  {32'hc0291434, 32'h3fc0168f} /* (22, 26, 0) {real, imag} */,
  {32'h3ec4bbc5, 32'h404dbded} /* (22, 25, 31) {real, imag} */,
  {32'hbfc94de0, 32'h406578ca} /* (22, 25, 30) {real, imag} */,
  {32'hbf1a48da, 32'hbfae5256} /* (22, 25, 29) {real, imag} */,
  {32'h3eb7338a, 32'h3fa79e44} /* (22, 25, 28) {real, imag} */,
  {32'h3f4e94c5, 32'h4001bac3} /* (22, 25, 27) {real, imag} */,
  {32'h3f7a8153, 32'h403145ee} /* (22, 25, 26) {real, imag} */,
  {32'hbf536a2b, 32'hbedbca99} /* (22, 25, 25) {real, imag} */,
  {32'hbf8ce558, 32'h3f0e7af9} /* (22, 25, 24) {real, imag} */,
  {32'h3ffdaec4, 32'h402c0bd2} /* (22, 25, 23) {real, imag} */,
  {32'hc00bc91e, 32'h408307b8} /* (22, 25, 22) {real, imag} */,
  {32'h3fabb16a, 32'hbf7e9b6f} /* (22, 25, 21) {real, imag} */,
  {32'hbfac5c3a, 32'hbf791f2f} /* (22, 25, 20) {real, imag} */,
  {32'h404475d6, 32'h3c3a4bc3} /* (22, 25, 19) {real, imag} */,
  {32'h3ec2efa4, 32'h3f84f9c9} /* (22, 25, 18) {real, imag} */,
  {32'hc0019500, 32'hbf8a02b7} /* (22, 25, 17) {real, imag} */,
  {32'hbec8173a, 32'h404c4e20} /* (22, 25, 16) {real, imag} */,
  {32'hbf27cda2, 32'hc04110df} /* (22, 25, 15) {real, imag} */,
  {32'h3f11209b, 32'h3e94030b} /* (22, 25, 14) {real, imag} */,
  {32'hbf4fde3b, 32'h40349082} /* (22, 25, 13) {real, imag} */,
  {32'hbf06d25b, 32'h3f4aeb29} /* (22, 25, 12) {real, imag} */,
  {32'hbedbe6cd, 32'h400b4ec1} /* (22, 25, 11) {real, imag} */,
  {32'h3e2cc0ed, 32'h3fd1b4af} /* (22, 25, 10) {real, imag} */,
  {32'h3fc5ff16, 32'h400dce63} /* (22, 25, 9) {real, imag} */,
  {32'h3f61500b, 32'h4086844f} /* (22, 25, 8) {real, imag} */,
  {32'h402b2d59, 32'h3fba38b3} /* (22, 25, 7) {real, imag} */,
  {32'h3f400b58, 32'h3f2ca8bc} /* (22, 25, 6) {real, imag} */,
  {32'h3ff52553, 32'hc01f03c3} /* (22, 25, 5) {real, imag} */,
  {32'h40332444, 32'hc00bfc07} /* (22, 25, 4) {real, imag} */,
  {32'hbfc60fce, 32'hbf09ea20} /* (22, 25, 3) {real, imag} */,
  {32'h3f140983, 32'hc03d14ac} /* (22, 25, 2) {real, imag} */,
  {32'hbfdfdbc3, 32'hc02090f5} /* (22, 25, 1) {real, imag} */,
  {32'h3fe552dd, 32'h4000af49} /* (22, 25, 0) {real, imag} */,
  {32'hbf6210f0, 32'hbfa19aa5} /* (22, 24, 31) {real, imag} */,
  {32'hc0302b1b, 32'h3fe5a293} /* (22, 24, 30) {real, imag} */,
  {32'h40459ec3, 32'h3f9926bc} /* (22, 24, 29) {real, imag} */,
  {32'h3f3539fb, 32'hc02b6639} /* (22, 24, 28) {real, imag} */,
  {32'h3faaf357, 32'h40010822} /* (22, 24, 27) {real, imag} */,
  {32'h404ff133, 32'hbfc06ccc} /* (22, 24, 26) {real, imag} */,
  {32'h408bc487, 32'h3e6ea931} /* (22, 24, 25) {real, imag} */,
  {32'hbed79700, 32'hc05acbd7} /* (22, 24, 24) {real, imag} */,
  {32'hc01ddfe9, 32'h3fab8e98} /* (22, 24, 23) {real, imag} */,
  {32'hbdc9859a, 32'h3ed3c894} /* (22, 24, 22) {real, imag} */,
  {32'h4044fe80, 32'h3eae749f} /* (22, 24, 21) {real, imag} */,
  {32'hc05b2368, 32'hbfcd1334} /* (22, 24, 20) {real, imag} */,
  {32'h3fab53d0, 32'hbfad830f} /* (22, 24, 19) {real, imag} */,
  {32'h40017313, 32'h4016d908} /* (22, 24, 18) {real, imag} */,
  {32'h3e42c791, 32'hbf989bf3} /* (22, 24, 17) {real, imag} */,
  {32'h3fd6669f, 32'hbfbb08fc} /* (22, 24, 16) {real, imag} */,
  {32'h3e1f6444, 32'h3fe8fba1} /* (22, 24, 15) {real, imag} */,
  {32'h3fc17d9c, 32'h3f3be9d0} /* (22, 24, 14) {real, imag} */,
  {32'h3e39256d, 32'h3fad19be} /* (22, 24, 13) {real, imag} */,
  {32'hc023cc80, 32'hbff856b7} /* (22, 24, 12) {real, imag} */,
  {32'h3dbe2885, 32'hbfa81ef7} /* (22, 24, 11) {real, imag} */,
  {32'hbf96ea19, 32'h3f07baca} /* (22, 24, 10) {real, imag} */,
  {32'hbe37e526, 32'hbf3b8d25} /* (22, 24, 9) {real, imag} */,
  {32'h3fbac5c4, 32'hbe75a383} /* (22, 24, 8) {real, imag} */,
  {32'hc039ec5d, 32'hbecfeaaa} /* (22, 24, 7) {real, imag} */,
  {32'hc0583d9e, 32'h3f88dd28} /* (22, 24, 6) {real, imag} */,
  {32'h4000d970, 32'h3ee01724} /* (22, 24, 5) {real, imag} */,
  {32'hbfcd77a8, 32'h40060ea8} /* (22, 24, 4) {real, imag} */,
  {32'hc0046efc, 32'hbf7ca0b3} /* (22, 24, 3) {real, imag} */,
  {32'hbf6f5b67, 32'hbfc883a1} /* (22, 24, 2) {real, imag} */,
  {32'hbec90470, 32'hbf1f56ef} /* (22, 24, 1) {real, imag} */,
  {32'h407c9133, 32'h3fba31ee} /* (22, 24, 0) {real, imag} */,
  {32'hbfee8b15, 32'hc009cbf3} /* (22, 23, 31) {real, imag} */,
  {32'hbe822e96, 32'hc0945261} /* (22, 23, 30) {real, imag} */,
  {32'h40175395, 32'hbfd3448b} /* (22, 23, 29) {real, imag} */,
  {32'h3fb15e18, 32'hbf9d64e3} /* (22, 23, 28) {real, imag} */,
  {32'hbeef6455, 32'hbf32a9ae} /* (22, 23, 27) {real, imag} */,
  {32'h3f22b18a, 32'h3f8bfb21} /* (22, 23, 26) {real, imag} */,
  {32'h403d7fff, 32'hc063ac1d} /* (22, 23, 25) {real, imag} */,
  {32'h40860e1a, 32'hbdf5774a} /* (22, 23, 24) {real, imag} */,
  {32'h3e768ae4, 32'hc032e8b6} /* (22, 23, 23) {real, imag} */,
  {32'h3f99a054, 32'h403f56ab} /* (22, 23, 22) {real, imag} */,
  {32'h3f7ce782, 32'h3fe662ad} /* (22, 23, 21) {real, imag} */,
  {32'h3f8dfe67, 32'hbdf2d8e7} /* (22, 23, 20) {real, imag} */,
  {32'hc04eebcb, 32'hbee49202} /* (22, 23, 19) {real, imag} */,
  {32'hbf340c7a, 32'hbe390c02} /* (22, 23, 18) {real, imag} */,
  {32'h3f83ac21, 32'h3dd5618e} /* (22, 23, 17) {real, imag} */,
  {32'hbe1a1bca, 32'hbfd90bd4} /* (22, 23, 16) {real, imag} */,
  {32'hbde6d90d, 32'hbfc1d743} /* (22, 23, 15) {real, imag} */,
  {32'hbfd0b506, 32'hbf08f070} /* (22, 23, 14) {real, imag} */,
  {32'hbf918c27, 32'hbe8cba51} /* (22, 23, 13) {real, imag} */,
  {32'hc03b82f1, 32'h3f8aaff8} /* (22, 23, 12) {real, imag} */,
  {32'hc000c1af, 32'h3f70abb3} /* (22, 23, 11) {real, imag} */,
  {32'hbfbd7f34, 32'hc06ace24} /* (22, 23, 10) {real, imag} */,
  {32'hbf886543, 32'hc01bb668} /* (22, 23, 9) {real, imag} */,
  {32'h3f5710e3, 32'h3c89197f} /* (22, 23, 8) {real, imag} */,
  {32'h3ef0acf2, 32'h3f083041} /* (22, 23, 7) {real, imag} */,
  {32'hbda418cb, 32'h400bd930} /* (22, 23, 6) {real, imag} */,
  {32'h3febc31d, 32'hc0131c6c} /* (22, 23, 5) {real, imag} */,
  {32'hbf1c00ec, 32'hbf3f3be7} /* (22, 23, 4) {real, imag} */,
  {32'h3efc3426, 32'hc0052a97} /* (22, 23, 3) {real, imag} */,
  {32'hbff380a4, 32'hbf9df8ff} /* (22, 23, 2) {real, imag} */,
  {32'h3f53e147, 32'hbf664910} /* (22, 23, 1) {real, imag} */,
  {32'h3dc20707, 32'h401e9c6c} /* (22, 23, 0) {real, imag} */,
  {32'h403851c9, 32'h3fdfd941} /* (22, 22, 31) {real, imag} */,
  {32'h3f9e3991, 32'h3fb4eb7b} /* (22, 22, 30) {real, imag} */,
  {32'h3fd26bad, 32'hbe7154fd} /* (22, 22, 29) {real, imag} */,
  {32'hc0122404, 32'h406b0370} /* (22, 22, 28) {real, imag} */,
  {32'hbebea6cc, 32'h3f06e482} /* (22, 22, 27) {real, imag} */,
  {32'h3fe84b95, 32'hc0508d57} /* (22, 22, 26) {real, imag} */,
  {32'hbfbba98d, 32'h3f7c069e} /* (22, 22, 25) {real, imag} */,
  {32'hbe7dd266, 32'hbff8d187} /* (22, 22, 24) {real, imag} */,
  {32'hc029bf98, 32'h3fb9313f} /* (22, 22, 23) {real, imag} */,
  {32'hc054ff42, 32'h3f2bb2f5} /* (22, 22, 22) {real, imag} */,
  {32'h40571001, 32'h40053009} /* (22, 22, 21) {real, imag} */,
  {32'h3dd41362, 32'h3fd50f0e} /* (22, 22, 20) {real, imag} */,
  {32'h3e270f30, 32'h3fc1124f} /* (22, 22, 19) {real, imag} */,
  {32'h3e914caa, 32'hc0349833} /* (22, 22, 18) {real, imag} */,
  {32'h402e0ac2, 32'h3f131343} /* (22, 22, 17) {real, imag} */,
  {32'hbfbf8ccd, 32'h3e5f92c9} /* (22, 22, 16) {real, imag} */,
  {32'h3f026efb, 32'h3fa53952} /* (22, 22, 15) {real, imag} */,
  {32'hbf2842ca, 32'hc02ecad7} /* (22, 22, 14) {real, imag} */,
  {32'h403513c0, 32'hbfae2b69} /* (22, 22, 13) {real, imag} */,
  {32'h3fb00f53, 32'h3ff0defe} /* (22, 22, 12) {real, imag} */,
  {32'h405b5f49, 32'hbd8ae73a} /* (22, 22, 11) {real, imag} */,
  {32'h3ebd19e4, 32'hc07cf4c1} /* (22, 22, 10) {real, imag} */,
  {32'h403cf4e5, 32'h4048bf4b} /* (22, 22, 9) {real, imag} */,
  {32'h401e5587, 32'h3ef46446} /* (22, 22, 8) {real, imag} */,
  {32'h3ee7358f, 32'hbf06d111} /* (22, 22, 7) {real, imag} */,
  {32'hbf8b9d5e, 32'h3f1dcdcf} /* (22, 22, 6) {real, imag} */,
  {32'h3f3fec26, 32'h40005c04} /* (22, 22, 5) {real, imag} */,
  {32'hbfbbe794, 32'hbfef80c1} /* (22, 22, 4) {real, imag} */,
  {32'h3fa6c51c, 32'hbf85a963} /* (22, 22, 3) {real, imag} */,
  {32'h3f847530, 32'h3e6810df} /* (22, 22, 2) {real, imag} */,
  {32'h3ff134e3, 32'hbfa80605} /* (22, 22, 1) {real, imag} */,
  {32'hbf5dec20, 32'hbd30a3d1} /* (22, 22, 0) {real, imag} */,
  {32'hbe0a8627, 32'h401513fa} /* (22, 21, 31) {real, imag} */,
  {32'h3db6850e, 32'hbe049052} /* (22, 21, 30) {real, imag} */,
  {32'hc0648e19, 32'hbeb1ee73} /* (22, 21, 29) {real, imag} */,
  {32'hc097ebbc, 32'h3e49f4a2} /* (22, 21, 28) {real, imag} */,
  {32'hbe30b894, 32'hc05afa83} /* (22, 21, 27) {real, imag} */,
  {32'h3e7d50c2, 32'h400d7e3e} /* (22, 21, 26) {real, imag} */,
  {32'hbec71054, 32'h405183a3} /* (22, 21, 25) {real, imag} */,
  {32'hbf0a94f4, 32'hc0cf6629} /* (22, 21, 24) {real, imag} */,
  {32'hbff12934, 32'hbfa8ec29} /* (22, 21, 23) {real, imag} */,
  {32'hbfbba844, 32'hbf094c9a} /* (22, 21, 22) {real, imag} */,
  {32'hc024a0c0, 32'hc01d568e} /* (22, 21, 21) {real, imag} */,
  {32'h3f1f14ee, 32'hbf14731a} /* (22, 21, 20) {real, imag} */,
  {32'h401603d0, 32'h3e6ea323} /* (22, 21, 19) {real, imag} */,
  {32'hbfb10537, 32'hbc18c3a8} /* (22, 21, 18) {real, imag} */,
  {32'h3efcd476, 32'h3ebb8e05} /* (22, 21, 17) {real, imag} */,
  {32'hbf88d3ca, 32'h40107fa5} /* (22, 21, 16) {real, imag} */,
  {32'h3fb5f98c, 32'hbf803581} /* (22, 21, 15) {real, imag} */,
  {32'hbfb31bd0, 32'hc028e9c7} /* (22, 21, 14) {real, imag} */,
  {32'h3fc94751, 32'h3f6787e0} /* (22, 21, 13) {real, imag} */,
  {32'h3ec2faea, 32'h404ad4c1} /* (22, 21, 12) {real, imag} */,
  {32'hc05fd1d6, 32'h40377047} /* (22, 21, 11) {real, imag} */,
  {32'hc08b41e1, 32'hc06104c8} /* (22, 21, 10) {real, imag} */,
  {32'hc01c4248, 32'hbfc7078e} /* (22, 21, 9) {real, imag} */,
  {32'hbff53f37, 32'hc091605e} /* (22, 21, 8) {real, imag} */,
  {32'h3f945bcc, 32'hbee5a884} /* (22, 21, 7) {real, imag} */,
  {32'hbf3b14d2, 32'hc029fb7f} /* (22, 21, 6) {real, imag} */,
  {32'hbfc0621f, 32'h3f8df519} /* (22, 21, 5) {real, imag} */,
  {32'h3e1fcb00, 32'h407fa7d4} /* (22, 21, 4) {real, imag} */,
  {32'h40591187, 32'hbf9b622f} /* (22, 21, 3) {real, imag} */,
  {32'h3debd6a2, 32'h40779052} /* (22, 21, 2) {real, imag} */,
  {32'hbb0215f2, 32'h4020c9c5} /* (22, 21, 1) {real, imag} */,
  {32'hbfeea6fa, 32'hbf1d1e02} /* (22, 21, 0) {real, imag} */,
  {32'h3e44c6bc, 32'h40240cb1} /* (22, 20, 31) {real, imag} */,
  {32'h4017bfcd, 32'h3f3c9eb6} /* (22, 20, 30) {real, imag} */,
  {32'hbeaeb71e, 32'hbf25b61a} /* (22, 20, 29) {real, imag} */,
  {32'hbf62c5eb, 32'h3ad7ed99} /* (22, 20, 28) {real, imag} */,
  {32'hc09d721f, 32'hc0030c53} /* (22, 20, 27) {real, imag} */,
  {32'hbfac7f26, 32'hbf148a2a} /* (22, 20, 26) {real, imag} */,
  {32'h4036ec43, 32'h402b280a} /* (22, 20, 25) {real, imag} */,
  {32'h3f90b405, 32'h407e5f85} /* (22, 20, 24) {real, imag} */,
  {32'h3ff6cbac, 32'hc0485842} /* (22, 20, 23) {real, imag} */,
  {32'h3f0b4b5d, 32'hc05cc0fc} /* (22, 20, 22) {real, imag} */,
  {32'h3fe67047, 32'h3f317b3b} /* (22, 20, 21) {real, imag} */,
  {32'h3fa77b0e, 32'hbe231724} /* (22, 20, 20) {real, imag} */,
  {32'h4028cadb, 32'h3fc4ec04} /* (22, 20, 19) {real, imag} */,
  {32'h40502467, 32'h3ee6c891} /* (22, 20, 18) {real, imag} */,
  {32'h3e2350f7, 32'hc05df816} /* (22, 20, 17) {real, imag} */,
  {32'hc01c6be1, 32'h3db65edf} /* (22, 20, 16) {real, imag} */,
  {32'h3e02a4a1, 32'h3faaf340} /* (22, 20, 15) {real, imag} */,
  {32'h3fa1830c, 32'hbcb46037} /* (22, 20, 14) {real, imag} */,
  {32'h4042156f, 32'h4019b692} /* (22, 20, 13) {real, imag} */,
  {32'hbd861c0b, 32'hbfae976a} /* (22, 20, 12) {real, imag} */,
  {32'hc029d234, 32'hbfae9ee3} /* (22, 20, 11) {real, imag} */,
  {32'hc027ac65, 32'h3e09d0d4} /* (22, 20, 10) {real, imag} */,
  {32'h3fb59e63, 32'hbf4618ed} /* (22, 20, 9) {real, imag} */,
  {32'hc03a0465, 32'h407a8e8c} /* (22, 20, 8) {real, imag} */,
  {32'hc002d927, 32'hbc0b90af} /* (22, 20, 7) {real, imag} */,
  {32'h3f99b4fe, 32'h3f769837} /* (22, 20, 6) {real, imag} */,
  {32'hbfcad4eb, 32'hc07d7550} /* (22, 20, 5) {real, imag} */,
  {32'h403e9f15, 32'h3e2d73fd} /* (22, 20, 4) {real, imag} */,
  {32'h3ff4b707, 32'hbf4da56b} /* (22, 20, 3) {real, imag} */,
  {32'h4024b266, 32'hbf3c231b} /* (22, 20, 2) {real, imag} */,
  {32'h3e988290, 32'hc01f4aa8} /* (22, 20, 1) {real, imag} */,
  {32'hc046768a, 32'hbc6f38ed} /* (22, 20, 0) {real, imag} */,
  {32'hbf4488c1, 32'h3fcd7066} /* (22, 19, 31) {real, imag} */,
  {32'h3f76e24d, 32'h3e885eb0} /* (22, 19, 30) {real, imag} */,
  {32'h3f1661ec, 32'hbf265447} /* (22, 19, 29) {real, imag} */,
  {32'hbf79e366, 32'hbea8d56e} /* (22, 19, 28) {real, imag} */,
  {32'h3fe41b62, 32'hbfb3712c} /* (22, 19, 27) {real, imag} */,
  {32'h3e98da25, 32'h3d4e2d80} /* (22, 19, 26) {real, imag} */,
  {32'h3fbce31b, 32'hbe6e6708} /* (22, 19, 25) {real, imag} */,
  {32'h3f76ad13, 32'h3f0f9137} /* (22, 19, 24) {real, imag} */,
  {32'h3e8346f2, 32'hc02410a2} /* (22, 19, 23) {real, imag} */,
  {32'h4049cc4a, 32'h3dbd38be} /* (22, 19, 22) {real, imag} */,
  {32'hbf91cbe6, 32'hbfc3572c} /* (22, 19, 21) {real, imag} */,
  {32'h401876e5, 32'h3ea2d722} /* (22, 19, 20) {real, imag} */,
  {32'hbfffad27, 32'h3ff7bbd1} /* (22, 19, 19) {real, imag} */,
  {32'hbfb6f36c, 32'h3f9664ec} /* (22, 19, 18) {real, imag} */,
  {32'h3dce66c4, 32'hc0336e9a} /* (22, 19, 17) {real, imag} */,
  {32'hbf8fbbb2, 32'h407e9809} /* (22, 19, 16) {real, imag} */,
  {32'hbf1423d3, 32'hbf2e36a8} /* (22, 19, 15) {real, imag} */,
  {32'hc006e442, 32'hc0849903} /* (22, 19, 14) {real, imag} */,
  {32'h400364a7, 32'hc008e64a} /* (22, 19, 13) {real, imag} */,
  {32'hc03b1880, 32'hc08a98a6} /* (22, 19, 12) {real, imag} */,
  {32'hbd285919, 32'h3e8a9ca0} /* (22, 19, 11) {real, imag} */,
  {32'h3e857859, 32'hbf32e44d} /* (22, 19, 10) {real, imag} */,
  {32'h3fea6268, 32'h3f4e3788} /* (22, 19, 9) {real, imag} */,
  {32'hbfda1776, 32'h3b853030} /* (22, 19, 8) {real, imag} */,
  {32'h3fa1a393, 32'h3edba50f} /* (22, 19, 7) {real, imag} */,
  {32'h3f72e428, 32'hbfb7df88} /* (22, 19, 6) {real, imag} */,
  {32'h4000282a, 32'hbe74c5d6} /* (22, 19, 5) {real, imag} */,
  {32'hbfc78914, 32'h3fe5c1af} /* (22, 19, 4) {real, imag} */,
  {32'hc02d110b, 32'h3f6d1e9b} /* (22, 19, 3) {real, imag} */,
  {32'h3fd3af73, 32'h3efd121f} /* (22, 19, 2) {real, imag} */,
  {32'h4004ae51, 32'h3f3f9be7} /* (22, 19, 1) {real, imag} */,
  {32'h3f4a081d, 32'hc03edc98} /* (22, 19, 0) {real, imag} */,
  {32'hc0329400, 32'hc05a3e43} /* (22, 18, 31) {real, imag} */,
  {32'hbf9daf8a, 32'h3d0a0ddc} /* (22, 18, 30) {real, imag} */,
  {32'h3fd37897, 32'h3dfe3d42} /* (22, 18, 29) {real, imag} */,
  {32'h3e4c821b, 32'hc02ea5ae} /* (22, 18, 28) {real, imag} */,
  {32'hbfb75ff1, 32'h3fba43eb} /* (22, 18, 27) {real, imag} */,
  {32'hbf0b2246, 32'h401d9800} /* (22, 18, 26) {real, imag} */,
  {32'h3f130675, 32'h400257d1} /* (22, 18, 25) {real, imag} */,
  {32'hbe5116ca, 32'h3f6f805b} /* (22, 18, 24) {real, imag} */,
  {32'hc03e3c34, 32'h3f832e1c} /* (22, 18, 23) {real, imag} */,
  {32'h3ee19e3a, 32'h4086bf73} /* (22, 18, 22) {real, imag} */,
  {32'hc01f290e, 32'h3f56e59b} /* (22, 18, 21) {real, imag} */,
  {32'h3fff33e0, 32'hbfd8bfbd} /* (22, 18, 20) {real, imag} */,
  {32'hbde23a87, 32'hbe8885ba} /* (22, 18, 19) {real, imag} */,
  {32'hbed78420, 32'hc0273fda} /* (22, 18, 18) {real, imag} */,
  {32'hbfb1b9e4, 32'hc011b52f} /* (22, 18, 17) {real, imag} */,
  {32'h3f82cb96, 32'h3e5cde0f} /* (22, 18, 16) {real, imag} */,
  {32'hbf95c28d, 32'h408676fb} /* (22, 18, 15) {real, imag} */,
  {32'hc00b1884, 32'h3e475150} /* (22, 18, 14) {real, imag} */,
  {32'hc00c2ab0, 32'h3e8503a9} /* (22, 18, 13) {real, imag} */,
  {32'h4066227c, 32'hbf8f48e3} /* (22, 18, 12) {real, imag} */,
  {32'h401a7f2e, 32'hbfa4e089} /* (22, 18, 11) {real, imag} */,
  {32'h403200da, 32'hbed919f3} /* (22, 18, 10) {real, imag} */,
  {32'h3fc3b4fc, 32'h402546e2} /* (22, 18, 9) {real, imag} */,
  {32'h3f08c5d7, 32'h3f2ea662} /* (22, 18, 8) {real, imag} */,
  {32'hbf8cb4c5, 32'h3fbff869} /* (22, 18, 7) {real, imag} */,
  {32'h3f8e73bb, 32'h3febb425} /* (22, 18, 6) {real, imag} */,
  {32'h3d58adf9, 32'hc00a2a74} /* (22, 18, 5) {real, imag} */,
  {32'h3fdb30d5, 32'hbe44ea03} /* (22, 18, 4) {real, imag} */,
  {32'hbfc7a4de, 32'h3f818954} /* (22, 18, 3) {real, imag} */,
  {32'h3ff32c9a, 32'hbe62015e} /* (22, 18, 2) {real, imag} */,
  {32'h3e22d61d, 32'hbe9f2dcf} /* (22, 18, 1) {real, imag} */,
  {32'hbf97d98e, 32'hbfab4e52} /* (22, 18, 0) {real, imag} */,
  {32'hbe832cb5, 32'h3f093f3b} /* (22, 17, 31) {real, imag} */,
  {32'h3e72fa52, 32'hbed9ea05} /* (22, 17, 30) {real, imag} */,
  {32'h3e977207, 32'h3ea4b5b0} /* (22, 17, 29) {real, imag} */,
  {32'h3f5ade3d, 32'hbdb7e922} /* (22, 17, 28) {real, imag} */,
  {32'h4036649c, 32'hbe36b818} /* (22, 17, 27) {real, imag} */,
  {32'hbeaa63c2, 32'hbe93182f} /* (22, 17, 26) {real, imag} */,
  {32'h3f73cc44, 32'hc01d1b80} /* (22, 17, 25) {real, imag} */,
  {32'h3ea6f73c, 32'hbdf9a6b5} /* (22, 17, 24) {real, imag} */,
  {32'h3ed865ff, 32'h4032919b} /* (22, 17, 23) {real, imag} */,
  {32'hbf4524f2, 32'hbf960b0e} /* (22, 17, 22) {real, imag} */,
  {32'h3fb457b1, 32'h403af092} /* (22, 17, 21) {real, imag} */,
  {32'hbefa1ef7, 32'hbfb72782} /* (22, 17, 20) {real, imag} */,
  {32'hbf03eee4, 32'h405e153d} /* (22, 17, 19) {real, imag} */,
  {32'hbfea0d2b, 32'hc0771734} /* (22, 17, 18) {real, imag} */,
  {32'hbed59b0a, 32'h3f86666b} /* (22, 17, 17) {real, imag} */,
  {32'h3f6d7c14, 32'hbf07fc11} /* (22, 17, 16) {real, imag} */,
  {32'hbea7915a, 32'h3f31af4d} /* (22, 17, 15) {real, imag} */,
  {32'h3f751aea, 32'h3fbe066c} /* (22, 17, 14) {real, imag} */,
  {32'h3fb148d5, 32'hc099b764} /* (22, 17, 13) {real, imag} */,
  {32'hbd9d5b7e, 32'h4018c0f2} /* (22, 17, 12) {real, imag} */,
  {32'hbf11971e, 32'hbfa7fec8} /* (22, 17, 11) {real, imag} */,
  {32'h4046b427, 32'hbed5f439} /* (22, 17, 10) {real, imag} */,
  {32'hc049fddc, 32'hbfe02144} /* (22, 17, 9) {real, imag} */,
  {32'hbdd7bc96, 32'hc035ad65} /* (22, 17, 8) {real, imag} */,
  {32'h4047d1f5, 32'h408fc273} /* (22, 17, 7) {real, imag} */,
  {32'hbf3f3df8, 32'h3f028c5f} /* (22, 17, 6) {real, imag} */,
  {32'hbfb8e0f7, 32'h3bbb7337} /* (22, 17, 5) {real, imag} */,
  {32'hbf34e70e, 32'h3e4abf96} /* (22, 17, 4) {real, imag} */,
  {32'h3f9889cc, 32'hbfd7119b} /* (22, 17, 3) {real, imag} */,
  {32'h3f9beb90, 32'hbf588d7e} /* (22, 17, 2) {real, imag} */,
  {32'hbe68475a, 32'hbf6808c5} /* (22, 17, 1) {real, imag} */,
  {32'h3dd8349d, 32'hc00dc4f1} /* (22, 17, 0) {real, imag} */,
  {32'h3fe54e1c, 32'hbf1b29c8} /* (22, 16, 31) {real, imag} */,
  {32'h3fb262c7, 32'h3f3047d8} /* (22, 16, 30) {real, imag} */,
  {32'h4000fac2, 32'hbfa8919b} /* (22, 16, 29) {real, imag} */,
  {32'h3ff7d1b9, 32'hbf5db462} /* (22, 16, 28) {real, imag} */,
  {32'h3f1182e9, 32'h3fa22bca} /* (22, 16, 27) {real, imag} */,
  {32'hbf1cfdd1, 32'hbf4ca268} /* (22, 16, 26) {real, imag} */,
  {32'hbd066b41, 32'h3e524078} /* (22, 16, 25) {real, imag} */,
  {32'hbfbe304e, 32'hbfab2491} /* (22, 16, 24) {real, imag} */,
  {32'h3f1f29db, 32'h3f402675} /* (22, 16, 23) {real, imag} */,
  {32'h3ebe931c, 32'hbbcdf030} /* (22, 16, 22) {real, imag} */,
  {32'h3df1ad81, 32'hbfd37660} /* (22, 16, 21) {real, imag} */,
  {32'h3df04954, 32'hbf76c7f0} /* (22, 16, 20) {real, imag} */,
  {32'hbfea9ca7, 32'hbef921a2} /* (22, 16, 19) {real, imag} */,
  {32'h3fcef83d, 32'hbfd9e69c} /* (22, 16, 18) {real, imag} */,
  {32'h3f81560f, 32'h3fd36cf0} /* (22, 16, 17) {real, imag} */,
  {32'hbf059ea7, 32'h3ecdd518} /* (22, 16, 16) {real, imag} */,
  {32'h3f7b244a, 32'hbfdb58d2} /* (22, 16, 15) {real, imag} */,
  {32'h3f96061f, 32'h3fad1c8a} /* (22, 16, 14) {real, imag} */,
  {32'h3f6c57f6, 32'hbfa7cf1b} /* (22, 16, 13) {real, imag} */,
  {32'hc0215c85, 32'hbfbe96e7} /* (22, 16, 12) {real, imag} */,
  {32'hbffac8b5, 32'h3d1d1d02} /* (22, 16, 11) {real, imag} */,
  {32'hbf567a52, 32'hbd126c80} /* (22, 16, 10) {real, imag} */,
  {32'h401d9812, 32'h3faa01e4} /* (22, 16, 9) {real, imag} */,
  {32'hbf5fe327, 32'h3ea943df} /* (22, 16, 8) {real, imag} */,
  {32'h3ecba60c, 32'hc07d8069} /* (22, 16, 7) {real, imag} */,
  {32'h3f8f04f7, 32'h3f6922a3} /* (22, 16, 6) {real, imag} */,
  {32'hbf5c280b, 32'hbfabe971} /* (22, 16, 5) {real, imag} */,
  {32'hc017c86f, 32'h3f042e72} /* (22, 16, 4) {real, imag} */,
  {32'hbfe257d7, 32'h3edccd64} /* (22, 16, 3) {real, imag} */,
  {32'h3e2a41c9, 32'h3ed262e0} /* (22, 16, 2) {real, imag} */,
  {32'hbfc66b06, 32'h3ecf27fe} /* (22, 16, 1) {real, imag} */,
  {32'h3fa6465c, 32'hbe7ebe3b} /* (22, 16, 0) {real, imag} */,
  {32'h3e29cc4c, 32'h3dbf4c01} /* (22, 15, 31) {real, imag} */,
  {32'h3d9271fe, 32'h3ff65b52} /* (22, 15, 30) {real, imag} */,
  {32'h3ec9b51b, 32'hbf72936a} /* (22, 15, 29) {real, imag} */,
  {32'hc006cc0f, 32'hc03b7f18} /* (22, 15, 28) {real, imag} */,
  {32'h3e92f5aa, 32'h3f716df4} /* (22, 15, 27) {real, imag} */,
  {32'hbef5ba00, 32'h3fdb33ff} /* (22, 15, 26) {real, imag} */,
  {32'h3ea4589e, 32'h3f16616e} /* (22, 15, 25) {real, imag} */,
  {32'hbe30a7ab, 32'h40191dac} /* (22, 15, 24) {real, imag} */,
  {32'h3e81b543, 32'hbfa6cad3} /* (22, 15, 23) {real, imag} */,
  {32'hc00df91a, 32'hbf9579cc} /* (22, 15, 22) {real, imag} */,
  {32'h3f480a64, 32'hbfbc894f} /* (22, 15, 21) {real, imag} */,
  {32'hbfa194d4, 32'h3eddd8bb} /* (22, 15, 20) {real, imag} */,
  {32'h3f3499b6, 32'hbfbcdd9c} /* (22, 15, 19) {real, imag} */,
  {32'h403a783e, 32'h3edebe5f} /* (22, 15, 18) {real, imag} */,
  {32'h3fc7d358, 32'hbc023cf1} /* (22, 15, 17) {real, imag} */,
  {32'hbe40db98, 32'h3d7e20d5} /* (22, 15, 16) {real, imag} */,
  {32'hbb404c97, 32'hbe1167b8} /* (22, 15, 15) {real, imag} */,
  {32'h3f6313b5, 32'h3fe84148} /* (22, 15, 14) {real, imag} */,
  {32'h3fc1d80d, 32'h40109f03} /* (22, 15, 13) {real, imag} */,
  {32'h3da87f80, 32'hc0300052} /* (22, 15, 12) {real, imag} */,
  {32'hbea924a2, 32'hbe7e72c5} /* (22, 15, 11) {real, imag} */,
  {32'hc019c248, 32'h3f35008c} /* (22, 15, 10) {real, imag} */,
  {32'h4082d8bc, 32'hb906addc} /* (22, 15, 9) {real, imag} */,
  {32'h3fa0af5b, 32'hbfba05b7} /* (22, 15, 8) {real, imag} */,
  {32'h3f1858a7, 32'hbfbcc9cd} /* (22, 15, 7) {real, imag} */,
  {32'h3ee1cddb, 32'hbf5803b9} /* (22, 15, 6) {real, imag} */,
  {32'hbf878d5d, 32'h3f62c8c4} /* (22, 15, 5) {real, imag} */,
  {32'h3ee18ec0, 32'hbec94b8d} /* (22, 15, 4) {real, imag} */,
  {32'hbe8f1427, 32'h3f87f69d} /* (22, 15, 3) {real, imag} */,
  {32'h3f1a3ee2, 32'h40214eb4} /* (22, 15, 2) {real, imag} */,
  {32'hbf3b55b7, 32'hbf3382b4} /* (22, 15, 1) {real, imag} */,
  {32'h3f7396ff, 32'h3e778b79} /* (22, 15, 0) {real, imag} */,
  {32'h4049e850, 32'hbe70ca74} /* (22, 14, 31) {real, imag} */,
  {32'h3d18b048, 32'hbfdfc853} /* (22, 14, 30) {real, imag} */,
  {32'h3f293cc5, 32'h3fb7be48} /* (22, 14, 29) {real, imag} */,
  {32'h3f14825b, 32'hbf73b947} /* (22, 14, 28) {real, imag} */,
  {32'h403ce435, 32'h3f9cd3d1} /* (22, 14, 27) {real, imag} */,
  {32'hbf66100a, 32'hbf8d6b06} /* (22, 14, 26) {real, imag} */,
  {32'h3e58fddd, 32'h3f778d12} /* (22, 14, 25) {real, imag} */,
  {32'h3f96414a, 32'h3f479230} /* (22, 14, 24) {real, imag} */,
  {32'hbfd1e03f, 32'h3f969ed3} /* (22, 14, 23) {real, imag} */,
  {32'h3fb965c9, 32'hc03f5dd6} /* (22, 14, 22) {real, imag} */,
  {32'hbe375c40, 32'h3fac9751} /* (22, 14, 21) {real, imag} */,
  {32'h4053d01f, 32'h40dfbb88} /* (22, 14, 20) {real, imag} */,
  {32'hbff0555c, 32'hbfa97618} /* (22, 14, 19) {real, imag} */,
  {32'h3f89d71b, 32'hbfba489e} /* (22, 14, 18) {real, imag} */,
  {32'hbf93cb52, 32'h3f534a9b} /* (22, 14, 17) {real, imag} */,
  {32'hbed0f266, 32'hbf27bf67} /* (22, 14, 16) {real, imag} */,
  {32'h3f5d6ced, 32'hbf8e23a4} /* (22, 14, 15) {real, imag} */,
  {32'hc04fc6c7, 32'hbf208e8b} /* (22, 14, 14) {real, imag} */,
  {32'h3eaf401c, 32'hbf866adf} /* (22, 14, 13) {real, imag} */,
  {32'hc0264530, 32'hbff712ef} /* (22, 14, 12) {real, imag} */,
  {32'hbfcb1c0e, 32'h3f4871ed} /* (22, 14, 11) {real, imag} */,
  {32'h3fe92726, 32'hc04c156c} /* (22, 14, 10) {real, imag} */,
  {32'h4030ee3e, 32'hbf9f7395} /* (22, 14, 9) {real, imag} */,
  {32'hbd9bead9, 32'hbf700863} /* (22, 14, 8) {real, imag} */,
  {32'h3f9f5090, 32'hbf5426e3} /* (22, 14, 7) {real, imag} */,
  {32'hbf83cb1f, 32'h3ee828d4} /* (22, 14, 6) {real, imag} */,
  {32'h3f971738, 32'hbfa0da58} /* (22, 14, 5) {real, imag} */,
  {32'h3ffd8dd0, 32'h3f8059fb} /* (22, 14, 4) {real, imag} */,
  {32'h3cd74114, 32'h3f29f410} /* (22, 14, 3) {real, imag} */,
  {32'h3e8f5dd1, 32'hc02041b4} /* (22, 14, 2) {real, imag} */,
  {32'hbcefd0ca, 32'h3f159e07} /* (22, 14, 1) {real, imag} */,
  {32'hbf581eb2, 32'h3fff58e1} /* (22, 14, 0) {real, imag} */,
  {32'h3fd1b436, 32'h3bad47d0} /* (22, 13, 31) {real, imag} */,
  {32'h4004b533, 32'hbf8c9bfb} /* (22, 13, 30) {real, imag} */,
  {32'hc01679a6, 32'hbd8613ca} /* (22, 13, 29) {real, imag} */,
  {32'hbfb5b003, 32'h3f7c3998} /* (22, 13, 28) {real, imag} */,
  {32'h3eb633ef, 32'hbc24c657} /* (22, 13, 27) {real, imag} */,
  {32'h40c7f964, 32'h4017dc00} /* (22, 13, 26) {real, imag} */,
  {32'h3fa9aebd, 32'h3fc24924} /* (22, 13, 25) {real, imag} */,
  {32'hbf7f9ad7, 32'hbebec6a3} /* (22, 13, 24) {real, imag} */,
  {32'hc038a006, 32'h3f5dc0fa} /* (22, 13, 23) {real, imag} */,
  {32'h3f97348e, 32'hc041c30b} /* (22, 13, 22) {real, imag} */,
  {32'hbfc58670, 32'h3f9a3360} /* (22, 13, 21) {real, imag} */,
  {32'hbfc6d23b, 32'h3fe8bbfa} /* (22, 13, 20) {real, imag} */,
  {32'h4002d379, 32'hc02cc9c2} /* (22, 13, 19) {real, imag} */,
  {32'h3e9fbf49, 32'hc0956c56} /* (22, 13, 18) {real, imag} */,
  {32'h3f7d290f, 32'hbfb4187e} /* (22, 13, 17) {real, imag} */,
  {32'h40279950, 32'h3fd2ad2d} /* (22, 13, 16) {real, imag} */,
  {32'h4032cb52, 32'h403ede15} /* (22, 13, 15) {real, imag} */,
  {32'h3f65ca62, 32'hc01a6031} /* (22, 13, 14) {real, imag} */,
  {32'hc0076683, 32'hbfb9619c} /* (22, 13, 13) {real, imag} */,
  {32'h3f085158, 32'hbf4d4aad} /* (22, 13, 12) {real, imag} */,
  {32'h3da8b993, 32'h4063cb5f} /* (22, 13, 11) {real, imag} */,
  {32'h4004efad, 32'h4035b7ac} /* (22, 13, 10) {real, imag} */,
  {32'hc00fa76b, 32'h404b008d} /* (22, 13, 9) {real, imag} */,
  {32'h3ed36c62, 32'hbfbc96ce} /* (22, 13, 8) {real, imag} */,
  {32'hc005b1f1, 32'hbfcd42e5} /* (22, 13, 7) {real, imag} */,
  {32'h3fc0f12a, 32'hbeff020a} /* (22, 13, 6) {real, imag} */,
  {32'hc0278752, 32'hc00f7318} /* (22, 13, 5) {real, imag} */,
  {32'h405def47, 32'h3e2613cd} /* (22, 13, 4) {real, imag} */,
  {32'h3fa878ec, 32'h3f6af79f} /* (22, 13, 3) {real, imag} */,
  {32'hbfecc115, 32'hbfc27318} /* (22, 13, 2) {real, imag} */,
  {32'hbee198f9, 32'hbf2fad6a} /* (22, 13, 1) {real, imag} */,
  {32'hbf41e102, 32'h3eb281e8} /* (22, 13, 0) {real, imag} */,
  {32'hbeb1cf46, 32'hc016486b} /* (22, 12, 31) {real, imag} */,
  {32'h3f60f55b, 32'hbe5fdb76} /* (22, 12, 30) {real, imag} */,
  {32'hc01e2492, 32'h3e6bcfd4} /* (22, 12, 29) {real, imag} */,
  {32'hbff22ec3, 32'h40192e0b} /* (22, 12, 28) {real, imag} */,
  {32'h3e2be6a5, 32'h3ccb9f0a} /* (22, 12, 27) {real, imag} */,
  {32'h40411f5d, 32'h40499e5d} /* (22, 12, 26) {real, imag} */,
  {32'hbfe83156, 32'hc01fa420} /* (22, 12, 25) {real, imag} */,
  {32'hbf032cec, 32'hbff44ad0} /* (22, 12, 24) {real, imag} */,
  {32'hbffed559, 32'hbfcc9a1b} /* (22, 12, 23) {real, imag} */,
  {32'hc03ae12a, 32'hbc3674b0} /* (22, 12, 22) {real, imag} */,
  {32'hbff1654a, 32'h3e1dc369} /* (22, 12, 21) {real, imag} */,
  {32'hc0355e83, 32'hc0214ae4} /* (22, 12, 20) {real, imag} */,
  {32'h3fc617bd, 32'h3e6e0644} /* (22, 12, 19) {real, imag} */,
  {32'h405938c7, 32'h40524923} /* (22, 12, 18) {real, imag} */,
  {32'hbf698aa2, 32'hc0004dc4} /* (22, 12, 17) {real, imag} */,
  {32'h40855895, 32'hbe93e847} /* (22, 12, 16) {real, imag} */,
  {32'hbecfc8a7, 32'hbdec02d6} /* (22, 12, 15) {real, imag} */,
  {32'hbfb63731, 32'h3f070cfd} /* (22, 12, 14) {real, imag} */,
  {32'h3e399146, 32'hbfd4d31f} /* (22, 12, 13) {real, imag} */,
  {32'hbffd0adc, 32'hbfd53e06} /* (22, 12, 12) {real, imag} */,
  {32'h3f8b8680, 32'h3fac079f} /* (22, 12, 11) {real, imag} */,
  {32'h3f393125, 32'h3f985e93} /* (22, 12, 10) {real, imag} */,
  {32'h3f23c5af, 32'hbfad035c} /* (22, 12, 9) {real, imag} */,
  {32'h3f825e25, 32'h3f5f90ac} /* (22, 12, 8) {real, imag} */,
  {32'h3fe97042, 32'h4039a65c} /* (22, 12, 7) {real, imag} */,
  {32'hbffb135b, 32'h3fc9daa2} /* (22, 12, 6) {real, imag} */,
  {32'hbe14772a, 32'h3e31e63b} /* (22, 12, 5) {real, imag} */,
  {32'h40118b8e, 32'h3eb41913} /* (22, 12, 4) {real, imag} */,
  {32'hc02e109b, 32'h3fad6aba} /* (22, 12, 3) {real, imag} */,
  {32'h3e0931c2, 32'h3faddf58} /* (22, 12, 2) {real, imag} */,
  {32'h3fba1edb, 32'hbecb8926} /* (22, 12, 1) {real, imag} */,
  {32'h3f2f33c9, 32'hc0013f34} /* (22, 12, 0) {real, imag} */,
  {32'hc02c6858, 32'hbfac2bb7} /* (22, 11, 31) {real, imag} */,
  {32'h3f8551c2, 32'h3f6ed28f} /* (22, 11, 30) {real, imag} */,
  {32'h3f4bf169, 32'h3db14f8f} /* (22, 11, 29) {real, imag} */,
  {32'hbed2ac37, 32'hbf3bc01f} /* (22, 11, 28) {real, imag} */,
  {32'hbfcc823a, 32'hbfecc789} /* (22, 11, 27) {real, imag} */,
  {32'h402f8977, 32'hc06d6c58} /* (22, 11, 26) {real, imag} */,
  {32'h3e186e77, 32'h3f57ab68} /* (22, 11, 25) {real, imag} */,
  {32'hbf462883, 32'hc0729b1f} /* (22, 11, 24) {real, imag} */,
  {32'h40783885, 32'h40437a7f} /* (22, 11, 23) {real, imag} */,
  {32'hbf467d89, 32'hbd508127} /* (22, 11, 22) {real, imag} */,
  {32'h40486c1f, 32'hc01e8334} /* (22, 11, 21) {real, imag} */,
  {32'hc0089143, 32'hbf472ad5} /* (22, 11, 20) {real, imag} */,
  {32'hbd8abfd0, 32'hc05fd6dc} /* (22, 11, 19) {real, imag} */,
  {32'hc04fc2c5, 32'h3f0b5642} /* (22, 11, 18) {real, imag} */,
  {32'h3f62d08e, 32'hbe0b9ab5} /* (22, 11, 17) {real, imag} */,
  {32'h4004f973, 32'hbfe1ad41} /* (22, 11, 16) {real, imag} */,
  {32'hbe36401c, 32'h3fd21a20} /* (22, 11, 15) {real, imag} */,
  {32'hbfdf5837, 32'hbfb088f3} /* (22, 11, 14) {real, imag} */,
  {32'h3fdc4e16, 32'h3feb5bbc} /* (22, 11, 13) {real, imag} */,
  {32'h3fcd9d13, 32'h3f82ff70} /* (22, 11, 12) {real, imag} */,
  {32'h3fb50009, 32'hbe9320f3} /* (22, 11, 11) {real, imag} */,
  {32'hbf7a2442, 32'hc018a46f} /* (22, 11, 10) {real, imag} */,
  {32'hbf5cce10, 32'h3f0ed739} /* (22, 11, 9) {real, imag} */,
  {32'hbf2795db, 32'h3f5691b3} /* (22, 11, 8) {real, imag} */,
  {32'hc02e3672, 32'h4009c9a5} /* (22, 11, 7) {real, imag} */,
  {32'hc04aef3a, 32'h3fb034f2} /* (22, 11, 6) {real, imag} */,
  {32'h3f7983ee, 32'hc07b681e} /* (22, 11, 5) {real, imag} */,
  {32'h3f064acc, 32'h3f73ed4e} /* (22, 11, 4) {real, imag} */,
  {32'h3f1dcf16, 32'hc04c7f11} /* (22, 11, 3) {real, imag} */,
  {32'hbffa4807, 32'h3e18c390} /* (22, 11, 2) {real, imag} */,
  {32'h3e289649, 32'h3f7daa8b} /* (22, 11, 1) {real, imag} */,
  {32'h40284cf8, 32'h3f9a95d5} /* (22, 11, 0) {real, imag} */,
  {32'h3f1446b3, 32'hbe6f2783} /* (22, 10, 31) {real, imag} */,
  {32'hbfbc8167, 32'hc001126b} /* (22, 10, 30) {real, imag} */,
  {32'hbfcf910b, 32'hbfa7517f} /* (22, 10, 29) {real, imag} */,
  {32'h3f9e172f, 32'hbe4de288} /* (22, 10, 28) {real, imag} */,
  {32'h3fb7b64b, 32'h3d4cfbce} /* (22, 10, 27) {real, imag} */,
  {32'hbf1554d7, 32'h3eb1ed69} /* (22, 10, 26) {real, imag} */,
  {32'h3e9ef75f, 32'hbeaab9e9} /* (22, 10, 25) {real, imag} */,
  {32'h3e8dcb9c, 32'h3fb82b5f} /* (22, 10, 24) {real, imag} */,
  {32'h3f589ca3, 32'h3ddef880} /* (22, 10, 23) {real, imag} */,
  {32'h3fafd3d6, 32'h3f36d014} /* (22, 10, 22) {real, imag} */,
  {32'hc03341ba, 32'h3e846ef4} /* (22, 10, 21) {real, imag} */,
  {32'h3eeaf063, 32'h3e6b4b8e} /* (22, 10, 20) {real, imag} */,
  {32'hc0184234, 32'h40840420} /* (22, 10, 19) {real, imag} */,
  {32'hbfad264a, 32'h3f3f5147} /* (22, 10, 18) {real, imag} */,
  {32'hbf5824ad, 32'h3f93c94c} /* (22, 10, 17) {real, imag} */,
  {32'hbed74ce8, 32'h3f6f29e2} /* (22, 10, 16) {real, imag} */,
  {32'h3e75c05d, 32'hc0091486} /* (22, 10, 15) {real, imag} */,
  {32'h3ffa4b8b, 32'h3f5d6290} /* (22, 10, 14) {real, imag} */,
  {32'hc0574f0c, 32'hbf13622e} /* (22, 10, 13) {real, imag} */,
  {32'hc0280541, 32'h3e8d4310} /* (22, 10, 12) {real, imag} */,
  {32'h3e6a0c74, 32'h3f165948} /* (22, 10, 11) {real, imag} */,
  {32'h3f6cee8a, 32'h40431901} /* (22, 10, 10) {real, imag} */,
  {32'hbfd638d1, 32'hbe060543} /* (22, 10, 9) {real, imag} */,
  {32'hbfb721df, 32'h4020f597} /* (22, 10, 8) {real, imag} */,
  {32'h3f659cb2, 32'hc0136d25} /* (22, 10, 7) {real, imag} */,
  {32'hbfffbaee, 32'h40717755} /* (22, 10, 6) {real, imag} */,
  {32'h3ecacabb, 32'h407770ce} /* (22, 10, 5) {real, imag} */,
  {32'h3f27ca0b, 32'hbff4a8cc} /* (22, 10, 4) {real, imag} */,
  {32'hbfce7db2, 32'hbe3409f7} /* (22, 10, 3) {real, imag} */,
  {32'h3f7f7917, 32'h3fae51b5} /* (22, 10, 2) {real, imag} */,
  {32'hbf9b5e24, 32'hbf857338} /* (22, 10, 1) {real, imag} */,
  {32'h3f63ceb4, 32'h401deaee} /* (22, 10, 0) {real, imag} */,
  {32'h3fbc5356, 32'h3f3fbf18} /* (22, 9, 31) {real, imag} */,
  {32'h40049cdd, 32'h40281c63} /* (22, 9, 30) {real, imag} */,
  {32'h3e6f3c23, 32'hc0057e98} /* (22, 9, 29) {real, imag} */,
  {32'h4032cc08, 32'h3e3adfa5} /* (22, 9, 28) {real, imag} */,
  {32'hbf4e52bc, 32'hbfdece17} /* (22, 9, 27) {real, imag} */,
  {32'hbfd9d52f, 32'h40216461} /* (22, 9, 26) {real, imag} */,
  {32'hc038d2a0, 32'hbfc19686} /* (22, 9, 25) {real, imag} */,
  {32'h3ec6ecbf, 32'h3fe72567} /* (22, 9, 24) {real, imag} */,
  {32'h401db943, 32'h3f4b79a5} /* (22, 9, 23) {real, imag} */,
  {32'hc02be764, 32'h3f3d098f} /* (22, 9, 22) {real, imag} */,
  {32'hc00e7109, 32'hc0128e3d} /* (22, 9, 21) {real, imag} */,
  {32'h40627641, 32'h3f073753} /* (22, 9, 20) {real, imag} */,
  {32'h3fe9f564, 32'h406a2feb} /* (22, 9, 19) {real, imag} */,
  {32'hbf86b1df, 32'h3f3f27f9} /* (22, 9, 18) {real, imag} */,
  {32'h3f71cc1d, 32'h3f9ba667} /* (22, 9, 17) {real, imag} */,
  {32'h3f909ec4, 32'hbfb196e3} /* (22, 9, 16) {real, imag} */,
  {32'h3fde932e, 32'hbf9aacc3} /* (22, 9, 15) {real, imag} */,
  {32'h40527cca, 32'h3db99568} /* (22, 9, 14) {real, imag} */,
  {32'hbf12ccb4, 32'hbe1f9681} /* (22, 9, 13) {real, imag} */,
  {32'h3fa0d68d, 32'h4099973f} /* (22, 9, 12) {real, imag} */,
  {32'h406342ba, 32'h3e39049e} /* (22, 9, 11) {real, imag} */,
  {32'h3fab9a44, 32'hc03400c9} /* (22, 9, 10) {real, imag} */,
  {32'hc098fc29, 32'hbc984f8d} /* (22, 9, 9) {real, imag} */,
  {32'hbed54421, 32'hbf425120} /* (22, 9, 8) {real, imag} */,
  {32'h3f6f1d77, 32'h3ffab64e} /* (22, 9, 7) {real, imag} */,
  {32'h403ebf20, 32'h3ea05656} /* (22, 9, 6) {real, imag} */,
  {32'hbfb78c08, 32'h40056b7a} /* (22, 9, 5) {real, imag} */,
  {32'hbfd83886, 32'h3fc4f66b} /* (22, 9, 4) {real, imag} */,
  {32'h3f8f0003, 32'hbf9fd23d} /* (22, 9, 3) {real, imag} */,
  {32'hc00c5e34, 32'hbf55ac02} /* (22, 9, 2) {real, imag} */,
  {32'h3e8da07c, 32'hc02dc880} /* (22, 9, 1) {real, imag} */,
  {32'hbdc5d7b9, 32'h3f21c875} /* (22, 9, 0) {real, imag} */,
  {32'hbdb00ea5, 32'h3fd8c730} /* (22, 8, 31) {real, imag} */,
  {32'h3efcf2a7, 32'hbf9ff7ac} /* (22, 8, 30) {real, imag} */,
  {32'h3f5945bb, 32'hc048c49a} /* (22, 8, 29) {real, imag} */,
  {32'h3ec7651c, 32'h400e0e19} /* (22, 8, 28) {real, imag} */,
  {32'hbf7960b7, 32'h4015995c} /* (22, 8, 27) {real, imag} */,
  {32'hc0468d62, 32'hc00d91d5} /* (22, 8, 26) {real, imag} */,
  {32'h3c64bf5c, 32'hbf26692d} /* (22, 8, 25) {real, imag} */,
  {32'h3f2d9fcb, 32'h3e585b32} /* (22, 8, 24) {real, imag} */,
  {32'h3ef3ec91, 32'hbf8489f2} /* (22, 8, 23) {real, imag} */,
  {32'hbf2c8826, 32'h3f548123} /* (22, 8, 22) {real, imag} */,
  {32'h3e9effdb, 32'hbe6d104e} /* (22, 8, 21) {real, imag} */,
  {32'hc0900306, 32'hbf8a4afa} /* (22, 8, 20) {real, imag} */,
  {32'hbfb8bdf0, 32'hbf08d211} /* (22, 8, 19) {real, imag} */,
  {32'h3f9379ac, 32'hbe892cd5} /* (22, 8, 18) {real, imag} */,
  {32'hc08740be, 32'h3cd6e610} /* (22, 8, 17) {real, imag} */,
  {32'h3eabfcf1, 32'hbe113f5e} /* (22, 8, 16) {real, imag} */,
  {32'h409c6375, 32'hbf66a685} /* (22, 8, 15) {real, imag} */,
  {32'h3f9c2e17, 32'h3f37798e} /* (22, 8, 14) {real, imag} */,
  {32'hbf048374, 32'h3fc1ad14} /* (22, 8, 13) {real, imag} */,
  {32'h3ffecc15, 32'h40446c0c} /* (22, 8, 12) {real, imag} */,
  {32'hbf04c1c0, 32'h3fcbcfb1} /* (22, 8, 11) {real, imag} */,
  {32'hbfaa4a90, 32'hc01d2aa9} /* (22, 8, 10) {real, imag} */,
  {32'h3f387817, 32'hbfa8c50c} /* (22, 8, 9) {real, imag} */,
  {32'hbf506504, 32'hbd3cf415} /* (22, 8, 8) {real, imag} */,
  {32'hc00a948e, 32'h403d4cf7} /* (22, 8, 7) {real, imag} */,
  {32'hc09d8db0, 32'h3e4bc4b2} /* (22, 8, 6) {real, imag} */,
  {32'h4080d1b7, 32'hc051590c} /* (22, 8, 5) {real, imag} */,
  {32'hbf0b399e, 32'hc004a878} /* (22, 8, 4) {real, imag} */,
  {32'h3f74ec4f, 32'h40588202} /* (22, 8, 3) {real, imag} */,
  {32'hbfb9213d, 32'hbff40c55} /* (22, 8, 2) {real, imag} */,
  {32'h40065e6c, 32'hbf32f4f8} /* (22, 8, 1) {real, imag} */,
  {32'hbe4daabc, 32'hbf1550c8} /* (22, 8, 0) {real, imag} */,
  {32'hbf8a3253, 32'hbf817a42} /* (22, 7, 31) {real, imag} */,
  {32'hbfb12df1, 32'h403e8797} /* (22, 7, 30) {real, imag} */,
  {32'hc0357fb4, 32'h402a2611} /* (22, 7, 29) {real, imag} */,
  {32'h3f9ba783, 32'h3dd45c8e} /* (22, 7, 28) {real, imag} */,
  {32'h4025c10b, 32'h404cf3ee} /* (22, 7, 27) {real, imag} */,
  {32'hc05bac33, 32'h3f49cacb} /* (22, 7, 26) {real, imag} */,
  {32'hbf9dc9b7, 32'hc02a6680} /* (22, 7, 25) {real, imag} */,
  {32'h3f6cfc47, 32'h3f0f2e5f} /* (22, 7, 24) {real, imag} */,
  {32'hbeacb4da, 32'hbf413873} /* (22, 7, 23) {real, imag} */,
  {32'h3f8360ed, 32'h4037b693} /* (22, 7, 22) {real, imag} */,
  {32'hbf85dbf5, 32'hc0057ce3} /* (22, 7, 21) {real, imag} */,
  {32'hbfb7f22f, 32'h3ec4f9d1} /* (22, 7, 20) {real, imag} */,
  {32'hc05a0d57, 32'h3f1bc88e} /* (22, 7, 19) {real, imag} */,
  {32'h3f38b9b1, 32'hbebca950} /* (22, 7, 18) {real, imag} */,
  {32'hbea2ce89, 32'hbd50dd05} /* (22, 7, 17) {real, imag} */,
  {32'hbf95f7c6, 32'h3f45dfa7} /* (22, 7, 16) {real, imag} */,
  {32'h3f096ec4, 32'h4016bc4a} /* (22, 7, 15) {real, imag} */,
  {32'h3e6a7dbe, 32'hc013e6a7} /* (22, 7, 14) {real, imag} */,
  {32'hbfaec064, 32'hbfa5d27c} /* (22, 7, 13) {real, imag} */,
  {32'h3f828bb5, 32'hbf9b66d6} /* (22, 7, 12) {real, imag} */,
  {32'hbfbbb7e7, 32'hbfb41dd4} /* (22, 7, 11) {real, imag} */,
  {32'hc02f1a34, 32'hc028bc69} /* (22, 7, 10) {real, imag} */,
  {32'hbd31ef64, 32'h40503571} /* (22, 7, 9) {real, imag} */,
  {32'hbfc030dc, 32'h3f000bf6} /* (22, 7, 8) {real, imag} */,
  {32'h3e081cab, 32'hc04b11d2} /* (22, 7, 7) {real, imag} */,
  {32'h40508566, 32'h404623a7} /* (22, 7, 6) {real, imag} */,
  {32'h404ca5d4, 32'hbf9a0104} /* (22, 7, 5) {real, imag} */,
  {32'h3e9aaa1e, 32'hbfa61775} /* (22, 7, 4) {real, imag} */,
  {32'h402cf930, 32'h3f51a532} /* (22, 7, 3) {real, imag} */,
  {32'h3f8cd5a2, 32'hbf49a274} /* (22, 7, 2) {real, imag} */,
  {32'h40326d7c, 32'h402f6d2a} /* (22, 7, 1) {real, imag} */,
  {32'hbf8d1d77, 32'hbfb3b0c9} /* (22, 7, 0) {real, imag} */,
  {32'h3f397361, 32'h3eb409fe} /* (22, 6, 31) {real, imag} */,
  {32'h3f071d4b, 32'h3e25a469} /* (22, 6, 30) {real, imag} */,
  {32'h40698d26, 32'hbf0c8199} /* (22, 6, 29) {real, imag} */,
  {32'hc06f6833, 32'hbf348c79} /* (22, 6, 28) {real, imag} */,
  {32'hc02373ee, 32'h406148fa} /* (22, 6, 27) {real, imag} */,
  {32'h3e0bd1a6, 32'hbd88fc34} /* (22, 6, 26) {real, imag} */,
  {32'h406fd052, 32'h4002e2ed} /* (22, 6, 25) {real, imag} */,
  {32'hbf1db47a, 32'hbf6e34b1} /* (22, 6, 24) {real, imag} */,
  {32'hbe51b4d0, 32'hbe9d6422} /* (22, 6, 23) {real, imag} */,
  {32'h3f5f7e72, 32'hbfdb357d} /* (22, 6, 22) {real, imag} */,
  {32'hbdf84f71, 32'hc0350a25} /* (22, 6, 21) {real, imag} */,
  {32'h3ff88123, 32'hbea57da1} /* (22, 6, 20) {real, imag} */,
  {32'h3f948627, 32'hbec4f340} /* (22, 6, 19) {real, imag} */,
  {32'hbee644fc, 32'h3fc059df} /* (22, 6, 18) {real, imag} */,
  {32'hbf98bd38, 32'h3daa34ae} /* (22, 6, 17) {real, imag} */,
  {32'hbeb235c6, 32'h3e8aa72a} /* (22, 6, 16) {real, imag} */,
  {32'h3fe58188, 32'hbee165db} /* (22, 6, 15) {real, imag} */,
  {32'hbf98adf0, 32'hbf15c33d} /* (22, 6, 14) {real, imag} */,
  {32'h408819d9, 32'h3fd8b7eb} /* (22, 6, 13) {real, imag} */,
  {32'h3f6d067b, 32'h4083e350} /* (22, 6, 12) {real, imag} */,
  {32'h3f1a5631, 32'h4030481a} /* (22, 6, 11) {real, imag} */,
  {32'h3fb162ef, 32'hbfd827b6} /* (22, 6, 10) {real, imag} */,
  {32'hbe9ee226, 32'h3efa82b8} /* (22, 6, 9) {real, imag} */,
  {32'h401e7779, 32'hbe68400f} /* (22, 6, 8) {real, imag} */,
  {32'h3f3ac312, 32'h3ecc5d64} /* (22, 6, 7) {real, imag} */,
  {32'h4000f523, 32'hbfce24c7} /* (22, 6, 6) {real, imag} */,
  {32'hc064ec50, 32'h3e858e74} /* (22, 6, 5) {real, imag} */,
  {32'hbeb791e9, 32'hbf608e00} /* (22, 6, 4) {real, imag} */,
  {32'hbe8f7632, 32'hc01ed2b9} /* (22, 6, 3) {real, imag} */,
  {32'hc0491000, 32'h3fe08a85} /* (22, 6, 2) {real, imag} */,
  {32'h3dd4c029, 32'hbf6085f6} /* (22, 6, 1) {real, imag} */,
  {32'h4013fb5f, 32'h4008aeaf} /* (22, 6, 0) {real, imag} */,
  {32'h3f6b758b, 32'hc015c892} /* (22, 5, 31) {real, imag} */,
  {32'h3d77b14c, 32'h3f80008a} /* (22, 5, 30) {real, imag} */,
  {32'h3f410bf0, 32'h4016ba7c} /* (22, 5, 29) {real, imag} */,
  {32'hc088d3e0, 32'h3f177fd7} /* (22, 5, 28) {real, imag} */,
  {32'h405acb1e, 32'h3f811965} /* (22, 5, 27) {real, imag} */,
  {32'h3fbe3b76, 32'hc03f312f} /* (22, 5, 26) {real, imag} */,
  {32'h3f40a913, 32'hbf9d8f26} /* (22, 5, 25) {real, imag} */,
  {32'hbfe06e81, 32'hbf236fdd} /* (22, 5, 24) {real, imag} */,
  {32'hbe5bb8a6, 32'hbf9e3d20} /* (22, 5, 23) {real, imag} */,
  {32'h3f5fea57, 32'h4060811a} /* (22, 5, 22) {real, imag} */,
  {32'h3f46c98e, 32'h3fb33a22} /* (22, 5, 21) {real, imag} */,
  {32'hbf041381, 32'h3fef5042} /* (22, 5, 20) {real, imag} */,
  {32'h3ef8fda0, 32'hbea71679} /* (22, 5, 19) {real, imag} */,
  {32'h402f1d55, 32'h3e4c1d49} /* (22, 5, 18) {real, imag} */,
  {32'h3eef720e, 32'h3c6c98f0} /* (22, 5, 17) {real, imag} */,
  {32'hc0176176, 32'hbf308956} /* (22, 5, 16) {real, imag} */,
  {32'hbe4abd5c, 32'hbf0acda9} /* (22, 5, 15) {real, imag} */,
  {32'h3f5d7d9d, 32'hbf8e4841} /* (22, 5, 14) {real, imag} */,
  {32'hbe62d1f7, 32'hbf2eb232} /* (22, 5, 13) {real, imag} */,
  {32'h3eec3a8f, 32'hbf79a45c} /* (22, 5, 12) {real, imag} */,
  {32'h400a9e51, 32'h3f579f57} /* (22, 5, 11) {real, imag} */,
  {32'hc0306c38, 32'hbeae15ec} /* (22, 5, 10) {real, imag} */,
  {32'h3fa8a679, 32'h3fd5c8b7} /* (22, 5, 9) {real, imag} */,
  {32'hbdb5f954, 32'h3eca823a} /* (22, 5, 8) {real, imag} */,
  {32'hbecd0a1f, 32'hbfd1c069} /* (22, 5, 7) {real, imag} */,
  {32'hbfb910e7, 32'h40022ac0} /* (22, 5, 6) {real, imag} */,
  {32'h3edfb491, 32'hc00ea6f3} /* (22, 5, 5) {real, imag} */,
  {32'h400d5673, 32'h4026498f} /* (22, 5, 4) {real, imag} */,
  {32'hc02d98e7, 32'h3fe97d78} /* (22, 5, 3) {real, imag} */,
  {32'hbfc08945, 32'hbeb651a0} /* (22, 5, 2) {real, imag} */,
  {32'hbffc1429, 32'h3ead76cd} /* (22, 5, 1) {real, imag} */,
  {32'h3fec85d7, 32'hbfd20dd2} /* (22, 5, 0) {real, imag} */,
  {32'h3fb931e5, 32'h3f5e7b61} /* (22, 4, 31) {real, imag} */,
  {32'h3e7a1e6e, 32'h401b86c2} /* (22, 4, 30) {real, imag} */,
  {32'hc00ff585, 32'h4026c586} /* (22, 4, 29) {real, imag} */,
  {32'h3e1d061d, 32'hc04c3cc1} /* (22, 4, 28) {real, imag} */,
  {32'hbf9fadd5, 32'h3f407440} /* (22, 4, 27) {real, imag} */,
  {32'hc05fd663, 32'hc075e57b} /* (22, 4, 26) {real, imag} */,
  {32'h3fc2bacc, 32'hbfbcd10c} /* (22, 4, 25) {real, imag} */,
  {32'h3fa9a75f, 32'h3e326ae0} /* (22, 4, 24) {real, imag} */,
  {32'hc016f291, 32'h3f341bee} /* (22, 4, 23) {real, imag} */,
  {32'hbe4e324a, 32'h402d3aa5} /* (22, 4, 22) {real, imag} */,
  {32'h40858f03, 32'h3ea27e98} /* (22, 4, 21) {real, imag} */,
  {32'hc0b7a8dd, 32'hc042cf8c} /* (22, 4, 20) {real, imag} */,
  {32'h3fb5ec17, 32'hbe6cdbf6} /* (22, 4, 19) {real, imag} */,
  {32'hbfbf7357, 32'hbf88dfd4} /* (22, 4, 18) {real, imag} */,
  {32'h3f84c619, 32'hbfc3cf03} /* (22, 4, 17) {real, imag} */,
  {32'hbf6fd324, 32'h3f0d8995} /* (22, 4, 16) {real, imag} */,
  {32'h3f58589e, 32'h3eb491c0} /* (22, 4, 15) {real, imag} */,
  {32'hbfe636c9, 32'hbf946642} /* (22, 4, 14) {real, imag} */,
  {32'h3f788fef, 32'hbf472f31} /* (22, 4, 13) {real, imag} */,
  {32'hbfafed0e, 32'h3f6a6340} /* (22, 4, 12) {real, imag} */,
  {32'h3ed525d2, 32'hbf87e1d2} /* (22, 4, 11) {real, imag} */,
  {32'h3cb0e54b, 32'h40013807} /* (22, 4, 10) {real, imag} */,
  {32'h3d995478, 32'h3fe9edd7} /* (22, 4, 9) {real, imag} */,
  {32'h40088c8e, 32'hbf9ed6e7} /* (22, 4, 8) {real, imag} */,
  {32'h3ff293fa, 32'hc002a851} /* (22, 4, 7) {real, imag} */,
  {32'hbd2d543b, 32'h3de1cfec} /* (22, 4, 6) {real, imag} */,
  {32'h3e60aeea, 32'h400442e0} /* (22, 4, 5) {real, imag} */,
  {32'hc0cd905f, 32'hbdc77034} /* (22, 4, 4) {real, imag} */,
  {32'h3d37a4be, 32'hbf6e666d} /* (22, 4, 3) {real, imag} */,
  {32'hbff0782d, 32'h4035e3dd} /* (22, 4, 2) {real, imag} */,
  {32'h3f62f05e, 32'hc001cebd} /* (22, 4, 1) {real, imag} */,
  {32'hbf016d31, 32'hbfd061ae} /* (22, 4, 0) {real, imag} */,
  {32'hc07375bd, 32'h40082344} /* (22, 3, 31) {real, imag} */,
  {32'hbf9ccab7, 32'h406b367b} /* (22, 3, 30) {real, imag} */,
  {32'hbe850959, 32'hbf550c50} /* (22, 3, 29) {real, imag} */,
  {32'h3fc6018c, 32'h3f8030fb} /* (22, 3, 28) {real, imag} */,
  {32'h3fb19bb3, 32'h3ffd024c} /* (22, 3, 27) {real, imag} */,
  {32'h3e92e248, 32'hbf87c10c} /* (22, 3, 26) {real, imag} */,
  {32'hbeca9f7f, 32'hbf616e66} /* (22, 3, 25) {real, imag} */,
  {32'h3eb4d0cb, 32'hc0940932} /* (22, 3, 24) {real, imag} */,
  {32'h3fba375b, 32'hbe4f4b7f} /* (22, 3, 23) {real, imag} */,
  {32'hc0770bcf, 32'hbfc7273e} /* (22, 3, 22) {real, imag} */,
  {32'hbfafb3d4, 32'hbf2317e7} /* (22, 3, 21) {real, imag} */,
  {32'h3f27e388, 32'hc0314a14} /* (22, 3, 20) {real, imag} */,
  {32'hbf1f313d, 32'hbf985513} /* (22, 3, 19) {real, imag} */,
  {32'hbf690c39, 32'hc0428a0a} /* (22, 3, 18) {real, imag} */,
  {32'h3cc754c5, 32'h3f85e220} /* (22, 3, 17) {real, imag} */,
  {32'h3fce048d, 32'h3fae0ffa} /* (22, 3, 16) {real, imag} */,
  {32'h3f497730, 32'hbf0c3f0c} /* (22, 3, 15) {real, imag} */,
  {32'hbf82c2a6, 32'h40255835} /* (22, 3, 14) {real, imag} */,
  {32'hbfabe1bf, 32'h3f1dfbd2} /* (22, 3, 13) {real, imag} */,
  {32'h40491993, 32'h3ec9e3a5} /* (22, 3, 12) {real, imag} */,
  {32'hbfb826c0, 32'h3f13d9c4} /* (22, 3, 11) {real, imag} */,
  {32'hbe336dc2, 32'h3f73b12c} /* (22, 3, 10) {real, imag} */,
  {32'h3fba1fd4, 32'hbfa70a26} /* (22, 3, 9) {real, imag} */,
  {32'hbf82d697, 32'h3f033314} /* (22, 3, 8) {real, imag} */,
  {32'hbfbfffda, 32'h3f48f322} /* (22, 3, 7) {real, imag} */,
  {32'h3f3b97f5, 32'hc07cdf92} /* (22, 3, 6) {real, imag} */,
  {32'hbfb327da, 32'hc0619aef} /* (22, 3, 5) {real, imag} */,
  {32'hbf548813, 32'hbebcd1f8} /* (22, 3, 4) {real, imag} */,
  {32'hc0008451, 32'h3e31621a} /* (22, 3, 3) {real, imag} */,
  {32'hbf3bb982, 32'h3ffbd3dd} /* (22, 3, 2) {real, imag} */,
  {32'hc0265a76, 32'h40100153} /* (22, 3, 1) {real, imag} */,
  {32'hc0203052, 32'h40630c80} /* (22, 3, 0) {real, imag} */,
  {32'h40190bd2, 32'h405497a5} /* (22, 2, 31) {real, imag} */,
  {32'hbeb20184, 32'h3f023292} /* (22, 2, 30) {real, imag} */,
  {32'h407fe443, 32'h3e68f325} /* (22, 2, 29) {real, imag} */,
  {32'h3f26aca7, 32'hc0e30dec} /* (22, 2, 28) {real, imag} */,
  {32'hbe534921, 32'hc01d1651} /* (22, 2, 27) {real, imag} */,
  {32'h3faf83a3, 32'h3fdcdee8} /* (22, 2, 26) {real, imag} */,
  {32'hbed8a7a5, 32'hbfebd391} /* (22, 2, 25) {real, imag} */,
  {32'hc03e9bbc, 32'hbfae29da} /* (22, 2, 24) {real, imag} */,
  {32'hbfe32c25, 32'h3e0de28a} /* (22, 2, 23) {real, imag} */,
  {32'h3e8c3f7f, 32'hbee8ec53} /* (22, 2, 22) {real, imag} */,
  {32'hbee5f106, 32'h3e72ec1b} /* (22, 2, 21) {real, imag} */,
  {32'hbfd395ae, 32'h402dd145} /* (22, 2, 20) {real, imag} */,
  {32'h3f30f373, 32'h3f936f36} /* (22, 2, 19) {real, imag} */,
  {32'h3f9cc296, 32'h40221db0} /* (22, 2, 18) {real, imag} */,
  {32'hbf72d12c, 32'h3eeebef3} /* (22, 2, 17) {real, imag} */,
  {32'h3edb7423, 32'hbc9fcb79} /* (22, 2, 16) {real, imag} */,
  {32'h3e9b55a8, 32'h3f2c35de} /* (22, 2, 15) {real, imag} */,
  {32'h4036106b, 32'hc00bcfd9} /* (22, 2, 14) {real, imag} */,
  {32'h3f1bc4a8, 32'hc0169f12} /* (22, 2, 13) {real, imag} */,
  {32'hbfc51771, 32'hbff47655} /* (22, 2, 12) {real, imag} */,
  {32'hbe078c0c, 32'h3f88ba3f} /* (22, 2, 11) {real, imag} */,
  {32'hbf73b0fa, 32'h40178c83} /* (22, 2, 10) {real, imag} */,
  {32'hbfb45ca7, 32'hbf8587dd} /* (22, 2, 9) {real, imag} */,
  {32'hc0077c8d, 32'hc08af7c0} /* (22, 2, 8) {real, imag} */,
  {32'h3ea4010a, 32'h4039901d} /* (22, 2, 7) {real, imag} */,
  {32'h3ea11706, 32'hbf815475} /* (22, 2, 6) {real, imag} */,
  {32'hc04b0a80, 32'hbfdb78e7} /* (22, 2, 5) {real, imag} */,
  {32'h3eb77618, 32'h4011790c} /* (22, 2, 4) {real, imag} */,
  {32'hbefd11a0, 32'h4057060c} /* (22, 2, 3) {real, imag} */,
  {32'hc0bfd73a, 32'h3e831296} /* (22, 2, 2) {real, imag} */,
  {32'h3f9ae4e7, 32'hc0323dc3} /* (22, 2, 1) {real, imag} */,
  {32'h40acaeb1, 32'h3f8fbba7} /* (22, 2, 0) {real, imag} */,
  {32'hc0583de1, 32'hbfc3d800} /* (22, 1, 31) {real, imag} */,
  {32'h4027ba79, 32'h407333e0} /* (22, 1, 30) {real, imag} */,
  {32'h3f85465d, 32'hc066cbb6} /* (22, 1, 29) {real, imag} */,
  {32'hbfc19935, 32'hbcda9c06} /* (22, 1, 28) {real, imag} */,
  {32'hbf6fb7af, 32'h40c83fdd} /* (22, 1, 27) {real, imag} */,
  {32'hbf633628, 32'h3ff832b8} /* (22, 1, 26) {real, imag} */,
  {32'hbf8e2b40, 32'hbfd1edb7} /* (22, 1, 25) {real, imag} */,
  {32'hbec60bcd, 32'h402f71d8} /* (22, 1, 24) {real, imag} */,
  {32'h3f4eb966, 32'hbec22ad4} /* (22, 1, 23) {real, imag} */,
  {32'h3fcebf8d, 32'h3fa89fce} /* (22, 1, 22) {real, imag} */,
  {32'h3f18caf5, 32'hbf0d0c41} /* (22, 1, 21) {real, imag} */,
  {32'h3e05a053, 32'h3f0b269a} /* (22, 1, 20) {real, imag} */,
  {32'h4012fa9e, 32'h40447a5b} /* (22, 1, 19) {real, imag} */,
  {32'hbf14df8e, 32'hbf2dc6c0} /* (22, 1, 18) {real, imag} */,
  {32'hbf6814f4, 32'hbfdf62da} /* (22, 1, 17) {real, imag} */,
  {32'h3f14caa0, 32'h3e1a9b5a} /* (22, 1, 16) {real, imag} */,
  {32'h3f8a9f7a, 32'h3f60c0bf} /* (22, 1, 15) {real, imag} */,
  {32'hbf9bd7c2, 32'hbf5d377f} /* (22, 1, 14) {real, imag} */,
  {32'hbf2fbc7e, 32'hbedd5b5f} /* (22, 1, 13) {real, imag} */,
  {32'hbfa9e635, 32'hbdde5f4b} /* (22, 1, 12) {real, imag} */,
  {32'h3f04dc08, 32'hbfe5ee1f} /* (22, 1, 11) {real, imag} */,
  {32'h3ef81ffa, 32'h3fd93b90} /* (22, 1, 10) {real, imag} */,
  {32'hc06080df, 32'hbf9d9471} /* (22, 1, 9) {real, imag} */,
  {32'hbf6a9a19, 32'hbfb404c2} /* (22, 1, 8) {real, imag} */,
  {32'h3eaa8ff9, 32'hc08c971f} /* (22, 1, 7) {real, imag} */,
  {32'h3fcf82f2, 32'h3fa7ebfa} /* (22, 1, 6) {real, imag} */,
  {32'h40af2bc6, 32'h3fdcc56d} /* (22, 1, 5) {real, imag} */,
  {32'hbfcc9ff5, 32'hbf1cd8cb} /* (22, 1, 4) {real, imag} */,
  {32'h40a1adbe, 32'h3c738e87} /* (22, 1, 3) {real, imag} */,
  {32'h3f905a44, 32'h40568bca} /* (22, 1, 2) {real, imag} */,
  {32'hc013519c, 32'hc09d3234} /* (22, 1, 1) {real, imag} */,
  {32'h4011481f, 32'hc0aff7c3} /* (22, 1, 0) {real, imag} */,
  {32'hc06c4dbd, 32'h40690ed4} /* (22, 0, 31) {real, imag} */,
  {32'h3fe19ba9, 32'h4041b0e9} /* (22, 0, 30) {real, imag} */,
  {32'hc0a20d8b, 32'h3e95d545} /* (22, 0, 29) {real, imag} */,
  {32'hbec3296a, 32'hbcdea6b0} /* (22, 0, 28) {real, imag} */,
  {32'hbf76bfa4, 32'hc022768b} /* (22, 0, 27) {real, imag} */,
  {32'h3eeb14b2, 32'hbe30681d} /* (22, 0, 26) {real, imag} */,
  {32'hc0020cfb, 32'hc06247bd} /* (22, 0, 25) {real, imag} */,
  {32'hc06e9456, 32'hbffc3910} /* (22, 0, 24) {real, imag} */,
  {32'h404915c8, 32'hc03db2fe} /* (22, 0, 23) {real, imag} */,
  {32'hbea95f87, 32'hbedb4452} /* (22, 0, 22) {real, imag} */,
  {32'hbe40b3cb, 32'h403ad638} /* (22, 0, 21) {real, imag} */,
  {32'h3e9c74e4, 32'h3faf3677} /* (22, 0, 20) {real, imag} */,
  {32'h3eae4200, 32'hc02339b0} /* (22, 0, 19) {real, imag} */,
  {32'hbf1740a7, 32'h3fbdc252} /* (22, 0, 18) {real, imag} */,
  {32'h3f678b61, 32'hbf5e8391} /* (22, 0, 17) {real, imag} */,
  {32'h3fc00d36, 32'hc044a113} /* (22, 0, 16) {real, imag} */,
  {32'h3f07571a, 32'h3fe5bd17} /* (22, 0, 15) {real, imag} */,
  {32'hbf33dc51, 32'h3ea843ae} /* (22, 0, 14) {real, imag} */,
  {32'hbfd6e878, 32'h400ad271} /* (22, 0, 13) {real, imag} */,
  {32'h401b723c, 32'hbeee5e66} /* (22, 0, 12) {real, imag} */,
  {32'h40051461, 32'h3fb514d9} /* (22, 0, 11) {real, imag} */,
  {32'hbf575956, 32'hbfd5904c} /* (22, 0, 10) {real, imag} */,
  {32'h40997dc7, 32'h3f1999ef} /* (22, 0, 9) {real, imag} */,
  {32'hbf3dda03, 32'hbf72551b} /* (22, 0, 8) {real, imag} */,
  {32'h3f8ef49a, 32'h3f4fe837} /* (22, 0, 7) {real, imag} */,
  {32'hc0149a7a, 32'h409bd375} /* (22, 0, 6) {real, imag} */,
  {32'h40d4245e, 32'h402a3fa4} /* (22, 0, 5) {real, imag} */,
  {32'h4063d4b2, 32'h4085e23c} /* (22, 0, 4) {real, imag} */,
  {32'hc03437b5, 32'h3ff36dd0} /* (22, 0, 3) {real, imag} */,
  {32'hbe5d3967, 32'h3f70e9d7} /* (22, 0, 2) {real, imag} */,
  {32'hbfbcbd1b, 32'hbf806b45} /* (22, 0, 1) {real, imag} */,
  {32'hbfa85644, 32'h3fa639ca} /* (22, 0, 0) {real, imag} */,
  {32'h41206b4f, 32'hbf84d39a} /* (21, 31, 31) {real, imag} */,
  {32'hc0e4c1a5, 32'h4007de89} /* (21, 31, 30) {real, imag} */,
  {32'h40181de8, 32'hbf53cb6b} /* (21, 31, 29) {real, imag} */,
  {32'h3fad4cf9, 32'hbfd64ac0} /* (21, 31, 28) {real, imag} */,
  {32'hc03890c4, 32'hbfa3ab52} /* (21, 31, 27) {real, imag} */,
  {32'h403aeecb, 32'h3f314612} /* (21, 31, 26) {real, imag} */,
  {32'hbfcb21e5, 32'h3f9db62c} /* (21, 31, 25) {real, imag} */,
  {32'hc082ae66, 32'hbffd345c} /* (21, 31, 24) {real, imag} */,
  {32'h4028900f, 32'h3f9fb47f} /* (21, 31, 23) {real, imag} */,
  {32'hbd811423, 32'hbf35fce1} /* (21, 31, 22) {real, imag} */,
  {32'hbfc61399, 32'h3e4aa935} /* (21, 31, 21) {real, imag} */,
  {32'hbe924442, 32'hbfc1bf1c} /* (21, 31, 20) {real, imag} */,
  {32'h3fbd872e, 32'h3f39e714} /* (21, 31, 19) {real, imag} */,
  {32'h4088fc43, 32'h3fe744ed} /* (21, 31, 18) {real, imag} */,
  {32'hbe59249e, 32'hbff5abbf} /* (21, 31, 17) {real, imag} */,
  {32'hbee7ce01, 32'h3f847826} /* (21, 31, 16) {real, imag} */,
  {32'h4036ae06, 32'h4007aae6} /* (21, 31, 15) {real, imag} */,
  {32'hbe3a74ac, 32'h3e58d53e} /* (21, 31, 14) {real, imag} */,
  {32'h3f295fbb, 32'h402911ac} /* (21, 31, 13) {real, imag} */,
  {32'h3f5475ea, 32'hc053aaa0} /* (21, 31, 12) {real, imag} */,
  {32'hbef461d7, 32'h3f100575} /* (21, 31, 11) {real, imag} */,
  {32'hbf040ed4, 32'h3ffda74e} /* (21, 31, 10) {real, imag} */,
  {32'hbe8a4378, 32'h3f5afe45} /* (21, 31, 9) {real, imag} */,
  {32'h3fad385e, 32'h40970be0} /* (21, 31, 8) {real, imag} */,
  {32'hbf53e957, 32'h40161357} /* (21, 31, 7) {real, imag} */,
  {32'hc01862f6, 32'hbf18e742} /* (21, 31, 6) {real, imag} */,
  {32'hc0a27ac4, 32'hc014f00f} /* (21, 31, 5) {real, imag} */,
  {32'h4000925a, 32'hc09c0f50} /* (21, 31, 4) {real, imag} */,
  {32'hbec2c814, 32'hbfe25dd3} /* (21, 31, 3) {real, imag} */,
  {32'hc088c9c8, 32'h3ed34f0a} /* (21, 31, 2) {real, imag} */,
  {32'h3fab1fcf, 32'h40545e40} /* (21, 31, 1) {real, imag} */,
  {32'h40cae1a2, 32'h3fa40baf} /* (21, 31, 0) {real, imag} */,
  {32'hbfd1a6c7, 32'hbf93fad1} /* (21, 30, 31) {real, imag} */,
  {32'h3f2fffd1, 32'h40a8d90f} /* (21, 30, 30) {real, imag} */,
  {32'hbf7e50f4, 32'h3d42d83d} /* (21, 30, 29) {real, imag} */,
  {32'hc002089d, 32'h3fbaa0e6} /* (21, 30, 28) {real, imag} */,
  {32'h40123ea6, 32'hbf065393} /* (21, 30, 27) {real, imag} */,
  {32'h3f6ed9a5, 32'h3fffe64e} /* (21, 30, 26) {real, imag} */,
  {32'h3fa78bfe, 32'hbfa8204b} /* (21, 30, 25) {real, imag} */,
  {32'hbf97f716, 32'hc066934f} /* (21, 30, 24) {real, imag} */,
  {32'hc0068ea7, 32'h402902c6} /* (21, 30, 23) {real, imag} */,
  {32'hc09f8aaf, 32'h3f031d29} /* (21, 30, 22) {real, imag} */,
  {32'h4000917d, 32'hc0453c17} /* (21, 30, 21) {real, imag} */,
  {32'h40932071, 32'hbe508b69} /* (21, 30, 20) {real, imag} */,
  {32'hbfdea654, 32'h3f1a3f8d} /* (21, 30, 19) {real, imag} */,
  {32'hbff81028, 32'h3eb58d4c} /* (21, 30, 18) {real, imag} */,
  {32'h3f587d0c, 32'h40399f35} /* (21, 30, 17) {real, imag} */,
  {32'h3b35d331, 32'hbf507b76} /* (21, 30, 16) {real, imag} */,
  {32'hbec11458, 32'hc0140693} /* (21, 30, 15) {real, imag} */,
  {32'hbf67c6ef, 32'hbe7738a4} /* (21, 30, 14) {real, imag} */,
  {32'h3fe3ffd1, 32'hbef5a885} /* (21, 30, 13) {real, imag} */,
  {32'hbf9e6b0e, 32'hc00775bd} /* (21, 30, 12) {real, imag} */,
  {32'h3e82da76, 32'h3f86a30c} /* (21, 30, 11) {real, imag} */,
  {32'h3ed6a724, 32'hbf9c9315} /* (21, 30, 10) {real, imag} */,
  {32'h403cda25, 32'hbe546a10} /* (21, 30, 9) {real, imag} */,
  {32'h3f07fbcc, 32'h40684a1d} /* (21, 30, 8) {real, imag} */,
  {32'hc03127cb, 32'hc09558ca} /* (21, 30, 7) {real, imag} */,
  {32'h3f351b61, 32'hc0057ebe} /* (21, 30, 6) {real, imag} */,
  {32'hbe3b92bd, 32'hbf3c4d6c} /* (21, 30, 5) {real, imag} */,
  {32'h3f127a9c, 32'h3e51d806} /* (21, 30, 4) {real, imag} */,
  {32'h3e8db507, 32'h3d133e04} /* (21, 30, 3) {real, imag} */,
  {32'h40cfdbd2, 32'h3eb9a1f9} /* (21, 30, 2) {real, imag} */,
  {32'hc0dde7e2, 32'hc0774c7a} /* (21, 30, 1) {real, imag} */,
  {32'hc064d99f, 32'hbe60e8f7} /* (21, 30, 0) {real, imag} */,
  {32'hbf7ca812, 32'hbfe1b321} /* (21, 29, 31) {real, imag} */,
  {32'hc07d042f, 32'h3e05ac81} /* (21, 29, 30) {real, imag} */,
  {32'hc04d6430, 32'h3fd8c081} /* (21, 29, 29) {real, imag} */,
  {32'hbf909028, 32'hbf83286b} /* (21, 29, 28) {real, imag} */,
  {32'hbf3589ff, 32'h3f629589} /* (21, 29, 27) {real, imag} */,
  {32'h3f6d054c, 32'h3f90c87e} /* (21, 29, 26) {real, imag} */,
  {32'h3f904625, 32'hbe1476d5} /* (21, 29, 25) {real, imag} */,
  {32'hbf8a6b1b, 32'hc02b442e} /* (21, 29, 24) {real, imag} */,
  {32'h4060cba1, 32'h3f3e06b3} /* (21, 29, 23) {real, imag} */,
  {32'hbff439ea, 32'h3e8d5878} /* (21, 29, 22) {real, imag} */,
  {32'h3ff24116, 32'hc012f167} /* (21, 29, 21) {real, imag} */,
  {32'hbfad19d0, 32'hc014b63f} /* (21, 29, 20) {real, imag} */,
  {32'h3fa11eb7, 32'h3f480516} /* (21, 29, 19) {real, imag} */,
  {32'h3ff6f097, 32'hbfb01e9f} /* (21, 29, 18) {real, imag} */,
  {32'hbf73b350, 32'h3f86d639} /* (21, 29, 17) {real, imag} */,
  {32'hc01192f5, 32'h3f0e3d21} /* (21, 29, 16) {real, imag} */,
  {32'h3f092744, 32'hbfab6932} /* (21, 29, 15) {real, imag} */,
  {32'hbfadb0b0, 32'hbf937ceb} /* (21, 29, 14) {real, imag} */,
  {32'hbfa3834d, 32'h3ebfe63a} /* (21, 29, 13) {real, imag} */,
  {32'hbfa057bd, 32'hc0857f6b} /* (21, 29, 12) {real, imag} */,
  {32'hc03c1de5, 32'h3f42eb9e} /* (21, 29, 11) {real, imag} */,
  {32'hc002f4ef, 32'h3f6397eb} /* (21, 29, 10) {real, imag} */,
  {32'h403063af, 32'h3fcbc745} /* (21, 29, 9) {real, imag} */,
  {32'hbe8ea97c, 32'h3ffe52ea} /* (21, 29, 8) {real, imag} */,
  {32'hbfedf34a, 32'h405bd519} /* (21, 29, 7) {real, imag} */,
  {32'hc0042671, 32'hc013c982} /* (21, 29, 6) {real, imag} */,
  {32'h3f9f362b, 32'h40909ae0} /* (21, 29, 5) {real, imag} */,
  {32'h3ff69c34, 32'h3fa54b53} /* (21, 29, 4) {real, imag} */,
  {32'h400a63c3, 32'hbfc65da5} /* (21, 29, 3) {real, imag} */,
  {32'hbf558be6, 32'h40905791} /* (21, 29, 2) {real, imag} */,
  {32'h3fb54741, 32'hc07c8032} /* (21, 29, 1) {real, imag} */,
  {32'h405f37f9, 32'hbfc8fa33} /* (21, 29, 0) {real, imag} */,
  {32'h4098d628, 32'hbd8ca88c} /* (21, 28, 31) {real, imag} */,
  {32'hc064cefb, 32'h40972fb3} /* (21, 28, 30) {real, imag} */,
  {32'h405abfbf, 32'h3f9e813b} /* (21, 28, 29) {real, imag} */,
  {32'h3f43eb6a, 32'hbff3cc68} /* (21, 28, 28) {real, imag} */,
  {32'hc01e8834, 32'hbfa777b0} /* (21, 28, 27) {real, imag} */,
  {32'hc066ff14, 32'hc017c864} /* (21, 28, 26) {real, imag} */,
  {32'h40862ecc, 32'h4019cad0} /* (21, 28, 25) {real, imag} */,
  {32'hbea0b66d, 32'h3f87dece} /* (21, 28, 24) {real, imag} */,
  {32'hbe150668, 32'h40655e30} /* (21, 28, 23) {real, imag} */,
  {32'h3e2832d7, 32'h400cc0fd} /* (21, 28, 22) {real, imag} */,
  {32'hc0205b87, 32'hbef9842c} /* (21, 28, 21) {real, imag} */,
  {32'hc02e7302, 32'hc00ed925} /* (21, 28, 20) {real, imag} */,
  {32'hc03d5931, 32'h3eed9433} /* (21, 28, 19) {real, imag} */,
  {32'hbe4d77dd, 32'hbfb8a10e} /* (21, 28, 18) {real, imag} */,
  {32'h3fefc660, 32'hbe61125a} /* (21, 28, 17) {real, imag} */,
  {32'hbe939bb3, 32'hbfeddea6} /* (21, 28, 16) {real, imag} */,
  {32'hbc413bbe, 32'h401a0724} /* (21, 28, 15) {real, imag} */,
  {32'h3e2b20ce, 32'h3fea8d65} /* (21, 28, 14) {real, imag} */,
  {32'h3fd95fd4, 32'h3f8571df} /* (21, 28, 13) {real, imag} */,
  {32'h3fd2d8da, 32'hbff70c57} /* (21, 28, 12) {real, imag} */,
  {32'hbd980a98, 32'hbf9a61d0} /* (21, 28, 11) {real, imag} */,
  {32'hc0540cab, 32'hbe498505} /* (21, 28, 10) {real, imag} */,
  {32'hbfd33170, 32'h3f77805f} /* (21, 28, 9) {real, imag} */,
  {32'h3ed8eb17, 32'hbf12b04d} /* (21, 28, 8) {real, imag} */,
  {32'hbf14df6d, 32'hc08f7186} /* (21, 28, 7) {real, imag} */,
  {32'h4004b748, 32'h3fbabcaa} /* (21, 28, 6) {real, imag} */,
  {32'hc08fdc85, 32'hc00d36ac} /* (21, 28, 5) {real, imag} */,
  {32'h3f02e598, 32'h3ff0b2f2} /* (21, 28, 4) {real, imag} */,
  {32'hbe82165c, 32'hbfe6a094} /* (21, 28, 3) {real, imag} */,
  {32'h3da6de0a, 32'h4040c515} /* (21, 28, 2) {real, imag} */,
  {32'h3ef2fb35, 32'hbf622a32} /* (21, 28, 1) {real, imag} */,
  {32'h3fbca97c, 32'h3f1c5702} /* (21, 28, 0) {real, imag} */,
  {32'hc0cfde39, 32'h400ec508} /* (21, 27, 31) {real, imag} */,
  {32'h400eab21, 32'h3f7e72b1} /* (21, 27, 30) {real, imag} */,
  {32'hbe020cc0, 32'h4011495a} /* (21, 27, 29) {real, imag} */,
  {32'hbf0db96f, 32'h4031cc62} /* (21, 27, 28) {real, imag} */,
  {32'h3f506413, 32'hc03d684a} /* (21, 27, 27) {real, imag} */,
  {32'hbf686a81, 32'h3f4e5870} /* (21, 27, 26) {real, imag} */,
  {32'hc0128b94, 32'h3ffbde9e} /* (21, 27, 25) {real, imag} */,
  {32'h4030f941, 32'hbf7ac793} /* (21, 27, 24) {real, imag} */,
  {32'h3fae60cf, 32'h403b7957} /* (21, 27, 23) {real, imag} */,
  {32'hbeb16946, 32'hbff1242b} /* (21, 27, 22) {real, imag} */,
  {32'h3ff3ff47, 32'hc037d502} /* (21, 27, 21) {real, imag} */,
  {32'hc0598c76, 32'h3e9864dc} /* (21, 27, 20) {real, imag} */,
  {32'hc017a706, 32'hbf9ebc3e} /* (21, 27, 19) {real, imag} */,
  {32'hbfd45e1d, 32'hbec041ca} /* (21, 27, 18) {real, imag} */,
  {32'h4016bccf, 32'h3f52a3fb} /* (21, 27, 17) {real, imag} */,
  {32'h3fea6f47, 32'h3dad585e} /* (21, 27, 16) {real, imag} */,
  {32'hbe3d883a, 32'hbea8509f} /* (21, 27, 15) {real, imag} */,
  {32'hbf839e61, 32'h3f4db962} /* (21, 27, 14) {real, imag} */,
  {32'hbf32ece2, 32'hc04b9f53} /* (21, 27, 13) {real, imag} */,
  {32'h3f82ce52, 32'hbf912def} /* (21, 27, 12) {real, imag} */,
  {32'h3fa2bee0, 32'h3ff3523a} /* (21, 27, 11) {real, imag} */,
  {32'hc022c9f7, 32'hbed8b16e} /* (21, 27, 10) {real, imag} */,
  {32'h3d97b5d8, 32'h3fe4c1ed} /* (21, 27, 9) {real, imag} */,
  {32'h3eeea292, 32'hbed7490a} /* (21, 27, 8) {real, imag} */,
  {32'hbfa37a0d, 32'hc00b2349} /* (21, 27, 7) {real, imag} */,
  {32'hbf1c9fde, 32'hbf0fed86} /* (21, 27, 6) {real, imag} */,
  {32'h3fec4949, 32'h3f960986} /* (21, 27, 5) {real, imag} */,
  {32'h3f845a37, 32'h4039cc84} /* (21, 27, 4) {real, imag} */,
  {32'h3e9c1be3, 32'hbd30678c} /* (21, 27, 3) {real, imag} */,
  {32'h3fd9d152, 32'hc01108c9} /* (21, 27, 2) {real, imag} */,
  {32'hc020077c, 32'hc05e5d75} /* (21, 27, 1) {real, imag} */,
  {32'hc0142e01, 32'hbf69279a} /* (21, 27, 0) {real, imag} */,
  {32'h4001f84b, 32'hbf52d613} /* (21, 26, 31) {real, imag} */,
  {32'hbe9c760a, 32'hbfdfb3d4} /* (21, 26, 30) {real, imag} */,
  {32'h3fd91974, 32'hbec68958} /* (21, 26, 29) {real, imag} */,
  {32'h401e9db7, 32'h3ff7aba0} /* (21, 26, 28) {real, imag} */,
  {32'h3fe23ff5, 32'h3f574563} /* (21, 26, 27) {real, imag} */,
  {32'hbff13e56, 32'hc01cdf96} /* (21, 26, 26) {real, imag} */,
  {32'hbff5512b, 32'h3f814a29} /* (21, 26, 25) {real, imag} */,
  {32'hc01f57df, 32'h3ea311cf} /* (21, 26, 24) {real, imag} */,
  {32'h4039d466, 32'hc0056b0b} /* (21, 26, 23) {real, imag} */,
  {32'hbe1c32cb, 32'hc09c1725} /* (21, 26, 22) {real, imag} */,
  {32'h3f3f4eef, 32'hc01f13f8} /* (21, 26, 21) {real, imag} */,
  {32'hbdbc56de, 32'hc0146082} /* (21, 26, 20) {real, imag} */,
  {32'hbf67447c, 32'hbefd710f} /* (21, 26, 19) {real, imag} */,
  {32'hbf353a97, 32'hbf75ba74} /* (21, 26, 18) {real, imag} */,
  {32'h3f0ce067, 32'h3f67a811} /* (21, 26, 17) {real, imag} */,
  {32'h3fc83131, 32'hbfde0c38} /* (21, 26, 16) {real, imag} */,
  {32'h3f970194, 32'h3ff52ec9} /* (21, 26, 15) {real, imag} */,
  {32'h3ffbf315, 32'hbfd2c8e3} /* (21, 26, 14) {real, imag} */,
  {32'hbfe7eee8, 32'h3ff8cdc7} /* (21, 26, 13) {real, imag} */,
  {32'h3ff2b7b4, 32'hc04b0aaf} /* (21, 26, 12) {real, imag} */,
  {32'hbf4e8969, 32'hbfb94286} /* (21, 26, 11) {real, imag} */,
  {32'h3e5e30d2, 32'h402b1332} /* (21, 26, 10) {real, imag} */,
  {32'h3f57e807, 32'h3ee172d2} /* (21, 26, 9) {real, imag} */,
  {32'hc065a4b5, 32'hc0205e9f} /* (21, 26, 8) {real, imag} */,
  {32'hbee5fda1, 32'h3f9a3f49} /* (21, 26, 7) {real, imag} */,
  {32'hbfff8755, 32'h3f8621a6} /* (21, 26, 6) {real, imag} */,
  {32'hc01ac7c0, 32'hbf84e087} /* (21, 26, 5) {real, imag} */,
  {32'h3fd8d137, 32'h3f53f608} /* (21, 26, 4) {real, imag} */,
  {32'hc02a9bbe, 32'h4010b18f} /* (21, 26, 3) {real, imag} */,
  {32'hbe795c78, 32'hbfb3d539} /* (21, 26, 2) {real, imag} */,
  {32'h40b78efd, 32'hbff6ba9a} /* (21, 26, 1) {real, imag} */,
  {32'hc070d5c4, 32'h3f2bb91e} /* (21, 26, 0) {real, imag} */,
  {32'h40896800, 32'h3f8c6d8f} /* (21, 25, 31) {real, imag} */,
  {32'hbcdd89a7, 32'hbe91ebe6} /* (21, 25, 30) {real, imag} */,
  {32'hbfa28867, 32'h406e4237} /* (21, 25, 29) {real, imag} */,
  {32'h3fe79009, 32'hbf77b9d6} /* (21, 25, 28) {real, imag} */,
  {32'hc00272df, 32'h408f6688} /* (21, 25, 27) {real, imag} */,
  {32'h4085617d, 32'h3deec9da} /* (21, 25, 26) {real, imag} */,
  {32'h3fb06c72, 32'hc03d3d64} /* (21, 25, 25) {real, imag} */,
  {32'h4031f627, 32'hbf434b65} /* (21, 25, 24) {real, imag} */,
  {32'h3f6f70cf, 32'h397e78f8} /* (21, 25, 23) {real, imag} */,
  {32'hbf23d677, 32'h3f910cac} /* (21, 25, 22) {real, imag} */,
  {32'h403a1907, 32'hc008e4a2} /* (21, 25, 21) {real, imag} */,
  {32'hbe76afc3, 32'h3d8d39c2} /* (21, 25, 20) {real, imag} */,
  {32'hc001a47d, 32'h402d0695} /* (21, 25, 19) {real, imag} */,
  {32'h3f464e0a, 32'h3fbac320} /* (21, 25, 18) {real, imag} */,
  {32'hbfb5b28b, 32'hc005233a} /* (21, 25, 17) {real, imag} */,
  {32'hc001d7be, 32'h3e465af5} /* (21, 25, 16) {real, imag} */,
  {32'h3f21e498, 32'hbf0188ee} /* (21, 25, 15) {real, imag} */,
  {32'hbec1c3a0, 32'h3f81cad2} /* (21, 25, 14) {real, imag} */,
  {32'hbf890f46, 32'hc06052bf} /* (21, 25, 13) {real, imag} */,
  {32'h4096dfa8, 32'hbfd4b642} /* (21, 25, 12) {real, imag} */,
  {32'hc02e825a, 32'h3e64a38e} /* (21, 25, 11) {real, imag} */,
  {32'h3e797008, 32'hc07db43f} /* (21, 25, 10) {real, imag} */,
  {32'hc038c07f, 32'h3f99dc3e} /* (21, 25, 9) {real, imag} */,
  {32'h400e1184, 32'h3ed003d6} /* (21, 25, 8) {real, imag} */,
  {32'hbedfac49, 32'h3f7124f4} /* (21, 25, 7) {real, imag} */,
  {32'hbfb2dd6a, 32'h3f990f96} /* (21, 25, 6) {real, imag} */,
  {32'hc04c0859, 32'hbf3ee9e8} /* (21, 25, 5) {real, imag} */,
  {32'h3d5bb6f3, 32'h3f9cb73c} /* (21, 25, 4) {real, imag} */,
  {32'h402bd3ad, 32'hc0745c28} /* (21, 25, 3) {real, imag} */,
  {32'hc00639c0, 32'h3e4b436b} /* (21, 25, 2) {real, imag} */,
  {32'h4074ca4d, 32'h3f7e1b77} /* (21, 25, 1) {real, imag} */,
  {32'hc0523611, 32'hbfaa0fd6} /* (21, 25, 0) {real, imag} */,
  {32'h3d948aa4, 32'h3f89e71d} /* (21, 24, 31) {real, imag} */,
  {32'hbfb92b4e, 32'hbc5ac838} /* (21, 24, 30) {real, imag} */,
  {32'h3f943f0d, 32'hbd27080e} /* (21, 24, 29) {real, imag} */,
  {32'hc00a5606, 32'hbfeb09ea} /* (21, 24, 28) {real, imag} */,
  {32'hbfa9bbd2, 32'hc012cb4c} /* (21, 24, 27) {real, imag} */,
  {32'hc061918a, 32'hbfdf0f92} /* (21, 24, 26) {real, imag} */,
  {32'h40434d19, 32'hbe353c20} /* (21, 24, 25) {real, imag} */,
  {32'h4051e72e, 32'h3e7dab3e} /* (21, 24, 24) {real, imag} */,
  {32'hbfc7fda6, 32'h3f2fde58} /* (21, 24, 23) {real, imag} */,
  {32'hbfff125c, 32'h3fbf64f1} /* (21, 24, 22) {real, imag} */,
  {32'hbed7b49b, 32'h3ffe4493} /* (21, 24, 21) {real, imag} */,
  {32'hbedd36b4, 32'hbfc21ab2} /* (21, 24, 20) {real, imag} */,
  {32'h3fc959ef, 32'hc0a0b63d} /* (21, 24, 19) {real, imag} */,
  {32'hbf931733, 32'hbf18fe43} /* (21, 24, 18) {real, imag} */,
  {32'hbfa7be59, 32'hbf2c8133} /* (21, 24, 17) {real, imag} */,
  {32'h3f6347a5, 32'h3d188e42} /* (21, 24, 16) {real, imag} */,
  {32'hbfa79d1e, 32'h3f9c2503} /* (21, 24, 15) {real, imag} */,
  {32'h400e1da0, 32'h3ff064b9} /* (21, 24, 14) {real, imag} */,
  {32'hbe024d93, 32'hbf06fcf7} /* (21, 24, 13) {real, imag} */,
  {32'hbe880eef, 32'h3fca28d2} /* (21, 24, 12) {real, imag} */,
  {32'h4092bf08, 32'hbe06f85e} /* (21, 24, 11) {real, imag} */,
  {32'h40856658, 32'hc006b1ad} /* (21, 24, 10) {real, imag} */,
  {32'hbef17046, 32'hc00a2e36} /* (21, 24, 9) {real, imag} */,
  {32'hbfd1c85e, 32'h3fee92b7} /* (21, 24, 8) {real, imag} */,
  {32'hc093e57d, 32'h3fc3597e} /* (21, 24, 7) {real, imag} */,
  {32'h3f0dd042, 32'h3f0156e2} /* (21, 24, 6) {real, imag} */,
  {32'h3e27e788, 32'h3ffd182f} /* (21, 24, 5) {real, imag} */,
  {32'h3ff040ca, 32'h40041b37} /* (21, 24, 4) {real, imag} */,
  {32'hbf8e72b2, 32'hbf5bcc39} /* (21, 24, 3) {real, imag} */,
  {32'hbfc34675, 32'hbf5f60e6} /* (21, 24, 2) {real, imag} */,
  {32'hbed1e88a, 32'h3fc50d44} /* (21, 24, 1) {real, imag} */,
  {32'h3f533ab1, 32'hbf762b7d} /* (21, 24, 0) {real, imag} */,
  {32'h409f3251, 32'hbec3ef9c} /* (21, 23, 31) {real, imag} */,
  {32'hbdb8f85c, 32'h40161168} /* (21, 23, 30) {real, imag} */,
  {32'h3e96484e, 32'h40280bd1} /* (21, 23, 29) {real, imag} */,
  {32'hbd8c66a2, 32'hbfb154fb} /* (21, 23, 28) {real, imag} */,
  {32'h3feb19a6, 32'h3f7067ee} /* (21, 23, 27) {real, imag} */,
  {32'h3f1d6da6, 32'hc00a6c5d} /* (21, 23, 26) {real, imag} */,
  {32'hbe4e6550, 32'hbf2c67eb} /* (21, 23, 25) {real, imag} */,
  {32'h401b2b48, 32'hbf02a021} /* (21, 23, 24) {real, imag} */,
  {32'hc0072b9d, 32'h3e8200ef} /* (21, 23, 23) {real, imag} */,
  {32'hbffa931a, 32'h3e06bb8f} /* (21, 23, 22) {real, imag} */,
  {32'hc01f1de0, 32'hbf281372} /* (21, 23, 21) {real, imag} */,
  {32'h3fbdd610, 32'hc0222ac7} /* (21, 23, 20) {real, imag} */,
  {32'h3f41b52b, 32'hc00800ab} /* (21, 23, 19) {real, imag} */,
  {32'hbfeba8f5, 32'hbf2b5c9e} /* (21, 23, 18) {real, imag} */,
  {32'hbfbf33a8, 32'h3eced4bb} /* (21, 23, 17) {real, imag} */,
  {32'h3f6745cb, 32'h3fd96933} /* (21, 23, 16) {real, imag} */,
  {32'hbf8a61b0, 32'h4087af4e} /* (21, 23, 15) {real, imag} */,
  {32'hbf558cc9, 32'hbe84ba23} /* (21, 23, 14) {real, imag} */,
  {32'h3f88574a, 32'hbf9752bf} /* (21, 23, 13) {real, imag} */,
  {32'hbf46dc88, 32'h3f8eef93} /* (21, 23, 12) {real, imag} */,
  {32'h3fa21831, 32'h3f9534e8} /* (21, 23, 11) {real, imag} */,
  {32'hc07690a9, 32'h4040391e} /* (21, 23, 10) {real, imag} */,
  {32'hc02025c9, 32'hbfe131c9} /* (21, 23, 9) {real, imag} */,
  {32'hc037efbf, 32'hc01b890d} /* (21, 23, 8) {real, imag} */,
  {32'h3ffe2e18, 32'hc02c0a1b} /* (21, 23, 7) {real, imag} */,
  {32'hbdc8c7ff, 32'h3f0979ce} /* (21, 23, 6) {real, imag} */,
  {32'hbfdfb7ad, 32'hc00102ff} /* (21, 23, 5) {real, imag} */,
  {32'hc04ef84a, 32'hbf009ef8} /* (21, 23, 4) {real, imag} */,
  {32'hc0028fab, 32'hbe601c48} /* (21, 23, 3) {real, imag} */,
  {32'h40096e6b, 32'hc002ca42} /* (21, 23, 2) {real, imag} */,
  {32'hc00a72e8, 32'h3eee4b1e} /* (21, 23, 1) {real, imag} */,
  {32'h40325ad0, 32'h40437eda} /* (21, 23, 0) {real, imag} */,
  {32'hc067df18, 32'hc014797a} /* (21, 22, 31) {real, imag} */,
  {32'hbfe6014d, 32'h3f3efff2} /* (21, 22, 30) {real, imag} */,
  {32'hbf56ce19, 32'hc0095724} /* (21, 22, 29) {real, imag} */,
  {32'hbf9b5e9c, 32'hbfac0757} /* (21, 22, 28) {real, imag} */,
  {32'hbf8e5fda, 32'h3fb40ea8} /* (21, 22, 27) {real, imag} */,
  {32'h3f59b8bb, 32'h3f585b72} /* (21, 22, 26) {real, imag} */,
  {32'h3f3a3e76, 32'h3dcaaa59} /* (21, 22, 25) {real, imag} */,
  {32'h3fbe059d, 32'h403622a6} /* (21, 22, 24) {real, imag} */,
  {32'hc02e5550, 32'h409b5cc6} /* (21, 22, 23) {real, imag} */,
  {32'h3fcf626b, 32'hc043db4d} /* (21, 22, 22) {real, imag} */,
  {32'h3f30d726, 32'h3ea651d6} /* (21, 22, 21) {real, imag} */,
  {32'h405506f2, 32'hbf2b473b} /* (21, 22, 20) {real, imag} */,
  {32'hc055514a, 32'h3fbc1784} /* (21, 22, 19) {real, imag} */,
  {32'h405d3c32, 32'hbfaceb75} /* (21, 22, 18) {real, imag} */,
  {32'hbe0d85c0, 32'hbef15fa1} /* (21, 22, 17) {real, imag} */,
  {32'hbe252814, 32'h3fa667e4} /* (21, 22, 16) {real, imag} */,
  {32'h3fb6049a, 32'h3e51f497} /* (21, 22, 15) {real, imag} */,
  {32'hc0096c94, 32'hc00cbd35} /* (21, 22, 14) {real, imag} */,
  {32'h3f3961a8, 32'h3f7618a4} /* (21, 22, 13) {real, imag} */,
  {32'hc0275ea1, 32'hbf84c2c8} /* (21, 22, 12) {real, imag} */,
  {32'h3f98169f, 32'hbf0b38c1} /* (21, 22, 11) {real, imag} */,
  {32'hbfd0e7f0, 32'h3d4c5904} /* (21, 22, 10) {real, imag} */,
  {32'hc096f2ba, 32'hc01f8404} /* (21, 22, 9) {real, imag} */,
  {32'h40be212d, 32'h409c66d9} /* (21, 22, 8) {real, imag} */,
  {32'hbe266f6a, 32'hc09e0088} /* (21, 22, 7) {real, imag} */,
  {32'hbf49ebbb, 32'h401c821d} /* (21, 22, 6) {real, imag} */,
  {32'h400c206d, 32'h3f795a1f} /* (21, 22, 5) {real, imag} */,
  {32'h3ef1d154, 32'hc0099466} /* (21, 22, 4) {real, imag} */,
  {32'h40121e3a, 32'h3fbc74fa} /* (21, 22, 3) {real, imag} */,
  {32'hbf5549a4, 32'h3f154948} /* (21, 22, 2) {real, imag} */,
  {32'hbee5d1c0, 32'hbe129e3a} /* (21, 22, 1) {real, imag} */,
  {32'hbf56ea16, 32'hc08a1edd} /* (21, 22, 0) {real, imag} */,
  {32'hbda77b81, 32'h3f535290} /* (21, 21, 31) {real, imag} */,
  {32'hbf80046f, 32'hbde5c42a} /* (21, 21, 30) {real, imag} */,
  {32'hc0447e9c, 32'hbf023503} /* (21, 21, 29) {real, imag} */,
  {32'hc06dd8a1, 32'hc074044f} /* (21, 21, 28) {real, imag} */,
  {32'hbecd51ff, 32'h3ef3a6d9} /* (21, 21, 27) {real, imag} */,
  {32'hbf2538d6, 32'h3fef03a3} /* (21, 21, 26) {real, imag} */,
  {32'hbdc6f15d, 32'h3eb5bfc6} /* (21, 21, 25) {real, imag} */,
  {32'h3eeea5fd, 32'hbf7f4d99} /* (21, 21, 24) {real, imag} */,
  {32'hbfdb6f59, 32'h3f87204e} /* (21, 21, 23) {real, imag} */,
  {32'h3f14663d, 32'h3fcc6b3e} /* (21, 21, 22) {real, imag} */,
  {32'hbdef3216, 32'hc06e0b4b} /* (21, 21, 21) {real, imag} */,
  {32'h4000173e, 32'hbf65af6c} /* (21, 21, 20) {real, imag} */,
  {32'hbf70072f, 32'h3f48b902} /* (21, 21, 19) {real, imag} */,
  {32'hbf71d263, 32'h4018e844} /* (21, 21, 18) {real, imag} */,
  {32'h3eb9e2f6, 32'hbf9050b9} /* (21, 21, 17) {real, imag} */,
  {32'hbf4fa3c0, 32'h3f7ae806} /* (21, 21, 16) {real, imag} */,
  {32'hbf099bde, 32'hc02c1c24} /* (21, 21, 15) {real, imag} */,
  {32'hc0661975, 32'h402a01ef} /* (21, 21, 14) {real, imag} */,
  {32'hbfbf0b3c, 32'h3f9356cf} /* (21, 21, 13) {real, imag} */,
  {32'hbfaf74c9, 32'h408ca1de} /* (21, 21, 12) {real, imag} */,
  {32'h3f5ded65, 32'h3fb4694f} /* (21, 21, 11) {real, imag} */,
  {32'h40054836, 32'h3fa7b376} /* (21, 21, 10) {real, imag} */,
  {32'hbf31fd9a, 32'h3e3bd98a} /* (21, 21, 9) {real, imag} */,
  {32'h40078cb1, 32'h3ff3131c} /* (21, 21, 8) {real, imag} */,
  {32'hc017e1f5, 32'h3fa09256} /* (21, 21, 7) {real, imag} */,
  {32'h3fb78b0b, 32'h401cc3d4} /* (21, 21, 6) {real, imag} */,
  {32'hbf3a6105, 32'h3fd70572} /* (21, 21, 5) {real, imag} */,
  {32'hbee45db7, 32'h3ef5b72e} /* (21, 21, 4) {real, imag} */,
  {32'hc00babd5, 32'hbf34306d} /* (21, 21, 3) {real, imag} */,
  {32'hbfef6388, 32'hc07fc043} /* (21, 21, 2) {real, imag} */,
  {32'hc08906a2, 32'hbf7e6603} /* (21, 21, 1) {real, imag} */,
  {32'hbf924a23, 32'h4015a117} /* (21, 21, 0) {real, imag} */,
  {32'hc012b468, 32'h4000ce3b} /* (21, 20, 31) {real, imag} */,
  {32'hc0093ae7, 32'hc01bef47} /* (21, 20, 30) {real, imag} */,
  {32'hbfa66bdd, 32'hbf23df64} /* (21, 20, 29) {real, imag} */,
  {32'h3f05724a, 32'hbe67668f} /* (21, 20, 28) {real, imag} */,
  {32'hbf8850bc, 32'h40067273} /* (21, 20, 27) {real, imag} */,
  {32'h3f253058, 32'h3e6b0dc7} /* (21, 20, 26) {real, imag} */,
  {32'h40335867, 32'h3eea0727} /* (21, 20, 25) {real, imag} */,
  {32'hbfdb9d08, 32'h3fc244b1} /* (21, 20, 24) {real, imag} */,
  {32'h3f07ad0d, 32'hbf29e3ad} /* (21, 20, 23) {real, imag} */,
  {32'h3f5c98c9, 32'hbd828133} /* (21, 20, 22) {real, imag} */,
  {32'hbf870c26, 32'h3f59269d} /* (21, 20, 21) {real, imag} */,
  {32'hbd17b16f, 32'h3f66aa35} /* (21, 20, 20) {real, imag} */,
  {32'h3f8887d2, 32'h406a0afc} /* (21, 20, 19) {real, imag} */,
  {32'h3e19084f, 32'hbfb9b5d4} /* (21, 20, 18) {real, imag} */,
  {32'hbf6242e5, 32'h401b14d2} /* (21, 20, 17) {real, imag} */,
  {32'hbef4b74e, 32'h3ddbb3dd} /* (21, 20, 16) {real, imag} */,
  {32'hbfa0335c, 32'h402d6f02} /* (21, 20, 15) {real, imag} */,
  {32'h4037db7a, 32'h407d2c5e} /* (21, 20, 14) {real, imag} */,
  {32'hc0132842, 32'hc03393c0} /* (21, 20, 13) {real, imag} */,
  {32'hbeedfdab, 32'h406fe19f} /* (21, 20, 12) {real, imag} */,
  {32'h3ec6f48f, 32'h405374ad} /* (21, 20, 11) {real, imag} */,
  {32'hc00792a8, 32'h403299ed} /* (21, 20, 10) {real, imag} */,
  {32'hbf80fbdb, 32'h3f812fe6} /* (21, 20, 9) {real, imag} */,
  {32'h3ef58bbd, 32'hc042b3f5} /* (21, 20, 8) {real, imag} */,
  {32'hbfece681, 32'hbfd5c6be} /* (21, 20, 7) {real, imag} */,
  {32'hc0008776, 32'hc050f2bb} /* (21, 20, 6) {real, imag} */,
  {32'h3fafa3d5, 32'h3fb5aa56} /* (21, 20, 5) {real, imag} */,
  {32'h3fdc02a4, 32'hbebf34b8} /* (21, 20, 4) {real, imag} */,
  {32'hbd0d7db0, 32'hbe25b892} /* (21, 20, 3) {real, imag} */,
  {32'hc0316679, 32'h3e65f308} /* (21, 20, 2) {real, imag} */,
  {32'h3fc64aa1, 32'hc0085727} /* (21, 20, 1) {real, imag} */,
  {32'h3e6f1eb1, 32'h3fca36ed} /* (21, 20, 0) {real, imag} */,
  {32'hbf825772, 32'hbeb837a7} /* (21, 19, 31) {real, imag} */,
  {32'hbf55d0ef, 32'hbfbd31e3} /* (21, 19, 30) {real, imag} */,
  {32'hc0004306, 32'h3e31e30f} /* (21, 19, 29) {real, imag} */,
  {32'h3f8928ba, 32'hbf840c4e} /* (21, 19, 28) {real, imag} */,
  {32'h3ebf280a, 32'h40181ddc} /* (21, 19, 27) {real, imag} */,
  {32'h3ff5350c, 32'hbd17fdc0} /* (21, 19, 26) {real, imag} */,
  {32'hbe43d348, 32'hbf19ddae} /* (21, 19, 25) {real, imag} */,
  {32'h3fba3564, 32'h3f4655e0} /* (21, 19, 24) {real, imag} */,
  {32'hbf49af94, 32'h3fe1b5e7} /* (21, 19, 23) {real, imag} */,
  {32'h3f09376d, 32'hbf540168} /* (21, 19, 22) {real, imag} */,
  {32'h3fa4fde9, 32'h4020a02a} /* (21, 19, 21) {real, imag} */,
  {32'h3fbb5c65, 32'h3fb0b2ed} /* (21, 19, 20) {real, imag} */,
  {32'hbebe8561, 32'h3fc42530} /* (21, 19, 19) {real, imag} */,
  {32'h3f2cc80f, 32'h3f312d81} /* (21, 19, 18) {real, imag} */,
  {32'hbf55dc86, 32'h3f968568} /* (21, 19, 17) {real, imag} */,
  {32'hbf49c893, 32'h3f30cc1f} /* (21, 19, 16) {real, imag} */,
  {32'hbfe52b87, 32'hbef296b2} /* (21, 19, 15) {real, imag} */,
  {32'h3d156ef7, 32'hc057c6fd} /* (21, 19, 14) {real, imag} */,
  {32'hbf13554d, 32'h3fc077d3} /* (21, 19, 13) {real, imag} */,
  {32'h3f794910, 32'hc00ac292} /* (21, 19, 12) {real, imag} */,
  {32'hbe05366e, 32'h3ed3608b} /* (21, 19, 11) {real, imag} */,
  {32'h40008981, 32'h40484377} /* (21, 19, 10) {real, imag} */,
  {32'h402e75ab, 32'hc0024a31} /* (21, 19, 9) {real, imag} */,
  {32'h3f282fb8, 32'hbe3f43c3} /* (21, 19, 8) {real, imag} */,
  {32'h4025bcc5, 32'h3f84ac4d} /* (21, 19, 7) {real, imag} */,
  {32'h3fa020e1, 32'hbf012953} /* (21, 19, 6) {real, imag} */,
  {32'hbf95621c, 32'hbfc7b2b2} /* (21, 19, 5) {real, imag} */,
  {32'hbf0d2e7d, 32'h3d3d19a4} /* (21, 19, 4) {real, imag} */,
  {32'h3f28789d, 32'hbfd74b47} /* (21, 19, 3) {real, imag} */,
  {32'h3f3adde9, 32'hc00e84c0} /* (21, 19, 2) {real, imag} */,
  {32'h3f5700f0, 32'h3fc52460} /* (21, 19, 1) {real, imag} */,
  {32'h3fee56d4, 32'hbf8fe7b6} /* (21, 19, 0) {real, imag} */,
  {32'hbfdbaaf2, 32'hc01a1f97} /* (21, 18, 31) {real, imag} */,
  {32'h3f8ad87e, 32'hbed13814} /* (21, 18, 30) {real, imag} */,
  {32'h3e0f7cf0, 32'h3fcbac0f} /* (21, 18, 29) {real, imag} */,
  {32'h3dec5466, 32'h3ea1f45a} /* (21, 18, 28) {real, imag} */,
  {32'h3e3d7d6d, 32'hc00f49e9} /* (21, 18, 27) {real, imag} */,
  {32'hbd072152, 32'h3f597190} /* (21, 18, 26) {real, imag} */,
  {32'hbfcc91b5, 32'h3e792c11} /* (21, 18, 25) {real, imag} */,
  {32'h3e147c1c, 32'h3f56d275} /* (21, 18, 24) {real, imag} */,
  {32'hbf6afd8e, 32'h3eec0126} /* (21, 18, 23) {real, imag} */,
  {32'hbfb489fa, 32'hbea8867e} /* (21, 18, 22) {real, imag} */,
  {32'hbe4b932c, 32'hc007b41e} /* (21, 18, 21) {real, imag} */,
  {32'h3e3f1539, 32'h3f8cc537} /* (21, 18, 20) {real, imag} */,
  {32'h40107f40, 32'hbf8c8bda} /* (21, 18, 19) {real, imag} */,
  {32'h3f482d1b, 32'h3f555a70} /* (21, 18, 18) {real, imag} */,
  {32'hbf7c3d50, 32'hbf98f5be} /* (21, 18, 17) {real, imag} */,
  {32'h40062259, 32'h4035ab7e} /* (21, 18, 16) {real, imag} */,
  {32'h3efdc52b, 32'hbf559def} /* (21, 18, 15) {real, imag} */,
  {32'h405095d3, 32'hbfdac6ef} /* (21, 18, 14) {real, imag} */,
  {32'h3f9dec76, 32'h3fdd4322} /* (21, 18, 13) {real, imag} */,
  {32'hbe7cb05f, 32'h3dc2f9a1} /* (21, 18, 12) {real, imag} */,
  {32'hbe290387, 32'hbe4d06b4} /* (21, 18, 11) {real, imag} */,
  {32'hc0914c44, 32'hbde65791} /* (21, 18, 10) {real, imag} */,
  {32'h3ff96ca6, 32'hbf9a19f7} /* (21, 18, 9) {real, imag} */,
  {32'hbfd53c65, 32'h4021b1db} /* (21, 18, 8) {real, imag} */,
  {32'hbd6dfbd0, 32'hbde8ab52} /* (21, 18, 7) {real, imag} */,
  {32'hbf5a5cdb, 32'hbe20b4c7} /* (21, 18, 6) {real, imag} */,
  {32'h3eed0bdc, 32'h3d197b12} /* (21, 18, 5) {real, imag} */,
  {32'hbf5a6aa6, 32'hbf74bd3e} /* (21, 18, 4) {real, imag} */,
  {32'h3f6b8ffb, 32'h3fe6232f} /* (21, 18, 3) {real, imag} */,
  {32'hbfa4a4b6, 32'hbfadd63e} /* (21, 18, 2) {real, imag} */,
  {32'hbe5b2e85, 32'h3fee0be7} /* (21, 18, 1) {real, imag} */,
  {32'hbeec714b, 32'h3fe007ad} /* (21, 18, 0) {real, imag} */,
  {32'h3f6a26c8, 32'hbf36886b} /* (21, 17, 31) {real, imag} */,
  {32'h3e2cf09b, 32'h3ccbbb12} /* (21, 17, 30) {real, imag} */,
  {32'hbd08861f, 32'hbfe8ee6d} /* (21, 17, 29) {real, imag} */,
  {32'h3e85f17e, 32'h3fd8735d} /* (21, 17, 28) {real, imag} */,
  {32'h3fc14131, 32'hbf9df864} /* (21, 17, 27) {real, imag} */,
  {32'hbf5293d7, 32'hbfa47fbb} /* (21, 17, 26) {real, imag} */,
  {32'h3f83afa5, 32'h3f5a5759} /* (21, 17, 25) {real, imag} */,
  {32'hbe0ba70c, 32'hbfec050c} /* (21, 17, 24) {real, imag} */,
  {32'hbf879099, 32'hbe0476ed} /* (21, 17, 23) {real, imag} */,
  {32'h3f81478b, 32'h3f869a87} /* (21, 17, 22) {real, imag} */,
  {32'h4038899b, 32'h4037a75d} /* (21, 17, 21) {real, imag} */,
  {32'h3f2ba702, 32'h3ec76247} /* (21, 17, 20) {real, imag} */,
  {32'hc02934b5, 32'h3f19289d} /* (21, 17, 19) {real, imag} */,
  {32'h3ecb01ac, 32'hbf739c94} /* (21, 17, 18) {real, imag} */,
  {32'hbf6a1370, 32'h3ecba7e8} /* (21, 17, 17) {real, imag} */,
  {32'hbfb9c564, 32'hbf085960} /* (21, 17, 16) {real, imag} */,
  {32'h3dd7a7e7, 32'h3ef75ce6} /* (21, 17, 15) {real, imag} */,
  {32'h3f074e39, 32'h3ff48117} /* (21, 17, 14) {real, imag} */,
  {32'h3f1aa5de, 32'h401aafb7} /* (21, 17, 13) {real, imag} */,
  {32'hbfbe72de, 32'h3f769fba} /* (21, 17, 12) {real, imag} */,
  {32'h3fd8e01e, 32'hc0080fbd} /* (21, 17, 11) {real, imag} */,
  {32'h3e85ffad, 32'hbf26d2b7} /* (21, 17, 10) {real, imag} */,
  {32'hbfb44c35, 32'h3efa7885} /* (21, 17, 9) {real, imag} */,
  {32'hc0423654, 32'hc01146c2} /* (21, 17, 8) {real, imag} */,
  {32'h3ed6efd4, 32'h3f339d59} /* (21, 17, 7) {real, imag} */,
  {32'h3e0b101b, 32'h3f0e77a5} /* (21, 17, 6) {real, imag} */,
  {32'hbe97dd9b, 32'hc005605f} /* (21, 17, 5) {real, imag} */,
  {32'hbebd155b, 32'h3df2455a} /* (21, 17, 4) {real, imag} */,
  {32'hbfa793e7, 32'hbf9b3b06} /* (21, 17, 3) {real, imag} */,
  {32'hbfac40cf, 32'hbe695ff6} /* (21, 17, 2) {real, imag} */,
  {32'h3fdf9015, 32'h3f6e6a00} /* (21, 17, 1) {real, imag} */,
  {32'h3f4180e1, 32'h3e0b031a} /* (21, 17, 0) {real, imag} */,
  {32'hbf2cbdb0, 32'h3f1ff262} /* (21, 16, 31) {real, imag} */,
  {32'h3eee991c, 32'hbf5973d2} /* (21, 16, 30) {real, imag} */,
  {32'h3f9d3176, 32'h3dc30b37} /* (21, 16, 29) {real, imag} */,
  {32'h3f6241c5, 32'h3dd33b76} /* (21, 16, 28) {real, imag} */,
  {32'hbfc45bd9, 32'hbf1e2642} /* (21, 16, 27) {real, imag} */,
  {32'h3e25e021, 32'hbfc8d1d6} /* (21, 16, 26) {real, imag} */,
  {32'h3fa0a7f5, 32'h40111045} /* (21, 16, 25) {real, imag} */,
  {32'h3f8ae2be, 32'h3ff10e60} /* (21, 16, 24) {real, imag} */,
  {32'hbd427509, 32'h403c4802} /* (21, 16, 23) {real, imag} */,
  {32'hbf3eb191, 32'h3f7f54e8} /* (21, 16, 22) {real, imag} */,
  {32'h3f507182, 32'h3fcc6e45} /* (21, 16, 21) {real, imag} */,
  {32'h3f26b087, 32'hbfa4ea3c} /* (21, 16, 20) {real, imag} */,
  {32'h4038fab3, 32'h3f86f750} /* (21, 16, 19) {real, imag} */,
  {32'h3cebd6e3, 32'h3ec80168} /* (21, 16, 18) {real, imag} */,
  {32'hbf70c087, 32'h3f9f13fc} /* (21, 16, 17) {real, imag} */,
  {32'h3ed1fee4, 32'hbda47fe8} /* (21, 16, 16) {real, imag} */,
  {32'h3f9c52cd, 32'h3e1dc05d} /* (21, 16, 15) {real, imag} */,
  {32'h3f038e8d, 32'hbef68f3b} /* (21, 16, 14) {real, imag} */,
  {32'hbf8af5e9, 32'hbf993f2d} /* (21, 16, 13) {real, imag} */,
  {32'hbf9d8f2b, 32'h3f901518} /* (21, 16, 12) {real, imag} */,
  {32'hbf8b0ec5, 32'hbfed9f24} /* (21, 16, 11) {real, imag} */,
  {32'hbed09cf9, 32'hbede6055} /* (21, 16, 10) {real, imag} */,
  {32'h408a8007, 32'hbef721a4} /* (21, 16, 9) {real, imag} */,
  {32'h3f965d9a, 32'h3f12eec1} /* (21, 16, 8) {real, imag} */,
  {32'hbeed29e2, 32'hbe7604cf} /* (21, 16, 7) {real, imag} */,
  {32'hbf9215d0, 32'h3f47f623} /* (21, 16, 6) {real, imag} */,
  {32'h3d330c01, 32'hc0062225} /* (21, 16, 5) {real, imag} */,
  {32'hbf590ea9, 32'hbde99a01} /* (21, 16, 4) {real, imag} */,
  {32'hbf4e9d25, 32'h3ef05a6e} /* (21, 16, 3) {real, imag} */,
  {32'hbd22a7b8, 32'hbdba06b4} /* (21, 16, 2) {real, imag} */,
  {32'hbda28af3, 32'hbf44160d} /* (21, 16, 1) {real, imag} */,
  {32'h3ff417fc, 32'hbecbf637} /* (21, 16, 0) {real, imag} */,
  {32'hbf80985e, 32'hbdb739f2} /* (21, 15, 31) {real, imag} */,
  {32'h408a33fb, 32'hbe764095} /* (21, 15, 30) {real, imag} */,
  {32'h3f51abe4, 32'h3fa3463a} /* (21, 15, 29) {real, imag} */,
  {32'h3e6c8c2e, 32'h3f8bdb90} /* (21, 15, 28) {real, imag} */,
  {32'h3f93d410, 32'h3f8a6b85} /* (21, 15, 27) {real, imag} */,
  {32'hbfefbc2c, 32'hbfd9e60d} /* (21, 15, 26) {real, imag} */,
  {32'hc025e906, 32'h3ecb032e} /* (21, 15, 25) {real, imag} */,
  {32'hbd8de0ac, 32'hbe86b1b5} /* (21, 15, 24) {real, imag} */,
  {32'hbff6992e, 32'h3fc0f88d} /* (21, 15, 23) {real, imag} */,
  {32'h3f04260e, 32'h3f67fd93} /* (21, 15, 22) {real, imag} */,
  {32'hc00ecb50, 32'hc021d7fa} /* (21, 15, 21) {real, imag} */,
  {32'h3e5550c3, 32'hbfb2df6c} /* (21, 15, 20) {real, imag} */,
  {32'hc028aada, 32'h3f8f113c} /* (21, 15, 19) {real, imag} */,
  {32'h3e406efe, 32'hbfa6f738} /* (21, 15, 18) {real, imag} */,
  {32'hbff262fd, 32'hbf46d9ed} /* (21, 15, 17) {real, imag} */,
  {32'hbfb5c8c1, 32'hbfc88451} /* (21, 15, 16) {real, imag} */,
  {32'hbff3e997, 32'h3dce3df3} /* (21, 15, 15) {real, imag} */,
  {32'h3fb65747, 32'hbdbf90bb} /* (21, 15, 14) {real, imag} */,
  {32'h3d613245, 32'h3e5bd4d9} /* (21, 15, 13) {real, imag} */,
  {32'hbef82465, 32'h3f7ac534} /* (21, 15, 12) {real, imag} */,
  {32'hc02b0e64, 32'h406de636} /* (21, 15, 11) {real, imag} */,
  {32'h3f2b951f, 32'h3c3f7b20} /* (21, 15, 10) {real, imag} */,
  {32'hbf951a84, 32'h3ff40730} /* (21, 15, 9) {real, imag} */,
  {32'hbff54931, 32'hbeacce54} /* (21, 15, 8) {real, imag} */,
  {32'h3f5b8e18, 32'hbfa9cf24} /* (21, 15, 7) {real, imag} */,
  {32'h3eaa4c75, 32'h3f86789c} /* (21, 15, 6) {real, imag} */,
  {32'hbf9a243a, 32'h3f4e6674} /* (21, 15, 5) {real, imag} */,
  {32'hbe1cd454, 32'h3fa206b1} /* (21, 15, 4) {real, imag} */,
  {32'hbe50bf7b, 32'hc02e992f} /* (21, 15, 3) {real, imag} */,
  {32'h3f8fb071, 32'hbf3f3881} /* (21, 15, 2) {real, imag} */,
  {32'h3f8751f7, 32'h3ef0c56d} /* (21, 15, 1) {real, imag} */,
  {32'hbf2fd553, 32'h3f8ae94e} /* (21, 15, 0) {real, imag} */,
  {32'h3f2e5186, 32'h3e61ce19} /* (21, 14, 31) {real, imag} */,
  {32'hbe891f0e, 32'hbf5f3577} /* (21, 14, 30) {real, imag} */,
  {32'h3ea9cad5, 32'h3ff005c0} /* (21, 14, 29) {real, imag} */,
  {32'h3de2f9b4, 32'hbee6cb95} /* (21, 14, 28) {real, imag} */,
  {32'hbfd6bef4, 32'hbe07d195} /* (21, 14, 27) {real, imag} */,
  {32'hbf585c2d, 32'hbd4145e2} /* (21, 14, 26) {real, imag} */,
  {32'hbf754a9a, 32'h3fb36279} /* (21, 14, 25) {real, imag} */,
  {32'h3f5894b3, 32'h3f875ac3} /* (21, 14, 24) {real, imag} */,
  {32'h4032844e, 32'h3fd4d877} /* (21, 14, 23) {real, imag} */,
  {32'h3ecf63b7, 32'hbfeea4ea} /* (21, 14, 22) {real, imag} */,
  {32'hbedcea16, 32'hc06094eb} /* (21, 14, 21) {real, imag} */,
  {32'h3fe988f5, 32'h40223ddb} /* (21, 14, 20) {real, imag} */,
  {32'hbfbd5ccf, 32'h3f65a586} /* (21, 14, 19) {real, imag} */,
  {32'h406895cf, 32'hbee41431} /* (21, 14, 18) {real, imag} */,
  {32'h4005d873, 32'hc00bca01} /* (21, 14, 17) {real, imag} */,
  {32'h401ab647, 32'h3f45ca7d} /* (21, 14, 16) {real, imag} */,
  {32'hbe35e345, 32'hbe99e265} /* (21, 14, 15) {real, imag} */,
  {32'h3f69a875, 32'hc0232c3a} /* (21, 14, 14) {real, imag} */,
  {32'h3f93eedf, 32'hc03797e0} /* (21, 14, 13) {real, imag} */,
  {32'hbfd3ac4e, 32'h3f35ac5c} /* (21, 14, 12) {real, imag} */,
  {32'hbf9fa6c1, 32'h3e84fd47} /* (21, 14, 11) {real, imag} */,
  {32'h3f604be6, 32'hc0580caa} /* (21, 14, 10) {real, imag} */,
  {32'h3df4b129, 32'hc06a31e8} /* (21, 14, 9) {real, imag} */,
  {32'hbffe0675, 32'hbf896687} /* (21, 14, 8) {real, imag} */,
  {32'h400c07ce, 32'h3e879bd9} /* (21, 14, 7) {real, imag} */,
  {32'h3dd4d6d9, 32'h3f6d03e4} /* (21, 14, 6) {real, imag} */,
  {32'hbf8c399f, 32'hbfe8b884} /* (21, 14, 5) {real, imag} */,
  {32'h3e6af56a, 32'h3f3b216c} /* (21, 14, 4) {real, imag} */,
  {32'hbeefb87e, 32'h3f0b0a65} /* (21, 14, 3) {real, imag} */,
  {32'h3ff5ba49, 32'hc02f7018} /* (21, 14, 2) {real, imag} */,
  {32'h3fa14081, 32'hbfee188e} /* (21, 14, 1) {real, imag} */,
  {32'h3f9ba926, 32'h3e9ecfd7} /* (21, 14, 0) {real, imag} */,
  {32'hbf5ed44d, 32'h3f056ac8} /* (21, 13, 31) {real, imag} */,
  {32'hbcea39a2, 32'h3f509738} /* (21, 13, 30) {real, imag} */,
  {32'hbedea681, 32'h3fe721d6} /* (21, 13, 29) {real, imag} */,
  {32'h3f722936, 32'hbf755e9c} /* (21, 13, 28) {real, imag} */,
  {32'h3e8f61ea, 32'hbfba80fc} /* (21, 13, 27) {real, imag} */,
  {32'h3fa95e3d, 32'hbfcf1a00} /* (21, 13, 26) {real, imag} */,
  {32'hbf72a1c6, 32'hc022ad7e} /* (21, 13, 25) {real, imag} */,
  {32'hbf04f19e, 32'h3fbe28b5} /* (21, 13, 24) {real, imag} */,
  {32'h404fc16d, 32'h40039138} /* (21, 13, 23) {real, imag} */,
  {32'hbf659b07, 32'h3f9b9983} /* (21, 13, 22) {real, imag} */,
  {32'hbf7cdf05, 32'hbe90d767} /* (21, 13, 21) {real, imag} */,
  {32'hbcb670a4, 32'hbf0bbcd9} /* (21, 13, 20) {real, imag} */,
  {32'h3ef7abe2, 32'h3fc24426} /* (21, 13, 19) {real, imag} */,
  {32'hc0053662, 32'h3ee2d883} /* (21, 13, 18) {real, imag} */,
  {32'h4005a8e9, 32'h3fa91469} /* (21, 13, 17) {real, imag} */,
  {32'h3ea521dc, 32'h3fde8fa9} /* (21, 13, 16) {real, imag} */,
  {32'hbf201932, 32'h402adee0} /* (21, 13, 15) {real, imag} */,
  {32'h3fc27f5a, 32'hbf0e149f} /* (21, 13, 14) {real, imag} */,
  {32'h3ea940ae, 32'h3eb9fe44} /* (21, 13, 13) {real, imag} */,
  {32'hbd61f916, 32'hc03774d1} /* (21, 13, 12) {real, imag} */,
  {32'hc0786e46, 32'h3fad36bc} /* (21, 13, 11) {real, imag} */,
  {32'h3f541ca5, 32'hc03b55ff} /* (21, 13, 10) {real, imag} */,
  {32'hc0909243, 32'hbfd73ba9} /* (21, 13, 9) {real, imag} */,
  {32'h3fb7f9a9, 32'h3f21dfc9} /* (21, 13, 8) {real, imag} */,
  {32'hb9ebebf3, 32'h3fadb042} /* (21, 13, 7) {real, imag} */,
  {32'hbf5fd561, 32'hc055f229} /* (21, 13, 6) {real, imag} */,
  {32'h3f69923f, 32'h3fe8f297} /* (21, 13, 5) {real, imag} */,
  {32'h404fc5fb, 32'h3fe31ff4} /* (21, 13, 4) {real, imag} */,
  {32'h4008cd23, 32'hc02bc49e} /* (21, 13, 3) {real, imag} */,
  {32'h3fe925e8, 32'hbe647b7f} /* (21, 13, 2) {real, imag} */,
  {32'h40361a10, 32'h3fdc8ab8} /* (21, 13, 1) {real, imag} */,
  {32'hbd9e6f6f, 32'h3f6db5ef} /* (21, 13, 0) {real, imag} */,
  {32'hbef7271a, 32'h3f9c0bf0} /* (21, 12, 31) {real, imag} */,
  {32'hbfa329b7, 32'hbf9e6d31} /* (21, 12, 30) {real, imag} */,
  {32'h401c666a, 32'h3e18105e} /* (21, 12, 29) {real, imag} */,
  {32'hbdccf729, 32'hbf4d46a2} /* (21, 12, 28) {real, imag} */,
  {32'hbf9d017e, 32'hc04b14ce} /* (21, 12, 27) {real, imag} */,
  {32'h3f1705d8, 32'hbf8dd5c5} /* (21, 12, 26) {real, imag} */,
  {32'h3fb4e413, 32'h3ff927c1} /* (21, 12, 25) {real, imag} */,
  {32'hc00e0bb7, 32'hbfbe3eca} /* (21, 12, 24) {real, imag} */,
  {32'hbd0d1265, 32'hbf4ac2de} /* (21, 12, 23) {real, imag} */,
  {32'hbf6b6393, 32'hc0a5c8a5} /* (21, 12, 22) {real, imag} */,
  {32'hbfaf077a, 32'h3f050232} /* (21, 12, 21) {real, imag} */,
  {32'h40175c1e, 32'h4003963d} /* (21, 12, 20) {real, imag} */,
  {32'h3fc08735, 32'h403bd07a} /* (21, 12, 19) {real, imag} */,
  {32'h402dbf7a, 32'h40232a07} /* (21, 12, 18) {real, imag} */,
  {32'hbfd33ba7, 32'h400d1e7c} /* (21, 12, 17) {real, imag} */,
  {32'hbfbb8585, 32'h3f6aa5f0} /* (21, 12, 16) {real, imag} */,
  {32'h3f922667, 32'hbfc6d972} /* (21, 12, 15) {real, imag} */,
  {32'hbff2f56e, 32'hbe39efd0} /* (21, 12, 14) {real, imag} */,
  {32'h401a9545, 32'hbfba1465} /* (21, 12, 13) {real, imag} */,
  {32'hbf9b9a82, 32'h403e0a63} /* (21, 12, 12) {real, imag} */,
  {32'h3fb7b7ec, 32'hbe7aced1} /* (21, 12, 11) {real, imag} */,
  {32'hc0920035, 32'hc01ddb73} /* (21, 12, 10) {real, imag} */,
  {32'hc0796a4d, 32'h3f8ee1e7} /* (21, 12, 9) {real, imag} */,
  {32'h3f06a0b3, 32'hbff006fe} /* (21, 12, 8) {real, imag} */,
  {32'h3eebeb70, 32'hbee2327e} /* (21, 12, 7) {real, imag} */,
  {32'hc04b56ff, 32'h3fb37cd2} /* (21, 12, 6) {real, imag} */,
  {32'h401749b4, 32'h3f4d1069} /* (21, 12, 5) {real, imag} */,
  {32'hbfa3adac, 32'h3f3c18d8} /* (21, 12, 4) {real, imag} */,
  {32'hbddc7645, 32'hbfa1ee35} /* (21, 12, 3) {real, imag} */,
  {32'h3faf6842, 32'hbea717d5} /* (21, 12, 2) {real, imag} */,
  {32'h3de8f94c, 32'hbed8affa} /* (21, 12, 1) {real, imag} */,
  {32'hc007e07f, 32'h3fbdb675} /* (21, 12, 0) {real, imag} */,
  {32'h3fdd0e7f, 32'hc0211964} /* (21, 11, 31) {real, imag} */,
  {32'h3fdb5ea8, 32'h3f4cac77} /* (21, 11, 30) {real, imag} */,
  {32'hc032076d, 32'h3facecee} /* (21, 11, 29) {real, imag} */,
  {32'h3fa51fad, 32'hbfe7fa96} /* (21, 11, 28) {real, imag} */,
  {32'h3f0fca19, 32'hbfd74209} /* (21, 11, 27) {real, imag} */,
  {32'hbfe48e3d, 32'h3fcee5ef} /* (21, 11, 26) {real, imag} */,
  {32'h4009cd1d, 32'h3d659cad} /* (21, 11, 25) {real, imag} */,
  {32'hbf599f70, 32'h3d9279fc} /* (21, 11, 24) {real, imag} */,
  {32'h4001af55, 32'h3ba7c68a} /* (21, 11, 23) {real, imag} */,
  {32'hbf9e8b02, 32'h3f89fa6c} /* (21, 11, 22) {real, imag} */,
  {32'hbfce288d, 32'h3f2a85cb} /* (21, 11, 21) {real, imag} */,
  {32'hbf5cfb27, 32'hc055817a} /* (21, 11, 20) {real, imag} */,
  {32'h3f98cfe1, 32'h3f8d67a8} /* (21, 11, 19) {real, imag} */,
  {32'hbf4b492c, 32'h3e8394ef} /* (21, 11, 18) {real, imag} */,
  {32'h3f91a4ee, 32'h3faa22f9} /* (21, 11, 17) {real, imag} */,
  {32'hc03988b0, 32'hbf2bad5a} /* (21, 11, 16) {real, imag} */,
  {32'hbfac4646, 32'h3e893628} /* (21, 11, 15) {real, imag} */,
  {32'h3f238cc9, 32'hc0412045} /* (21, 11, 14) {real, imag} */,
  {32'h3f952d5f, 32'h3f80119b} /* (21, 11, 13) {real, imag} */,
  {32'h3ea04607, 32'hbf7f5c0d} /* (21, 11, 12) {real, imag} */,
  {32'h3f3ae74f, 32'hbcd4d463} /* (21, 11, 11) {real, imag} */,
  {32'h3c43e698, 32'hbf559711} /* (21, 11, 10) {real, imag} */,
  {32'h3f52848a, 32'hc041d91b} /* (21, 11, 9) {real, imag} */,
  {32'hc082256a, 32'h3fdc2df1} /* (21, 11, 8) {real, imag} */,
  {32'h3fda0558, 32'h408c08d7} /* (21, 11, 7) {real, imag} */,
  {32'h4019be4d, 32'hbf6d2101} /* (21, 11, 6) {real, imag} */,
  {32'hbf233742, 32'hbf5ca0ad} /* (21, 11, 5) {real, imag} */,
  {32'hc00fe600, 32'hbe00fc6d} /* (21, 11, 4) {real, imag} */,
  {32'h3f90de44, 32'h4082a857} /* (21, 11, 3) {real, imag} */,
  {32'h3e8a59f4, 32'h3f335ea3} /* (21, 11, 2) {real, imag} */,
  {32'hbfede088, 32'hc072fd80} /* (21, 11, 1) {real, imag} */,
  {32'hc05451b4, 32'hbdd798fc} /* (21, 11, 0) {real, imag} */,
  {32'hbdc51524, 32'h3f1dd81e} /* (21, 10, 31) {real, imag} */,
  {32'hbe42963b, 32'h3edf0e8e} /* (21, 10, 30) {real, imag} */,
  {32'h3f54e69d, 32'h3d4e4934} /* (21, 10, 29) {real, imag} */,
  {32'hbf9ea46b, 32'h3de9000b} /* (21, 10, 28) {real, imag} */,
  {32'hc015b03d, 32'h3f6d8f64} /* (21, 10, 27) {real, imag} */,
  {32'h4019d641, 32'hbfbc5da6} /* (21, 10, 26) {real, imag} */,
  {32'h3fc6ee77, 32'h3e224946} /* (21, 10, 25) {real, imag} */,
  {32'h4025fe29, 32'hc018bd47} /* (21, 10, 24) {real, imag} */,
  {32'hbfbd60a1, 32'h40853799} /* (21, 10, 23) {real, imag} */,
  {32'h400fb9a2, 32'hbb4c04ca} /* (21, 10, 22) {real, imag} */,
  {32'h4051a0fe, 32'h3de223a4} /* (21, 10, 21) {real, imag} */,
  {32'hc01919cf, 32'h3d92ef76} /* (21, 10, 20) {real, imag} */,
  {32'h3bec1200, 32'hc04707d4} /* (21, 10, 19) {real, imag} */,
  {32'hbfd1dadb, 32'hc079542e} /* (21, 10, 18) {real, imag} */,
  {32'hbdeadb31, 32'hc0386358} /* (21, 10, 17) {real, imag} */,
  {32'hbfd695ae, 32'h3e90e20d} /* (21, 10, 16) {real, imag} */,
  {32'hbf8f23ab, 32'hbc2d3de3} /* (21, 10, 15) {real, imag} */,
  {32'h40d7ca0c, 32'h400cbd9c} /* (21, 10, 14) {real, imag} */,
  {32'hbfc6462f, 32'hbf391e10} /* (21, 10, 13) {real, imag} */,
  {32'hbfd25fcf, 32'h3f515bc3} /* (21, 10, 12) {real, imag} */,
  {32'hbea4bb34, 32'h40682d15} /* (21, 10, 11) {real, imag} */,
  {32'hc011c1ed, 32'h3ea6cf04} /* (21, 10, 10) {real, imag} */,
  {32'hbf919346, 32'hc0a6873f} /* (21, 10, 9) {real, imag} */,
  {32'h406c8806, 32'hbef488bf} /* (21, 10, 8) {real, imag} */,
  {32'h40123e14, 32'hbe8b0d30} /* (21, 10, 7) {real, imag} */,
  {32'h400168e9, 32'hbfde995a} /* (21, 10, 6) {real, imag} */,
  {32'h4016321d, 32'hc00c3fe2} /* (21, 10, 5) {real, imag} */,
  {32'hc05d51f3, 32'hbf88c92e} /* (21, 10, 4) {real, imag} */,
  {32'hbf3bc425, 32'hbf82b209} /* (21, 10, 3) {real, imag} */,
  {32'h3e67205a, 32'h3fa1b924} /* (21, 10, 2) {real, imag} */,
  {32'h3e037d99, 32'h40508ad0} /* (21, 10, 1) {real, imag} */,
  {32'h3e6ddb65, 32'hbf4af8b7} /* (21, 10, 0) {real, imag} */,
  {32'hbfc19b09, 32'hbf9a80ec} /* (21, 9, 31) {real, imag} */,
  {32'hbfd62560, 32'hbed7b142} /* (21, 9, 30) {real, imag} */,
  {32'hbf010d53, 32'hc02ad08a} /* (21, 9, 29) {real, imag} */,
  {32'hbf1cd483, 32'h3f8cb578} /* (21, 9, 28) {real, imag} */,
  {32'hc007dfb1, 32'h4024a849} /* (21, 9, 27) {real, imag} */,
  {32'h3fb89bb5, 32'hbf76f4e5} /* (21, 9, 26) {real, imag} */,
  {32'h3f5bc071, 32'hbf9d0564} /* (21, 9, 25) {real, imag} */,
  {32'h402aad4a, 32'hc00ca745} /* (21, 9, 24) {real, imag} */,
  {32'h403251e5, 32'hbd8bfb28} /* (21, 9, 23) {real, imag} */,
  {32'h3e9f364a, 32'hbfc54be8} /* (21, 9, 22) {real, imag} */,
  {32'h3f424f2f, 32'h401499be} /* (21, 9, 21) {real, imag} */,
  {32'hbe487a3c, 32'h3f899311} /* (21, 9, 20) {real, imag} */,
  {32'h3e8a601e, 32'hbedf405f} /* (21, 9, 19) {real, imag} */,
  {32'h3ed69248, 32'hbe88f270} /* (21, 9, 18) {real, imag} */,
  {32'hbfa0b9d1, 32'hbf8b70a6} /* (21, 9, 17) {real, imag} */,
  {32'h3f9fa886, 32'hbf8adfe5} /* (21, 9, 16) {real, imag} */,
  {32'h3f40eb31, 32'h3f27ee3d} /* (21, 9, 15) {real, imag} */,
  {32'hc017b1c5, 32'hbe779884} /* (21, 9, 14) {real, imag} */,
  {32'hbff844ac, 32'h3f6b3a49} /* (21, 9, 13) {real, imag} */,
  {32'h3f2fd20a, 32'hbeec2c46} /* (21, 9, 12) {real, imag} */,
  {32'hc00ed613, 32'hbfe2d323} /* (21, 9, 11) {real, imag} */,
  {32'h40679e88, 32'h3fbaa108} /* (21, 9, 10) {real, imag} */,
  {32'h3ff2ceaa, 32'h3f95ce5f} /* (21, 9, 9) {real, imag} */,
  {32'h3fb1157f, 32'hbf9ada10} /* (21, 9, 8) {real, imag} */,
  {32'hc040e8cf, 32'hbfa6f180} /* (21, 9, 7) {real, imag} */,
  {32'h4012de66, 32'h400bb805} /* (21, 9, 6) {real, imag} */,
  {32'hbfff847f, 32'h3f50157f} /* (21, 9, 5) {real, imag} */,
  {32'hbfad79be, 32'h3f4c5cb3} /* (21, 9, 4) {real, imag} */,
  {32'h3ff9e434, 32'h3f50bcd7} /* (21, 9, 3) {real, imag} */,
  {32'hc089a4a9, 32'hc038df42} /* (21, 9, 2) {real, imag} */,
  {32'hbea189e9, 32'hbf3aa165} /* (21, 9, 1) {real, imag} */,
  {32'h3f5030f3, 32'h3f59839d} /* (21, 9, 0) {real, imag} */,
  {32'hbfe77675, 32'hc0313b07} /* (21, 8, 31) {real, imag} */,
  {32'h4039fa80, 32'hc015f877} /* (21, 8, 30) {real, imag} */,
  {32'h3f293640, 32'h3df639e2} /* (21, 8, 29) {real, imag} */,
  {32'h3feba00a, 32'h3f82c415} /* (21, 8, 28) {real, imag} */,
  {32'hbd9ec6ae, 32'hbf0ec493} /* (21, 8, 27) {real, imag} */,
  {32'h4092ace4, 32'h3f299312} /* (21, 8, 26) {real, imag} */,
  {32'h3fea5f36, 32'hc03b3f77} /* (21, 8, 25) {real, imag} */,
  {32'h3f5c39d6, 32'h3fe60143} /* (21, 8, 24) {real, imag} */,
  {32'hc071b6ce, 32'hbfcb1f17} /* (21, 8, 23) {real, imag} */,
  {32'hbf8c29a8, 32'hc01dccc4} /* (21, 8, 22) {real, imag} */,
  {32'hc0064ff7, 32'h3ee5eed4} /* (21, 8, 21) {real, imag} */,
  {32'hbf16c34c, 32'h3fa015a9} /* (21, 8, 20) {real, imag} */,
  {32'h400dd31e, 32'h3f264dc6} /* (21, 8, 19) {real, imag} */,
  {32'hbc72ff3e, 32'h3d7fead0} /* (21, 8, 18) {real, imag} */,
  {32'h3f7f651e, 32'h3eec671b} /* (21, 8, 17) {real, imag} */,
  {32'h3ffbc800, 32'hc00379a4} /* (21, 8, 16) {real, imag} */,
  {32'hbef6bbde, 32'h3ea7f38c} /* (21, 8, 15) {real, imag} */,
  {32'hbfc7af11, 32'h3fa9ebf1} /* (21, 8, 14) {real, imag} */,
  {32'h3f9d2f63, 32'h4034ca8a} /* (21, 8, 13) {real, imag} */,
  {32'hbfd5d893, 32'h3ed85da3} /* (21, 8, 12) {real, imag} */,
  {32'hbf277434, 32'hbec13ac8} /* (21, 8, 11) {real, imag} */,
  {32'h3fe28a2e, 32'hbf79a4cd} /* (21, 8, 10) {real, imag} */,
  {32'hbf291fbf, 32'hbf3b2c57} /* (21, 8, 9) {real, imag} */,
  {32'hc02e0f36, 32'h3f8d5f38} /* (21, 8, 8) {real, imag} */,
  {32'hbfee4717, 32'h404a005a} /* (21, 8, 7) {real, imag} */,
  {32'hc01f6497, 32'h3e304998} /* (21, 8, 6) {real, imag} */,
  {32'h4020c6ab, 32'h4005f7bf} /* (21, 8, 5) {real, imag} */,
  {32'h3ec1d27c, 32'hc02607da} /* (21, 8, 4) {real, imag} */,
  {32'h3fed146a, 32'h3fe78c4c} /* (21, 8, 3) {real, imag} */,
  {32'hc0352fbf, 32'hbf8d7557} /* (21, 8, 2) {real, imag} */,
  {32'hbf8a53dd, 32'h3e8b5795} /* (21, 8, 1) {real, imag} */,
  {32'hc028da7b, 32'hc0781ce6} /* (21, 8, 0) {real, imag} */,
  {32'hbfcf234a, 32'hbe3ceaf1} /* (21, 7, 31) {real, imag} */,
  {32'h3ebd8765, 32'h400d4bd3} /* (21, 7, 30) {real, imag} */,
  {32'hbeb10af1, 32'hbf05de76} /* (21, 7, 29) {real, imag} */,
  {32'h3fbc1b6f, 32'hbf7b4082} /* (21, 7, 28) {real, imag} */,
  {32'h3faa0a14, 32'h4050b501} /* (21, 7, 27) {real, imag} */,
  {32'hbff55492, 32'h40607e35} /* (21, 7, 26) {real, imag} */,
  {32'h3c77e64d, 32'hbfbaafa0} /* (21, 7, 25) {real, imag} */,
  {32'h40093f74, 32'h3fa333b4} /* (21, 7, 24) {real, imag} */,
  {32'hbfca6c59, 32'h3f6ff27d} /* (21, 7, 23) {real, imag} */,
  {32'h400b4ff4, 32'h4010af1f} /* (21, 7, 22) {real, imag} */,
  {32'h3e93e995, 32'hbf927bd0} /* (21, 7, 21) {real, imag} */,
  {32'hbc402298, 32'hc0148868} /* (21, 7, 20) {real, imag} */,
  {32'hbe305aa2, 32'h3f285b46} /* (21, 7, 19) {real, imag} */,
  {32'hbf542ffe, 32'hbe840576} /* (21, 7, 18) {real, imag} */,
  {32'hbfa87da8, 32'hc05b0ad6} /* (21, 7, 17) {real, imag} */,
  {32'h3c1b5c3e, 32'hbe2e4d97} /* (21, 7, 16) {real, imag} */,
  {32'h3fc48983, 32'hbfd0e187} /* (21, 7, 15) {real, imag} */,
  {32'hc027e368, 32'h3fe8397b} /* (21, 7, 14) {real, imag} */,
  {32'h3fc4e97c, 32'hbe96f887} /* (21, 7, 13) {real, imag} */,
  {32'h3ff9f5e6, 32'h40343801} /* (21, 7, 12) {real, imag} */,
  {32'hbe970d7a, 32'h3f664686} /* (21, 7, 11) {real, imag} */,
  {32'hbf8dba55, 32'hbfcac671} /* (21, 7, 10) {real, imag} */,
  {32'hbf88ca4b, 32'h3fd8de9a} /* (21, 7, 9) {real, imag} */,
  {32'h3f62445d, 32'hbfd50788} /* (21, 7, 8) {real, imag} */,
  {32'hbf801648, 32'hbf8c1dc2} /* (21, 7, 7) {real, imag} */,
  {32'hc019c08e, 32'hbf82fcc0} /* (21, 7, 6) {real, imag} */,
  {32'hbf69233d, 32'h3f95f1f6} /* (21, 7, 5) {real, imag} */,
  {32'hbe1911d6, 32'h3f1e1283} /* (21, 7, 4) {real, imag} */,
  {32'hbf7d5297, 32'hbfdb692b} /* (21, 7, 3) {real, imag} */,
  {32'hbd57cdce, 32'h3f3d7d17} /* (21, 7, 2) {real, imag} */,
  {32'h3faee9a2, 32'hbeab8811} /* (21, 7, 1) {real, imag} */,
  {32'h402da826, 32'hbf9d155c} /* (21, 7, 0) {real, imag} */,
  {32'hbf4ee889, 32'hbf83b6d5} /* (21, 6, 31) {real, imag} */,
  {32'hbf39d5e2, 32'h3fbfce76} /* (21, 6, 30) {real, imag} */,
  {32'hbfc1f9f6, 32'hbf73f99b} /* (21, 6, 29) {real, imag} */,
  {32'hbf489226, 32'h3f8b891a} /* (21, 6, 28) {real, imag} */,
  {32'hc01fdad9, 32'h3fe06dd5} /* (21, 6, 27) {real, imag} */,
  {32'h3ff3c7da, 32'h3f6f921f} /* (21, 6, 26) {real, imag} */,
  {32'hbe8970be, 32'hbe48885a} /* (21, 6, 25) {real, imag} */,
  {32'h3fd04e4b, 32'h40258abc} /* (21, 6, 24) {real, imag} */,
  {32'h408e64c6, 32'hc0170aae} /* (21, 6, 23) {real, imag} */,
  {32'hbe83a1d5, 32'hbffe6399} /* (21, 6, 22) {real, imag} */,
  {32'hbfa04c97, 32'hbf8d7eb7} /* (21, 6, 21) {real, imag} */,
  {32'h3faa35f3, 32'h3f0d7a07} /* (21, 6, 20) {real, imag} */,
  {32'h3f974f0b, 32'hbfc6dc76} /* (21, 6, 19) {real, imag} */,
  {32'h3f7266ca, 32'h4033b1f9} /* (21, 6, 18) {real, imag} */,
  {32'hc0105395, 32'h3dee13bd} /* (21, 6, 17) {real, imag} */,
  {32'hbf83ed89, 32'hbf1abcc5} /* (21, 6, 16) {real, imag} */,
  {32'h3fce4aec, 32'hbfb7972f} /* (21, 6, 15) {real, imag} */,
  {32'hbfd7acbd, 32'h404459eb} /* (21, 6, 14) {real, imag} */,
  {32'hbfb65090, 32'hbfa330b8} /* (21, 6, 13) {real, imag} */,
  {32'hbfe9e36a, 32'hbf805d12} /* (21, 6, 12) {real, imag} */,
  {32'h401fde3a, 32'hc02834bb} /* (21, 6, 11) {real, imag} */,
  {32'h3eb9e07c, 32'h3e89484b} /* (21, 6, 10) {real, imag} */,
  {32'hbed45004, 32'h3fcade5b} /* (21, 6, 9) {real, imag} */,
  {32'hbf31d009, 32'hbf054ec7} /* (21, 6, 8) {real, imag} */,
  {32'h401e4945, 32'h3ff17769} /* (21, 6, 7) {real, imag} */,
  {32'h3f8ba47b, 32'h3f3ad1c9} /* (21, 6, 6) {real, imag} */,
  {32'h3f7e8e95, 32'h3e032cc2} /* (21, 6, 5) {real, imag} */,
  {32'h401ea4b3, 32'hc0183878} /* (21, 6, 4) {real, imag} */,
  {32'hbfc437fe, 32'hc0212fd7} /* (21, 6, 3) {real, imag} */,
  {32'hc0424c84, 32'h40814888} /* (21, 6, 2) {real, imag} */,
  {32'h3f13ffe0, 32'h40115396} /* (21, 6, 1) {real, imag} */,
  {32'h3fe89fa9, 32'hbffe36d9} /* (21, 6, 0) {real, imag} */,
  {32'hbfa278ea, 32'hbe6ec5bf} /* (21, 5, 31) {real, imag} */,
  {32'h3f5bfd40, 32'h40c81473} /* (21, 5, 30) {real, imag} */,
  {32'h3ecaa699, 32'hbf27117f} /* (21, 5, 29) {real, imag} */,
  {32'hbf9ae26f, 32'h3f88c8f0} /* (21, 5, 28) {real, imag} */,
  {32'hbf2d5ede, 32'h402688e7} /* (21, 5, 27) {real, imag} */,
  {32'hbec2dffb, 32'hc0388d54} /* (21, 5, 26) {real, imag} */,
  {32'hbf81058c, 32'hc00541ce} /* (21, 5, 25) {real, imag} */,
  {32'h4010b269, 32'h3f726876} /* (21, 5, 24) {real, imag} */,
  {32'h3fb1239d, 32'hbefca579} /* (21, 5, 23) {real, imag} */,
  {32'hbfc8f11c, 32'h3fbef702} /* (21, 5, 22) {real, imag} */,
  {32'hbf501f22, 32'hbf8e129c} /* (21, 5, 21) {real, imag} */,
  {32'h3f896299, 32'h3e494646} /* (21, 5, 20) {real, imag} */,
  {32'h3fa7cc68, 32'h3f264d32} /* (21, 5, 19) {real, imag} */,
  {32'hbeb4563d, 32'h3d2ee610} /* (21, 5, 18) {real, imag} */,
  {32'hbf81989c, 32'hbdc697ef} /* (21, 5, 17) {real, imag} */,
  {32'h3f8de73f, 32'hbe31052b} /* (21, 5, 16) {real, imag} */,
  {32'h4022bf37, 32'hc032b069} /* (21, 5, 15) {real, imag} */,
  {32'h3f07d474, 32'hbfa816ed} /* (21, 5, 14) {real, imag} */,
  {32'h3f0982a6, 32'h3f74a8dc} /* (21, 5, 13) {real, imag} */,
  {32'hbf6fda95, 32'hbf8e8fd7} /* (21, 5, 12) {real, imag} */,
  {32'h3e22f85c, 32'hbfcf3278} /* (21, 5, 11) {real, imag} */,
  {32'h3f12ed63, 32'h402a7645} /* (21, 5, 10) {real, imag} */,
  {32'h3fc19e79, 32'hbf1c8a02} /* (21, 5, 9) {real, imag} */,
  {32'h403c8678, 32'hc00ba7ba} /* (21, 5, 8) {real, imag} */,
  {32'hbf721d35, 32'h4073ab55} /* (21, 5, 7) {real, imag} */,
  {32'hc009dd13, 32'hbf483e96} /* (21, 5, 6) {real, imag} */,
  {32'h409e58d0, 32'hbcc8abc0} /* (21, 5, 5) {real, imag} */,
  {32'h3f46c7bb, 32'h3b2d54c4} /* (21, 5, 4) {real, imag} */,
  {32'hbf833dcd, 32'h3fe8ff2d} /* (21, 5, 3) {real, imag} */,
  {32'hc0205958, 32'h3f8f8026} /* (21, 5, 2) {real, imag} */,
  {32'hbf78dcca, 32'hc05e1db4} /* (21, 5, 1) {real, imag} */,
  {32'hc00bf33f, 32'hc07bab26} /* (21, 5, 0) {real, imag} */,
  {32'hbeaaae75, 32'hbf8c4df0} /* (21, 4, 31) {real, imag} */,
  {32'hc038a00a, 32'hbfbab1a2} /* (21, 4, 30) {real, imag} */,
  {32'h40215f82, 32'h40c8eaad} /* (21, 4, 29) {real, imag} */,
  {32'hbe92b84b, 32'h3eb1e73a} /* (21, 4, 28) {real, imag} */,
  {32'h3f47aa35, 32'hbf83aab5} /* (21, 4, 27) {real, imag} */,
  {32'hbef32d36, 32'h3fb03a64} /* (21, 4, 26) {real, imag} */,
  {32'h3f9393b5, 32'h4024a071} /* (21, 4, 25) {real, imag} */,
  {32'hc00916d9, 32'hbf40303d} /* (21, 4, 24) {real, imag} */,
  {32'hc0380ff5, 32'h3d9a7091} /* (21, 4, 23) {real, imag} */,
  {32'hbf1b7678, 32'h3eaf19ad} /* (21, 4, 22) {real, imag} */,
  {32'h3f952543, 32'h3f21c53a} /* (21, 4, 21) {real, imag} */,
  {32'h3f9c17eb, 32'h3cd9a37d} /* (21, 4, 20) {real, imag} */,
  {32'hbff91a98, 32'hc00dec83} /* (21, 4, 19) {real, imag} */,
  {32'hbff51eac, 32'h3ef3a6fb} /* (21, 4, 18) {real, imag} */,
  {32'hbdb639d4, 32'h3f1baa11} /* (21, 4, 17) {real, imag} */,
  {32'h3fc65444, 32'hc01d21b7} /* (21, 4, 16) {real, imag} */,
  {32'hbfb336a1, 32'h3f6819f9} /* (21, 4, 15) {real, imag} */,
  {32'h3e6c4241, 32'hc014ad45} /* (21, 4, 14) {real, imag} */,
  {32'h3fc53a46, 32'h3e87f9be} /* (21, 4, 13) {real, imag} */,
  {32'hbf7c08f7, 32'hbd3beb02} /* (21, 4, 12) {real, imag} */,
  {32'hbe219331, 32'h3ece53c7} /* (21, 4, 11) {real, imag} */,
  {32'h3fdcb2db, 32'h40149bb1} /* (21, 4, 10) {real, imag} */,
  {32'h3f74b8d5, 32'h3fc9bbe3} /* (21, 4, 9) {real, imag} */,
  {32'hc02a1d49, 32'hc010fbe4} /* (21, 4, 8) {real, imag} */,
  {32'hbea9d152, 32'h3ebd99b6} /* (21, 4, 7) {real, imag} */,
  {32'h40310f3c, 32'h3ff3be31} /* (21, 4, 6) {real, imag} */,
  {32'h3f179caf, 32'h3fe5291f} /* (21, 4, 5) {real, imag} */,
  {32'hbf6e99b9, 32'h3f17f5ea} /* (21, 4, 4) {real, imag} */,
  {32'hbf168378, 32'h400dfd6e} /* (21, 4, 3) {real, imag} */,
  {32'h4080b98a, 32'h3fa2c832} /* (21, 4, 2) {real, imag} */,
  {32'h40251210, 32'hbe89a83f} /* (21, 4, 1) {real, imag} */,
  {32'h3dd1aaa8, 32'h3ce1bf18} /* (21, 4, 0) {real, imag} */,
  {32'hbfa6026e, 32'h3fabbd61} /* (21, 3, 31) {real, imag} */,
  {32'hbf173548, 32'hc0a27ce9} /* (21, 3, 30) {real, imag} */,
  {32'h3f83957a, 32'hbf2a578b} /* (21, 3, 29) {real, imag} */,
  {32'h3f00c68d, 32'h3f8740e5} /* (21, 3, 28) {real, imag} */,
  {32'h3fa85e94, 32'h3fbe2077} /* (21, 3, 27) {real, imag} */,
  {32'hbfade4da, 32'h3ff2a325} /* (21, 3, 26) {real, imag} */,
  {32'h3efcc359, 32'hc0801f8d} /* (21, 3, 25) {real, imag} */,
  {32'hbf9d3e5b, 32'hbf8899cd} /* (21, 3, 24) {real, imag} */,
  {32'hc03aff3b, 32'hbf1c1796} /* (21, 3, 23) {real, imag} */,
  {32'h4053f38d, 32'hbe3b7bc2} /* (21, 3, 22) {real, imag} */,
  {32'hbf099d38, 32'h3f1c3599} /* (21, 3, 21) {real, imag} */,
  {32'h3ea1ee2a, 32'h3eb25c1d} /* (21, 3, 20) {real, imag} */,
  {32'h40494c70, 32'h3f5409d6} /* (21, 3, 19) {real, imag} */,
  {32'hc01d6236, 32'hbef5cca6} /* (21, 3, 18) {real, imag} */,
  {32'h3f60e435, 32'h3efd576f} /* (21, 3, 17) {real, imag} */,
  {32'h40099b8e, 32'h40683d14} /* (21, 3, 16) {real, imag} */,
  {32'hbfdb0a9e, 32'h3fdb2446} /* (21, 3, 15) {real, imag} */,
  {32'h3f0204b1, 32'h3de6bd76} /* (21, 3, 14) {real, imag} */,
  {32'h3f6191b7, 32'hbf7e3f42} /* (21, 3, 13) {real, imag} */,
  {32'hbfef3af6, 32'h402160c9} /* (21, 3, 12) {real, imag} */,
  {32'hbfa51f87, 32'h3e92572b} /* (21, 3, 11) {real, imag} */,
  {32'h3fb56989, 32'hbd0cad65} /* (21, 3, 10) {real, imag} */,
  {32'hbe2c7502, 32'h3fcca917} /* (21, 3, 9) {real, imag} */,
  {32'hbf8762d6, 32'hc03c14cc} /* (21, 3, 8) {real, imag} */,
  {32'hbe3bdabf, 32'hbfa4b883} /* (21, 3, 7) {real, imag} */,
  {32'h3fa2e90c, 32'h3ecc368e} /* (21, 3, 6) {real, imag} */,
  {32'h40505f52, 32'h4001d162} /* (21, 3, 5) {real, imag} */,
  {32'h3ea4c835, 32'h3ff31295} /* (21, 3, 4) {real, imag} */,
  {32'hbf7c124b, 32'h3ede4d2d} /* (21, 3, 3) {real, imag} */,
  {32'h4006b267, 32'hc082c047} /* (21, 3, 2) {real, imag} */,
  {32'h3f23713e, 32'h40663582} /* (21, 3, 1) {real, imag} */,
  {32'h3f42c461, 32'hbfd6417d} /* (21, 3, 0) {real, imag} */,
  {32'hc0e5e651, 32'hc0385c2b} /* (21, 2, 31) {real, imag} */,
  {32'h40ce527a, 32'h40570112} /* (21, 2, 30) {real, imag} */,
  {32'hc0531f70, 32'hbf89e528} /* (21, 2, 29) {real, imag} */,
  {32'hbfd7a324, 32'h3feba21c} /* (21, 2, 28) {real, imag} */,
  {32'h3ca342ec, 32'h3f173b72} /* (21, 2, 27) {real, imag} */,
  {32'hbfe53fd2, 32'hbeb2b38f} /* (21, 2, 26) {real, imag} */,
  {32'h401ea008, 32'hbe98dcf5} /* (21, 2, 25) {real, imag} */,
  {32'h3ff0e6cf, 32'h3f361612} /* (21, 2, 24) {real, imag} */,
  {32'hc008b163, 32'hbe664720} /* (21, 2, 23) {real, imag} */,
  {32'h3e13c68c, 32'h3f60b813} /* (21, 2, 22) {real, imag} */,
  {32'hbf29312b, 32'h3fcc6859} /* (21, 2, 21) {real, imag} */,
  {32'hc07a3c42, 32'hbf40a828} /* (21, 2, 20) {real, imag} */,
  {32'h3fe9605b, 32'hbf17097e} /* (21, 2, 19) {real, imag} */,
  {32'h3e465f8f, 32'hbf19c5c5} /* (21, 2, 18) {real, imag} */,
  {32'h3dfc6892, 32'h3fc34112} /* (21, 2, 17) {real, imag} */,
  {32'h3e396810, 32'hbf5f404f} /* (21, 2, 16) {real, imag} */,
  {32'h3ffe40fe, 32'hbfc9ceaf} /* (21, 2, 15) {real, imag} */,
  {32'h3f8ab6ef, 32'h400cb573} /* (21, 2, 14) {real, imag} */,
  {32'h3f99dbcd, 32'hc00d20bf} /* (21, 2, 13) {real, imag} */,
  {32'h3f3bef51, 32'h3f755526} /* (21, 2, 12) {real, imag} */,
  {32'hbf015a47, 32'h40143a9c} /* (21, 2, 11) {real, imag} */,
  {32'h4067aea7, 32'hbfd7793e} /* (21, 2, 10) {real, imag} */,
  {32'h400011e6, 32'h3f531346} /* (21, 2, 9) {real, imag} */,
  {32'h3fb713c1, 32'h3fd51014} /* (21, 2, 8) {real, imag} */,
  {32'h3f3875f0, 32'h3ff3d1ad} /* (21, 2, 7) {real, imag} */,
  {32'h3f876722, 32'h409ab441} /* (21, 2, 6) {real, imag} */,
  {32'hbf8ca14a, 32'h3f81892f} /* (21, 2, 5) {real, imag} */,
  {32'h405c2168, 32'hbfe952fb} /* (21, 2, 4) {real, imag} */,
  {32'hbfadb355, 32'h4014893c} /* (21, 2, 3) {real, imag} */,
  {32'h408cb9d4, 32'h3e767f08} /* (21, 2, 2) {real, imag} */,
  {32'hc017d342, 32'hc02f2403} /* (21, 2, 1) {real, imag} */,
  {32'hbf9aa279, 32'hc0821432} /* (21, 2, 0) {real, imag} */,
  {32'h402ddff7, 32'h3f9d6480} /* (21, 1, 31) {real, imag} */,
  {32'h3fb0dd0e, 32'hc0985605} /* (21, 1, 30) {real, imag} */,
  {32'h4001c368, 32'h401509b6} /* (21, 1, 29) {real, imag} */,
  {32'h3a089aef, 32'h404ec705} /* (21, 1, 28) {real, imag} */,
  {32'hbf267b66, 32'hc084381d} /* (21, 1, 27) {real, imag} */,
  {32'h401ddf82, 32'hbfca6630} /* (21, 1, 26) {real, imag} */,
  {32'h3f2a2d00, 32'h3fbe33af} /* (21, 1, 25) {real, imag} */,
  {32'hbfe09173, 32'h3d2d9d22} /* (21, 1, 24) {real, imag} */,
  {32'h40346c75, 32'hc03f3a4f} /* (21, 1, 23) {real, imag} */,
  {32'h3f94d4c4, 32'h402cef25} /* (21, 1, 22) {real, imag} */,
  {32'hc020162f, 32'h3fd3e53b} /* (21, 1, 21) {real, imag} */,
  {32'hc0225ee3, 32'hbf04801f} /* (21, 1, 20) {real, imag} */,
  {32'h3f8aeb02, 32'h401e6750} /* (21, 1, 19) {real, imag} */,
  {32'hc02ad555, 32'hbd35ae47} /* (21, 1, 18) {real, imag} */,
  {32'h3fceaf83, 32'h3fab20e7} /* (21, 1, 17) {real, imag} */,
  {32'h3f1ebaee, 32'hbf3088d2} /* (21, 1, 16) {real, imag} */,
  {32'h3f5b8332, 32'hbfe1e5d1} /* (21, 1, 15) {real, imag} */,
  {32'hbefb475a, 32'hc043df99} /* (21, 1, 14) {real, imag} */,
  {32'h4019a6a4, 32'hbf9c9810} /* (21, 1, 13) {real, imag} */,
  {32'hbd8f2125, 32'hbf05d54f} /* (21, 1, 12) {real, imag} */,
  {32'h3f1ac058, 32'hc051e020} /* (21, 1, 11) {real, imag} */,
  {32'hc02fa291, 32'hbff3ec37} /* (21, 1, 10) {real, imag} */,
  {32'hc0152c14, 32'h3fb848c1} /* (21, 1, 9) {real, imag} */,
  {32'h3fb2f58c, 32'hbf1f4fc9} /* (21, 1, 8) {real, imag} */,
  {32'h40478fc3, 32'h400295ad} /* (21, 1, 7) {real, imag} */,
  {32'h3fff5d0f, 32'hbf605648} /* (21, 1, 6) {real, imag} */,
  {32'hbf9bdb95, 32'h3f524e95} /* (21, 1, 5) {real, imag} */,
  {32'hc06d7c55, 32'h4086522e} /* (21, 1, 4) {real, imag} */,
  {32'hbe3879a0, 32'hbfaa4256} /* (21, 1, 3) {real, imag} */,
  {32'hc0224b97, 32'hc1112e0f} /* (21, 1, 2) {real, imag} */,
  {32'h40a48cfd, 32'h40babc42} /* (21, 1, 1) {real, imag} */,
  {32'h409c9c9d, 32'h40fb8d1d} /* (21, 1, 0) {real, imag} */,
  {32'h40a302b6, 32'h402ec925} /* (21, 0, 31) {real, imag} */,
  {32'hbf91f44e, 32'h409baedb} /* (21, 0, 30) {real, imag} */,
  {32'h3fa9a847, 32'h3da83f92} /* (21, 0, 29) {real, imag} */,
  {32'h40390405, 32'h3f022669} /* (21, 0, 28) {real, imag} */,
  {32'h3fa88b87, 32'hbfda968b} /* (21, 0, 27) {real, imag} */,
  {32'hbf9636ae, 32'h3eae3df9} /* (21, 0, 26) {real, imag} */,
  {32'h3fc91117, 32'h4026aa7a} /* (21, 0, 25) {real, imag} */,
  {32'hbfb26c67, 32'hbf63d9a4} /* (21, 0, 24) {real, imag} */,
  {32'hbfc8817d, 32'h3fdfc8f6} /* (21, 0, 23) {real, imag} */,
  {32'hbf6d346d, 32'h3f0aa7b9} /* (21, 0, 22) {real, imag} */,
  {32'hbee0a41d, 32'h3f86f5d9} /* (21, 0, 21) {real, imag} */,
  {32'h3f0fac48, 32'h3fc0e668} /* (21, 0, 20) {real, imag} */,
  {32'hc01543e0, 32'h3ff8fd3d} /* (21, 0, 19) {real, imag} */,
  {32'h3d8dd622, 32'h406ba86e} /* (21, 0, 18) {real, imag} */,
  {32'hbf6294db, 32'hbf1e354e} /* (21, 0, 17) {real, imag} */,
  {32'h3f5d8d92, 32'h3f973574} /* (21, 0, 16) {real, imag} */,
  {32'hbf59dc98, 32'h3fdb4f82} /* (21, 0, 15) {real, imag} */,
  {32'h3f5a4a53, 32'h3ebedea8} /* (21, 0, 14) {real, imag} */,
  {32'hbf74d1a2, 32'h3ec3865f} /* (21, 0, 13) {real, imag} */,
  {32'h3f6b7c4a, 32'h3f0d8289} /* (21, 0, 12) {real, imag} */,
  {32'h3f5786da, 32'hbfede211} /* (21, 0, 11) {real, imag} */,
  {32'hbf53d1b6, 32'hbfde753f} /* (21, 0, 10) {real, imag} */,
  {32'hc037921e, 32'hc075a332} /* (21, 0, 9) {real, imag} */,
  {32'h408d1cc1, 32'hc0d7b5e2} /* (21, 0, 8) {real, imag} */,
  {32'hbf125de9, 32'hbed12ea8} /* (21, 0, 7) {real, imag} */,
  {32'h3f8cfe43, 32'h3ecb5782} /* (21, 0, 6) {real, imag} */,
  {32'hc0375c99, 32'h400cbb08} /* (21, 0, 5) {real, imag} */,
  {32'h3f28e0fe, 32'h3f213ad3} /* (21, 0, 4) {real, imag} */,
  {32'h3fb14fca, 32'hc088222d} /* (21, 0, 3) {real, imag} */,
  {32'h408e33fc, 32'hbed6407a} /* (21, 0, 2) {real, imag} */,
  {32'h403b2e35, 32'h40a67a93} /* (21, 0, 1) {real, imag} */,
  {32'h4094392b, 32'h402b81b0} /* (21, 0, 0) {real, imag} */,
  {32'h3f88e6e3, 32'hbc7f6f40} /* (20, 31, 31) {real, imag} */,
  {32'h400d5587, 32'h3fcc1124} /* (20, 31, 30) {real, imag} */,
  {32'h3fc8b5a5, 32'hbfb1eb00} /* (20, 31, 29) {real, imag} */,
  {32'hc06959f4, 32'hbf2b9f14} /* (20, 31, 28) {real, imag} */,
  {32'hbeb041a4, 32'hc0281ea9} /* (20, 31, 27) {real, imag} */,
  {32'hbe9b6a59, 32'hc01a6eac} /* (20, 31, 26) {real, imag} */,
  {32'hbf1a5f26, 32'hbfc5e4ac} /* (20, 31, 25) {real, imag} */,
  {32'h40302fff, 32'hbfc78066} /* (20, 31, 24) {real, imag} */,
  {32'hbf9ed500, 32'hbf81ce74} /* (20, 31, 23) {real, imag} */,
  {32'hbf327edf, 32'h3fc2277d} /* (20, 31, 22) {real, imag} */,
  {32'h3fc50994, 32'h400c6ed7} /* (20, 31, 21) {real, imag} */,
  {32'hbfe05357, 32'hbfc58625} /* (20, 31, 20) {real, imag} */,
  {32'h3fd84387, 32'h3f30dd3f} /* (20, 31, 19) {real, imag} */,
  {32'h3e10b2bf, 32'h3e795db6} /* (20, 31, 18) {real, imag} */,
  {32'h3ec65d0e, 32'hbf5e8d3d} /* (20, 31, 17) {real, imag} */,
  {32'h3fa9a920, 32'hbeccb87b} /* (20, 31, 16) {real, imag} */,
  {32'h3fabb085, 32'h3f02bdd9} /* (20, 31, 15) {real, imag} */,
  {32'hbf4d1c74, 32'h3e984437} /* (20, 31, 14) {real, imag} */,
  {32'h3d8a8ca6, 32'h3fc86757} /* (20, 31, 13) {real, imag} */,
  {32'hc0022e3a, 32'h400676a3} /* (20, 31, 12) {real, imag} */,
  {32'h3f3c4f9c, 32'hbf70a06c} /* (20, 31, 11) {real, imag} */,
  {32'hbf50bbd2, 32'hbffe8608} /* (20, 31, 10) {real, imag} */,
  {32'h3f499a36, 32'h3f1cb28c} /* (20, 31, 9) {real, imag} */,
  {32'hbf65f51f, 32'hbfbe32a7} /* (20, 31, 8) {real, imag} */,
  {32'h3f4e3952, 32'hbeec5c11} /* (20, 31, 7) {real, imag} */,
  {32'hbff79a61, 32'h3fa77511} /* (20, 31, 6) {real, imag} */,
  {32'hc04352a0, 32'h3f3839c0} /* (20, 31, 5) {real, imag} */,
  {32'hc05721c9, 32'hbfd63ebf} /* (20, 31, 4) {real, imag} */,
  {32'h3e9c6fa6, 32'hbd415fe3} /* (20, 31, 3) {real, imag} */,
  {32'h402a2e88, 32'h3f175360} /* (20, 31, 2) {real, imag} */,
  {32'hbfab8a9f, 32'h3c382ecc} /* (20, 31, 1) {real, imag} */,
  {32'h4008c1e6, 32'hbe0dbdf0} /* (20, 31, 0) {real, imag} */,
  {32'h3fce5582, 32'hc039435c} /* (20, 30, 31) {real, imag} */,
  {32'hbf78a9c6, 32'hc01e8d08} /* (20, 30, 30) {real, imag} */,
  {32'h3f7ada9b, 32'h3fe4b5a6} /* (20, 30, 29) {real, imag} */,
  {32'hbe4edb86, 32'h4014c007} /* (20, 30, 28) {real, imag} */,
  {32'hbf79b789, 32'hbf92019c} /* (20, 30, 27) {real, imag} */,
  {32'h403d5a6e, 32'hc014f162} /* (20, 30, 26) {real, imag} */,
  {32'h3ef95b07, 32'h407444ba} /* (20, 30, 25) {real, imag} */,
  {32'hc0037745, 32'h40419849} /* (20, 30, 24) {real, imag} */,
  {32'h3de329d9, 32'h400ae267} /* (20, 30, 23) {real, imag} */,
  {32'hbfc8fe2f, 32'h3fa60e4c} /* (20, 30, 22) {real, imag} */,
  {32'h3f2d9c3d, 32'h3f4be5bf} /* (20, 30, 21) {real, imag} */,
  {32'hc0347969, 32'hbfa65353} /* (20, 30, 20) {real, imag} */,
  {32'h3fb49cbd, 32'h3e9eb972} /* (20, 30, 19) {real, imag} */,
  {32'h3f713faf, 32'h40408275} /* (20, 30, 18) {real, imag} */,
  {32'hbf228023, 32'h3f270d47} /* (20, 30, 17) {real, imag} */,
  {32'h3ea94a27, 32'h3e6f35e8} /* (20, 30, 16) {real, imag} */,
  {32'h401f878f, 32'hbf9510de} /* (20, 30, 15) {real, imag} */,
  {32'hc00b70fe, 32'hc010620f} /* (20, 30, 14) {real, imag} */,
  {32'hbf7f723d, 32'h3f966ca6} /* (20, 30, 13) {real, imag} */,
  {32'h3d8b3bf5, 32'h3fd84507} /* (20, 30, 12) {real, imag} */,
  {32'h3eca87d9, 32'hc0709cda} /* (20, 30, 11) {real, imag} */,
  {32'hc00799a9, 32'h400abb6d} /* (20, 30, 10) {real, imag} */,
  {32'hbfff5adf, 32'h3e710394} /* (20, 30, 9) {real, imag} */,
  {32'h3f76ec04, 32'hc00df0a4} /* (20, 30, 8) {real, imag} */,
  {32'h3e8abad0, 32'h3f088b96} /* (20, 30, 7) {real, imag} */,
  {32'hc0874c12, 32'h3f822b0d} /* (20, 30, 6) {real, imag} */,
  {32'h40034cc7, 32'hbeb9a7d2} /* (20, 30, 5) {real, imag} */,
  {32'h3fbfb0da, 32'h3f92548e} /* (20, 30, 4) {real, imag} */,
  {32'hbfcf12e3, 32'hbfe50ac9} /* (20, 30, 3) {real, imag} */,
  {32'hbf61fcec, 32'hbf7bd3ef} /* (20, 30, 2) {real, imag} */,
  {32'h3dac474e, 32'h402c9139} /* (20, 30, 1) {real, imag} */,
  {32'hbf424646, 32'hbf14e922} /* (20, 30, 0) {real, imag} */,
  {32'hbf72485c, 32'h3fa9fd36} /* (20, 29, 31) {real, imag} */,
  {32'h402b599a, 32'h3f0c9970} /* (20, 29, 30) {real, imag} */,
  {32'hc061cab9, 32'hbfec3c28} /* (20, 29, 29) {real, imag} */,
  {32'h3f2d2d22, 32'h3e57bbae} /* (20, 29, 28) {real, imag} */,
  {32'h3e81ca2d, 32'hc00419c6} /* (20, 29, 27) {real, imag} */,
  {32'hbf1f20bc, 32'h4049b5e3} /* (20, 29, 26) {real, imag} */,
  {32'hbfb038de, 32'h3f981aa7} /* (20, 29, 25) {real, imag} */,
  {32'h3f9db46a, 32'hbe78340e} /* (20, 29, 24) {real, imag} */,
  {32'hbd4b455a, 32'h40384f3a} /* (20, 29, 23) {real, imag} */,
  {32'h3dc00796, 32'hbfaac7be} /* (20, 29, 22) {real, imag} */,
  {32'h403664d5, 32'h3cadfcb6} /* (20, 29, 21) {real, imag} */,
  {32'hbe02e0d2, 32'h3ee312ae} /* (20, 29, 20) {real, imag} */,
  {32'h3e4ee5e9, 32'hbe152e94} /* (20, 29, 19) {real, imag} */,
  {32'hbfdb2a4d, 32'h3dd59ae7} /* (20, 29, 18) {real, imag} */,
  {32'h3ffc3e31, 32'hc029b8d6} /* (20, 29, 17) {real, imag} */,
  {32'h3d92112d, 32'hbfc99ff7} /* (20, 29, 16) {real, imag} */,
  {32'hbf7dc35d, 32'hbfb9b6de} /* (20, 29, 15) {real, imag} */,
  {32'h3fd2c13f, 32'hbea08ccb} /* (20, 29, 14) {real, imag} */,
  {32'h3fba5958, 32'hbf1ac303} /* (20, 29, 13) {real, imag} */,
  {32'h3f5a8c4d, 32'h3f6d0ac6} /* (20, 29, 12) {real, imag} */,
  {32'h40525502, 32'hc017bf80} /* (20, 29, 11) {real, imag} */,
  {32'h3f9423d2, 32'h3e7c1963} /* (20, 29, 10) {real, imag} */,
  {32'h3e4225a4, 32'hbee559da} /* (20, 29, 9) {real, imag} */,
  {32'h3f40cdf3, 32'h3f03564f} /* (20, 29, 8) {real, imag} */,
  {32'hbee9a6c1, 32'h3f978a46} /* (20, 29, 7) {real, imag} */,
  {32'h3f81dd1e, 32'h3edcd278} /* (20, 29, 6) {real, imag} */,
  {32'hbfadd8de, 32'h3f2ae5da} /* (20, 29, 5) {real, imag} */,
  {32'hbfb1a083, 32'hc040b8a8} /* (20, 29, 4) {real, imag} */,
  {32'h3fb9425c, 32'h3f90bad8} /* (20, 29, 3) {real, imag} */,
  {32'hbfe19be8, 32'hbee7a972} /* (20, 29, 2) {real, imag} */,
  {32'h404a734b, 32'h3f823454} /* (20, 29, 1) {real, imag} */,
  {32'h3fc8f89a, 32'hbcdcd572} /* (20, 29, 0) {real, imag} */,
  {32'h3fd33fe9, 32'hbce466d0} /* (20, 28, 31) {real, imag} */,
  {32'h3e7c9985, 32'hc01d3901} /* (20, 28, 30) {real, imag} */,
  {32'h3fe8ee78, 32'hbf84aa7b} /* (20, 28, 29) {real, imag} */,
  {32'hbf90a112, 32'h3f032f17} /* (20, 28, 28) {real, imag} */,
  {32'hbf3c1074, 32'hc053928b} /* (20, 28, 27) {real, imag} */,
  {32'h3f66ef2f, 32'h3f9168e2} /* (20, 28, 26) {real, imag} */,
  {32'hbdd8e6b2, 32'h3fa00466} /* (20, 28, 25) {real, imag} */,
  {32'h404c08f7, 32'hbf42f251} /* (20, 28, 24) {real, imag} */,
  {32'h3fa2da65, 32'h3f9a52e4} /* (20, 28, 23) {real, imag} */,
  {32'h3fc1b747, 32'hbf8fca49} /* (20, 28, 22) {real, imag} */,
  {32'h3f103b26, 32'hc04b2eac} /* (20, 28, 21) {real, imag} */,
  {32'h3db989a1, 32'hbef9e80f} /* (20, 28, 20) {real, imag} */,
  {32'h3c8d087b, 32'h3ec7c17c} /* (20, 28, 19) {real, imag} */,
  {32'h3de92f93, 32'hbe8b04f3} /* (20, 28, 18) {real, imag} */,
  {32'h3e986cca, 32'h400154b4} /* (20, 28, 17) {real, imag} */,
  {32'h3e2a3758, 32'h3f479526} /* (20, 28, 16) {real, imag} */,
  {32'hbbd4998d, 32'hbdf796a5} /* (20, 28, 15) {real, imag} */,
  {32'hbeefc9e4, 32'h4071ce35} /* (20, 28, 14) {real, imag} */,
  {32'hc011a5e3, 32'hbf7f8585} /* (20, 28, 13) {real, imag} */,
  {32'hc0286788, 32'hbfa20209} /* (20, 28, 12) {real, imag} */,
  {32'h406186b9, 32'h3eb21419} /* (20, 28, 11) {real, imag} */,
  {32'hbf8999eb, 32'hbf8e79c7} /* (20, 28, 10) {real, imag} */,
  {32'h4017c7fd, 32'h3f322b80} /* (20, 28, 9) {real, imag} */,
  {32'h3f4d8bca, 32'hbf67341e} /* (20, 28, 8) {real, imag} */,
  {32'hbf3ca5a8, 32'hbe42904a} /* (20, 28, 7) {real, imag} */,
  {32'h3f462836, 32'h3f0b4c6d} /* (20, 28, 6) {real, imag} */,
  {32'h3fb6d2dd, 32'h3f59475f} /* (20, 28, 5) {real, imag} */,
  {32'hc0184694, 32'hc067c80f} /* (20, 28, 4) {real, imag} */,
  {32'hc039f364, 32'hbfebf440} /* (20, 28, 3) {real, imag} */,
  {32'h3f406762, 32'h402ad6c4} /* (20, 28, 2) {real, imag} */,
  {32'h3e989e6a, 32'h3f0f8922} /* (20, 28, 1) {real, imag} */,
  {32'hc022a435, 32'h3fa3dc1e} /* (20, 28, 0) {real, imag} */,
  {32'h3fc48926, 32'h4032e290} /* (20, 27, 31) {real, imag} */,
  {32'hc064e193, 32'h405a58ea} /* (20, 27, 30) {real, imag} */,
  {32'hbf16b030, 32'hc072983e} /* (20, 27, 29) {real, imag} */,
  {32'hbf267282, 32'h3f215094} /* (20, 27, 28) {real, imag} */,
  {32'hbfe149bf, 32'hbf6afc48} /* (20, 27, 27) {real, imag} */,
  {32'hc09c61dc, 32'h3eca85bd} /* (20, 27, 26) {real, imag} */,
  {32'h4039fb0c, 32'hbf08fa03} /* (20, 27, 25) {real, imag} */,
  {32'hbf8903ba, 32'hc01bd864} /* (20, 27, 24) {real, imag} */,
  {32'hbf6affcf, 32'hbf91e0c0} /* (20, 27, 23) {real, imag} */,
  {32'h3f1919eb, 32'h3e656db9} /* (20, 27, 22) {real, imag} */,
  {32'h401c046c, 32'h3f320a98} /* (20, 27, 21) {real, imag} */,
  {32'h4035c874, 32'hbff11c40} /* (20, 27, 20) {real, imag} */,
  {32'hbed16b71, 32'h400ec0b8} /* (20, 27, 19) {real, imag} */,
  {32'h3fb74b8c, 32'h3fd73a7e} /* (20, 27, 18) {real, imag} */,
  {32'hbff2867e, 32'h3ffad4ce} /* (20, 27, 17) {real, imag} */,
  {32'h3e5fbe59, 32'hbef76083} /* (20, 27, 16) {real, imag} */,
  {32'h401e10b9, 32'hbf900563} /* (20, 27, 15) {real, imag} */,
  {32'hbe5c12b3, 32'h40124dd9} /* (20, 27, 14) {real, imag} */,
  {32'h3e3c747e, 32'h3f6c55cc} /* (20, 27, 13) {real, imag} */,
  {32'hc073d7e6, 32'h3f28e908} /* (20, 27, 12) {real, imag} */,
  {32'hbfb5ebca, 32'h3fb16615} /* (20, 27, 11) {real, imag} */,
  {32'h3ff6409e, 32'hc0af30d0} /* (20, 27, 10) {real, imag} */,
  {32'hc0927f5b, 32'hbfec55e8} /* (20, 27, 9) {real, imag} */,
  {32'hbe93a6bd, 32'h403aa7ff} /* (20, 27, 8) {real, imag} */,
  {32'h3eed4340, 32'h401570ff} /* (20, 27, 7) {real, imag} */,
  {32'h4010b6bd, 32'hbfa15a67} /* (20, 27, 6) {real, imag} */,
  {32'hbfa2bf12, 32'h3f531cf2} /* (20, 27, 5) {real, imag} */,
  {32'h3f907caa, 32'hc00a0833} /* (20, 27, 4) {real, imag} */,
  {32'h3ed4a938, 32'hc06dc03d} /* (20, 27, 3) {real, imag} */,
  {32'h3fcc72ca, 32'hbeba528a} /* (20, 27, 2) {real, imag} */,
  {32'h40008b5a, 32'h4019bd99} /* (20, 27, 1) {real, imag} */,
  {32'hbf6d011d, 32'h3f8266de} /* (20, 27, 0) {real, imag} */,
  {32'hc0010780, 32'h3ffc2d41} /* (20, 26, 31) {real, imag} */,
  {32'h3fec6c83, 32'hbffc75d5} /* (20, 26, 30) {real, imag} */,
  {32'h3ede7837, 32'hbe944ad3} /* (20, 26, 29) {real, imag} */,
  {32'h3f14f106, 32'h3dc3c8dd} /* (20, 26, 28) {real, imag} */,
  {32'hc061b7e0, 32'h3f04e562} /* (20, 26, 27) {real, imag} */,
  {32'h4018619a, 32'h3f169bf2} /* (20, 26, 26) {real, imag} */,
  {32'hc01c909c, 32'hbf1ecd9f} /* (20, 26, 25) {real, imag} */,
  {32'h3f10724e, 32'hbf9bf8ad} /* (20, 26, 24) {real, imag} */,
  {32'h3f269043, 32'hbf7f986c} /* (20, 26, 23) {real, imag} */,
  {32'h3fafd7d7, 32'hbe514aa9} /* (20, 26, 22) {real, imag} */,
  {32'hc03a5a4b, 32'h3d119ab4} /* (20, 26, 21) {real, imag} */,
  {32'hbf2ec99c, 32'h3f6f0b45} /* (20, 26, 20) {real, imag} */,
  {32'h3f98e002, 32'hbe4a63ce} /* (20, 26, 19) {real, imag} */,
  {32'h3f22720e, 32'hc035c5a3} /* (20, 26, 18) {real, imag} */,
  {32'h3eea9c46, 32'h3e0c2d9e} /* (20, 26, 17) {real, imag} */,
  {32'hbf1cbb02, 32'hbf00fd46} /* (20, 26, 16) {real, imag} */,
  {32'hbfe15c8d, 32'hbe3809fb} /* (20, 26, 15) {real, imag} */,
  {32'h3f59feb2, 32'h3f93ffbf} /* (20, 26, 14) {real, imag} */,
  {32'h3f9361d1, 32'hc0003763} /* (20, 26, 13) {real, imag} */,
  {32'hbf6b37be, 32'h3fd968f5} /* (20, 26, 12) {real, imag} */,
  {32'h3f7becd5, 32'hbfd74261} /* (20, 26, 11) {real, imag} */,
  {32'h3fcf2a29, 32'hbe1f7fdb} /* (20, 26, 10) {real, imag} */,
  {32'h3f25dfda, 32'hbfcd5946} /* (20, 26, 9) {real, imag} */,
  {32'hc03cc10c, 32'h401825a2} /* (20, 26, 8) {real, imag} */,
  {32'h3d12ce04, 32'hbfe74235} /* (20, 26, 7) {real, imag} */,
  {32'h3fbfefe9, 32'h403593e1} /* (20, 26, 6) {real, imag} */,
  {32'h3f8340e3, 32'h3fd22f6d} /* (20, 26, 5) {real, imag} */,
  {32'hbf68e345, 32'h3f86f7f6} /* (20, 26, 4) {real, imag} */,
  {32'hc0092a5c, 32'h3eed1535} /* (20, 26, 3) {real, imag} */,
  {32'h3f68096a, 32'hbff84dca} /* (20, 26, 2) {real, imag} */,
  {32'h3fa1c29f, 32'h401d5b98} /* (20, 26, 1) {real, imag} */,
  {32'hbfddf40e, 32'hbff7b456} /* (20, 26, 0) {real, imag} */,
  {32'hc00d10f4, 32'hbffc5d0c} /* (20, 25, 31) {real, imag} */,
  {32'hc007d201, 32'hc0118c4a} /* (20, 25, 30) {real, imag} */,
  {32'h3fd56dd6, 32'h3ff3eaf3} /* (20, 25, 29) {real, imag} */,
  {32'h3ed77ac6, 32'h3fee76ff} /* (20, 25, 28) {real, imag} */,
  {32'h3f5ca7fa, 32'h3e4bb56e} /* (20, 25, 27) {real, imag} */,
  {32'hbfe3fccb, 32'hbf6ec713} /* (20, 25, 26) {real, imag} */,
  {32'hbf936138, 32'h3f9c0509} /* (20, 25, 25) {real, imag} */,
  {32'h401fbe62, 32'h3f194b0b} /* (20, 25, 24) {real, imag} */,
  {32'hbfbf57a3, 32'h3e3668f4} /* (20, 25, 23) {real, imag} */,
  {32'hbfc0db66, 32'hbf9d9670} /* (20, 25, 22) {real, imag} */,
  {32'hc02107df, 32'hbe9a164e} /* (20, 25, 21) {real, imag} */,
  {32'h4052830c, 32'hbf5d9140} /* (20, 25, 20) {real, imag} */,
  {32'hbe355215, 32'h3fea9572} /* (20, 25, 19) {real, imag} */,
  {32'h3fd3fa65, 32'h3fc83961} /* (20, 25, 18) {real, imag} */,
  {32'h3f9b4b43, 32'hbfc30ed3} /* (20, 25, 17) {real, imag} */,
  {32'h4005ed5a, 32'h403eef9a} /* (20, 25, 16) {real, imag} */,
  {32'hbf018ddd, 32'h3fbfa66d} /* (20, 25, 15) {real, imag} */,
  {32'hc06974c7, 32'h3ec64aaa} /* (20, 25, 14) {real, imag} */,
  {32'h3f621fed, 32'hbd09c997} /* (20, 25, 13) {real, imag} */,
  {32'hbf5a15f1, 32'hbfb91a42} /* (20, 25, 12) {real, imag} */,
  {32'h3f21ec92, 32'h4006cf7c} /* (20, 25, 11) {real, imag} */,
  {32'h3f2b94b6, 32'h3f9d819d} /* (20, 25, 10) {real, imag} */,
  {32'h40842474, 32'hbe298107} /* (20, 25, 9) {real, imag} */,
  {32'hbffa4101, 32'hc045bf51} /* (20, 25, 8) {real, imag} */,
  {32'hbfc3bca9, 32'h3ff76edc} /* (20, 25, 7) {real, imag} */,
  {32'hc0135c0f, 32'h3f3dbabe} /* (20, 25, 6) {real, imag} */,
  {32'h3fb0d042, 32'hc03a4232} /* (20, 25, 5) {real, imag} */,
  {32'h3f93fd5f, 32'hbfa44649} /* (20, 25, 4) {real, imag} */,
  {32'h3f263049, 32'h3fbb7dae} /* (20, 25, 3) {real, imag} */,
  {32'hbe1edd95, 32'h3f3bff19} /* (20, 25, 2) {real, imag} */,
  {32'h3fb6676d, 32'hbf76033b} /* (20, 25, 1) {real, imag} */,
  {32'h3fd8faaa, 32'h404fed1c} /* (20, 25, 0) {real, imag} */,
  {32'h3e12cb44, 32'h3f1c58c9} /* (20, 24, 31) {real, imag} */,
  {32'h405db04f, 32'h400e60a2} /* (20, 24, 30) {real, imag} */,
  {32'h4035c874, 32'hbfa39a89} /* (20, 24, 29) {real, imag} */,
  {32'h402a4d3b, 32'h3f8b125e} /* (20, 24, 28) {real, imag} */,
  {32'h3f378914, 32'hbfb4bb25} /* (20, 24, 27) {real, imag} */,
  {32'h40069077, 32'hbe7774dc} /* (20, 24, 26) {real, imag} */,
  {32'h400e24ab, 32'hbf7ab8ac} /* (20, 24, 25) {real, imag} */,
  {32'hbecd896e, 32'hbfb52feb} /* (20, 24, 24) {real, imag} */,
  {32'hc02c5c66, 32'h3f9b4ec9} /* (20, 24, 23) {real, imag} */,
  {32'hbfa75b11, 32'h3f11d415} /* (20, 24, 22) {real, imag} */,
  {32'h3f234298, 32'hbdd98936} /* (20, 24, 21) {real, imag} */,
  {32'h40266fad, 32'h3f7cda85} /* (20, 24, 20) {real, imag} */,
  {32'h3fadd750, 32'h3f33c075} /* (20, 24, 19) {real, imag} */,
  {32'hbf9d6d81, 32'hc0114813} /* (20, 24, 18) {real, imag} */,
  {32'hbeb8073d, 32'hbfa83e56} /* (20, 24, 17) {real, imag} */,
  {32'hbf4aeadb, 32'hc011d567} /* (20, 24, 16) {real, imag} */,
  {32'h3f6ec3b8, 32'hbf83b9f4} /* (20, 24, 15) {real, imag} */,
  {32'h3f1ee021, 32'h3f0a6607} /* (20, 24, 14) {real, imag} */,
  {32'hbf7b35fe, 32'h3ecc875c} /* (20, 24, 13) {real, imag} */,
  {32'h3e722b6e, 32'hbdf55a55} /* (20, 24, 12) {real, imag} */,
  {32'h3e104349, 32'hbdfabeb7} /* (20, 24, 11) {real, imag} */,
  {32'hbff9a9d2, 32'h3ef48c00} /* (20, 24, 10) {real, imag} */,
  {32'h3dc3e983, 32'hbf937a11} /* (20, 24, 9) {real, imag} */,
  {32'hbef13d6f, 32'hc0244269} /* (20, 24, 8) {real, imag} */,
  {32'h3faacda1, 32'h3ec7b355} /* (20, 24, 7) {real, imag} */,
  {32'h3ee98aff, 32'hbfe825bc} /* (20, 24, 6) {real, imag} */,
  {32'hc00a6fef, 32'hbe8643ab} /* (20, 24, 5) {real, imag} */,
  {32'h3faa8367, 32'hbf588590} /* (20, 24, 4) {real, imag} */,
  {32'hbf8e2801, 32'hbf7db5c9} /* (20, 24, 3) {real, imag} */,
  {32'hbff070a9, 32'h4004c3b4} /* (20, 24, 2) {real, imag} */,
  {32'hbf5a1dda, 32'hbfeade83} /* (20, 24, 1) {real, imag} */,
  {32'h3f034000, 32'h3d8ec137} /* (20, 24, 0) {real, imag} */,
  {32'hc0708f0d, 32'h3fd19d44} /* (20, 23, 31) {real, imag} */,
  {32'hbf0a5037, 32'h3ee44d2c} /* (20, 23, 30) {real, imag} */,
  {32'hbfab0b3d, 32'h404e546a} /* (20, 23, 29) {real, imag} */,
  {32'hbfd0767e, 32'hbf80ef85} /* (20, 23, 28) {real, imag} */,
  {32'h405839de, 32'h3fd6a5bf} /* (20, 23, 27) {real, imag} */,
  {32'h3fdb3324, 32'h3f160293} /* (20, 23, 26) {real, imag} */,
  {32'hbfc6fdba, 32'h3ec6e3ed} /* (20, 23, 25) {real, imag} */,
  {32'hbfba0627, 32'h3e93b85f} /* (20, 23, 24) {real, imag} */,
  {32'hbfb0e3b9, 32'h3f7a8c1f} /* (20, 23, 23) {real, imag} */,
  {32'hc01986bb, 32'hbfd3bf31} /* (20, 23, 22) {real, imag} */,
  {32'h3f5d7720, 32'hc0603f07} /* (20, 23, 21) {real, imag} */,
  {32'hbfbb50c9, 32'h3f1f9274} /* (20, 23, 20) {real, imag} */,
  {32'hc017dfbd, 32'hbfbb1acc} /* (20, 23, 19) {real, imag} */,
  {32'hbf9ab209, 32'hc0488f7a} /* (20, 23, 18) {real, imag} */,
  {32'hbf906f97, 32'hbf1ecf79} /* (20, 23, 17) {real, imag} */,
  {32'h3ec67b46, 32'hbf57eb2c} /* (20, 23, 16) {real, imag} */,
  {32'h3e346baf, 32'h3ff90358} /* (20, 23, 15) {real, imag} */,
  {32'h3e9a4dcf, 32'h3f01acf4} /* (20, 23, 14) {real, imag} */,
  {32'h40367ecd, 32'h3f8e503e} /* (20, 23, 13) {real, imag} */,
  {32'hbf31ad54, 32'h3fbeaac0} /* (20, 23, 12) {real, imag} */,
  {32'hbe37c96d, 32'h3ea351d0} /* (20, 23, 11) {real, imag} */,
  {32'hbef2cef3, 32'h3edd8b62} /* (20, 23, 10) {real, imag} */,
  {32'hc0850b75, 32'hc001dd52} /* (20, 23, 9) {real, imag} */,
  {32'h3facef0c, 32'hbf524124} /* (20, 23, 8) {real, imag} */,
  {32'hbf1e55b5, 32'h403f2222} /* (20, 23, 7) {real, imag} */,
  {32'hbe459573, 32'hbdf7a872} /* (20, 23, 6) {real, imag} */,
  {32'hbe1e6095, 32'hbf8c3d84} /* (20, 23, 5) {real, imag} */,
  {32'h3de961e0, 32'hbf5bcbb7} /* (20, 23, 4) {real, imag} */,
  {32'h3f5439a7, 32'hbfb7285f} /* (20, 23, 3) {real, imag} */,
  {32'h3e00e999, 32'hc08e209e} /* (20, 23, 2) {real, imag} */,
  {32'hbfb67aef, 32'hbf9490d7} /* (20, 23, 1) {real, imag} */,
  {32'h3ef3b4b2, 32'h3fdbebc3} /* (20, 23, 0) {real, imag} */,
  {32'hbfa54dcd, 32'h401de49d} /* (20, 22, 31) {real, imag} */,
  {32'h3fc092fb, 32'hbf74c236} /* (20, 22, 30) {real, imag} */,
  {32'hc03b388c, 32'h3f9115ef} /* (20, 22, 29) {real, imag} */,
  {32'h401ab7ad, 32'h3f40ed81} /* (20, 22, 28) {real, imag} */,
  {32'hbfc4dbe6, 32'hbfc01e74} /* (20, 22, 27) {real, imag} */,
  {32'hc081171b, 32'h3f541278} /* (20, 22, 26) {real, imag} */,
  {32'hbf7ac57b, 32'h3fa73ee8} /* (20, 22, 25) {real, imag} */,
  {32'hbe83165e, 32'h3f8e2eee} /* (20, 22, 24) {real, imag} */,
  {32'hc0153672, 32'h3e2850a5} /* (20, 22, 23) {real, imag} */,
  {32'hbedf6e4c, 32'hbf226fd3} /* (20, 22, 22) {real, imag} */,
  {32'hbf272fa6, 32'h3d36a3b2} /* (20, 22, 21) {real, imag} */,
  {32'hc01f32d1, 32'hc0538daa} /* (20, 22, 20) {real, imag} */,
  {32'hbfafe83f, 32'hbd4598f5} /* (20, 22, 19) {real, imag} */,
  {32'h40a7542e, 32'h3fb605a4} /* (20, 22, 18) {real, imag} */,
  {32'h4049b8b8, 32'hc04fe67b} /* (20, 22, 17) {real, imag} */,
  {32'hbfb0d33f, 32'hbe37b6e0} /* (20, 22, 16) {real, imag} */,
  {32'hbedd057b, 32'h3baf5c9b} /* (20, 22, 15) {real, imag} */,
  {32'hc0244066, 32'h3fd542b2} /* (20, 22, 14) {real, imag} */,
  {32'h400eed35, 32'hbfc53f1e} /* (20, 22, 13) {real, imag} */,
  {32'h3f308b5f, 32'h3f611dd4} /* (20, 22, 12) {real, imag} */,
  {32'h3fd026b8, 32'hbdcd44bf} /* (20, 22, 11) {real, imag} */,
  {32'h3f7a0a57, 32'h3e6f257e} /* (20, 22, 10) {real, imag} */,
  {32'h3e7f4eb1, 32'h3fce8f31} /* (20, 22, 9) {real, imag} */,
  {32'hbfab611f, 32'h40086432} /* (20, 22, 8) {real, imag} */,
  {32'h3e583a26, 32'h3f70fa4b} /* (20, 22, 7) {real, imag} */,
  {32'hc014f1cb, 32'h3e6b2ecf} /* (20, 22, 6) {real, imag} */,
  {32'hbf330825, 32'hc07a452f} /* (20, 22, 5) {real, imag} */,
  {32'h3f16ee62, 32'h3ef316a6} /* (20, 22, 4) {real, imag} */,
  {32'hbebd3cf4, 32'h3f99591a} /* (20, 22, 3) {real, imag} */,
  {32'hbedecf38, 32'hbf559ddd} /* (20, 22, 2) {real, imag} */,
  {32'hc00214f3, 32'hbec91c52} /* (20, 22, 1) {real, imag} */,
  {32'hbf314444, 32'h3f172a66} /* (20, 22, 0) {real, imag} */,
  {32'hbe5ba1c6, 32'h3f38645d} /* (20, 21, 31) {real, imag} */,
  {32'h401a659c, 32'hbfc4d913} /* (20, 21, 30) {real, imag} */,
  {32'h403a6a17, 32'hbfcb26af} /* (20, 21, 29) {real, imag} */,
  {32'h3e1259b6, 32'h3f69a7b1} /* (20, 21, 28) {real, imag} */,
  {32'h3ef71dde, 32'hbf91d6db} /* (20, 21, 27) {real, imag} */,
  {32'hc067109f, 32'hbdf94e45} /* (20, 21, 26) {real, imag} */,
  {32'hc0040cf5, 32'hbfd63479} /* (20, 21, 25) {real, imag} */,
  {32'h4020d5c3, 32'hbfba3023} /* (20, 21, 24) {real, imag} */,
  {32'h4095d4ae, 32'hc0866ad3} /* (20, 21, 23) {real, imag} */,
  {32'hc03af8fb, 32'h3f3b3951} /* (20, 21, 22) {real, imag} */,
  {32'h3f2283c0, 32'hbf947792} /* (20, 21, 21) {real, imag} */,
  {32'h402d8c4f, 32'h3f272085} /* (20, 21, 20) {real, imag} */,
  {32'hbfc4bf51, 32'h3e894e1f} /* (20, 21, 19) {real, imag} */,
  {32'h3fb5b406, 32'hbfcb0163} /* (20, 21, 18) {real, imag} */,
  {32'hbf70ac81, 32'h400daaa9} /* (20, 21, 17) {real, imag} */,
  {32'h3e941d7c, 32'hbfc02c9e} /* (20, 21, 16) {real, imag} */,
  {32'hbe4d47fc, 32'h3f839b31} /* (20, 21, 15) {real, imag} */,
  {32'h3fddada8, 32'h3eed6f10} /* (20, 21, 14) {real, imag} */,
  {32'hbe81fc22, 32'hc05efddf} /* (20, 21, 13) {real, imag} */,
  {32'h4070927a, 32'hc0394cbf} /* (20, 21, 12) {real, imag} */,
  {32'h400fce49, 32'h400c240c} /* (20, 21, 11) {real, imag} */,
  {32'h4046791b, 32'hbf923cc3} /* (20, 21, 10) {real, imag} */,
  {32'hbf81d346, 32'hbef56ef7} /* (20, 21, 9) {real, imag} */,
  {32'h3f126521, 32'h401a5a9f} /* (20, 21, 8) {real, imag} */,
  {32'h408108bf, 32'h3ea2bf5f} /* (20, 21, 7) {real, imag} */,
  {32'h3f784c89, 32'h3e315bfa} /* (20, 21, 6) {real, imag} */,
  {32'h3f094f89, 32'hbfcbc111} /* (20, 21, 5) {real, imag} */,
  {32'hbfef6cea, 32'hbf023bce} /* (20, 21, 4) {real, imag} */,
  {32'h3fd68f45, 32'h3f7790a9} /* (20, 21, 3) {real, imag} */,
  {32'hc02a587e, 32'h3f99edf4} /* (20, 21, 2) {real, imag} */,
  {32'h3f09371e, 32'h400a3a31} /* (20, 21, 1) {real, imag} */,
  {32'hbf0ae548, 32'h4032bcf6} /* (20, 21, 0) {real, imag} */,
  {32'hbf373c8c, 32'h3f6b6c7b} /* (20, 20, 31) {real, imag} */,
  {32'hbec8c877, 32'h3fe1330d} /* (20, 20, 30) {real, imag} */,
  {32'h4041e546, 32'hc01919cf} /* (20, 20, 29) {real, imag} */,
  {32'hbf35fc58, 32'h3e98941d} /* (20, 20, 28) {real, imag} */,
  {32'h40060571, 32'h3fa338aa} /* (20, 20, 27) {real, imag} */,
  {32'hbec050b8, 32'h40769b75} /* (20, 20, 26) {real, imag} */,
  {32'hbee031be, 32'hbf0534c1} /* (20, 20, 25) {real, imag} */,
  {32'hbf74fbef, 32'hbe54f0e2} /* (20, 20, 24) {real, imag} */,
  {32'h409d855e, 32'h403a521b} /* (20, 20, 23) {real, imag} */,
  {32'hc00f083d, 32'hc05bc8eb} /* (20, 20, 22) {real, imag} */,
  {32'hbdc39445, 32'h3ff18ca1} /* (20, 20, 21) {real, imag} */,
  {32'hc06ea7c4, 32'h3fc5f4f4} /* (20, 20, 20) {real, imag} */,
  {32'hc01ce977, 32'h3e1a3e83} /* (20, 20, 19) {real, imag} */,
  {32'hc0019e27, 32'h400c02c3} /* (20, 20, 18) {real, imag} */,
  {32'h3fa55409, 32'h3faa9d65} /* (20, 20, 17) {real, imag} */,
  {32'h401cbca5, 32'hbf921c15} /* (20, 20, 16) {real, imag} */,
  {32'hbfbe876d, 32'h3e49bcef} /* (20, 20, 15) {real, imag} */,
  {32'hc030fa65, 32'hbf172d66} /* (20, 20, 14) {real, imag} */,
  {32'hbfbaf1f2, 32'h40077ac1} /* (20, 20, 13) {real, imag} */,
  {32'h3eb11e9f, 32'hbfe56224} /* (20, 20, 12) {real, imag} */,
  {32'h3cb41ef0, 32'hbcf222ea} /* (20, 20, 11) {real, imag} */,
  {32'h3fb10c91, 32'h3fffb21b} /* (20, 20, 10) {real, imag} */,
  {32'hbfc4ea4f, 32'h3fdf2169} /* (20, 20, 9) {real, imag} */,
  {32'h3f4c6b67, 32'h3fc53b3e} /* (20, 20, 8) {real, imag} */,
  {32'hbeaab354, 32'h3fefa64f} /* (20, 20, 7) {real, imag} */,
  {32'h3f0197a2, 32'h3fd411f5} /* (20, 20, 6) {real, imag} */,
  {32'hbf1adf75, 32'h3f915cad} /* (20, 20, 5) {real, imag} */,
  {32'hc00cb56f, 32'hbf4ee717} /* (20, 20, 4) {real, imag} */,
  {32'h4004ecaa, 32'hc0055d11} /* (20, 20, 3) {real, imag} */,
  {32'h3e80b3c2, 32'h3f70fa74} /* (20, 20, 2) {real, imag} */,
  {32'hbf9cf633, 32'hc0063484} /* (20, 20, 1) {real, imag} */,
  {32'h40295a6f, 32'hc08729c3} /* (20, 20, 0) {real, imag} */,
  {32'hbf95fe39, 32'hc00f57db} /* (20, 19, 31) {real, imag} */,
  {32'hbee45358, 32'h3f1221ba} /* (20, 19, 30) {real, imag} */,
  {32'h3e945014, 32'h3ffaf401} /* (20, 19, 29) {real, imag} */,
  {32'hbfa00a1c, 32'h40441b7e} /* (20, 19, 28) {real, imag} */,
  {32'h4096f567, 32'h3f16e7b9} /* (20, 19, 27) {real, imag} */,
  {32'h3e88a4f6, 32'hbea70d50} /* (20, 19, 26) {real, imag} */,
  {32'h3fb49727, 32'h3f818ab4} /* (20, 19, 25) {real, imag} */,
  {32'h4008858a, 32'h3d892e22} /* (20, 19, 24) {real, imag} */,
  {32'h401e23ca, 32'hbe2abb57} /* (20, 19, 23) {real, imag} */,
  {32'h3f23eedb, 32'h3fd4214c} /* (20, 19, 22) {real, imag} */,
  {32'h40252f6f, 32'hc0061470} /* (20, 19, 21) {real, imag} */,
  {32'hbe848ae0, 32'h3fe0170e} /* (20, 19, 20) {real, imag} */,
  {32'hbe76b5e8, 32'hbec06895} /* (20, 19, 19) {real, imag} */,
  {32'hbf771f1f, 32'h3eb87b44} /* (20, 19, 18) {real, imag} */,
  {32'hbf9421d9, 32'hbf974416} /* (20, 19, 17) {real, imag} */,
  {32'hc02a11ba, 32'hbf0a21d0} /* (20, 19, 16) {real, imag} */,
  {32'hbf89d200, 32'h3fae348d} /* (20, 19, 15) {real, imag} */,
  {32'hc01f549f, 32'hc01827df} /* (20, 19, 14) {real, imag} */,
  {32'hbfdf40fa, 32'hbf7903a5} /* (20, 19, 13) {real, imag} */,
  {32'hbebf6773, 32'hc046b167} /* (20, 19, 12) {real, imag} */,
  {32'h406d3527, 32'hbe810a5f} /* (20, 19, 11) {real, imag} */,
  {32'h3e64195b, 32'hbebcb788} /* (20, 19, 10) {real, imag} */,
  {32'h3faf5f47, 32'h3f628b0f} /* (20, 19, 9) {real, imag} */,
  {32'h3fc686c5, 32'hbd9753e2} /* (20, 19, 8) {real, imag} */,
  {32'h3e7d3b45, 32'hbeee89c6} /* (20, 19, 7) {real, imag} */,
  {32'hbf9715b7, 32'hc0444c45} /* (20, 19, 6) {real, imag} */,
  {32'hc0160970, 32'hc033612d} /* (20, 19, 5) {real, imag} */,
  {32'hbf41d0e6, 32'h3e25b63d} /* (20, 19, 4) {real, imag} */,
  {32'hc03e3e7d, 32'hc0428389} /* (20, 19, 3) {real, imag} */,
  {32'h3fd72be4, 32'hbf515754} /* (20, 19, 2) {real, imag} */,
  {32'hc02c0579, 32'h3f25da9e} /* (20, 19, 1) {real, imag} */,
  {32'h400cec7f, 32'hbe503136} /* (20, 19, 0) {real, imag} */,
  {32'h3eca8ee3, 32'h3e8b0c63} /* (20, 18, 31) {real, imag} */,
  {32'h3faa6259, 32'h3f7c4ec0} /* (20, 18, 30) {real, imag} */,
  {32'hbfbaf525, 32'h3dada517} /* (20, 18, 29) {real, imag} */,
  {32'hc01d59f0, 32'hbfe76d2b} /* (20, 18, 28) {real, imag} */,
  {32'hbf973665, 32'h40934b76} /* (20, 18, 27) {real, imag} */,
  {32'hbf87da4f, 32'h4002a569} /* (20, 18, 26) {real, imag} */,
  {32'hc0826b3d, 32'h3de5b106} /* (20, 18, 25) {real, imag} */,
  {32'h3f5f3b1c, 32'hbdfd3135} /* (20, 18, 24) {real, imag} */,
  {32'hc02a1c2b, 32'hbfb91066} /* (20, 18, 23) {real, imag} */,
  {32'hbf81819c, 32'hbf8fa31e} /* (20, 18, 22) {real, imag} */,
  {32'h3fb8e01a, 32'hbf97ef20} /* (20, 18, 21) {real, imag} */,
  {32'h3e728038, 32'hbf960282} /* (20, 18, 20) {real, imag} */,
  {32'h3fe9b6b2, 32'hbfebe771} /* (20, 18, 19) {real, imag} */,
  {32'h3fd90387, 32'h406eb69a} /* (20, 18, 18) {real, imag} */,
  {32'h4091ce37, 32'h4041802a} /* (20, 18, 17) {real, imag} */,
  {32'hbf119345, 32'h40116ef4} /* (20, 18, 16) {real, imag} */,
  {32'hbf307fc3, 32'hbf5a5ff6} /* (20, 18, 15) {real, imag} */,
  {32'h3e83a305, 32'hbe384be8} /* (20, 18, 14) {real, imag} */,
  {32'h4014d0bb, 32'h40007a47} /* (20, 18, 13) {real, imag} */,
  {32'h40267253, 32'h3f83e160} /* (20, 18, 12) {real, imag} */,
  {32'h4059893c, 32'h3fef379b} /* (20, 18, 11) {real, imag} */,
  {32'hc0821b83, 32'hbe161651} /* (20, 18, 10) {real, imag} */,
  {32'hc01ad171, 32'hbf7d4db5} /* (20, 18, 9) {real, imag} */,
  {32'hbe3d98f6, 32'hbf46d18f} /* (20, 18, 8) {real, imag} */,
  {32'hbfa17348, 32'hbebaa10f} /* (20, 18, 7) {real, imag} */,
  {32'hc03fef6a, 32'hbf99230d} /* (20, 18, 6) {real, imag} */,
  {32'h3dbaa385, 32'h3ffc648a} /* (20, 18, 5) {real, imag} */,
  {32'h404845f9, 32'h3d5ba71e} /* (20, 18, 4) {real, imag} */,
  {32'h3e9d1181, 32'hbe8afa69} /* (20, 18, 3) {real, imag} */,
  {32'hbfbf4465, 32'hbfc080c5} /* (20, 18, 2) {real, imag} */,
  {32'hbfcaa632, 32'h3f863b1a} /* (20, 18, 1) {real, imag} */,
  {32'hbe86f147, 32'hbf8e6d70} /* (20, 18, 0) {real, imag} */,
  {32'h3e8fb452, 32'hbf54503a} /* (20, 17, 31) {real, imag} */,
  {32'h3de3f83b, 32'hbe945530} /* (20, 17, 30) {real, imag} */,
  {32'hbf429e0a, 32'hbd813a4b} /* (20, 17, 29) {real, imag} */,
  {32'hbff63321, 32'h400ba828} /* (20, 17, 28) {real, imag} */,
  {32'hbf7dabd1, 32'hbfc179bb} /* (20, 17, 27) {real, imag} */,
  {32'h3e9845de, 32'h404c058e} /* (20, 17, 26) {real, imag} */,
  {32'h3e96f053, 32'hbfb53dbd} /* (20, 17, 25) {real, imag} */,
  {32'h3f1bfad5, 32'h401d043f} /* (20, 17, 24) {real, imag} */,
  {32'hbe22222d, 32'hbf15f434} /* (20, 17, 23) {real, imag} */,
  {32'hc01e0c5c, 32'h3e727fde} /* (20, 17, 22) {real, imag} */,
  {32'h3f130728, 32'hc00dac11} /* (20, 17, 21) {real, imag} */,
  {32'h3f5f9209, 32'h4074ee95} /* (20, 17, 20) {real, imag} */,
  {32'h40229a95, 32'h3fe83aca} /* (20, 17, 19) {real, imag} */,
  {32'hbf1767a6, 32'hbeb7ab6e} /* (20, 17, 18) {real, imag} */,
  {32'hbf048156, 32'h3fa07be2} /* (20, 17, 17) {real, imag} */,
  {32'hbe56fdb3, 32'hbf526464} /* (20, 17, 16) {real, imag} */,
  {32'h3fe08baa, 32'hc0379828} /* (20, 17, 15) {real, imag} */,
  {32'h3f8f7b45, 32'h3f5ecf11} /* (20, 17, 14) {real, imag} */,
  {32'h3ed0b70f, 32'hbea1700d} /* (20, 17, 13) {real, imag} */,
  {32'hc0b07864, 32'hbee245ee} /* (20, 17, 12) {real, imag} */,
  {32'hbfdd7160, 32'hbf8c6fee} /* (20, 17, 11) {real, imag} */,
  {32'h3dd5e219, 32'h3f449978} /* (20, 17, 10) {real, imag} */,
  {32'h407dc0f5, 32'h3e4a5996} /* (20, 17, 9) {real, imag} */,
  {32'h401950fc, 32'hbf74ed77} /* (20, 17, 8) {real, imag} */,
  {32'hbf59509b, 32'hbf9b4496} /* (20, 17, 7) {real, imag} */,
  {32'hbf27d347, 32'hbfde5093} /* (20, 17, 6) {real, imag} */,
  {32'hbf54a706, 32'hbed843fe} /* (20, 17, 5) {real, imag} */,
  {32'h3f67a170, 32'hbeb16c01} /* (20, 17, 4) {real, imag} */,
  {32'h3fb908cc, 32'h3ea86160} /* (20, 17, 3) {real, imag} */,
  {32'h3f4e47c1, 32'hbf807a16} /* (20, 17, 2) {real, imag} */,
  {32'h3f82bc03, 32'h3f2e4b04} /* (20, 17, 1) {real, imag} */,
  {32'h3fe05b1b, 32'hbd1a311e} /* (20, 17, 0) {real, imag} */,
  {32'h3f2529cf, 32'h3d00e017} /* (20, 16, 31) {real, imag} */,
  {32'hbe8b5bee, 32'hbf3dd707} /* (20, 16, 30) {real, imag} */,
  {32'hbfdd63c1, 32'h3ea39bad} /* (20, 16, 29) {real, imag} */,
  {32'hbce569f3, 32'hbf94e02c} /* (20, 16, 28) {real, imag} */,
  {32'h3c3080e3, 32'hbf681d90} /* (20, 16, 27) {real, imag} */,
  {32'hc00ebe0b, 32'h3fb71fcf} /* (20, 16, 26) {real, imag} */,
  {32'h3ea90121, 32'h3fe0c467} /* (20, 16, 25) {real, imag} */,
  {32'hbe514099, 32'h3feaf68d} /* (20, 16, 24) {real, imag} */,
  {32'h3fc23be7, 32'hbff3cfe6} /* (20, 16, 23) {real, imag} */,
  {32'hbf8238a3, 32'hbed6269f} /* (20, 16, 22) {real, imag} */,
  {32'h3e3ef911, 32'hbc910b05} /* (20, 16, 21) {real, imag} */,
  {32'hbfef3e28, 32'h3f1cde93} /* (20, 16, 20) {real, imag} */,
  {32'hc02bdce6, 32'hc0042b6c} /* (20, 16, 19) {real, imag} */,
  {32'hbfc52942, 32'hbf3aa457} /* (20, 16, 18) {real, imag} */,
  {32'hbfe3a9ad, 32'hc0095252} /* (20, 16, 17) {real, imag} */,
  {32'hbfc1df6b, 32'hbe4c9cc8} /* (20, 16, 16) {real, imag} */,
  {32'h3f8111e2, 32'hbfef683a} /* (20, 16, 15) {real, imag} */,
  {32'h3f51f7f0, 32'h3f4c1a65} /* (20, 16, 14) {real, imag} */,
  {32'hc03fa6da, 32'hc0209f0e} /* (20, 16, 13) {real, imag} */,
  {32'h40323e11, 32'h3d9dbb6e} /* (20, 16, 12) {real, imag} */,
  {32'h402bbc3a, 32'h3f5edddb} /* (20, 16, 11) {real, imag} */,
  {32'hbe502012, 32'h3fafdf01} /* (20, 16, 10) {real, imag} */,
  {32'h3f830de3, 32'hbec1d4e7} /* (20, 16, 9) {real, imag} */,
  {32'hbfe8aa4f, 32'h3f807358} /* (20, 16, 8) {real, imag} */,
  {32'h3f090236, 32'hbf65c0c7} /* (20, 16, 7) {real, imag} */,
  {32'hbf1618e0, 32'h3f7c7489} /* (20, 16, 6) {real, imag} */,
  {32'h3e43e027, 32'hc005f5d8} /* (20, 16, 5) {real, imag} */,
  {32'hc0045fd3, 32'h3f52b3ed} /* (20, 16, 4) {real, imag} */,
  {32'hbf8c45bb, 32'hbfa365ac} /* (20, 16, 3) {real, imag} */,
  {32'h3ff2a6f4, 32'hc01452a9} /* (20, 16, 2) {real, imag} */,
  {32'h3f2bd5ba, 32'h3fc505db} /* (20, 16, 1) {real, imag} */,
  {32'h3f0abea4, 32'h3e3f69e3} /* (20, 16, 0) {real, imag} */,
  {32'hbf265b59, 32'h403d077e} /* (20, 15, 31) {real, imag} */,
  {32'h3f0b78c5, 32'hbf09d159} /* (20, 15, 30) {real, imag} */,
  {32'h3f8cb042, 32'h3f711a82} /* (20, 15, 29) {real, imag} */,
  {32'hbed1794e, 32'hbc51137b} /* (20, 15, 28) {real, imag} */,
  {32'hbfb00ee9, 32'hc0098dda} /* (20, 15, 27) {real, imag} */,
  {32'h409965a7, 32'h3f82d5bf} /* (20, 15, 26) {real, imag} */,
  {32'h4014e15a, 32'h3f0d8a31} /* (20, 15, 25) {real, imag} */,
  {32'h3c9a6d5a, 32'h4058a489} /* (20, 15, 24) {real, imag} */,
  {32'hbf99d544, 32'hc014febb} /* (20, 15, 23) {real, imag} */,
  {32'hbf7e69a2, 32'hbf48d81c} /* (20, 15, 22) {real, imag} */,
  {32'hbf289f01, 32'hbf27fb2e} /* (20, 15, 21) {real, imag} */,
  {32'hbe450c16, 32'hbf4e608e} /* (20, 15, 20) {real, imag} */,
  {32'hbf6fe58c, 32'hbfa705cb} /* (20, 15, 19) {real, imag} */,
  {32'h403dc201, 32'hbfa53030} /* (20, 15, 18) {real, imag} */,
  {32'h3fc38680, 32'h3f68160a} /* (20, 15, 17) {real, imag} */,
  {32'hbe3398f9, 32'hbd9fdcd7} /* (20, 15, 16) {real, imag} */,
  {32'hbe25b574, 32'h3eb8c881} /* (20, 15, 15) {real, imag} */,
  {32'hbf04ba9e, 32'hbf2af483} /* (20, 15, 14) {real, imag} */,
  {32'h3f84a4b7, 32'hbedafa6e} /* (20, 15, 13) {real, imag} */,
  {32'h3fa42bd7, 32'hbf864ae4} /* (20, 15, 12) {real, imag} */,
  {32'h3f4b36d3, 32'h3f93a560} /* (20, 15, 11) {real, imag} */,
  {32'h4017b767, 32'hc02d21dd} /* (20, 15, 10) {real, imag} */,
  {32'hc04ac0f5, 32'h400c18c4} /* (20, 15, 9) {real, imag} */,
  {32'hbf0e07ca, 32'hbf27c2f8} /* (20, 15, 8) {real, imag} */,
  {32'hbfd2625e, 32'h400e196c} /* (20, 15, 7) {real, imag} */,
  {32'h3e2e31c5, 32'hc0508e94} /* (20, 15, 6) {real, imag} */,
  {32'h3f1076bc, 32'hbf1ad45c} /* (20, 15, 5) {real, imag} */,
  {32'h3fba5641, 32'hc0371b7d} /* (20, 15, 4) {real, imag} */,
  {32'hbf922855, 32'h3e21dc96} /* (20, 15, 3) {real, imag} */,
  {32'h40102cde, 32'h3f0abc52} /* (20, 15, 2) {real, imag} */,
  {32'hbdd82d2e, 32'h3ea95ddf} /* (20, 15, 1) {real, imag} */,
  {32'hbe98e0ce, 32'h3fdfebaf} /* (20, 15, 0) {real, imag} */,
  {32'h4001f8cb, 32'h3e1995f4} /* (20, 14, 31) {real, imag} */,
  {32'hbf68a7ac, 32'hc03768e5} /* (20, 14, 30) {real, imag} */,
  {32'hbf631cfa, 32'hbf24b9b6} /* (20, 14, 29) {real, imag} */,
  {32'h3de36833, 32'h3fe38b7b} /* (20, 14, 28) {real, imag} */,
  {32'h3f852203, 32'hbf906fe2} /* (20, 14, 27) {real, imag} */,
  {32'hbeda4206, 32'h406ca04a} /* (20, 14, 26) {real, imag} */,
  {32'h3f9b2fe5, 32'hbf1f8e88} /* (20, 14, 25) {real, imag} */,
  {32'hbf12ee71, 32'h3fa09f3a} /* (20, 14, 24) {real, imag} */,
  {32'h405e2676, 32'h3f481baf} /* (20, 14, 23) {real, imag} */,
  {32'h403f7356, 32'hc05c7be4} /* (20, 14, 22) {real, imag} */,
  {32'hc0157be1, 32'h3fd08331} /* (20, 14, 21) {real, imag} */,
  {32'hc042034d, 32'hbefd7aff} /* (20, 14, 20) {real, imag} */,
  {32'h4028c5f0, 32'hc041dd30} /* (20, 14, 19) {real, imag} */,
  {32'hbf54f018, 32'h408ab0d7} /* (20, 14, 18) {real, imag} */,
  {32'hc048af3c, 32'h3f760916} /* (20, 14, 17) {real, imag} */,
  {32'hc0281794, 32'h3f009579} /* (20, 14, 16) {real, imag} */,
  {32'hbe0c09eb, 32'h3fac2e4c} /* (20, 14, 15) {real, imag} */,
  {32'hbfd45b3d, 32'h4087fbd8} /* (20, 14, 14) {real, imag} */,
  {32'h3f1c9412, 32'hc003dbec} /* (20, 14, 13) {real, imag} */,
  {32'hbfedbbff, 32'h3e94e180} /* (20, 14, 12) {real, imag} */,
  {32'h3ffa9d8f, 32'hbffb2d37} /* (20, 14, 11) {real, imag} */,
  {32'hc06136d6, 32'h402912dd} /* (20, 14, 10) {real, imag} */,
  {32'h3f1ea82c, 32'hc0192d24} /* (20, 14, 9) {real, imag} */,
  {32'hbe4e8f41, 32'h3f01555d} /* (20, 14, 8) {real, imag} */,
  {32'h3f6be1d4, 32'h3eb706c8} /* (20, 14, 7) {real, imag} */,
  {32'h3d60cd61, 32'hbe993f72} /* (20, 14, 6) {real, imag} */,
  {32'hbf4c9cc6, 32'hbfd6fffa} /* (20, 14, 5) {real, imag} */,
  {32'h3f804535, 32'h3f8bec81} /* (20, 14, 4) {real, imag} */,
  {32'h403ffe8b, 32'h3f8e1c9d} /* (20, 14, 3) {real, imag} */,
  {32'hbfb1008c, 32'h3c21e5d3} /* (20, 14, 2) {real, imag} */,
  {32'h3f22f672, 32'hbf6c16c9} /* (20, 14, 1) {real, imag} */,
  {32'h3f8d035b, 32'hbfeccbf7} /* (20, 14, 0) {real, imag} */,
  {32'h3faf2de7, 32'hc0008c9c} /* (20, 13, 31) {real, imag} */,
  {32'h40225349, 32'hbfcc53ec} /* (20, 13, 30) {real, imag} */,
  {32'hbd0bc284, 32'h3ff87f30} /* (20, 13, 29) {real, imag} */,
  {32'h3efb1933, 32'h3eb9e83f} /* (20, 13, 28) {real, imag} */,
  {32'hbf8829ee, 32'h3fc38690} /* (20, 13, 27) {real, imag} */,
  {32'hc009e29c, 32'h403b30f5} /* (20, 13, 26) {real, imag} */,
  {32'hbebb1cdc, 32'h3eb51690} /* (20, 13, 25) {real, imag} */,
  {32'hc01fd145, 32'hc0555d0c} /* (20, 13, 24) {real, imag} */,
  {32'hbf90f216, 32'hbe3a9aa3} /* (20, 13, 23) {real, imag} */,
  {32'hbd86df7b, 32'hbed5eb44} /* (20, 13, 22) {real, imag} */,
  {32'hbfd450e1, 32'h3f23fb04} /* (20, 13, 21) {real, imag} */,
  {32'h4053ad46, 32'hbf93df98} /* (20, 13, 20) {real, imag} */,
  {32'h3fccc05a, 32'h3df8a4ef} /* (20, 13, 19) {real, imag} */,
  {32'h3f5463bc, 32'hbfb147c8} /* (20, 13, 18) {real, imag} */,
  {32'hbfcb475d, 32'h3f02999c} /* (20, 13, 17) {real, imag} */,
  {32'hbf725cdc, 32'h3f023a15} /* (20, 13, 16) {real, imag} */,
  {32'h3fef02c6, 32'h3e89ffbd} /* (20, 13, 15) {real, imag} */,
  {32'h3f83989e, 32'hbf4b0909} /* (20, 13, 14) {real, imag} */,
  {32'h3d360781, 32'hc0222e50} /* (20, 13, 13) {real, imag} */,
  {32'h3f24a0ad, 32'h3fa8144a} /* (20, 13, 12) {real, imag} */,
  {32'h3e55ccd1, 32'hc0000efe} /* (20, 13, 11) {real, imag} */,
  {32'h40a47bd1, 32'h406c24b8} /* (20, 13, 10) {real, imag} */,
  {32'hc046523c, 32'hbd1e0cee} /* (20, 13, 9) {real, imag} */,
  {32'hbf201674, 32'h3c9e6b9e} /* (20, 13, 8) {real, imag} */,
  {32'hbf313b96, 32'h3fd47a8a} /* (20, 13, 7) {real, imag} */,
  {32'h3f9235a4, 32'h408c313a} /* (20, 13, 6) {real, imag} */,
  {32'h3d3b97bb, 32'hc06d5839} /* (20, 13, 5) {real, imag} */,
  {32'h3fe80a22, 32'hc036ff78} /* (20, 13, 4) {real, imag} */,
  {32'h3fc6c438, 32'h3ff4bbac} /* (20, 13, 3) {real, imag} */,
  {32'hbe9a21e5, 32'hc014432a} /* (20, 13, 2) {real, imag} */,
  {32'h3f11e5bb, 32'h3ef9d52e} /* (20, 13, 1) {real, imag} */,
  {32'hbe01ab71, 32'h40321a55} /* (20, 13, 0) {real, imag} */,
  {32'h3fed8861, 32'h3f7f460e} /* (20, 12, 31) {real, imag} */,
  {32'h3ecbbda3, 32'hbe9e8a03} /* (20, 12, 30) {real, imag} */,
  {32'h3fd51dd9, 32'hbf67d6d7} /* (20, 12, 29) {real, imag} */,
  {32'h3f9fa606, 32'hc03c9b4f} /* (20, 12, 28) {real, imag} */,
  {32'hc0a25162, 32'hbe299506} /* (20, 12, 27) {real, imag} */,
  {32'hbf492fae, 32'hbe674648} /* (20, 12, 26) {real, imag} */,
  {32'h3fa380b4, 32'hc0513992} /* (20, 12, 25) {real, imag} */,
  {32'hbf91079a, 32'h402a2a73} /* (20, 12, 24) {real, imag} */,
  {32'hc02d4b37, 32'h3eb49ea0} /* (20, 12, 23) {real, imag} */,
  {32'hbfbf6323, 32'h40d92c77} /* (20, 12, 22) {real, imag} */,
  {32'h402456f2, 32'hbdc683b1} /* (20, 12, 21) {real, imag} */,
  {32'h3f31460a, 32'hc09e2580} /* (20, 12, 20) {real, imag} */,
  {32'h40000c0e, 32'hbf060037} /* (20, 12, 19) {real, imag} */,
  {32'h3dbb61f5, 32'hbfd58787} /* (20, 12, 18) {real, imag} */,
  {32'hbfa7af62, 32'h3f329bab} /* (20, 12, 17) {real, imag} */,
  {32'hbf45ec5e, 32'hbec178e2} /* (20, 12, 16) {real, imag} */,
  {32'h3fb2ca3e, 32'hc004b91c} /* (20, 12, 15) {real, imag} */,
  {32'hbfe791f2, 32'hbfe64d6e} /* (20, 12, 14) {real, imag} */,
  {32'h3fe079d6, 32'hbf7a8fc4} /* (20, 12, 13) {real, imag} */,
  {32'h404e570b, 32'hbfa46307} /* (20, 12, 12) {real, imag} */,
  {32'hc042d8b7, 32'hbfb44acb} /* (20, 12, 11) {real, imag} */,
  {32'h3e620893, 32'h3ec95777} /* (20, 12, 10) {real, imag} */,
  {32'h3fcc84b5, 32'hbf813d2a} /* (20, 12, 9) {real, imag} */,
  {32'hc08107bc, 32'hbe1adae1} /* (20, 12, 8) {real, imag} */,
  {32'hbecba4a3, 32'h3fcb954a} /* (20, 12, 7) {real, imag} */,
  {32'h3fc89cf1, 32'h3ec18edf} /* (20, 12, 6) {real, imag} */,
  {32'h3fcddf16, 32'hbf1b6258} /* (20, 12, 5) {real, imag} */,
  {32'hbfd8071a, 32'hbe045b21} /* (20, 12, 4) {real, imag} */,
  {32'h3fcb420b, 32'h40048403} /* (20, 12, 3) {real, imag} */,
  {32'hbf162136, 32'h40908909} /* (20, 12, 2) {real, imag} */,
  {32'h3fbd0add, 32'h3fa5a5aa} /* (20, 12, 1) {real, imag} */,
  {32'hbe128460, 32'hbf598984} /* (20, 12, 0) {real, imag} */,
  {32'h3fa85bcb, 32'hbfc7a285} /* (20, 11, 31) {real, imag} */,
  {32'h3fd3816e, 32'h40132395} /* (20, 11, 30) {real, imag} */,
  {32'hbcb44756, 32'hbff59807} /* (20, 11, 29) {real, imag} */,
  {32'h3f80b937, 32'h40589461} /* (20, 11, 28) {real, imag} */,
  {32'h4033f85c, 32'h3fa83b92} /* (20, 11, 27) {real, imag} */,
  {32'hc017fbdd, 32'hbfc055f7} /* (20, 11, 26) {real, imag} */,
  {32'h4045b4e8, 32'h3fe5f36b} /* (20, 11, 25) {real, imag} */,
  {32'hbfe75fdd, 32'hbeee877c} /* (20, 11, 24) {real, imag} */,
  {32'h3f90abcf, 32'h3fd914e9} /* (20, 11, 23) {real, imag} */,
  {32'hc040b3fb, 32'hc079b743} /* (20, 11, 22) {real, imag} */,
  {32'hbfd7059a, 32'h3f304f91} /* (20, 11, 21) {real, imag} */,
  {32'h3fc5bcdb, 32'h3fc745ba} /* (20, 11, 20) {real, imag} */,
  {32'h3fcf0d43, 32'hbf553332} /* (20, 11, 19) {real, imag} */,
  {32'hbdcffaf0, 32'hbf8bb87a} /* (20, 11, 18) {real, imag} */,
  {32'h3f0e5e18, 32'hbf5ff3c3} /* (20, 11, 17) {real, imag} */,
  {32'h3d539b9c, 32'h3f161b55} /* (20, 11, 16) {real, imag} */,
  {32'hbfc2ac5f, 32'h3d677150} /* (20, 11, 15) {real, imag} */,
  {32'h3e5012f7, 32'h4001c318} /* (20, 11, 14) {real, imag} */,
  {32'hc03a52ab, 32'h404851ce} /* (20, 11, 13) {real, imag} */,
  {32'hc02e0748, 32'h401d143f} /* (20, 11, 12) {real, imag} */,
  {32'h400c89d4, 32'hc070fbd3} /* (20, 11, 11) {real, imag} */,
  {32'hbdd6d806, 32'hbfe41515} /* (20, 11, 10) {real, imag} */,
  {32'h402c37e0, 32'hc015b7d2} /* (20, 11, 9) {real, imag} */,
  {32'h400ff4dc, 32'hbfbef08c} /* (20, 11, 8) {real, imag} */,
  {32'hc03c3087, 32'h3f50c036} /* (20, 11, 7) {real, imag} */,
  {32'hbe0801d2, 32'h3f0ddcf6} /* (20, 11, 6) {real, imag} */,
  {32'hc0192ce6, 32'hbfa13f2d} /* (20, 11, 5) {real, imag} */,
  {32'h3fe95e1c, 32'h3f0df359} /* (20, 11, 4) {real, imag} */,
  {32'hbf9f638d, 32'h3fc09dfa} /* (20, 11, 3) {real, imag} */,
  {32'h3fa2b3fa, 32'h3ef87f0b} /* (20, 11, 2) {real, imag} */,
  {32'h3f1a279d, 32'hbfa536c2} /* (20, 11, 1) {real, imag} */,
  {32'h3ee6b147, 32'h3f0fdb89} /* (20, 11, 0) {real, imag} */,
  {32'hbeafe728, 32'hc0518868} /* (20, 10, 31) {real, imag} */,
  {32'h40317ff4, 32'hbe3c16b3} /* (20, 10, 30) {real, imag} */,
  {32'h40474c6c, 32'h3fa57442} /* (20, 10, 29) {real, imag} */,
  {32'hbe10e74c, 32'h3fdaed98} /* (20, 10, 28) {real, imag} */,
  {32'h3fe6b7ab, 32'hbf111498} /* (20, 10, 27) {real, imag} */,
  {32'h3fd35737, 32'h405b7784} /* (20, 10, 26) {real, imag} */,
  {32'hbf896959, 32'h3fa5ba82} /* (20, 10, 25) {real, imag} */,
  {32'hc00728ff, 32'h3ebf3568} /* (20, 10, 24) {real, imag} */,
  {32'h3f456b61, 32'hbdee141e} /* (20, 10, 23) {real, imag} */,
  {32'hbfc56a2f, 32'hbf3396de} /* (20, 10, 22) {real, imag} */,
  {32'hbfbbe448, 32'hc00d613e} /* (20, 10, 21) {real, imag} */,
  {32'hc0240904, 32'h3f66da9d} /* (20, 10, 20) {real, imag} */,
  {32'hbf4304b2, 32'hbed97482} /* (20, 10, 19) {real, imag} */,
  {32'h3e430285, 32'hbf8cc265} /* (20, 10, 18) {real, imag} */,
  {32'h3fa3808d, 32'h3ffa907d} /* (20, 10, 17) {real, imag} */,
  {32'h3ff5a745, 32'hc06101d0} /* (20, 10, 16) {real, imag} */,
  {32'hbf19d1e3, 32'h3e1972fc} /* (20, 10, 15) {real, imag} */,
  {32'hc0042e7e, 32'hbf604428} /* (20, 10, 14) {real, imag} */,
  {32'hbec58dbe, 32'h3f22b557} /* (20, 10, 13) {real, imag} */,
  {32'h3f042e83, 32'hbf0e1aaf} /* (20, 10, 12) {real, imag} */,
  {32'h3ff9fd79, 32'h3d565956} /* (20, 10, 11) {real, imag} */,
  {32'h40246315, 32'hc068c343} /* (20, 10, 10) {real, imag} */,
  {32'hbc1a73fe, 32'h3f10ce72} /* (20, 10, 9) {real, imag} */,
  {32'h3fd42b4c, 32'h3fa5469c} /* (20, 10, 8) {real, imag} */,
  {32'h400a20dd, 32'hc012d7b1} /* (20, 10, 7) {real, imag} */,
  {32'hbe395746, 32'hbf896ce0} /* (20, 10, 6) {real, imag} */,
  {32'h3f601b2f, 32'h405cfd22} /* (20, 10, 5) {real, imag} */,
  {32'h3fcf89fe, 32'h3f9de663} /* (20, 10, 4) {real, imag} */,
  {32'hc0a8f58e, 32'h3f27790f} /* (20, 10, 3) {real, imag} */,
  {32'h401dc9b2, 32'h3ca9325e} /* (20, 10, 2) {real, imag} */,
  {32'hc02d40f7, 32'hbde06018} /* (20, 10, 1) {real, imag} */,
  {32'hbe402dbb, 32'hc02677c2} /* (20, 10, 0) {real, imag} */,
  {32'hbffc706a, 32'hbf29ba2e} /* (20, 9, 31) {real, imag} */,
  {32'h3fcfff49, 32'h3f707ef2} /* (20, 9, 30) {real, imag} */,
  {32'hbe757597, 32'hbea71633} /* (20, 9, 29) {real, imag} */,
  {32'hbf6e051b, 32'hc014a646} /* (20, 9, 28) {real, imag} */,
  {32'hbd9007c4, 32'hc01f188c} /* (20, 9, 27) {real, imag} */,
  {32'hbf15812e, 32'hc00bbd13} /* (20, 9, 26) {real, imag} */,
  {32'h3fae62f5, 32'h3f25ea80} /* (20, 9, 25) {real, imag} */,
  {32'hbe1ff9b9, 32'hbf079d47} /* (20, 9, 24) {real, imag} */,
  {32'h3f280a6b, 32'h3f77728c} /* (20, 9, 23) {real, imag} */,
  {32'h3ed11ffa, 32'hbc3d4c60} /* (20, 9, 22) {real, imag} */,
  {32'hbf2779bb, 32'h3f8490eb} /* (20, 9, 21) {real, imag} */,
  {32'hbf490462, 32'h407f7605} /* (20, 9, 20) {real, imag} */,
  {32'h4037df22, 32'hc011a829} /* (20, 9, 19) {real, imag} */,
  {32'h3f2085de, 32'h3feb3b71} /* (20, 9, 18) {real, imag} */,
  {32'hbf21fc06, 32'h3eac4071} /* (20, 9, 17) {real, imag} */,
  {32'h3e6c1117, 32'hbfbef189} /* (20, 9, 16) {real, imag} */,
  {32'hbf031162, 32'h3fb53561} /* (20, 9, 15) {real, imag} */,
  {32'h3f8ca945, 32'h40408828} /* (20, 9, 14) {real, imag} */,
  {32'hbeea3c64, 32'hc0824a3c} /* (20, 9, 13) {real, imag} */,
  {32'h4067ea49, 32'h3fce8079} /* (20, 9, 12) {real, imag} */,
  {32'h400b6520, 32'h3f8dff7b} /* (20, 9, 11) {real, imag} */,
  {32'hbf8111a1, 32'h3fc83b35} /* (20, 9, 10) {real, imag} */,
  {32'hbfdfd3cf, 32'h3f9bc7b6} /* (20, 9, 9) {real, imag} */,
  {32'hbff2e9b5, 32'h3fc4ae6b} /* (20, 9, 8) {real, imag} */,
  {32'h3f1bbde3, 32'hbf352d3e} /* (20, 9, 7) {real, imag} */,
  {32'h3e839b7b, 32'hc041fb1d} /* (20, 9, 6) {real, imag} */,
  {32'h4075b5ab, 32'h3fc2accf} /* (20, 9, 5) {real, imag} */,
  {32'hc00fc45b, 32'h3fa5729d} /* (20, 9, 4) {real, imag} */,
  {32'h3fa79f4b, 32'hbfe1e93a} /* (20, 9, 3) {real, imag} */,
  {32'hbf7bc307, 32'h3d9a20ae} /* (20, 9, 2) {real, imag} */,
  {32'hbf12e421, 32'h4080a40b} /* (20, 9, 1) {real, imag} */,
  {32'hc002456d, 32'hc001a142} /* (20, 9, 0) {real, imag} */,
  {32'hbf8e8727, 32'hbe1b72bd} /* (20, 8, 31) {real, imag} */,
  {32'hbfb5873d, 32'hbfd1831b} /* (20, 8, 30) {real, imag} */,
  {32'hc0201642, 32'h3e98109a} /* (20, 8, 29) {real, imag} */,
  {32'h3fbf35cf, 32'hbf4392da} /* (20, 8, 28) {real, imag} */,
  {32'h3f1a445b, 32'hbf47c0d9} /* (20, 8, 27) {real, imag} */,
  {32'h3dc46363, 32'h3ebf2758} /* (20, 8, 26) {real, imag} */,
  {32'hbf759b33, 32'h3f87ee7e} /* (20, 8, 25) {real, imag} */,
  {32'hbf0b017d, 32'hc05c489e} /* (20, 8, 24) {real, imag} */,
  {32'h3fac76a8, 32'h3fbc7409} /* (20, 8, 23) {real, imag} */,
  {32'h3eee08ff, 32'hc0359582} /* (20, 8, 22) {real, imag} */,
  {32'h3f4d703f, 32'h4031fcbb} /* (20, 8, 21) {real, imag} */,
  {32'h3e66aeef, 32'hbf959640} /* (20, 8, 20) {real, imag} */,
  {32'h3ee6965f, 32'hbe9671e5} /* (20, 8, 19) {real, imag} */,
  {32'h3e4cb5ae, 32'hbfc9c3e3} /* (20, 8, 18) {real, imag} */,
  {32'hbf004c7f, 32'h3ed08236} /* (20, 8, 17) {real, imag} */,
  {32'h3f3c0c17, 32'h3f329603} /* (20, 8, 16) {real, imag} */,
  {32'h3f1bfc9a, 32'hbf42b4fe} /* (20, 8, 15) {real, imag} */,
  {32'hc0181875, 32'h4018b43e} /* (20, 8, 14) {real, imag} */,
  {32'h40962234, 32'hbf08ec1b} /* (20, 8, 13) {real, imag} */,
  {32'h40557013, 32'hc081590c} /* (20, 8, 12) {real, imag} */,
  {32'hbf2c155d, 32'h3ff6a43c} /* (20, 8, 11) {real, imag} */,
  {32'hc09071da, 32'hc064fafa} /* (20, 8, 10) {real, imag} */,
  {32'hbcb75507, 32'hbfab7943} /* (20, 8, 9) {real, imag} */,
  {32'hbb6b258f, 32'hc02333b4} /* (20, 8, 8) {real, imag} */,
  {32'hc0536a38, 32'h3e1607db} /* (20, 8, 7) {real, imag} */,
  {32'h3f7741c3, 32'hc073b581} /* (20, 8, 6) {real, imag} */,
  {32'hbf3c0d97, 32'h406f8b0c} /* (20, 8, 5) {real, imag} */,
  {32'hc002eac2, 32'hbfcdac38} /* (20, 8, 4) {real, imag} */,
  {32'h3f8e558e, 32'hc0871654} /* (20, 8, 3) {real, imag} */,
  {32'hbf8dd066, 32'hbf42f672} /* (20, 8, 2) {real, imag} */,
  {32'h3f1b54f4, 32'h3f804f9b} /* (20, 8, 1) {real, imag} */,
  {32'h406ebcf4, 32'hbe25a5e2} /* (20, 8, 0) {real, imag} */,
  {32'h3f0a9506, 32'h403da33f} /* (20, 7, 31) {real, imag} */,
  {32'hbf2427b1, 32'hbe85bc84} /* (20, 7, 30) {real, imag} */,
  {32'hc0006f24, 32'h406ff3e6} /* (20, 7, 29) {real, imag} */,
  {32'hbe756771, 32'hbf9c6da0} /* (20, 7, 28) {real, imag} */,
  {32'h3d8ac1c2, 32'h3f838d28} /* (20, 7, 27) {real, imag} */,
  {32'h3fea54c7, 32'hc06e6f20} /* (20, 7, 26) {real, imag} */,
  {32'h3f8b47be, 32'h3fdfacb5} /* (20, 7, 25) {real, imag} */,
  {32'h3f0b2098, 32'h3f41343c} /* (20, 7, 24) {real, imag} */,
  {32'hbfddafae, 32'h3f72d25e} /* (20, 7, 23) {real, imag} */,
  {32'h3fd4fc8a, 32'h3ff71eb0} /* (20, 7, 22) {real, imag} */,
  {32'h3e8010d2, 32'h3fc7c573} /* (20, 7, 21) {real, imag} */,
  {32'h3ef015f5, 32'hbf1c3a04} /* (20, 7, 20) {real, imag} */,
  {32'hbeb0f837, 32'hbe4e6461} /* (20, 7, 19) {real, imag} */,
  {32'h400e8f0b, 32'h3e73b03b} /* (20, 7, 18) {real, imag} */,
  {32'hbfb15f30, 32'hbed60e27} /* (20, 7, 17) {real, imag} */,
  {32'hc017cc6c, 32'h3df61074} /* (20, 7, 16) {real, imag} */,
  {32'hbf8dfd73, 32'h3fabaae1} /* (20, 7, 15) {real, imag} */,
  {32'h401d5de9, 32'h3f7fd037} /* (20, 7, 14) {real, imag} */,
  {32'hbe91cade, 32'h40250f97} /* (20, 7, 13) {real, imag} */,
  {32'hbfac9207, 32'hbf37ee51} /* (20, 7, 12) {real, imag} */,
  {32'h3ec433b9, 32'h3f175f86} /* (20, 7, 11) {real, imag} */,
  {32'hbfec8db3, 32'h4006af4b} /* (20, 7, 10) {real, imag} */,
  {32'h401e0b23, 32'h3fb27d6e} /* (20, 7, 9) {real, imag} */,
  {32'hbfe21c87, 32'h4071f08b} /* (20, 7, 8) {real, imag} */,
  {32'h3f1c3181, 32'hbf2695f8} /* (20, 7, 7) {real, imag} */,
  {32'h40278247, 32'hbfd119a7} /* (20, 7, 6) {real, imag} */,
  {32'hc023a366, 32'hbfded2a8} /* (20, 7, 5) {real, imag} */,
  {32'hbf97acf1, 32'hbf8a011c} /* (20, 7, 4) {real, imag} */,
  {32'hbeca7ea4, 32'hbf4d4516} /* (20, 7, 3) {real, imag} */,
  {32'h402476d2, 32'hbf092fe3} /* (20, 7, 2) {real, imag} */,
  {32'h3fa32e66, 32'hbfdbdaf3} /* (20, 7, 1) {real, imag} */,
  {32'hbfd58b62, 32'hbfb5f782} /* (20, 7, 0) {real, imag} */,
  {32'hbfaa0cbb, 32'h3f08cde2} /* (20, 6, 31) {real, imag} */,
  {32'hc0756c00, 32'hbf947e50} /* (20, 6, 30) {real, imag} */,
  {32'h3f8e87d6, 32'hc020817b} /* (20, 6, 29) {real, imag} */,
  {32'h3fc8ce81, 32'h3efa17f0} /* (20, 6, 28) {real, imag} */,
  {32'h401d5eef, 32'h3f318257} /* (20, 6, 27) {real, imag} */,
  {32'hc084394e, 32'h3f56be4d} /* (20, 6, 26) {real, imag} */,
  {32'h3f4ff034, 32'h3f57148b} /* (20, 6, 25) {real, imag} */,
  {32'h4031dd4c, 32'hbf8b70fb} /* (20, 6, 24) {real, imag} */,
  {32'hbfa5eee3, 32'hbf887ab3} /* (20, 6, 23) {real, imag} */,
  {32'h3ee79523, 32'h3fff9486} /* (20, 6, 22) {real, imag} */,
  {32'hbf3c901a, 32'h3fa7f6aa} /* (20, 6, 21) {real, imag} */,
  {32'hbf7053ca, 32'hc024ce4c} /* (20, 6, 20) {real, imag} */,
  {32'h4032dacb, 32'h3e1545dd} /* (20, 6, 19) {real, imag} */,
  {32'h3ee4fefb, 32'hc012ec89} /* (20, 6, 18) {real, imag} */,
  {32'h3fc33686, 32'h3f78fa83} /* (20, 6, 17) {real, imag} */,
  {32'hbd8b7b59, 32'h3f59cc7b} /* (20, 6, 16) {real, imag} */,
  {32'hbfbe24e8, 32'hbfd1966a} /* (20, 6, 15) {real, imag} */,
  {32'h3fefdd36, 32'hbd8c7160} /* (20, 6, 14) {real, imag} */,
  {32'h3f52a280, 32'h3f65b811} /* (20, 6, 13) {real, imag} */,
  {32'h3fe41644, 32'hbf9b9bad} /* (20, 6, 12) {real, imag} */,
  {32'hbf61b187, 32'h3e823514} /* (20, 6, 11) {real, imag} */,
  {32'h3f1a7cc2, 32'h3ed3e339} /* (20, 6, 10) {real, imag} */,
  {32'hbfe11ebe, 32'hbf9803f9} /* (20, 6, 9) {real, imag} */,
  {32'hbfe39220, 32'hbf92be5c} /* (20, 6, 8) {real, imag} */,
  {32'h405ab3bf, 32'h3dbbf1a9} /* (20, 6, 7) {real, imag} */,
  {32'h3e3b2f4a, 32'h3f989242} /* (20, 6, 6) {real, imag} */,
  {32'h3e778a0c, 32'hbf878b64} /* (20, 6, 5) {real, imag} */,
  {32'hbf2ca3dc, 32'h4073154d} /* (20, 6, 4) {real, imag} */,
  {32'h40329c15, 32'hbf910e56} /* (20, 6, 3) {real, imag} */,
  {32'h3f9d136c, 32'hbd28bd1f} /* (20, 6, 2) {real, imag} */,
  {32'hbfac2b45, 32'hc02f1c1f} /* (20, 6, 1) {real, imag} */,
  {32'hbec6219a, 32'hbe959412} /* (20, 6, 0) {real, imag} */,
  {32'h3f918d6d, 32'hbd5e6d0d} /* (20, 5, 31) {real, imag} */,
  {32'h3e063e45, 32'hbf1031cf} /* (20, 5, 30) {real, imag} */,
  {32'hc033ce62, 32'hbfdf6244} /* (20, 5, 29) {real, imag} */,
  {32'hbf80f8b2, 32'h3e3998f5} /* (20, 5, 28) {real, imag} */,
  {32'h3f5f9e9f, 32'h3fd03172} /* (20, 5, 27) {real, imag} */,
  {32'hbf14720f, 32'h40344ea8} /* (20, 5, 26) {real, imag} */,
  {32'hbf634473, 32'h3ee745a0} /* (20, 5, 25) {real, imag} */,
  {32'hc056dcea, 32'hbf790597} /* (20, 5, 24) {real, imag} */,
  {32'h40077c28, 32'h40533c57} /* (20, 5, 23) {real, imag} */,
  {32'hbf6c48d1, 32'hbebaf89f} /* (20, 5, 22) {real, imag} */,
  {32'hc004d13c, 32'hc073f2b1} /* (20, 5, 21) {real, imag} */,
  {32'hbeb81324, 32'h40054147} /* (20, 5, 20) {real, imag} */,
  {32'h3f3b69fd, 32'hbf3d08b9} /* (20, 5, 19) {real, imag} */,
  {32'hbfb33a99, 32'h3f1b57d3} /* (20, 5, 18) {real, imag} */,
  {32'h3f34d7bc, 32'h3de3fee8} /* (20, 5, 17) {real, imag} */,
  {32'hbfdd5939, 32'h3eacf1d8} /* (20, 5, 16) {real, imag} */,
  {32'hbe65ee37, 32'h3fc20f72} /* (20, 5, 15) {real, imag} */,
  {32'h3e06f591, 32'h3f52e916} /* (20, 5, 14) {real, imag} */,
  {32'h3e5df4a1, 32'h3fb1194c} /* (20, 5, 13) {real, imag} */,
  {32'hbe197aa5, 32'hbf829bd8} /* (20, 5, 12) {real, imag} */,
  {32'h40154bfe, 32'h3f03113c} /* (20, 5, 11) {real, imag} */,
  {32'hbfb8f875, 32'hbeffda43} /* (20, 5, 10) {real, imag} */,
  {32'hc006e7ce, 32'h3fc88063} /* (20, 5, 9) {real, imag} */,
  {32'hbe2966ec, 32'hc057ac12} /* (20, 5, 8) {real, imag} */,
  {32'h400f9332, 32'hbfffac1e} /* (20, 5, 7) {real, imag} */,
  {32'hbfe9aff0, 32'h3fade756} /* (20, 5, 6) {real, imag} */,
  {32'hbfe2c7af, 32'h401e6a55} /* (20, 5, 5) {real, imag} */,
  {32'hbf01f52e, 32'h401149bf} /* (20, 5, 4) {real, imag} */,
  {32'hbf81a7b6, 32'hbeeed2a6} /* (20, 5, 3) {real, imag} */,
  {32'hbfbeab12, 32'hbba6dcf5} /* (20, 5, 2) {real, imag} */,
  {32'h3f93b6cf, 32'h400f80a2} /* (20, 5, 1) {real, imag} */,
  {32'h3f9e5285, 32'h3f2a5b82} /* (20, 5, 0) {real, imag} */,
  {32'h3f69dc05, 32'hbeab84dd} /* (20, 4, 31) {real, imag} */,
  {32'h3fc0fdfe, 32'hbfa65a87} /* (20, 4, 30) {real, imag} */,
  {32'hc01bcc4a, 32'h3e52d956} /* (20, 4, 29) {real, imag} */,
  {32'hbf5765d8, 32'hbeea82cb} /* (20, 4, 28) {real, imag} */,
  {32'h3cd26528, 32'h405c09a1} /* (20, 4, 27) {real, imag} */,
  {32'h4015ed4f, 32'h3f95b10c} /* (20, 4, 26) {real, imag} */,
  {32'h3f1eb2dd, 32'h3e9880d0} /* (20, 4, 25) {real, imag} */,
  {32'hc023f797, 32'hc024cfea} /* (20, 4, 24) {real, imag} */,
  {32'h40104a83, 32'hbf8863ec} /* (20, 4, 23) {real, imag} */,
  {32'h3fbfb096, 32'hbfed7e91} /* (20, 4, 22) {real, imag} */,
  {32'hc066fa13, 32'hbf712fe4} /* (20, 4, 21) {real, imag} */,
  {32'hbfbf9734, 32'h3f12524b} /* (20, 4, 20) {real, imag} */,
  {32'h3f2c3640, 32'hbe2ed077} /* (20, 4, 19) {real, imag} */,
  {32'h3f1f0c2c, 32'h40306c07} /* (20, 4, 18) {real, imag} */,
  {32'h3f574873, 32'hbfaaabe1} /* (20, 4, 17) {real, imag} */,
  {32'hbec1b1cb, 32'h3ef51fca} /* (20, 4, 16) {real, imag} */,
  {32'h3f67a946, 32'hbf2b57f6} /* (20, 4, 15) {real, imag} */,
  {32'h3fa40293, 32'hbe9ad510} /* (20, 4, 14) {real, imag} */,
  {32'hbfd69bc0, 32'hbfc8c46d} /* (20, 4, 13) {real, imag} */,
  {32'h3fa49e7a, 32'h3e522390} /* (20, 4, 12) {real, imag} */,
  {32'hbe93e3f6, 32'hbf4b3618} /* (20, 4, 11) {real, imag} */,
  {32'hc06cd84e, 32'hbff78efc} /* (20, 4, 10) {real, imag} */,
  {32'h3ef01ccf, 32'h4059acc6} /* (20, 4, 9) {real, imag} */,
  {32'hbfbf8a65, 32'h3f6ccd61} /* (20, 4, 8) {real, imag} */,
  {32'h3ee1d115, 32'h40000a1b} /* (20, 4, 7) {real, imag} */,
  {32'hbdfab129, 32'hbf6f6817} /* (20, 4, 6) {real, imag} */,
  {32'hc016ef47, 32'h3e7c64f9} /* (20, 4, 5) {real, imag} */,
  {32'h3ede4271, 32'hbf967aff} /* (20, 4, 4) {real, imag} */,
  {32'hbf034a98, 32'h3ffe966c} /* (20, 4, 3) {real, imag} */,
  {32'hc0008d7d, 32'hbf8f8212} /* (20, 4, 2) {real, imag} */,
  {32'hbf200783, 32'hbf6ad6d3} /* (20, 4, 1) {real, imag} */,
  {32'h3f1f386a, 32'hc0008e0b} /* (20, 4, 0) {real, imag} */,
  {32'h3f3a4129, 32'h4030a671} /* (20, 3, 31) {real, imag} */,
  {32'h3f926d01, 32'hbf468f35} /* (20, 3, 30) {real, imag} */,
  {32'hbf35df50, 32'h4099ecdc} /* (20, 3, 29) {real, imag} */,
  {32'h3fd24078, 32'hc02db80c} /* (20, 3, 28) {real, imag} */,
  {32'hbf97b651, 32'h3ea891ad} /* (20, 3, 27) {real, imag} */,
  {32'h3e8c103a, 32'h3fc6d3da} /* (20, 3, 26) {real, imag} */,
  {32'h3f945b3c, 32'h405ab407} /* (20, 3, 25) {real, imag} */,
  {32'hbfda5028, 32'h3ed1a5d8} /* (20, 3, 24) {real, imag} */,
  {32'hbee8be94, 32'hbd3ce824} /* (20, 3, 23) {real, imag} */,
  {32'hc0309cc5, 32'hbfa4ec57} /* (20, 3, 22) {real, imag} */,
  {32'h3adb17d8, 32'h3f40f567} /* (20, 3, 21) {real, imag} */,
  {32'h3fd54999, 32'h3f1ecb03} /* (20, 3, 20) {real, imag} */,
  {32'hbf47c8f3, 32'h3f75001f} /* (20, 3, 19) {real, imag} */,
  {32'hbf58b9a7, 32'h3fda278c} /* (20, 3, 18) {real, imag} */,
  {32'hbdf17ff5, 32'h3f153b8a} /* (20, 3, 17) {real, imag} */,
  {32'h3ea72d25, 32'hbf17c891} /* (20, 3, 16) {real, imag} */,
  {32'hc00e9726, 32'hc0202454} /* (20, 3, 15) {real, imag} */,
  {32'h3ed6ee6f, 32'hbe8de53e} /* (20, 3, 14) {real, imag} */,
  {32'hc0386609, 32'hbf8be949} /* (20, 3, 13) {real, imag} */,
  {32'hbf2128fe, 32'h40237b9b} /* (20, 3, 12) {real, imag} */,
  {32'hbee0aa15, 32'hbe5ecaca} /* (20, 3, 11) {real, imag} */,
  {32'hbecaa01b, 32'hc05fdafd} /* (20, 3, 10) {real, imag} */,
  {32'h3fc0b84c, 32'h3f9b510e} /* (20, 3, 9) {real, imag} */,
  {32'h40063d5c, 32'hbfbec654} /* (20, 3, 8) {real, imag} */,
  {32'hbe7cabf5, 32'h3f99d7b7} /* (20, 3, 7) {real, imag} */,
  {32'hbe24f9a9, 32'hbe0fff0d} /* (20, 3, 6) {real, imag} */,
  {32'h3e8b88d1, 32'hbf2251c8} /* (20, 3, 5) {real, imag} */,
  {32'h3fe60eac, 32'h3fc606c1} /* (20, 3, 4) {real, imag} */,
  {32'h3ffe5b77, 32'h400c60db} /* (20, 3, 3) {real, imag} */,
  {32'h4005eaf3, 32'h3f4da739} /* (20, 3, 2) {real, imag} */,
  {32'h3ef3b9c0, 32'hc0a34614} /* (20, 3, 1) {real, imag} */,
  {32'h3eed901c, 32'h3e7dfc2e} /* (20, 3, 0) {real, imag} */,
  {32'h3fdc1830, 32'hc0a31230} /* (20, 2, 31) {real, imag} */,
  {32'hbf748537, 32'hbdc3fb60} /* (20, 2, 30) {real, imag} */,
  {32'h40432d51, 32'h40052cc1} /* (20, 2, 29) {real, imag} */,
  {32'h3d70608b, 32'h401003d9} /* (20, 2, 28) {real, imag} */,
  {32'h3fb54a8e, 32'h3f800d31} /* (20, 2, 27) {real, imag} */,
  {32'h3fb94a0b, 32'hbf75cf09} /* (20, 2, 26) {real, imag} */,
  {32'h4084d19e, 32'h3f5df565} /* (20, 2, 25) {real, imag} */,
  {32'hbebfd46c, 32'h3e1c3ae9} /* (20, 2, 24) {real, imag} */,
  {32'hbf32a676, 32'hbfab55cd} /* (20, 2, 23) {real, imag} */,
  {32'hbdaf0a77, 32'hbec9862f} /* (20, 2, 22) {real, imag} */,
  {32'hbdec559b, 32'hbf8b4a9f} /* (20, 2, 21) {real, imag} */,
  {32'h3f21f1a8, 32'h3e3e4814} /* (20, 2, 20) {real, imag} */,
  {32'hbf6ff8ce, 32'hbe5ada41} /* (20, 2, 19) {real, imag} */,
  {32'h3fc2849b, 32'h3faae9f2} /* (20, 2, 18) {real, imag} */,
  {32'h3f8619d6, 32'h3fa17f75} /* (20, 2, 17) {real, imag} */,
  {32'hbf7590ba, 32'h3f9e4966} /* (20, 2, 16) {real, imag} */,
  {32'hbf852081, 32'hbeb23713} /* (20, 2, 15) {real, imag} */,
  {32'hbfef57c9, 32'hbf8144ab} /* (20, 2, 14) {real, imag} */,
  {32'hbf4822bf, 32'h3efdb01f} /* (20, 2, 13) {real, imag} */,
  {32'h4058abb9, 32'hc018998c} /* (20, 2, 12) {real, imag} */,
  {32'hc0054e60, 32'hbed60041} /* (20, 2, 11) {real, imag} */,
  {32'hbf062f74, 32'hbe63489f} /* (20, 2, 10) {real, imag} */,
  {32'h3fe0d7fe, 32'hbee4fd5a} /* (20, 2, 9) {real, imag} */,
  {32'h3fa39cd9, 32'hbed54fe1} /* (20, 2, 8) {real, imag} */,
  {32'h3fe4549b, 32'hc014a118} /* (20, 2, 7) {real, imag} */,
  {32'h3f7c7eeb, 32'h3e22ae1c} /* (20, 2, 6) {real, imag} */,
  {32'h3fc443dd, 32'h3f70d5df} /* (20, 2, 5) {real, imag} */,
  {32'h3eb73e12, 32'h3f42c140} /* (20, 2, 4) {real, imag} */,
  {32'h3fd7b40f, 32'hbfaf0664} /* (20, 2, 3) {real, imag} */,
  {32'hc01323ab, 32'hbf4a1eb7} /* (20, 2, 2) {real, imag} */,
  {32'hbf5a4b5f, 32'h3ef661fc} /* (20, 2, 1) {real, imag} */,
  {32'h3f0907e4, 32'h3fcb7206} /* (20, 2, 0) {real, imag} */,
  {32'hbfb7e887, 32'h3ebda4ea} /* (20, 1, 31) {real, imag} */,
  {32'hbe1389bb, 32'hbf434144} /* (20, 1, 30) {real, imag} */,
  {32'h3fa398ab, 32'hbf110027} /* (20, 1, 29) {real, imag} */,
  {32'hbfa003cf, 32'h3e85d632} /* (20, 1, 28) {real, imag} */,
  {32'h400d385f, 32'h3fbb7db6} /* (20, 1, 27) {real, imag} */,
  {32'h3f4f2ae7, 32'hbfd11fd7} /* (20, 1, 26) {real, imag} */,
  {32'hbf613532, 32'hbf473900} /* (20, 1, 25) {real, imag} */,
  {32'h3fd00779, 32'hbeee4179} /* (20, 1, 24) {real, imag} */,
  {32'h4030353e, 32'hbe429bb6} /* (20, 1, 23) {real, imag} */,
  {32'h402fe66c, 32'h3f0babba} /* (20, 1, 22) {real, imag} */,
  {32'hbfaf7141, 32'hc08d86cf} /* (20, 1, 21) {real, imag} */,
  {32'h3f325091, 32'h3f06b9ea} /* (20, 1, 20) {real, imag} */,
  {32'h3fe647d7, 32'hc0536300} /* (20, 1, 19) {real, imag} */,
  {32'h3d12c71d, 32'hbd8cb836} /* (20, 1, 18) {real, imag} */,
  {32'hc016d070, 32'hc0024d60} /* (20, 1, 17) {real, imag} */,
  {32'hbb65d508, 32'h3f83f9c5} /* (20, 1, 16) {real, imag} */,
  {32'hbf6cbdac, 32'hbec5a969} /* (20, 1, 15) {real, imag} */,
  {32'h401bda2d, 32'hbf541e5c} /* (20, 1, 14) {real, imag} */,
  {32'h3eeb5468, 32'hbffaadee} /* (20, 1, 13) {real, imag} */,
  {32'h3e295be1, 32'h3eec99ab} /* (20, 1, 12) {real, imag} */,
  {32'h40602b63, 32'h3f724f7e} /* (20, 1, 11) {real, imag} */,
  {32'hc00c2906, 32'h3f6995d6} /* (20, 1, 10) {real, imag} */,
  {32'hbee9764b, 32'hbf28ee77} /* (20, 1, 9) {real, imag} */,
  {32'hbfdda269, 32'hbf1da6f0} /* (20, 1, 8) {real, imag} */,
  {32'h3ff28215, 32'hc0608b89} /* (20, 1, 7) {real, imag} */,
  {32'hc0475e0b, 32'h3da474d5} /* (20, 1, 6) {real, imag} */,
  {32'hbf0796c6, 32'hbf2104a0} /* (20, 1, 5) {real, imag} */,
  {32'h3dd25a15, 32'h401dddca} /* (20, 1, 4) {real, imag} */,
  {32'hbfb617dd, 32'h3f846d04} /* (20, 1, 3) {real, imag} */,
  {32'hc047278d, 32'hbe8a880b} /* (20, 1, 2) {real, imag} */,
  {32'hc0353655, 32'hbf6c2883} /* (20, 1, 1) {real, imag} */,
  {32'h3fd3f4f3, 32'hbfb0827a} /* (20, 1, 0) {real, imag} */,
  {32'h3ed627e2, 32'h3fd78dc6} /* (20, 0, 31) {real, imag} */,
  {32'hbf80ea4a, 32'hc010e22c} /* (20, 0, 30) {real, imag} */,
  {32'hc019341b, 32'hbed24ddb} /* (20, 0, 29) {real, imag} */,
  {32'h3fad0d11, 32'h3f5f9cba} /* (20, 0, 28) {real, imag} */,
  {32'hc0106c4f, 32'h3eca04a9} /* (20, 0, 27) {real, imag} */,
  {32'h4093aa2b, 32'hc00bc0a3} /* (20, 0, 26) {real, imag} */,
  {32'hbf1e5af9, 32'h3e4613f1} /* (20, 0, 25) {real, imag} */,
  {32'h3fcb0c0a, 32'h3ea4cb91} /* (20, 0, 24) {real, imag} */,
  {32'h40528817, 32'h40443fd5} /* (20, 0, 23) {real, imag} */,
  {32'h3f4d741b, 32'h400667d6} /* (20, 0, 22) {real, imag} */,
  {32'h3f045e72, 32'h3fb5ac5e} /* (20, 0, 21) {real, imag} */,
  {32'hbff2f38e, 32'h3febb336} /* (20, 0, 20) {real, imag} */,
  {32'hbef7d602, 32'h3f833efe} /* (20, 0, 19) {real, imag} */,
  {32'h3fafb135, 32'h3f2da643} /* (20, 0, 18) {real, imag} */,
  {32'h3eb858e2, 32'hbfe1bb52} /* (20, 0, 17) {real, imag} */,
  {32'hbe435355, 32'h3ee851c1} /* (20, 0, 16) {real, imag} */,
  {32'hbeeb5e17, 32'h3f269a52} /* (20, 0, 15) {real, imag} */,
  {32'h3de21874, 32'hc024b3b3} /* (20, 0, 14) {real, imag} */,
  {32'h3f2a932c, 32'h4057eda3} /* (20, 0, 13) {real, imag} */,
  {32'h3f0215d5, 32'h3fa7046b} /* (20, 0, 12) {real, imag} */,
  {32'hc037ffef, 32'hbe1d6dbe} /* (20, 0, 11) {real, imag} */,
  {32'h3f8ef3e4, 32'h3e78263b} /* (20, 0, 10) {real, imag} */,
  {32'hbf8f6c2b, 32'hbfa3ec82} /* (20, 0, 9) {real, imag} */,
  {32'h406225d9, 32'hc0027d4a} /* (20, 0, 8) {real, imag} */,
  {32'hbe913aee, 32'hbfe87782} /* (20, 0, 7) {real, imag} */,
  {32'h3fbfebcd, 32'h3feafe26} /* (20, 0, 6) {real, imag} */,
  {32'h404e8951, 32'h407b4beb} /* (20, 0, 5) {real, imag} */,
  {32'h3c306939, 32'hbf97cb17} /* (20, 0, 4) {real, imag} */,
  {32'h3ef90143, 32'h3eac0c34} /* (20, 0, 3) {real, imag} */,
  {32'hbffc9831, 32'h3f503040} /* (20, 0, 2) {real, imag} */,
  {32'hbe8bf94f, 32'hbe16ccc1} /* (20, 0, 1) {real, imag} */,
  {32'hbfa13490, 32'h3feb4004} /* (20, 0, 0) {real, imag} */,
  {32'hc02f143b, 32'h3e4f21ec} /* (19, 31, 31) {real, imag} */,
  {32'hbf22766c, 32'hc01bd976} /* (19, 31, 30) {real, imag} */,
  {32'h3f34f383, 32'h3fa6a455} /* (19, 31, 29) {real, imag} */,
  {32'hbef04e4b, 32'hbfda43ac} /* (19, 31, 28) {real, imag} */,
  {32'hbf68337f, 32'hbeb4016f} /* (19, 31, 27) {real, imag} */,
  {32'h3fcf8fd5, 32'hbe9a1776} /* (19, 31, 26) {real, imag} */,
  {32'hbfd7d06a, 32'h3ea6a295} /* (19, 31, 25) {real, imag} */,
  {32'hbf4a644a, 32'hbe261d30} /* (19, 31, 24) {real, imag} */,
  {32'hbfb90cb1, 32'h40a2682e} /* (19, 31, 23) {real, imag} */,
  {32'h3f8b99b8, 32'hbf1c411d} /* (19, 31, 22) {real, imag} */,
  {32'h4090042d, 32'h3e57b685} /* (19, 31, 21) {real, imag} */,
  {32'hbf69a8ef, 32'h3f62ade9} /* (19, 31, 20) {real, imag} */,
  {32'h3f1c7ead, 32'h3ea37ae2} /* (19, 31, 19) {real, imag} */,
  {32'h3e9c93a4, 32'h3fcbcb22} /* (19, 31, 18) {real, imag} */,
  {32'hbed44af6, 32'hbf75638a} /* (19, 31, 17) {real, imag} */,
  {32'h4007f799, 32'h405c7144} /* (19, 31, 16) {real, imag} */,
  {32'hbfd8a9eb, 32'h3e48fc8e} /* (19, 31, 15) {real, imag} */,
  {32'h3eb2d486, 32'hbf7549cb} /* (19, 31, 14) {real, imag} */,
  {32'h3f8753c5, 32'hbdf1dee6} /* (19, 31, 13) {real, imag} */,
  {32'hc066d15e, 32'hbee91c83} /* (19, 31, 12) {real, imag} */,
  {32'hbfb4f54c, 32'hbf0a6624} /* (19, 31, 11) {real, imag} */,
  {32'h3f97d99d, 32'hbeb031ef} /* (19, 31, 10) {real, imag} */,
  {32'h3f3fd089, 32'hc00a1f28} /* (19, 31, 9) {real, imag} */,
  {32'h400a21f2, 32'hc025278e} /* (19, 31, 8) {real, imag} */,
  {32'h3f25fdee, 32'hbfbc35c2} /* (19, 31, 7) {real, imag} */,
  {32'h3f641856, 32'hbe3c644f} /* (19, 31, 6) {real, imag} */,
  {32'hbf4e480e, 32'hc01dff43} /* (19, 31, 5) {real, imag} */,
  {32'h3f459bc3, 32'h3e0ca201} /* (19, 31, 4) {real, imag} */,
  {32'h407ed389, 32'hbed0b449} /* (19, 31, 3) {real, imag} */,
  {32'h3fc2ecdc, 32'hbf8d7499} /* (19, 31, 2) {real, imag} */,
  {32'h402262d6, 32'hbf40a034} /* (19, 31, 1) {real, imag} */,
  {32'h3fe7ff12, 32'hbf4ef287} /* (19, 31, 0) {real, imag} */,
  {32'h3fb7d2ab, 32'h4074c0c2} /* (19, 30, 31) {real, imag} */,
  {32'hbf92ac44, 32'hc013ea78} /* (19, 30, 30) {real, imag} */,
  {32'h3f834024, 32'h3eac8c61} /* (19, 30, 29) {real, imag} */,
  {32'h3ebfce07, 32'hc035740e} /* (19, 30, 28) {real, imag} */,
  {32'hbf87ebb6, 32'h402cfb89} /* (19, 30, 27) {real, imag} */,
  {32'hc0123416, 32'h3fbfd488} /* (19, 30, 26) {real, imag} */,
  {32'hbf7b5cac, 32'h3fd5f7cb} /* (19, 30, 25) {real, imag} */,
  {32'hc051c68a, 32'hc003112c} /* (19, 30, 24) {real, imag} */,
  {32'hbfd22f14, 32'h3f441fbb} /* (19, 30, 23) {real, imag} */,
  {32'hbf332ffd, 32'hbe9f697f} /* (19, 30, 22) {real, imag} */,
  {32'h3e112ffd, 32'hbfcb6f41} /* (19, 30, 21) {real, imag} */,
  {32'hc000e0cb, 32'h40129e02} /* (19, 30, 20) {real, imag} */,
  {32'hbe2669e4, 32'h3ffd7e34} /* (19, 30, 19) {real, imag} */,
  {32'h3f92baef, 32'hc01e400c} /* (19, 30, 18) {real, imag} */,
  {32'h3fe548b6, 32'h3f9f1b56} /* (19, 30, 17) {real, imag} */,
  {32'h3f275e41, 32'hbe1abbdf} /* (19, 30, 16) {real, imag} */,
  {32'hbe82d4d9, 32'h3f3ee339} /* (19, 30, 15) {real, imag} */,
  {32'h400245d6, 32'hbfd3a507} /* (19, 30, 14) {real, imag} */,
  {32'hbf7dc12e, 32'hbf42e472} /* (19, 30, 13) {real, imag} */,
  {32'hbece1432, 32'hbf58010f} /* (19, 30, 12) {real, imag} */,
  {32'hc0224b80, 32'hbf7695e8} /* (19, 30, 11) {real, imag} */,
  {32'hc0174af6, 32'h3f2ed9f9} /* (19, 30, 10) {real, imag} */,
  {32'h3f887a21, 32'hc0227a14} /* (19, 30, 9) {real, imag} */,
  {32'hc00d9236, 32'h4012484c} /* (19, 30, 8) {real, imag} */,
  {32'h3fd767eb, 32'h3f3ff10e} /* (19, 30, 7) {real, imag} */,
  {32'hbea50518, 32'h405c286e} /* (19, 30, 6) {real, imag} */,
  {32'hc025c19d, 32'hbe4812f8} /* (19, 30, 5) {real, imag} */,
  {32'h40213ab3, 32'hbf731676} /* (19, 30, 4) {real, imag} */,
  {32'h40654440, 32'h3f91b5bd} /* (19, 30, 3) {real, imag} */,
  {32'h40189c0d, 32'hc04bf6ac} /* (19, 30, 2) {real, imag} */,
  {32'hbf83cb0c, 32'hbf982026} /* (19, 30, 1) {real, imag} */,
  {32'h40248d38, 32'hbf15ce9b} /* (19, 30, 0) {real, imag} */,
  {32'hbf91de9e, 32'h3f880cc7} /* (19, 29, 31) {real, imag} */,
  {32'hbfb73a16, 32'hbf16494f} /* (19, 29, 30) {real, imag} */,
  {32'hbf74c1cf, 32'h3e0d785c} /* (19, 29, 29) {real, imag} */,
  {32'h3fdc208d, 32'hbf916241} /* (19, 29, 28) {real, imag} */,
  {32'hbf229048, 32'hbf997c0d} /* (19, 29, 27) {real, imag} */,
  {32'hbf0792bd, 32'hbefc7d7f} /* (19, 29, 26) {real, imag} */,
  {32'h3ecb1292, 32'hbfd99de1} /* (19, 29, 25) {real, imag} */,
  {32'hbf27904f, 32'hc0666253} /* (19, 29, 24) {real, imag} */,
  {32'h3ff0ead8, 32'h3f27882d} /* (19, 29, 23) {real, imag} */,
  {32'h3e802b7e, 32'hbfd75631} /* (19, 29, 22) {real, imag} */,
  {32'hbff34ae9, 32'hbeb75671} /* (19, 29, 21) {real, imag} */,
  {32'h3f11e9a7, 32'hbf28ed63} /* (19, 29, 20) {real, imag} */,
  {32'h3f033ab8, 32'hc00c9ee2} /* (19, 29, 19) {real, imag} */,
  {32'hc0415085, 32'h3f381f3b} /* (19, 29, 18) {real, imag} */,
  {32'h3f0e0ac2, 32'h3f1ec444} /* (19, 29, 17) {real, imag} */,
  {32'hbf79d807, 32'h3ebc6559} /* (19, 29, 16) {real, imag} */,
  {32'hbf7842bd, 32'hbdfa5757} /* (19, 29, 15) {real, imag} */,
  {32'hbe9de14b, 32'hbfcbe46f} /* (19, 29, 14) {real, imag} */,
  {32'hbd383792, 32'hbffe2f27} /* (19, 29, 13) {real, imag} */,
  {32'hbfd0fd63, 32'hbf537382} /* (19, 29, 12) {real, imag} */,
  {32'hbe9e3a90, 32'h3e82d19d} /* (19, 29, 11) {real, imag} */,
  {32'h3f38a998, 32'h4016f5e4} /* (19, 29, 10) {real, imag} */,
  {32'h3eea9f93, 32'h3d94841a} /* (19, 29, 9) {real, imag} */,
  {32'hbf36c356, 32'hbc70c214} /* (19, 29, 8) {real, imag} */,
  {32'h3fd9c80c, 32'hbe1b9f5b} /* (19, 29, 7) {real, imag} */,
  {32'hbe5d0b71, 32'hc0316017} /* (19, 29, 6) {real, imag} */,
  {32'hbdcd6359, 32'h3f381db6} /* (19, 29, 5) {real, imag} */,
  {32'h3f5c925f, 32'h3eee4fb1} /* (19, 29, 4) {real, imag} */,
  {32'hbf0c03d6, 32'h402efc89} /* (19, 29, 3) {real, imag} */,
  {32'hbfa1a81d, 32'h3fa79b23} /* (19, 29, 2) {real, imag} */,
  {32'hbf1a7842, 32'hbf097b7d} /* (19, 29, 1) {real, imag} */,
  {32'hbfd84f38, 32'h3c2452e7} /* (19, 29, 0) {real, imag} */,
  {32'h3f2d201d, 32'hbfcacd2e} /* (19, 28, 31) {real, imag} */,
  {32'h3fb1c3c0, 32'h3ded8590} /* (19, 28, 30) {real, imag} */,
  {32'hbe2104a1, 32'hbfb6598e} /* (19, 28, 29) {real, imag} */,
  {32'hc00166fa, 32'hc08efde1} /* (19, 28, 28) {real, imag} */,
  {32'h3de7b84e, 32'h400550d2} /* (19, 28, 27) {real, imag} */,
  {32'hbe50513b, 32'h3f3eefc3} /* (19, 28, 26) {real, imag} */,
  {32'h3f7984fb, 32'h3f4ab943} /* (19, 28, 25) {real, imag} */,
  {32'hbc8c022f, 32'h40268f1a} /* (19, 28, 24) {real, imag} */,
  {32'h3f298d74, 32'h3c9b8c57} /* (19, 28, 23) {real, imag} */,
  {32'hbf918ada, 32'hbfedf3f0} /* (19, 28, 22) {real, imag} */,
  {32'h3e87c2f0, 32'h3fa45970} /* (19, 28, 21) {real, imag} */,
  {32'hbd5cfd2f, 32'h3fa0f563} /* (19, 28, 20) {real, imag} */,
  {32'h400554bb, 32'hbfcb21d8} /* (19, 28, 19) {real, imag} */,
  {32'h3ec0d176, 32'hbf289496} /* (19, 28, 18) {real, imag} */,
  {32'hbe5f330f, 32'hbec80b1b} /* (19, 28, 17) {real, imag} */,
  {32'h3f6e1cd1, 32'hbe9e2942} /* (19, 28, 16) {real, imag} */,
  {32'hbf91525f, 32'hbf796df4} /* (19, 28, 15) {real, imag} */,
  {32'h3e09e542, 32'h4039ad84} /* (19, 28, 14) {real, imag} */,
  {32'h3f68ad1c, 32'h3f3098dc} /* (19, 28, 13) {real, imag} */,
  {32'hbfbb29a3, 32'h3f4b5269} /* (19, 28, 12) {real, imag} */,
  {32'h3eec4060, 32'hbf1a2f4b} /* (19, 28, 11) {real, imag} */,
  {32'h3f237385, 32'h3e9b9326} /* (19, 28, 10) {real, imag} */,
  {32'h3f544f22, 32'h3fe04af2} /* (19, 28, 9) {real, imag} */,
  {32'h3f690ed0, 32'h3f516cb9} /* (19, 28, 8) {real, imag} */,
  {32'h3f389705, 32'h3f4f9e41} /* (19, 28, 7) {real, imag} */,
  {32'hbe122b31, 32'hbface116} /* (19, 28, 6) {real, imag} */,
  {32'hbfd19c68, 32'h3ff28d11} /* (19, 28, 5) {real, imag} */,
  {32'h3fce1d81, 32'h3fd79b52} /* (19, 28, 4) {real, imag} */,
  {32'h3f8bcae2, 32'hbeeff98f} /* (19, 28, 3) {real, imag} */,
  {32'hbfaa2afd, 32'hc0145d43} /* (19, 28, 2) {real, imag} */,
  {32'h3f26cdf2, 32'h3fdce42d} /* (19, 28, 1) {real, imag} */,
  {32'h3f57d80a, 32'h401c6833} /* (19, 28, 0) {real, imag} */,
  {32'hbfab5413, 32'hbfee8417} /* (19, 27, 31) {real, imag} */,
  {32'h3e35d7e1, 32'hc0277c61} /* (19, 27, 30) {real, imag} */,
  {32'h40709f2f, 32'hbecbe447} /* (19, 27, 29) {real, imag} */,
  {32'h3f57beca, 32'hbe086c00} /* (19, 27, 28) {real, imag} */,
  {32'h3e2fa555, 32'hbada68e1} /* (19, 27, 27) {real, imag} */,
  {32'h40b0332c, 32'hbe1601a8} /* (19, 27, 26) {real, imag} */,
  {32'hc08cda59, 32'h40188e12} /* (19, 27, 25) {real, imag} */,
  {32'h40301ed7, 32'h3f8d2f6d} /* (19, 27, 24) {real, imag} */,
  {32'hbfd8c696, 32'hbe8904c4} /* (19, 27, 23) {real, imag} */,
  {32'hbf7aa3bb, 32'h3ec8e78b} /* (19, 27, 22) {real, imag} */,
  {32'hc0714c9d, 32'h3fc55bfe} /* (19, 27, 21) {real, imag} */,
  {32'hbfbd67a4, 32'h3fe0064d} /* (19, 27, 20) {real, imag} */,
  {32'h3f03c398, 32'h3f30870d} /* (19, 27, 19) {real, imag} */,
  {32'h40025853, 32'h3d92e46e} /* (19, 27, 18) {real, imag} */,
  {32'h3e5f6051, 32'hbf9f9914} /* (19, 27, 17) {real, imag} */,
  {32'h3fe8e2ab, 32'hbf18c676} /* (19, 27, 16) {real, imag} */,
  {32'hbf991ebf, 32'hbf3a9619} /* (19, 27, 15) {real, imag} */,
  {32'hbeea2f3e, 32'h3ee9ae43} /* (19, 27, 14) {real, imag} */,
  {32'hc0085a9a, 32'h3f201f61} /* (19, 27, 13) {real, imag} */,
  {32'hbeff8c18, 32'h3fa49b34} /* (19, 27, 12) {real, imag} */,
  {32'hc073f807, 32'hc00a7406} /* (19, 27, 11) {real, imag} */,
  {32'hc06e59a6, 32'h403cff64} /* (19, 27, 10) {real, imag} */,
  {32'h3d411437, 32'hbf45ea5e} /* (19, 27, 9) {real, imag} */,
  {32'hc00c1fa3, 32'hbfebe8ea} /* (19, 27, 8) {real, imag} */,
  {32'hbfd8ad18, 32'h3f6db43e} /* (19, 27, 7) {real, imag} */,
  {32'h3db14a91, 32'hbf4bc184} /* (19, 27, 6) {real, imag} */,
  {32'hbf827f03, 32'hbddc344f} /* (19, 27, 5) {real, imag} */,
  {32'hbf8b7d65, 32'hbfba37ed} /* (19, 27, 4) {real, imag} */,
  {32'hbf5ed454, 32'h3fe24350} /* (19, 27, 3) {real, imag} */,
  {32'h3fc425dd, 32'h4000a02c} /* (19, 27, 2) {real, imag} */,
  {32'h3e9df34d, 32'h3fc79c9a} /* (19, 27, 1) {real, imag} */,
  {32'h401307d8, 32'h3f28c4b8} /* (19, 27, 0) {real, imag} */,
  {32'h3dd11308, 32'h3ef2c552} /* (19, 26, 31) {real, imag} */,
  {32'h4048ba89, 32'h3fcf02d7} /* (19, 26, 30) {real, imag} */,
  {32'hbfcf8705, 32'h3e4bf5e2} /* (19, 26, 29) {real, imag} */,
  {32'hbfc0af12, 32'h3ee594c9} /* (19, 26, 28) {real, imag} */,
  {32'h402dd21b, 32'hbeb99221} /* (19, 26, 27) {real, imag} */,
  {32'h3fb16526, 32'hc042d155} /* (19, 26, 26) {real, imag} */,
  {32'hbf1b1131, 32'hbff58259} /* (19, 26, 25) {real, imag} */,
  {32'hc0123c29, 32'h3f8ca6dc} /* (19, 26, 24) {real, imag} */,
  {32'h3fec594e, 32'h3fd68576} /* (19, 26, 23) {real, imag} */,
  {32'hbf62d741, 32'h40056fbd} /* (19, 26, 22) {real, imag} */,
  {32'hbfe25e40, 32'hc01477e1} /* (19, 26, 21) {real, imag} */,
  {32'h3f2f94bc, 32'h3f5df98c} /* (19, 26, 20) {real, imag} */,
  {32'h3f95c385, 32'hbf2d2c32} /* (19, 26, 19) {real, imag} */,
  {32'h4002352a, 32'hbde82ff1} /* (19, 26, 18) {real, imag} */,
  {32'hc00b16b2, 32'h404346ca} /* (19, 26, 17) {real, imag} */,
  {32'hbf27fd27, 32'hbebc62a3} /* (19, 26, 16) {real, imag} */,
  {32'hbff1f211, 32'hbe946595} /* (19, 26, 15) {real, imag} */,
  {32'h3fd44997, 32'h3fcf8dc3} /* (19, 26, 14) {real, imag} */,
  {32'h4007ab9c, 32'hc08b60be} /* (19, 26, 13) {real, imag} */,
  {32'hbe5bf036, 32'h3e4ae801} /* (19, 26, 12) {real, imag} */,
  {32'h3f129ffd, 32'hbf24134a} /* (19, 26, 11) {real, imag} */,
  {32'hbf504b96, 32'hbd9e6e5c} /* (19, 26, 10) {real, imag} */,
  {32'h401ac73a, 32'h401786f6} /* (19, 26, 9) {real, imag} */,
  {32'hc02cadfe, 32'h40b56797} /* (19, 26, 8) {real, imag} */,
  {32'hbedb604c, 32'hbfb0d238} /* (19, 26, 7) {real, imag} */,
  {32'hbfb1ac2d, 32'h40252143} /* (19, 26, 6) {real, imag} */,
  {32'h3f4a48bb, 32'h3feca2cc} /* (19, 26, 5) {real, imag} */,
  {32'hbf447f03, 32'hbfe5a1b6} /* (19, 26, 4) {real, imag} */,
  {32'h3f285495, 32'h3f879f68} /* (19, 26, 3) {real, imag} */,
  {32'hbfb8e03a, 32'hc01a8681} /* (19, 26, 2) {real, imag} */,
  {32'hc00d90d1, 32'hbf2fa8e4} /* (19, 26, 1) {real, imag} */,
  {32'h3f972bce, 32'hbf977ee5} /* (19, 26, 0) {real, imag} */,
  {32'h400a54cf, 32'hbf4f8662} /* (19, 25, 31) {real, imag} */,
  {32'hc05606da, 32'hbf906d0e} /* (19, 25, 30) {real, imag} */,
  {32'hbf2931b7, 32'hbea7d3be} /* (19, 25, 29) {real, imag} */,
  {32'h3f19002d, 32'h3ed8e2b8} /* (19, 25, 28) {real, imag} */,
  {32'hbe7a7918, 32'hc02f817a} /* (19, 25, 27) {real, imag} */,
  {32'h3f13642a, 32'hbf93ec52} /* (19, 25, 26) {real, imag} */,
  {32'h405845a3, 32'h408696dc} /* (19, 25, 25) {real, imag} */,
  {32'hbe8bfc60, 32'h3fe4aef6} /* (19, 25, 24) {real, imag} */,
  {32'hbd9345c3, 32'hc081cc57} /* (19, 25, 23) {real, imag} */,
  {32'hbf29e6fb, 32'hc0016ce5} /* (19, 25, 22) {real, imag} */,
  {32'hbfa43007, 32'h40347249} /* (19, 25, 21) {real, imag} */,
  {32'h3f8ac1fd, 32'hbf94f8e2} /* (19, 25, 20) {real, imag} */,
  {32'h3e4c8573, 32'hbee9d413} /* (19, 25, 19) {real, imag} */,
  {32'h3f13cd23, 32'h4016f46f} /* (19, 25, 18) {real, imag} */,
  {32'h3eaf7b10, 32'hbef59fcb} /* (19, 25, 17) {real, imag} */,
  {32'h40021f9d, 32'hbfa05372} /* (19, 25, 16) {real, imag} */,
  {32'hbe0e2f76, 32'h3ca7175c} /* (19, 25, 15) {real, imag} */,
  {32'h3fb052eb, 32'h3f81482b} /* (19, 25, 14) {real, imag} */,
  {32'hc043bc1e, 32'h3dbdb9da} /* (19, 25, 13) {real, imag} */,
  {32'hc000da1a, 32'hbe83a415} /* (19, 25, 12) {real, imag} */,
  {32'h4038e56c, 32'hc00e3212} /* (19, 25, 11) {real, imag} */,
  {32'h3f89e65d, 32'h3f98b75d} /* (19, 25, 10) {real, imag} */,
  {32'hbf125002, 32'h3fac41c1} /* (19, 25, 9) {real, imag} */,
  {32'hbdd8dcdf, 32'hbf1f21ba} /* (19, 25, 8) {real, imag} */,
  {32'hbfedbb0d, 32'hbf3c2eb9} /* (19, 25, 7) {real, imag} */,
  {32'hbc13e87f, 32'h3fe4dba6} /* (19, 25, 6) {real, imag} */,
  {32'hbfeb69ae, 32'h3f78da98} /* (19, 25, 5) {real, imag} */,
  {32'h3f22ca7a, 32'h3f44dbfb} /* (19, 25, 4) {real, imag} */,
  {32'hbf3d6d43, 32'h3daa6315} /* (19, 25, 3) {real, imag} */,
  {32'hbed2b684, 32'h3f99179d} /* (19, 25, 2) {real, imag} */,
  {32'h3f9a0939, 32'h3f6796dc} /* (19, 25, 1) {real, imag} */,
  {32'hc018a51c, 32'h3f7eb79b} /* (19, 25, 0) {real, imag} */,
  {32'h3eabf47a, 32'h3d95bdd2} /* (19, 24, 31) {real, imag} */,
  {32'h3e6c0c4a, 32'h40059c9b} /* (19, 24, 30) {real, imag} */,
  {32'hc04fa65d, 32'hbf612851} /* (19, 24, 29) {real, imag} */,
  {32'hbbb96907, 32'hc01a7133} /* (19, 24, 28) {real, imag} */,
  {32'hbfba8927, 32'hbfe2b499} /* (19, 24, 27) {real, imag} */,
  {32'hbfacf580, 32'h3f78c3cc} /* (19, 24, 26) {real, imag} */,
  {32'hbec28b77, 32'h3e539820} /* (19, 24, 25) {real, imag} */,
  {32'h3d884931, 32'h3fdbb3f4} /* (19, 24, 24) {real, imag} */,
  {32'hbfc4cc84, 32'hbfe75624} /* (19, 24, 23) {real, imag} */,
  {32'h402c9384, 32'h405734ca} /* (19, 24, 22) {real, imag} */,
  {32'hbe9bbfee, 32'h402c6f11} /* (19, 24, 21) {real, imag} */,
  {32'h3ec371d0, 32'hc0152cab} /* (19, 24, 20) {real, imag} */,
  {32'hbfa386d9, 32'hc0158260} /* (19, 24, 19) {real, imag} */,
  {32'hbff649b4, 32'h3fa755e2} /* (19, 24, 18) {real, imag} */,
  {32'h3f31f6e7, 32'hbf30bda6} /* (19, 24, 17) {real, imag} */,
  {32'h3c80a0fb, 32'hbcc4e8c1} /* (19, 24, 16) {real, imag} */,
  {32'hbe998c83, 32'h3fa9ea8d} /* (19, 24, 15) {real, imag} */,
  {32'h3e910145, 32'hbe9953bb} /* (19, 24, 14) {real, imag} */,
  {32'hbfcaae43, 32'h402671da} /* (19, 24, 13) {real, imag} */,
  {32'h3de33229, 32'hc0112e18} /* (19, 24, 12) {real, imag} */,
  {32'hc05d2f68, 32'hbf46b1e7} /* (19, 24, 11) {real, imag} */,
  {32'h3f744da6, 32'hbfa25abe} /* (19, 24, 10) {real, imag} */,
  {32'h3f0b8017, 32'h406bbd88} /* (19, 24, 9) {real, imag} */,
  {32'h3f05ab6a, 32'h3ea51bca} /* (19, 24, 8) {real, imag} */,
  {32'hbf85a304, 32'hbf507ae3} /* (19, 24, 7) {real, imag} */,
  {32'h4032897b, 32'h3f9f025d} /* (19, 24, 6) {real, imag} */,
  {32'h3f62a1fd, 32'hbee5f01d} /* (19, 24, 5) {real, imag} */,
  {32'h400d5161, 32'h40021caf} /* (19, 24, 4) {real, imag} */,
  {32'h403c77c9, 32'h40207ec1} /* (19, 24, 3) {real, imag} */,
  {32'hc02afbc6, 32'hbf95d4ea} /* (19, 24, 2) {real, imag} */,
  {32'h40022526, 32'h3f0b90c0} /* (19, 24, 1) {real, imag} */,
  {32'h40254c0a, 32'h3f9adad2} /* (19, 24, 0) {real, imag} */,
  {32'h402ae57e, 32'h3ed2c271} /* (19, 23, 31) {real, imag} */,
  {32'hc0258bf0, 32'h3eb08897} /* (19, 23, 30) {real, imag} */,
  {32'hbfe72e27, 32'h3fb88718} /* (19, 23, 29) {real, imag} */,
  {32'h3eb3cbdc, 32'h3f5c279b} /* (19, 23, 28) {real, imag} */,
  {32'hc044201a, 32'hc00f5374} /* (19, 23, 27) {real, imag} */,
  {32'hc00cd02f, 32'hbf9c877f} /* (19, 23, 26) {real, imag} */,
  {32'hbf8a5d6a, 32'hbf22cfaf} /* (19, 23, 25) {real, imag} */,
  {32'h40339858, 32'hbf92f4c2} /* (19, 23, 24) {real, imag} */,
  {32'h40451674, 32'h3dfd8d80} /* (19, 23, 23) {real, imag} */,
  {32'hc02b8a45, 32'hbd91c9d6} /* (19, 23, 22) {real, imag} */,
  {32'h3f24d7bc, 32'h3ee65785} /* (19, 23, 21) {real, imag} */,
  {32'hbd36ed29, 32'h400cdf11} /* (19, 23, 20) {real, imag} */,
  {32'hbe5e3601, 32'h3eb5a0eb} /* (19, 23, 19) {real, imag} */,
  {32'hbfbd9904, 32'h3f878673} /* (19, 23, 18) {real, imag} */,
  {32'h3fad855a, 32'hc000a674} /* (19, 23, 17) {real, imag} */,
  {32'h3f1c2661, 32'h3f678fd9} /* (19, 23, 16) {real, imag} */,
  {32'hbf00d6e3, 32'hbfe70ca6} /* (19, 23, 15) {real, imag} */,
  {32'hc0347085, 32'hbeb69091} /* (19, 23, 14) {real, imag} */,
  {32'hbf1a9bd0, 32'hbf10eb1a} /* (19, 23, 13) {real, imag} */,
  {32'h3f3b4ada, 32'h40b97782} /* (19, 23, 12) {real, imag} */,
  {32'h4089b701, 32'h3f847c62} /* (19, 23, 11) {real, imag} */,
  {32'h3fd48a44, 32'hc03af0ea} /* (19, 23, 10) {real, imag} */,
  {32'h3fe4ece5, 32'h40512c40} /* (19, 23, 9) {real, imag} */,
  {32'h3f031fe9, 32'h40820a6e} /* (19, 23, 8) {real, imag} */,
  {32'hbf621b8d, 32'h3fda0bbb} /* (19, 23, 7) {real, imag} */,
  {32'hc05e5538, 32'hbfe94258} /* (19, 23, 6) {real, imag} */,
  {32'h3e3b2643, 32'hc0054ae6} /* (19, 23, 5) {real, imag} */,
  {32'hbfc0f4d0, 32'hbfa459cc} /* (19, 23, 4) {real, imag} */,
  {32'hbe1f37ed, 32'hc0982a76} /* (19, 23, 3) {real, imag} */,
  {32'h3ebb4c94, 32'h3fddb6fe} /* (19, 23, 2) {real, imag} */,
  {32'hc0060f5b, 32'h40704b5c} /* (19, 23, 1) {real, imag} */,
  {32'hbfaa57ec, 32'hbe88b47a} /* (19, 23, 0) {real, imag} */,
  {32'hbf4af6e6, 32'h3f59c725} /* (19, 22, 31) {real, imag} */,
  {32'hbfbf7c0d, 32'hbfd81d65} /* (19, 22, 30) {real, imag} */,
  {32'h3fbd2040, 32'h3cdea7cc} /* (19, 22, 29) {real, imag} */,
  {32'hbf95b8e1, 32'h407d2e5e} /* (19, 22, 28) {real, imag} */,
  {32'hbea43f6b, 32'hc0633d74} /* (19, 22, 27) {real, imag} */,
  {32'hbf54e5a4, 32'hc04a9e3c} /* (19, 22, 26) {real, imag} */,
  {32'h3fcdbe99, 32'h3f8a217a} /* (19, 22, 25) {real, imag} */,
  {32'h3fec8ba9, 32'hbf922d42} /* (19, 22, 24) {real, imag} */,
  {32'hbffc29a3, 32'h3ffebd03} /* (19, 22, 23) {real, imag} */,
  {32'h3e2bfcdd, 32'h3f5f0040} /* (19, 22, 22) {real, imag} */,
  {32'h3fc231a1, 32'h3de19939} /* (19, 22, 21) {real, imag} */,
  {32'hc06f36cd, 32'h3f699f52} /* (19, 22, 20) {real, imag} */,
  {32'h404d7484, 32'h3fcf4732} /* (19, 22, 19) {real, imag} */,
  {32'hbfcd52ce, 32'h3e4b3c1e} /* (19, 22, 18) {real, imag} */,
  {32'hbeef3738, 32'hbebefdfd} /* (19, 22, 17) {real, imag} */,
  {32'h400d7380, 32'h3f24fc67} /* (19, 22, 16) {real, imag} */,
  {32'hbea42b22, 32'h4021c2ee} /* (19, 22, 15) {real, imag} */,
  {32'hbf4660ce, 32'hc00c9df1} /* (19, 22, 14) {real, imag} */,
  {32'h3ffb0c36, 32'h403de546} /* (19, 22, 13) {real, imag} */,
  {32'h3f1f362d, 32'hc0562599} /* (19, 22, 12) {real, imag} */,
  {32'h3fc85fa8, 32'hc094cd68} /* (19, 22, 11) {real, imag} */,
  {32'hbf53e341, 32'h402a7d53} /* (19, 22, 10) {real, imag} */,
  {32'h3f53728b, 32'h400ca96d} /* (19, 22, 9) {real, imag} */,
  {32'h3f1d94f2, 32'h403549df} /* (19, 22, 8) {real, imag} */,
  {32'h3fff0210, 32'hbf4df922} /* (19, 22, 7) {real, imag} */,
  {32'h3e3925a8, 32'hbf940af7} /* (19, 22, 6) {real, imag} */,
  {32'h408d6831, 32'h3f26396e} /* (19, 22, 5) {real, imag} */,
  {32'hc0997d10, 32'h3feaccb9} /* (19, 22, 4) {real, imag} */,
  {32'hc00193c1, 32'h3ec1d886} /* (19, 22, 3) {real, imag} */,
  {32'hc00f549b, 32'hbe180029} /* (19, 22, 2) {real, imag} */,
  {32'h3fd5df99, 32'hbfd7784c} /* (19, 22, 1) {real, imag} */,
  {32'h3fb4f637, 32'h404e2337} /* (19, 22, 0) {real, imag} */,
  {32'hbe7d1e0c, 32'h4030e11e} /* (19, 21, 31) {real, imag} */,
  {32'h3f61d6c5, 32'hbf860ac2} /* (19, 21, 30) {real, imag} */,
  {32'h4028502b, 32'h4015a05c} /* (19, 21, 29) {real, imag} */,
  {32'hbf043c7b, 32'hbe640b7a} /* (19, 21, 28) {real, imag} */,
  {32'hc08e8da5, 32'hbf68d3a1} /* (19, 21, 27) {real, imag} */,
  {32'hc0946d3b, 32'hbed970a0} /* (19, 21, 26) {real, imag} */,
  {32'h3d4dafc1, 32'hbf4a0d2a} /* (19, 21, 25) {real, imag} */,
  {32'hbfcc70b4, 32'h403c162c} /* (19, 21, 24) {real, imag} */,
  {32'hbf9f0cb6, 32'hc02819d8} /* (19, 21, 23) {real, imag} */,
  {32'hbe672b65, 32'hbfc046f8} /* (19, 21, 22) {real, imag} */,
  {32'h40235a64, 32'h4070dcb5} /* (19, 21, 21) {real, imag} */,
  {32'h3fa7d286, 32'hc02703d1} /* (19, 21, 20) {real, imag} */,
  {32'h3fd50e94, 32'hbebc220e} /* (19, 21, 19) {real, imag} */,
  {32'h3f0d85b0, 32'hbf0b2515} /* (19, 21, 18) {real, imag} */,
  {32'hbf737054, 32'h3f816476} /* (19, 21, 17) {real, imag} */,
  {32'hbf85087e, 32'hbf252377} /* (19, 21, 16) {real, imag} */,
  {32'h3fe6c289, 32'h3fcf8b69} /* (19, 21, 15) {real, imag} */,
  {32'h402a3b6d, 32'hbf86985a} /* (19, 21, 14) {real, imag} */,
  {32'h3de559ad, 32'hbfb158e9} /* (19, 21, 13) {real, imag} */,
  {32'h404645ec, 32'hbdcf8046} /* (19, 21, 12) {real, imag} */,
  {32'hc0259ab9, 32'h3e8dbd41} /* (19, 21, 11) {real, imag} */,
  {32'hc01b1335, 32'h3fccee60} /* (19, 21, 10) {real, imag} */,
  {32'hc0bb86a6, 32'hbebf3d3e} /* (19, 21, 9) {real, imag} */,
  {32'hbf7c3765, 32'hbe875ea7} /* (19, 21, 8) {real, imag} */,
  {32'hc00225d9, 32'h40040c5b} /* (19, 21, 7) {real, imag} */,
  {32'h3f2fde4e, 32'hbf6815b6} /* (19, 21, 6) {real, imag} */,
  {32'h3f704311, 32'hbc9ccfcd} /* (19, 21, 5) {real, imag} */,
  {32'h3f281d7f, 32'h3f0795e9} /* (19, 21, 4) {real, imag} */,
  {32'hbf489c71, 32'hbf234598} /* (19, 21, 3) {real, imag} */,
  {32'h3f2db778, 32'h3f64d3fe} /* (19, 21, 2) {real, imag} */,
  {32'h3ee19ea7, 32'hbec691a5} /* (19, 21, 1) {real, imag} */,
  {32'hbf2b8aae, 32'hbf9fe013} /* (19, 21, 0) {real, imag} */,
  {32'h401b7dfa, 32'hbfadb0ef} /* (19, 20, 31) {real, imag} */,
  {32'h3fc927fa, 32'h3f2fe65a} /* (19, 20, 30) {real, imag} */,
  {32'h3e9df65a, 32'h40760909} /* (19, 20, 29) {real, imag} */,
  {32'hc0623927, 32'hbf570449} /* (19, 20, 28) {real, imag} */,
  {32'hbf84deee, 32'hbe229aa6} /* (19, 20, 27) {real, imag} */,
  {32'hbeb0fa30, 32'hbea41465} /* (19, 20, 26) {real, imag} */,
  {32'h3fae155b, 32'hbe8e1909} /* (19, 20, 25) {real, imag} */,
  {32'hbee2a07b, 32'h3fff0568} /* (19, 20, 24) {real, imag} */,
  {32'hbe583f65, 32'hbe4a2231} /* (19, 20, 23) {real, imag} */,
  {32'hbedaa8e8, 32'hbea37902} /* (19, 20, 22) {real, imag} */,
  {32'h404c7f5b, 32'h3f13a5e0} /* (19, 20, 21) {real, imag} */,
  {32'h40552f89, 32'hbf487b8e} /* (19, 20, 20) {real, imag} */,
  {32'hbfa76d94, 32'h3f4e547a} /* (19, 20, 19) {real, imag} */,
  {32'h3f8d457d, 32'hbe09753e} /* (19, 20, 18) {real, imag} */,
  {32'h3f8bf1b8, 32'h406eea54} /* (19, 20, 17) {real, imag} */,
  {32'hbf00a307, 32'hbf762eb9} /* (19, 20, 16) {real, imag} */,
  {32'h3f7b5c52, 32'hbff01bca} /* (19, 20, 15) {real, imag} */,
  {32'hbfdb175d, 32'hbfa34eea} /* (19, 20, 14) {real, imag} */,
  {32'hbea9a16c, 32'h3fdeeb59} /* (19, 20, 13) {real, imag} */,
  {32'h3fb0b3ef, 32'hbf470bda} /* (19, 20, 12) {real, imag} */,
  {32'h402ca14e, 32'h40115f64} /* (19, 20, 11) {real, imag} */,
  {32'h3ffad3c9, 32'hbe59c2a9} /* (19, 20, 10) {real, imag} */,
  {32'h3fef5214, 32'hbc081609} /* (19, 20, 9) {real, imag} */,
  {32'hbfe53bdd, 32'h3de56009} /* (19, 20, 8) {real, imag} */,
  {32'h408bc49c, 32'h3e6e3f76} /* (19, 20, 7) {real, imag} */,
  {32'hc049b980, 32'hbe84cbdb} /* (19, 20, 6) {real, imag} */,
  {32'h3f751ad7, 32'hbffa035f} /* (19, 20, 5) {real, imag} */,
  {32'h3f71683f, 32'h3f1a72a3} /* (19, 20, 4) {real, imag} */,
  {32'h3e3a74c8, 32'h3f15cbe3} /* (19, 20, 3) {real, imag} */,
  {32'hbfe8bc01, 32'hbf736ed4} /* (19, 20, 2) {real, imag} */,
  {32'h3df9ce5f, 32'h3ecef558} /* (19, 20, 1) {real, imag} */,
  {32'hbfbfe181, 32'hbf969a3a} /* (19, 20, 0) {real, imag} */,
  {32'h3fd97e4e, 32'hbe08820d} /* (19, 19, 31) {real, imag} */,
  {32'h3fadc6f4, 32'h3fc7b3ec} /* (19, 19, 30) {real, imag} */,
  {32'h3f80efc8, 32'hbf0dcac4} /* (19, 19, 29) {real, imag} */,
  {32'h3e9e5014, 32'h3fb84e8d} /* (19, 19, 28) {real, imag} */,
  {32'h3fb4a374, 32'hbfc436bc} /* (19, 19, 27) {real, imag} */,
  {32'h4074bc1c, 32'h400d7979} /* (19, 19, 26) {real, imag} */,
  {32'h3f602965, 32'hc003fb9f} /* (19, 19, 25) {real, imag} */,
  {32'hc03df95f, 32'h3fae26e4} /* (19, 19, 24) {real, imag} */,
  {32'hbfe8f661, 32'h3ddeffdc} /* (19, 19, 23) {real, imag} */,
  {32'h3f936d78, 32'h3f048822} /* (19, 19, 22) {real, imag} */,
  {32'hc0164bf9, 32'h3e80efa1} /* (19, 19, 21) {real, imag} */,
  {32'hbea4e538, 32'hbf96091e} /* (19, 19, 20) {real, imag} */,
  {32'h4065a4eb, 32'h3dc3b4ed} /* (19, 19, 19) {real, imag} */,
  {32'hbfb03540, 32'h3ffe24bb} /* (19, 19, 18) {real, imag} */,
  {32'hbfb9a974, 32'hc00c8f15} /* (19, 19, 17) {real, imag} */,
  {32'h3fa10963, 32'h3fedd0f6} /* (19, 19, 16) {real, imag} */,
  {32'hbed82108, 32'h3e749a28} /* (19, 19, 15) {real, imag} */,
  {32'hbf2d29af, 32'h3f601dec} /* (19, 19, 14) {real, imag} */,
  {32'hbfde6fce, 32'h3f90b982} /* (19, 19, 13) {real, imag} */,
  {32'h3f50847b, 32'h4001b31c} /* (19, 19, 12) {real, imag} */,
  {32'hbfa314b3, 32'hc00993b6} /* (19, 19, 11) {real, imag} */,
  {32'hbfa31857, 32'hc00e8f7d} /* (19, 19, 10) {real, imag} */,
  {32'hc0467609, 32'h3fc82641} /* (19, 19, 9) {real, imag} */,
  {32'h4024f532, 32'hbfe2133d} /* (19, 19, 8) {real, imag} */,
  {32'hbf553842, 32'h3fbb4369} /* (19, 19, 7) {real, imag} */,
  {32'h3f4a93e5, 32'hc0315689} /* (19, 19, 6) {real, imag} */,
  {32'h3dde66eb, 32'h404ace5c} /* (19, 19, 5) {real, imag} */,
  {32'hbfd9f33b, 32'h3f9e772f} /* (19, 19, 4) {real, imag} */,
  {32'hc033113e, 32'h402b0751} /* (19, 19, 3) {real, imag} */,
  {32'h401f3a67, 32'hbe862cb9} /* (19, 19, 2) {real, imag} */,
  {32'hbfe1c129, 32'hbfbf4de9} /* (19, 19, 1) {real, imag} */,
  {32'hc0074a2b, 32'h3fac5356} /* (19, 19, 0) {real, imag} */,
  {32'hbd977fe2, 32'hbfba3804} /* (19, 18, 31) {real, imag} */,
  {32'hbf7b1a8c, 32'hbe88a067} /* (19, 18, 30) {real, imag} */,
  {32'h3f3f06af, 32'h3f498a12} /* (19, 18, 29) {real, imag} */,
  {32'hbf882183, 32'h3f449f52} /* (19, 18, 28) {real, imag} */,
  {32'h3f883a57, 32'h3eadb709} /* (19, 18, 27) {real, imag} */,
  {32'h3efc260b, 32'h3f2293b1} /* (19, 18, 26) {real, imag} */,
  {32'h3f2baa71, 32'h3f813474} /* (19, 18, 25) {real, imag} */,
  {32'h3ff87ec6, 32'h3fe8c47a} /* (19, 18, 24) {real, imag} */,
  {32'hbf59376c, 32'hbf3626dd} /* (19, 18, 23) {real, imag} */,
  {32'hbfe6239c, 32'h3f43f5ce} /* (19, 18, 22) {real, imag} */,
  {32'h3feb6b28, 32'hbfafd231} /* (19, 18, 21) {real, imag} */,
  {32'h3ecec165, 32'h3fa2ea9a} /* (19, 18, 20) {real, imag} */,
  {32'hbe3d624e, 32'h4013b136} /* (19, 18, 19) {real, imag} */,
  {32'h3f1ea056, 32'hbfd4be8c} /* (19, 18, 18) {real, imag} */,
  {32'hbdf5c81d, 32'h3f49a37f} /* (19, 18, 17) {real, imag} */,
  {32'h3f56e660, 32'hbff3598d} /* (19, 18, 16) {real, imag} */,
  {32'h3ea8f39e, 32'h3f5c4203} /* (19, 18, 15) {real, imag} */,
  {32'hbd8637b3, 32'hbd72a82e} /* (19, 18, 14) {real, imag} */,
  {32'hc02677ae, 32'h3f312a25} /* (19, 18, 13) {real, imag} */,
  {32'h3f9a852d, 32'h3fc5c3a6} /* (19, 18, 12) {real, imag} */,
  {32'h3fac868e, 32'h4017b78d} /* (19, 18, 11) {real, imag} */,
  {32'h3fbd116e, 32'h3eebf94a} /* (19, 18, 10) {real, imag} */,
  {32'h400901e3, 32'hbfc06b3b} /* (19, 18, 9) {real, imag} */,
  {32'hbe35a9ac, 32'hbeafb979} /* (19, 18, 8) {real, imag} */,
  {32'hbd5bf6e9, 32'h3fcc26c5} /* (19, 18, 7) {real, imag} */,
  {32'hbe09f012, 32'hbff0a386} /* (19, 18, 6) {real, imag} */,
  {32'hbf9fd329, 32'h3d54d256} /* (19, 18, 5) {real, imag} */,
  {32'hbf963353, 32'h3d54ea70} /* (19, 18, 4) {real, imag} */,
  {32'h3fff4a89, 32'hbfb42bb6} /* (19, 18, 3) {real, imag} */,
  {32'h3f6353d8, 32'h401740c0} /* (19, 18, 2) {real, imag} */,
  {32'hbff3e427, 32'hbe947c78} /* (19, 18, 1) {real, imag} */,
  {32'h3fe2d336, 32'h3fd7f5dd} /* (19, 18, 0) {real, imag} */,
  {32'hbf80db8b, 32'h3f4745ab} /* (19, 17, 31) {real, imag} */,
  {32'hbdbeca8f, 32'h3fc103fd} /* (19, 17, 30) {real, imag} */,
  {32'hbfd27acd, 32'hbfe5f0c9} /* (19, 17, 29) {real, imag} */,
  {32'h3fd022c6, 32'hbf39e560} /* (19, 17, 28) {real, imag} */,
  {32'h3fc2c4ee, 32'h3f9d03ff} /* (19, 17, 27) {real, imag} */,
  {32'hbfa6db22, 32'hbf880834} /* (19, 17, 26) {real, imag} */,
  {32'hbfcac17a, 32'h3fc1bb31} /* (19, 17, 25) {real, imag} */,
  {32'h3e89d2f3, 32'hbda0d87f} /* (19, 17, 24) {real, imag} */,
  {32'hc037dd7f, 32'h3f56c9bd} /* (19, 17, 23) {real, imag} */,
  {32'h3ff0f5ba, 32'hbf1d9928} /* (19, 17, 22) {real, imag} */,
  {32'h3fa0f7f3, 32'hc0305a14} /* (19, 17, 21) {real, imag} */,
  {32'h3f874344, 32'hbf885b96} /* (19, 17, 20) {real, imag} */,
  {32'hbedf579c, 32'hbfba6c64} /* (19, 17, 19) {real, imag} */,
  {32'h3fac567d, 32'h3f2e8b4a} /* (19, 17, 18) {real, imag} */,
  {32'hbf94466c, 32'h40263210} /* (19, 17, 17) {real, imag} */,
  {32'h3fbd2dce, 32'h3f4f5cbc} /* (19, 17, 16) {real, imag} */,
  {32'h3f028724, 32'hbfb1db63} /* (19, 17, 15) {real, imag} */,
  {32'hbf5c2129, 32'hbe649832} /* (19, 17, 14) {real, imag} */,
  {32'h3ee6e1e4, 32'hbfb0f647} /* (19, 17, 13) {real, imag} */,
  {32'hc008e09c, 32'hbfb9ae5a} /* (19, 17, 12) {real, imag} */,
  {32'h3f6c1846, 32'hbf8e3129} /* (19, 17, 11) {real, imag} */,
  {32'hbfb6bf5e, 32'hbe7b4f0e} /* (19, 17, 10) {real, imag} */,
  {32'hbca6ca54, 32'hbdc7d157} /* (19, 17, 9) {real, imag} */,
  {32'h3f5465dc, 32'hbf231496} /* (19, 17, 8) {real, imag} */,
  {32'hbef0a80a, 32'hbf871cea} /* (19, 17, 7) {real, imag} */,
  {32'hbf18a1de, 32'h3f3dcf7e} /* (19, 17, 6) {real, imag} */,
  {32'h3f7eb95d, 32'hbee6d227} /* (19, 17, 5) {real, imag} */,
  {32'h400a8685, 32'h3e01a3e7} /* (19, 17, 4) {real, imag} */,
  {32'h3f58ed2a, 32'hbefaddba} /* (19, 17, 3) {real, imag} */,
  {32'h3da8a69a, 32'h3df73aaa} /* (19, 17, 2) {real, imag} */,
  {32'hbf9854c8, 32'h3f43a710} /* (19, 17, 1) {real, imag} */,
  {32'h3ffc6568, 32'h3ebaed0b} /* (19, 17, 0) {real, imag} */,
  {32'hbf6ff833, 32'hbeecdc92} /* (19, 16, 31) {real, imag} */,
  {32'h4003dc6c, 32'h3fc2f38c} /* (19, 16, 30) {real, imag} */,
  {32'h3e554fb9, 32'h3f42fe85} /* (19, 16, 29) {real, imag} */,
  {32'hbe3ddd05, 32'h3f8b9da8} /* (19, 16, 28) {real, imag} */,
  {32'h3d9fa8f6, 32'h3fd47da6} /* (19, 16, 27) {real, imag} */,
  {32'h3f1dd661, 32'h3fb7864f} /* (19, 16, 26) {real, imag} */,
  {32'hbf1c8f39, 32'hbff7e58f} /* (19, 16, 25) {real, imag} */,
  {32'hbe8447c4, 32'hbec05fd9} /* (19, 16, 24) {real, imag} */,
  {32'h4020162c, 32'hbf914218} /* (19, 16, 23) {real, imag} */,
  {32'hbf0d57c0, 32'h3f76732d} /* (19, 16, 22) {real, imag} */,
  {32'hbee026f1, 32'h40029e39} /* (19, 16, 21) {real, imag} */,
  {32'hc010e3fb, 32'hbdd69703} /* (19, 16, 20) {real, imag} */,
  {32'hbfce3366, 32'hbd3ee92f} /* (19, 16, 19) {real, imag} */,
  {32'hbf8d6e5a, 32'hbefe03c4} /* (19, 16, 18) {real, imag} */,
  {32'h3f1b60f5, 32'h3f166301} /* (19, 16, 17) {real, imag} */,
  {32'hbf20bb1f, 32'h3f9a96fe} /* (19, 16, 16) {real, imag} */,
  {32'hbe0791e9, 32'h3f1b8bd0} /* (19, 16, 15) {real, imag} */,
  {32'hbc253161, 32'hc0577551} /* (19, 16, 14) {real, imag} */,
  {32'h40085193, 32'hbf7956e4} /* (19, 16, 13) {real, imag} */,
  {32'h3ee3fb54, 32'hbe5af1d4} /* (19, 16, 12) {real, imag} */,
  {32'h4008460d, 32'h3f31ba2e} /* (19, 16, 11) {real, imag} */,
  {32'hbfc34321, 32'h400f59ac} /* (19, 16, 10) {real, imag} */,
  {32'hbf7434f2, 32'hc0316357} /* (19, 16, 9) {real, imag} */,
  {32'hbf2f73c0, 32'h3f5c451e} /* (19, 16, 8) {real, imag} */,
  {32'hbedbf7b9, 32'hc0313432} /* (19, 16, 7) {real, imag} */,
  {32'h3f86ebaa, 32'hbe4b0fec} /* (19, 16, 6) {real, imag} */,
  {32'h3fc94ff9, 32'hc00c07e5} /* (19, 16, 5) {real, imag} */,
  {32'h3cf3009b, 32'hbf9cacf9} /* (19, 16, 4) {real, imag} */,
  {32'hbf9680d5, 32'hbf071950} /* (19, 16, 3) {real, imag} */,
  {32'h3fcaa806, 32'hbfe73e4a} /* (19, 16, 2) {real, imag} */,
  {32'h3f0ff3c9, 32'hbd189fa1} /* (19, 16, 1) {real, imag} */,
  {32'h3f3885e1, 32'h3f780bfb} /* (19, 16, 0) {real, imag} */,
  {32'hbe3dcdf9, 32'hbfaf6cf6} /* (19, 15, 31) {real, imag} */,
  {32'hbd0c06b6, 32'hbec8438b} /* (19, 15, 30) {real, imag} */,
  {32'hc0268ab0, 32'hbf186a94} /* (19, 15, 29) {real, imag} */,
  {32'hbf7a70fa, 32'h3f96271c} /* (19, 15, 28) {real, imag} */,
  {32'hbf07d166, 32'hbe9c7114} /* (19, 15, 27) {real, imag} */,
  {32'hbf83a557, 32'h3e5e8b25} /* (19, 15, 26) {real, imag} */,
  {32'h3fdd05be, 32'hbf0575fe} /* (19, 15, 25) {real, imag} */,
  {32'h3f16db45, 32'hbfa48eaa} /* (19, 15, 24) {real, imag} */,
  {32'h3f2434da, 32'h3f47abd7} /* (19, 15, 23) {real, imag} */,
  {32'h3fb01ac3, 32'h3d78c2c4} /* (19, 15, 22) {real, imag} */,
  {32'h3fda5035, 32'h3da43e5a} /* (19, 15, 21) {real, imag} */,
  {32'h3e6ceb2a, 32'h3f98cae2} /* (19, 15, 20) {real, imag} */,
  {32'hbec48254, 32'h3d1b9b56} /* (19, 15, 19) {real, imag} */,
  {32'hbf80a0de, 32'h3c70b1e5} /* (19, 15, 18) {real, imag} */,
  {32'hc036d731, 32'h3d1ea616} /* (19, 15, 17) {real, imag} */,
  {32'hbf857067, 32'hbf94f879} /* (19, 15, 16) {real, imag} */,
  {32'h3ec5152c, 32'hbe74e783} /* (19, 15, 15) {real, imag} */,
  {32'h401351d7, 32'hbe0d49af} /* (19, 15, 14) {real, imag} */,
  {32'h3fbf2634, 32'h3fd189df} /* (19, 15, 13) {real, imag} */,
  {32'hbf6b3b1c, 32'h3eac2688} /* (19, 15, 12) {real, imag} */,
  {32'h3f0a4dc9, 32'h3d9d5ccf} /* (19, 15, 11) {real, imag} */,
  {32'h3f845b5c, 32'h3dc495dc} /* (19, 15, 10) {real, imag} */,
  {32'hbf2a19ec, 32'hbf4ff088} /* (19, 15, 9) {real, imag} */,
  {32'h3e8852d8, 32'h3fa6c178} /* (19, 15, 8) {real, imag} */,
  {32'hbf40c055, 32'hbf45da1a} /* (19, 15, 7) {real, imag} */,
  {32'hbf4032f7, 32'h3f1af2f5} /* (19, 15, 6) {real, imag} */,
  {32'hbe44ea1e, 32'hbfc5c89f} /* (19, 15, 5) {real, imag} */,
  {32'h3f8ec325, 32'hbef06e27} /* (19, 15, 4) {real, imag} */,
  {32'h3efe6433, 32'hc062a024} /* (19, 15, 3) {real, imag} */,
  {32'h3f57503a, 32'h3fe04e83} /* (19, 15, 2) {real, imag} */,
  {32'hbf237886, 32'hbe552452} /* (19, 15, 1) {real, imag} */,
  {32'h3f46ced1, 32'h3e41b3c8} /* (19, 15, 0) {real, imag} */,
  {32'h3d2d682d, 32'h3f000194} /* (19, 14, 31) {real, imag} */,
  {32'hc02b976e, 32'hbf138f63} /* (19, 14, 30) {real, imag} */,
  {32'hc013810f, 32'hc0031a23} /* (19, 14, 29) {real, imag} */,
  {32'h3fca4a76, 32'hbda439fc} /* (19, 14, 28) {real, imag} */,
  {32'h3f835aa0, 32'h3f8fecc5} /* (19, 14, 27) {real, imag} */,
  {32'h3ea233de, 32'hc00452e2} /* (19, 14, 26) {real, imag} */,
  {32'hbe4445f8, 32'hc01c3efa} /* (19, 14, 25) {real, imag} */,
  {32'hbf2f9ebb, 32'h40086762} /* (19, 14, 24) {real, imag} */,
  {32'hbfcbe129, 32'h3f948145} /* (19, 14, 23) {real, imag} */,
  {32'h3f40cac3, 32'hc01ebcb2} /* (19, 14, 22) {real, imag} */,
  {32'hc05e0a65, 32'hc0179fcf} /* (19, 14, 21) {real, imag} */,
  {32'hbfc3b41c, 32'h3fab2d64} /* (19, 14, 20) {real, imag} */,
  {32'h3f238c42, 32'h3fad1cae} /* (19, 14, 19) {real, imag} */,
  {32'hc0138fbd, 32'h3fec5fc5} /* (19, 14, 18) {real, imag} */,
  {32'h3f46cc17, 32'hbfab0647} /* (19, 14, 17) {real, imag} */,
  {32'h3fdbcfac, 32'hc00b32b7} /* (19, 14, 16) {real, imag} */,
  {32'h3f07807c, 32'hbdc11487} /* (19, 14, 15) {real, imag} */,
  {32'hbe50b200, 32'h3fa7be6e} /* (19, 14, 14) {real, imag} */,
  {32'hbfa5fef5, 32'hbfa32849} /* (19, 14, 13) {real, imag} */,
  {32'hbfcd16fe, 32'h3f439c14} /* (19, 14, 12) {real, imag} */,
  {32'h3e29de31, 32'h3ed90493} /* (19, 14, 11) {real, imag} */,
  {32'hc0bbd7bc, 32'hbf1d7e9a} /* (19, 14, 10) {real, imag} */,
  {32'h3f8a0fe2, 32'hc01b58e3} /* (19, 14, 9) {real, imag} */,
  {32'h40193025, 32'h4014f584} /* (19, 14, 8) {real, imag} */,
  {32'h401d00c6, 32'h402c482e} /* (19, 14, 7) {real, imag} */,
  {32'h3ffad4e1, 32'h3ec8396b} /* (19, 14, 6) {real, imag} */,
  {32'hbf68b3e3, 32'h40173fd6} /* (19, 14, 5) {real, imag} */,
  {32'h3ea38a97, 32'hbf438e22} /* (19, 14, 4) {real, imag} */,
  {32'hbfe30497, 32'h3f026881} /* (19, 14, 3) {real, imag} */,
  {32'h3ee9ad22, 32'h3fa87307} /* (19, 14, 2) {real, imag} */,
  {32'hbe73f42e, 32'h3fb3014b} /* (19, 14, 1) {real, imag} */,
  {32'hbeae6f2f, 32'h3f949a4a} /* (19, 14, 0) {real, imag} */,
  {32'h3f45979b, 32'h3ff3b7ea} /* (19, 13, 31) {real, imag} */,
  {32'h3f3d35d2, 32'hbf2532f0} /* (19, 13, 30) {real, imag} */,
  {32'hc040e9a1, 32'h3f82214a} /* (19, 13, 29) {real, imag} */,
  {32'hc00e3b89, 32'h3f4bd277} /* (19, 13, 28) {real, imag} */,
  {32'hbf0985d8, 32'h3e9675c6} /* (19, 13, 27) {real, imag} */,
  {32'h3eb36d49, 32'h3dceed45} /* (19, 13, 26) {real, imag} */,
  {32'h3e98a113, 32'hc026248a} /* (19, 13, 25) {real, imag} */,
  {32'hbec5755b, 32'h401ae52c} /* (19, 13, 24) {real, imag} */,
  {32'h3fa9c1a6, 32'h3fae7845} /* (19, 13, 23) {real, imag} */,
  {32'hbdcf7ad6, 32'h40123641} /* (19, 13, 22) {real, imag} */,
  {32'h3fc67818, 32'hc04494d1} /* (19, 13, 21) {real, imag} */,
  {32'hbf78f7fd, 32'hbf9cb760} /* (19, 13, 20) {real, imag} */,
  {32'hbde17dc0, 32'h3fe687e9} /* (19, 13, 19) {real, imag} */,
  {32'hc012e86d, 32'hbeddab12} /* (19, 13, 18) {real, imag} */,
  {32'hbed70870, 32'h3e95b68d} /* (19, 13, 17) {real, imag} */,
  {32'hbf5af67e, 32'hbf8a2583} /* (19, 13, 16) {real, imag} */,
  {32'h40515ae3, 32'h3f52bc0a} /* (19, 13, 15) {real, imag} */,
  {32'hbfc3db61, 32'h401218c3} /* (19, 13, 14) {real, imag} */,
  {32'h3f2c5fc4, 32'h3c7e2968} /* (19, 13, 13) {real, imag} */,
  {32'hbea6095b, 32'hbc938828} /* (19, 13, 12) {real, imag} */,
  {32'hc00bf900, 32'hbdd36021} /* (19, 13, 11) {real, imag} */,
  {32'hbf3ae4b2, 32'hbf11c999} /* (19, 13, 10) {real, imag} */,
  {32'h3ee05e4d, 32'hbfd9e257} /* (19, 13, 9) {real, imag} */,
  {32'h3f3696b9, 32'h3f6cb34b} /* (19, 13, 8) {real, imag} */,
  {32'hc02a591a, 32'h3fa44010} /* (19, 13, 7) {real, imag} */,
  {32'h3fc66bc3, 32'hbf7a1418} /* (19, 13, 6) {real, imag} */,
  {32'hc02436ac, 32'h3fa53524} /* (19, 13, 5) {real, imag} */,
  {32'h3f4f0c68, 32'h3eec9da3} /* (19, 13, 4) {real, imag} */,
  {32'h3ed8166b, 32'hbf1e9bf1} /* (19, 13, 3) {real, imag} */,
  {32'hbe33bd2b, 32'h3e957a55} /* (19, 13, 2) {real, imag} */,
  {32'hbdfcfd58, 32'h3fac982b} /* (19, 13, 1) {real, imag} */,
  {32'hbf933048, 32'h3fae7eac} /* (19, 13, 0) {real, imag} */,
  {32'hbf5c55e2, 32'h3f7635b9} /* (19, 12, 31) {real, imag} */,
  {32'hbf52eb1b, 32'hbfe3473c} /* (19, 12, 30) {real, imag} */,
  {32'h402ae09a, 32'h3dd7c69a} /* (19, 12, 29) {real, imag} */,
  {32'hbf0419d9, 32'hbf64e045} /* (19, 12, 28) {real, imag} */,
  {32'hc01eef89, 32'h3f97d24e} /* (19, 12, 27) {real, imag} */,
  {32'h40636ecf, 32'hbee31699} /* (19, 12, 26) {real, imag} */,
  {32'hbe64c248, 32'hbf8469b5} /* (19, 12, 25) {real, imag} */,
  {32'h3fd0a68a, 32'h3f93aee0} /* (19, 12, 24) {real, imag} */,
  {32'hbf011c04, 32'h3fae3da3} /* (19, 12, 23) {real, imag} */,
  {32'hbfce5e24, 32'hbf9bc9ed} /* (19, 12, 22) {real, imag} */,
  {32'hbfc29bd1, 32'hc050b69e} /* (19, 12, 21) {real, imag} */,
  {32'h3fe20a7f, 32'hbe78b6e6} /* (19, 12, 20) {real, imag} */,
  {32'h3e4b886d, 32'hbf7068fd} /* (19, 12, 19) {real, imag} */,
  {32'h3f96b06c, 32'h3f154edc} /* (19, 12, 18) {real, imag} */,
  {32'h3fe10d94, 32'h3fa26324} /* (19, 12, 17) {real, imag} */,
  {32'h3f576731, 32'h3f2bdbb2} /* (19, 12, 16) {real, imag} */,
  {32'h3f01d1d2, 32'h3f9f6df6} /* (19, 12, 15) {real, imag} */,
  {32'hbe2ecb74, 32'hc00e015b} /* (19, 12, 14) {real, imag} */,
  {32'h3f6e77b4, 32'h3fb30f0c} /* (19, 12, 13) {real, imag} */,
  {32'hbf0cd96b, 32'h3e906ea9} /* (19, 12, 12) {real, imag} */,
  {32'hbf5eaa59, 32'hbfd92540} /* (19, 12, 11) {real, imag} */,
  {32'h4039039c, 32'h3fa7869b} /* (19, 12, 10) {real, imag} */,
  {32'h3fc24ae2, 32'hbf8537eb} /* (19, 12, 9) {real, imag} */,
  {32'hbf71328d, 32'hbf2ddcfe} /* (19, 12, 8) {real, imag} */,
  {32'h3fac4d7e, 32'h4083f835} /* (19, 12, 7) {real, imag} */,
  {32'hbfabc57c, 32'hbcea22f9} /* (19, 12, 6) {real, imag} */,
  {32'h3f93d534, 32'h3e561239} /* (19, 12, 5) {real, imag} */,
  {32'hbfeba1f5, 32'h3e116c39} /* (19, 12, 4) {real, imag} */,
  {32'h3ff41e99, 32'hbf48c0eb} /* (19, 12, 3) {real, imag} */,
  {32'hbfbb940c, 32'h3ed885b8} /* (19, 12, 2) {real, imag} */,
  {32'hbf88a583, 32'h3ea655b4} /* (19, 12, 1) {real, imag} */,
  {32'hbf23a953, 32'hbf8b44af} /* (19, 12, 0) {real, imag} */,
  {32'h3d75cc5b, 32'h3ef4c4d9} /* (19, 11, 31) {real, imag} */,
  {32'h3fe52ec4, 32'h3e675589} /* (19, 11, 30) {real, imag} */,
  {32'h3f81bcbe, 32'hbd955671} /* (19, 11, 29) {real, imag} */,
  {32'h3d1b1c2c, 32'hbfa765fe} /* (19, 11, 28) {real, imag} */,
  {32'hbf2f0dfa, 32'hbf8350bc} /* (19, 11, 27) {real, imag} */,
  {32'h3f882ee1, 32'h40abe9ec} /* (19, 11, 26) {real, imag} */,
  {32'hc0350b4f, 32'hbddc3fed} /* (19, 11, 25) {real, imag} */,
  {32'h400ed26e, 32'h3fcd03d9} /* (19, 11, 24) {real, imag} */,
  {32'h3fba2f74, 32'h400ab74c} /* (19, 11, 23) {real, imag} */,
  {32'hbf2f59f9, 32'hbf81a9e0} /* (19, 11, 22) {real, imag} */,
  {32'h3f1c8841, 32'hc06bca9d} /* (19, 11, 21) {real, imag} */,
  {32'h3ff4ce83, 32'hbf262235} /* (19, 11, 20) {real, imag} */,
  {32'h406ac0f3, 32'hbefecb1a} /* (19, 11, 19) {real, imag} */,
  {32'hbe8f7c1f, 32'h3f952d6c} /* (19, 11, 18) {real, imag} */,
  {32'hbfe0ce3e, 32'h40013f04} /* (19, 11, 17) {real, imag} */,
  {32'hbeb1b03a, 32'hbf84b4f9} /* (19, 11, 16) {real, imag} */,
  {32'h3da40425, 32'h3ed55bb5} /* (19, 11, 15) {real, imag} */,
  {32'h3f09b1d8, 32'hbf984ce3} /* (19, 11, 14) {real, imag} */,
  {32'hc01c3ed8, 32'hbf1c3af7} /* (19, 11, 13) {real, imag} */,
  {32'h3e8223c6, 32'h4007a0a8} /* (19, 11, 12) {real, imag} */,
  {32'h4053cdca, 32'h3facda74} /* (19, 11, 11) {real, imag} */,
  {32'hbeee8998, 32'h3ec57de0} /* (19, 11, 10) {real, imag} */,
  {32'hbdfc744a, 32'h3dddf18c} /* (19, 11, 9) {real, imag} */,
  {32'hbf80530a, 32'hc0022742} /* (19, 11, 8) {real, imag} */,
  {32'h4055da5c, 32'hbdceffa3} /* (19, 11, 7) {real, imag} */,
  {32'hc00bacc7, 32'hbf3bb078} /* (19, 11, 6) {real, imag} */,
  {32'hbef2aab1, 32'h402e53fe} /* (19, 11, 5) {real, imag} */,
  {32'h3ed98103, 32'h3ccde61f} /* (19, 11, 4) {real, imag} */,
  {32'h40758a6b, 32'hc07559be} /* (19, 11, 3) {real, imag} */,
  {32'hbf69f417, 32'hc068d311} /* (19, 11, 2) {real, imag} */,
  {32'hbdebf633, 32'hbf58659c} /* (19, 11, 1) {real, imag} */,
  {32'hbe90bead, 32'h3e0ba29d} /* (19, 11, 0) {real, imag} */,
  {32'hc000eb2c, 32'h3f81c1c7} /* (19, 10, 31) {real, imag} */,
  {32'hbfb65988, 32'h3d563b9e} /* (19, 10, 30) {real, imag} */,
  {32'h3fc4ac77, 32'h3d899b15} /* (19, 10, 29) {real, imag} */,
  {32'h3fa25a21, 32'h3fcb312f} /* (19, 10, 28) {real, imag} */,
  {32'h3ffece93, 32'hc00419e8} /* (19, 10, 27) {real, imag} */,
  {32'hc049f214, 32'hc0153c08} /* (19, 10, 26) {real, imag} */,
  {32'h3f54260a, 32'hbff48446} /* (19, 10, 25) {real, imag} */,
  {32'h3f12f01b, 32'hbed22d13} /* (19, 10, 24) {real, imag} */,
  {32'h3fae7ec8, 32'hbe10b62f} /* (19, 10, 23) {real, imag} */,
  {32'h3fc90a29, 32'hbe5ec26c} /* (19, 10, 22) {real, imag} */,
  {32'hc00e9055, 32'hc00542fe} /* (19, 10, 21) {real, imag} */,
  {32'h3f2abf6c, 32'hbf637970} /* (19, 10, 20) {real, imag} */,
  {32'hbff96347, 32'h3ec92b28} /* (19, 10, 19) {real, imag} */,
  {32'h3f8b574d, 32'h402a823e} /* (19, 10, 18) {real, imag} */,
  {32'hc013758b, 32'h3f66260d} /* (19, 10, 17) {real, imag} */,
  {32'hbf19dfc3, 32'hbc14cedd} /* (19, 10, 16) {real, imag} */,
  {32'hbf1fd9f1, 32'hbd8d74ec} /* (19, 10, 15) {real, imag} */,
  {32'h3e987bed, 32'hc08cc98a} /* (19, 10, 14) {real, imag} */,
  {32'h3fe57acc, 32'hbf0f9460} /* (19, 10, 13) {real, imag} */,
  {32'h3f055f30, 32'hc04b430a} /* (19, 10, 12) {real, imag} */,
  {32'hc0a0d07c, 32'hbef33680} /* (19, 10, 11) {real, imag} */,
  {32'hc051a0cf, 32'h3fe78265} /* (19, 10, 10) {real, imag} */,
  {32'h3f138e67, 32'h4051795f} /* (19, 10, 9) {real, imag} */,
  {32'h401c4b6d, 32'h3f022060} /* (19, 10, 8) {real, imag} */,
  {32'hbfcd0069, 32'h3f24714c} /* (19, 10, 7) {real, imag} */,
  {32'hbf028ee2, 32'hbf5cd0f4} /* (19, 10, 6) {real, imag} */,
  {32'hbf548591, 32'hbf6d566b} /* (19, 10, 5) {real, imag} */,
  {32'h3e914bd5, 32'h3fbda0d5} /* (19, 10, 4) {real, imag} */,
  {32'h3ff9f9c6, 32'h3fcf8540} /* (19, 10, 3) {real, imag} */,
  {32'hbf7054c5, 32'h3f0553fe} /* (19, 10, 2) {real, imag} */,
  {32'hbf1d459e, 32'hc00abd72} /* (19, 10, 1) {real, imag} */,
  {32'h3feada62, 32'h3ffabfb5} /* (19, 10, 0) {real, imag} */,
  {32'h3f835112, 32'hc02e41ff} /* (19, 9, 31) {real, imag} */,
  {32'h4031b6a8, 32'h3fcef66e} /* (19, 9, 30) {real, imag} */,
  {32'hbe5a34fb, 32'h3f4aabec} /* (19, 9, 29) {real, imag} */,
  {32'h3e27a190, 32'hbd09ee74} /* (19, 9, 28) {real, imag} */,
  {32'h400abcee, 32'hbf997643} /* (19, 9, 27) {real, imag} */,
  {32'hbf5badd3, 32'h40734be4} /* (19, 9, 26) {real, imag} */,
  {32'h3f4de0ca, 32'hbfc8b86c} /* (19, 9, 25) {real, imag} */,
  {32'hbe86cbb3, 32'hc01429cc} /* (19, 9, 24) {real, imag} */,
  {32'hc0040494, 32'h3ffd8222} /* (19, 9, 23) {real, imag} */,
  {32'hbf11fd85, 32'h4010011a} /* (19, 9, 22) {real, imag} */,
  {32'h400aadde, 32'h407f6599} /* (19, 9, 21) {real, imag} */,
  {32'h3e407775, 32'h3f2655b5} /* (19, 9, 20) {real, imag} */,
  {32'h408cb313, 32'hbfbecbfb} /* (19, 9, 19) {real, imag} */,
  {32'hc0208e79, 32'hc083fc26} /* (19, 9, 18) {real, imag} */,
  {32'hc0190014, 32'h3eaa8ee8} /* (19, 9, 17) {real, imag} */,
  {32'hbfa5a0a6, 32'h3fb2159f} /* (19, 9, 16) {real, imag} */,
  {32'hbfc85edf, 32'h3ec91a28} /* (19, 9, 15) {real, imag} */,
  {32'h3f98aabf, 32'hbf0890ea} /* (19, 9, 14) {real, imag} */,
  {32'h3f126178, 32'hbbbb8de3} /* (19, 9, 13) {real, imag} */,
  {32'h3ccb8c60, 32'h403502ad} /* (19, 9, 12) {real, imag} */,
  {32'h3f7d83f7, 32'hbf0f2889} /* (19, 9, 11) {real, imag} */,
  {32'h3d7f093e, 32'hbe0c4140} /* (19, 9, 10) {real, imag} */,
  {32'hbf1da512, 32'hc02c41df} /* (19, 9, 9) {real, imag} */,
  {32'h3f94855e, 32'h408d5266} /* (19, 9, 8) {real, imag} */,
  {32'hbf3c60e7, 32'h3f5555ec} /* (19, 9, 7) {real, imag} */,
  {32'h3f109a31, 32'h4070cbe1} /* (19, 9, 6) {real, imag} */,
  {32'hbfeb414e, 32'hbda934ca} /* (19, 9, 5) {real, imag} */,
  {32'h3f046593, 32'h3f5cd0f7} /* (19, 9, 4) {real, imag} */,
  {32'h3f9d368a, 32'hbe38b741} /* (19, 9, 3) {real, imag} */,
  {32'h3ed2a0c2, 32'hc00803b9} /* (19, 9, 2) {real, imag} */,
  {32'hc001e325, 32'hc0381a1a} /* (19, 9, 1) {real, imag} */,
  {32'hbefef943, 32'hbfad98f3} /* (19, 9, 0) {real, imag} */,
  {32'hbede5528, 32'h4003af7d} /* (19, 8, 31) {real, imag} */,
  {32'h3f85b4db, 32'h3fb0119f} /* (19, 8, 30) {real, imag} */,
  {32'hbe84368d, 32'h3e930abd} /* (19, 8, 29) {real, imag} */,
  {32'h4005a25b, 32'hc008bb97} /* (19, 8, 28) {real, imag} */,
  {32'hbf7a2724, 32'hbf5b6795} /* (19, 8, 27) {real, imag} */,
  {32'h3f090b7b, 32'hbf8725da} /* (19, 8, 26) {real, imag} */,
  {32'hbf772111, 32'h400c2330} /* (19, 8, 25) {real, imag} */,
  {32'h3f66824c, 32'h3ff82c36} /* (19, 8, 24) {real, imag} */,
  {32'h3f76234b, 32'hbf0b3a56} /* (19, 8, 23) {real, imag} */,
  {32'hbf8fd421, 32'hbf12fe5c} /* (19, 8, 22) {real, imag} */,
  {32'h3ed56f74, 32'hbf173496} /* (19, 8, 21) {real, imag} */,
  {32'hbf4c54c0, 32'hbfab6e09} /* (19, 8, 20) {real, imag} */,
  {32'h3ffb3670, 32'h408e5b74} /* (19, 8, 19) {real, imag} */,
  {32'h3e98394b, 32'hbfad6dea} /* (19, 8, 18) {real, imag} */,
  {32'h3f38eb89, 32'hbf58a271} /* (19, 8, 17) {real, imag} */,
  {32'hbdeb2d30, 32'hbf4d63b2} /* (19, 8, 16) {real, imag} */,
  {32'hc010b464, 32'hbe2c432e} /* (19, 8, 15) {real, imag} */,
  {32'h3ec5ae7e, 32'hc038d761} /* (19, 8, 14) {real, imag} */,
  {32'hbfa37834, 32'h3fb93a0e} /* (19, 8, 13) {real, imag} */,
  {32'hbfccb8d9, 32'h3df5e3ee} /* (19, 8, 12) {real, imag} */,
  {32'h403a1f72, 32'h400f910b} /* (19, 8, 11) {real, imag} */,
  {32'h3ee00def, 32'h3fa3a700} /* (19, 8, 10) {real, imag} */,
  {32'hbf563b5d, 32'h3f29db63} /* (19, 8, 9) {real, imag} */,
  {32'h40939bbc, 32'h3ee6e0e1} /* (19, 8, 8) {real, imag} */,
  {32'h3e70104b, 32'h3ec3b6bc} /* (19, 8, 7) {real, imag} */,
  {32'hbfbd4312, 32'hbffe50aa} /* (19, 8, 6) {real, imag} */,
  {32'hbd997626, 32'h3ffac31f} /* (19, 8, 5) {real, imag} */,
  {32'hbe910c86, 32'hbf79ab2a} /* (19, 8, 4) {real, imag} */,
  {32'hbfa9e043, 32'hbec79c04} /* (19, 8, 3) {real, imag} */,
  {32'hc0014a6f, 32'h3fd347b6} /* (19, 8, 2) {real, imag} */,
  {32'hbf2657a0, 32'hbd52db8b} /* (19, 8, 1) {real, imag} */,
  {32'h3f0293ba, 32'h3f2a190b} /* (19, 8, 0) {real, imag} */,
  {32'hbf9debd9, 32'hbf134d54} /* (19, 7, 31) {real, imag} */,
  {32'h3deb1db7, 32'hc047a9b4} /* (19, 7, 30) {real, imag} */,
  {32'hbe9b615e, 32'h404e9027} /* (19, 7, 29) {real, imag} */,
  {32'hbdcbc391, 32'h3e874311} /* (19, 7, 28) {real, imag} */,
  {32'hbfc9c89f, 32'hc065e5bc} /* (19, 7, 27) {real, imag} */,
  {32'hbebb8dd3, 32'h3fb921b2} /* (19, 7, 26) {real, imag} */,
  {32'h4042ea35, 32'h400601f6} /* (19, 7, 25) {real, imag} */,
  {32'hbff4463c, 32'h3fd276fd} /* (19, 7, 24) {real, imag} */,
  {32'h3d3cf253, 32'h3eb8ee35} /* (19, 7, 23) {real, imag} */,
  {32'h406b60bc, 32'hbf3059ce} /* (19, 7, 22) {real, imag} */,
  {32'h3fe48ff9, 32'hbfda3c1c} /* (19, 7, 21) {real, imag} */,
  {32'h3ef6a463, 32'hc00a68ba} /* (19, 7, 20) {real, imag} */,
  {32'h3fa8d75e, 32'hc0383439} /* (19, 7, 19) {real, imag} */,
  {32'h3f3a0807, 32'h3ee11498} /* (19, 7, 18) {real, imag} */,
  {32'hbf855535, 32'hbe93177b} /* (19, 7, 17) {real, imag} */,
  {32'h3f241a50, 32'h3f225f1f} /* (19, 7, 16) {real, imag} */,
  {32'h3f318348, 32'hbdd1115b} /* (19, 7, 15) {real, imag} */,
  {32'hbf2d21bf, 32'h3fb2ae55} /* (19, 7, 14) {real, imag} */,
  {32'h3f85fa31, 32'hbea8f0f6} /* (19, 7, 13) {real, imag} */,
  {32'h40108c00, 32'h401db4a6} /* (19, 7, 12) {real, imag} */,
  {32'h3f039d20, 32'h3f90e26a} /* (19, 7, 11) {real, imag} */,
  {32'h3ffcb52e, 32'hbf2b87ee} /* (19, 7, 10) {real, imag} */,
  {32'h3fa8c0b6, 32'hbf8ecb1a} /* (19, 7, 9) {real, imag} */,
  {32'h3e864f1a, 32'hbed9412e} /* (19, 7, 8) {real, imag} */,
  {32'hc0085214, 32'h3f092a69} /* (19, 7, 7) {real, imag} */,
  {32'hbf6d6bbe, 32'hc046944d} /* (19, 7, 6) {real, imag} */,
  {32'hc020f95d, 32'hbe4b289e} /* (19, 7, 5) {real, imag} */,
  {32'h3f37e1a9, 32'h3fbf5c5e} /* (19, 7, 4) {real, imag} */,
  {32'hbfa2c4f9, 32'hbee35204} /* (19, 7, 3) {real, imag} */,
  {32'hc0926d36, 32'h3f8da410} /* (19, 7, 2) {real, imag} */,
  {32'hbf881d0d, 32'hbf1203ba} /* (19, 7, 1) {real, imag} */,
  {32'h3f5bccdf, 32'h3f1bec7e} /* (19, 7, 0) {real, imag} */,
  {32'h403217d7, 32'hc0336ce9} /* (19, 6, 31) {real, imag} */,
  {32'h3f2cbe54, 32'hbf38c539} /* (19, 6, 30) {real, imag} */,
  {32'h40036281, 32'hbfaafc99} /* (19, 6, 29) {real, imag} */,
  {32'hbf304605, 32'h3f916529} /* (19, 6, 28) {real, imag} */,
  {32'h3ebc335f, 32'h3f0a3dd8} /* (19, 6, 27) {real, imag} */,
  {32'hbfb8c8b7, 32'hbf8ec327} /* (19, 6, 26) {real, imag} */,
  {32'h3f652444, 32'h40210e59} /* (19, 6, 25) {real, imag} */,
  {32'h3d883b3c, 32'hc02038fb} /* (19, 6, 24) {real, imag} */,
  {32'h3fc3d318, 32'h3fd502c8} /* (19, 6, 23) {real, imag} */,
  {32'hc02c05b5, 32'h3eb293af} /* (19, 6, 22) {real, imag} */,
  {32'h3fbc9430, 32'h3f411cd4} /* (19, 6, 21) {real, imag} */,
  {32'h3f43f133, 32'hbd9b5cf1} /* (19, 6, 20) {real, imag} */,
  {32'hbf6d6404, 32'hbf43d20c} /* (19, 6, 19) {real, imag} */,
  {32'h3f6cf7d0, 32'h3fce541a} /* (19, 6, 18) {real, imag} */,
  {32'h3f29d381, 32'h40030d48} /* (19, 6, 17) {real, imag} */,
  {32'h3f06ff5b, 32'h40050ebe} /* (19, 6, 16) {real, imag} */,
  {32'hbf8d5abf, 32'hbfd6e089} /* (19, 6, 15) {real, imag} */,
  {32'hc0857c87, 32'h401ccdcb} /* (19, 6, 14) {real, imag} */,
  {32'h3f06c96f, 32'h3f823e39} /* (19, 6, 13) {real, imag} */,
  {32'h3fd8fd13, 32'h3f832d61} /* (19, 6, 12) {real, imag} */,
  {32'h3fcb16e6, 32'h40090d79} /* (19, 6, 11) {real, imag} */,
  {32'hbf14c43a, 32'hbf183dc8} /* (19, 6, 10) {real, imag} */,
  {32'hc060d929, 32'hbfe27258} /* (19, 6, 9) {real, imag} */,
  {32'hbe9c5a90, 32'h3f82febe} /* (19, 6, 8) {real, imag} */,
  {32'hc0383d42, 32'hbf2b3fce} /* (19, 6, 7) {real, imag} */,
  {32'hc0191ea7, 32'h3e2a0e17} /* (19, 6, 6) {real, imag} */,
  {32'h3f85bd92, 32'hbfe73392} /* (19, 6, 5) {real, imag} */,
  {32'h3f986231, 32'hbee17696} /* (19, 6, 4) {real, imag} */,
  {32'hbfadf627, 32'hbfbb1a00} /* (19, 6, 3) {real, imag} */,
  {32'hbfd33b26, 32'hbf95cfb5} /* (19, 6, 2) {real, imag} */,
  {32'h400ca8ea, 32'hc044238f} /* (19, 6, 1) {real, imag} */,
  {32'h3d53f41a, 32'h4003807d} /* (19, 6, 0) {real, imag} */,
  {32'h3f237f33, 32'hbfdda81e} /* (19, 5, 31) {real, imag} */,
  {32'hbfc4fdb8, 32'hbf4eaf14} /* (19, 5, 30) {real, imag} */,
  {32'hbe9cc80f, 32'hbf4ff48a} /* (19, 5, 29) {real, imag} */,
  {32'hbd27e359, 32'h4068b32c} /* (19, 5, 28) {real, imag} */,
  {32'hc013d293, 32'h3fa1503a} /* (19, 5, 27) {real, imag} */,
  {32'h4003822a, 32'hbf3c5e2a} /* (19, 5, 26) {real, imag} */,
  {32'hbfd81ef2, 32'h3ecc1bfe} /* (19, 5, 25) {real, imag} */,
  {32'hc0066bd6, 32'h3fd1692a} /* (19, 5, 24) {real, imag} */,
  {32'hc0330aec, 32'h3f20edec} /* (19, 5, 23) {real, imag} */,
  {32'h3e037307, 32'hc02c6d53} /* (19, 5, 22) {real, imag} */,
  {32'h4047f8fa, 32'hbc9d0982} /* (19, 5, 21) {real, imag} */,
  {32'hbeccf355, 32'hbfbbc49b} /* (19, 5, 20) {real, imag} */,
  {32'hbf178001, 32'hbef75b5b} /* (19, 5, 19) {real, imag} */,
  {32'hc01721c4, 32'hc04bd86b} /* (19, 5, 18) {real, imag} */,
  {32'h3f3c61a8, 32'hc02c0fc2} /* (19, 5, 17) {real, imag} */,
  {32'h3ee9bb01, 32'hbfad1683} /* (19, 5, 16) {real, imag} */,
  {32'hbf1c64e0, 32'h3ee30bfb} /* (19, 5, 15) {real, imag} */,
  {32'hc00a1b70, 32'h3f2310a5} /* (19, 5, 14) {real, imag} */,
  {32'h3eb96862, 32'h3fb164b1} /* (19, 5, 13) {real, imag} */,
  {32'h3ed2e465, 32'hbf753ccd} /* (19, 5, 12) {real, imag} */,
  {32'h3f02861d, 32'hbf99397f} /* (19, 5, 11) {real, imag} */,
  {32'h4042520b, 32'hbf9a84ec} /* (19, 5, 10) {real, imag} */,
  {32'h402825c3, 32'h3d9c62f7} /* (19, 5, 9) {real, imag} */,
  {32'hc07d655a, 32'h3f651364} /* (19, 5, 8) {real, imag} */,
  {32'hc043d8d1, 32'h3e293f47} /* (19, 5, 7) {real, imag} */,
  {32'h3ea68e7a, 32'hc015b32a} /* (19, 5, 6) {real, imag} */,
  {32'h40285685, 32'h3ffbe71c} /* (19, 5, 5) {real, imag} */,
  {32'hbff9c7a0, 32'h3f675c9c} /* (19, 5, 4) {real, imag} */,
  {32'h4023c5c4, 32'hbf76e7a8} /* (19, 5, 3) {real, imag} */,
  {32'h3e932ddc, 32'hbd8f60d4} /* (19, 5, 2) {real, imag} */,
  {32'h3f1b382c, 32'h40261133} /* (19, 5, 1) {real, imag} */,
  {32'hbfeb117c, 32'h3f9dc393} /* (19, 5, 0) {real, imag} */,
  {32'h3f318107, 32'hbf95acbe} /* (19, 4, 31) {real, imag} */,
  {32'hc05e57e2, 32'h4000dff6} /* (19, 4, 30) {real, imag} */,
  {32'h3d855dac, 32'h3f87f1a6} /* (19, 4, 29) {real, imag} */,
  {32'h3f853523, 32'h3e1b1393} /* (19, 4, 28) {real, imag} */,
  {32'h3e0fefe6, 32'h3dca351d} /* (19, 4, 27) {real, imag} */,
  {32'hbf860d01, 32'h400d7c88} /* (19, 4, 26) {real, imag} */,
  {32'h404ab81f, 32'hbfb115c8} /* (19, 4, 25) {real, imag} */,
  {32'h3fcbc0c5, 32'hc0199400} /* (19, 4, 24) {real, imag} */,
  {32'hc009defe, 32'hbf0cd779} /* (19, 4, 23) {real, imag} */,
  {32'h402a6c2f, 32'hc0145b6b} /* (19, 4, 22) {real, imag} */,
  {32'h3fc06290, 32'hbfd8dabb} /* (19, 4, 21) {real, imag} */,
  {32'hc067cf31, 32'h3e06a32d} /* (19, 4, 20) {real, imag} */,
  {32'hc043e36e, 32'h4014e6ae} /* (19, 4, 19) {real, imag} */,
  {32'hbf91c6db, 32'h402a2d8f} /* (19, 4, 18) {real, imag} */,
  {32'h3f5c8079, 32'hbf7098ed} /* (19, 4, 17) {real, imag} */,
  {32'h3f42487b, 32'h3f5c9da4} /* (19, 4, 16) {real, imag} */,
  {32'hbfd08462, 32'h3ffccd6f} /* (19, 4, 15) {real, imag} */,
  {32'h3facf103, 32'h3f7c5f50} /* (19, 4, 14) {real, imag} */,
  {32'hbe07d7d4, 32'h3fa6a208} /* (19, 4, 13) {real, imag} */,
  {32'hbf9b5818, 32'h40192717} /* (19, 4, 12) {real, imag} */,
  {32'hc01c0ebb, 32'h40155bd6} /* (19, 4, 11) {real, imag} */,
  {32'h3fa52772, 32'hbe8e6396} /* (19, 4, 10) {real, imag} */,
  {32'hbd8fe2cc, 32'hc00a7694} /* (19, 4, 9) {real, imag} */,
  {32'h3f104bf6, 32'h3f2649ec} /* (19, 4, 8) {real, imag} */,
  {32'h3e64e239, 32'h3f47f661} /* (19, 4, 7) {real, imag} */,
  {32'hbfb6cd7a, 32'hbf449f0a} /* (19, 4, 6) {real, imag} */,
  {32'hbf5154d4, 32'h3f67840a} /* (19, 4, 5) {real, imag} */,
  {32'h3f2ea902, 32'hbfc69aea} /* (19, 4, 4) {real, imag} */,
  {32'hbfb8d0a2, 32'h3fbbb737} /* (19, 4, 3) {real, imag} */,
  {32'h3fca7b9d, 32'hc069ce15} /* (19, 4, 2) {real, imag} */,
  {32'hbd099138, 32'h40667871} /* (19, 4, 1) {real, imag} */,
  {32'hc00d0987, 32'hbdfa706b} /* (19, 4, 0) {real, imag} */,
  {32'hbd872f9c, 32'hbfffecc2} /* (19, 3, 31) {real, imag} */,
  {32'h3f2c8bc4, 32'h401bbeb5} /* (19, 3, 30) {real, imag} */,
  {32'hbdda91ce, 32'hc020b40d} /* (19, 3, 29) {real, imag} */,
  {32'h3e9a6d24, 32'hc004c063} /* (19, 3, 28) {real, imag} */,
  {32'hbfcf71f7, 32'h3f6981eb} /* (19, 3, 27) {real, imag} */,
  {32'h3f23adfe, 32'h3f813d8b} /* (19, 3, 26) {real, imag} */,
  {32'h3f924d37, 32'h3fa337b1} /* (19, 3, 25) {real, imag} */,
  {32'hbfb5a16e, 32'h3f1d85a9} /* (19, 3, 24) {real, imag} */,
  {32'h3f1a1a52, 32'h3f807460} /* (19, 3, 23) {real, imag} */,
  {32'hc002fe60, 32'h4006de93} /* (19, 3, 22) {real, imag} */,
  {32'hc02b195f, 32'h3ff37214} /* (19, 3, 21) {real, imag} */,
  {32'h3e015286, 32'hbf95955c} /* (19, 3, 20) {real, imag} */,
  {32'hbf159321, 32'h3ffe0073} /* (19, 3, 19) {real, imag} */,
  {32'hbf556262, 32'h3faa388c} /* (19, 3, 18) {real, imag} */,
  {32'hbf655a0f, 32'hbfcbdd9d} /* (19, 3, 17) {real, imag} */,
  {32'hbfb99bf3, 32'hbfdcad23} /* (19, 3, 16) {real, imag} */,
  {32'h3d885361, 32'hbfd6fbcd} /* (19, 3, 15) {real, imag} */,
  {32'hbe46fcfe, 32'hc044965f} /* (19, 3, 14) {real, imag} */,
  {32'h3f964bb4, 32'h40362592} /* (19, 3, 13) {real, imag} */,
  {32'h4022aba4, 32'hc0288f1f} /* (19, 3, 12) {real, imag} */,
  {32'hc011b8f8, 32'h3f025f71} /* (19, 3, 11) {real, imag} */,
  {32'h3fec9a34, 32'hbed9f288} /* (19, 3, 10) {real, imag} */,
  {32'h3ea9e1b3, 32'hbec27f2b} /* (19, 3, 9) {real, imag} */,
  {32'h400e1d7c, 32'h400dabf9} /* (19, 3, 8) {real, imag} */,
  {32'hbf4fc6a7, 32'hbf4cf577} /* (19, 3, 7) {real, imag} */,
  {32'h40896e94, 32'hbf6ba95c} /* (19, 3, 6) {real, imag} */,
  {32'h3dad3d8d, 32'h3eacd4e5} /* (19, 3, 5) {real, imag} */,
  {32'hbffe29a0, 32'h3fe6db48} /* (19, 3, 4) {real, imag} */,
  {32'hbfa5244d, 32'h3d204964} /* (19, 3, 3) {real, imag} */,
  {32'hbff0673c, 32'h3f38f065} /* (19, 3, 2) {real, imag} */,
  {32'h3fdd4bdd, 32'hbf96ae68} /* (19, 3, 1) {real, imag} */,
  {32'h3ebf3eb5, 32'hbf88494d} /* (19, 3, 0) {real, imag} */,
  {32'h3effd838, 32'h3f722086} /* (19, 2, 31) {real, imag} */,
  {32'h3f3315c4, 32'h4053ea2b} /* (19, 2, 30) {real, imag} */,
  {32'h3f43bfc4, 32'hbfefc689} /* (19, 2, 29) {real, imag} */,
  {32'hbf6b0955, 32'hbfd613d4} /* (19, 2, 28) {real, imag} */,
  {32'hbfe7c642, 32'hbfd80312} /* (19, 2, 27) {real, imag} */,
  {32'hc05f7d8a, 32'h3e7e3163} /* (19, 2, 26) {real, imag} */,
  {32'hbfa05bbc, 32'h405b2b21} /* (19, 2, 25) {real, imag} */,
  {32'h40068fc2, 32'hbff514ce} /* (19, 2, 24) {real, imag} */,
  {32'hbf86fa20, 32'hc013f16c} /* (19, 2, 23) {real, imag} */,
  {32'h401cbddf, 32'hbe502065} /* (19, 2, 22) {real, imag} */,
  {32'h4039c234, 32'hbfcf5390} /* (19, 2, 21) {real, imag} */,
  {32'hbf027857, 32'h3f914281} /* (19, 2, 20) {real, imag} */,
  {32'hbfc68e8e, 32'h3f648dd5} /* (19, 2, 19) {real, imag} */,
  {32'h3e5facd3, 32'hbebc6d4a} /* (19, 2, 18) {real, imag} */,
  {32'h3f07d194, 32'hbe7ea1dc} /* (19, 2, 17) {real, imag} */,
  {32'hbfa35fda, 32'hbffefc0a} /* (19, 2, 16) {real, imag} */,
  {32'h3f118474, 32'h3ef1a3c3} /* (19, 2, 15) {real, imag} */,
  {32'hbf782684, 32'hbfa983b4} /* (19, 2, 14) {real, imag} */,
  {32'h3d353410, 32'hbfc6aec9} /* (19, 2, 13) {real, imag} */,
  {32'h4019f84e, 32'hbf53bb8f} /* (19, 2, 12) {real, imag} */,
  {32'hbeff58d7, 32'hbea01119} /* (19, 2, 11) {real, imag} */,
  {32'h400bd7db, 32'hbfb60958} /* (19, 2, 10) {real, imag} */,
  {32'h3f5f9e4f, 32'h3f84548b} /* (19, 2, 9) {real, imag} */,
  {32'hbe67bafb, 32'hbdbb9ccc} /* (19, 2, 8) {real, imag} */,
  {32'h3e2714a9, 32'h40089e36} /* (19, 2, 7) {real, imag} */,
  {32'hbeca0764, 32'hc000fbff} /* (19, 2, 6) {real, imag} */,
  {32'h3f3e3fac, 32'hbdd35f49} /* (19, 2, 5) {real, imag} */,
  {32'h3ed1fe4e, 32'h3f5f6810} /* (19, 2, 4) {real, imag} */,
  {32'hbf909032, 32'h3d099eba} /* (19, 2, 3) {real, imag} */,
  {32'h3f81e39c, 32'hbfb4e074} /* (19, 2, 2) {real, imag} */,
  {32'hbf8f1f45, 32'h40056b4b} /* (19, 2, 1) {real, imag} */,
  {32'hbfc4e39d, 32'h3f34589e} /* (19, 2, 0) {real, imag} */,
  {32'h3f2ef35a, 32'h3ee2f513} /* (19, 1, 31) {real, imag} */,
  {32'h3ff71f03, 32'h3e8d60e0} /* (19, 1, 30) {real, imag} */,
  {32'hc01ed3c0, 32'hbfaa5300} /* (19, 1, 29) {real, imag} */,
  {32'h3e35aae4, 32'h3f401dbd} /* (19, 1, 28) {real, imag} */,
  {32'h3f9d75a7, 32'h40487447} /* (19, 1, 27) {real, imag} */,
  {32'h3f444f7d, 32'h405a95d1} /* (19, 1, 26) {real, imag} */,
  {32'hbfa0271c, 32'hbe642e89} /* (19, 1, 25) {real, imag} */,
  {32'hbdb9545b, 32'hbed0e0b9} /* (19, 1, 24) {real, imag} */,
  {32'hbef8bb2f, 32'hc064a2e2} /* (19, 1, 23) {real, imag} */,
  {32'h3d967cb9, 32'hc01ed1ce} /* (19, 1, 22) {real, imag} */,
  {32'hbfb5ecaf, 32'h3fcde70d} /* (19, 1, 21) {real, imag} */,
  {32'h3ff1c961, 32'h3ff1d33a} /* (19, 1, 20) {real, imag} */,
  {32'hbd169314, 32'h3e8fdd21} /* (19, 1, 19) {real, imag} */,
  {32'h3e2fb7e5, 32'hbf4cd226} /* (19, 1, 18) {real, imag} */,
  {32'h3fa4da85, 32'h3f11d487} /* (19, 1, 17) {real, imag} */,
  {32'hbe6262a8, 32'h3f2f44b7} /* (19, 1, 16) {real, imag} */,
  {32'h3f6e564c, 32'hbe539b0b} /* (19, 1, 15) {real, imag} */,
  {32'hbd839fd4, 32'h3fbc7c48} /* (19, 1, 14) {real, imag} */,
  {32'hc012248d, 32'hbf828752} /* (19, 1, 13) {real, imag} */,
  {32'hbf2ec150, 32'hbfc13e4b} /* (19, 1, 12) {real, imag} */,
  {32'h3f1e5676, 32'hc079fe77} /* (19, 1, 11) {real, imag} */,
  {32'h3f5b1b7c, 32'h4009d831} /* (19, 1, 10) {real, imag} */,
  {32'hbfb197d5, 32'h3f8473dc} /* (19, 1, 9) {real, imag} */,
  {32'h3fff4c8f, 32'h3fd48c05} /* (19, 1, 8) {real, imag} */,
  {32'hbfbb2c7a, 32'hbe9f72b6} /* (19, 1, 7) {real, imag} */,
  {32'h3cd2a8b6, 32'h3fbdd617} /* (19, 1, 6) {real, imag} */,
  {32'hc028e4ec, 32'hbf833175} /* (19, 1, 5) {real, imag} */,
  {32'h40148d9e, 32'h3ef5a9ba} /* (19, 1, 4) {real, imag} */,
  {32'hbf0573fd, 32'hbf86df1e} /* (19, 1, 3) {real, imag} */,
  {32'hbf4ad4a2, 32'h3df1b2d4} /* (19, 1, 2) {real, imag} */,
  {32'hbea0a70e, 32'h3fa972ed} /* (19, 1, 1) {real, imag} */,
  {32'h3f41c080, 32'hbf286788} /* (19, 1, 0) {real, imag} */,
  {32'h3f459184, 32'h403aceef} /* (19, 0, 31) {real, imag} */,
  {32'hbe97d10c, 32'h3fb1fa94} /* (19, 0, 30) {real, imag} */,
  {32'h3fdce0fe, 32'h3fb5c528} /* (19, 0, 29) {real, imag} */,
  {32'h3f9407a7, 32'h401e3167} /* (19, 0, 28) {real, imag} */,
  {32'h3dc7bdbf, 32'h3f8ee409} /* (19, 0, 27) {real, imag} */,
  {32'hc0160973, 32'h3facb501} /* (19, 0, 26) {real, imag} */,
  {32'hbf2e55e9, 32'hbfb0cd75} /* (19, 0, 25) {real, imag} */,
  {32'hbfb158f0, 32'hbe69df8a} /* (19, 0, 24) {real, imag} */,
  {32'h3d9a6281, 32'h3f86ff59} /* (19, 0, 23) {real, imag} */,
  {32'hc0077c1f, 32'h3faaa56f} /* (19, 0, 22) {real, imag} */,
  {32'h3f61efb8, 32'hbf71d034} /* (19, 0, 21) {real, imag} */,
  {32'h3f130ef1, 32'h3ef3fef0} /* (19, 0, 20) {real, imag} */,
  {32'h3f0eb28f, 32'hbee95a10} /* (19, 0, 19) {real, imag} */,
  {32'h3d26f8f6, 32'hbe0acad4} /* (19, 0, 18) {real, imag} */,
  {32'hbe702583, 32'h3e83d7cf} /* (19, 0, 17) {real, imag} */,
  {32'hc0101cdb, 32'hc00d34d1} /* (19, 0, 16) {real, imag} */,
  {32'h3fea22f4, 32'h3f1b8138} /* (19, 0, 15) {real, imag} */,
  {32'h3e7112b4, 32'hbf3008c5} /* (19, 0, 14) {real, imag} */,
  {32'hbffedce4, 32'hbf7d5a94} /* (19, 0, 13) {real, imag} */,
  {32'hbfd0895a, 32'hbef1c6e8} /* (19, 0, 12) {real, imag} */,
  {32'h4085d3b0, 32'h3fc6840e} /* (19, 0, 11) {real, imag} */,
  {32'hbfa1de18, 32'hc0394282} /* (19, 0, 10) {real, imag} */,
  {32'h4060cd5d, 32'h3e989d7a} /* (19, 0, 9) {real, imag} */,
  {32'hc003ad94, 32'hc01e3624} /* (19, 0, 8) {real, imag} */,
  {32'hbfd7437a, 32'h3e964c45} /* (19, 0, 7) {real, imag} */,
  {32'hbf9868eb, 32'h3f915ec2} /* (19, 0, 6) {real, imag} */,
  {32'hbfb6217e, 32'h3e8caa03} /* (19, 0, 5) {real, imag} */,
  {32'h3ec7640b, 32'hc013245d} /* (19, 0, 4) {real, imag} */,
  {32'h3ecdea9b, 32'h404a69d5} /* (19, 0, 3) {real, imag} */,
  {32'h40023ce4, 32'hbfd673ce} /* (19, 0, 2) {real, imag} */,
  {32'hbff1a0c9, 32'hbee70613} /* (19, 0, 1) {real, imag} */,
  {32'hbe7ff58c, 32'h3d3ae56e} /* (19, 0, 0) {real, imag} */,
  {32'hc0d3b970, 32'h4044ea7d} /* (18, 31, 31) {real, imag} */,
  {32'h40898cca, 32'hbe787ee6} /* (18, 31, 30) {real, imag} */,
  {32'hbeead71e, 32'hbf0af515} /* (18, 31, 29) {real, imag} */,
  {32'hbfabcfbf, 32'hc00f47ad} /* (18, 31, 28) {real, imag} */,
  {32'hbe854b3d, 32'hbe857007} /* (18, 31, 27) {real, imag} */,
  {32'hbf0e2a67, 32'h3fcb2a48} /* (18, 31, 26) {real, imag} */,
  {32'h3f80bc36, 32'hbbaf7bdd} /* (18, 31, 25) {real, imag} */,
  {32'hbf01db57, 32'h3f3b1b7a} /* (18, 31, 24) {real, imag} */,
  {32'h40361ac9, 32'hbeec06b1} /* (18, 31, 23) {real, imag} */,
  {32'h3f8a64eb, 32'hc0272f91} /* (18, 31, 22) {real, imag} */,
  {32'h3f8f9e27, 32'h3f5348fb} /* (18, 31, 21) {real, imag} */,
  {32'hbd1623d0, 32'h3f2b703f} /* (18, 31, 20) {real, imag} */,
  {32'h3fee71a8, 32'h3f610b67} /* (18, 31, 19) {real, imag} */,
  {32'hbfbeef32, 32'hbfc99d5b} /* (18, 31, 18) {real, imag} */,
  {32'hbfdc3ef5, 32'h40004dc3} /* (18, 31, 17) {real, imag} */,
  {32'h3d386da8, 32'h3dbf91e9} /* (18, 31, 16) {real, imag} */,
  {32'h3e7c95c3, 32'h401a0c57} /* (18, 31, 15) {real, imag} */,
  {32'h3edbc00d, 32'h3d99c303} /* (18, 31, 14) {real, imag} */,
  {32'h3f07d063, 32'h3e9e3b29} /* (18, 31, 13) {real, imag} */,
  {32'hbfbfd66d, 32'h3f70eed4} /* (18, 31, 12) {real, imag} */,
  {32'h3fb93fed, 32'hbf962adb} /* (18, 31, 11) {real, imag} */,
  {32'h3f1c49ff, 32'hbf57e0a7} /* (18, 31, 10) {real, imag} */,
  {32'h3f55aff0, 32'h3fdc7844} /* (18, 31, 9) {real, imag} */,
  {32'hc052b399, 32'hbffd2a60} /* (18, 31, 8) {real, imag} */,
  {32'h3f9ebe9e, 32'hbfb81023} /* (18, 31, 7) {real, imag} */,
  {32'h3f023574, 32'h3d3b0fce} /* (18, 31, 6) {real, imag} */,
  {32'h400d61fa, 32'h40511bbc} /* (18, 31, 5) {real, imag} */,
  {32'hbf958401, 32'h3fe1a489} /* (18, 31, 4) {real, imag} */,
  {32'h3efe46a8, 32'h3fa8e31e} /* (18, 31, 3) {real, imag} */,
  {32'h40558d32, 32'h3f99ed72} /* (18, 31, 2) {real, imag} */,
  {32'hc09bfa6e, 32'hc04d330b} /* (18, 31, 1) {real, imag} */,
  {32'hc08991b1, 32'hbf03be47} /* (18, 31, 0) {real, imag} */,
  {32'h3fd90ab7, 32'hbe57653d} /* (18, 30, 31) {real, imag} */,
  {32'hbf65ca1c, 32'hc00343a3} /* (18, 30, 30) {real, imag} */,
  {32'hb980113f, 32'hbfdca0f8} /* (18, 30, 29) {real, imag} */,
  {32'h3f3b11cf, 32'hbf4000c8} /* (18, 30, 28) {real, imag} */,
  {32'h4043cc49, 32'h3feae7d8} /* (18, 30, 27) {real, imag} */,
  {32'h3f02d062, 32'h3f5e4585} /* (18, 30, 26) {real, imag} */,
  {32'h3fa8ab10, 32'hbc7200e1} /* (18, 30, 25) {real, imag} */,
  {32'h3f921ff6, 32'h3de96992} /* (18, 30, 24) {real, imag} */,
  {32'h3feb97d6, 32'hbf50e2de} /* (18, 30, 23) {real, imag} */,
  {32'hc01460fb, 32'hbf81e13a} /* (18, 30, 22) {real, imag} */,
  {32'h3ffde9a3, 32'h400f5c5b} /* (18, 30, 21) {real, imag} */,
  {32'hc03637b0, 32'h3ee5ffbb} /* (18, 30, 20) {real, imag} */,
  {32'h3ead31e1, 32'hc0499a82} /* (18, 30, 19) {real, imag} */,
  {32'hbfb1ad74, 32'h40158fe9} /* (18, 30, 18) {real, imag} */,
  {32'h3fc4c13e, 32'hbf77421c} /* (18, 30, 17) {real, imag} */,
  {32'h3f84611e, 32'h3de2e9c2} /* (18, 30, 16) {real, imag} */,
  {32'h3f4f7f4b, 32'h3eba2678} /* (18, 30, 15) {real, imag} */,
  {32'hbf83f2e8, 32'h401625e0} /* (18, 30, 14) {real, imag} */,
  {32'h3eb6ffd0, 32'h3efae771} /* (18, 30, 13) {real, imag} */,
  {32'hbe30ea3c, 32'h3d4f678c} /* (18, 30, 12) {real, imag} */,
  {32'hbfb91d08, 32'hbfeb14cc} /* (18, 30, 11) {real, imag} */,
  {32'h3fec1a75, 32'hbdaf978f} /* (18, 30, 10) {real, imag} */,
  {32'h3d20d476, 32'hbf6593ce} /* (18, 30, 9) {real, imag} */,
  {32'hbfb4f19a, 32'hc06831e2} /* (18, 30, 8) {real, imag} */,
  {32'hbfbb0830, 32'h3edf0d00} /* (18, 30, 7) {real, imag} */,
  {32'h400ed288, 32'h3e8b9a71} /* (18, 30, 6) {real, imag} */,
  {32'h3f2defeb, 32'hc003f152} /* (18, 30, 5) {real, imag} */,
  {32'h3f6b989a, 32'h3f80336c} /* (18, 30, 4) {real, imag} */,
  {32'h3f523d10, 32'h4005b64e} /* (18, 30, 3) {real, imag} */,
  {32'hc0ac02d5, 32'hc0413826} /* (18, 30, 2) {real, imag} */,
  {32'h40d75171, 32'hbf4b4f32} /* (18, 30, 1) {real, imag} */,
  {32'h40427640, 32'hbf3cb94c} /* (18, 30, 0) {real, imag} */,
  {32'hbf514f08, 32'h3f8b11f1} /* (18, 29, 31) {real, imag} */,
  {32'hbe23e316, 32'h3de64992} /* (18, 29, 30) {real, imag} */,
  {32'h3dc99dcc, 32'h3fb6f636} /* (18, 29, 29) {real, imag} */,
  {32'h4016dfe9, 32'h3f95a515} /* (18, 29, 28) {real, imag} */,
  {32'h3ff46435, 32'h3f30b28d} /* (18, 29, 27) {real, imag} */,
  {32'h3ebcbeb1, 32'hbf2f310a} /* (18, 29, 26) {real, imag} */,
  {32'h3f149048, 32'h3f62b416} /* (18, 29, 25) {real, imag} */,
  {32'h3f4134d6, 32'hbcc56c8f} /* (18, 29, 24) {real, imag} */,
  {32'hbf9a0cab, 32'hbf0985ef} /* (18, 29, 23) {real, imag} */,
  {32'hbb72ea3b, 32'h3ff3d36b} /* (18, 29, 22) {real, imag} */,
  {32'hbf8745e1, 32'hbec5af00} /* (18, 29, 21) {real, imag} */,
  {32'hbfcc8eda, 32'hbfb37c17} /* (18, 29, 20) {real, imag} */,
  {32'hbea44045, 32'hbfdd6bb4} /* (18, 29, 19) {real, imag} */,
  {32'hbf8e51d1, 32'h3ec6b439} /* (18, 29, 18) {real, imag} */,
  {32'h402663e2, 32'hbf7417b7} /* (18, 29, 17) {real, imag} */,
  {32'h3fdd8320, 32'hbdb59e46} /* (18, 29, 16) {real, imag} */,
  {32'hbfc94eec, 32'h3f63cb04} /* (18, 29, 15) {real, imag} */,
  {32'hbfc60700, 32'hbfe81581} /* (18, 29, 14) {real, imag} */,
  {32'h3f38bb48, 32'h3f231307} /* (18, 29, 13) {real, imag} */,
  {32'hbd78826d, 32'h3f82945e} /* (18, 29, 12) {real, imag} */,
  {32'h3fab6233, 32'h3fb117c8} /* (18, 29, 11) {real, imag} */,
  {32'hbf176d5a, 32'hbf7ab9d0} /* (18, 29, 10) {real, imag} */,
  {32'h3fec21aa, 32'h3f93fc4c} /* (18, 29, 9) {real, imag} */,
  {32'h3f7c54b0, 32'h3e83044d} /* (18, 29, 8) {real, imag} */,
  {32'h3ee60668, 32'hc035f507} /* (18, 29, 7) {real, imag} */,
  {32'hbdbf0c83, 32'h3f7ea94c} /* (18, 29, 6) {real, imag} */,
  {32'hbb24c975, 32'h3feaa16c} /* (18, 29, 5) {real, imag} */,
  {32'hbf44abaf, 32'h3f04f7ae} /* (18, 29, 4) {real, imag} */,
  {32'hc04cf2cf, 32'hc0008afb} /* (18, 29, 3) {real, imag} */,
  {32'h3f98d785, 32'hbec769d3} /* (18, 29, 2) {real, imag} */,
  {32'h401532fc, 32'h3feac4e1} /* (18, 29, 1) {real, imag} */,
  {32'h3f5221b7, 32'h3ebaa896} /* (18, 29, 0) {real, imag} */,
  {32'hc08ce35d, 32'hc001837a} /* (18, 28, 31) {real, imag} */,
  {32'h3f2c2b49, 32'hbf14edf5} /* (18, 28, 30) {real, imag} */,
  {32'h3f1a080e, 32'hbe7a406c} /* (18, 28, 29) {real, imag} */,
  {32'h3e65d8dc, 32'h3ead1469} /* (18, 28, 28) {real, imag} */,
  {32'h3feea5f8, 32'h3fbd4399} /* (18, 28, 27) {real, imag} */,
  {32'hbf06c884, 32'h3daddf93} /* (18, 28, 26) {real, imag} */,
  {32'hbf8dd23e, 32'hbfa49d12} /* (18, 28, 25) {real, imag} */,
  {32'h3e607231, 32'hbe227bef} /* (18, 28, 24) {real, imag} */,
  {32'hbf3f9db2, 32'hbe277c17} /* (18, 28, 23) {real, imag} */,
  {32'h40068ba9, 32'hbe3e4860} /* (18, 28, 22) {real, imag} */,
  {32'hc03ab7d1, 32'h3ff1d9da} /* (18, 28, 21) {real, imag} */,
  {32'hbf17b579, 32'hbfb963fd} /* (18, 28, 20) {real, imag} */,
  {32'hbf178568, 32'hbfabcc16} /* (18, 28, 19) {real, imag} */,
  {32'hbef3f528, 32'hbec246ff} /* (18, 28, 18) {real, imag} */,
  {32'h3f8b9b26, 32'h3e234d75} /* (18, 28, 17) {real, imag} */,
  {32'hbe825e60, 32'h3e2373c4} /* (18, 28, 16) {real, imag} */,
  {32'hbda0b828, 32'hbdc47ec7} /* (18, 28, 15) {real, imag} */,
  {32'h3f5d1cbf, 32'hbffba84e} /* (18, 28, 14) {real, imag} */,
  {32'hbf76d3a9, 32'hc02e923a} /* (18, 28, 13) {real, imag} */,
  {32'h4027bdd6, 32'hbfcbe0b8} /* (18, 28, 12) {real, imag} */,
  {32'hbeb714f1, 32'h3f43af9e} /* (18, 28, 11) {real, imag} */,
  {32'h3d9c102f, 32'hbfbfeb01} /* (18, 28, 10) {real, imag} */,
  {32'h3f5c7975, 32'h3d178f7d} /* (18, 28, 9) {real, imag} */,
  {32'h3f9e1247, 32'h3f7a0477} /* (18, 28, 8) {real, imag} */,
  {32'h3f35dd3d, 32'h3f8873f9} /* (18, 28, 7) {real, imag} */,
  {32'h3f366d2f, 32'h3c0cdf0b} /* (18, 28, 6) {real, imag} */,
  {32'hbf504d70, 32'h3fd1d7b1} /* (18, 28, 5) {real, imag} */,
  {32'h3e0c2313, 32'hbee53753} /* (18, 28, 4) {real, imag} */,
  {32'h3f4424d7, 32'h4013f8cc} /* (18, 28, 3) {real, imag} */,
  {32'h3f6a416a, 32'h3fceb700} /* (18, 28, 2) {real, imag} */,
  {32'hbffa3342, 32'h402216a7} /* (18, 28, 1) {real, imag} */,
  {32'h3ef877a9, 32'h3f84a29f} /* (18, 28, 0) {real, imag} */,
  {32'hbe246ae2, 32'hc05fcd2b} /* (18, 27, 31) {real, imag} */,
  {32'hbf002a83, 32'h3efc40b1} /* (18, 27, 30) {real, imag} */,
  {32'hbd11998d, 32'h3f88a7f4} /* (18, 27, 29) {real, imag} */,
  {32'h3ee53edb, 32'hc0055348} /* (18, 27, 28) {real, imag} */,
  {32'h400d63f3, 32'hbfae1619} /* (18, 27, 27) {real, imag} */,
  {32'hbeb3f132, 32'hbf533212} /* (18, 27, 26) {real, imag} */,
  {32'hbe3db293, 32'h3f4d5f0b} /* (18, 27, 25) {real, imag} */,
  {32'hbf3641ff, 32'hbfb899c3} /* (18, 27, 24) {real, imag} */,
  {32'h3fb55b0e, 32'h408003bb} /* (18, 27, 23) {real, imag} */,
  {32'hbf084c5f, 32'hbee7379b} /* (18, 27, 22) {real, imag} */,
  {32'h3fb0c9e9, 32'h3e17d07b} /* (18, 27, 21) {real, imag} */,
  {32'h3fcaae01, 32'hbf80fb22} /* (18, 27, 20) {real, imag} */,
  {32'h3f9c7e73, 32'h3f571ad8} /* (18, 27, 19) {real, imag} */,
  {32'h3ff22bc8, 32'hbf8bdef5} /* (18, 27, 18) {real, imag} */,
  {32'hbfa601ac, 32'hbf7f4e4d} /* (18, 27, 17) {real, imag} */,
  {32'h3ff43fd9, 32'hbfb78c2d} /* (18, 27, 16) {real, imag} */,
  {32'hc02eaa38, 32'h3cc67969} /* (18, 27, 15) {real, imag} */,
  {32'hbffa44be, 32'hbfd5886d} /* (18, 27, 14) {real, imag} */,
  {32'h3fa8bb77, 32'hbfa066ed} /* (18, 27, 13) {real, imag} */,
  {32'hbfce5561, 32'hbf726062} /* (18, 27, 12) {real, imag} */,
  {32'hbfddb845, 32'hbe127d14} /* (18, 27, 11) {real, imag} */,
  {32'hc01155c8, 32'h3fb06b6e} /* (18, 27, 10) {real, imag} */,
  {32'h3faeb454, 32'h3f5fe959} /* (18, 27, 9) {real, imag} */,
  {32'hbf9e43ae, 32'hc0312f5c} /* (18, 27, 8) {real, imag} */,
  {32'h3fd04142, 32'h3fa75ba4} /* (18, 27, 7) {real, imag} */,
  {32'hbdbd1019, 32'hbfb269e7} /* (18, 27, 6) {real, imag} */,
  {32'hc001ee96, 32'hbed00173} /* (18, 27, 5) {real, imag} */,
  {32'h401053be, 32'h3f0e4005} /* (18, 27, 4) {real, imag} */,
  {32'hbf3935fb, 32'hbfaeccb6} /* (18, 27, 3) {real, imag} */,
  {32'hbdd576a4, 32'h401ecd31} /* (18, 27, 2) {real, imag} */,
  {32'hbf398a48, 32'h3f5753ff} /* (18, 27, 1) {real, imag} */,
  {32'h4066416e, 32'hc07a28a6} /* (18, 27, 0) {real, imag} */,
  {32'h3e0cbb17, 32'h3fd71e07} /* (18, 26, 31) {real, imag} */,
  {32'hbe29b2c7, 32'hbf351699} /* (18, 26, 30) {real, imag} */,
  {32'h3fa9ec5d, 32'hbfcacd55} /* (18, 26, 29) {real, imag} */,
  {32'h3f98bb4e, 32'h3fad8d0e} /* (18, 26, 28) {real, imag} */,
  {32'hbf335dd3, 32'h3f6281e1} /* (18, 26, 27) {real, imag} */,
  {32'h3ef066b2, 32'hc000b35b} /* (18, 26, 26) {real, imag} */,
  {32'h3f80ba74, 32'h3fa6adb4} /* (18, 26, 25) {real, imag} */,
  {32'hbf895ecd, 32'h3feabf81} /* (18, 26, 24) {real, imag} */,
  {32'hc0868857, 32'hbfe9ce4a} /* (18, 26, 23) {real, imag} */,
  {32'h3e578ace, 32'hbf99fd3b} /* (18, 26, 22) {real, imag} */,
  {32'hbfedc6d1, 32'hbee60829} /* (18, 26, 21) {real, imag} */,
  {32'hbf6f3bc7, 32'hbede3510} /* (18, 26, 20) {real, imag} */,
  {32'h3e64f96d, 32'hbfdf8c15} /* (18, 26, 19) {real, imag} */,
  {32'hbf49ec6f, 32'h3f8c59fe} /* (18, 26, 18) {real, imag} */,
  {32'h3fad3053, 32'hbfdc3ca6} /* (18, 26, 17) {real, imag} */,
  {32'hbfb3f030, 32'h3f6024b3} /* (18, 26, 16) {real, imag} */,
  {32'h3f7d36e8, 32'h3ebcc1c1} /* (18, 26, 15) {real, imag} */,
  {32'hbf84d1b8, 32'hbee5371a} /* (18, 26, 14) {real, imag} */,
  {32'h3f90d80c, 32'h3ec66b6c} /* (18, 26, 13) {real, imag} */,
  {32'h40027723, 32'h3efa3be7} /* (18, 26, 12) {real, imag} */,
  {32'h3eaa3b2f, 32'hbf873238} /* (18, 26, 11) {real, imag} */,
  {32'hbfa54ed6, 32'h401cc0f3} /* (18, 26, 10) {real, imag} */,
  {32'h3fcfa3c1, 32'hbfcc4791} /* (18, 26, 9) {real, imag} */,
  {32'hbeaa2a60, 32'h3d599590} /* (18, 26, 8) {real, imag} */,
  {32'hbf44e543, 32'h4004b01f} /* (18, 26, 7) {real, imag} */,
  {32'h3fc1dd15, 32'h3eacc719} /* (18, 26, 6) {real, imag} */,
  {32'h3f1f5ea5, 32'hc014e0fc} /* (18, 26, 5) {real, imag} */,
  {32'h3f7b0b17, 32'hbf1c3ac1} /* (18, 26, 4) {real, imag} */,
  {32'hc05245d6, 32'h3fbf0023} /* (18, 26, 3) {real, imag} */,
  {32'h4009e262, 32'hbfc06662} /* (18, 26, 2) {real, imag} */,
  {32'h3f741c49, 32'hbf8706b2} /* (18, 26, 1) {real, imag} */,
  {32'h400db0fb, 32'h3f8bc8a4} /* (18, 26, 0) {real, imag} */,
  {32'hc02ea316, 32'h3fe3709a} /* (18, 25, 31) {real, imag} */,
  {32'h3fe26e94, 32'hbfb1032f} /* (18, 25, 30) {real, imag} */,
  {32'h3fb026f3, 32'hbf398413} /* (18, 25, 29) {real, imag} */,
  {32'h3f65f31e, 32'hc0795d78} /* (18, 25, 28) {real, imag} */,
  {32'h3fb2297c, 32'hbf8d5201} /* (18, 25, 27) {real, imag} */,
  {32'h3fab27c1, 32'hbf7b0c5a} /* (18, 25, 26) {real, imag} */,
  {32'hbee8ee54, 32'h3f0e54c7} /* (18, 25, 25) {real, imag} */,
  {32'hbfa7a6c0, 32'h406b9686} /* (18, 25, 24) {real, imag} */,
  {32'hc0008c1e, 32'h3e9cecaf} /* (18, 25, 23) {real, imag} */,
  {32'h40176105, 32'hc00d3c1b} /* (18, 25, 22) {real, imag} */,
  {32'hbf31474b, 32'h405f84d6} /* (18, 25, 21) {real, imag} */,
  {32'hc0074f6d, 32'hbfbe5848} /* (18, 25, 20) {real, imag} */,
  {32'h3ffa456b, 32'hbd129cf4} /* (18, 25, 19) {real, imag} */,
  {32'hc024eb87, 32'h3f22a373} /* (18, 25, 18) {real, imag} */,
  {32'h3f1a0a51, 32'h3fb776d4} /* (18, 25, 17) {real, imag} */,
  {32'hbe7bf387, 32'h3fb229b4} /* (18, 25, 16) {real, imag} */,
  {32'h3eab22bd, 32'hbdee0b9f} /* (18, 25, 15) {real, imag} */,
  {32'h3d62d9ad, 32'hbf6747a7} /* (18, 25, 14) {real, imag} */,
  {32'hbe8e999b, 32'h3e9f4194} /* (18, 25, 13) {real, imag} */,
  {32'hbf515479, 32'h3f08962a} /* (18, 25, 12) {real, imag} */,
  {32'hbe58e12b, 32'h4019f060} /* (18, 25, 11) {real, imag} */,
  {32'hbf9e62ff, 32'h402201af} /* (18, 25, 10) {real, imag} */,
  {32'hbe8f35d0, 32'hbf719118} /* (18, 25, 9) {real, imag} */,
  {32'h3f7859d9, 32'h3fd178ab} /* (18, 25, 8) {real, imag} */,
  {32'hc01a099f, 32'hbf942947} /* (18, 25, 7) {real, imag} */,
  {32'h3f8ca600, 32'hc0265125} /* (18, 25, 6) {real, imag} */,
  {32'hbfc22866, 32'hbfd6fd9f} /* (18, 25, 5) {real, imag} */,
  {32'h401e4257, 32'h40664093} /* (18, 25, 4) {real, imag} */,
  {32'h3f6a27ad, 32'hbf69266e} /* (18, 25, 3) {real, imag} */,
  {32'hc01f96f7, 32'h3f85d7f5} /* (18, 25, 2) {real, imag} */,
  {32'h3f981c49, 32'h3f43cdfa} /* (18, 25, 1) {real, imag} */,
  {32'hbfa19a10, 32'h3f1b3ac5} /* (18, 25, 0) {real, imag} */,
  {32'h3fd8ea26, 32'h3d14d7d0} /* (18, 24, 31) {real, imag} */,
  {32'h3f791b92, 32'hbe1fe80e} /* (18, 24, 30) {real, imag} */,
  {32'hbe8ee50e, 32'h3f7eb7a4} /* (18, 24, 29) {real, imag} */,
  {32'hbf8bc52d, 32'h3fa51111} /* (18, 24, 28) {real, imag} */,
  {32'hbe688f9c, 32'h3fafe299} /* (18, 24, 27) {real, imag} */,
  {32'hc0099c5a, 32'h3fe98800} /* (18, 24, 26) {real, imag} */,
  {32'hbf00227d, 32'hbea79593} /* (18, 24, 25) {real, imag} */,
  {32'hc03f4f8d, 32'hbf1887e0} /* (18, 24, 24) {real, imag} */,
  {32'hbfb8972c, 32'h4042cdf6} /* (18, 24, 23) {real, imag} */,
  {32'h3f302c78, 32'h3e8becf8} /* (18, 24, 22) {real, imag} */,
  {32'hc081490a, 32'h3edec9b2} /* (18, 24, 21) {real, imag} */,
  {32'hbf5fce37, 32'h3fab5030} /* (18, 24, 20) {real, imag} */,
  {32'hbe58597f, 32'hbffc0592} /* (18, 24, 19) {real, imag} */,
  {32'hbe999326, 32'hbfd54e71} /* (18, 24, 18) {real, imag} */,
  {32'hbf28e34f, 32'h3f836ae5} /* (18, 24, 17) {real, imag} */,
  {32'hc0115996, 32'hbe09ecc3} /* (18, 24, 16) {real, imag} */,
  {32'hbe7cbdeb, 32'h3f09d1a6} /* (18, 24, 15) {real, imag} */,
  {32'h40081720, 32'hbd126184} /* (18, 24, 14) {real, imag} */,
  {32'hbfcda153, 32'hbff2eb7c} /* (18, 24, 13) {real, imag} */,
  {32'h3ff5c34d, 32'h3ffc96f9} /* (18, 24, 12) {real, imag} */,
  {32'hbed9f408, 32'h3ec74ef0} /* (18, 24, 11) {real, imag} */,
  {32'hbfde4df7, 32'h3ffb9d02} /* (18, 24, 10) {real, imag} */,
  {32'hbf99be02, 32'h40257be3} /* (18, 24, 9) {real, imag} */,
  {32'h3ee09548, 32'hbff2f28f} /* (18, 24, 8) {real, imag} */,
  {32'h3fc808fd, 32'h3ff37dfc} /* (18, 24, 7) {real, imag} */,
  {32'h3ff9d10f, 32'hbd2e67dd} /* (18, 24, 6) {real, imag} */,
  {32'h3e56062d, 32'h3fcd0117} /* (18, 24, 5) {real, imag} */,
  {32'hbdfca5a7, 32'hbfe29cf3} /* (18, 24, 4) {real, imag} */,
  {32'hbcf05fdc, 32'h3fe7232d} /* (18, 24, 3) {real, imag} */,
  {32'hbf0b55c6, 32'hbf10120e} /* (18, 24, 2) {real, imag} */,
  {32'h40263b0e, 32'hc03891ed} /* (18, 24, 1) {real, imag} */,
  {32'hbe232ee2, 32'hbe1e30c9} /* (18, 24, 0) {real, imag} */,
  {32'hbf4c83f7, 32'h3fbf7f45} /* (18, 23, 31) {real, imag} */,
  {32'hbebddb34, 32'h3e027193} /* (18, 23, 30) {real, imag} */,
  {32'hbfc8947d, 32'hbe2ff21b} /* (18, 23, 29) {real, imag} */,
  {32'hbfcb4d8f, 32'hbfbe7f6d} /* (18, 23, 28) {real, imag} */,
  {32'h3fac4b67, 32'hbe6bc165} /* (18, 23, 27) {real, imag} */,
  {32'hbf9a15dc, 32'hbcf48009} /* (18, 23, 26) {real, imag} */,
  {32'h3f1c3685, 32'h3f83da8d} /* (18, 23, 25) {real, imag} */,
  {32'h3e14fb4d, 32'hbffdc5ab} /* (18, 23, 24) {real, imag} */,
  {32'hbff0ab16, 32'h3f6ae771} /* (18, 23, 23) {real, imag} */,
  {32'h400aac15, 32'h3f593572} /* (18, 23, 22) {real, imag} */,
  {32'hbe1d8aae, 32'hc03fdb17} /* (18, 23, 21) {real, imag} */,
  {32'hbf13aa48, 32'hc0393fab} /* (18, 23, 20) {real, imag} */,
  {32'hc016cd8d, 32'h3feffa74} /* (18, 23, 19) {real, imag} */,
  {32'h3fc12456, 32'hc0078939} /* (18, 23, 18) {real, imag} */,
  {32'hbe49ed91, 32'h401d5373} /* (18, 23, 17) {real, imag} */,
  {32'h3ffb52fa, 32'h3fec4250} /* (18, 23, 16) {real, imag} */,
  {32'hbfff5631, 32'hbe8a5e67} /* (18, 23, 15) {real, imag} */,
  {32'hbeb1c269, 32'h3f71d3c5} /* (18, 23, 14) {real, imag} */,
  {32'h3f37393d, 32'h3fd180d0} /* (18, 23, 13) {real, imag} */,
  {32'hbf63055a, 32'hbfe82029} /* (18, 23, 12) {real, imag} */,
  {32'hbfd4ce6e, 32'hbf127c9f} /* (18, 23, 11) {real, imag} */,
  {32'h4034ac3e, 32'h3feb6b62} /* (18, 23, 10) {real, imag} */,
  {32'h3f92f6b9, 32'hbe151908} /* (18, 23, 9) {real, imag} */,
  {32'hbe6ad0ed, 32'h3f9f358d} /* (18, 23, 8) {real, imag} */,
  {32'h3f2af826, 32'h3e573b91} /* (18, 23, 7) {real, imag} */,
  {32'h3fc4fc04, 32'h3f7c3527} /* (18, 23, 6) {real, imag} */,
  {32'hc05d1e3e, 32'hbfbe6b75} /* (18, 23, 5) {real, imag} */,
  {32'hc08a7887, 32'h3ff5f75f} /* (18, 23, 4) {real, imag} */,
  {32'hbf6e5df8, 32'hc02ef19a} /* (18, 23, 3) {real, imag} */,
  {32'h3fca9fdf, 32'h3f6dc5b3} /* (18, 23, 2) {real, imag} */,
  {32'h40019da6, 32'h3f82826b} /* (18, 23, 1) {real, imag} */,
  {32'h3f7a8384, 32'h3fa368b9} /* (18, 23, 0) {real, imag} */,
  {32'hc004c24c, 32'hc0381a9d} /* (18, 22, 31) {real, imag} */,
  {32'hc0024e07, 32'h3c5bbc6b} /* (18, 22, 30) {real, imag} */,
  {32'hba614f0d, 32'hbf1981e1} /* (18, 22, 29) {real, imag} */,
  {32'h3e59bef5, 32'h40085a25} /* (18, 22, 28) {real, imag} */,
  {32'h3f09824c, 32'hbee1444f} /* (18, 22, 27) {real, imag} */,
  {32'h3fc659a3, 32'h3f5d7cbe} /* (18, 22, 26) {real, imag} */,
  {32'h4005b5ed, 32'hbf0b3f53} /* (18, 22, 25) {real, imag} */,
  {32'hbfbfe9cd, 32'h3f291346} /* (18, 22, 24) {real, imag} */,
  {32'h3e4ec128, 32'h3ec861e8} /* (18, 22, 23) {real, imag} */,
  {32'h407d84bf, 32'hbf18359d} /* (18, 22, 22) {real, imag} */,
  {32'h3fbcca73, 32'hbf48899d} /* (18, 22, 21) {real, imag} */,
  {32'h3e3dcde6, 32'h3fc0fa02} /* (18, 22, 20) {real, imag} */,
  {32'hbff119ca, 32'h40a69ace} /* (18, 22, 19) {real, imag} */,
  {32'hc00a61a0, 32'hc03a9329} /* (18, 22, 18) {real, imag} */,
  {32'h3f50a9bb, 32'h3fb8b5f1} /* (18, 22, 17) {real, imag} */,
  {32'hc04c49a8, 32'h3f09c0cd} /* (18, 22, 16) {real, imag} */,
  {32'hc0423759, 32'hbfb3cc64} /* (18, 22, 15) {real, imag} */,
  {32'hbe172c1c, 32'h40040cf2} /* (18, 22, 14) {real, imag} */,
  {32'h404fb919, 32'h3fbd0b17} /* (18, 22, 13) {real, imag} */,
  {32'h3f2c3df7, 32'hbfbbf155} /* (18, 22, 12) {real, imag} */,
  {32'hbe17f8f4, 32'h4009e654} /* (18, 22, 11) {real, imag} */,
  {32'hc003228c, 32'h40458191} /* (18, 22, 10) {real, imag} */,
  {32'hbf0190b7, 32'h3f0097c8} /* (18, 22, 9) {real, imag} */,
  {32'hbe85258e, 32'hbd0d21dc} /* (18, 22, 8) {real, imag} */,
  {32'h3e81e079, 32'hbe532327} /* (18, 22, 7) {real, imag} */,
  {32'h4095ff39, 32'hbf06cd2e} /* (18, 22, 6) {real, imag} */,
  {32'h3bbaa991, 32'hbf4fd0ab} /* (18, 22, 5) {real, imag} */,
  {32'hbf307d0b, 32'hbf32660e} /* (18, 22, 4) {real, imag} */,
  {32'hbf7b3299, 32'h3c982cb9} /* (18, 22, 3) {real, imag} */,
  {32'h402167fa, 32'hbfbd558c} /* (18, 22, 2) {real, imag} */,
  {32'hbf267017, 32'h3fb14fd8} /* (18, 22, 1) {real, imag} */,
  {32'h401396b3, 32'h3e047c3c} /* (18, 22, 0) {real, imag} */,
  {32'h3d8c16d3, 32'h3cf3e7f6} /* (18, 21, 31) {real, imag} */,
  {32'hbf9eafeb, 32'h403e80ca} /* (18, 21, 30) {real, imag} */,
  {32'hbe1f91b3, 32'h3ffa2b4d} /* (18, 21, 29) {real, imag} */,
  {32'hbfa2ba31, 32'h401ae27f} /* (18, 21, 28) {real, imag} */,
  {32'hbf9df577, 32'h3e43ae0c} /* (18, 21, 27) {real, imag} */,
  {32'h401eda7e, 32'hbeb8cd7a} /* (18, 21, 26) {real, imag} */,
  {32'h3fbeb044, 32'hbf26e553} /* (18, 21, 25) {real, imag} */,
  {32'h400931dd, 32'hc01c4fb3} /* (18, 21, 24) {real, imag} */,
  {32'hbea51d58, 32'hbf4b51d1} /* (18, 21, 23) {real, imag} */,
  {32'hbe182785, 32'h3edf6d29} /* (18, 21, 22) {real, imag} */,
  {32'h4086ffd9, 32'h3f79131b} /* (18, 21, 21) {real, imag} */,
  {32'h3f2f1b1c, 32'hbf27ecc9} /* (18, 21, 20) {real, imag} */,
  {32'h3fb354ff, 32'h4038dc40} /* (18, 21, 19) {real, imag} */,
  {32'h3f827e22, 32'h3fe46ab0} /* (18, 21, 18) {real, imag} */,
  {32'hbfce7000, 32'h3f9ff7c2} /* (18, 21, 17) {real, imag} */,
  {32'hc003979d, 32'hc04653c8} /* (18, 21, 16) {real, imag} */,
  {32'hbf4ab750, 32'h407aa1d3} /* (18, 21, 15) {real, imag} */,
  {32'h3f657f5c, 32'hc0161928} /* (18, 21, 14) {real, imag} */,
  {32'hbf353aa5, 32'hc0845ef1} /* (18, 21, 13) {real, imag} */,
  {32'h3f424d8d, 32'hc01ad640} /* (18, 21, 12) {real, imag} */,
  {32'h3fadb7b4, 32'h3fdbe64b} /* (18, 21, 11) {real, imag} */,
  {32'h3f2b8ecc, 32'h3ec2ccc9} /* (18, 21, 10) {real, imag} */,
  {32'hbe034ce1, 32'h3fd90143} /* (18, 21, 9) {real, imag} */,
  {32'h3ed40961, 32'hc00203f4} /* (18, 21, 8) {real, imag} */,
  {32'hbf2eef27, 32'hbfd47cd1} /* (18, 21, 7) {real, imag} */,
  {32'hbf8c8d7f, 32'h3f29f1bd} /* (18, 21, 6) {real, imag} */,
  {32'h3f64db9e, 32'hc02edd1b} /* (18, 21, 5) {real, imag} */,
  {32'h3eab734b, 32'h3fb855bf} /* (18, 21, 4) {real, imag} */,
  {32'h4009c3d8, 32'hbf6de63c} /* (18, 21, 3) {real, imag} */,
  {32'hbe65c16c, 32'h3f3b7570} /* (18, 21, 2) {real, imag} */,
  {32'hbf36f32f, 32'hbf5dc943} /* (18, 21, 1) {real, imag} */,
  {32'hbd8a83c6, 32'hbf9a7a33} /* (18, 21, 0) {real, imag} */,
  {32'h3f6e5381, 32'h3fc547c2} /* (18, 20, 31) {real, imag} */,
  {32'hbe69f9cc, 32'h3fb3b7e1} /* (18, 20, 30) {real, imag} */,
  {32'h3eeb56f8, 32'h3ebe1422} /* (18, 20, 29) {real, imag} */,
  {32'h3fef4657, 32'hbdef05e5} /* (18, 20, 28) {real, imag} */,
  {32'hc00c0bbf, 32'hbdd1f7ed} /* (18, 20, 27) {real, imag} */,
  {32'h3e1c59e6, 32'h3f9eef3c} /* (18, 20, 26) {real, imag} */,
  {32'h3fa820a7, 32'h3fd36f33} /* (18, 20, 25) {real, imag} */,
  {32'hc07eadad, 32'h3f8ef92b} /* (18, 20, 24) {real, imag} */,
  {32'hbf854ce4, 32'hbe2d9eae} /* (18, 20, 23) {real, imag} */,
  {32'h40885007, 32'h3f583995} /* (18, 20, 22) {real, imag} */,
  {32'hbfc0b2d9, 32'hc010ef99} /* (18, 20, 21) {real, imag} */,
  {32'h3f288079, 32'hbf42ae02} /* (18, 20, 20) {real, imag} */,
  {32'hbf9c8e8e, 32'h3e53ee4f} /* (18, 20, 19) {real, imag} */,
  {32'hbf9c5943, 32'h40969592} /* (18, 20, 18) {real, imag} */,
  {32'hc026191b, 32'hbfe31f6b} /* (18, 20, 17) {real, imag} */,
  {32'hbd66da48, 32'hbfe7ab46} /* (18, 20, 16) {real, imag} */,
  {32'hbe60bcd3, 32'hbe66f59a} /* (18, 20, 15) {real, imag} */,
  {32'h3f20de66, 32'h3e8c6c3d} /* (18, 20, 14) {real, imag} */,
  {32'hbf4f6896, 32'h3ed90862} /* (18, 20, 13) {real, imag} */,
  {32'hc02418fe, 32'hbfac6c28} /* (18, 20, 12) {real, imag} */,
  {32'h3f397ab4, 32'h3fd0cfec} /* (18, 20, 11) {real, imag} */,
  {32'h3f5b5715, 32'h4017a4d3} /* (18, 20, 10) {real, imag} */,
  {32'h3f92669a, 32'hc018e40d} /* (18, 20, 9) {real, imag} */,
  {32'h3f161995, 32'hbf85b3f1} /* (18, 20, 8) {real, imag} */,
  {32'h3f9951bc, 32'h3d147233} /* (18, 20, 7) {real, imag} */,
  {32'hbf95b239, 32'hbfeaef01} /* (18, 20, 6) {real, imag} */,
  {32'h40181399, 32'hbe80898d} /* (18, 20, 5) {real, imag} */,
  {32'h3fad269d, 32'hc0810a9d} /* (18, 20, 4) {real, imag} */,
  {32'hc0697cac, 32'h3f9580cd} /* (18, 20, 3) {real, imag} */,
  {32'hbfb3ae27, 32'h3e137bd4} /* (18, 20, 2) {real, imag} */,
  {32'hbf78086c, 32'h3f9848c1} /* (18, 20, 1) {real, imag} */,
  {32'hbe6051aa, 32'h4053b23b} /* (18, 20, 0) {real, imag} */,
  {32'h3f094f20, 32'h3d86002c} /* (18, 19, 31) {real, imag} */,
  {32'hbeb11214, 32'hc0148061} /* (18, 19, 30) {real, imag} */,
  {32'hbf61fd27, 32'hbf9eb666} /* (18, 19, 29) {real, imag} */,
  {32'hbd12dc8e, 32'hbf579859} /* (18, 19, 28) {real, imag} */,
  {32'h3fc251ce, 32'h3fa32a23} /* (18, 19, 27) {real, imag} */,
  {32'hbfdcd479, 32'h3f215909} /* (18, 19, 26) {real, imag} */,
  {32'hc035c2e4, 32'h3eac0c6c} /* (18, 19, 25) {real, imag} */,
  {32'hbfe70b99, 32'h3f7928fd} /* (18, 19, 24) {real, imag} */,
  {32'hbea17c42, 32'hc04f3b60} /* (18, 19, 23) {real, imag} */,
  {32'hbfbda832, 32'h3e7546aa} /* (18, 19, 22) {real, imag} */,
  {32'h3f113551, 32'h3fabe13c} /* (18, 19, 21) {real, imag} */,
  {32'h4067c4b5, 32'h3f033f9c} /* (18, 19, 20) {real, imag} */,
  {32'h4010b4e9, 32'h4047921c} /* (18, 19, 19) {real, imag} */,
  {32'hbfa0edc0, 32'hbf421174} /* (18, 19, 18) {real, imag} */,
  {32'h3ff6fec7, 32'hbf140633} /* (18, 19, 17) {real, imag} */,
  {32'hbf0ed44d, 32'h3e90eb96} /* (18, 19, 16) {real, imag} */,
  {32'hbf832404, 32'hc01c60bc} /* (18, 19, 15) {real, imag} */,
  {32'h3e9d2a62, 32'hbf45f0e6} /* (18, 19, 14) {real, imag} */,
  {32'h3df6b70f, 32'h3f0d42fc} /* (18, 19, 13) {real, imag} */,
  {32'h401ee7c6, 32'h3ff23b7f} /* (18, 19, 12) {real, imag} */,
  {32'hc0079e30, 32'hbf9549bc} /* (18, 19, 11) {real, imag} */,
  {32'h406b583a, 32'h3fe019dc} /* (18, 19, 10) {real, imag} */,
  {32'hbed70a20, 32'hc0899333} /* (18, 19, 9) {real, imag} */,
  {32'hc0202a56, 32'hbdb873ef} /* (18, 19, 8) {real, imag} */,
  {32'h3fe89112, 32'h3fb9dda3} /* (18, 19, 7) {real, imag} */,
  {32'hbf988220, 32'h400cb3a7} /* (18, 19, 6) {real, imag} */,
  {32'h3f6b71e2, 32'hbf0aa162} /* (18, 19, 5) {real, imag} */,
  {32'h3dfd3612, 32'h3fa82269} /* (18, 19, 4) {real, imag} */,
  {32'hbefd8afe, 32'h3dcf3266} /* (18, 19, 3) {real, imag} */,
  {32'h3fde86b1, 32'hbff30754} /* (18, 19, 2) {real, imag} */,
  {32'h3f385e0d, 32'h3da42ae1} /* (18, 19, 1) {real, imag} */,
  {32'hc062458e, 32'h3f89a6e8} /* (18, 19, 0) {real, imag} */,
  {32'h3f58f2ed, 32'h3f1a8d91} /* (18, 18, 31) {real, imag} */,
  {32'h3f3f5514, 32'hbe8c4fd5} /* (18, 18, 30) {real, imag} */,
  {32'hbf81023a, 32'h3faadb91} /* (18, 18, 29) {real, imag} */,
  {32'hbf534bd9, 32'hbfe19a1e} /* (18, 18, 28) {real, imag} */,
  {32'h3f138d90, 32'h3f84f39a} /* (18, 18, 27) {real, imag} */,
  {32'h403503c6, 32'hbf807330} /* (18, 18, 26) {real, imag} */,
  {32'hbf3245fd, 32'h3f7a93c0} /* (18, 18, 25) {real, imag} */,
  {32'hc01f8691, 32'hbf370cf6} /* (18, 18, 24) {real, imag} */,
  {32'h3e70a583, 32'hc0710eda} /* (18, 18, 23) {real, imag} */,
  {32'h3e57f7ec, 32'hbf0bb0e9} /* (18, 18, 22) {real, imag} */,
  {32'h400a13e5, 32'h3fd17df6} /* (18, 18, 21) {real, imag} */,
  {32'h3f0e3cf2, 32'h3f9130cd} /* (18, 18, 20) {real, imag} */,
  {32'h3fa15b45, 32'h4041b9b1} /* (18, 18, 19) {real, imag} */,
  {32'hbe8964a5, 32'h3fc66ce5} /* (18, 18, 18) {real, imag} */,
  {32'h3e8a5624, 32'h3f1cc200} /* (18, 18, 17) {real, imag} */,
  {32'hbf27525e, 32'h3ff6d98e} /* (18, 18, 16) {real, imag} */,
  {32'h3f45dd1e, 32'hbf8985d9} /* (18, 18, 15) {real, imag} */,
  {32'h3fe3425d, 32'hbf5f9600} /* (18, 18, 14) {real, imag} */,
  {32'h3e133717, 32'hbf4eae4f} /* (18, 18, 13) {real, imag} */,
  {32'hbf1c9fb0, 32'h40011038} /* (18, 18, 12) {real, imag} */,
  {32'h3fc298b1, 32'h3e8ecee2} /* (18, 18, 11) {real, imag} */,
  {32'hbf58954a, 32'hbe62f968} /* (18, 18, 10) {real, imag} */,
  {32'hbfe815fc, 32'h4055a19f} /* (18, 18, 9) {real, imag} */,
  {32'h3feec533, 32'h3fa9eeb2} /* (18, 18, 8) {real, imag} */,
  {32'hbf078ac4, 32'h3ae048cd} /* (18, 18, 7) {real, imag} */,
  {32'h3ee175be, 32'h3fe12760} /* (18, 18, 6) {real, imag} */,
  {32'h4031420c, 32'hc000c7a3} /* (18, 18, 5) {real, imag} */,
  {32'h3f2f675f, 32'h3e8b4d10} /* (18, 18, 4) {real, imag} */,
  {32'hbe87f262, 32'hbf1a2ac5} /* (18, 18, 3) {real, imag} */,
  {32'hbef109aa, 32'h3fcfe955} /* (18, 18, 2) {real, imag} */,
  {32'h3db4b031, 32'hbf948356} /* (18, 18, 1) {real, imag} */,
  {32'hbd8cf1a1, 32'h3e1e999f} /* (18, 18, 0) {real, imag} */,
  {32'h3fa64cee, 32'h3f1982f1} /* (18, 17, 31) {real, imag} */,
  {32'h3e8d252e, 32'hc01200c8} /* (18, 17, 30) {real, imag} */,
  {32'h3f26fd54, 32'hbe679da7} /* (18, 17, 29) {real, imag} */,
  {32'h3f9e89a6, 32'hbfd7d600} /* (18, 17, 28) {real, imag} */,
  {32'hbebe1fcb, 32'h3e48df82} /* (18, 17, 27) {real, imag} */,
  {32'h401466f6, 32'h3ff22070} /* (18, 17, 26) {real, imag} */,
  {32'h3f4bab99, 32'h3d2e1abf} /* (18, 17, 25) {real, imag} */,
  {32'hbeff0a7f, 32'hc04fbf86} /* (18, 17, 24) {real, imag} */,
  {32'h3f58dd14, 32'h3e775b8d} /* (18, 17, 23) {real, imag} */,
  {32'h3fc0d96b, 32'h3e60f8db} /* (18, 17, 22) {real, imag} */,
  {32'hbfe788d8, 32'h402aa2a3} /* (18, 17, 21) {real, imag} */,
  {32'hbfd4c7b2, 32'h3e4e03be} /* (18, 17, 20) {real, imag} */,
  {32'hbffc3c23, 32'hc02172e6} /* (18, 17, 19) {real, imag} */,
  {32'h3f6c6a91, 32'h4011188f} /* (18, 17, 18) {real, imag} */,
  {32'h3f7490b2, 32'h3fb08eef} /* (18, 17, 17) {real, imag} */,
  {32'hbe9dbf05, 32'h400e840d} /* (18, 17, 16) {real, imag} */,
  {32'h3e590001, 32'hbeeb3180} /* (18, 17, 15) {real, imag} */,
  {32'h3ec7d260, 32'hbe710a51} /* (18, 17, 14) {real, imag} */,
  {32'hbfb75ece, 32'hbf4c2615} /* (18, 17, 13) {real, imag} */,
  {32'h3eac0723, 32'h3f985685} /* (18, 17, 12) {real, imag} */,
  {32'h3fed1062, 32'hbfe36b19} /* (18, 17, 11) {real, imag} */,
  {32'h403214b1, 32'h400d01a3} /* (18, 17, 10) {real, imag} */,
  {32'hbeda0937, 32'hbfb72050} /* (18, 17, 9) {real, imag} */,
  {32'hbfaf0778, 32'h3f74226b} /* (18, 17, 8) {real, imag} */,
  {32'h3f3c2923, 32'hbf54d46f} /* (18, 17, 7) {real, imag} */,
  {32'hbfa3fc1c, 32'hbec698d4} /* (18, 17, 6) {real, imag} */,
  {32'h3f6b07e4, 32'h3e6c8fe6} /* (18, 17, 5) {real, imag} */,
  {32'hbfe7146e, 32'hbe107643} /* (18, 17, 4) {real, imag} */,
  {32'h3fb0f17d, 32'h3f90cc4f} /* (18, 17, 3) {real, imag} */,
  {32'h3caf2f6e, 32'h3e8f3e45} /* (18, 17, 2) {real, imag} */,
  {32'hbf5f6e48, 32'h40082c39} /* (18, 17, 1) {real, imag} */,
  {32'hbfe197d9, 32'h3f486185} /* (18, 17, 0) {real, imag} */,
  {32'h3e11f954, 32'h401a63ef} /* (18, 16, 31) {real, imag} */,
  {32'hbf8e311a, 32'hbfea6114} /* (18, 16, 30) {real, imag} */,
  {32'h3f4a98a2, 32'h3f17edab} /* (18, 16, 29) {real, imag} */,
  {32'h3f2c963d, 32'hbd69c942} /* (18, 16, 28) {real, imag} */,
  {32'h3fabfea1, 32'hbf8a90d3} /* (18, 16, 27) {real, imag} */,
  {32'hbe3e1168, 32'hbf0d9ea1} /* (18, 16, 26) {real, imag} */,
  {32'hbf02412e, 32'h3e9019c9} /* (18, 16, 25) {real, imag} */,
  {32'hbedd48f0, 32'hbee649c6} /* (18, 16, 24) {real, imag} */,
  {32'h3eb46a87, 32'h3f72180f} /* (18, 16, 23) {real, imag} */,
  {32'hbe5914c3, 32'h405901c4} /* (18, 16, 22) {real, imag} */,
  {32'hbef1ac77, 32'h3dadd828} /* (18, 16, 21) {real, imag} */,
  {32'h3f4d2559, 32'hbf0b62de} /* (18, 16, 20) {real, imag} */,
  {32'hbfb71ac9, 32'h3f5fe7db} /* (18, 16, 19) {real, imag} */,
  {32'h3f0d301f, 32'h3ef8ead5} /* (18, 16, 18) {real, imag} */,
  {32'h3d9fcff8, 32'hbee6d48a} /* (18, 16, 17) {real, imag} */,
  {32'h3dbbde8d, 32'h3f464312} /* (18, 16, 16) {real, imag} */,
  {32'hbe6656c2, 32'h3eb6d73c} /* (18, 16, 15) {real, imag} */,
  {32'hbfd37524, 32'hbfa5bf81} /* (18, 16, 14) {real, imag} */,
  {32'h3ff182cd, 32'hc0020e37} /* (18, 16, 13) {real, imag} */,
  {32'h3fa9e4c2, 32'hbd9cd32a} /* (18, 16, 12) {real, imag} */,
  {32'hbd7d0712, 32'h3eb870fe} /* (18, 16, 11) {real, imag} */,
  {32'h3f6d77bf, 32'h3fa84976} /* (18, 16, 10) {real, imag} */,
  {32'h3f8578be, 32'hbf7c4d6a} /* (18, 16, 9) {real, imag} */,
  {32'hbf426a4b, 32'h3f1eded6} /* (18, 16, 8) {real, imag} */,
  {32'h3f83af5e, 32'h3fb15bb5} /* (18, 16, 7) {real, imag} */,
  {32'hbfb59547, 32'hbfa39ff0} /* (18, 16, 6) {real, imag} */,
  {32'hbec58124, 32'hbf890f4a} /* (18, 16, 5) {real, imag} */,
  {32'h3f5ef34b, 32'hbf88c775} /* (18, 16, 4) {real, imag} */,
  {32'hbed63e41, 32'h3f3b24c0} /* (18, 16, 3) {real, imag} */,
  {32'hbf072aff, 32'h3f48558c} /* (18, 16, 2) {real, imag} */,
  {32'hbf03a6dd, 32'hbdedb29f} /* (18, 16, 1) {real, imag} */,
  {32'h3ed49494, 32'hbea8fb26} /* (18, 16, 0) {real, imag} */,
  {32'h3ef0f618, 32'h3ee8b31d} /* (18, 15, 31) {real, imag} */,
  {32'h3f1cc71a, 32'hbf2926f8} /* (18, 15, 30) {real, imag} */,
  {32'h3fff0af1, 32'h3e8ca0d1} /* (18, 15, 29) {real, imag} */,
  {32'h3f43b80a, 32'h40365a70} /* (18, 15, 28) {real, imag} */,
  {32'hbd8e4fd8, 32'hbf1a3193} /* (18, 15, 27) {real, imag} */,
  {32'h3f84ec83, 32'hc0272f75} /* (18, 15, 26) {real, imag} */,
  {32'hbfd7bcaf, 32'hbe5a3b65} /* (18, 15, 25) {real, imag} */,
  {32'h3f6e60ad, 32'hbfb4ce6b} /* (18, 15, 24) {real, imag} */,
  {32'h3f39a58a, 32'hbf960b58} /* (18, 15, 23) {real, imag} */,
  {32'h3fd22c39, 32'h3fb43836} /* (18, 15, 22) {real, imag} */,
  {32'hbfb0559d, 32'h3d16d2ec} /* (18, 15, 21) {real, imag} */,
  {32'hbf8782f4, 32'h3f8d7d00} /* (18, 15, 20) {real, imag} */,
  {32'hbf6c90e4, 32'hc032b94a} /* (18, 15, 19) {real, imag} */,
  {32'h3f5b4391, 32'hbecc9cce} /* (18, 15, 18) {real, imag} */,
  {32'hbf177b39, 32'h3fadc64f} /* (18, 15, 17) {real, imag} */,
  {32'h3f07586a, 32'hbf82c1fc} /* (18, 15, 16) {real, imag} */,
  {32'hc00b7dd9, 32'hbf7eb10b} /* (18, 15, 15) {real, imag} */,
  {32'hc0063375, 32'hc03ad93e} /* (18, 15, 14) {real, imag} */,
  {32'hbfef74ed, 32'h3e534d13} /* (18, 15, 13) {real, imag} */,
  {32'hbf8d122b, 32'hc0a1b7cd} /* (18, 15, 12) {real, imag} */,
  {32'hbfe1c515, 32'hbf7c51a8} /* (18, 15, 11) {real, imag} */,
  {32'h404450bf, 32'h3ebd4c3d} /* (18, 15, 10) {real, imag} */,
  {32'h40246d28, 32'h3fbd039a} /* (18, 15, 9) {real, imag} */,
  {32'h3f47bf98, 32'h3f45cd01} /* (18, 15, 8) {real, imag} */,
  {32'hbf95d5dd, 32'hbf959a77} /* (18, 15, 7) {real, imag} */,
  {32'hbf15e6bf, 32'hbd6a4dbb} /* (18, 15, 6) {real, imag} */,
  {32'h3eea52bb, 32'h3f5677e5} /* (18, 15, 5) {real, imag} */,
  {32'hbfbbdd4b, 32'h3f5f10ca} /* (18, 15, 4) {real, imag} */,
  {32'h3f323739, 32'h3e87fdfd} /* (18, 15, 3) {real, imag} */,
  {32'hbf576529, 32'h3f12a7c3} /* (18, 15, 2) {real, imag} */,
  {32'hbfb60dbd, 32'hbe6bf1cf} /* (18, 15, 1) {real, imag} */,
  {32'h3f0541e6, 32'h3e1d72f8} /* (18, 15, 0) {real, imag} */,
  {32'hbde11275, 32'h3fdf079e} /* (18, 14, 31) {real, imag} */,
  {32'h3f8a3318, 32'h3f216cdb} /* (18, 14, 30) {real, imag} */,
  {32'hbf4260d3, 32'h3f84f40c} /* (18, 14, 29) {real, imag} */,
  {32'h40274549, 32'h3f521645} /* (18, 14, 28) {real, imag} */,
  {32'hbf32a698, 32'hbcfabfb0} /* (18, 14, 27) {real, imag} */,
  {32'hbfc5d1ed, 32'h3f362b77} /* (18, 14, 26) {real, imag} */,
  {32'hbfbc2ad3, 32'h3ecfe114} /* (18, 14, 25) {real, imag} */,
  {32'hbe41bcb6, 32'hbf161530} /* (18, 14, 24) {real, imag} */,
  {32'hbfceb65f, 32'h3e322770} /* (18, 14, 23) {real, imag} */,
  {32'hc026ade1, 32'hbf09edfb} /* (18, 14, 22) {real, imag} */,
  {32'hbf04c868, 32'hc02365a1} /* (18, 14, 21) {real, imag} */,
  {32'hc02cfb50, 32'hc02518e2} /* (18, 14, 20) {real, imag} */,
  {32'hc0507069, 32'h400f9dd8} /* (18, 14, 19) {real, imag} */,
  {32'hbfc686a2, 32'hbf6a505e} /* (18, 14, 18) {real, imag} */,
  {32'h3f5c4240, 32'hbf3f7537} /* (18, 14, 17) {real, imag} */,
  {32'h3fb6a584, 32'hbe963dc6} /* (18, 14, 16) {real, imag} */,
  {32'h3ef3e47a, 32'h3f811ae3} /* (18, 14, 15) {real, imag} */,
  {32'h3ef3b773, 32'h3f12afde} /* (18, 14, 14) {real, imag} */,
  {32'h3fe19ce5, 32'hc02a94a0} /* (18, 14, 13) {real, imag} */,
  {32'h3fd1118c, 32'h402dc919} /* (18, 14, 12) {real, imag} */,
  {32'h400c2994, 32'h3e203568} /* (18, 14, 11) {real, imag} */,
  {32'h4063fc87, 32'hbeadc08b} /* (18, 14, 10) {real, imag} */,
  {32'hc07882b6, 32'hc02e269a} /* (18, 14, 9) {real, imag} */,
  {32'h3f09ddee, 32'h3f296cff} /* (18, 14, 8) {real, imag} */,
  {32'h400e5de7, 32'h3f824f8e} /* (18, 14, 7) {real, imag} */,
  {32'h3f4dcd45, 32'h3ea6787f} /* (18, 14, 6) {real, imag} */,
  {32'h3e400aa6, 32'hc0035be6} /* (18, 14, 5) {real, imag} */,
  {32'hbe8d3c34, 32'h3f4a5422} /* (18, 14, 4) {real, imag} */,
  {32'h3e450a0c, 32'hbff6d351} /* (18, 14, 3) {real, imag} */,
  {32'h3e26f9a2, 32'hbf16b42e} /* (18, 14, 2) {real, imag} */,
  {32'h3e17d4e6, 32'h3f907715} /* (18, 14, 1) {real, imag} */,
  {32'hbf01228a, 32'h3f08ae7b} /* (18, 14, 0) {real, imag} */,
  {32'hbff3d768, 32'h3f2ede0c} /* (18, 13, 31) {real, imag} */,
  {32'hbeb32683, 32'hbbddffcc} /* (18, 13, 30) {real, imag} */,
  {32'h3f805452, 32'h3f395b9d} /* (18, 13, 29) {real, imag} */,
  {32'h3e3bd225, 32'hbf9a90f0} /* (18, 13, 28) {real, imag} */,
  {32'hbf1f78ca, 32'hbfb118a4} /* (18, 13, 27) {real, imag} */,
  {32'h3fd016fa, 32'hbfda72bc} /* (18, 13, 26) {real, imag} */,
  {32'hbfdd94fb, 32'h3fc638e0} /* (18, 13, 25) {real, imag} */,
  {32'hbf32a31e, 32'hbfc09f08} /* (18, 13, 24) {real, imag} */,
  {32'h3d8c2b2c, 32'hbf3d9c91} /* (18, 13, 23) {real, imag} */,
  {32'h3f6ee650, 32'h3d4f1177} /* (18, 13, 22) {real, imag} */,
  {32'hbe2f9bbd, 32'hbff828d2} /* (18, 13, 21) {real, imag} */,
  {32'hbf161f8e, 32'h3dee962e} /* (18, 13, 20) {real, imag} */,
  {32'hc034ed86, 32'hbefbef07} /* (18, 13, 19) {real, imag} */,
  {32'hbff9a52c, 32'h3ebeca9e} /* (18, 13, 18) {real, imag} */,
  {32'h3f89af47, 32'h3f6b9d69} /* (18, 13, 17) {real, imag} */,
  {32'hbfebf84e, 32'hbf82f440} /* (18, 13, 16) {real, imag} */,
  {32'h3f8a2e70, 32'hbe414f59} /* (18, 13, 15) {real, imag} */,
  {32'h4024d21b, 32'h3fadf3f9} /* (18, 13, 14) {real, imag} */,
  {32'h400403eb, 32'h3f2c7d69} /* (18, 13, 13) {real, imag} */,
  {32'hc03ef542, 32'h400b5aeb} /* (18, 13, 12) {real, imag} */,
  {32'hc00ba7fa, 32'h3f6a5c07} /* (18, 13, 11) {real, imag} */,
  {32'h3ee04eb6, 32'h3fea3553} /* (18, 13, 10) {real, imag} */,
  {32'h3f007dd5, 32'hbff27535} /* (18, 13, 9) {real, imag} */,
  {32'h400394b3, 32'h4007eecb} /* (18, 13, 8) {real, imag} */,
  {32'hbfac1801, 32'h3ed99ffb} /* (18, 13, 7) {real, imag} */,
  {32'hc023c6e3, 32'h4029bdf6} /* (18, 13, 6) {real, imag} */,
  {32'h3f27a967, 32'h3fe0372a} /* (18, 13, 5) {real, imag} */,
  {32'h3fb27894, 32'h3ebc306e} /* (18, 13, 4) {real, imag} */,
  {32'hbfec6bfa, 32'h4003b1e2} /* (18, 13, 3) {real, imag} */,
  {32'hc000f17d, 32'h3cf480f1} /* (18, 13, 2) {real, imag} */,
  {32'h3f60f38c, 32'hbf9c2014} /* (18, 13, 1) {real, imag} */,
  {32'hbff547f6, 32'hbfe55025} /* (18, 13, 0) {real, imag} */,
  {32'h3f33b336, 32'h3f76d34c} /* (18, 12, 31) {real, imag} */,
  {32'hbfc36013, 32'hbf2365a3} /* (18, 12, 30) {real, imag} */,
  {32'h3fc635b0, 32'h3e81655e} /* (18, 12, 29) {real, imag} */,
  {32'hc02d08e6, 32'hbfc1468b} /* (18, 12, 28) {real, imag} */,
  {32'hbfb4bcbf, 32'hc01951c4} /* (18, 12, 27) {real, imag} */,
  {32'h3e35034a, 32'hbe310f4f} /* (18, 12, 26) {real, imag} */,
  {32'h401c04af, 32'hc023f99c} /* (18, 12, 25) {real, imag} */,
  {32'h4020b955, 32'hbcc04e8d} /* (18, 12, 24) {real, imag} */,
  {32'h3fb8e4b2, 32'h400c2a19} /* (18, 12, 23) {real, imag} */,
  {32'hc0517044, 32'hc04e6652} /* (18, 12, 22) {real, imag} */,
  {32'h3f14fed8, 32'hc02e5561} /* (18, 12, 21) {real, imag} */,
  {32'h3fd6c01f, 32'h3fa22fb1} /* (18, 12, 20) {real, imag} */,
  {32'h3f20afac, 32'hbe691261} /* (18, 12, 19) {real, imag} */,
  {32'h3e75edd3, 32'hc00222fc} /* (18, 12, 18) {real, imag} */,
  {32'hbed2113c, 32'h3df1f671} /* (18, 12, 17) {real, imag} */,
  {32'hbd524f4d, 32'h3f8092ec} /* (18, 12, 16) {real, imag} */,
  {32'h4048c396, 32'h3f2cf768} /* (18, 12, 15) {real, imag} */,
  {32'hbfd9de1e, 32'h3f61a66e} /* (18, 12, 14) {real, imag} */,
  {32'h3f33dbea, 32'h3edfd44d} /* (18, 12, 13) {real, imag} */,
  {32'h3fcd3eb5, 32'h3fac9755} /* (18, 12, 12) {real, imag} */,
  {32'hc0bf2a67, 32'h3f724dcc} /* (18, 12, 11) {real, imag} */,
  {32'h3f79de28, 32'hbfd5495f} /* (18, 12, 10) {real, imag} */,
  {32'hbf9e5f45, 32'h3e4d765b} /* (18, 12, 9) {real, imag} */,
  {32'hbfb2d4a4, 32'hbfa1886d} /* (18, 12, 8) {real, imag} */,
  {32'hc000dc34, 32'hbef7bc6b} /* (18, 12, 7) {real, imag} */,
  {32'hbf7b8989, 32'hbf0087dd} /* (18, 12, 6) {real, imag} */,
  {32'hc070ffa2, 32'hc00b03d0} /* (18, 12, 5) {real, imag} */,
  {32'h3ee56289, 32'h3f901cc3} /* (18, 12, 4) {real, imag} */,
  {32'hbfd8eaec, 32'h3f971fe7} /* (18, 12, 3) {real, imag} */,
  {32'h40104f75, 32'h3f85b21b} /* (18, 12, 2) {real, imag} */,
  {32'hbf72e530, 32'h3f1a0a2f} /* (18, 12, 1) {real, imag} */,
  {32'h3fb947a7, 32'hbdf45269} /* (18, 12, 0) {real, imag} */,
  {32'h3fdd552f, 32'h3f4669d4} /* (18, 11, 31) {real, imag} */,
  {32'h3ea7c99e, 32'h400d4c46} /* (18, 11, 30) {real, imag} */,
  {32'hbfa14cce, 32'hbe8fd4ad} /* (18, 11, 29) {real, imag} */,
  {32'h3b9cd32e, 32'hbfe17ae7} /* (18, 11, 28) {real, imag} */,
  {32'hbffb0c69, 32'h3ea967ef} /* (18, 11, 27) {real, imag} */,
  {32'h3e407d30, 32'h3fbb4752} /* (18, 11, 26) {real, imag} */,
  {32'hbec3225d, 32'hbf54aecd} /* (18, 11, 25) {real, imag} */,
  {32'hbceffc39, 32'h4007aebb} /* (18, 11, 24) {real, imag} */,
  {32'h3e0aa6b4, 32'h3e297a35} /* (18, 11, 23) {real, imag} */,
  {32'h40789ab1, 32'h3f95e2ae} /* (18, 11, 22) {real, imag} */,
  {32'hbfd29562, 32'hbe694d6b} /* (18, 11, 21) {real, imag} */,
  {32'h4003f188, 32'hc00edd88} /* (18, 11, 20) {real, imag} */,
  {32'hc00033ed, 32'h408b6964} /* (18, 11, 19) {real, imag} */,
  {32'h4038e1ad, 32'h3fc6089a} /* (18, 11, 18) {real, imag} */,
  {32'hc022a286, 32'hbf2ed7d0} /* (18, 11, 17) {real, imag} */,
  {32'h3e11e4ec, 32'h3fd7c304} /* (18, 11, 16) {real, imag} */,
  {32'h40056fa7, 32'h3f667795} /* (18, 11, 15) {real, imag} */,
  {32'hbfe91475, 32'hc0514a68} /* (18, 11, 14) {real, imag} */,
  {32'h3f5564ca, 32'h401a3ab0} /* (18, 11, 13) {real, imag} */,
  {32'hbf01056d, 32'hbd323af9} /* (18, 11, 12) {real, imag} */,
  {32'h401d05e5, 32'h3f411d73} /* (18, 11, 11) {real, imag} */,
  {32'hc03c613a, 32'hc03bc71f} /* (18, 11, 10) {real, imag} */,
  {32'hbf2027f5, 32'hbfcd198f} /* (18, 11, 9) {real, imag} */,
  {32'h406582cc, 32'h3f066a8d} /* (18, 11, 8) {real, imag} */,
  {32'h3efb5458, 32'h3fdd6ad6} /* (18, 11, 7) {real, imag} */,
  {32'h3f7edcae, 32'hbe51b83f} /* (18, 11, 6) {real, imag} */,
  {32'h4058099e, 32'h4014aad3} /* (18, 11, 5) {real, imag} */,
  {32'h400a6086, 32'hc02e1de9} /* (18, 11, 4) {real, imag} */,
  {32'h4038de62, 32'h40162163} /* (18, 11, 3) {real, imag} */,
  {32'hbf67382d, 32'h3e55bf44} /* (18, 11, 2) {real, imag} */,
  {32'h400ed8a8, 32'hc00e393e} /* (18, 11, 1) {real, imag} */,
  {32'hbf0464db, 32'h3fb06139} /* (18, 11, 0) {real, imag} */,
  {32'h4024e3e8, 32'hbf6b6b79} /* (18, 10, 31) {real, imag} */,
  {32'h400fc1a6, 32'h3fc90fe6} /* (18, 10, 30) {real, imag} */,
  {32'hbf00cf44, 32'hbe53d251} /* (18, 10, 29) {real, imag} */,
  {32'hc06cd0d3, 32'hbf1a0655} /* (18, 10, 28) {real, imag} */,
  {32'hc024e275, 32'hbe9cc57a} /* (18, 10, 27) {real, imag} */,
  {32'h3e1e1f1a, 32'h3f8c7cd9} /* (18, 10, 26) {real, imag} */,
  {32'h3fbbf9ec, 32'h3fabc9a1} /* (18, 10, 25) {real, imag} */,
  {32'hc012b02e, 32'hbde4ec57} /* (18, 10, 24) {real, imag} */,
  {32'h3fad402d, 32'h3e8a03cc} /* (18, 10, 23) {real, imag} */,
  {32'hc02367d5, 32'hbfaacd54} /* (18, 10, 22) {real, imag} */,
  {32'h3ffa1a8d, 32'h3fa80f6b} /* (18, 10, 21) {real, imag} */,
  {32'h4058f1e2, 32'hbebc1501} /* (18, 10, 20) {real, imag} */,
  {32'h3e8eedaa, 32'h3f4806ef} /* (18, 10, 19) {real, imag} */,
  {32'h3fb3ac65, 32'h3f46a95e} /* (18, 10, 18) {real, imag} */,
  {32'h3f6edf34, 32'h3faab0d6} /* (18, 10, 17) {real, imag} */,
  {32'h3fea7ea9, 32'hbe37e70c} /* (18, 10, 16) {real, imag} */,
  {32'hbda68e2c, 32'hbf897884} /* (18, 10, 15) {real, imag} */,
  {32'h3db75319, 32'h3f53073d} /* (18, 10, 14) {real, imag} */,
  {32'h404271b4, 32'h3c58cc69} /* (18, 10, 13) {real, imag} */,
  {32'h3f9af22f, 32'hbfb9df1a} /* (18, 10, 12) {real, imag} */,
  {32'h3f9cc8cf, 32'hc0a08d91} /* (18, 10, 11) {real, imag} */,
  {32'h3f99d184, 32'hbf746caa} /* (18, 10, 10) {real, imag} */,
  {32'h3f496009, 32'hbf2120b3} /* (18, 10, 9) {real, imag} */,
  {32'h3f37a133, 32'hbee53a8e} /* (18, 10, 8) {real, imag} */,
  {32'hbff7c681, 32'hbfa5dded} /* (18, 10, 7) {real, imag} */,
  {32'h3f9504e8, 32'hc0133d10} /* (18, 10, 6) {real, imag} */,
  {32'h3ff7aefd, 32'hbed7d140} /* (18, 10, 5) {real, imag} */,
  {32'hbfa3ebdb, 32'hbfaaf527} /* (18, 10, 4) {real, imag} */,
  {32'hbdb80f39, 32'h40099f5a} /* (18, 10, 3) {real, imag} */,
  {32'hbe9b6216, 32'h3e9d8aa6} /* (18, 10, 2) {real, imag} */,
  {32'hbe9e16b1, 32'h3e8ce1f2} /* (18, 10, 1) {real, imag} */,
  {32'h3fbfd123, 32'hbfafaa60} /* (18, 10, 0) {real, imag} */,
  {32'h3f7ece34, 32'hbf5fdade} /* (18, 9, 31) {real, imag} */,
  {32'hbeb684a2, 32'hc0462097} /* (18, 9, 30) {real, imag} */,
  {32'hc017fd09, 32'hbf8fcc75} /* (18, 9, 29) {real, imag} */,
  {32'h400c39a6, 32'hbea0a593} /* (18, 9, 28) {real, imag} */,
  {32'h400efd5e, 32'hbf4a68d3} /* (18, 9, 27) {real, imag} */,
  {32'h3f81aee7, 32'hbf006b68} /* (18, 9, 26) {real, imag} */,
  {32'h4010e302, 32'h3f83db31} /* (18, 9, 25) {real, imag} */,
  {32'h3e2bb97a, 32'hc0406c70} /* (18, 9, 24) {real, imag} */,
  {32'hbf07e7f4, 32'hbf9355d9} /* (18, 9, 23) {real, imag} */,
  {32'hbf622f3e, 32'h3f4148f9} /* (18, 9, 22) {real, imag} */,
  {32'hbfadb98c, 32'hbe273981} /* (18, 9, 21) {real, imag} */,
  {32'h3e402d55, 32'h3f8ec9bd} /* (18, 9, 20) {real, imag} */,
  {32'h3faec888, 32'h3f23bdba} /* (18, 9, 19) {real, imag} */,
  {32'h40027d02, 32'h3f1ded62} /* (18, 9, 18) {real, imag} */,
  {32'h3fc37955, 32'h3fb6017d} /* (18, 9, 17) {real, imag} */,
  {32'hbef4d866, 32'h40062631} /* (18, 9, 16) {real, imag} */,
  {32'h3f41d606, 32'hbe9261e0} /* (18, 9, 15) {real, imag} */,
  {32'hbee1d024, 32'hbeaa2cb0} /* (18, 9, 14) {real, imag} */,
  {32'h3c3cefc3, 32'h3eb6e0a6} /* (18, 9, 13) {real, imag} */,
  {32'hbf64e0f3, 32'h3f41bff8} /* (18, 9, 12) {real, imag} */,
  {32'hbf6a85dd, 32'h3fc11ef2} /* (18, 9, 11) {real, imag} */,
  {32'h3f968033, 32'h4073aeb7} /* (18, 9, 10) {real, imag} */,
  {32'hbf4927c7, 32'h3fabd8fd} /* (18, 9, 9) {real, imag} */,
  {32'h3f934fff, 32'hbf58e950} /* (18, 9, 8) {real, imag} */,
  {32'h3e485989, 32'hbf983d7a} /* (18, 9, 7) {real, imag} */,
  {32'h401c5e5f, 32'hbf8223b5} /* (18, 9, 6) {real, imag} */,
  {32'hc0085920, 32'h3d7f91af} /* (18, 9, 5) {real, imag} */,
  {32'hc05b12fb, 32'h4001a8c8} /* (18, 9, 4) {real, imag} */,
  {32'h3fc4da23, 32'hbf19e898} /* (18, 9, 3) {real, imag} */,
  {32'hc00095f2, 32'h3f5faf7f} /* (18, 9, 2) {real, imag} */,
  {32'hbf859edc, 32'h3e334be4} /* (18, 9, 1) {real, imag} */,
  {32'hbf565ad7, 32'hbfdc73b9} /* (18, 9, 0) {real, imag} */,
  {32'h3ec21586, 32'h3fd84a84} /* (18, 8, 31) {real, imag} */,
  {32'hbf95d973, 32'h3f7bb9e0} /* (18, 8, 30) {real, imag} */,
  {32'h3f27935f, 32'h3e2bdd32} /* (18, 8, 29) {real, imag} */,
  {32'h3f446d82, 32'hc01bd700} /* (18, 8, 28) {real, imag} */,
  {32'hbfe8ce88, 32'hbf0ee0c9} /* (18, 8, 27) {real, imag} */,
  {32'hbf4584a8, 32'h3f57b428} /* (18, 8, 26) {real, imag} */,
  {32'hbf6d3311, 32'hbf1e1c4e} /* (18, 8, 25) {real, imag} */,
  {32'hc03b380e, 32'hbf9442dd} /* (18, 8, 24) {real, imag} */,
  {32'h3f23e217, 32'hbfc1c5c8} /* (18, 8, 23) {real, imag} */,
  {32'h3f577dc6, 32'hc0011dcc} /* (18, 8, 22) {real, imag} */,
  {32'h3f20a9a6, 32'hbfa306b3} /* (18, 8, 21) {real, imag} */,
  {32'hbdd2ebe4, 32'hc07b4002} /* (18, 8, 20) {real, imag} */,
  {32'h4094d11c, 32'h4006a223} /* (18, 8, 19) {real, imag} */,
  {32'hbf68108e, 32'h3ff41a7d} /* (18, 8, 18) {real, imag} */,
  {32'hbf62ee12, 32'hbfc440c5} /* (18, 8, 17) {real, imag} */,
  {32'h3faa471e, 32'hbd8f1b97} /* (18, 8, 16) {real, imag} */,
  {32'hbf2e02e2, 32'h3f7ae7af} /* (18, 8, 15) {real, imag} */,
  {32'h3e9ab0ae, 32'hbf72b8f4} /* (18, 8, 14) {real, imag} */,
  {32'hc029fd26, 32'hc00a84dd} /* (18, 8, 13) {real, imag} */,
  {32'hbfb0c84e, 32'hbfc1e514} /* (18, 8, 12) {real, imag} */,
  {32'h3e841ee2, 32'hbf9c6f71} /* (18, 8, 11) {real, imag} */,
  {32'hc0074c48, 32'hbf415fba} /* (18, 8, 10) {real, imag} */,
  {32'h3f69639c, 32'hbf9613db} /* (18, 8, 9) {real, imag} */,
  {32'h3ead3312, 32'h407a2093} /* (18, 8, 8) {real, imag} */,
  {32'h3fba3131, 32'h3fbb1e0e} /* (18, 8, 7) {real, imag} */,
  {32'h3e74f7a2, 32'h403cb7de} /* (18, 8, 6) {real, imag} */,
  {32'h3ff83570, 32'h3ff24b62} /* (18, 8, 5) {real, imag} */,
  {32'hbf901748, 32'h3fa30fbf} /* (18, 8, 4) {real, imag} */,
  {32'hc002bf6a, 32'hbed4932f} /* (18, 8, 3) {real, imag} */,
  {32'hc036bd04, 32'hbf2ba0bd} /* (18, 8, 2) {real, imag} */,
  {32'h3fbeadf6, 32'h3fddcc89} /* (18, 8, 1) {real, imag} */,
  {32'h3f1e5721, 32'h3dc88d38} /* (18, 8, 0) {real, imag} */,
  {32'h3fab096e, 32'hbf3fd247} /* (18, 7, 31) {real, imag} */,
  {32'h40409320, 32'hc0312ef3} /* (18, 7, 30) {real, imag} */,
  {32'hc002b561, 32'hbf5bbbed} /* (18, 7, 29) {real, imag} */,
  {32'h3e41be8b, 32'h3f93cef1} /* (18, 7, 28) {real, imag} */,
  {32'hbf4e208f, 32'hbff06c34} /* (18, 7, 27) {real, imag} */,
  {32'hbec92e25, 32'h3fcf55ca} /* (18, 7, 26) {real, imag} */,
  {32'hc0386d1a, 32'h3f6724cd} /* (18, 7, 25) {real, imag} */,
  {32'hbe7b02df, 32'hbeda3d97} /* (18, 7, 24) {real, imag} */,
  {32'h3e30cf5d, 32'hbfd0bd49} /* (18, 7, 23) {real, imag} */,
  {32'h3f13cbc0, 32'hbe998aa2} /* (18, 7, 22) {real, imag} */,
  {32'h402ba77e, 32'h3e89c25f} /* (18, 7, 21) {real, imag} */,
  {32'h3ebd1121, 32'hbc90dced} /* (18, 7, 20) {real, imag} */,
  {32'h4033bca6, 32'hbf8bf77c} /* (18, 7, 19) {real, imag} */,
  {32'hbe6a8938, 32'hbee5dfc1} /* (18, 7, 18) {real, imag} */,
  {32'hc0030a72, 32'hbf0c2010} /* (18, 7, 17) {real, imag} */,
  {32'h3eef612a, 32'hbf2899c3} /* (18, 7, 16) {real, imag} */,
  {32'hbfbac42a, 32'h3fd6539b} /* (18, 7, 15) {real, imag} */,
  {32'hbf11a87b, 32'hbfdd4e2d} /* (18, 7, 14) {real, imag} */,
  {32'h3d11e014, 32'h3f8928a4} /* (18, 7, 13) {real, imag} */,
  {32'hbf4604d1, 32'h3db6b968} /* (18, 7, 12) {real, imag} */,
  {32'h3d07c622, 32'hbf095a84} /* (18, 7, 11) {real, imag} */,
  {32'h40231683, 32'h3ed1c766} /* (18, 7, 10) {real, imag} */,
  {32'hbeeceaac, 32'hbfe3fa7d} /* (18, 7, 9) {real, imag} */,
  {32'hbf34ea51, 32'h3ebf6193} /* (18, 7, 8) {real, imag} */,
  {32'h3f159d4d, 32'hbf66c2d9} /* (18, 7, 7) {real, imag} */,
  {32'hbfc185c1, 32'hbe26deab} /* (18, 7, 6) {real, imag} */,
  {32'h40039643, 32'h4007c89b} /* (18, 7, 5) {real, imag} */,
  {32'h3eacaa94, 32'h3ea63309} /* (18, 7, 4) {real, imag} */,
  {32'h3f8af3c5, 32'hbfc2d666} /* (18, 7, 3) {real, imag} */,
  {32'h3f8883a8, 32'hbff6e8d6} /* (18, 7, 2) {real, imag} */,
  {32'hc038a073, 32'hbfcaed3f} /* (18, 7, 1) {real, imag} */,
  {32'hbf3d7b39, 32'hbf804248} /* (18, 7, 0) {real, imag} */,
  {32'h3ea3bba3, 32'hbfa76f4e} /* (18, 6, 31) {real, imag} */,
  {32'hbfe1e314, 32'hbdaca3fc} /* (18, 6, 30) {real, imag} */,
  {32'h3eef35cc, 32'hc00a4338} /* (18, 6, 29) {real, imag} */,
  {32'hbf9579f1, 32'h3cc46f32} /* (18, 6, 28) {real, imag} */,
  {32'h3fbc2390, 32'hbd89fc94} /* (18, 6, 27) {real, imag} */,
  {32'hbf07ab44, 32'h3e7cbb6b} /* (18, 6, 26) {real, imag} */,
  {32'h3f2a98bf, 32'hbe427b53} /* (18, 6, 25) {real, imag} */,
  {32'h3f917095, 32'h3f33f61a} /* (18, 6, 24) {real, imag} */,
  {32'hbeb4e332, 32'h3f9890ef} /* (18, 6, 23) {real, imag} */,
  {32'h3fdca29c, 32'hbf6ca5f4} /* (18, 6, 22) {real, imag} */,
  {32'hbf3aff73, 32'h3f91dc31} /* (18, 6, 21) {real, imag} */,
  {32'h3f2425dc, 32'h3f80dfae} /* (18, 6, 20) {real, imag} */,
  {32'hbf9dc677, 32'h3df1b4dd} /* (18, 6, 19) {real, imag} */,
  {32'hbf84fc47, 32'hbf8ae316} /* (18, 6, 18) {real, imag} */,
  {32'h3f74e743, 32'h3fb60aab} /* (18, 6, 17) {real, imag} */,
  {32'h4016a967, 32'hbf971649} /* (18, 6, 16) {real, imag} */,
  {32'hbe619acb, 32'h3f59138f} /* (18, 6, 15) {real, imag} */,
  {32'hbfe71b60, 32'h4049eb27} /* (18, 6, 14) {real, imag} */,
  {32'hbe1cf528, 32'hbf0a1d55} /* (18, 6, 13) {real, imag} */,
  {32'hbf70af3c, 32'hbf5d32b2} /* (18, 6, 12) {real, imag} */,
  {32'h3fcb8713, 32'h3f1f912b} /* (18, 6, 11) {real, imag} */,
  {32'h40265984, 32'h3fd3c420} /* (18, 6, 10) {real, imag} */,
  {32'hbef2d64b, 32'hbf98548b} /* (18, 6, 9) {real, imag} */,
  {32'h3f8430ca, 32'hbef4e2c4} /* (18, 6, 8) {real, imag} */,
  {32'h3f847d62, 32'h4000d662} /* (18, 6, 7) {real, imag} */,
  {32'hc03104da, 32'h3e7aed1d} /* (18, 6, 6) {real, imag} */,
  {32'hbe324767, 32'hbea71695} /* (18, 6, 5) {real, imag} */,
  {32'h3f386fd8, 32'hbf01b69e} /* (18, 6, 4) {real, imag} */,
  {32'hbf877797, 32'h3ff827db} /* (18, 6, 3) {real, imag} */,
  {32'h3f96b4d3, 32'hbfb0256e} /* (18, 6, 2) {real, imag} */,
  {32'h3f62760e, 32'hbd472edf} /* (18, 6, 1) {real, imag} */,
  {32'hbffad8dd, 32'hbfc50e77} /* (18, 6, 0) {real, imag} */,
  {32'h4025f766, 32'h401d855f} /* (18, 5, 31) {real, imag} */,
  {32'hbfae68d9, 32'hbe92d6fa} /* (18, 5, 30) {real, imag} */,
  {32'h3f24f4a0, 32'hbe1b9b32} /* (18, 5, 29) {real, imag} */,
  {32'h40336357, 32'h3f46bb9c} /* (18, 5, 28) {real, imag} */,
  {32'hbfa2ce58, 32'hc01fec49} /* (18, 5, 27) {real, imag} */,
  {32'hbeb28631, 32'hbfc8d1f0} /* (18, 5, 26) {real, imag} */,
  {32'h3fac5b9e, 32'h3e5bbf08} /* (18, 5, 25) {real, imag} */,
  {32'h3fac5c80, 32'h40050aff} /* (18, 5, 24) {real, imag} */,
  {32'hbe1bafa2, 32'hbf59826b} /* (18, 5, 23) {real, imag} */,
  {32'h400ec146, 32'h3f1bd3b0} /* (18, 5, 22) {real, imag} */,
  {32'h3ebf410c, 32'h3f8b2be5} /* (18, 5, 21) {real, imag} */,
  {32'hc0260357, 32'h3ffe3de8} /* (18, 5, 20) {real, imag} */,
  {32'hc0192919, 32'h3fa59d4d} /* (18, 5, 19) {real, imag} */,
  {32'hbf153ccb, 32'hbf1145ae} /* (18, 5, 18) {real, imag} */,
  {32'h401d2be8, 32'h403f93ae} /* (18, 5, 17) {real, imag} */,
  {32'h3f6c4b7b, 32'h3e8ee9cd} /* (18, 5, 16) {real, imag} */,
  {32'h3f23bb36, 32'h3ef7ef0d} /* (18, 5, 15) {real, imag} */,
  {32'h3d348ff9, 32'hbf9d91ef} /* (18, 5, 14) {real, imag} */,
  {32'h3f2ba5d4, 32'h3f1a306a} /* (18, 5, 13) {real, imag} */,
  {32'hc023a877, 32'h40150e4c} /* (18, 5, 12) {real, imag} */,
  {32'hc02175fe, 32'hc0416785} /* (18, 5, 11) {real, imag} */,
  {32'hbf44b7ef, 32'h3e91cfe5} /* (18, 5, 10) {real, imag} */,
  {32'hc063cc93, 32'h3fc7dae1} /* (18, 5, 9) {real, imag} */,
  {32'hbcd5986e, 32'hbec82817} /* (18, 5, 8) {real, imag} */,
  {32'hbecd4ade, 32'h3fdba501} /* (18, 5, 7) {real, imag} */,
  {32'h3fbfe5cc, 32'h3f986996} /* (18, 5, 6) {real, imag} */,
  {32'hbf9597cc, 32'hbf5a12ea} /* (18, 5, 5) {real, imag} */,
  {32'h3e88fba6, 32'hbe7ec093} /* (18, 5, 4) {real, imag} */,
  {32'hbfa94193, 32'hbfea7b29} /* (18, 5, 3) {real, imag} */,
  {32'hbec92072, 32'hc0866939} /* (18, 5, 2) {real, imag} */,
  {32'h3edce174, 32'hbd99ec12} /* (18, 5, 1) {real, imag} */,
  {32'h3fd57dde, 32'hbff0a8dd} /* (18, 5, 0) {real, imag} */,
  {32'hc0013e50, 32'hc01328f3} /* (18, 4, 31) {real, imag} */,
  {32'hbbfc783c, 32'h3f3dde7b} /* (18, 4, 30) {real, imag} */,
  {32'h40214a95, 32'h3fae1233} /* (18, 4, 29) {real, imag} */,
  {32'hc05bf039, 32'h402ea756} /* (18, 4, 28) {real, imag} */,
  {32'h405d63dd, 32'h3f8f3f25} /* (18, 4, 27) {real, imag} */,
  {32'hbe66b9e0, 32'hbe64b950} /* (18, 4, 26) {real, imag} */,
  {32'hbf96d50a, 32'h3f78031d} /* (18, 4, 25) {real, imag} */,
  {32'h400d5bcb, 32'h3e3252b3} /* (18, 4, 24) {real, imag} */,
  {32'hc02aae93, 32'hbe0e95db} /* (18, 4, 23) {real, imag} */,
  {32'hbd68fa29, 32'hbefec91e} /* (18, 4, 22) {real, imag} */,
  {32'hbf865334, 32'hc0267db5} /* (18, 4, 21) {real, imag} */,
  {32'hbf9b8738, 32'h3ff83c86} /* (18, 4, 20) {real, imag} */,
  {32'hbf13b6fc, 32'hbdf3c73e} /* (18, 4, 19) {real, imag} */,
  {32'hc02ee98d, 32'h3fba2b7d} /* (18, 4, 18) {real, imag} */,
  {32'h3e16c384, 32'hbf4823d2} /* (18, 4, 17) {real, imag} */,
  {32'hbf2af7e6, 32'hbe8bf860} /* (18, 4, 16) {real, imag} */,
  {32'h3fe6f0d9, 32'hbf0b4243} /* (18, 4, 15) {real, imag} */,
  {32'hbf89dbe1, 32'hbe7c4284} /* (18, 4, 14) {real, imag} */,
  {32'hc023ada2, 32'hbf4380bc} /* (18, 4, 13) {real, imag} */,
  {32'h3f74d6ff, 32'h3e0fe423} /* (18, 4, 12) {real, imag} */,
  {32'hbff83b33, 32'hbe449646} /* (18, 4, 11) {real, imag} */,
  {32'h3de189af, 32'h4031e200} /* (18, 4, 10) {real, imag} */,
  {32'hbed2c60e, 32'hbf125e67} /* (18, 4, 9) {real, imag} */,
  {32'h3fd3b5b2, 32'h409ea28c} /* (18, 4, 8) {real, imag} */,
  {32'hc0588763, 32'hbfd78adf} /* (18, 4, 7) {real, imag} */,
  {32'h3f50fe21, 32'h3ffa7f29} /* (18, 4, 6) {real, imag} */,
  {32'hbe1a1b53, 32'h3fdf00e0} /* (18, 4, 5) {real, imag} */,
  {32'h3feeb736, 32'hbe0f7d9b} /* (18, 4, 4) {real, imag} */,
  {32'h4017cfb0, 32'hbf11a96b} /* (18, 4, 3) {real, imag} */,
  {32'h4036aba6, 32'hbfbe0d1f} /* (18, 4, 2) {real, imag} */,
  {32'hbfcb3a94, 32'hc07dc960} /* (18, 4, 1) {real, imag} */,
  {32'hbf932926, 32'h3f2c38bc} /* (18, 4, 0) {real, imag} */,
  {32'hbeba672a, 32'hbf945ce4} /* (18, 3, 31) {real, imag} */,
  {32'h3f8f2d41, 32'h3e1041c2} /* (18, 3, 30) {real, imag} */,
  {32'hc01a0a64, 32'h3fffe960} /* (18, 3, 29) {real, imag} */,
  {32'hbfc55812, 32'hbd8642c5} /* (18, 3, 28) {real, imag} */,
  {32'h3ebb7cee, 32'hbf3dd477} /* (18, 3, 27) {real, imag} */,
  {32'h4052fea4, 32'hbdfe4a17} /* (18, 3, 26) {real, imag} */,
  {32'hbf68e8cd, 32'hc03ded2c} /* (18, 3, 25) {real, imag} */,
  {32'h3eb5f92f, 32'h3f9759fe} /* (18, 3, 24) {real, imag} */,
  {32'hbf12abe1, 32'hbf2f6847} /* (18, 3, 23) {real, imag} */,
  {32'hbfef2446, 32'hbffe8695} /* (18, 3, 22) {real, imag} */,
  {32'h3ef1b9ff, 32'hbdbae815} /* (18, 3, 21) {real, imag} */,
  {32'hbec7bc38, 32'h3f621bff} /* (18, 3, 20) {real, imag} */,
  {32'h3e9ab749, 32'h3f64ecd2} /* (18, 3, 19) {real, imag} */,
  {32'h40315954, 32'h3d1d1a0a} /* (18, 3, 18) {real, imag} */,
  {32'hbf9692d2, 32'hbfc21083} /* (18, 3, 17) {real, imag} */,
  {32'h3f0ad788, 32'hbf73a11c} /* (18, 3, 16) {real, imag} */,
  {32'h4028743d, 32'h4019fc20} /* (18, 3, 15) {real, imag} */,
  {32'h3ee47fda, 32'h3f278543} /* (18, 3, 14) {real, imag} */,
  {32'h400496a0, 32'hbf16156f} /* (18, 3, 13) {real, imag} */,
  {32'hc018fbd3, 32'hbf9c1815} /* (18, 3, 12) {real, imag} */,
  {32'hbe4ddbd1, 32'hbfc7373e} /* (18, 3, 11) {real, imag} */,
  {32'h3f9f7818, 32'hbe11af33} /* (18, 3, 10) {real, imag} */,
  {32'hbf8ec073, 32'h3feefb32} /* (18, 3, 9) {real, imag} */,
  {32'hc030c8a1, 32'h3f2921ba} /* (18, 3, 8) {real, imag} */,
  {32'h404cce03, 32'hbfe47ebc} /* (18, 3, 7) {real, imag} */,
  {32'hbe35ec4e, 32'h3e561716} /* (18, 3, 6) {real, imag} */,
  {32'hbf9a9446, 32'hbfe0691d} /* (18, 3, 5) {real, imag} */,
  {32'h3c81a768, 32'h3f622609} /* (18, 3, 4) {real, imag} */,
  {32'h3f067d33, 32'h4022204b} /* (18, 3, 3) {real, imag} */,
  {32'h3f83f546, 32'h3f82ec5b} /* (18, 3, 2) {real, imag} */,
  {32'hc01dfb7b, 32'h3d9e1800} /* (18, 3, 1) {real, imag} */,
  {32'hbfb24d58, 32'hbfbd1608} /* (18, 3, 0) {real, imag} */,
  {32'h40ab856b, 32'h4006cad8} /* (18, 2, 31) {real, imag} */,
  {32'hc0684acd, 32'hbe9493c7} /* (18, 2, 30) {real, imag} */,
  {32'h40023a9d, 32'h3f88360c} /* (18, 2, 29) {real, imag} */,
  {32'h400a5bc7, 32'hbf880333} /* (18, 2, 28) {real, imag} */,
  {32'hbf9cfabb, 32'hbf017e05} /* (18, 2, 27) {real, imag} */,
  {32'h3f3522b6, 32'hbed24c77} /* (18, 2, 26) {real, imag} */,
  {32'hbf87826f, 32'hbf5c27e8} /* (18, 2, 25) {real, imag} */,
  {32'hbfc79a92, 32'hbe10eb83} /* (18, 2, 24) {real, imag} */,
  {32'h40188c17, 32'h3f081b8f} /* (18, 2, 23) {real, imag} */,
  {32'h3ff0c7fe, 32'h400b3000} /* (18, 2, 22) {real, imag} */,
  {32'hbfa89251, 32'hbf1832e6} /* (18, 2, 21) {real, imag} */,
  {32'h40088dba, 32'h3f51b19e} /* (18, 2, 20) {real, imag} */,
  {32'hbdf12b1b, 32'hbf84ee64} /* (18, 2, 19) {real, imag} */,
  {32'hbd463cc2, 32'hc007b646} /* (18, 2, 18) {real, imag} */,
  {32'hbfeb53cd, 32'hbf4bd02e} /* (18, 2, 17) {real, imag} */,
  {32'hbfb2644a, 32'h3f1d9c09} /* (18, 2, 16) {real, imag} */,
  {32'hbe910184, 32'h3eb63d6b} /* (18, 2, 15) {real, imag} */,
  {32'h3f4db245, 32'h3e64d18b} /* (18, 2, 14) {real, imag} */,
  {32'hc0482179, 32'hbf0d9449} /* (18, 2, 13) {real, imag} */,
  {32'hbeafa363, 32'hbe9e907c} /* (18, 2, 12) {real, imag} */,
  {32'hbe990b5f, 32'hbf7a1821} /* (18, 2, 11) {real, imag} */,
  {32'h4026d91a, 32'h3ec56334} /* (18, 2, 10) {real, imag} */,
  {32'h3d224423, 32'h3f8a9b3a} /* (18, 2, 9) {real, imag} */,
  {32'hc0024e98, 32'h3f331ab1} /* (18, 2, 8) {real, imag} */,
  {32'h3f8ead60, 32'hbfa1f9e5} /* (18, 2, 7) {real, imag} */,
  {32'hbf8cb089, 32'h3e19b3f1} /* (18, 2, 6) {real, imag} */,
  {32'hbfdcf19b, 32'hbfd5e926} /* (18, 2, 5) {real, imag} */,
  {32'hbde84ad6, 32'hbfec1935} /* (18, 2, 4) {real, imag} */,
  {32'hbe5031b4, 32'hbf2ab9aa} /* (18, 2, 3) {real, imag} */,
  {32'hc060b778, 32'hbf2fdf06} /* (18, 2, 2) {real, imag} */,
  {32'h40b0771d, 32'h3ec8a1ff} /* (18, 2, 1) {real, imag} */,
  {32'h4020173e, 32'hbed7527e} /* (18, 2, 0) {real, imag} */,
  {32'hc07df3ac, 32'hbf5b45ef} /* (18, 1, 31) {real, imag} */,
  {32'h3fb36a21, 32'h3f6a462c} /* (18, 1, 30) {real, imag} */,
  {32'h3f476487, 32'hbb450ef7} /* (18, 1, 29) {real, imag} */,
  {32'hbcce9749, 32'hbf6324c3} /* (18, 1, 28) {real, imag} */,
  {32'h3fac482e, 32'hbf76e5d0} /* (18, 1, 27) {real, imag} */,
  {32'hbefa11f4, 32'hc022fd0e} /* (18, 1, 26) {real, imag} */,
  {32'h3fd9f702, 32'h3f373ca5} /* (18, 1, 25) {real, imag} */,
  {32'h3e30dc6b, 32'h4007adc3} /* (18, 1, 24) {real, imag} */,
  {32'h3f436756, 32'h3f8c0629} /* (18, 1, 23) {real, imag} */,
  {32'hc03d1811, 32'h3f8a35fd} /* (18, 1, 22) {real, imag} */,
  {32'h404b576b, 32'hbd15e57d} /* (18, 1, 21) {real, imag} */,
  {32'hbf201953, 32'h3c78240c} /* (18, 1, 20) {real, imag} */,
  {32'hbff006a7, 32'h3e7881b0} /* (18, 1, 19) {real, imag} */,
  {32'h3ed0ca3e, 32'h3f476807} /* (18, 1, 18) {real, imag} */,
  {32'hbf8f8dcd, 32'hbf40516f} /* (18, 1, 17) {real, imag} */,
  {32'h3ed6632f, 32'h3fe42260} /* (18, 1, 16) {real, imag} */,
  {32'hbfb3aeef, 32'h3ec25e89} /* (18, 1, 15) {real, imag} */,
  {32'h3fb8d597, 32'hbd0a3b4c} /* (18, 1, 14) {real, imag} */,
  {32'h3ef543c7, 32'hbf4a4e3f} /* (18, 1, 13) {real, imag} */,
  {32'h3f2e963d, 32'hbe88fbb5} /* (18, 1, 12) {real, imag} */,
  {32'h400de8a0, 32'h4023fe13} /* (18, 1, 11) {real, imag} */,
  {32'h4023710e, 32'hbf87ab50} /* (18, 1, 10) {real, imag} */,
  {32'h3f679673, 32'h3f9fe3ee} /* (18, 1, 9) {real, imag} */,
  {32'h3e0f1b7c, 32'h401b419d} /* (18, 1, 8) {real, imag} */,
  {32'hc04c61cc, 32'h3f69af87} /* (18, 1, 7) {real, imag} */,
  {32'hbf1d7c9e, 32'h3ffa526a} /* (18, 1, 6) {real, imag} */,
  {32'hbfcefb5c, 32'h3f2668ae} /* (18, 1, 5) {real, imag} */,
  {32'hbe66489a, 32'hbf6056a8} /* (18, 1, 4) {real, imag} */,
  {32'h3fd0fea4, 32'hbfa9e29c} /* (18, 1, 3) {real, imag} */,
  {32'h3f6c3eab, 32'h4055b25b} /* (18, 1, 2) {real, imag} */,
  {32'hc0b00dcb, 32'hbfa46337} /* (18, 1, 1) {real, imag} */,
  {32'hc03c4dbd, 32'h3e0fb841} /* (18, 1, 0) {real, imag} */,
  {32'hbfc2025c, 32'h405bc53f} /* (18, 0, 31) {real, imag} */,
  {32'h403a7e8a, 32'hbf541e48} /* (18, 0, 30) {real, imag} */,
  {32'hc013d3bb, 32'h3efd7ea7} /* (18, 0, 29) {real, imag} */,
  {32'hbf97ba16, 32'hbd3ebf79} /* (18, 0, 28) {real, imag} */,
  {32'h3d5f5beb, 32'hbe3d9de2} /* (18, 0, 27) {real, imag} */,
  {32'hbf8473bd, 32'h3f3366be} /* (18, 0, 26) {real, imag} */,
  {32'hbfec47c9, 32'h3db15c6b} /* (18, 0, 25) {real, imag} */,
  {32'hbfca1147, 32'hbe7184b8} /* (18, 0, 24) {real, imag} */,
  {32'h3f9e5b2a, 32'h40863a11} /* (18, 0, 23) {real, imag} */,
  {32'hbf7fec6a, 32'hbff87ce1} /* (18, 0, 22) {real, imag} */,
  {32'h3e98ef32, 32'hbfe0571e} /* (18, 0, 21) {real, imag} */,
  {32'h3f626239, 32'hbd306639} /* (18, 0, 20) {real, imag} */,
  {32'hbf93ec11, 32'hbf4ed9bb} /* (18, 0, 19) {real, imag} */,
  {32'h3f1982f7, 32'hbf2dbcbf} /* (18, 0, 18) {real, imag} */,
  {32'h3f69a5ca, 32'hc02e482e} /* (18, 0, 17) {real, imag} */,
  {32'hbfa6ba06, 32'h3f8bbece} /* (18, 0, 16) {real, imag} */,
  {32'h3ee40a0c, 32'hbdc55b19} /* (18, 0, 15) {real, imag} */,
  {32'hbf84f327, 32'h3ead51c1} /* (18, 0, 14) {real, imag} */,
  {32'h3d8271dd, 32'hbfa0f6a5} /* (18, 0, 13) {real, imag} */,
  {32'hbca740b3, 32'hbdfab48c} /* (18, 0, 12) {real, imag} */,
  {32'h3f77379d, 32'h3ee38d3e} /* (18, 0, 11) {real, imag} */,
  {32'h3e5294f0, 32'hbf3d4601} /* (18, 0, 10) {real, imag} */,
  {32'h40167802, 32'h3fd38a71} /* (18, 0, 9) {real, imag} */,
  {32'hbfed6d0e, 32'h3f784581} /* (18, 0, 8) {real, imag} */,
  {32'h3ffe8523, 32'hc047c1f0} /* (18, 0, 7) {real, imag} */,
  {32'hc0112a53, 32'hc03b0452} /* (18, 0, 6) {real, imag} */,
  {32'h3ff37a52, 32'h3d2e893b} /* (18, 0, 5) {real, imag} */,
  {32'h401bf50c, 32'h3ec09f4b} /* (18, 0, 4) {real, imag} */,
  {32'h3f52be18, 32'h3fe637ab} /* (18, 0, 3) {real, imag} */,
  {32'h3f14056c, 32'hbf81543c} /* (18, 0, 2) {real, imag} */,
  {32'hbf7935ec, 32'hbfd9163a} /* (18, 0, 1) {real, imag} */,
  {32'hbff4f8bc, 32'hbfd9fdda} /* (18, 0, 0) {real, imag} */,
  {32'h40511ec0, 32'hbf47af05} /* (17, 31, 31) {real, imag} */,
  {32'hbff8ee7d, 32'h3ff7be5a} /* (17, 31, 30) {real, imag} */,
  {32'hbf7b3fb3, 32'h3f0dc7c0} /* (17, 31, 29) {real, imag} */,
  {32'h3f5384b5, 32'hbf86d8b1} /* (17, 31, 28) {real, imag} */,
  {32'hbfe902bc, 32'hbf26e949} /* (17, 31, 27) {real, imag} */,
  {32'h3e3462e3, 32'hbf198541} /* (17, 31, 26) {real, imag} */,
  {32'h3f2efc71, 32'hbfaf30d4} /* (17, 31, 25) {real, imag} */,
  {32'hbf8992d8, 32'h3f2f6d9d} /* (17, 31, 24) {real, imag} */,
  {32'h3fe49559, 32'hbfd22377} /* (17, 31, 23) {real, imag} */,
  {32'h3f6a5460, 32'h3f81e409} /* (17, 31, 22) {real, imag} */,
  {32'h3f7c6cdb, 32'hbfcfefcc} /* (17, 31, 21) {real, imag} */,
  {32'h3f868d92, 32'h3fd7cc09} /* (17, 31, 20) {real, imag} */,
  {32'h3f779cff, 32'h3f10c976} /* (17, 31, 19) {real, imag} */,
  {32'h3e8491ac, 32'h3fd378a6} /* (17, 31, 18) {real, imag} */,
  {32'h3f113aa0, 32'h3eb8c647} /* (17, 31, 17) {real, imag} */,
  {32'hc0034712, 32'h4000e57c} /* (17, 31, 16) {real, imag} */,
  {32'h3e18dd58, 32'h3f39df0c} /* (17, 31, 15) {real, imag} */,
  {32'h3ec9f78d, 32'h3f0560de} /* (17, 31, 14) {real, imag} */,
  {32'hbf30d1db, 32'h3faa4b7b} /* (17, 31, 13) {real, imag} */,
  {32'h3fca1ac8, 32'hbfe84b99} /* (17, 31, 12) {real, imag} */,
  {32'h3e097fb3, 32'h3f25382a} /* (17, 31, 11) {real, imag} */,
  {32'h3e5e0f22, 32'hbf39c547} /* (17, 31, 10) {real, imag} */,
  {32'h403b888f, 32'hbf8d85c5} /* (17, 31, 9) {real, imag} */,
  {32'hbec8381a, 32'hbfcf6765} /* (17, 31, 8) {real, imag} */,
  {32'h3f40767d, 32'hbc1c503e} /* (17, 31, 7) {real, imag} */,
  {32'hbf9956ac, 32'hbe6e1e42} /* (17, 31, 6) {real, imag} */,
  {32'h3f08202b, 32'h3dd92afe} /* (17, 31, 5) {real, imag} */,
  {32'h3ef53360, 32'h3d1fe423} /* (17, 31, 4) {real, imag} */,
  {32'h3f77752d, 32'hbf1172f4} /* (17, 31, 3) {real, imag} */,
  {32'hbf707c4e, 32'hbf517b55} /* (17, 31, 2) {real, imag} */,
  {32'h3fe97c8d, 32'hbed97682} /* (17, 31, 1) {real, imag} */,
  {32'h3fb21377, 32'hbf8d27de} /* (17, 31, 0) {real, imag} */,
  {32'hbfe42a7c, 32'h3fbcff38} /* (17, 30, 31) {real, imag} */,
  {32'h3f8fbb0c, 32'h3f79cad9} /* (17, 30, 30) {real, imag} */,
  {32'hc01ef885, 32'hbf71852d} /* (17, 30, 29) {real, imag} */,
  {32'hbf3e190d, 32'hbc4eaa38} /* (17, 30, 28) {real, imag} */,
  {32'h3f80c55f, 32'h3f2d20a9} /* (17, 30, 27) {real, imag} */,
  {32'hbeba85a6, 32'h40397ae6} /* (17, 30, 26) {real, imag} */,
  {32'hbe55d896, 32'h3d0c9f60} /* (17, 30, 25) {real, imag} */,
  {32'hbf5a9ebe, 32'hbf0aad17} /* (17, 30, 24) {real, imag} */,
  {32'h3e215173, 32'hbf5a637e} /* (17, 30, 23) {real, imag} */,
  {32'hbe615a55, 32'hbf2fe733} /* (17, 30, 22) {real, imag} */,
  {32'h3e48b437, 32'h3fa59665} /* (17, 30, 21) {real, imag} */,
  {32'h3f8eba1a, 32'h3f869e44} /* (17, 30, 20) {real, imag} */,
  {32'h3d9298a6, 32'hbff2d967} /* (17, 30, 19) {real, imag} */,
  {32'hbfcea1e0, 32'h3f171ec0} /* (17, 30, 18) {real, imag} */,
  {32'hbf349d0f, 32'hbef7123b} /* (17, 30, 17) {real, imag} */,
  {32'h3eb5d6c9, 32'h3fda4df2} /* (17, 30, 16) {real, imag} */,
  {32'h3f5a34e4, 32'h3fda48aa} /* (17, 30, 15) {real, imag} */,
  {32'h3e626030, 32'h3f1cedc7} /* (17, 30, 14) {real, imag} */,
  {32'h3f0061ba, 32'hbff02c3c} /* (17, 30, 13) {real, imag} */,
  {32'hbf9305c7, 32'hbd354849} /* (17, 30, 12) {real, imag} */,
  {32'hbe4f5e38, 32'h405a7516} /* (17, 30, 11) {real, imag} */,
  {32'h3f235030, 32'h3f64e082} /* (17, 30, 10) {real, imag} */,
  {32'hbfd705bc, 32'h400ce850} /* (17, 30, 9) {real, imag} */,
  {32'hbf24e76a, 32'h3fbf9a3c} /* (17, 30, 8) {real, imag} */,
  {32'hbeb9e570, 32'hbfe70d50} /* (17, 30, 7) {real, imag} */,
  {32'h3ed994a0, 32'hc03e4912} /* (17, 30, 6) {real, imag} */,
  {32'h3ff92aa3, 32'hbf624b3a} /* (17, 30, 5) {real, imag} */,
  {32'hbe86e6d2, 32'h3f78e638} /* (17, 30, 4) {real, imag} */,
  {32'h3fa1569a, 32'hbf06214c} /* (17, 30, 3) {real, imag} */,
  {32'hbf9a774b, 32'h3e7edf65} /* (17, 30, 2) {real, imag} */,
  {32'hbf68f536, 32'h3eb5260c} /* (17, 30, 1) {real, imag} */,
  {32'h3e95acad, 32'hc027179d} /* (17, 30, 0) {real, imag} */,
  {32'h3fd08d6d, 32'hbeaf8868} /* (17, 29, 31) {real, imag} */,
  {32'hbe6140ac, 32'hbe1dbd86} /* (17, 29, 30) {real, imag} */,
  {32'h3e8c9b83, 32'hbf841797} /* (17, 29, 29) {real, imag} */,
  {32'h3edeb1b2, 32'hbd821171} /* (17, 29, 28) {real, imag} */,
  {32'h3fe5a4c1, 32'h3d85a8e1} /* (17, 29, 27) {real, imag} */,
  {32'h3dd41898, 32'hbf92978c} /* (17, 29, 26) {real, imag} */,
  {32'h3e6afeb3, 32'h3f665b6c} /* (17, 29, 25) {real, imag} */,
  {32'h3fb4937d, 32'h3f447277} /* (17, 29, 24) {real, imag} */,
  {32'hbf98d5a2, 32'hbd81d472} /* (17, 29, 23) {real, imag} */,
  {32'hbfec291b, 32'hc034d193} /* (17, 29, 22) {real, imag} */,
  {32'hbf767706, 32'hbf89afb8} /* (17, 29, 21) {real, imag} */,
  {32'h3fc5009b, 32'h3fda6e98} /* (17, 29, 20) {real, imag} */,
  {32'h3f5f5b7b, 32'hc0053bff} /* (17, 29, 19) {real, imag} */,
  {32'hbf900fd1, 32'hbf83d2d9} /* (17, 29, 18) {real, imag} */,
  {32'h3d80f20d, 32'h3f68b90d} /* (17, 29, 17) {real, imag} */,
  {32'hbee929ae, 32'hbe3e2a38} /* (17, 29, 16) {real, imag} */,
  {32'h4012507e, 32'hbfb7a88a} /* (17, 29, 15) {real, imag} */,
  {32'h3f266a5e, 32'h3f5a1032} /* (17, 29, 14) {real, imag} */,
  {32'hc025907d, 32'hbe3017eb} /* (17, 29, 13) {real, imag} */,
  {32'hbfe939ee, 32'hbf3e2ac2} /* (17, 29, 12) {real, imag} */,
  {32'hc05b4c07, 32'hbfb02398} /* (17, 29, 11) {real, imag} */,
  {32'h3fd5ed76, 32'h3e3798ef} /* (17, 29, 10) {real, imag} */,
  {32'h3eeef134, 32'hbd78a5e0} /* (17, 29, 9) {real, imag} */,
  {32'hbf6d8b2f, 32'h3f8b2f29} /* (17, 29, 8) {real, imag} */,
  {32'hbf7c71da, 32'hbfcb9736} /* (17, 29, 7) {real, imag} */,
  {32'h3f978c70, 32'hbf4dfd64} /* (17, 29, 6) {real, imag} */,
  {32'h40113cc6, 32'hbeabb745} /* (17, 29, 5) {real, imag} */,
  {32'hbe7918cb, 32'h3ddb17b2} /* (17, 29, 4) {real, imag} */,
  {32'h3cba7973, 32'h3fdc3379} /* (17, 29, 3) {real, imag} */,
  {32'hbff0bbb3, 32'h400c67fa} /* (17, 29, 2) {real, imag} */,
  {32'h3f634e23, 32'hbe2b3fc6} /* (17, 29, 1) {real, imag} */,
  {32'hbfc5f499, 32'hbf2f00af} /* (17, 29, 0) {real, imag} */,
  {32'h3dd68806, 32'h3ff57b23} /* (17, 28, 31) {real, imag} */,
  {32'hbbae8008, 32'h40004d6a} /* (17, 28, 30) {real, imag} */,
  {32'hbe2830e9, 32'h40103f78} /* (17, 28, 29) {real, imag} */,
  {32'h3faa7c7d, 32'hbff2d255} /* (17, 28, 28) {real, imag} */,
  {32'h3fb56660, 32'hbed5127d} /* (17, 28, 27) {real, imag} */,
  {32'hbd17fbb9, 32'h3fad4d90} /* (17, 28, 26) {real, imag} */,
  {32'hbf8ce9f0, 32'hbf4d43e1} /* (17, 28, 25) {real, imag} */,
  {32'hbf690a2f, 32'h3ece6f1b} /* (17, 28, 24) {real, imag} */,
  {32'hbf602572, 32'hbcbc3f54} /* (17, 28, 23) {real, imag} */,
  {32'hc0746db0, 32'h3f03cb88} /* (17, 28, 22) {real, imag} */,
  {32'h3fe2f5f0, 32'h400d7554} /* (17, 28, 21) {real, imag} */,
  {32'hbf5b3d42, 32'hc02bba8f} /* (17, 28, 20) {real, imag} */,
  {32'h3fe1b1a6, 32'h3e62cc86} /* (17, 28, 19) {real, imag} */,
  {32'h3f305ce7, 32'h3f09a88e} /* (17, 28, 18) {real, imag} */,
  {32'h3f1c6287, 32'hbf896326} /* (17, 28, 17) {real, imag} */,
  {32'h3ee9a3a6, 32'hbf5f3902} /* (17, 28, 16) {real, imag} */,
  {32'h3eeddef8, 32'h402f0c0e} /* (17, 28, 15) {real, imag} */,
  {32'h3f35ff73, 32'hbfc751db} /* (17, 28, 14) {real, imag} */,
  {32'hbf8bf166, 32'h3ecb6975} /* (17, 28, 13) {real, imag} */,
  {32'h3ec5d48d, 32'h40063596} /* (17, 28, 12) {real, imag} */,
  {32'h3d74941e, 32'hbff4f0fa} /* (17, 28, 11) {real, imag} */,
  {32'h3fa4c152, 32'h3dc1a8fb} /* (17, 28, 10) {real, imag} */,
  {32'h3ecbb8d8, 32'h3e666deb} /* (17, 28, 9) {real, imag} */,
  {32'hbd5064eb, 32'h3f7b2505} /* (17, 28, 8) {real, imag} */,
  {32'h4053fec8, 32'hbfbff6aa} /* (17, 28, 7) {real, imag} */,
  {32'hbfad67b7, 32'h3fd3c0ec} /* (17, 28, 6) {real, imag} */,
  {32'h3e680104, 32'h3eb6bc20} /* (17, 28, 5) {real, imag} */,
  {32'h3f158a9c, 32'h3fcf734a} /* (17, 28, 4) {real, imag} */,
  {32'hbe4a0dfb, 32'hbd8cee3b} /* (17, 28, 3) {real, imag} */,
  {32'hbd179372, 32'hbfe2e454} /* (17, 28, 2) {real, imag} */,
  {32'h3ec716f6, 32'hbff6c87c} /* (17, 28, 1) {real, imag} */,
  {32'hc02641f7, 32'hbf163fee} /* (17, 28, 0) {real, imag} */,
  {32'h40021842, 32'h3ed994c6} /* (17, 27, 31) {real, imag} */,
  {32'hbf2ff800, 32'hbfd336a5} /* (17, 27, 30) {real, imag} */,
  {32'h3f648615, 32'hbfefecbf} /* (17, 27, 29) {real, imag} */,
  {32'h4032b8c2, 32'h3f9cb962} /* (17, 27, 28) {real, imag} */,
  {32'hbfb4e33f, 32'h3f4affe5} /* (17, 27, 27) {real, imag} */,
  {32'hbe421711, 32'hbf0a89d7} /* (17, 27, 26) {real, imag} */,
  {32'h3f90dd03, 32'h3f895e91} /* (17, 27, 25) {real, imag} */,
  {32'h3f480d4f, 32'h3fc2930a} /* (17, 27, 24) {real, imag} */,
  {32'hbeaea8e6, 32'h3f9d38cb} /* (17, 27, 23) {real, imag} */,
  {32'hbf5e7cf6, 32'hbea51453} /* (17, 27, 22) {real, imag} */,
  {32'h3fde8c78, 32'hbfbf9953} /* (17, 27, 21) {real, imag} */,
  {32'h3ec3d7f6, 32'h3e97249b} /* (17, 27, 20) {real, imag} */,
  {32'hc00ba6d5, 32'hbf287f53} /* (17, 27, 19) {real, imag} */,
  {32'hbf86a1b3, 32'h3fdb1b70} /* (17, 27, 18) {real, imag} */,
  {32'h3de4579f, 32'hbee75335} /* (17, 27, 17) {real, imag} */,
  {32'hbf2a2ae4, 32'hbe9b5bd7} /* (17, 27, 16) {real, imag} */,
  {32'h3ebbbd94, 32'h3f9f8610} /* (17, 27, 15) {real, imag} */,
  {32'h3e4fdd5e, 32'hbf2734c6} /* (17, 27, 14) {real, imag} */,
  {32'hbf3d5626, 32'hbc9d8f7c} /* (17, 27, 13) {real, imag} */,
  {32'hbf17a806, 32'hbfdefa78} /* (17, 27, 12) {real, imag} */,
  {32'h3f180f4e, 32'hbed8df3f} /* (17, 27, 11) {real, imag} */,
  {32'h3d9853c8, 32'hbf59cb93} /* (17, 27, 10) {real, imag} */,
  {32'hbf743c27, 32'hbff6f2e7} /* (17, 27, 9) {real, imag} */,
  {32'hbf2c3305, 32'h3ec2d032} /* (17, 27, 8) {real, imag} */,
  {32'h3f7635ae, 32'hbff95e66} /* (17, 27, 7) {real, imag} */,
  {32'h4011a322, 32'h4039bcf4} /* (17, 27, 6) {real, imag} */,
  {32'h3f9ed175, 32'h3dec67df} /* (17, 27, 5) {real, imag} */,
  {32'h3f92d028, 32'hbeda007b} /* (17, 27, 4) {real, imag} */,
  {32'h3de34343, 32'hc031e6f2} /* (17, 27, 3) {real, imag} */,
  {32'h3f15a499, 32'hbf813716} /* (17, 27, 2) {real, imag} */,
  {32'h3fa7d94e, 32'h3dc77e45} /* (17, 27, 1) {real, imag} */,
  {32'h3f5d5622, 32'h3fa4903c} /* (17, 27, 0) {real, imag} */,
  {32'hbf5cb6f7, 32'hbf86598b} /* (17, 26, 31) {real, imag} */,
  {32'h3f235d0a, 32'h3f13981d} /* (17, 26, 30) {real, imag} */,
  {32'h3f780143, 32'h3f7c6ac7} /* (17, 26, 29) {real, imag} */,
  {32'h3fe85193, 32'hbe15d9f0} /* (17, 26, 28) {real, imag} */,
  {32'hbf325478, 32'hbf2c2bf0} /* (17, 26, 27) {real, imag} */,
  {32'hbfb932e6, 32'hbe0a1a79} /* (17, 26, 26) {real, imag} */,
  {32'h3eb6842a, 32'h3eb11a1d} /* (17, 26, 25) {real, imag} */,
  {32'hc0958613, 32'h3fea7693} /* (17, 26, 24) {real, imag} */,
  {32'hbeb755e4, 32'h40255697} /* (17, 26, 23) {real, imag} */,
  {32'h3d0d58a5, 32'hc030295e} /* (17, 26, 22) {real, imag} */,
  {32'h4006314f, 32'hbefc303e} /* (17, 26, 21) {real, imag} */,
  {32'hbfd806e8, 32'hbea42ecc} /* (17, 26, 20) {real, imag} */,
  {32'h3f8b7800, 32'hbfb25135} /* (17, 26, 19) {real, imag} */,
  {32'h402f6297, 32'h4005d2b5} /* (17, 26, 18) {real, imag} */,
  {32'hbdc91d3c, 32'h3e8a91d2} /* (17, 26, 17) {real, imag} */,
  {32'hbf07c162, 32'h3f0ff7f9} /* (17, 26, 16) {real, imag} */,
  {32'h3d0d74bb, 32'hbfa435bb} /* (17, 26, 15) {real, imag} */,
  {32'h3fa946af, 32'hbf7b91be} /* (17, 26, 14) {real, imag} */,
  {32'hbbd6bfd5, 32'h3fd39c02} /* (17, 26, 13) {real, imag} */,
  {32'hbeaf73d6, 32'h3f079037} /* (17, 26, 12) {real, imag} */,
  {32'h3f853853, 32'hbf98b66a} /* (17, 26, 11) {real, imag} */,
  {32'h402426e7, 32'hc010adf9} /* (17, 26, 10) {real, imag} */,
  {32'hbfaba9db, 32'h3deed12d} /* (17, 26, 9) {real, imag} */,
  {32'hbe704ee7, 32'h3fbc5eb2} /* (17, 26, 8) {real, imag} */,
  {32'hbe9c4273, 32'hbf94626b} /* (17, 26, 7) {real, imag} */,
  {32'h40466fa3, 32'hbda5294c} /* (17, 26, 6) {real, imag} */,
  {32'h3f17bd33, 32'h4019fa50} /* (17, 26, 5) {real, imag} */,
  {32'h3fa56795, 32'hbedba797} /* (17, 26, 4) {real, imag} */,
  {32'h3f1ec538, 32'hbe42eb43} /* (17, 26, 3) {real, imag} */,
  {32'h3dd027a7, 32'hbfac0cf6} /* (17, 26, 2) {real, imag} */,
  {32'hbf359da5, 32'hbeafdd15} /* (17, 26, 1) {real, imag} */,
  {32'hbf6efa69, 32'h3e672eef} /* (17, 26, 0) {real, imag} */,
  {32'h3ecbd200, 32'hc001bb38} /* (17, 25, 31) {real, imag} */,
  {32'h4023cada, 32'hbfa08160} /* (17, 25, 30) {real, imag} */,
  {32'h3f1e0f48, 32'h3e162578} /* (17, 25, 29) {real, imag} */,
  {32'h3f60e258, 32'h400e8f58} /* (17, 25, 28) {real, imag} */,
  {32'h4018f556, 32'hbda79710} /* (17, 25, 27) {real, imag} */,
  {32'hc01929af, 32'hbdbebd31} /* (17, 25, 26) {real, imag} */,
  {32'h3cd44dd7, 32'hbf91661e} /* (17, 25, 25) {real, imag} */,
  {32'hbf80c4ae, 32'h3ded44e0} /* (17, 25, 24) {real, imag} */,
  {32'h4003595f, 32'hbf9c54b7} /* (17, 25, 23) {real, imag} */,
  {32'h3fa8c5f5, 32'h402d3c02} /* (17, 25, 22) {real, imag} */,
  {32'h3f1d1d49, 32'hbf92fb41} /* (17, 25, 21) {real, imag} */,
  {32'hbf11b708, 32'h3fd07671} /* (17, 25, 20) {real, imag} */,
  {32'hbe940d52, 32'h3e21c7c6} /* (17, 25, 19) {real, imag} */,
  {32'hbf413d63, 32'h3f50ec13} /* (17, 25, 18) {real, imag} */,
  {32'h3f8a4495, 32'h3ee21f1d} /* (17, 25, 17) {real, imag} */,
  {32'h3e19b40d, 32'hbeedaea8} /* (17, 25, 16) {real, imag} */,
  {32'h3e3135da, 32'h3fc7f132} /* (17, 25, 15) {real, imag} */,
  {32'h3f2501dc, 32'hbf63d132} /* (17, 25, 14) {real, imag} */,
  {32'h404cfa0c, 32'hc00d9d29} /* (17, 25, 13) {real, imag} */,
  {32'h3fa22f4a, 32'h3f0f3db1} /* (17, 25, 12) {real, imag} */,
  {32'h3f212b0b, 32'hc0148f35} /* (17, 25, 11) {real, imag} */,
  {32'hc02187c4, 32'hbe3d41a7} /* (17, 25, 10) {real, imag} */,
  {32'hbf0d0d0c, 32'h3f91be1c} /* (17, 25, 9) {real, imag} */,
  {32'hbf113ba3, 32'h3d8de30f} /* (17, 25, 8) {real, imag} */,
  {32'hbf0ae046, 32'h3fe09af0} /* (17, 25, 7) {real, imag} */,
  {32'hc031e533, 32'hbeebad37} /* (17, 25, 6) {real, imag} */,
  {32'h3ea7c769, 32'h3d6b12c6} /* (17, 25, 5) {real, imag} */,
  {32'hbf0d6b78, 32'hbec4e1b4} /* (17, 25, 4) {real, imag} */,
  {32'hbe82d762, 32'h3f884dca} /* (17, 25, 3) {real, imag} */,
  {32'h3fd277ba, 32'hbf8581fe} /* (17, 25, 2) {real, imag} */,
  {32'hbfb283f5, 32'hc0292203} /* (17, 25, 1) {real, imag} */,
  {32'hbcf65638, 32'hbf5ad7c3} /* (17, 25, 0) {real, imag} */,
  {32'hc0204067, 32'h3ef0642c} /* (17, 24, 31) {real, imag} */,
  {32'hbf530dbc, 32'h3f8cd77e} /* (17, 24, 30) {real, imag} */,
  {32'h3f4186ff, 32'hbf09b42f} /* (17, 24, 29) {real, imag} */,
  {32'h40304003, 32'h3fb1ba58} /* (17, 24, 28) {real, imag} */,
  {32'h3ef07e2a, 32'hbf802760} /* (17, 24, 27) {real, imag} */,
  {32'hbde93bdd, 32'h3ff3ab0d} /* (17, 24, 26) {real, imag} */,
  {32'hc00aa1d7, 32'hbf3fcdde} /* (17, 24, 25) {real, imag} */,
  {32'hbf4102ba, 32'hbfd12a94} /* (17, 24, 24) {real, imag} */,
  {32'hbf81034d, 32'hbf995ac0} /* (17, 24, 23) {real, imag} */,
  {32'h3e9490d1, 32'hc023fda5} /* (17, 24, 22) {real, imag} */,
  {32'h3f3ec1e3, 32'h3f9723ba} /* (17, 24, 21) {real, imag} */,
  {32'hc002a394, 32'hbfbced59} /* (17, 24, 20) {real, imag} */,
  {32'h3f5af744, 32'h3fbd0446} /* (17, 24, 19) {real, imag} */,
  {32'h400eebb5, 32'h3f2d0998} /* (17, 24, 18) {real, imag} */,
  {32'hbf15b2b9, 32'hbf35e82b} /* (17, 24, 17) {real, imag} */,
  {32'h3fd605cf, 32'hc006c2d5} /* (17, 24, 16) {real, imag} */,
  {32'hbf2f0b56, 32'hbe524342} /* (17, 24, 15) {real, imag} */,
  {32'h3d829e20, 32'h3f58d678} /* (17, 24, 14) {real, imag} */,
  {32'hbe9d191e, 32'hbeb7347f} /* (17, 24, 13) {real, imag} */,
  {32'h402adb74, 32'hbf804e27} /* (17, 24, 12) {real, imag} */,
  {32'h3f8182ec, 32'hbee5e11e} /* (17, 24, 11) {real, imag} */,
  {32'h40283bd5, 32'hbf7ec185} /* (17, 24, 10) {real, imag} */,
  {32'hbf9ba4b9, 32'hc00c7eeb} /* (17, 24, 9) {real, imag} */,
  {32'hbf7dc052, 32'h3ffe8f63} /* (17, 24, 8) {real, imag} */,
  {32'hbf9cd591, 32'h3fba7fe9} /* (17, 24, 7) {real, imag} */,
  {32'h3ffdba9d, 32'hbfd24c30} /* (17, 24, 6) {real, imag} */,
  {32'h3f7d36d1, 32'hbf989a90} /* (17, 24, 5) {real, imag} */,
  {32'h3fcc16b1, 32'hc024024a} /* (17, 24, 4) {real, imag} */,
  {32'h3d90db44, 32'h3fc18cd1} /* (17, 24, 3) {real, imag} */,
  {32'hbc33f99e, 32'h3e405812} /* (17, 24, 2) {real, imag} */,
  {32'h3ebb9430, 32'h3f01584e} /* (17, 24, 1) {real, imag} */,
  {32'hc00c5ef2, 32'hbda3951c} /* (17, 24, 0) {real, imag} */,
  {32'h3fad3d25, 32'hbf881d68} /* (17, 23, 31) {real, imag} */,
  {32'h3f08a465, 32'h3fddef9c} /* (17, 23, 30) {real, imag} */,
  {32'h3f8e3304, 32'h3f6cd11a} /* (17, 23, 29) {real, imag} */,
  {32'hbeb6f2cc, 32'h3fb8962d} /* (17, 23, 28) {real, imag} */,
  {32'h3d99db9a, 32'h3f62b68c} /* (17, 23, 27) {real, imag} */,
  {32'h3f5288ae, 32'hc042b90f} /* (17, 23, 26) {real, imag} */,
  {32'h3f9a67c0, 32'h3e86a3f4} /* (17, 23, 25) {real, imag} */,
  {32'hc030eac2, 32'h3fac0093} /* (17, 23, 24) {real, imag} */,
  {32'h3fc5e4ea, 32'hc044d7a9} /* (17, 23, 23) {real, imag} */,
  {32'h40a21176, 32'h3fc5fa82} /* (17, 23, 22) {real, imag} */,
  {32'hbfb9c1e1, 32'h3f8f0399} /* (17, 23, 21) {real, imag} */,
  {32'hc024f651, 32'h3f481bbe} /* (17, 23, 20) {real, imag} */,
  {32'h3f36bde7, 32'hbfbdd018} /* (17, 23, 19) {real, imag} */,
  {32'hbfb6ebb5, 32'hc0389686} /* (17, 23, 18) {real, imag} */,
  {32'hbfc57c84, 32'h3fc8cac5} /* (17, 23, 17) {real, imag} */,
  {32'hbf9bccc3, 32'h3f3fb4ef} /* (17, 23, 16) {real, imag} */,
  {32'hbf75dfff, 32'h3f3b5ac3} /* (17, 23, 15) {real, imag} */,
  {32'h3d7b0c7b, 32'hbf67ce9a} /* (17, 23, 14) {real, imag} */,
  {32'hbe972fbc, 32'hbf4a24d0} /* (17, 23, 13) {real, imag} */,
  {32'hbda4c377, 32'hbfd7f5fa} /* (17, 23, 12) {real, imag} */,
  {32'hc066e4b5, 32'hbfdaec09} /* (17, 23, 11) {real, imag} */,
  {32'h4035d26f, 32'h40611c8d} /* (17, 23, 10) {real, imag} */,
  {32'h3f68ef4b, 32'hbfb0ad67} /* (17, 23, 9) {real, imag} */,
  {32'hc030d404, 32'hbff48199} /* (17, 23, 8) {real, imag} */,
  {32'hbf107692, 32'hbd50c231} /* (17, 23, 7) {real, imag} */,
  {32'h3e9179c8, 32'h3f0dfbaf} /* (17, 23, 6) {real, imag} */,
  {32'h4010c440, 32'hbf21f712} /* (17, 23, 5) {real, imag} */,
  {32'h3cde9d9e, 32'h3f80cddc} /* (17, 23, 4) {real, imag} */,
  {32'hbef92fb9, 32'hbeabf1f7} /* (17, 23, 3) {real, imag} */,
  {32'h3d95bfeb, 32'h3f2df189} /* (17, 23, 2) {real, imag} */,
  {32'h3dd60c17, 32'hbf80ff19} /* (17, 23, 1) {real, imag} */,
  {32'h3ebd4a2c, 32'hbd87d0a0} /* (17, 23, 0) {real, imag} */,
  {32'hbf4780f8, 32'hbf0f4819} /* (17, 22, 31) {real, imag} */,
  {32'h3e35066f, 32'h3f535d62} /* (17, 22, 30) {real, imag} */,
  {32'h3d0bf12f, 32'h3f0a7b98} /* (17, 22, 29) {real, imag} */,
  {32'hbf09cc7c, 32'hc002af5d} /* (17, 22, 28) {real, imag} */,
  {32'h3eae187d, 32'h3f88e980} /* (17, 22, 27) {real, imag} */,
  {32'h3faee526, 32'hbfdde08c} /* (17, 22, 26) {real, imag} */,
  {32'hbf6646d9, 32'hbf06d65e} /* (17, 22, 25) {real, imag} */,
  {32'hbfbf3972, 32'hbf1dc051} /* (17, 22, 24) {real, imag} */,
  {32'h3faa0cdc, 32'h3f1caf45} /* (17, 22, 23) {real, imag} */,
  {32'hbe7609b9, 32'hc02451c6} /* (17, 22, 22) {real, imag} */,
  {32'hbf3c92eb, 32'hbe854c91} /* (17, 22, 21) {real, imag} */,
  {32'hbedfce88, 32'hbff92f50} /* (17, 22, 20) {real, imag} */,
  {32'h3fab3c24, 32'h40301054} /* (17, 22, 19) {real, imag} */,
  {32'hbf6aedfc, 32'h3fc7794d} /* (17, 22, 18) {real, imag} */,
  {32'hbf9fb915, 32'h39f5034f} /* (17, 22, 17) {real, imag} */,
  {32'h3f9e5c0c, 32'h3f433aa2} /* (17, 22, 16) {real, imag} */,
  {32'hbfbc2dd2, 32'hbee4d273} /* (17, 22, 15) {real, imag} */,
  {32'hbfc5c551, 32'hbf34f63f} /* (17, 22, 14) {real, imag} */,
  {32'h3f81c1e8, 32'h3e8bb785} /* (17, 22, 13) {real, imag} */,
  {32'h3fdc15fc, 32'hbfc618e7} /* (17, 22, 12) {real, imag} */,
  {32'h3e37731c, 32'hbe20a966} /* (17, 22, 11) {real, imag} */,
  {32'hc08441c2, 32'h3f99f0f8} /* (17, 22, 10) {real, imag} */,
  {32'h3ff946e7, 32'h4043e999} /* (17, 22, 9) {real, imag} */,
  {32'hbf4a9c2d, 32'hbf576ce0} /* (17, 22, 8) {real, imag} */,
  {32'hbf814f3a, 32'h40230f28} /* (17, 22, 7) {real, imag} */,
  {32'h3ee1d165, 32'hbfacec80} /* (17, 22, 6) {real, imag} */,
  {32'h3ed12325, 32'hbfe4557b} /* (17, 22, 5) {real, imag} */,
  {32'h3e3ef23f, 32'hbf1f0c25} /* (17, 22, 4) {real, imag} */,
  {32'hbefb5f9a, 32'h3f278ea5} /* (17, 22, 3) {real, imag} */,
  {32'h40000ffc, 32'h3f474254} /* (17, 22, 2) {real, imag} */,
  {32'h3ebe31df, 32'hbf8f7d11} /* (17, 22, 1) {real, imag} */,
  {32'hbf877d26, 32'h3d3dd9af} /* (17, 22, 0) {real, imag} */,
  {32'h3f97baea, 32'hbeff5def} /* (17, 21, 31) {real, imag} */,
  {32'h3e9a2d46, 32'hbe8319df} /* (17, 21, 30) {real, imag} */,
  {32'hbc32bfd6, 32'h3f452b86} /* (17, 21, 29) {real, imag} */,
  {32'hbf8400b5, 32'h400239cc} /* (17, 21, 28) {real, imag} */,
  {32'h3ffc03bb, 32'h3f8cb294} /* (17, 21, 27) {real, imag} */,
  {32'h3fed63c3, 32'hbedfd32b} /* (17, 21, 26) {real, imag} */,
  {32'h3fd7d298, 32'hbe9d646e} /* (17, 21, 25) {real, imag} */,
  {32'hc01fb69d, 32'h400bd21d} /* (17, 21, 24) {real, imag} */,
  {32'h3fe21964, 32'h3e8631f8} /* (17, 21, 23) {real, imag} */,
  {32'hbda1fbc0, 32'hbf02ca73} /* (17, 21, 22) {real, imag} */,
  {32'hbe9ed564, 32'hbe16bb8e} /* (17, 21, 21) {real, imag} */,
  {32'hbfbe6dda, 32'hc03e2198} /* (17, 21, 20) {real, imag} */,
  {32'h3f4e9ca7, 32'h3f3bbb43} /* (17, 21, 19) {real, imag} */,
  {32'h3fb9c087, 32'h3ca8524b} /* (17, 21, 18) {real, imag} */,
  {32'h3ed875c3, 32'h3e8f87b9} /* (17, 21, 17) {real, imag} */,
  {32'h3fd49f9d, 32'h40204059} /* (17, 21, 16) {real, imag} */,
  {32'h3e4fb0e9, 32'h3f8bdf5d} /* (17, 21, 15) {real, imag} */,
  {32'h3f23edac, 32'h3e30ba42} /* (17, 21, 14) {real, imag} */,
  {32'hbf26970b, 32'hc04dd0f5} /* (17, 21, 13) {real, imag} */,
  {32'h3fcf7a34, 32'h3ea4ef30} /* (17, 21, 12) {real, imag} */,
  {32'hbfcbe7d6, 32'h3e8c58cc} /* (17, 21, 11) {real, imag} */,
  {32'hc04368b2, 32'h3ddba86b} /* (17, 21, 10) {real, imag} */,
  {32'hbffa2d4f, 32'hbfa3b680} /* (17, 21, 9) {real, imag} */,
  {32'hbefbf9dc, 32'hbfd75cf7} /* (17, 21, 8) {real, imag} */,
  {32'h400fd44c, 32'h3f576ab8} /* (17, 21, 7) {real, imag} */,
  {32'hbecefc1f, 32'hbd5a3489} /* (17, 21, 6) {real, imag} */,
  {32'hbf2f1284, 32'h3c76992c} /* (17, 21, 5) {real, imag} */,
  {32'hbfb410d6, 32'h3e5279d4} /* (17, 21, 4) {real, imag} */,
  {32'h3f9bdd8d, 32'hbfa7c11d} /* (17, 21, 3) {real, imag} */,
  {32'h3e35ec1c, 32'h3f250c5f} /* (17, 21, 2) {real, imag} */,
  {32'hbdd07711, 32'hbfb0e1e6} /* (17, 21, 1) {real, imag} */,
  {32'h3f0be871, 32'hbf9c09ac} /* (17, 21, 0) {real, imag} */,
  {32'h3f9002f0, 32'h3ec10439} /* (17, 20, 31) {real, imag} */,
  {32'h3fcea723, 32'h3f8c0494} /* (17, 20, 30) {real, imag} */,
  {32'h3f263f8f, 32'hbd57c749} /* (17, 20, 29) {real, imag} */,
  {32'hbfae3142, 32'h3f3f9018} /* (17, 20, 28) {real, imag} */,
  {32'hbfb278b1, 32'h3f1b6c7f} /* (17, 20, 27) {real, imag} */,
  {32'h3f435f1a, 32'hbe8fd109} /* (17, 20, 26) {real, imag} */,
  {32'hbfad1628, 32'h3f563def} /* (17, 20, 25) {real, imag} */,
  {32'h3fe35e09, 32'h3ed41abe} /* (17, 20, 24) {real, imag} */,
  {32'hbfa12c67, 32'hbf919de3} /* (17, 20, 23) {real, imag} */,
  {32'hc003d7fd, 32'h3fa1dc66} /* (17, 20, 22) {real, imag} */,
  {32'hbe14d744, 32'hbf289cb4} /* (17, 20, 21) {real, imag} */,
  {32'hbd69df9d, 32'hbf954007} /* (17, 20, 20) {real, imag} */,
  {32'h3d8d5b65, 32'h3e2e446f} /* (17, 20, 19) {real, imag} */,
  {32'hbfbfa723, 32'hbf45a9ee} /* (17, 20, 18) {real, imag} */,
  {32'hbe975d36, 32'h3e4c615f} /* (17, 20, 17) {real, imag} */,
  {32'hbf39dcd8, 32'hbfb8dbb8} /* (17, 20, 16) {real, imag} */,
  {32'h3d4f05d1, 32'hc071c512} /* (17, 20, 15) {real, imag} */,
  {32'hbfcf3310, 32'h3c531847} /* (17, 20, 14) {real, imag} */,
  {32'hbf8ef5b7, 32'hbfb40197} /* (17, 20, 13) {real, imag} */,
  {32'h3fa16104, 32'h4040abaa} /* (17, 20, 12) {real, imag} */,
  {32'hbf074c66, 32'hbfa35863} /* (17, 20, 11) {real, imag} */,
  {32'h4006c83b, 32'hbf8c32d0} /* (17, 20, 10) {real, imag} */,
  {32'h3fa1d28d, 32'h3fc11ce8} /* (17, 20, 9) {real, imag} */,
  {32'hbed0107a, 32'hbff67126} /* (17, 20, 8) {real, imag} */,
  {32'hbf49a285, 32'h3fa0e150} /* (17, 20, 7) {real, imag} */,
  {32'h3fab1f41, 32'hbd7b627b} /* (17, 20, 6) {real, imag} */,
  {32'h4020abf1, 32'hbf3b8e51} /* (17, 20, 5) {real, imag} */,
  {32'h3f221a34, 32'hbf523211} /* (17, 20, 4) {real, imag} */,
  {32'hbf0c149f, 32'h3fb5423f} /* (17, 20, 3) {real, imag} */,
  {32'h3f7a5f6a, 32'h3e671479} /* (17, 20, 2) {real, imag} */,
  {32'h40521d81, 32'h3d873841} /* (17, 20, 1) {real, imag} */,
  {32'hbfe919db, 32'hbf983312} /* (17, 20, 0) {real, imag} */,
  {32'hbfd38ad5, 32'hbd8d15a6} /* (17, 19, 31) {real, imag} */,
  {32'hc0642a50, 32'hbea9d4f0} /* (17, 19, 30) {real, imag} */,
  {32'h3f504942, 32'h3edc1c8b} /* (17, 19, 29) {real, imag} */,
  {32'hbd6e79b0, 32'h3fc34751} /* (17, 19, 28) {real, imag} */,
  {32'h3d7396e3, 32'hbf682e73} /* (17, 19, 27) {real, imag} */,
  {32'h3f761154, 32'h4006c4ee} /* (17, 19, 26) {real, imag} */,
  {32'hbf0ea01b, 32'h3f1ae39f} /* (17, 19, 25) {real, imag} */,
  {32'hbf3d1c68, 32'hbfe9f1f9} /* (17, 19, 24) {real, imag} */,
  {32'h400befd9, 32'h40089207} /* (17, 19, 23) {real, imag} */,
  {32'hbf8ea908, 32'hbed16994} /* (17, 19, 22) {real, imag} */,
  {32'h3ff5af9c, 32'h3f9a14ce} /* (17, 19, 21) {real, imag} */,
  {32'hc02d59b1, 32'hbf7e3321} /* (17, 19, 20) {real, imag} */,
  {32'hc01f1e0f, 32'hbf99515d} /* (17, 19, 19) {real, imag} */,
  {32'hbf44e223, 32'hc0580dc2} /* (17, 19, 18) {real, imag} */,
  {32'h404cb7dc, 32'h3f9ecc8f} /* (17, 19, 17) {real, imag} */,
  {32'h3f40feec, 32'hbde96145} /* (17, 19, 16) {real, imag} */,
  {32'hbf61f115, 32'hbfc7bd4c} /* (17, 19, 15) {real, imag} */,
  {32'hbdbb8691, 32'hc028c3c8} /* (17, 19, 14) {real, imag} */,
  {32'hc01f1735, 32'h3f9b2411} /* (17, 19, 13) {real, imag} */,
  {32'hbf4df0fa, 32'hbf738c78} /* (17, 19, 12) {real, imag} */,
  {32'hbfb6a79f, 32'h3eba72f3} /* (17, 19, 11) {real, imag} */,
  {32'h3ecc6795, 32'h3ffcf389} /* (17, 19, 10) {real, imag} */,
  {32'hc019f1d1, 32'h3ed7653a} /* (17, 19, 9) {real, imag} */,
  {32'hbe44e2b5, 32'hbfcd620b} /* (17, 19, 8) {real, imag} */,
  {32'hbf84cf29, 32'hbf10bf81} /* (17, 19, 7) {real, imag} */,
  {32'h3f4b3170, 32'h3f399954} /* (17, 19, 6) {real, imag} */,
  {32'h3ee86266, 32'h3f46e29e} /* (17, 19, 5) {real, imag} */,
  {32'h3fe3e333, 32'hbe99ec60} /* (17, 19, 4) {real, imag} */,
  {32'h3ba5ccd3, 32'h3f928a17} /* (17, 19, 3) {real, imag} */,
  {32'h3e41a2c5, 32'h3ff3efcd} /* (17, 19, 2) {real, imag} */,
  {32'hbfb64e74, 32'hbf3e2124} /* (17, 19, 1) {real, imag} */,
  {32'h3ec059e0, 32'hbf881b32} /* (17, 19, 0) {real, imag} */,
  {32'h3f1581e5, 32'hbdae8ea7} /* (17, 18, 31) {real, imag} */,
  {32'hbfd0f96f, 32'hbdcc51f1} /* (17, 18, 30) {real, imag} */,
  {32'hc00c5f10, 32'h3e457107} /* (17, 18, 29) {real, imag} */,
  {32'h3f64bb65, 32'h3fac4e49} /* (17, 18, 28) {real, imag} */,
  {32'hbf16399e, 32'h400d0354} /* (17, 18, 27) {real, imag} */,
  {32'hbe442a96, 32'hbee99ba8} /* (17, 18, 26) {real, imag} */,
  {32'h3f11f96b, 32'h3f3246fb} /* (17, 18, 25) {real, imag} */,
  {32'h3d463271, 32'h3f474438} /* (17, 18, 24) {real, imag} */,
  {32'h3fc896dc, 32'hc028e5b1} /* (17, 18, 23) {real, imag} */,
  {32'hbf8629b3, 32'hbfbec190} /* (17, 18, 22) {real, imag} */,
  {32'hbf91815b, 32'h3f8bdd56} /* (17, 18, 21) {real, imag} */,
  {32'h3fea7b96, 32'h3f540dc1} /* (17, 18, 20) {real, imag} */,
  {32'h3ed97a86, 32'hbfa4f4f8} /* (17, 18, 19) {real, imag} */,
  {32'hbf4cc461, 32'hbf51ee42} /* (17, 18, 18) {real, imag} */,
  {32'h3f838c8a, 32'h3f57b36c} /* (17, 18, 17) {real, imag} */,
  {32'hbf9436ec, 32'h40392c68} /* (17, 18, 16) {real, imag} */,
  {32'hbf954ea5, 32'h3f33d0e1} /* (17, 18, 15) {real, imag} */,
  {32'hbeabe2d7, 32'hc016cce8} /* (17, 18, 14) {real, imag} */,
  {32'hbe9e00fd, 32'h3fcfbdfd} /* (17, 18, 13) {real, imag} */,
  {32'hbffa47c4, 32'h3f0cdb72} /* (17, 18, 12) {real, imag} */,
  {32'hbea28f52, 32'hbd95a785} /* (17, 18, 11) {real, imag} */,
  {32'hbea11d23, 32'h3f16ca66} /* (17, 18, 10) {real, imag} */,
  {32'h3ff00672, 32'h3d11992c} /* (17, 18, 9) {real, imag} */,
  {32'h3c46abe8, 32'hbff35a72} /* (17, 18, 8) {real, imag} */,
  {32'hbfbe31a9, 32'h3f8b3d7a} /* (17, 18, 7) {real, imag} */,
  {32'hbf719a57, 32'h3f9e9e2d} /* (17, 18, 6) {real, imag} */,
  {32'h3f036c51, 32'h400c970e} /* (17, 18, 5) {real, imag} */,
  {32'hbe4b9d03, 32'hbf69fb6c} /* (17, 18, 4) {real, imag} */,
  {32'h3f4c7450, 32'h3ebc7a7e} /* (17, 18, 3) {real, imag} */,
  {32'hbea865ce, 32'hc0111660} /* (17, 18, 2) {real, imag} */,
  {32'h3de7c1b5, 32'hbedac20f} /* (17, 18, 1) {real, imag} */,
  {32'h3fc3a815, 32'h4008487d} /* (17, 18, 0) {real, imag} */,
  {32'hbe88a4af, 32'hbf8a64d6} /* (17, 17, 31) {real, imag} */,
  {32'hbf389339, 32'hbf2d2713} /* (17, 17, 30) {real, imag} */,
  {32'hbda79712, 32'h3e2a6a0f} /* (17, 17, 29) {real, imag} */,
  {32'h3ee2c9ca, 32'h3b3b4718} /* (17, 17, 28) {real, imag} */,
  {32'h3f38d8c5, 32'h3fbfb675} /* (17, 17, 27) {real, imag} */,
  {32'h3f09ca02, 32'hc0200bab} /* (17, 17, 26) {real, imag} */,
  {32'hbed3772f, 32'h3f13ca60} /* (17, 17, 25) {real, imag} */,
  {32'h3e5ddb7c, 32'h3f46e9a3} /* (17, 17, 24) {real, imag} */,
  {32'hbeb936c1, 32'hbf0ecb63} /* (17, 17, 23) {real, imag} */,
  {32'h40106f63, 32'hbfe84fcc} /* (17, 17, 22) {real, imag} */,
  {32'hbfcffed4, 32'hbf9137b2} /* (17, 17, 21) {real, imag} */,
  {32'h4007bf40, 32'hc0035647} /* (17, 17, 20) {real, imag} */,
  {32'h3f44afcf, 32'hbf3e0379} /* (17, 17, 19) {real, imag} */,
  {32'h3fc88157, 32'h3f7231e9} /* (17, 17, 18) {real, imag} */,
  {32'h3f11e700, 32'hc011a27f} /* (17, 17, 17) {real, imag} */,
  {32'h3ea87420, 32'h3d54109e} /* (17, 17, 16) {real, imag} */,
  {32'h3f2b9dee, 32'h3f40017d} /* (17, 17, 15) {real, imag} */,
  {32'h3f140607, 32'hc0044865} /* (17, 17, 14) {real, imag} */,
  {32'h3f0c30c8, 32'hbf662bd1} /* (17, 17, 13) {real, imag} */,
  {32'h4006bc8d, 32'h3f1ea21e} /* (17, 17, 12) {real, imag} */,
  {32'hbfca4d88, 32'h3fed7d75} /* (17, 17, 11) {real, imag} */,
  {32'hbf941632, 32'h3ec55b8a} /* (17, 17, 10) {real, imag} */,
  {32'h3e2e3c78, 32'hbf80eb96} /* (17, 17, 9) {real, imag} */,
  {32'h3eb003e1, 32'h3f7b24fd} /* (17, 17, 8) {real, imag} */,
  {32'h3fa6b95b, 32'hbfeef3d1} /* (17, 17, 7) {real, imag} */,
  {32'hbeae9ac4, 32'hbf2cf335} /* (17, 17, 6) {real, imag} */,
  {32'h3fb4522b, 32'hbf831669} /* (17, 17, 5) {real, imag} */,
  {32'h3f0438df, 32'h3f53ef1e} /* (17, 17, 4) {real, imag} */,
  {32'h3f1756f2, 32'hbf2ac46d} /* (17, 17, 3) {real, imag} */,
  {32'hbda808a2, 32'hbe1f295f} /* (17, 17, 2) {real, imag} */,
  {32'hbe4716d9, 32'h3f28e0ec} /* (17, 17, 1) {real, imag} */,
  {32'hbe51b948, 32'h3edb8a09} /* (17, 17, 0) {real, imag} */,
  {32'h3ef86493, 32'hbf093b34} /* (17, 16, 31) {real, imag} */,
  {32'h3ed4646e, 32'hbf345219} /* (17, 16, 30) {real, imag} */,
  {32'h3e91331c, 32'h3fbe2009} /* (17, 16, 29) {real, imag} */,
  {32'h3e9960aa, 32'hbf104c73} /* (17, 16, 28) {real, imag} */,
  {32'h3f9cb468, 32'hbfe1f0e2} /* (17, 16, 27) {real, imag} */,
  {32'h3fada164, 32'h3e84bf07} /* (17, 16, 26) {real, imag} */,
  {32'hbf01d9b4, 32'h3f4a7a59} /* (17, 16, 25) {real, imag} */,
  {32'h3fd58bd4, 32'h3f0bd83e} /* (17, 16, 24) {real, imag} */,
  {32'hbfabfbf6, 32'hbed05d3a} /* (17, 16, 23) {real, imag} */,
  {32'h3f2d3b0f, 32'hc048c6ab} /* (17, 16, 22) {real, imag} */,
  {32'h3f032379, 32'h404a3ec7} /* (17, 16, 21) {real, imag} */,
  {32'hbfa5e1f1, 32'h3fc3f12d} /* (17, 16, 20) {real, imag} */,
  {32'hbfd0ce89, 32'h3f70d3d8} /* (17, 16, 19) {real, imag} */,
  {32'hbfcc4354, 32'hbfee2f3d} /* (17, 16, 18) {real, imag} */,
  {32'hbee7db82, 32'h3e0d04b4} /* (17, 16, 17) {real, imag} */,
  {32'h3f09eccd, 32'hbe07173b} /* (17, 16, 16) {real, imag} */,
  {32'hbef4b215, 32'hbdf0fcee} /* (17, 16, 15) {real, imag} */,
  {32'hbebd16fc, 32'hbe9a5c26} /* (17, 16, 14) {real, imag} */,
  {32'h3fda4479, 32'h3fbdbd4f} /* (17, 16, 13) {real, imag} */,
  {32'h3f548705, 32'hbf7ca1e0} /* (17, 16, 12) {real, imag} */,
  {32'hbf00ffed, 32'hbe15344e} /* (17, 16, 11) {real, imag} */,
  {32'h40679505, 32'h4005af35} /* (17, 16, 10) {real, imag} */,
  {32'hbd89138b, 32'h4033ee4e} /* (17, 16, 9) {real, imag} */,
  {32'hbf86259c, 32'h3f7b9aa5} /* (17, 16, 8) {real, imag} */,
  {32'hbf6fdf5a, 32'hbd5ae745} /* (17, 16, 7) {real, imag} */,
  {32'hbf4a970a, 32'hbfa8501c} /* (17, 16, 6) {real, imag} */,
  {32'hbf1f4fad, 32'h3f6c237d} /* (17, 16, 5) {real, imag} */,
  {32'hbfa19092, 32'h3f568133} /* (17, 16, 4) {real, imag} */,
  {32'hbf00faed, 32'h3fc9df37} /* (17, 16, 3) {real, imag} */,
  {32'hbe74be81, 32'h3e68f6df} /* (17, 16, 2) {real, imag} */,
  {32'hbf8fcb91, 32'h3c43f24b} /* (17, 16, 1) {real, imag} */,
  {32'h3e87912a, 32'hbf147917} /* (17, 16, 0) {real, imag} */,
  {32'h3f3aa1c0, 32'hbfcb3911} /* (17, 15, 31) {real, imag} */,
  {32'hbf0bb2d3, 32'h3e7adb79} /* (17, 15, 30) {real, imag} */,
  {32'h3f35ed42, 32'h3d46bcae} /* (17, 15, 29) {real, imag} */,
  {32'hbe88d8af, 32'hbe113eeb} /* (17, 15, 28) {real, imag} */,
  {32'h3d1c43fe, 32'h3e679f2d} /* (17, 15, 27) {real, imag} */,
  {32'h3f494566, 32'h3ea46778} /* (17, 15, 26) {real, imag} */,
  {32'hc0156461, 32'h3ec64132} /* (17, 15, 25) {real, imag} */,
  {32'hbecd6073, 32'h3ed0898d} /* (17, 15, 24) {real, imag} */,
  {32'hbf0dbf8e, 32'h3ef711fd} /* (17, 15, 23) {real, imag} */,
  {32'hc01b6603, 32'hbeef8fce} /* (17, 15, 22) {real, imag} */,
  {32'hbf7e4f95, 32'h3ee499b1} /* (17, 15, 21) {real, imag} */,
  {32'h4086ae75, 32'hbfda8d42} /* (17, 15, 20) {real, imag} */,
  {32'h3f88ebbb, 32'hbffc49ba} /* (17, 15, 19) {real, imag} */,
  {32'h3fa68fa9, 32'h3e5f0950} /* (17, 15, 18) {real, imag} */,
  {32'h3fd4df10, 32'h3f2b384d} /* (17, 15, 17) {real, imag} */,
  {32'h3fbb0b88, 32'h3ee515be} /* (17, 15, 16) {real, imag} */,
  {32'h3f2d6686, 32'h3f2d2985} /* (17, 15, 15) {real, imag} */,
  {32'hc00fa97e, 32'h3ed80984} /* (17, 15, 14) {real, imag} */,
  {32'hbe503562, 32'h3e9d7e23} /* (17, 15, 13) {real, imag} */,
  {32'hbf6573cd, 32'hbeeab455} /* (17, 15, 12) {real, imag} */,
  {32'hbf237865, 32'hbf044da4} /* (17, 15, 11) {real, imag} */,
  {32'hbe2e41db, 32'hc037320c} /* (17, 15, 10) {real, imag} */,
  {32'hc018d817, 32'hbe5735ce} /* (17, 15, 9) {real, imag} */,
  {32'h3d5803e5, 32'h3fbca45a} /* (17, 15, 8) {real, imag} */,
  {32'hbddb760c, 32'hbf8ab28d} /* (17, 15, 7) {real, imag} */,
  {32'h3f013a85, 32'hbf1be958} /* (17, 15, 6) {real, imag} */,
  {32'h3d6db068, 32'h3fab368f} /* (17, 15, 5) {real, imag} */,
  {32'hbc883c33, 32'h3f0a0189} /* (17, 15, 4) {real, imag} */,
  {32'h3d8fac24, 32'hbf3eedd9} /* (17, 15, 3) {real, imag} */,
  {32'h3f459058, 32'hbe05b820} /* (17, 15, 2) {real, imag} */,
  {32'hbf491c66, 32'hbfa1ebe7} /* (17, 15, 1) {real, imag} */,
  {32'hbda5e566, 32'hbf994b53} /* (17, 15, 0) {real, imag} */,
  {32'h4002fbab, 32'hbf484660} /* (17, 14, 31) {real, imag} */,
  {32'h3fce0736, 32'h3f2e3983} /* (17, 14, 30) {real, imag} */,
  {32'hbf717369, 32'h3f7ae1fc} /* (17, 14, 29) {real, imag} */,
  {32'hbdff37b3, 32'h3f858a4c} /* (17, 14, 28) {real, imag} */,
  {32'h400f85f1, 32'hbfa916ad} /* (17, 14, 27) {real, imag} */,
  {32'h3f82e67a, 32'h3ffe363d} /* (17, 14, 26) {real, imag} */,
  {32'h402b5083, 32'h40018a88} /* (17, 14, 25) {real, imag} */,
  {32'h3dadb7df, 32'h3faa0d35} /* (17, 14, 24) {real, imag} */,
  {32'hbf9d7c03, 32'h3fb83bb6} /* (17, 14, 23) {real, imag} */,
  {32'h3f266544, 32'h40147e59} /* (17, 14, 22) {real, imag} */,
  {32'h3e5074d9, 32'h402f2346} /* (17, 14, 21) {real, imag} */,
  {32'h3e8cb6a3, 32'h3def2b7f} /* (17, 14, 20) {real, imag} */,
  {32'hbf14c2d6, 32'hbe3ff145} /* (17, 14, 19) {real, imag} */,
  {32'hbf8de6d0, 32'hbfb0ec08} /* (17, 14, 18) {real, imag} */,
  {32'h3f696000, 32'hbf0864bc} /* (17, 14, 17) {real, imag} */,
  {32'hbf9409b4, 32'h3f39c46d} /* (17, 14, 16) {real, imag} */,
  {32'hc06d59cb, 32'hbfd94931} /* (17, 14, 15) {real, imag} */,
  {32'h3f907ed9, 32'h3ed7ad48} /* (17, 14, 14) {real, imag} */,
  {32'hc0741b59, 32'hc000ab8b} /* (17, 14, 13) {real, imag} */,
  {32'hbe45ecf3, 32'hc02ba0fe} /* (17, 14, 12) {real, imag} */,
  {32'h400fa60c, 32'hbf5a48e1} /* (17, 14, 11) {real, imag} */,
  {32'hbe855a89, 32'h3fbaf4b0} /* (17, 14, 10) {real, imag} */,
  {32'hbf124101, 32'h3e8d2981} /* (17, 14, 9) {real, imag} */,
  {32'h3f9748d6, 32'h3fb2ae5d} /* (17, 14, 8) {real, imag} */,
  {32'h4062f1f0, 32'hbd95ce8a} /* (17, 14, 7) {real, imag} */,
  {32'h3fffcd49, 32'hbe9e4032} /* (17, 14, 6) {real, imag} */,
  {32'h3eaed351, 32'hbf014ca6} /* (17, 14, 5) {real, imag} */,
  {32'h3fc47fbe, 32'hbfc0bbb8} /* (17, 14, 4) {real, imag} */,
  {32'hbe3af8c6, 32'hbe6921df} /* (17, 14, 3) {real, imag} */,
  {32'h3fc53dac, 32'hbf1a4c90} /* (17, 14, 2) {real, imag} */,
  {32'h3e6e6c19, 32'hbdb63b47} /* (17, 14, 1) {real, imag} */,
  {32'h3c1a3ae0, 32'h3f7a54e1} /* (17, 14, 0) {real, imag} */,
  {32'h3f36b338, 32'h3ec8d049} /* (17, 13, 31) {real, imag} */,
  {32'hbf904c04, 32'hbf209d44} /* (17, 13, 30) {real, imag} */,
  {32'hbf94c86a, 32'hbf420701} /* (17, 13, 29) {real, imag} */,
  {32'hbf237542, 32'hbff80ce8} /* (17, 13, 28) {real, imag} */,
  {32'h3f36ecf8, 32'h3febc7b1} /* (17, 13, 27) {real, imag} */,
  {32'h3ec8a7af, 32'hbe9cf5de} /* (17, 13, 26) {real, imag} */,
  {32'h3f83452d, 32'h3e97e3ec} /* (17, 13, 25) {real, imag} */,
  {32'h3ff7eb60, 32'hbfc2207b} /* (17, 13, 24) {real, imag} */,
  {32'h3f8df10b, 32'hbf411431} /* (17, 13, 23) {real, imag} */,
  {32'h3f1d4e25, 32'hc0334e00} /* (17, 13, 22) {real, imag} */,
  {32'h3fb68174, 32'h3dde077a} /* (17, 13, 21) {real, imag} */,
  {32'h3c87dfe1, 32'hbf742cdb} /* (17, 13, 20) {real, imag} */,
  {32'hc02013d6, 32'h40808730} /* (17, 13, 19) {real, imag} */,
  {32'hbfb79ff7, 32'h3f859161} /* (17, 13, 18) {real, imag} */,
  {32'hc0322d8d, 32'h3f929f5b} /* (17, 13, 17) {real, imag} */,
  {32'h3ecafbf8, 32'h3ed689cd} /* (17, 13, 16) {real, imag} */,
  {32'h3fdd5f44, 32'hbfc63948} /* (17, 13, 15) {real, imag} */,
  {32'hc0302bfe, 32'hc00f83a3} /* (17, 13, 14) {real, imag} */,
  {32'h3ea27233, 32'h3f70758c} /* (17, 13, 13) {real, imag} */,
  {32'hbecdef43, 32'hc034e5ce} /* (17, 13, 12) {real, imag} */,
  {32'hbf1ba8e3, 32'hbf76ce27} /* (17, 13, 11) {real, imag} */,
  {32'hbef181ca, 32'hbf7a8113} /* (17, 13, 10) {real, imag} */,
  {32'hbfc40de5, 32'h3e4a9699} /* (17, 13, 9) {real, imag} */,
  {32'h3feadde4, 32'h3f2775b4} /* (17, 13, 8) {real, imag} */,
  {32'h3f618bce, 32'h3e93d20d} /* (17, 13, 7) {real, imag} */,
  {32'h3f11e974, 32'hc037adf5} /* (17, 13, 6) {real, imag} */,
  {32'hbe615c93, 32'hbf7ace13} /* (17, 13, 5) {real, imag} */,
  {32'hbc212c0f, 32'hbfb5568d} /* (17, 13, 4) {real, imag} */,
  {32'hbeb946f8, 32'h3f90983a} /* (17, 13, 3) {real, imag} */,
  {32'h3f2a7329, 32'h3ffda5fc} /* (17, 13, 2) {real, imag} */,
  {32'h3fd645f2, 32'h3f658874} /* (17, 13, 1) {real, imag} */,
  {32'hbe6591e2, 32'hbeda4732} /* (17, 13, 0) {real, imag} */,
  {32'hbf97861c, 32'h3fc345d1} /* (17, 12, 31) {real, imag} */,
  {32'hbfa3ad86, 32'h3f3a9312} /* (17, 12, 30) {real, imag} */,
  {32'hbf4dd065, 32'hbe640b4e} /* (17, 12, 29) {real, imag} */,
  {32'hbf8ea24e, 32'h3fa8a217} /* (17, 12, 28) {real, imag} */,
  {32'hbfaf3e41, 32'hbfc9a6fb} /* (17, 12, 27) {real, imag} */,
  {32'h3f884501, 32'hbec3928c} /* (17, 12, 26) {real, imag} */,
  {32'hbf9e9125, 32'hbe007c84} /* (17, 12, 25) {real, imag} */,
  {32'hbfa26b4c, 32'hbdb71eac} /* (17, 12, 24) {real, imag} */,
  {32'hbaa6ac0e, 32'hbfdd4bca} /* (17, 12, 23) {real, imag} */,
  {32'h3f82d34e, 32'hbfbdf315} /* (17, 12, 22) {real, imag} */,
  {32'h404004c6, 32'hbf77338f} /* (17, 12, 21) {real, imag} */,
  {32'hc09b70af, 32'h3fc4ea60} /* (17, 12, 20) {real, imag} */,
  {32'h3fbba89b, 32'hbf96882b} /* (17, 12, 19) {real, imag} */,
  {32'h401367d6, 32'hc0148b21} /* (17, 12, 18) {real, imag} */,
  {32'h3f678ff0, 32'hbf11f83a} /* (17, 12, 17) {real, imag} */,
  {32'h3fd2c2d2, 32'h3f8fd482} /* (17, 12, 16) {real, imag} */,
  {32'h3f6d29ab, 32'h4020eaf2} /* (17, 12, 15) {real, imag} */,
  {32'h401b688c, 32'h3f67637e} /* (17, 12, 14) {real, imag} */,
  {32'hbee3e42a, 32'h3fee35c6} /* (17, 12, 13) {real, imag} */,
  {32'h3f25cec0, 32'hc02c9f0f} /* (17, 12, 12) {real, imag} */,
  {32'h3ef3b137, 32'h3decc12b} /* (17, 12, 11) {real, imag} */,
  {32'h3fc1df46, 32'hbf5ce81d} /* (17, 12, 10) {real, imag} */,
  {32'h3f524c85, 32'hc021691c} /* (17, 12, 9) {real, imag} */,
  {32'h4039aa56, 32'hc012e219} /* (17, 12, 8) {real, imag} */,
  {32'hbf4d9027, 32'h3feeb509} /* (17, 12, 7) {real, imag} */,
  {32'hbe41c5be, 32'h3f2b4940} /* (17, 12, 6) {real, imag} */,
  {32'hbeb924f8, 32'hbf7d5afe} /* (17, 12, 5) {real, imag} */,
  {32'h3f872a91, 32'h3fdd36c0} /* (17, 12, 4) {real, imag} */,
  {32'h3f244917, 32'h3ef6b977} /* (17, 12, 3) {real, imag} */,
  {32'h3fe4087d, 32'h3f62c8d7} /* (17, 12, 2) {real, imag} */,
  {32'hbf99ed61, 32'hbf98864c} /* (17, 12, 1) {real, imag} */,
  {32'h3f110e34, 32'hbf5674d4} /* (17, 12, 0) {real, imag} */,
  {32'h3ec2ff01, 32'h3f55f42a} /* (17, 11, 31) {real, imag} */,
  {32'h3f902a0e, 32'h4066eedf} /* (17, 11, 30) {real, imag} */,
  {32'h3ec8204f, 32'h3ecde30e} /* (17, 11, 29) {real, imag} */,
  {32'h3f0fa4df, 32'hbf7f3b90} /* (17, 11, 28) {real, imag} */,
  {32'hbf00384f, 32'h3ff7324f} /* (17, 11, 27) {real, imag} */,
  {32'hc000352a, 32'h3f742695} /* (17, 11, 26) {real, imag} */,
  {32'hbf760699, 32'hbf86e425} /* (17, 11, 25) {real, imag} */,
  {32'hbe6d41ac, 32'h3f8f7d28} /* (17, 11, 24) {real, imag} */,
  {32'hbfaab9b3, 32'hc0255688} /* (17, 11, 23) {real, imag} */,
  {32'h3feee609, 32'hbeb97fa9} /* (17, 11, 22) {real, imag} */,
  {32'hbf5e095b, 32'h40021d7a} /* (17, 11, 21) {real, imag} */,
  {32'h4024bbe0, 32'hbf196451} /* (17, 11, 20) {real, imag} */,
  {32'hc02b4862, 32'hbf9c97b6} /* (17, 11, 19) {real, imag} */,
  {32'hbe960288, 32'hbeb04bb0} /* (17, 11, 18) {real, imag} */,
  {32'hbfca2ee8, 32'h3efaaec1} /* (17, 11, 17) {real, imag} */,
  {32'hbfadd9a6, 32'h3f996283} /* (17, 11, 16) {real, imag} */,
  {32'h3fcf0d3f, 32'h3fdb3d56} /* (17, 11, 15) {real, imag} */,
  {32'h40005e6c, 32'h4001989c} /* (17, 11, 14) {real, imag} */,
  {32'h3fa662f2, 32'hbda87792} /* (17, 11, 13) {real, imag} */,
  {32'hbe344454, 32'h40464e1c} /* (17, 11, 12) {real, imag} */,
  {32'hc00d74e8, 32'hbf95a725} /* (17, 11, 11) {real, imag} */,
  {32'hbd9d73f1, 32'hbf772093} /* (17, 11, 10) {real, imag} */,
  {32'h3d626fb6, 32'h3f516278} /* (17, 11, 9) {real, imag} */,
  {32'hbee3458c, 32'hbf291b76} /* (17, 11, 8) {real, imag} */,
  {32'hbfbe7fb4, 32'hc018b55c} /* (17, 11, 7) {real, imag} */,
  {32'hbf82b41c, 32'hbf88a972} /* (17, 11, 6) {real, imag} */,
  {32'h3ffb5aa0, 32'h402f3a40} /* (17, 11, 5) {real, imag} */,
  {32'h3faf4d94, 32'hc01d0233} /* (17, 11, 4) {real, imag} */,
  {32'hbf6cc9ab, 32'h3f20759c} /* (17, 11, 3) {real, imag} */,
  {32'hbcaefe83, 32'hbfbf5582} /* (17, 11, 2) {real, imag} */,
  {32'hbff053de, 32'h3dbb6b1d} /* (17, 11, 1) {real, imag} */,
  {32'h3eda960c, 32'hbf873f38} /* (17, 11, 0) {real, imag} */,
  {32'h3e52efe2, 32'h3f9f103d} /* (17, 10, 31) {real, imag} */,
  {32'h3ec884a5, 32'hbfdb3285} /* (17, 10, 30) {real, imag} */,
  {32'h3f2cb1a2, 32'hbe6ed326} /* (17, 10, 29) {real, imag} */,
  {32'h3fd8f8fd, 32'hbf993279} /* (17, 10, 28) {real, imag} */,
  {32'h400e594a, 32'h3fc2a71a} /* (17, 10, 27) {real, imag} */,
  {32'h3d7f8939, 32'hbe9c8c92} /* (17, 10, 26) {real, imag} */,
  {32'h3fa12691, 32'hbf58bc30} /* (17, 10, 25) {real, imag} */,
  {32'hc0047b19, 32'hbf13302a} /* (17, 10, 24) {real, imag} */,
  {32'hbfb06ad3, 32'hc01ca688} /* (17, 10, 23) {real, imag} */,
  {32'h3f667264, 32'h3e9c89c6} /* (17, 10, 22) {real, imag} */,
  {32'h3fe07b5e, 32'h3e694cd0} /* (17, 10, 21) {real, imag} */,
  {32'hc00a06f4, 32'h3edfdaab} /* (17, 10, 20) {real, imag} */,
  {32'hc021b13a, 32'hbf20677a} /* (17, 10, 19) {real, imag} */,
  {32'h402b6fcc, 32'hbfa76968} /* (17, 10, 18) {real, imag} */,
  {32'h4034486e, 32'h3ff2f32e} /* (17, 10, 17) {real, imag} */,
  {32'h3fb67368, 32'h3efe9fe5} /* (17, 10, 16) {real, imag} */,
  {32'hbfbfb75f, 32'hbd7629c3} /* (17, 10, 15) {real, imag} */,
  {32'h3f76240d, 32'h3f7f2a24} /* (17, 10, 14) {real, imag} */,
  {32'h40284891, 32'h3f3b3618} /* (17, 10, 13) {real, imag} */,
  {32'hbfa12f6c, 32'hc023eabd} /* (17, 10, 12) {real, imag} */,
  {32'hbfd4f4f2, 32'h3e2441d1} /* (17, 10, 11) {real, imag} */,
  {32'h3fe99186, 32'hc0310435} /* (17, 10, 10) {real, imag} */,
  {32'hbef600f6, 32'hbfe52368} /* (17, 10, 9) {real, imag} */,
  {32'hbeea3e6a, 32'h3f8348de} /* (17, 10, 8) {real, imag} */,
  {32'hbf512ff4, 32'h4007ea7c} /* (17, 10, 7) {real, imag} */,
  {32'h3f0a0bcf, 32'hbfaec373} /* (17, 10, 6) {real, imag} */,
  {32'hbf88b499, 32'hbf84538c} /* (17, 10, 5) {real, imag} */,
  {32'h3f79c698, 32'h40411eb5} /* (17, 10, 4) {real, imag} */,
  {32'h3e9ca8c3, 32'h3ef02eba} /* (17, 10, 3) {real, imag} */,
  {32'hbfa12fd6, 32'hbf31e0db} /* (17, 10, 2) {real, imag} */,
  {32'hc0a168a4, 32'h3f883929} /* (17, 10, 1) {real, imag} */,
  {32'h3ec39a73, 32'h3f9c7423} /* (17, 10, 0) {real, imag} */,
  {32'hbdc0a9d3, 32'hbf18a91e} /* (17, 9, 31) {real, imag} */,
  {32'h3e8c05b3, 32'hbf97ac95} /* (17, 9, 30) {real, imag} */,
  {32'hbfd8bf5d, 32'h4011b535} /* (17, 9, 29) {real, imag} */,
  {32'hbfad7319, 32'hbf2fdcdf} /* (17, 9, 28) {real, imag} */,
  {32'h3e8e58ea, 32'hbf5c1b05} /* (17, 9, 27) {real, imag} */,
  {32'hbf3caa6b, 32'h3f03922b} /* (17, 9, 26) {real, imag} */,
  {32'h3fd3698b, 32'h3e330166} /* (17, 9, 25) {real, imag} */,
  {32'h3f9a637e, 32'h40946110} /* (17, 9, 24) {real, imag} */,
  {32'h400eb05f, 32'hc00c3925} /* (17, 9, 23) {real, imag} */,
  {32'hbf91a43b, 32'h3f9fb80c} /* (17, 9, 22) {real, imag} */,
  {32'h40074aa1, 32'hbdd49621} /* (17, 9, 21) {real, imag} */,
  {32'hbe695686, 32'hbfcaef65} /* (17, 9, 20) {real, imag} */,
  {32'hc003c96d, 32'h404c3427} /* (17, 9, 19) {real, imag} */,
  {32'hbf9d1dca, 32'hc0036d7d} /* (17, 9, 18) {real, imag} */,
  {32'hbf97e7a7, 32'hbe7d59f7} /* (17, 9, 17) {real, imag} */,
  {32'hbf6f2d32, 32'h3f437a3e} /* (17, 9, 16) {real, imag} */,
  {32'h3ec706df, 32'h3f0e53b4} /* (17, 9, 15) {real, imag} */,
  {32'h3e777e6c, 32'h3f748674} /* (17, 9, 14) {real, imag} */,
  {32'hbdb273bf, 32'hbf18759b} /* (17, 9, 13) {real, imag} */,
  {32'h3f0fbfb2, 32'h3fba5c3e} /* (17, 9, 12) {real, imag} */,
  {32'hbea0c14d, 32'hbf423fdc} /* (17, 9, 11) {real, imag} */,
  {32'hbfffc5f9, 32'hbfcf3ab8} /* (17, 9, 10) {real, imag} */,
  {32'h3e09f72b, 32'h3f99d682} /* (17, 9, 9) {real, imag} */,
  {32'h3e2bb564, 32'h3dbbd58a} /* (17, 9, 8) {real, imag} */,
  {32'hbefbac38, 32'hbf4394c8} /* (17, 9, 7) {real, imag} */,
  {32'h3ef9e79a, 32'h3f164b81} /* (17, 9, 6) {real, imag} */,
  {32'h3f820ddc, 32'hbf80daea} /* (17, 9, 5) {real, imag} */,
  {32'hc01460d2, 32'h3fbd8dae} /* (17, 9, 4) {real, imag} */,
  {32'hbf954576, 32'hbffea266} /* (17, 9, 3) {real, imag} */,
  {32'h400cdf2e, 32'hbf1399e3} /* (17, 9, 2) {real, imag} */,
  {32'hbfac91e6, 32'hbe64c335} /* (17, 9, 1) {real, imag} */,
  {32'hbd975491, 32'h401e988c} /* (17, 9, 0) {real, imag} */,
  {32'hbf04591d, 32'hbf2f1940} /* (17, 8, 31) {real, imag} */,
  {32'hbf0de9c1, 32'h3fd67364} /* (17, 8, 30) {real, imag} */,
  {32'h3e3545c2, 32'hbea6c3cf} /* (17, 8, 29) {real, imag} */,
  {32'hbf993d34, 32'h40305e31} /* (17, 8, 28) {real, imag} */,
  {32'hbd466ade, 32'hbffc5edc} /* (17, 8, 27) {real, imag} */,
  {32'h3f106920, 32'h3e5e117a} /* (17, 8, 26) {real, imag} */,
  {32'hbefdaca4, 32'h3d6657a1} /* (17, 8, 25) {real, imag} */,
  {32'h3ff32954, 32'h3dd79bc1} /* (17, 8, 24) {real, imag} */,
  {32'h3e8c9591, 32'h3fd6c6ca} /* (17, 8, 23) {real, imag} */,
  {32'hbe04462f, 32'hbfadf115} /* (17, 8, 22) {real, imag} */,
  {32'h3fd13bf4, 32'hc0187536} /* (17, 8, 21) {real, imag} */,
  {32'h3fb0f01d, 32'hbf83f527} /* (17, 8, 20) {real, imag} */,
  {32'h3fcb47d4, 32'h3ff0d25a} /* (17, 8, 19) {real, imag} */,
  {32'hbfcb798f, 32'h3ff347e3} /* (17, 8, 18) {real, imag} */,
  {32'hbd5881bc, 32'hc031ebc0} /* (17, 8, 17) {real, imag} */,
  {32'h3f73193c, 32'hc00b9326} /* (17, 8, 16) {real, imag} */,
  {32'h3eb31995, 32'hbeec46be} /* (17, 8, 15) {real, imag} */,
  {32'h3eff5ae2, 32'h3f839c58} /* (17, 8, 14) {real, imag} */,
  {32'hbe81eeea, 32'hbf48b28f} /* (17, 8, 13) {real, imag} */,
  {32'h3faf4c4a, 32'hbf3559b7} /* (17, 8, 12) {real, imag} */,
  {32'hbf4101d5, 32'hbf481eac} /* (17, 8, 11) {real, imag} */,
  {32'h3e6f889f, 32'hbf2a291f} /* (17, 8, 10) {real, imag} */,
  {32'hbf46f498, 32'h3f1193a1} /* (17, 8, 9) {real, imag} */,
  {32'hbeb5b6a7, 32'h3e9532b8} /* (17, 8, 8) {real, imag} */,
  {32'h3f44a863, 32'hbff383c2} /* (17, 8, 7) {real, imag} */,
  {32'hbda1db43, 32'h3f9cb0d9} /* (17, 8, 6) {real, imag} */,
  {32'hbfc32585, 32'hbfdd94dc} /* (17, 8, 5) {real, imag} */,
  {32'h3f9b990c, 32'h3f6c6c7e} /* (17, 8, 4) {real, imag} */,
  {32'h3f997bba, 32'h3f596ac0} /* (17, 8, 3) {real, imag} */,
  {32'h3dacbfa6, 32'hbf8852b9} /* (17, 8, 2) {real, imag} */,
  {32'hbf81e573, 32'h3feb7810} /* (17, 8, 1) {real, imag} */,
  {32'h39ae2682, 32'h3f291de5} /* (17, 8, 0) {real, imag} */,
  {32'hbfc3204f, 32'h3fa4f957} /* (17, 7, 31) {real, imag} */,
  {32'h3ea1e604, 32'h3f596184} /* (17, 7, 30) {real, imag} */,
  {32'h3ee2f05e, 32'h3f85d651} /* (17, 7, 29) {real, imag} */,
  {32'h3fb4a9f4, 32'h3bdf28dc} /* (17, 7, 28) {real, imag} */,
  {32'hbef94953, 32'hbe6d6bef} /* (17, 7, 27) {real, imag} */,
  {32'hbfc190f6, 32'h3ee2f3ac} /* (17, 7, 26) {real, imag} */,
  {32'hbfaa790d, 32'h3eba1656} /* (17, 7, 25) {real, imag} */,
  {32'hbe94ef6f, 32'hbf89b8a1} /* (17, 7, 24) {real, imag} */,
  {32'hbff43708, 32'h3ec7e39f} /* (17, 7, 23) {real, imag} */,
  {32'h3e8c45a9, 32'h3f22ced2} /* (17, 7, 22) {real, imag} */,
  {32'h3f36442e, 32'hc0410c2c} /* (17, 7, 21) {real, imag} */,
  {32'hbeed439e, 32'h3fc737d0} /* (17, 7, 20) {real, imag} */,
  {32'h3ed68818, 32'h3d21fe99} /* (17, 7, 19) {real, imag} */,
  {32'hc02ceffe, 32'hbfd6cee4} /* (17, 7, 18) {real, imag} */,
  {32'hbf2f476d, 32'h3f2dbada} /* (17, 7, 17) {real, imag} */,
  {32'hbfbc8c91, 32'hc0244974} /* (17, 7, 16) {real, imag} */,
  {32'hbff48f99, 32'hbfc718d5} /* (17, 7, 15) {real, imag} */,
  {32'hbf8bfd5b, 32'hbfadebbc} /* (17, 7, 14) {real, imag} */,
  {32'h40227c45, 32'h3c258bbe} /* (17, 7, 13) {real, imag} */,
  {32'hbe8ea5ec, 32'h3fcd73c1} /* (17, 7, 12) {real, imag} */,
  {32'hbfe489dc, 32'hbfd63edf} /* (17, 7, 11) {real, imag} */,
  {32'hc013e3a1, 32'h3dc56fd8} /* (17, 7, 10) {real, imag} */,
  {32'hbf705542, 32'h402c0172} /* (17, 7, 9) {real, imag} */,
  {32'h3f92c3f0, 32'hbf4926af} /* (17, 7, 8) {real, imag} */,
  {32'h400bc770, 32'h3fb35f9d} /* (17, 7, 7) {real, imag} */,
  {32'hbf860526, 32'hbf125c02} /* (17, 7, 6) {real, imag} */,
  {32'h3e88b9d8, 32'h3f18070f} /* (17, 7, 5) {real, imag} */,
  {32'hbee82a0d, 32'hbf9b3534} /* (17, 7, 4) {real, imag} */,
  {32'h3fd6b64d, 32'hbe67b80a} /* (17, 7, 3) {real, imag} */,
  {32'h3ec6a77b, 32'hbfd2f873} /* (17, 7, 2) {real, imag} */,
  {32'h3ecdbee3, 32'h3ecc4608} /* (17, 7, 1) {real, imag} */,
  {32'hc01f6bd4, 32'hbf3b728c} /* (17, 7, 0) {real, imag} */,
  {32'hc04f342d, 32'hbd7ba6c1} /* (17, 6, 31) {real, imag} */,
  {32'h3e826e00, 32'hbf6fe16a} /* (17, 6, 30) {real, imag} */,
  {32'h3fb09952, 32'hbeab757c} /* (17, 6, 29) {real, imag} */,
  {32'h3f450f1e, 32'h3e6ad09b} /* (17, 6, 28) {real, imag} */,
  {32'h3f8e6fa3, 32'h3f0cd824} /* (17, 6, 27) {real, imag} */,
  {32'hbf873945, 32'h3e147957} /* (17, 6, 26) {real, imag} */,
  {32'h3edf6d60, 32'hbf082cea} /* (17, 6, 25) {real, imag} */,
  {32'h3fa01f49, 32'h40180b19} /* (17, 6, 24) {real, imag} */,
  {32'h3e9f063c, 32'hbf8781e3} /* (17, 6, 23) {real, imag} */,
  {32'hbfc5deff, 32'h3fcb8d0d} /* (17, 6, 22) {real, imag} */,
  {32'hbc1abed5, 32'h3e65ad6d} /* (17, 6, 21) {real, imag} */,
  {32'hc02c86ba, 32'h40297de4} /* (17, 6, 20) {real, imag} */,
  {32'hc01fcdea, 32'h3dd8c48e} /* (17, 6, 19) {real, imag} */,
  {32'hbf6f4963, 32'hbe6eeda9} /* (17, 6, 18) {real, imag} */,
  {32'h3f457d4a, 32'h3e9b7e1e} /* (17, 6, 17) {real, imag} */,
  {32'h3f299518, 32'hbf5c7930} /* (17, 6, 16) {real, imag} */,
  {32'hbeb775fe, 32'h3f85b5d2} /* (17, 6, 15) {real, imag} */,
  {32'hc0071b0d, 32'hc00cab05} /* (17, 6, 14) {real, imag} */,
  {32'h3e4c4615, 32'h3e51202d} /* (17, 6, 13) {real, imag} */,
  {32'hbfdffc9c, 32'hbfa23b60} /* (17, 6, 12) {real, imag} */,
  {32'h3f860ee8, 32'h400b44fa} /* (17, 6, 11) {real, imag} */,
  {32'hbedeca67, 32'hbdbb6b38} /* (17, 6, 10) {real, imag} */,
  {32'h3ffee693, 32'h3f2e1f8d} /* (17, 6, 9) {real, imag} */,
  {32'h3dfeaaf4, 32'h3f9ed0fd} /* (17, 6, 8) {real, imag} */,
  {32'hbf89ad43, 32'h3feb85ae} /* (17, 6, 7) {real, imag} */,
  {32'h3f2c3123, 32'h3e85da05} /* (17, 6, 6) {real, imag} */,
  {32'hbef49c49, 32'hbe358ec6} /* (17, 6, 5) {real, imag} */,
  {32'hc0064ee7, 32'hbef2384d} /* (17, 6, 4) {real, imag} */,
  {32'h3f63f237, 32'h3e41dab4} /* (17, 6, 3) {real, imag} */,
  {32'hbfb3c8c8, 32'h3fd20771} /* (17, 6, 2) {real, imag} */,
  {32'h3a9314cd, 32'hbf0fb2aa} /* (17, 6, 1) {real, imag} */,
  {32'hbffb3fbf, 32'h3fda8879} /* (17, 6, 0) {real, imag} */,
  {32'hbdb27c76, 32'h3e9dbe6f} /* (17, 5, 31) {real, imag} */,
  {32'h3fa1ad12, 32'hbf8f1a01} /* (17, 5, 30) {real, imag} */,
  {32'h3f0c7ed5, 32'h3f2eeb31} /* (17, 5, 29) {real, imag} */,
  {32'h3ea972c8, 32'hbfa26716} /* (17, 5, 28) {real, imag} */,
  {32'hbfaf863a, 32'hbd924427} /* (17, 5, 27) {real, imag} */,
  {32'h3e1e3969, 32'h3fd1784c} /* (17, 5, 26) {real, imag} */,
  {32'hbe039fdb, 32'hc00548e2} /* (17, 5, 25) {real, imag} */,
  {32'h3fde42bf, 32'hbf8055f7} /* (17, 5, 24) {real, imag} */,
  {32'h3c92b71e, 32'h3e5f2e0f} /* (17, 5, 23) {real, imag} */,
  {32'h3f8b239e, 32'hbfff5cee} /* (17, 5, 22) {real, imag} */,
  {32'hbf3d4e88, 32'hbe6e40f5} /* (17, 5, 21) {real, imag} */,
  {32'hbf7b4933, 32'h3ea1590d} /* (17, 5, 20) {real, imag} */,
  {32'h3e7f7b2c, 32'h3ef7a03a} /* (17, 5, 19) {real, imag} */,
  {32'h3e08f03b, 32'hbe2e9747} /* (17, 5, 18) {real, imag} */,
  {32'h3e6bf582, 32'hbf4df6ea} /* (17, 5, 17) {real, imag} */,
  {32'h3fe0b149, 32'hbf71bfa3} /* (17, 5, 16) {real, imag} */,
  {32'h3fea689f, 32'hbf5dc04a} /* (17, 5, 15) {real, imag} */,
  {32'h3fd13e74, 32'hbf71684f} /* (17, 5, 14) {real, imag} */,
  {32'hbf0c3b70, 32'h3e00a1da} /* (17, 5, 13) {real, imag} */,
  {32'hbeaddb9d, 32'hbf140586} /* (17, 5, 12) {real, imag} */,
  {32'hc02bc89c, 32'h403e461a} /* (17, 5, 11) {real, imag} */,
  {32'h3f2d5616, 32'h3fc47db8} /* (17, 5, 10) {real, imag} */,
  {32'h3f4f7dbf, 32'hbd41ad40} /* (17, 5, 9) {real, imag} */,
  {32'hbf3e4940, 32'hbf937181} /* (17, 5, 8) {real, imag} */,
  {32'hbf6a2747, 32'h3f8fd17a} /* (17, 5, 7) {real, imag} */,
  {32'hc00cae83, 32'hc00cb1eb} /* (17, 5, 6) {real, imag} */,
  {32'h3f73de44, 32'hbfcca47c} /* (17, 5, 5) {real, imag} */,
  {32'hbf6b9ae7, 32'h3f163cfd} /* (17, 5, 4) {real, imag} */,
  {32'h3f1d99de, 32'hbff7fcdc} /* (17, 5, 3) {real, imag} */,
  {32'h40177dd4, 32'h4016be88} /* (17, 5, 2) {real, imag} */,
  {32'hbfb50ba0, 32'hc02ad701} /* (17, 5, 1) {real, imag} */,
  {32'h3f562bf3, 32'hbf78089c} /* (17, 5, 0) {real, imag} */,
  {32'h3df99af2, 32'h3e0264d7} /* (17, 4, 31) {real, imag} */,
  {32'hbf9863a5, 32'hbfb1c81a} /* (17, 4, 30) {real, imag} */,
  {32'h4017a694, 32'hbf40edd3} /* (17, 4, 29) {real, imag} */,
  {32'h3e809714, 32'h4004b35c} /* (17, 4, 28) {real, imag} */,
  {32'h3f1a1014, 32'h3f978fde} /* (17, 4, 27) {real, imag} */,
  {32'h3f49c430, 32'hbf58a704} /* (17, 4, 26) {real, imag} */,
  {32'h3f21cc83, 32'h4002087f} /* (17, 4, 25) {real, imag} */,
  {32'h3ed431f0, 32'hbfaf3538} /* (17, 4, 24) {real, imag} */,
  {32'h3f87f9d4, 32'h3d901729} /* (17, 4, 23) {real, imag} */,
  {32'hbfc2aab3, 32'h3f40decf} /* (17, 4, 22) {real, imag} */,
  {32'hbeb64280, 32'h3d8c646c} /* (17, 4, 21) {real, imag} */,
  {32'hbf457c99, 32'hbff9f845} /* (17, 4, 20) {real, imag} */,
  {32'hbe57f9db, 32'hbebf02dd} /* (17, 4, 19) {real, imag} */,
  {32'h3fbae6bc, 32'hbce2f6cd} /* (17, 4, 18) {real, imag} */,
  {32'h3f11e03d, 32'hbf424b24} /* (17, 4, 17) {real, imag} */,
  {32'hbdc30125, 32'hbe97691a} /* (17, 4, 16) {real, imag} */,
  {32'hbe3994e5, 32'h3faf2839} /* (17, 4, 15) {real, imag} */,
  {32'hbf2c4ad9, 32'hbf989797} /* (17, 4, 14) {real, imag} */,
  {32'h3fd42cc0, 32'hbfc785a5} /* (17, 4, 13) {real, imag} */,
  {32'h3fb90d64, 32'h3cdf9e13} /* (17, 4, 12) {real, imag} */,
  {32'h3f57d638, 32'h3fb5d421} /* (17, 4, 11) {real, imag} */,
  {32'h3f420e3b, 32'hbe1ef4f5} /* (17, 4, 10) {real, imag} */,
  {32'h3e375cc2, 32'h3f8e0b2a} /* (17, 4, 9) {real, imag} */,
  {32'hbef5bbfa, 32'hbf920887} /* (17, 4, 8) {real, imag} */,
  {32'hbeb60508, 32'h401c893e} /* (17, 4, 7) {real, imag} */,
  {32'h3efa42ea, 32'hbf4e7310} /* (17, 4, 6) {real, imag} */,
  {32'hc04f1b10, 32'hbdf5d809} /* (17, 4, 5) {real, imag} */,
  {32'hbcce5924, 32'hc0086918} /* (17, 4, 4) {real, imag} */,
  {32'hbfee8894, 32'h3ee65f43} /* (17, 4, 3) {real, imag} */,
  {32'h3fd7d5e3, 32'h3f5c0fe5} /* (17, 4, 2) {real, imag} */,
  {32'hbf887e3a, 32'hbf1c928c} /* (17, 4, 1) {real, imag} */,
  {32'h3f5dfad5, 32'h3f0d5cc3} /* (17, 4, 0) {real, imag} */,
  {32'h3f1370bf, 32'hbe7a4608} /* (17, 3, 31) {real, imag} */,
  {32'hbf593557, 32'hbfa9a733} /* (17, 3, 30) {real, imag} */,
  {32'hbeed75e2, 32'hbfcc05f0} /* (17, 3, 29) {real, imag} */,
  {32'hbf3d970a, 32'hbfa28870} /* (17, 3, 28) {real, imag} */,
  {32'hbecf3196, 32'h3f237ec6} /* (17, 3, 27) {real, imag} */,
  {32'h3f2fd084, 32'h3d944532} /* (17, 3, 26) {real, imag} */,
  {32'hbf2e4787, 32'hbf5b0ad4} /* (17, 3, 25) {real, imag} */,
  {32'h3f204924, 32'h3ed41e99} /* (17, 3, 24) {real, imag} */,
  {32'hbff07a28, 32'hbf8ff85a} /* (17, 3, 23) {real, imag} */,
  {32'hbffd21d8, 32'h3efb86be} /* (17, 3, 22) {real, imag} */,
  {32'h3fd2967c, 32'h3fec994f} /* (17, 3, 21) {real, imag} */,
  {32'hbf0ac1ef, 32'h3fde78db} /* (17, 3, 20) {real, imag} */,
  {32'h3f6f92a0, 32'hbd452245} /* (17, 3, 19) {real, imag} */,
  {32'hbfcc04ae, 32'h3fad75af} /* (17, 3, 18) {real, imag} */,
  {32'h3f8905be, 32'h3eb010ba} /* (17, 3, 17) {real, imag} */,
  {32'h3fc49285, 32'hbec4a2d9} /* (17, 3, 16) {real, imag} */,
  {32'hbdbc5097, 32'hbf705e46} /* (17, 3, 15) {real, imag} */,
  {32'hbfebc910, 32'h3f6bff82} /* (17, 3, 14) {real, imag} */,
  {32'h3fbf2923, 32'hbe900cd9} /* (17, 3, 13) {real, imag} */,
  {32'hbe4c385f, 32'hc01217a0} /* (17, 3, 12) {real, imag} */,
  {32'h3fd73834, 32'hbf233678} /* (17, 3, 11) {real, imag} */,
  {32'hbfa71b8a, 32'h400cd184} /* (17, 3, 10) {real, imag} */,
  {32'hbf918a82, 32'hbf56443c} /* (17, 3, 9) {real, imag} */,
  {32'h401ffe57, 32'hbf459a64} /* (17, 3, 8) {real, imag} */,
  {32'hbf7200f5, 32'h3fc353d9} /* (17, 3, 7) {real, imag} */,
  {32'hbf466943, 32'h3fc6b178} /* (17, 3, 6) {real, imag} */,
  {32'h3fb9722c, 32'hbea04591} /* (17, 3, 5) {real, imag} */,
  {32'hbf88b849, 32'hbd4ead9c} /* (17, 3, 4) {real, imag} */,
  {32'hbdb214fb, 32'h3fa5bbca} /* (17, 3, 3) {real, imag} */,
  {32'hbe160cd1, 32'hbf8e1901} /* (17, 3, 2) {real, imag} */,
  {32'h3f01f624, 32'h3fb85fa7} /* (17, 3, 1) {real, imag} */,
  {32'h3ff86cdd, 32'h3f291748} /* (17, 3, 0) {real, imag} */,
  {32'h3d008666, 32'hbfe280bc} /* (17, 2, 31) {real, imag} */,
  {32'h3f41915a, 32'hbd0d90fb} /* (17, 2, 30) {real, imag} */,
  {32'h3fa5294a, 32'h3f98404c} /* (17, 2, 29) {real, imag} */,
  {32'hbf06f112, 32'h3f18bc6b} /* (17, 2, 28) {real, imag} */,
  {32'hbfac4a4e, 32'hbe1c67c8} /* (17, 2, 27) {real, imag} */,
  {32'hbe47db9d, 32'h3f4792f0} /* (17, 2, 26) {real, imag} */,
  {32'hbf497764, 32'hbdc10890} /* (17, 2, 25) {real, imag} */,
  {32'h3fe3b23a, 32'h3f4fe9fb} /* (17, 2, 24) {real, imag} */,
  {32'h3d014839, 32'h403774a2} /* (17, 2, 23) {real, imag} */,
  {32'hbe6a38f4, 32'h3fe9786b} /* (17, 2, 22) {real, imag} */,
  {32'hc03262a3, 32'hbeca34f2} /* (17, 2, 21) {real, imag} */,
  {32'h3f37a9cc, 32'hbd96ca50} /* (17, 2, 20) {real, imag} */,
  {32'h3d98e0fb, 32'hbf3a8ce5} /* (17, 2, 19) {real, imag} */,
  {32'h3d17cee8, 32'h3f414db0} /* (17, 2, 18) {real, imag} */,
  {32'hbf41319e, 32'hbfcfa97d} /* (17, 2, 17) {real, imag} */,
  {32'h3f9ec299, 32'h3f54f496} /* (17, 2, 16) {real, imag} */,
  {32'h3f80e86e, 32'h3f664da0} /* (17, 2, 15) {real, imag} */,
  {32'hbfca0610, 32'hbfa8a7d7} /* (17, 2, 14) {real, imag} */,
  {32'hbf07238d, 32'h3e66084d} /* (17, 2, 13) {real, imag} */,
  {32'h3f362f52, 32'hbf35a23b} /* (17, 2, 12) {real, imag} */,
  {32'h3f57609d, 32'h3f7389f9} /* (17, 2, 11) {real, imag} */,
  {32'h3fb18439, 32'hbf1c9b37} /* (17, 2, 10) {real, imag} */,
  {32'hbf2ab9e5, 32'hbfb36e2b} /* (17, 2, 9) {real, imag} */,
  {32'h3faaba90, 32'h3e75a233} /* (17, 2, 8) {real, imag} */,
  {32'hbfa83419, 32'hbf38f3f2} /* (17, 2, 7) {real, imag} */,
  {32'h3f078ceb, 32'h3f4321e0} /* (17, 2, 6) {real, imag} */,
  {32'hbfb55a5b, 32'h3f040791} /* (17, 2, 5) {real, imag} */,
  {32'h3eeeb3be, 32'h3f9b3c8f} /* (17, 2, 4) {real, imag} */,
  {32'hbf53af39, 32'h3f33baf4} /* (17, 2, 3) {real, imag} */,
  {32'h402f9dc4, 32'h3fc8d9aa} /* (17, 2, 2) {real, imag} */,
  {32'h3d8be3a9, 32'hbf8dfaa4} /* (17, 2, 1) {real, imag} */,
  {32'hbe96e111, 32'hbf8b6b41} /* (17, 2, 0) {real, imag} */,
  {32'h400e6349, 32'hbfd5ef51} /* (17, 1, 31) {real, imag} */,
  {32'hbed99beb, 32'h400e31dd} /* (17, 1, 30) {real, imag} */,
  {32'h3c82cef3, 32'hbf56007c} /* (17, 1, 29) {real, imag} */,
  {32'h3d36aaff, 32'hbfa0dd99} /* (17, 1, 28) {real, imag} */,
  {32'h3f903d07, 32'h3fdd53cb} /* (17, 1, 27) {real, imag} */,
  {32'hbf00bcab, 32'hc014775c} /* (17, 1, 26) {real, imag} */,
  {32'h4018d82f, 32'hbff9250a} /* (17, 1, 25) {real, imag} */,
  {32'hbe417e70, 32'h400d11be} /* (17, 1, 24) {real, imag} */,
  {32'h3f84c5ff, 32'h400aed9e} /* (17, 1, 23) {real, imag} */,
  {32'h3e00cf5d, 32'hbe4ac89a} /* (17, 1, 22) {real, imag} */,
  {32'h3fb238be, 32'h3ec56bc5} /* (17, 1, 21) {real, imag} */,
  {32'h40580e32, 32'hbe3730f8} /* (17, 1, 20) {real, imag} */,
  {32'h3e8035e9, 32'hbe3163cc} /* (17, 1, 19) {real, imag} */,
  {32'hbf2b7ec9, 32'h3e409ea2} /* (17, 1, 18) {real, imag} */,
  {32'h3fe00f12, 32'hbfeaac91} /* (17, 1, 17) {real, imag} */,
  {32'h3cdf7016, 32'hbd014a39} /* (17, 1, 16) {real, imag} */,
  {32'hbf4d1485, 32'hbf9f1b26} /* (17, 1, 15) {real, imag} */,
  {32'hbf8f4a50, 32'h3f43e234} /* (17, 1, 14) {real, imag} */,
  {32'hbedaebba, 32'hbfbc585f} /* (17, 1, 13) {real, imag} */,
  {32'h3f666742, 32'h3f72c5a6} /* (17, 1, 12) {real, imag} */,
  {32'hbe542699, 32'h3fc0363a} /* (17, 1, 11) {real, imag} */,
  {32'h3f89260e, 32'hbfef1c15} /* (17, 1, 10) {real, imag} */,
  {32'hbf52c46a, 32'hbfcfced6} /* (17, 1, 9) {real, imag} */,
  {32'hbf86353b, 32'h3ea1bd36} /* (17, 1, 8) {real, imag} */,
  {32'h3f741f78, 32'h3f2199f2} /* (17, 1, 7) {real, imag} */,
  {32'hbe388719, 32'hbfcae9d8} /* (17, 1, 6) {real, imag} */,
  {32'hc037eb6a, 32'hbfd4ba44} /* (17, 1, 5) {real, imag} */,
  {32'h3f3d8caa, 32'hbf731b47} /* (17, 1, 4) {real, imag} */,
  {32'hbf958e79, 32'hc072430c} /* (17, 1, 3) {real, imag} */,
  {32'hbffb9a3d, 32'hbf68dc30} /* (17, 1, 2) {real, imag} */,
  {32'h3f8ddb01, 32'h3f76c711} /* (17, 1, 1) {real, imag} */,
  {32'h3d06068c, 32'h3f5f05f7} /* (17, 1, 0) {real, imag} */,
  {32'hbf754673, 32'h3ec821b1} /* (17, 0, 31) {real, imag} */,
  {32'h3c381615, 32'h3a300204} /* (17, 0, 30) {real, imag} */,
  {32'hbfc45292, 32'h3ffcfd67} /* (17, 0, 29) {real, imag} */,
  {32'hbfdb7095, 32'h3eb22468} /* (17, 0, 28) {real, imag} */,
  {32'hbe4c6b6a, 32'h3e69d500} /* (17, 0, 27) {real, imag} */,
  {32'h3f4d3e85, 32'hbeea1d6e} /* (17, 0, 26) {real, imag} */,
  {32'h3f4446cd, 32'h401571dc} /* (17, 0, 25) {real, imag} */,
  {32'h404d5e9c, 32'h3f926da6} /* (17, 0, 24) {real, imag} */,
  {32'h3d8c6d3a, 32'hc00e82f2} /* (17, 0, 23) {real, imag} */,
  {32'hbf26770d, 32'hbf5abacc} /* (17, 0, 22) {real, imag} */,
  {32'hbf81315e, 32'hbfe361d2} /* (17, 0, 21) {real, imag} */,
  {32'h3f4ba22a, 32'hbe6641f6} /* (17, 0, 20) {real, imag} */,
  {32'h4007e254, 32'hbf26f718} /* (17, 0, 19) {real, imag} */,
  {32'hbfb6ad6a, 32'h3f4785bf} /* (17, 0, 18) {real, imag} */,
  {32'hbd497a38, 32'h3f816bef} /* (17, 0, 17) {real, imag} */,
  {32'h3f19bb43, 32'hbead3075} /* (17, 0, 16) {real, imag} */,
  {32'h3f0ea30c, 32'hbf8a7803} /* (17, 0, 15) {real, imag} */,
  {32'h4049f3cf, 32'h3f010efb} /* (17, 0, 14) {real, imag} */,
  {32'hbfc42213, 32'hc006f0d2} /* (17, 0, 13) {real, imag} */,
  {32'h3e90eed7, 32'h3f44e3d5} /* (17, 0, 12) {real, imag} */,
  {32'hbf3a5626, 32'hbee5e02a} /* (17, 0, 11) {real, imag} */,
  {32'h3f95d059, 32'h3f496e6d} /* (17, 0, 10) {real, imag} */,
  {32'h3f50deda, 32'hbf473f58} /* (17, 0, 9) {real, imag} */,
  {32'hbfaeed9f, 32'h3c19556c} /* (17, 0, 8) {real, imag} */,
  {32'h3f1c58c2, 32'hbe1c26f3} /* (17, 0, 7) {real, imag} */,
  {32'hbf05f859, 32'h3f8625f1} /* (17, 0, 6) {real, imag} */,
  {32'hbf370a9f, 32'hbf72b8d9} /* (17, 0, 5) {real, imag} */,
  {32'hbfe514ad, 32'h3f81f94e} /* (17, 0, 4) {real, imag} */,
  {32'hbec0ba3a, 32'h3ff1d194} /* (17, 0, 3) {real, imag} */,
  {32'h3efb4f57, 32'hbf9ddb2c} /* (17, 0, 2) {real, imag} */,
  {32'h3dc8437d, 32'h4010d8a0} /* (17, 0, 1) {real, imag} */,
  {32'h3f32920e, 32'hbf71358b} /* (17, 0, 0) {real, imag} */,
  {32'hbe4f5ee5, 32'h3afde438} /* (16, 31, 31) {real, imag} */,
  {32'hbf525e6a, 32'hbfa5852b} /* (16, 31, 30) {real, imag} */,
  {32'hbedb507a, 32'h3f91ea45} /* (16, 31, 29) {real, imag} */,
  {32'hbfe4a6fe, 32'h3f411c83} /* (16, 31, 28) {real, imag} */,
  {32'h3fad2841, 32'h3ec7d2bb} /* (16, 31, 27) {real, imag} */,
  {32'h3e8a5470, 32'hbedf3643} /* (16, 31, 26) {real, imag} */,
  {32'hbe9f1a5d, 32'h3ec72279} /* (16, 31, 25) {real, imag} */,
  {32'h3dd9cf7f, 32'h3db04dc8} /* (16, 31, 24) {real, imag} */,
  {32'h3f8de299, 32'h3fbcac11} /* (16, 31, 23) {real, imag} */,
  {32'hbfeeb48c, 32'hbf16f076} /* (16, 31, 22) {real, imag} */,
  {32'hbeee653d, 32'h400009f7} /* (16, 31, 21) {real, imag} */,
  {32'h3e51cb50, 32'h3f6e6ff2} /* (16, 31, 20) {real, imag} */,
  {32'h3eef3160, 32'hbfd9192c} /* (16, 31, 19) {real, imag} */,
  {32'hbd4127f2, 32'hbeb2458b} /* (16, 31, 18) {real, imag} */,
  {32'h3d9616b9, 32'hbbe1ba61} /* (16, 31, 17) {real, imag} */,
  {32'h3e00f0fc, 32'hbf9090d9} /* (16, 31, 16) {real, imag} */,
  {32'hbdb92454, 32'h3ce68a89} /* (16, 31, 15) {real, imag} */,
  {32'h3f119517, 32'hbf05c3e8} /* (16, 31, 14) {real, imag} */,
  {32'h3f5416e0, 32'h3f8d26e7} /* (16, 31, 13) {real, imag} */,
  {32'hc0138540, 32'h3de08795} /* (16, 31, 12) {real, imag} */,
  {32'hbf4e0358, 32'hbe66959a} /* (16, 31, 11) {real, imag} */,
  {32'hbf74bebd, 32'hbf20016f} /* (16, 31, 10) {real, imag} */,
  {32'hbf2da598, 32'h3e7eac86} /* (16, 31, 9) {real, imag} */,
  {32'hbe50a3a8, 32'h3f81fd71} /* (16, 31, 8) {real, imag} */,
  {32'hbe0e1c56, 32'h3db79849} /* (16, 31, 7) {real, imag} */,
  {32'h3f15915b, 32'hbf75e42e} /* (16, 31, 6) {real, imag} */,
  {32'hbe043dbf, 32'h3fadfb23} /* (16, 31, 5) {real, imag} */,
  {32'h3d9816f6, 32'h3d9f17ba} /* (16, 31, 4) {real, imag} */,
  {32'h3ecf393a, 32'hbfb96afd} /* (16, 31, 3) {real, imag} */,
  {32'hbf1b10cc, 32'hbfbd0080} /* (16, 31, 2) {real, imag} */,
  {32'h3f2a469f, 32'hbf9e0196} /* (16, 31, 1) {real, imag} */,
  {32'h3f805e94, 32'h3ea769a9} /* (16, 31, 0) {real, imag} */,
  {32'hbfc6d9e9, 32'hbf12a3af} /* (16, 30, 31) {real, imag} */,
  {32'hbf04ab9f, 32'hbf30b39f} /* (16, 30, 30) {real, imag} */,
  {32'hbf2b66ba, 32'h3f55954d} /* (16, 30, 29) {real, imag} */,
  {32'hbef0dd36, 32'hbfb30aaf} /* (16, 30, 28) {real, imag} */,
  {32'h3fb6a836, 32'h3e811004} /* (16, 30, 27) {real, imag} */,
  {32'h3ed49852, 32'hbfb9dd2e} /* (16, 30, 26) {real, imag} */,
  {32'hbebaca04, 32'hbd818fc8} /* (16, 30, 25) {real, imag} */,
  {32'hbf5d6854, 32'hbf85e826} /* (16, 30, 24) {real, imag} */,
  {32'hbd0fcb66, 32'hbe742233} /* (16, 30, 23) {real, imag} */,
  {32'h3fedb83e, 32'hbe8b766b} /* (16, 30, 22) {real, imag} */,
  {32'h401243cc, 32'hbf72144c} /* (16, 30, 21) {real, imag} */,
  {32'hbd78f5ac, 32'h3f8756a0} /* (16, 30, 20) {real, imag} */,
  {32'hbf80fd51, 32'h3e6cd2d9} /* (16, 30, 19) {real, imag} */,
  {32'hbef9e34a, 32'h3ef09ccb} /* (16, 30, 18) {real, imag} */,
  {32'hbf7e096c, 32'h3f30cb2a} /* (16, 30, 17) {real, imag} */,
  {32'h3d856b61, 32'h3e5ecb6d} /* (16, 30, 16) {real, imag} */,
  {32'hbe948e26, 32'hbfe0646f} /* (16, 30, 15) {real, imag} */,
  {32'hbd1282cb, 32'h3f120c33} /* (16, 30, 14) {real, imag} */,
  {32'hc01d1d22, 32'hbfee0490} /* (16, 30, 13) {real, imag} */,
  {32'hbe2c862a, 32'hbea53cee} /* (16, 30, 12) {real, imag} */,
  {32'h3f146084, 32'hbe6db50d} /* (16, 30, 11) {real, imag} */,
  {32'hc0362897, 32'hbf40f171} /* (16, 30, 10) {real, imag} */,
  {32'h3fbcb5a0, 32'h3f52fc27} /* (16, 30, 9) {real, imag} */,
  {32'h3ef307f9, 32'hbf974d22} /* (16, 30, 8) {real, imag} */,
  {32'hbb8d60a1, 32'h3f6c511c} /* (16, 30, 7) {real, imag} */,
  {32'h3e9c19ad, 32'hbeefb723} /* (16, 30, 6) {real, imag} */,
  {32'hbf686d9d, 32'h3af5929e} /* (16, 30, 5) {real, imag} */,
  {32'h3f21cbc9, 32'h3eb064ce} /* (16, 30, 4) {real, imag} */,
  {32'hbf26e2f7, 32'h3f34faf3} /* (16, 30, 3) {real, imag} */,
  {32'h3f6a5e85, 32'hbeac98cc} /* (16, 30, 2) {real, imag} */,
  {32'h3d12906e, 32'h3ec6ecb4} /* (16, 30, 1) {real, imag} */,
  {32'h3d8ead56, 32'hbe8dc88d} /* (16, 30, 0) {real, imag} */,
  {32'hbfe5fc66, 32'hbf949405} /* (16, 29, 31) {real, imag} */,
  {32'h3e736e70, 32'h3fbf95e1} /* (16, 29, 30) {real, imag} */,
  {32'hbf8fdbf5, 32'hbe84fe8a} /* (16, 29, 29) {real, imag} */,
  {32'hbe41a8a7, 32'h3f02d235} /* (16, 29, 28) {real, imag} */,
  {32'h3f7ed4e4, 32'hbf0ace45} /* (16, 29, 27) {real, imag} */,
  {32'hbecbf76c, 32'h3f18531a} /* (16, 29, 26) {real, imag} */,
  {32'h3e587921, 32'hbfeab37c} /* (16, 29, 25) {real, imag} */,
  {32'h3f5816a6, 32'h3e585c10} /* (16, 29, 24) {real, imag} */,
  {32'hbf7923c5, 32'h3f85d18f} /* (16, 29, 23) {real, imag} */,
  {32'h3fa47ecf, 32'h3e32ea78} /* (16, 29, 22) {real, imag} */,
  {32'h40090b0d, 32'hc0200d2a} /* (16, 29, 21) {real, imag} */,
  {32'h3ddae87b, 32'h3f528286} /* (16, 29, 20) {real, imag} */,
  {32'hbf0c38e3, 32'h402954ad} /* (16, 29, 19) {real, imag} */,
  {32'h3f358d66, 32'h3fd15669} /* (16, 29, 18) {real, imag} */,
  {32'hbf4a6b10, 32'hbf871365} /* (16, 29, 17) {real, imag} */,
  {32'hbdd8b902, 32'hbeef3335} /* (16, 29, 16) {real, imag} */,
  {32'h3fc56e5b, 32'h3f672ccd} /* (16, 29, 15) {real, imag} */,
  {32'hbfe59f7f, 32'h3e5ac2ff} /* (16, 29, 14) {real, imag} */,
  {32'h3f5140b0, 32'h3ee1fa37} /* (16, 29, 13) {real, imag} */,
  {32'hbf3f0dbc, 32'hbf378b65} /* (16, 29, 12) {real, imag} */,
  {32'hbfa0bb84, 32'hbef4999f} /* (16, 29, 11) {real, imag} */,
  {32'h3f622a09, 32'hbd3c5058} /* (16, 29, 10) {real, imag} */,
  {32'hbe87c95e, 32'h3f2b1257} /* (16, 29, 9) {real, imag} */,
  {32'hbf020d27, 32'h3fb076a9} /* (16, 29, 8) {real, imag} */,
  {32'hbfb8a978, 32'h3f499372} /* (16, 29, 7) {real, imag} */,
  {32'h3f6c2cbc, 32'h3f2ad22b} /* (16, 29, 6) {real, imag} */,
  {32'hbe8f2f86, 32'h3f79be9c} /* (16, 29, 5) {real, imag} */,
  {32'h3fc10dd1, 32'hbf0cb92e} /* (16, 29, 4) {real, imag} */,
  {32'hbfbd2d67, 32'hbffadf08} /* (16, 29, 3) {real, imag} */,
  {32'hbef971f5, 32'h3f1df3d1} /* (16, 29, 2) {real, imag} */,
  {32'hbff2a3d2, 32'hbf92f748} /* (16, 29, 1) {real, imag} */,
  {32'hbeaad7d0, 32'h3d3c728b} /* (16, 29, 0) {real, imag} */,
  {32'h3bf4c2f0, 32'h3f31504d} /* (16, 28, 31) {real, imag} */,
  {32'hbe7d79b0, 32'hc0013560} /* (16, 28, 30) {real, imag} */,
  {32'h3f86a0cb, 32'h3e7e349c} /* (16, 28, 29) {real, imag} */,
  {32'h3f41050e, 32'h400ab187} /* (16, 28, 28) {real, imag} */,
  {32'h3f08d3a3, 32'hbf8bd079} /* (16, 28, 27) {real, imag} */,
  {32'hbfb8e8a7, 32'hbf35d13c} /* (16, 28, 26) {real, imag} */,
  {32'hbf99b0c8, 32'hbf2da2aa} /* (16, 28, 25) {real, imag} */,
  {32'h3f366194, 32'h3f6babfc} /* (16, 28, 24) {real, imag} */,
  {32'h3f561869, 32'hbfa3e169} /* (16, 28, 23) {real, imag} */,
  {32'h3f8b15fd, 32'hc03b67a1} /* (16, 28, 22) {real, imag} */,
  {32'hbf9fd026, 32'h3fdeca42} /* (16, 28, 21) {real, imag} */,
  {32'h3f87a042, 32'h3f6b0687} /* (16, 28, 20) {real, imag} */,
  {32'hbf42041d, 32'hbf9ee31f} /* (16, 28, 19) {real, imag} */,
  {32'h3f9f3443, 32'h3ed74d5d} /* (16, 28, 18) {real, imag} */,
  {32'hbfb36337, 32'h3f655fbe} /* (16, 28, 17) {real, imag} */,
  {32'hbde23ff9, 32'h3f8d1be8} /* (16, 28, 16) {real, imag} */,
  {32'hc0194ae6, 32'hc0223e34} /* (16, 28, 15) {real, imag} */,
  {32'hbfce5079, 32'h3e9cfda4} /* (16, 28, 14) {real, imag} */,
  {32'hbeb046ed, 32'h3f2e77eb} /* (16, 28, 13) {real, imag} */,
  {32'h3eb44a3e, 32'h3fefe21c} /* (16, 28, 12) {real, imag} */,
  {32'h3f146252, 32'hbf2715dc} /* (16, 28, 11) {real, imag} */,
  {32'h3ec52fde, 32'hbf529033} /* (16, 28, 10) {real, imag} */,
  {32'h400131f8, 32'h3e43553a} /* (16, 28, 9) {real, imag} */,
  {32'hbf8b7d9e, 32'hbe8b5ff8} /* (16, 28, 8) {real, imag} */,
  {32'h3fb5c7db, 32'h3f83143f} /* (16, 28, 7) {real, imag} */,
  {32'h3f9c91d7, 32'h3db4fedf} /* (16, 28, 6) {real, imag} */,
  {32'hbedcdd58, 32'hbfc930a0} /* (16, 28, 5) {real, imag} */,
  {32'hbff35c29, 32'hbe8c48fe} /* (16, 28, 4) {real, imag} */,
  {32'hbd24cc3c, 32'hbe9964f9} /* (16, 28, 3) {real, imag} */,
  {32'hbf37eab3, 32'hbf9fc1a7} /* (16, 28, 2) {real, imag} */,
  {32'h3f62657b, 32'h400ccab8} /* (16, 28, 1) {real, imag} */,
  {32'hbf51b94f, 32'h3f2880f1} /* (16, 28, 0) {real, imag} */,
  {32'hbf0f97f1, 32'h3f29b130} /* (16, 27, 31) {real, imag} */,
  {32'hbf9effce, 32'hbe92957a} /* (16, 27, 30) {real, imag} */,
  {32'h3f58591d, 32'hbfb66cfc} /* (16, 27, 29) {real, imag} */,
  {32'hbe8b0c93, 32'h3fb7b6f8} /* (16, 27, 28) {real, imag} */,
  {32'hbe4c8dd4, 32'hbffffa16} /* (16, 27, 27) {real, imag} */,
  {32'hbe002223, 32'hbf1c6d6c} /* (16, 27, 26) {real, imag} */,
  {32'hbede1e2d, 32'hbf0f5d6d} /* (16, 27, 25) {real, imag} */,
  {32'h3fbe34bf, 32'h3eef9a31} /* (16, 27, 24) {real, imag} */,
  {32'hbf496480, 32'hbf721a1d} /* (16, 27, 23) {real, imag} */,
  {32'h3eda3d67, 32'hbca0770b} /* (16, 27, 22) {real, imag} */,
  {32'h3fdb8b36, 32'hbf196083} /* (16, 27, 21) {real, imag} */,
  {32'hbf3b8062, 32'h3ee30373} /* (16, 27, 20) {real, imag} */,
  {32'hbe0a05a2, 32'hbecf484c} /* (16, 27, 19) {real, imag} */,
  {32'h3f3de5ed, 32'hbf213088} /* (16, 27, 18) {real, imag} */,
  {32'h3eb7f0ec, 32'hbfe7952a} /* (16, 27, 17) {real, imag} */,
  {32'h3d83466c, 32'h3f173c09} /* (16, 27, 16) {real, imag} */,
  {32'hbf435afa, 32'hbdb668c5} /* (16, 27, 15) {real, imag} */,
  {32'hbfa13402, 32'h3e6a7978} /* (16, 27, 14) {real, imag} */,
  {32'h3e8dcbb7, 32'h3ffa15c4} /* (16, 27, 13) {real, imag} */,
  {32'hbfed6845, 32'h3e632879} /* (16, 27, 12) {real, imag} */,
  {32'h3f12d504, 32'h3fb83f29} /* (16, 27, 11) {real, imag} */,
  {32'h3f0c7772, 32'hbd3c0f2d} /* (16, 27, 10) {real, imag} */,
  {32'h3d18ffd3, 32'h3f28f975} /* (16, 27, 9) {real, imag} */,
  {32'h3f68d353, 32'hbe8e72b3} /* (16, 27, 8) {real, imag} */,
  {32'hbcb89da4, 32'hbdf2f694} /* (16, 27, 7) {real, imag} */,
  {32'hbf2ce2ec, 32'hbf6939ec} /* (16, 27, 6) {real, imag} */,
  {32'hbf126670, 32'hbf7a3950} /* (16, 27, 5) {real, imag} */,
  {32'h3ee8e4ae, 32'hbf616ff8} /* (16, 27, 4) {real, imag} */,
  {32'h3fb05d62, 32'h3c2fbe81} /* (16, 27, 3) {real, imag} */,
  {32'hbe8b8da7, 32'hbff519b5} /* (16, 27, 2) {real, imag} */,
  {32'hbe996a02, 32'h3f37bd09} /* (16, 27, 1) {real, imag} */,
  {32'hbe6f81a5, 32'h3fa42237} /* (16, 27, 0) {real, imag} */,
  {32'hbfad9650, 32'h4002aa2f} /* (16, 26, 31) {real, imag} */,
  {32'hbf1c9518, 32'h3f169f70} /* (16, 26, 30) {real, imag} */,
  {32'hbdf31a93, 32'hbf91f9aa} /* (16, 26, 29) {real, imag} */,
  {32'h3f7750d5, 32'hbd2a4bbb} /* (16, 26, 28) {real, imag} */,
  {32'h3fd081ff, 32'hbee9ccf7} /* (16, 26, 27) {real, imag} */,
  {32'h3ed10fe4, 32'h3f3be682} /* (16, 26, 26) {real, imag} */,
  {32'hbf397af8, 32'hbf99571c} /* (16, 26, 25) {real, imag} */,
  {32'h3ffcc9e2, 32'h3e0b5949} /* (16, 26, 24) {real, imag} */,
  {32'h3ed21950, 32'h3f9411a9} /* (16, 26, 23) {real, imag} */,
  {32'hbfb329fa, 32'hbdaee7f1} /* (16, 26, 22) {real, imag} */,
  {32'h3fbfab7d, 32'h401f6483} /* (16, 26, 21) {real, imag} */,
  {32'h3f4ef2b8, 32'h3e292d47} /* (16, 26, 20) {real, imag} */,
  {32'hbd1f232b, 32'h3ed8e24a} /* (16, 26, 19) {real, imag} */,
  {32'h3ee56818, 32'hbeb1d60f} /* (16, 26, 18) {real, imag} */,
  {32'h3f9d623a, 32'hbf55309a} /* (16, 26, 17) {real, imag} */,
  {32'hbdb1c068, 32'h3bedd744} /* (16, 26, 16) {real, imag} */,
  {32'hbf0fa3e0, 32'h3fd36074} /* (16, 26, 15) {real, imag} */,
  {32'hbf1f8a48, 32'h3f9a8703} /* (16, 26, 14) {real, imag} */,
  {32'h3fb9193e, 32'h3fb9509b} /* (16, 26, 13) {real, imag} */,
  {32'h3fec7647, 32'hbf74a6a8} /* (16, 26, 12) {real, imag} */,
  {32'h3f57f53f, 32'h3f2a9e50} /* (16, 26, 11) {real, imag} */,
  {32'h3ed844fa, 32'h3fc98ba4} /* (16, 26, 10) {real, imag} */,
  {32'hbf7149d7, 32'h3e1abc02} /* (16, 26, 9) {real, imag} */,
  {32'h3f696e5e, 32'hbe4ff717} /* (16, 26, 8) {real, imag} */,
  {32'hbf9ca9cf, 32'h3fa16415} /* (16, 26, 7) {real, imag} */,
  {32'hbf83dd4e, 32'h3d1a5586} /* (16, 26, 6) {real, imag} */,
  {32'hbf8dbcd9, 32'hbfa456ce} /* (16, 26, 5) {real, imag} */,
  {32'hbfbc623b, 32'hbd21a9f1} /* (16, 26, 4) {real, imag} */,
  {32'hbf22027e, 32'hbfcc7e2f} /* (16, 26, 3) {real, imag} */,
  {32'h3f122d10, 32'hbf84d518} /* (16, 26, 2) {real, imag} */,
  {32'hbf59cb6d, 32'h3ef90db4} /* (16, 26, 1) {real, imag} */,
  {32'h3de8cc59, 32'h3fa96b66} /* (16, 26, 0) {real, imag} */,
  {32'h3f64a5b4, 32'h3ca52d7e} /* (16, 25, 31) {real, imag} */,
  {32'hbf5b38ad, 32'hbda1c9a6} /* (16, 25, 30) {real, imag} */,
  {32'hbe54c55d, 32'hbfc01631} /* (16, 25, 29) {real, imag} */,
  {32'hbfc02ff3, 32'hbf857430} /* (16, 25, 28) {real, imag} */,
  {32'hbf33a5f8, 32'hc00744f6} /* (16, 25, 27) {real, imag} */,
  {32'h3dbdd7d8, 32'hbee367c5} /* (16, 25, 26) {real, imag} */,
  {32'hbff6351c, 32'h3e1c00cb} /* (16, 25, 25) {real, imag} */,
  {32'h3eb54fb1, 32'h3f1e0512} /* (16, 25, 24) {real, imag} */,
  {32'hbe3c101f, 32'h40021f4e} /* (16, 25, 23) {real, imag} */,
  {32'hbee3aeba, 32'h3f116c92} /* (16, 25, 22) {real, imag} */,
  {32'h3ec24501, 32'hbbf18c38} /* (16, 25, 21) {real, imag} */,
  {32'hbded0ce0, 32'hbfd32062} /* (16, 25, 20) {real, imag} */,
  {32'hbf913b57, 32'hbf53d509} /* (16, 25, 19) {real, imag} */,
  {32'h3f582973, 32'hbf87b15c} /* (16, 25, 18) {real, imag} */,
  {32'h3e44ead7, 32'h3f1d336d} /* (16, 25, 17) {real, imag} */,
  {32'hbf519b41, 32'hbf85553d} /* (16, 25, 16) {real, imag} */,
  {32'hbee6c9b2, 32'h3f739b92} /* (16, 25, 15) {real, imag} */,
  {32'h3d91088c, 32'hbe61c08f} /* (16, 25, 14) {real, imag} */,
  {32'hbef78e8e, 32'h3f20c077} /* (16, 25, 13) {real, imag} */,
  {32'hbf828ab0, 32'h3f5bd0e2} /* (16, 25, 12) {real, imag} */,
  {32'h3fa05403, 32'h3e04a6a4} /* (16, 25, 11) {real, imag} */,
  {32'hc00c818c, 32'h3fbb9fed} /* (16, 25, 10) {real, imag} */,
  {32'h3f10fbc7, 32'h3cff5002} /* (16, 25, 9) {real, imag} */,
  {32'hbf0b06e4, 32'hbd3d12ea} /* (16, 25, 8) {real, imag} */,
  {32'hbfacf73b, 32'hbf5a8376} /* (16, 25, 7) {real, imag} */,
  {32'h3f57a354, 32'h3f0f18cb} /* (16, 25, 6) {real, imag} */,
  {32'h3ed2e4b7, 32'hbf0e05b9} /* (16, 25, 5) {real, imag} */,
  {32'hbf1e30fa, 32'h3e222650} /* (16, 25, 4) {real, imag} */,
  {32'hbf12fafb, 32'hbf244ca8} /* (16, 25, 3) {real, imag} */,
  {32'hbd3d9cee, 32'hbf3faccc} /* (16, 25, 2) {real, imag} */,
  {32'hbeaf3902, 32'h3f5bda08} /* (16, 25, 1) {real, imag} */,
  {32'h3e889c94, 32'hbfb3389b} /* (16, 25, 0) {real, imag} */,
  {32'hbf635952, 32'hbfdaae1f} /* (16, 24, 31) {real, imag} */,
  {32'hbf10addb, 32'hbfa6f36b} /* (16, 24, 30) {real, imag} */,
  {32'hbfcc42ee, 32'hbf929e8a} /* (16, 24, 29) {real, imag} */,
  {32'hbf7c276f, 32'h3ff3e754} /* (16, 24, 28) {real, imag} */,
  {32'h3fdc629e, 32'h3fe46f04} /* (16, 24, 27) {real, imag} */,
  {32'h3fc9ce86, 32'h40031045} /* (16, 24, 26) {real, imag} */,
  {32'h3f3c5b74, 32'hbf4af19e} /* (16, 24, 25) {real, imag} */,
  {32'hc0000c69, 32'h3ea0ee95} /* (16, 24, 24) {real, imag} */,
  {32'hbeacce7e, 32'hc0434bf3} /* (16, 24, 23) {real, imag} */,
  {32'hbf9f88d6, 32'hbf9138b6} /* (16, 24, 22) {real, imag} */,
  {32'hbeff02f7, 32'h3f596a31} /* (16, 24, 21) {real, imag} */,
  {32'h3fc8a03b, 32'hbf111809} /* (16, 24, 20) {real, imag} */,
  {32'hbfc262b1, 32'hbea6cd81} /* (16, 24, 19) {real, imag} */,
  {32'h3e5ef322, 32'hbddc3574} /* (16, 24, 18) {real, imag} */,
  {32'h3f11a36d, 32'hbde90e06} /* (16, 24, 17) {real, imag} */,
  {32'hbfdf913d, 32'hbde7a005} /* (16, 24, 16) {real, imag} */,
  {32'h3fe00bf8, 32'hbf5278a4} /* (16, 24, 15) {real, imag} */,
  {32'h3cdbb781, 32'h401d6e72} /* (16, 24, 14) {real, imag} */,
  {32'h3f0ac0c5, 32'hbf990185} /* (16, 24, 13) {real, imag} */,
  {32'h3f8a07f2, 32'h3f1ce123} /* (16, 24, 12) {real, imag} */,
  {32'hbf6f1c88, 32'h3f8a8d23} /* (16, 24, 11) {real, imag} */,
  {32'hbfa06117, 32'hbfa4b259} /* (16, 24, 10) {real, imag} */,
  {32'h3e8498a5, 32'h3fb11e4b} /* (16, 24, 9) {real, imag} */,
  {32'h3f94c44f, 32'hbe965870} /* (16, 24, 8) {real, imag} */,
  {32'hbd6829ce, 32'hbede5ff7} /* (16, 24, 7) {real, imag} */,
  {32'hbf9237ed, 32'h3e4bd2b7} /* (16, 24, 6) {real, imag} */,
  {32'hbf6fa4e3, 32'hbf4577bc} /* (16, 24, 5) {real, imag} */,
  {32'h3e55f090, 32'h3f99b92f} /* (16, 24, 4) {real, imag} */,
  {32'hbfdc294a, 32'h3c7d29e9} /* (16, 24, 3) {real, imag} */,
  {32'hbd0562bd, 32'h3fd9c82e} /* (16, 24, 2) {real, imag} */,
  {32'h3fda7f86, 32'hc01b5f8c} /* (16, 24, 1) {real, imag} */,
  {32'hbf07da02, 32'hbe911e1d} /* (16, 24, 0) {real, imag} */,
  {32'hbfa7fd73, 32'hbf750e1f} /* (16, 23, 31) {real, imag} */,
  {32'h3f19f314, 32'hbffbf92d} /* (16, 23, 30) {real, imag} */,
  {32'h3fcb13d9, 32'hbf887de1} /* (16, 23, 29) {real, imag} */,
  {32'hbd94835e, 32'h3f0177b7} /* (16, 23, 28) {real, imag} */,
  {32'h3dcc0b20, 32'h3f8bc103} /* (16, 23, 27) {real, imag} */,
  {32'h3fdce571, 32'hbf13c03f} /* (16, 23, 26) {real, imag} */,
  {32'h3f529ac8, 32'hbe390768} /* (16, 23, 25) {real, imag} */,
  {32'hbfec6086, 32'hc021c55f} /* (16, 23, 24) {real, imag} */,
  {32'h3f0e0396, 32'h3f551e71} /* (16, 23, 23) {real, imag} */,
  {32'hbfe30434, 32'h3dfd72c7} /* (16, 23, 22) {real, imag} */,
  {32'hbfb73093, 32'hbf4ec302} /* (16, 23, 21) {real, imag} */,
  {32'h3f0f156c, 32'h3f9a92eb} /* (16, 23, 20) {real, imag} */,
  {32'hbf11d4da, 32'h3fdf2524} /* (16, 23, 19) {real, imag} */,
  {32'hc046729c, 32'hbdf6b56e} /* (16, 23, 18) {real, imag} */,
  {32'h3ec32560, 32'hc01e494d} /* (16, 23, 17) {real, imag} */,
  {32'hbfb07b8d, 32'h3f3e41a1} /* (16, 23, 16) {real, imag} */,
  {32'hbe67cbf7, 32'hbf4f286b} /* (16, 23, 15) {real, imag} */,
  {32'h400b376c, 32'h3d5f25e0} /* (16, 23, 14) {real, imag} */,
  {32'hc05de14c, 32'h3fb6cb11} /* (16, 23, 13) {real, imag} */,
  {32'h3e42327f, 32'hc0381e04} /* (16, 23, 12) {real, imag} */,
  {32'hc0222fe3, 32'hbfeba4d5} /* (16, 23, 11) {real, imag} */,
  {32'h3d11c510, 32'hc01d4428} /* (16, 23, 10) {real, imag} */,
  {32'hbf91ce16, 32'hbf22f3c0} /* (16, 23, 9) {real, imag} */,
  {32'hbffed027, 32'h3fb44eb6} /* (16, 23, 8) {real, imag} */,
  {32'h3f2d9337, 32'hbf1a6f0b} /* (16, 23, 7) {real, imag} */,
  {32'h3dab0b8a, 32'h3f52054a} /* (16, 23, 6) {real, imag} */,
  {32'h3fc414ce, 32'h3f63809c} /* (16, 23, 5) {real, imag} */,
  {32'hbf476391, 32'h3dfc36dd} /* (16, 23, 4) {real, imag} */,
  {32'hbf9a6978, 32'hbeaedc79} /* (16, 23, 3) {real, imag} */,
  {32'hbfb6ade5, 32'hbf99b1bf} /* (16, 23, 2) {real, imag} */,
  {32'h3fc451d3, 32'hc0051999} /* (16, 23, 1) {real, imag} */,
  {32'h3ccff897, 32'hbfb1d5e9} /* (16, 23, 0) {real, imag} */,
  {32'hbfd58dbe, 32'h3f504385} /* (16, 22, 31) {real, imag} */,
  {32'hbed149fa, 32'hbf8e525f} /* (16, 22, 30) {real, imag} */,
  {32'hbff8b181, 32'h3dc79247} /* (16, 22, 29) {real, imag} */,
  {32'hbf380c7f, 32'h3fbcedfe} /* (16, 22, 28) {real, imag} */,
  {32'hbe0528d2, 32'hbf8e4d3c} /* (16, 22, 27) {real, imag} */,
  {32'h3e3f965a, 32'hc04b004e} /* (16, 22, 26) {real, imag} */,
  {32'h3e2c0012, 32'hbf3b3cf4} /* (16, 22, 25) {real, imag} */,
  {32'h3f3d5fad, 32'h3f94ae46} /* (16, 22, 24) {real, imag} */,
  {32'hc0037ca8, 32'hbf8e5818} /* (16, 22, 23) {real, imag} */,
  {32'hbe94cf41, 32'hbed3d230} /* (16, 22, 22) {real, imag} */,
  {32'h40393936, 32'h3f9255e2} /* (16, 22, 21) {real, imag} */,
  {32'h3f0083b2, 32'h3ff41371} /* (16, 22, 20) {real, imag} */,
  {32'h3fae1459, 32'hbfc97905} /* (16, 22, 19) {real, imag} */,
  {32'hbe7783b0, 32'hbfe041f2} /* (16, 22, 18) {real, imag} */,
  {32'hbe318f09, 32'hbf4a4da3} /* (16, 22, 17) {real, imag} */,
  {32'hbcfdb28d, 32'hbfdcb57e} /* (16, 22, 16) {real, imag} */,
  {32'h3ea8e5f4, 32'h3fb97f12} /* (16, 22, 15) {real, imag} */,
  {32'hbf347f2d, 32'hbf8e515f} /* (16, 22, 14) {real, imag} */,
  {32'hbd3885ac, 32'hc004c7e1} /* (16, 22, 13) {real, imag} */,
  {32'h40028de0, 32'h3f3a4a96} /* (16, 22, 12) {real, imag} */,
  {32'hbe85ec53, 32'h406483f2} /* (16, 22, 11) {real, imag} */,
  {32'h3f238cbf, 32'h3f70eddb} /* (16, 22, 10) {real, imag} */,
  {32'h3f58eaf7, 32'hbfb96035} /* (16, 22, 9) {real, imag} */,
  {32'hbf48140c, 32'h3f5fbe49} /* (16, 22, 8) {real, imag} */,
  {32'hbfb2f34f, 32'h3f355cc0} /* (16, 22, 7) {real, imag} */,
  {32'hbf553d33, 32'h4008ee36} /* (16, 22, 6) {real, imag} */,
  {32'h3f141843, 32'hbf605f4b} /* (16, 22, 5) {real, imag} */,
  {32'hc004e02c, 32'h3ec74d8c} /* (16, 22, 4) {real, imag} */,
  {32'hbfa973bf, 32'hbf33a8c0} /* (16, 22, 3) {real, imag} */,
  {32'hbee476f5, 32'h3f5edf62} /* (16, 22, 2) {real, imag} */,
  {32'hbeef5b61, 32'hbf872caa} /* (16, 22, 1) {real, imag} */,
  {32'h400f8ac3, 32'h3fbe9a9c} /* (16, 22, 0) {real, imag} */,
  {32'hbeb972a0, 32'hbf8bb050} /* (16, 21, 31) {real, imag} */,
  {32'h3fcd2933, 32'hbed68030} /* (16, 21, 30) {real, imag} */,
  {32'hbf6aaaed, 32'hc027f217} /* (16, 21, 29) {real, imag} */,
  {32'h3ddd665e, 32'hbff4f6bf} /* (16, 21, 28) {real, imag} */,
  {32'hbf2eb6b6, 32'h3f75da70} /* (16, 21, 27) {real, imag} */,
  {32'hbd2271f7, 32'h3eb2ca56} /* (16, 21, 26) {real, imag} */,
  {32'h3fe1f979, 32'hbdc9d1e8} /* (16, 21, 25) {real, imag} */,
  {32'hbf9bd54e, 32'h3f993b43} /* (16, 21, 24) {real, imag} */,
  {32'hbfc485eb, 32'hbfd1f611} /* (16, 21, 23) {real, imag} */,
  {32'hbf65bf28, 32'hc0141e2d} /* (16, 21, 22) {real, imag} */,
  {32'h3d8391f4, 32'h3fd7f880} /* (16, 21, 21) {real, imag} */,
  {32'h3d49b25f, 32'hbf617dae} /* (16, 21, 20) {real, imag} */,
  {32'hbfc0d10a, 32'hbf8900d1} /* (16, 21, 19) {real, imag} */,
  {32'h4055ef2a, 32'hc022498b} /* (16, 21, 18) {real, imag} */,
  {32'h3f8ef4a9, 32'h3dd948db} /* (16, 21, 17) {real, imag} */,
  {32'hbf39c917, 32'hbccbcd20} /* (16, 21, 16) {real, imag} */,
  {32'hbf5926a7, 32'hbf88f004} /* (16, 21, 15) {real, imag} */,
  {32'hbec17eba, 32'h3e6929a3} /* (16, 21, 14) {real, imag} */,
  {32'h3f0e6716, 32'hbe90b4ee} /* (16, 21, 13) {real, imag} */,
  {32'hbfc45638, 32'hbc9bd488} /* (16, 21, 12) {real, imag} */,
  {32'hbe8a9db5, 32'h3f6c53c5} /* (16, 21, 11) {real, imag} */,
  {32'h3e0aed7e, 32'h3f45737d} /* (16, 21, 10) {real, imag} */,
  {32'h3f5d6a0b, 32'h3d0ac571} /* (16, 21, 9) {real, imag} */,
  {32'h3f7171ba, 32'hbfba90c7} /* (16, 21, 8) {real, imag} */,
  {32'h3fa15c62, 32'h3f200cfc} /* (16, 21, 7) {real, imag} */,
  {32'h3f8c3275, 32'h3fbbad07} /* (16, 21, 6) {real, imag} */,
  {32'h3f1965ac, 32'h3eb87031} /* (16, 21, 5) {real, imag} */,
  {32'h3c585202, 32'hbe95e467} /* (16, 21, 4) {real, imag} */,
  {32'hbfe86aa6, 32'h3fa5ec88} /* (16, 21, 3) {real, imag} */,
  {32'hbef9acd7, 32'hbf3b20e5} /* (16, 21, 2) {real, imag} */,
  {32'hbf04f0e9, 32'hbe943399} /* (16, 21, 1) {real, imag} */,
  {32'hbe4a0d55, 32'h3fb78007} /* (16, 21, 0) {real, imag} */,
  {32'hbf9fa23f, 32'h3f82f2a3} /* (16, 20, 31) {real, imag} */,
  {32'hbf690a1e, 32'hbf88f65b} /* (16, 20, 30) {real, imag} */,
  {32'h3f5b230f, 32'hbd114101} /* (16, 20, 29) {real, imag} */,
  {32'hbdb81314, 32'hc01681c2} /* (16, 20, 28) {real, imag} */,
  {32'hbf0dd929, 32'hbfc2b038} /* (16, 20, 27) {real, imag} */,
  {32'hbf12561a, 32'hbe2c7ab0} /* (16, 20, 26) {real, imag} */,
  {32'h4044ce30, 32'hbfffc461} /* (16, 20, 25) {real, imag} */,
  {32'h3d3160c6, 32'hc0811370} /* (16, 20, 24) {real, imag} */,
  {32'hbf164d62, 32'hbfe01da1} /* (16, 20, 23) {real, imag} */,
  {32'h3e7148a0, 32'h3f5a9259} /* (16, 20, 22) {real, imag} */,
  {32'hc0582c17, 32'hbedacd86} /* (16, 20, 21) {real, imag} */,
  {32'h400c4e04, 32'h3f092c49} /* (16, 20, 20) {real, imag} */,
  {32'h401eeaee, 32'hbf7dcbc8} /* (16, 20, 19) {real, imag} */,
  {32'hbf5f547b, 32'h400accad} /* (16, 20, 18) {real, imag} */,
  {32'hc010a45f, 32'h3f4f590d} /* (16, 20, 17) {real, imag} */,
  {32'hbf4e7340, 32'hbe822c5e} /* (16, 20, 16) {real, imag} */,
  {32'hbeb34aa2, 32'h3ea13553} /* (16, 20, 15) {real, imag} */,
  {32'hbeea6dd7, 32'hc018c4ea} /* (16, 20, 14) {real, imag} */,
  {32'h3fa683df, 32'hc0362fe3} /* (16, 20, 13) {real, imag} */,
  {32'h3f48bef6, 32'h404fd052} /* (16, 20, 12) {real, imag} */,
  {32'h3f6422e5, 32'h3d172e8a} /* (16, 20, 11) {real, imag} */,
  {32'h3fdbb401, 32'hbc19fc35} /* (16, 20, 10) {real, imag} */,
  {32'hc01e33c7, 32'hbf6b1c86} /* (16, 20, 9) {real, imag} */,
  {32'hbe183123, 32'hbf5677bb} /* (16, 20, 8) {real, imag} */,
  {32'hbfd1e3af, 32'hbff336f4} /* (16, 20, 7) {real, imag} */,
  {32'hbf8f078a, 32'h3edef0e6} /* (16, 20, 6) {real, imag} */,
  {32'hbfd8b445, 32'h3dfc9c46} /* (16, 20, 5) {real, imag} */,
  {32'h400600e9, 32'hbf23ef8e} /* (16, 20, 4) {real, imag} */,
  {32'h3d156dc6, 32'h3fde57d6} /* (16, 20, 3) {real, imag} */,
  {32'hbd83e3b3, 32'hbfa248a2} /* (16, 20, 2) {real, imag} */,
  {32'hbf78bc87, 32'h3d64dd81} /* (16, 20, 1) {real, imag} */,
  {32'h401e1236, 32'h3f8a42bf} /* (16, 20, 0) {real, imag} */,
  {32'h3ffa7bd4, 32'hc026cf55} /* (16, 19, 31) {real, imag} */,
  {32'h3fd96b1d, 32'h3fd4852a} /* (16, 19, 30) {real, imag} */,
  {32'h3f5b465a, 32'h3e064f57} /* (16, 19, 29) {real, imag} */,
  {32'hc00f7e39, 32'hbfd83021} /* (16, 19, 28) {real, imag} */,
  {32'h3f54e615, 32'h3f630505} /* (16, 19, 27) {real, imag} */,
  {32'h3fd1ea90, 32'h3f3472f9} /* (16, 19, 26) {real, imag} */,
  {32'hbf87ff16, 32'h3ec7a9b2} /* (16, 19, 25) {real, imag} */,
  {32'h3f92eb5a, 32'hbe94f23d} /* (16, 19, 24) {real, imag} */,
  {32'h3e947118, 32'hbf8e107b} /* (16, 19, 23) {real, imag} */,
  {32'h3f37f4de, 32'h3fe4ab10} /* (16, 19, 22) {real, imag} */,
  {32'hbf87c2eb, 32'h400919b4} /* (16, 19, 21) {real, imag} */,
  {32'hc00044d8, 32'hbee97b1f} /* (16, 19, 20) {real, imag} */,
  {32'hbf8b53a7, 32'hc0784a6e} /* (16, 19, 19) {real, imag} */,
  {32'hbc975fee, 32'h3a70e159} /* (16, 19, 18) {real, imag} */,
  {32'hbf963353, 32'h40548b3c} /* (16, 19, 17) {real, imag} */,
  {32'h3febdb3a, 32'hbf0759c4} /* (16, 19, 16) {real, imag} */,
  {32'h3e78c5c5, 32'hbf3968ac} /* (16, 19, 15) {real, imag} */,
  {32'h3f969ea0, 32'h3daf2992} /* (16, 19, 14) {real, imag} */,
  {32'hbfa3cda3, 32'h3f8c31d0} /* (16, 19, 13) {real, imag} */,
  {32'hbf52679b, 32'h3f979f0e} /* (16, 19, 12) {real, imag} */,
  {32'h4026a699, 32'h3ffeb182} /* (16, 19, 11) {real, imag} */,
  {32'hbf06b0ec, 32'hbf2949b6} /* (16, 19, 10) {real, imag} */,
  {32'hbfc43000, 32'h3ed056c2} /* (16, 19, 9) {real, imag} */,
  {32'h3f2e47f0, 32'hbf9cab4f} /* (16, 19, 8) {real, imag} */,
  {32'h401469fb, 32'hc08d14f3} /* (16, 19, 7) {real, imag} */,
  {32'hc004688f, 32'h3e0f2d11} /* (16, 19, 6) {real, imag} */,
  {32'hbfffc1e6, 32'h3efd577a} /* (16, 19, 5) {real, imag} */,
  {32'hbfb75088, 32'h3e9a3da7} /* (16, 19, 4) {real, imag} */,
  {32'h3fcdb830, 32'h3e06aea2} /* (16, 19, 3) {real, imag} */,
  {32'h4006caf2, 32'hbe0c42af} /* (16, 19, 2) {real, imag} */,
  {32'hbf97b9f3, 32'h4011c704} /* (16, 19, 1) {real, imag} */,
  {32'hbc5055e2, 32'hbf09b690} /* (16, 19, 0) {real, imag} */,
  {32'hbf0fdcf3, 32'hbff6a37c} /* (16, 18, 31) {real, imag} */,
  {32'hbfdd6319, 32'hbf196f39} /* (16, 18, 30) {real, imag} */,
  {32'h3fe18476, 32'hbf7517ea} /* (16, 18, 29) {real, imag} */,
  {32'hbfaaeca9, 32'hbf392a2b} /* (16, 18, 28) {real, imag} */,
  {32'hbee1ccb2, 32'h3fae831c} /* (16, 18, 27) {real, imag} */,
  {32'hbfaf4d5a, 32'hbf50d547} /* (16, 18, 26) {real, imag} */,
  {32'hbedccdc7, 32'h3fcb1ddb} /* (16, 18, 25) {real, imag} */,
  {32'hc0602727, 32'h3f7d5ca7} /* (16, 18, 24) {real, imag} */,
  {32'h3f941943, 32'h3e76f951} /* (16, 18, 23) {real, imag} */,
  {32'hbfb208c6, 32'h3eb09059} /* (16, 18, 22) {real, imag} */,
  {32'hbee3b68c, 32'hbffa8877} /* (16, 18, 21) {real, imag} */,
  {32'h3eda943b, 32'h400d65fa} /* (16, 18, 20) {real, imag} */,
  {32'h3f8f4efd, 32'h3f3b2e39} /* (16, 18, 19) {real, imag} */,
  {32'h4001672b, 32'h3ef323ab} /* (16, 18, 18) {real, imag} */,
  {32'h3f33bd21, 32'hc00e3b2b} /* (16, 18, 17) {real, imag} */,
  {32'hbf3c02f2, 32'h3fd297f2} /* (16, 18, 16) {real, imag} */,
  {32'h3fa22ca1, 32'hbe24fe43} /* (16, 18, 15) {real, imag} */,
  {32'hbf7305da, 32'hbf86756b} /* (16, 18, 14) {real, imag} */,
  {32'hbf538abd, 32'hbfa0b7da} /* (16, 18, 13) {real, imag} */,
  {32'h3f52ef8b, 32'hbf3e2260} /* (16, 18, 12) {real, imag} */,
  {32'hbf48a94b, 32'h3f6a560f} /* (16, 18, 11) {real, imag} */,
  {32'hbfd99258, 32'h3dd4b4c9} /* (16, 18, 10) {real, imag} */,
  {32'hbdebf69c, 32'h3ec36549} /* (16, 18, 9) {real, imag} */,
  {32'hbf30c383, 32'h3f5901e5} /* (16, 18, 8) {real, imag} */,
  {32'h3fc5d033, 32'h3f63d2e3} /* (16, 18, 7) {real, imag} */,
  {32'h3eba2928, 32'h3f0b8f3a} /* (16, 18, 6) {real, imag} */,
  {32'h3ee611da, 32'h3f8704c0} /* (16, 18, 5) {real, imag} */,
  {32'h3f83ebe4, 32'h3febb359} /* (16, 18, 4) {real, imag} */,
  {32'hbd6625f2, 32'hbefb3a2f} /* (16, 18, 3) {real, imag} */,
  {32'h3ecfe43b, 32'h3e97a596} /* (16, 18, 2) {real, imag} */,
  {32'h3e50f9c2, 32'h3f7a58f6} /* (16, 18, 1) {real, imag} */,
  {32'h3fc181f1, 32'hbf1f2c18} /* (16, 18, 0) {real, imag} */,
  {32'hbdefc591, 32'h3fb9d62c} /* (16, 17, 31) {real, imag} */,
  {32'hbf7e8fd8, 32'h3f6d3cf7} /* (16, 17, 30) {real, imag} */,
  {32'h3f10c267, 32'hbe960e76} /* (16, 17, 29) {real, imag} */,
  {32'h3f5d2215, 32'h3f3788db} /* (16, 17, 28) {real, imag} */,
  {32'hbf77d7cb, 32'h3f3f6c2b} /* (16, 17, 27) {real, imag} */,
  {32'hbf7a43cf, 32'hbf4e65a6} /* (16, 17, 26) {real, imag} */,
  {32'h3e0d3c83, 32'hc00503a9} /* (16, 17, 25) {real, imag} */,
  {32'h3e22df8a, 32'hbf197b0a} /* (16, 17, 24) {real, imag} */,
  {32'hbf578e05, 32'hbe2f4f1d} /* (16, 17, 23) {real, imag} */,
  {32'hbea898ce, 32'hbf3ba9c1} /* (16, 17, 22) {real, imag} */,
  {32'h3f670333, 32'h40075337} /* (16, 17, 21) {real, imag} */,
  {32'h3d4123a7, 32'h3e8e4ab1} /* (16, 17, 20) {real, imag} */,
  {32'h3f8aa759, 32'hbe7e2d76} /* (16, 17, 19) {real, imag} */,
  {32'hc0022e4c, 32'h3f54bd4d} /* (16, 17, 18) {real, imag} */,
  {32'hbfab277b, 32'h3e993ddc} /* (16, 17, 17) {real, imag} */,
  {32'h3f7e4f98, 32'h3ecb4c70} /* (16, 17, 16) {real, imag} */,
  {32'hbef2c9ba, 32'h3f9ba8bc} /* (16, 17, 15) {real, imag} */,
  {32'hbef9c176, 32'h3f952c12} /* (16, 17, 14) {real, imag} */,
  {32'hbef3125e, 32'hc00afeec} /* (16, 17, 13) {real, imag} */,
  {32'hbf4885f7, 32'h3f27d9cd} /* (16, 17, 12) {real, imag} */,
  {32'h3f053790, 32'hbfa82624} /* (16, 17, 11) {real, imag} */,
  {32'h3eaf18f4, 32'hbc8872ea} /* (16, 17, 10) {real, imag} */,
  {32'h3fd7f161, 32'hbe577d02} /* (16, 17, 9) {real, imag} */,
  {32'h3f3b4fd6, 32'h3fb0af5f} /* (16, 17, 8) {real, imag} */,
  {32'hbfbccfe1, 32'h3ed82e6c} /* (16, 17, 7) {real, imag} */,
  {32'hbe12b417, 32'hbf413610} /* (16, 17, 6) {real, imag} */,
  {32'h3fd2479f, 32'h3f60729c} /* (16, 17, 5) {real, imag} */,
  {32'hbfd3d6b5, 32'hbfaf2170} /* (16, 17, 4) {real, imag} */,
  {32'hbf14f8f4, 32'hbd3169ab} /* (16, 17, 3) {real, imag} */,
  {32'hbfacf781, 32'hbed956bf} /* (16, 17, 2) {real, imag} */,
  {32'h3f381435, 32'hbfa35107} /* (16, 17, 1) {real, imag} */,
  {32'hbff0f4fb, 32'h3f4c8c64} /* (16, 17, 0) {real, imag} */,
  {32'hbf0629a8, 32'hbf1819d2} /* (16, 16, 31) {real, imag} */,
  {32'h3f0e7f12, 32'hbe85a012} /* (16, 16, 30) {real, imag} */,
  {32'hc0343621, 32'h3ec674fb} /* (16, 16, 29) {real, imag} */,
  {32'h3f24d3e6, 32'h3fa92885} /* (16, 16, 28) {real, imag} */,
  {32'h3e078fcb, 32'hbe7840ae} /* (16, 16, 27) {real, imag} */,
  {32'h3ea71ed6, 32'hbe61c0ea} /* (16, 16, 26) {real, imag} */,
  {32'h3f68e4d2, 32'h3f318ab1} /* (16, 16, 25) {real, imag} */,
  {32'hbe20d034, 32'h3e3ec59b} /* (16, 16, 24) {real, imag} */,
  {32'hbd6c79a0, 32'h3e81cdc7} /* (16, 16, 23) {real, imag} */,
  {32'hbe90cc39, 32'hbe8bed28} /* (16, 16, 22) {real, imag} */,
  {32'h3f39ba90, 32'hbe54197b} /* (16, 16, 21) {real, imag} */,
  {32'h3d259a65, 32'hbf9c8b6d} /* (16, 16, 20) {real, imag} */,
  {32'h3fbf7c3c, 32'h3fa2f255} /* (16, 16, 19) {real, imag} */,
  {32'hbf2ab019, 32'hbf3eeef4} /* (16, 16, 18) {real, imag} */,
  {32'h3f651750, 32'hbf3803fb} /* (16, 16, 17) {real, imag} */,
  {32'hbffa903d, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h3f651750, 32'h3f3803fb} /* (16, 16, 15) {real, imag} */,
  {32'hbf2ab019, 32'h3f3eeef4} /* (16, 16, 14) {real, imag} */,
  {32'h3fbf7c3c, 32'hbfa2f255} /* (16, 16, 13) {real, imag} */,
  {32'h3d259a65, 32'h3f9c8b6d} /* (16, 16, 12) {real, imag} */,
  {32'h3f39ba90, 32'h3e54197b} /* (16, 16, 11) {real, imag} */,
  {32'hbe90cc39, 32'h3e8bed28} /* (16, 16, 10) {real, imag} */,
  {32'hbd6c79a0, 32'hbe81cdc7} /* (16, 16, 9) {real, imag} */,
  {32'hbe20d034, 32'hbe3ec59b} /* (16, 16, 8) {real, imag} */,
  {32'h3f68e4d2, 32'hbf318ab1} /* (16, 16, 7) {real, imag} */,
  {32'h3ea71ed6, 32'h3e61c0ea} /* (16, 16, 6) {real, imag} */,
  {32'h3e078fcb, 32'h3e7840ae} /* (16, 16, 5) {real, imag} */,
  {32'h3f24d3e6, 32'hbfa92885} /* (16, 16, 4) {real, imag} */,
  {32'hc0343621, 32'hbec674fb} /* (16, 16, 3) {real, imag} */,
  {32'h3f0e7f12, 32'h3e85a012} /* (16, 16, 2) {real, imag} */,
  {32'hbf0629a8, 32'h3f1819d2} /* (16, 16, 1) {real, imag} */,
  {32'h3f80a32a, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h3f381435, 32'h3fa35107} /* (16, 15, 31) {real, imag} */,
  {32'hbfacf781, 32'h3ed956bf} /* (16, 15, 30) {real, imag} */,
  {32'hbf14f8f4, 32'h3d3169ab} /* (16, 15, 29) {real, imag} */,
  {32'hbfd3d6b5, 32'h3faf2170} /* (16, 15, 28) {real, imag} */,
  {32'h3fd2479f, 32'hbf60729c} /* (16, 15, 27) {real, imag} */,
  {32'hbe12b417, 32'h3f413610} /* (16, 15, 26) {real, imag} */,
  {32'hbfbccfe1, 32'hbed82e6c} /* (16, 15, 25) {real, imag} */,
  {32'h3f3b4fd6, 32'hbfb0af5f} /* (16, 15, 24) {real, imag} */,
  {32'h3fd7f161, 32'h3e577d02} /* (16, 15, 23) {real, imag} */,
  {32'h3eaf18f4, 32'h3c8872ea} /* (16, 15, 22) {real, imag} */,
  {32'h3f053790, 32'h3fa82624} /* (16, 15, 21) {real, imag} */,
  {32'hbf4885f7, 32'hbf27d9cd} /* (16, 15, 20) {real, imag} */,
  {32'hbef3125e, 32'h400afeec} /* (16, 15, 19) {real, imag} */,
  {32'hbef9c176, 32'hbf952c12} /* (16, 15, 18) {real, imag} */,
  {32'hbef2c9ba, 32'hbf9ba8bc} /* (16, 15, 17) {real, imag} */,
  {32'h3f7e4f98, 32'hbecb4c70} /* (16, 15, 16) {real, imag} */,
  {32'hbfab277b, 32'hbe993ddc} /* (16, 15, 15) {real, imag} */,
  {32'hc0022e4c, 32'hbf54bd4d} /* (16, 15, 14) {real, imag} */,
  {32'h3f8aa759, 32'h3e7e2d76} /* (16, 15, 13) {real, imag} */,
  {32'h3d4123a7, 32'hbe8e4ab1} /* (16, 15, 12) {real, imag} */,
  {32'h3f670333, 32'hc0075337} /* (16, 15, 11) {real, imag} */,
  {32'hbea898ce, 32'h3f3ba9c1} /* (16, 15, 10) {real, imag} */,
  {32'hbf578e05, 32'h3e2f4f1d} /* (16, 15, 9) {real, imag} */,
  {32'h3e22df8a, 32'h3f197b0a} /* (16, 15, 8) {real, imag} */,
  {32'h3e0d3c83, 32'h400503a9} /* (16, 15, 7) {real, imag} */,
  {32'hbf7a43cf, 32'h3f4e65a6} /* (16, 15, 6) {real, imag} */,
  {32'hbf77d7cb, 32'hbf3f6c2b} /* (16, 15, 5) {real, imag} */,
  {32'h3f5d2215, 32'hbf3788db} /* (16, 15, 4) {real, imag} */,
  {32'h3f10c267, 32'h3e960e76} /* (16, 15, 3) {real, imag} */,
  {32'hbf7e8fd8, 32'hbf6d3cf7} /* (16, 15, 2) {real, imag} */,
  {32'hbdefc591, 32'hbfb9d62c} /* (16, 15, 1) {real, imag} */,
  {32'hbff0f4fb, 32'hbf4c8c64} /* (16, 15, 0) {real, imag} */,
  {32'h3e50f9c2, 32'hbf7a58f6} /* (16, 14, 31) {real, imag} */,
  {32'h3ecfe43b, 32'hbe97a596} /* (16, 14, 30) {real, imag} */,
  {32'hbd6625f2, 32'h3efb3a2f} /* (16, 14, 29) {real, imag} */,
  {32'h3f83ebe4, 32'hbfebb359} /* (16, 14, 28) {real, imag} */,
  {32'h3ee611da, 32'hbf8704c0} /* (16, 14, 27) {real, imag} */,
  {32'h3eba2928, 32'hbf0b8f3a} /* (16, 14, 26) {real, imag} */,
  {32'h3fc5d033, 32'hbf63d2e3} /* (16, 14, 25) {real, imag} */,
  {32'hbf30c383, 32'hbf5901e5} /* (16, 14, 24) {real, imag} */,
  {32'hbdebf69c, 32'hbec36549} /* (16, 14, 23) {real, imag} */,
  {32'hbfd99258, 32'hbdd4b4c9} /* (16, 14, 22) {real, imag} */,
  {32'hbf48a94b, 32'hbf6a560f} /* (16, 14, 21) {real, imag} */,
  {32'h3f52ef8b, 32'h3f3e2260} /* (16, 14, 20) {real, imag} */,
  {32'hbf538abd, 32'h3fa0b7da} /* (16, 14, 19) {real, imag} */,
  {32'hbf7305da, 32'h3f86756b} /* (16, 14, 18) {real, imag} */,
  {32'h3fa22ca1, 32'h3e24fe43} /* (16, 14, 17) {real, imag} */,
  {32'hbf3c02f2, 32'hbfd297f2} /* (16, 14, 16) {real, imag} */,
  {32'h3f33bd21, 32'h400e3b2b} /* (16, 14, 15) {real, imag} */,
  {32'h4001672b, 32'hbef323ab} /* (16, 14, 14) {real, imag} */,
  {32'h3f8f4efd, 32'hbf3b2e39} /* (16, 14, 13) {real, imag} */,
  {32'h3eda943b, 32'hc00d65fa} /* (16, 14, 12) {real, imag} */,
  {32'hbee3b68c, 32'h3ffa8877} /* (16, 14, 11) {real, imag} */,
  {32'hbfb208c6, 32'hbeb09059} /* (16, 14, 10) {real, imag} */,
  {32'h3f941943, 32'hbe76f951} /* (16, 14, 9) {real, imag} */,
  {32'hc0602727, 32'hbf7d5ca7} /* (16, 14, 8) {real, imag} */,
  {32'hbedccdc7, 32'hbfcb1ddb} /* (16, 14, 7) {real, imag} */,
  {32'hbfaf4d5a, 32'h3f50d547} /* (16, 14, 6) {real, imag} */,
  {32'hbee1ccb2, 32'hbfae831c} /* (16, 14, 5) {real, imag} */,
  {32'hbfaaeca9, 32'h3f392a2b} /* (16, 14, 4) {real, imag} */,
  {32'h3fe18476, 32'h3f7517ea} /* (16, 14, 3) {real, imag} */,
  {32'hbfdd6319, 32'h3f196f39} /* (16, 14, 2) {real, imag} */,
  {32'hbf0fdcf3, 32'h3ff6a37c} /* (16, 14, 1) {real, imag} */,
  {32'h3fc181f1, 32'h3f1f2c18} /* (16, 14, 0) {real, imag} */,
  {32'hbf97b9f3, 32'hc011c704} /* (16, 13, 31) {real, imag} */,
  {32'h4006caf2, 32'h3e0c42af} /* (16, 13, 30) {real, imag} */,
  {32'h3fcdb830, 32'hbe06aea2} /* (16, 13, 29) {real, imag} */,
  {32'hbfb75088, 32'hbe9a3da7} /* (16, 13, 28) {real, imag} */,
  {32'hbfffc1e6, 32'hbefd577a} /* (16, 13, 27) {real, imag} */,
  {32'hc004688f, 32'hbe0f2d11} /* (16, 13, 26) {real, imag} */,
  {32'h401469fb, 32'h408d14f3} /* (16, 13, 25) {real, imag} */,
  {32'h3f2e47f0, 32'h3f9cab4f} /* (16, 13, 24) {real, imag} */,
  {32'hbfc43000, 32'hbed056c2} /* (16, 13, 23) {real, imag} */,
  {32'hbf06b0ec, 32'h3f2949b6} /* (16, 13, 22) {real, imag} */,
  {32'h4026a699, 32'hbffeb182} /* (16, 13, 21) {real, imag} */,
  {32'hbf52679b, 32'hbf979f0e} /* (16, 13, 20) {real, imag} */,
  {32'hbfa3cda3, 32'hbf8c31d0} /* (16, 13, 19) {real, imag} */,
  {32'h3f969ea0, 32'hbdaf2992} /* (16, 13, 18) {real, imag} */,
  {32'h3e78c5c5, 32'h3f3968ac} /* (16, 13, 17) {real, imag} */,
  {32'h3febdb3a, 32'h3f0759c4} /* (16, 13, 16) {real, imag} */,
  {32'hbf963353, 32'hc0548b3c} /* (16, 13, 15) {real, imag} */,
  {32'hbc975fee, 32'hba70e159} /* (16, 13, 14) {real, imag} */,
  {32'hbf8b53a7, 32'h40784a6e} /* (16, 13, 13) {real, imag} */,
  {32'hc00044d8, 32'h3ee97b1f} /* (16, 13, 12) {real, imag} */,
  {32'hbf87c2eb, 32'hc00919b4} /* (16, 13, 11) {real, imag} */,
  {32'h3f37f4de, 32'hbfe4ab10} /* (16, 13, 10) {real, imag} */,
  {32'h3e947118, 32'h3f8e107b} /* (16, 13, 9) {real, imag} */,
  {32'h3f92eb5a, 32'h3e94f23d} /* (16, 13, 8) {real, imag} */,
  {32'hbf87ff16, 32'hbec7a9b2} /* (16, 13, 7) {real, imag} */,
  {32'h3fd1ea90, 32'hbf3472f9} /* (16, 13, 6) {real, imag} */,
  {32'h3f54e615, 32'hbf630505} /* (16, 13, 5) {real, imag} */,
  {32'hc00f7e39, 32'h3fd83021} /* (16, 13, 4) {real, imag} */,
  {32'h3f5b465a, 32'hbe064f57} /* (16, 13, 3) {real, imag} */,
  {32'h3fd96b1d, 32'hbfd4852a} /* (16, 13, 2) {real, imag} */,
  {32'h3ffa7bd4, 32'h4026cf55} /* (16, 13, 1) {real, imag} */,
  {32'hbc5055e2, 32'h3f09b690} /* (16, 13, 0) {real, imag} */,
  {32'hbf78bc87, 32'hbd64dd81} /* (16, 12, 31) {real, imag} */,
  {32'hbd83e3b3, 32'h3fa248a2} /* (16, 12, 30) {real, imag} */,
  {32'h3d156dc6, 32'hbfde57d6} /* (16, 12, 29) {real, imag} */,
  {32'h400600e9, 32'h3f23ef8e} /* (16, 12, 28) {real, imag} */,
  {32'hbfd8b445, 32'hbdfc9c46} /* (16, 12, 27) {real, imag} */,
  {32'hbf8f078a, 32'hbedef0e6} /* (16, 12, 26) {real, imag} */,
  {32'hbfd1e3af, 32'h3ff336f4} /* (16, 12, 25) {real, imag} */,
  {32'hbe183123, 32'h3f5677bb} /* (16, 12, 24) {real, imag} */,
  {32'hc01e33c7, 32'h3f6b1c86} /* (16, 12, 23) {real, imag} */,
  {32'h3fdbb401, 32'h3c19fc35} /* (16, 12, 22) {real, imag} */,
  {32'h3f6422e5, 32'hbd172e8a} /* (16, 12, 21) {real, imag} */,
  {32'h3f48bef6, 32'hc04fd052} /* (16, 12, 20) {real, imag} */,
  {32'h3fa683df, 32'h40362fe3} /* (16, 12, 19) {real, imag} */,
  {32'hbeea6dd7, 32'h4018c4ea} /* (16, 12, 18) {real, imag} */,
  {32'hbeb34aa2, 32'hbea13553} /* (16, 12, 17) {real, imag} */,
  {32'hbf4e7340, 32'h3e822c5e} /* (16, 12, 16) {real, imag} */,
  {32'hc010a45f, 32'hbf4f590d} /* (16, 12, 15) {real, imag} */,
  {32'hbf5f547b, 32'hc00accad} /* (16, 12, 14) {real, imag} */,
  {32'h401eeaee, 32'h3f7dcbc8} /* (16, 12, 13) {real, imag} */,
  {32'h400c4e04, 32'hbf092c49} /* (16, 12, 12) {real, imag} */,
  {32'hc0582c17, 32'h3edacd86} /* (16, 12, 11) {real, imag} */,
  {32'h3e7148a0, 32'hbf5a9259} /* (16, 12, 10) {real, imag} */,
  {32'hbf164d62, 32'h3fe01da1} /* (16, 12, 9) {real, imag} */,
  {32'h3d3160c6, 32'h40811370} /* (16, 12, 8) {real, imag} */,
  {32'h4044ce30, 32'h3fffc461} /* (16, 12, 7) {real, imag} */,
  {32'hbf12561a, 32'h3e2c7ab0} /* (16, 12, 6) {real, imag} */,
  {32'hbf0dd929, 32'h3fc2b038} /* (16, 12, 5) {real, imag} */,
  {32'hbdb81314, 32'h401681c2} /* (16, 12, 4) {real, imag} */,
  {32'h3f5b230f, 32'h3d114101} /* (16, 12, 3) {real, imag} */,
  {32'hbf690a1e, 32'h3f88f65b} /* (16, 12, 2) {real, imag} */,
  {32'hbf9fa23f, 32'hbf82f2a3} /* (16, 12, 1) {real, imag} */,
  {32'h401e1236, 32'hbf8a42bf} /* (16, 12, 0) {real, imag} */,
  {32'hbf04f0e9, 32'h3e943399} /* (16, 11, 31) {real, imag} */,
  {32'hbef9acd7, 32'h3f3b20e5} /* (16, 11, 30) {real, imag} */,
  {32'hbfe86aa6, 32'hbfa5ec88} /* (16, 11, 29) {real, imag} */,
  {32'h3c585202, 32'h3e95e467} /* (16, 11, 28) {real, imag} */,
  {32'h3f1965ac, 32'hbeb87031} /* (16, 11, 27) {real, imag} */,
  {32'h3f8c3275, 32'hbfbbad07} /* (16, 11, 26) {real, imag} */,
  {32'h3fa15c62, 32'hbf200cfc} /* (16, 11, 25) {real, imag} */,
  {32'h3f7171ba, 32'h3fba90c7} /* (16, 11, 24) {real, imag} */,
  {32'h3f5d6a0b, 32'hbd0ac571} /* (16, 11, 23) {real, imag} */,
  {32'h3e0aed7e, 32'hbf45737d} /* (16, 11, 22) {real, imag} */,
  {32'hbe8a9db5, 32'hbf6c53c5} /* (16, 11, 21) {real, imag} */,
  {32'hbfc45638, 32'h3c9bd488} /* (16, 11, 20) {real, imag} */,
  {32'h3f0e6716, 32'h3e90b4ee} /* (16, 11, 19) {real, imag} */,
  {32'hbec17eba, 32'hbe6929a3} /* (16, 11, 18) {real, imag} */,
  {32'hbf5926a7, 32'h3f88f004} /* (16, 11, 17) {real, imag} */,
  {32'hbf39c917, 32'h3ccbcd20} /* (16, 11, 16) {real, imag} */,
  {32'h3f8ef4a9, 32'hbdd948db} /* (16, 11, 15) {real, imag} */,
  {32'h4055ef2a, 32'h4022498b} /* (16, 11, 14) {real, imag} */,
  {32'hbfc0d10a, 32'h3f8900d1} /* (16, 11, 13) {real, imag} */,
  {32'h3d49b25f, 32'h3f617dae} /* (16, 11, 12) {real, imag} */,
  {32'h3d8391f4, 32'hbfd7f880} /* (16, 11, 11) {real, imag} */,
  {32'hbf65bf28, 32'h40141e2d} /* (16, 11, 10) {real, imag} */,
  {32'hbfc485eb, 32'h3fd1f611} /* (16, 11, 9) {real, imag} */,
  {32'hbf9bd54e, 32'hbf993b43} /* (16, 11, 8) {real, imag} */,
  {32'h3fe1f979, 32'h3dc9d1e8} /* (16, 11, 7) {real, imag} */,
  {32'hbd2271f7, 32'hbeb2ca56} /* (16, 11, 6) {real, imag} */,
  {32'hbf2eb6b6, 32'hbf75da70} /* (16, 11, 5) {real, imag} */,
  {32'h3ddd665e, 32'h3ff4f6bf} /* (16, 11, 4) {real, imag} */,
  {32'hbf6aaaed, 32'h4027f217} /* (16, 11, 3) {real, imag} */,
  {32'h3fcd2933, 32'h3ed68030} /* (16, 11, 2) {real, imag} */,
  {32'hbeb972a0, 32'h3f8bb050} /* (16, 11, 1) {real, imag} */,
  {32'hbe4a0d55, 32'hbfb78007} /* (16, 11, 0) {real, imag} */,
  {32'hbeef5b61, 32'h3f872caa} /* (16, 10, 31) {real, imag} */,
  {32'hbee476f5, 32'hbf5edf62} /* (16, 10, 30) {real, imag} */,
  {32'hbfa973bf, 32'h3f33a8c0} /* (16, 10, 29) {real, imag} */,
  {32'hc004e02c, 32'hbec74d8c} /* (16, 10, 28) {real, imag} */,
  {32'h3f141843, 32'h3f605f4b} /* (16, 10, 27) {real, imag} */,
  {32'hbf553d33, 32'hc008ee36} /* (16, 10, 26) {real, imag} */,
  {32'hbfb2f34f, 32'hbf355cc0} /* (16, 10, 25) {real, imag} */,
  {32'hbf48140c, 32'hbf5fbe49} /* (16, 10, 24) {real, imag} */,
  {32'h3f58eaf7, 32'h3fb96035} /* (16, 10, 23) {real, imag} */,
  {32'h3f238cbf, 32'hbf70eddb} /* (16, 10, 22) {real, imag} */,
  {32'hbe85ec53, 32'hc06483f2} /* (16, 10, 21) {real, imag} */,
  {32'h40028de0, 32'hbf3a4a96} /* (16, 10, 20) {real, imag} */,
  {32'hbd3885ac, 32'h4004c7e1} /* (16, 10, 19) {real, imag} */,
  {32'hbf347f2d, 32'h3f8e515f} /* (16, 10, 18) {real, imag} */,
  {32'h3ea8e5f4, 32'hbfb97f12} /* (16, 10, 17) {real, imag} */,
  {32'hbcfdb28d, 32'h3fdcb57e} /* (16, 10, 16) {real, imag} */,
  {32'hbe318f09, 32'h3f4a4da3} /* (16, 10, 15) {real, imag} */,
  {32'hbe7783b0, 32'h3fe041f2} /* (16, 10, 14) {real, imag} */,
  {32'h3fae1459, 32'h3fc97905} /* (16, 10, 13) {real, imag} */,
  {32'h3f0083b2, 32'hbff41371} /* (16, 10, 12) {real, imag} */,
  {32'h40393936, 32'hbf9255e2} /* (16, 10, 11) {real, imag} */,
  {32'hbe94cf41, 32'h3ed3d230} /* (16, 10, 10) {real, imag} */,
  {32'hc0037ca8, 32'h3f8e5818} /* (16, 10, 9) {real, imag} */,
  {32'h3f3d5fad, 32'hbf94ae46} /* (16, 10, 8) {real, imag} */,
  {32'h3e2c0012, 32'h3f3b3cf4} /* (16, 10, 7) {real, imag} */,
  {32'h3e3f965a, 32'h404b004e} /* (16, 10, 6) {real, imag} */,
  {32'hbe0528d2, 32'h3f8e4d3c} /* (16, 10, 5) {real, imag} */,
  {32'hbf380c7f, 32'hbfbcedfe} /* (16, 10, 4) {real, imag} */,
  {32'hbff8b181, 32'hbdc79247} /* (16, 10, 3) {real, imag} */,
  {32'hbed149fa, 32'h3f8e525f} /* (16, 10, 2) {real, imag} */,
  {32'hbfd58dbe, 32'hbf504385} /* (16, 10, 1) {real, imag} */,
  {32'h400f8ac3, 32'hbfbe9a9c} /* (16, 10, 0) {real, imag} */,
  {32'h3fc451d3, 32'h40051999} /* (16, 9, 31) {real, imag} */,
  {32'hbfb6ade5, 32'h3f99b1bf} /* (16, 9, 30) {real, imag} */,
  {32'hbf9a6978, 32'h3eaedc79} /* (16, 9, 29) {real, imag} */,
  {32'hbf476391, 32'hbdfc36dd} /* (16, 9, 28) {real, imag} */,
  {32'h3fc414ce, 32'hbf63809c} /* (16, 9, 27) {real, imag} */,
  {32'h3dab0b8a, 32'hbf52054a} /* (16, 9, 26) {real, imag} */,
  {32'h3f2d9337, 32'h3f1a6f0b} /* (16, 9, 25) {real, imag} */,
  {32'hbffed027, 32'hbfb44eb6} /* (16, 9, 24) {real, imag} */,
  {32'hbf91ce16, 32'h3f22f3c0} /* (16, 9, 23) {real, imag} */,
  {32'h3d11c510, 32'h401d4428} /* (16, 9, 22) {real, imag} */,
  {32'hc0222fe3, 32'h3feba4d5} /* (16, 9, 21) {real, imag} */,
  {32'h3e42327f, 32'h40381e04} /* (16, 9, 20) {real, imag} */,
  {32'hc05de14c, 32'hbfb6cb11} /* (16, 9, 19) {real, imag} */,
  {32'h400b376c, 32'hbd5f25e0} /* (16, 9, 18) {real, imag} */,
  {32'hbe67cbf7, 32'h3f4f286b} /* (16, 9, 17) {real, imag} */,
  {32'hbfb07b8d, 32'hbf3e41a1} /* (16, 9, 16) {real, imag} */,
  {32'h3ec32560, 32'h401e494d} /* (16, 9, 15) {real, imag} */,
  {32'hc046729c, 32'h3df6b56e} /* (16, 9, 14) {real, imag} */,
  {32'hbf11d4da, 32'hbfdf2524} /* (16, 9, 13) {real, imag} */,
  {32'h3f0f156c, 32'hbf9a92eb} /* (16, 9, 12) {real, imag} */,
  {32'hbfb73093, 32'h3f4ec302} /* (16, 9, 11) {real, imag} */,
  {32'hbfe30434, 32'hbdfd72c7} /* (16, 9, 10) {real, imag} */,
  {32'h3f0e0396, 32'hbf551e71} /* (16, 9, 9) {real, imag} */,
  {32'hbfec6086, 32'h4021c55f} /* (16, 9, 8) {real, imag} */,
  {32'h3f529ac8, 32'h3e390768} /* (16, 9, 7) {real, imag} */,
  {32'h3fdce571, 32'h3f13c03f} /* (16, 9, 6) {real, imag} */,
  {32'h3dcc0b20, 32'hbf8bc103} /* (16, 9, 5) {real, imag} */,
  {32'hbd94835e, 32'hbf0177b7} /* (16, 9, 4) {real, imag} */,
  {32'h3fcb13d9, 32'h3f887de1} /* (16, 9, 3) {real, imag} */,
  {32'h3f19f314, 32'h3ffbf92d} /* (16, 9, 2) {real, imag} */,
  {32'hbfa7fd73, 32'h3f750e1f} /* (16, 9, 1) {real, imag} */,
  {32'h3ccff897, 32'h3fb1d5e9} /* (16, 9, 0) {real, imag} */,
  {32'h3fda7f86, 32'h401b5f8c} /* (16, 8, 31) {real, imag} */,
  {32'hbd0562bd, 32'hbfd9c82e} /* (16, 8, 30) {real, imag} */,
  {32'hbfdc294a, 32'hbc7d29e9} /* (16, 8, 29) {real, imag} */,
  {32'h3e55f090, 32'hbf99b92f} /* (16, 8, 28) {real, imag} */,
  {32'hbf6fa4e3, 32'h3f4577bc} /* (16, 8, 27) {real, imag} */,
  {32'hbf9237ed, 32'hbe4bd2b7} /* (16, 8, 26) {real, imag} */,
  {32'hbd6829ce, 32'h3ede5ff7} /* (16, 8, 25) {real, imag} */,
  {32'h3f94c44f, 32'h3e965870} /* (16, 8, 24) {real, imag} */,
  {32'h3e8498a5, 32'hbfb11e4b} /* (16, 8, 23) {real, imag} */,
  {32'hbfa06117, 32'h3fa4b259} /* (16, 8, 22) {real, imag} */,
  {32'hbf6f1c88, 32'hbf8a8d23} /* (16, 8, 21) {real, imag} */,
  {32'h3f8a07f2, 32'hbf1ce123} /* (16, 8, 20) {real, imag} */,
  {32'h3f0ac0c5, 32'h3f990185} /* (16, 8, 19) {real, imag} */,
  {32'h3cdbb781, 32'hc01d6e72} /* (16, 8, 18) {real, imag} */,
  {32'h3fe00bf8, 32'h3f5278a4} /* (16, 8, 17) {real, imag} */,
  {32'hbfdf913d, 32'h3de7a005} /* (16, 8, 16) {real, imag} */,
  {32'h3f11a36d, 32'h3de90e06} /* (16, 8, 15) {real, imag} */,
  {32'h3e5ef322, 32'h3ddc3574} /* (16, 8, 14) {real, imag} */,
  {32'hbfc262b1, 32'h3ea6cd81} /* (16, 8, 13) {real, imag} */,
  {32'h3fc8a03b, 32'h3f111809} /* (16, 8, 12) {real, imag} */,
  {32'hbeff02f7, 32'hbf596a31} /* (16, 8, 11) {real, imag} */,
  {32'hbf9f88d6, 32'h3f9138b6} /* (16, 8, 10) {real, imag} */,
  {32'hbeacce7e, 32'h40434bf3} /* (16, 8, 9) {real, imag} */,
  {32'hc0000c69, 32'hbea0ee95} /* (16, 8, 8) {real, imag} */,
  {32'h3f3c5b74, 32'h3f4af19e} /* (16, 8, 7) {real, imag} */,
  {32'h3fc9ce86, 32'hc0031045} /* (16, 8, 6) {real, imag} */,
  {32'h3fdc629e, 32'hbfe46f04} /* (16, 8, 5) {real, imag} */,
  {32'hbf7c276f, 32'hbff3e754} /* (16, 8, 4) {real, imag} */,
  {32'hbfcc42ee, 32'h3f929e8a} /* (16, 8, 3) {real, imag} */,
  {32'hbf10addb, 32'h3fa6f36b} /* (16, 8, 2) {real, imag} */,
  {32'hbf635952, 32'h3fdaae1f} /* (16, 8, 1) {real, imag} */,
  {32'hbf07da02, 32'h3e911e1d} /* (16, 8, 0) {real, imag} */,
  {32'hbeaf3902, 32'hbf5bda08} /* (16, 7, 31) {real, imag} */,
  {32'hbd3d9cee, 32'h3f3faccc} /* (16, 7, 30) {real, imag} */,
  {32'hbf12fafb, 32'h3f244ca8} /* (16, 7, 29) {real, imag} */,
  {32'hbf1e30fa, 32'hbe222650} /* (16, 7, 28) {real, imag} */,
  {32'h3ed2e4b7, 32'h3f0e05b9} /* (16, 7, 27) {real, imag} */,
  {32'h3f57a354, 32'hbf0f18cb} /* (16, 7, 26) {real, imag} */,
  {32'hbfacf73b, 32'h3f5a8376} /* (16, 7, 25) {real, imag} */,
  {32'hbf0b06e4, 32'h3d3d12ea} /* (16, 7, 24) {real, imag} */,
  {32'h3f10fbc7, 32'hbcff5002} /* (16, 7, 23) {real, imag} */,
  {32'hc00c818c, 32'hbfbb9fed} /* (16, 7, 22) {real, imag} */,
  {32'h3fa05403, 32'hbe04a6a4} /* (16, 7, 21) {real, imag} */,
  {32'hbf828ab0, 32'hbf5bd0e2} /* (16, 7, 20) {real, imag} */,
  {32'hbef78e8e, 32'hbf20c077} /* (16, 7, 19) {real, imag} */,
  {32'h3d91088c, 32'h3e61c08f} /* (16, 7, 18) {real, imag} */,
  {32'hbee6c9b2, 32'hbf739b92} /* (16, 7, 17) {real, imag} */,
  {32'hbf519b41, 32'h3f85553d} /* (16, 7, 16) {real, imag} */,
  {32'h3e44ead7, 32'hbf1d336d} /* (16, 7, 15) {real, imag} */,
  {32'h3f582973, 32'h3f87b15c} /* (16, 7, 14) {real, imag} */,
  {32'hbf913b57, 32'h3f53d509} /* (16, 7, 13) {real, imag} */,
  {32'hbded0ce0, 32'h3fd32062} /* (16, 7, 12) {real, imag} */,
  {32'h3ec24501, 32'h3bf18c38} /* (16, 7, 11) {real, imag} */,
  {32'hbee3aeba, 32'hbf116c92} /* (16, 7, 10) {real, imag} */,
  {32'hbe3c101f, 32'hc0021f4e} /* (16, 7, 9) {real, imag} */,
  {32'h3eb54fb1, 32'hbf1e0512} /* (16, 7, 8) {real, imag} */,
  {32'hbff6351c, 32'hbe1c00cb} /* (16, 7, 7) {real, imag} */,
  {32'h3dbdd7d8, 32'h3ee367c5} /* (16, 7, 6) {real, imag} */,
  {32'hbf33a5f8, 32'h400744f6} /* (16, 7, 5) {real, imag} */,
  {32'hbfc02ff3, 32'h3f857430} /* (16, 7, 4) {real, imag} */,
  {32'hbe54c55d, 32'h3fc01631} /* (16, 7, 3) {real, imag} */,
  {32'hbf5b38ad, 32'h3da1c9a6} /* (16, 7, 2) {real, imag} */,
  {32'h3f64a5b4, 32'hbca52d7e} /* (16, 7, 1) {real, imag} */,
  {32'h3e889c94, 32'h3fb3389b} /* (16, 7, 0) {real, imag} */,
  {32'hbf59cb6d, 32'hbef90db4} /* (16, 6, 31) {real, imag} */,
  {32'h3f122d10, 32'h3f84d518} /* (16, 6, 30) {real, imag} */,
  {32'hbf22027e, 32'h3fcc7e2f} /* (16, 6, 29) {real, imag} */,
  {32'hbfbc623b, 32'h3d21a9f1} /* (16, 6, 28) {real, imag} */,
  {32'hbf8dbcd9, 32'h3fa456ce} /* (16, 6, 27) {real, imag} */,
  {32'hbf83dd4e, 32'hbd1a5586} /* (16, 6, 26) {real, imag} */,
  {32'hbf9ca9cf, 32'hbfa16415} /* (16, 6, 25) {real, imag} */,
  {32'h3f696e5e, 32'h3e4ff717} /* (16, 6, 24) {real, imag} */,
  {32'hbf7149d7, 32'hbe1abc02} /* (16, 6, 23) {real, imag} */,
  {32'h3ed844fa, 32'hbfc98ba4} /* (16, 6, 22) {real, imag} */,
  {32'h3f57f53f, 32'hbf2a9e50} /* (16, 6, 21) {real, imag} */,
  {32'h3fec7647, 32'h3f74a6a8} /* (16, 6, 20) {real, imag} */,
  {32'h3fb9193e, 32'hbfb9509b} /* (16, 6, 19) {real, imag} */,
  {32'hbf1f8a48, 32'hbf9a8703} /* (16, 6, 18) {real, imag} */,
  {32'hbf0fa3e0, 32'hbfd36074} /* (16, 6, 17) {real, imag} */,
  {32'hbdb1c068, 32'hbbedd744} /* (16, 6, 16) {real, imag} */,
  {32'h3f9d623a, 32'h3f55309a} /* (16, 6, 15) {real, imag} */,
  {32'h3ee56818, 32'h3eb1d60f} /* (16, 6, 14) {real, imag} */,
  {32'hbd1f232b, 32'hbed8e24a} /* (16, 6, 13) {real, imag} */,
  {32'h3f4ef2b8, 32'hbe292d47} /* (16, 6, 12) {real, imag} */,
  {32'h3fbfab7d, 32'hc01f6483} /* (16, 6, 11) {real, imag} */,
  {32'hbfb329fa, 32'h3daee7f1} /* (16, 6, 10) {real, imag} */,
  {32'h3ed21950, 32'hbf9411a9} /* (16, 6, 9) {real, imag} */,
  {32'h3ffcc9e2, 32'hbe0b5949} /* (16, 6, 8) {real, imag} */,
  {32'hbf397af8, 32'h3f99571c} /* (16, 6, 7) {real, imag} */,
  {32'h3ed10fe4, 32'hbf3be682} /* (16, 6, 6) {real, imag} */,
  {32'h3fd081ff, 32'h3ee9ccf7} /* (16, 6, 5) {real, imag} */,
  {32'h3f7750d5, 32'h3d2a4bbb} /* (16, 6, 4) {real, imag} */,
  {32'hbdf31a93, 32'h3f91f9aa} /* (16, 6, 3) {real, imag} */,
  {32'hbf1c9518, 32'hbf169f70} /* (16, 6, 2) {real, imag} */,
  {32'hbfad9650, 32'hc002aa2f} /* (16, 6, 1) {real, imag} */,
  {32'h3de8cc59, 32'hbfa96b66} /* (16, 6, 0) {real, imag} */,
  {32'hbe996a02, 32'hbf37bd09} /* (16, 5, 31) {real, imag} */,
  {32'hbe8b8da7, 32'h3ff519b5} /* (16, 5, 30) {real, imag} */,
  {32'h3fb05d62, 32'hbc2fbe81} /* (16, 5, 29) {real, imag} */,
  {32'h3ee8e4ae, 32'h3f616ff8} /* (16, 5, 28) {real, imag} */,
  {32'hbf126670, 32'h3f7a3950} /* (16, 5, 27) {real, imag} */,
  {32'hbf2ce2ec, 32'h3f6939ec} /* (16, 5, 26) {real, imag} */,
  {32'hbcb89da4, 32'h3df2f694} /* (16, 5, 25) {real, imag} */,
  {32'h3f68d353, 32'h3e8e72b3} /* (16, 5, 24) {real, imag} */,
  {32'h3d18ffd3, 32'hbf28f975} /* (16, 5, 23) {real, imag} */,
  {32'h3f0c7772, 32'h3d3c0f2d} /* (16, 5, 22) {real, imag} */,
  {32'h3f12d504, 32'hbfb83f29} /* (16, 5, 21) {real, imag} */,
  {32'hbfed6845, 32'hbe632879} /* (16, 5, 20) {real, imag} */,
  {32'h3e8dcbb7, 32'hbffa15c4} /* (16, 5, 19) {real, imag} */,
  {32'hbfa13402, 32'hbe6a7978} /* (16, 5, 18) {real, imag} */,
  {32'hbf435afa, 32'h3db668c5} /* (16, 5, 17) {real, imag} */,
  {32'h3d83466c, 32'hbf173c09} /* (16, 5, 16) {real, imag} */,
  {32'h3eb7f0ec, 32'h3fe7952a} /* (16, 5, 15) {real, imag} */,
  {32'h3f3de5ed, 32'h3f213088} /* (16, 5, 14) {real, imag} */,
  {32'hbe0a05a2, 32'h3ecf484c} /* (16, 5, 13) {real, imag} */,
  {32'hbf3b8062, 32'hbee30373} /* (16, 5, 12) {real, imag} */,
  {32'h3fdb8b36, 32'h3f196083} /* (16, 5, 11) {real, imag} */,
  {32'h3eda3d67, 32'h3ca0770b} /* (16, 5, 10) {real, imag} */,
  {32'hbf496480, 32'h3f721a1d} /* (16, 5, 9) {real, imag} */,
  {32'h3fbe34bf, 32'hbeef9a31} /* (16, 5, 8) {real, imag} */,
  {32'hbede1e2d, 32'h3f0f5d6d} /* (16, 5, 7) {real, imag} */,
  {32'hbe002223, 32'h3f1c6d6c} /* (16, 5, 6) {real, imag} */,
  {32'hbe4c8dd4, 32'h3ffffa16} /* (16, 5, 5) {real, imag} */,
  {32'hbe8b0c93, 32'hbfb7b6f8} /* (16, 5, 4) {real, imag} */,
  {32'h3f58591d, 32'h3fb66cfc} /* (16, 5, 3) {real, imag} */,
  {32'hbf9effce, 32'h3e92957a} /* (16, 5, 2) {real, imag} */,
  {32'hbf0f97f1, 32'hbf29b130} /* (16, 5, 1) {real, imag} */,
  {32'hbe6f81a5, 32'hbfa42237} /* (16, 5, 0) {real, imag} */,
  {32'h3f62657b, 32'hc00ccab8} /* (16, 4, 31) {real, imag} */,
  {32'hbf37eab3, 32'h3f9fc1a7} /* (16, 4, 30) {real, imag} */,
  {32'hbd24cc3c, 32'h3e9964f9} /* (16, 4, 29) {real, imag} */,
  {32'hbff35c29, 32'h3e8c48fe} /* (16, 4, 28) {real, imag} */,
  {32'hbedcdd58, 32'h3fc930a0} /* (16, 4, 27) {real, imag} */,
  {32'h3f9c91d7, 32'hbdb4fedf} /* (16, 4, 26) {real, imag} */,
  {32'h3fb5c7db, 32'hbf83143f} /* (16, 4, 25) {real, imag} */,
  {32'hbf8b7d9e, 32'h3e8b5ff8} /* (16, 4, 24) {real, imag} */,
  {32'h400131f8, 32'hbe43553a} /* (16, 4, 23) {real, imag} */,
  {32'h3ec52fde, 32'h3f529033} /* (16, 4, 22) {real, imag} */,
  {32'h3f146252, 32'h3f2715dc} /* (16, 4, 21) {real, imag} */,
  {32'h3eb44a3e, 32'hbfefe21c} /* (16, 4, 20) {real, imag} */,
  {32'hbeb046ed, 32'hbf2e77eb} /* (16, 4, 19) {real, imag} */,
  {32'hbfce5079, 32'hbe9cfda4} /* (16, 4, 18) {real, imag} */,
  {32'hc0194ae6, 32'h40223e34} /* (16, 4, 17) {real, imag} */,
  {32'hbde23ff9, 32'hbf8d1be8} /* (16, 4, 16) {real, imag} */,
  {32'hbfb36337, 32'hbf655fbe} /* (16, 4, 15) {real, imag} */,
  {32'h3f9f3443, 32'hbed74d5d} /* (16, 4, 14) {real, imag} */,
  {32'hbf42041d, 32'h3f9ee31f} /* (16, 4, 13) {real, imag} */,
  {32'h3f87a042, 32'hbf6b0687} /* (16, 4, 12) {real, imag} */,
  {32'hbf9fd026, 32'hbfdeca42} /* (16, 4, 11) {real, imag} */,
  {32'h3f8b15fd, 32'h403b67a1} /* (16, 4, 10) {real, imag} */,
  {32'h3f561869, 32'h3fa3e169} /* (16, 4, 9) {real, imag} */,
  {32'h3f366194, 32'hbf6babfc} /* (16, 4, 8) {real, imag} */,
  {32'hbf99b0c8, 32'h3f2da2aa} /* (16, 4, 7) {real, imag} */,
  {32'hbfb8e8a7, 32'h3f35d13c} /* (16, 4, 6) {real, imag} */,
  {32'h3f08d3a3, 32'h3f8bd079} /* (16, 4, 5) {real, imag} */,
  {32'h3f41050e, 32'hc00ab187} /* (16, 4, 4) {real, imag} */,
  {32'h3f86a0cb, 32'hbe7e349c} /* (16, 4, 3) {real, imag} */,
  {32'hbe7d79b0, 32'h40013560} /* (16, 4, 2) {real, imag} */,
  {32'h3bf4c2f0, 32'hbf31504d} /* (16, 4, 1) {real, imag} */,
  {32'hbf51b94f, 32'hbf2880f1} /* (16, 4, 0) {real, imag} */,
  {32'hbff2a3d2, 32'h3f92f748} /* (16, 3, 31) {real, imag} */,
  {32'hbef971f5, 32'hbf1df3d1} /* (16, 3, 30) {real, imag} */,
  {32'hbfbd2d67, 32'h3ffadf08} /* (16, 3, 29) {real, imag} */,
  {32'h3fc10dd1, 32'h3f0cb92e} /* (16, 3, 28) {real, imag} */,
  {32'hbe8f2f86, 32'hbf79be9c} /* (16, 3, 27) {real, imag} */,
  {32'h3f6c2cbc, 32'hbf2ad22b} /* (16, 3, 26) {real, imag} */,
  {32'hbfb8a978, 32'hbf499372} /* (16, 3, 25) {real, imag} */,
  {32'hbf020d27, 32'hbfb076a9} /* (16, 3, 24) {real, imag} */,
  {32'hbe87c95e, 32'hbf2b1257} /* (16, 3, 23) {real, imag} */,
  {32'h3f622a09, 32'h3d3c5058} /* (16, 3, 22) {real, imag} */,
  {32'hbfa0bb84, 32'h3ef4999f} /* (16, 3, 21) {real, imag} */,
  {32'hbf3f0dbc, 32'h3f378b65} /* (16, 3, 20) {real, imag} */,
  {32'h3f5140b0, 32'hbee1fa37} /* (16, 3, 19) {real, imag} */,
  {32'hbfe59f7f, 32'hbe5ac2ff} /* (16, 3, 18) {real, imag} */,
  {32'h3fc56e5b, 32'hbf672ccd} /* (16, 3, 17) {real, imag} */,
  {32'hbdd8b902, 32'h3eef3335} /* (16, 3, 16) {real, imag} */,
  {32'hbf4a6b10, 32'h3f871365} /* (16, 3, 15) {real, imag} */,
  {32'h3f358d66, 32'hbfd15669} /* (16, 3, 14) {real, imag} */,
  {32'hbf0c38e3, 32'hc02954ad} /* (16, 3, 13) {real, imag} */,
  {32'h3ddae87b, 32'hbf528286} /* (16, 3, 12) {real, imag} */,
  {32'h40090b0d, 32'h40200d2a} /* (16, 3, 11) {real, imag} */,
  {32'h3fa47ecf, 32'hbe32ea78} /* (16, 3, 10) {real, imag} */,
  {32'hbf7923c5, 32'hbf85d18f} /* (16, 3, 9) {real, imag} */,
  {32'h3f5816a6, 32'hbe585c10} /* (16, 3, 8) {real, imag} */,
  {32'h3e587921, 32'h3feab37c} /* (16, 3, 7) {real, imag} */,
  {32'hbecbf76c, 32'hbf18531a} /* (16, 3, 6) {real, imag} */,
  {32'h3f7ed4e4, 32'h3f0ace45} /* (16, 3, 5) {real, imag} */,
  {32'hbe41a8a7, 32'hbf02d235} /* (16, 3, 4) {real, imag} */,
  {32'hbf8fdbf5, 32'h3e84fe8a} /* (16, 3, 3) {real, imag} */,
  {32'h3e736e70, 32'hbfbf95e1} /* (16, 3, 2) {real, imag} */,
  {32'hbfe5fc66, 32'h3f949405} /* (16, 3, 1) {real, imag} */,
  {32'hbeaad7d0, 32'hbd3c728b} /* (16, 3, 0) {real, imag} */,
  {32'h3d12906e, 32'hbec6ecb4} /* (16, 2, 31) {real, imag} */,
  {32'h3f6a5e85, 32'h3eac98cc} /* (16, 2, 30) {real, imag} */,
  {32'hbf26e2f7, 32'hbf34faf3} /* (16, 2, 29) {real, imag} */,
  {32'h3f21cbc9, 32'hbeb064ce} /* (16, 2, 28) {real, imag} */,
  {32'hbf686d9d, 32'hbaf5929e} /* (16, 2, 27) {real, imag} */,
  {32'h3e9c19ad, 32'h3eefb723} /* (16, 2, 26) {real, imag} */,
  {32'hbb8d60a1, 32'hbf6c511c} /* (16, 2, 25) {real, imag} */,
  {32'h3ef307f9, 32'h3f974d22} /* (16, 2, 24) {real, imag} */,
  {32'h3fbcb5a0, 32'hbf52fc27} /* (16, 2, 23) {real, imag} */,
  {32'hc0362897, 32'h3f40f171} /* (16, 2, 22) {real, imag} */,
  {32'h3f146084, 32'h3e6db50d} /* (16, 2, 21) {real, imag} */,
  {32'hbe2c862a, 32'h3ea53cee} /* (16, 2, 20) {real, imag} */,
  {32'hc01d1d22, 32'h3fee0490} /* (16, 2, 19) {real, imag} */,
  {32'hbd1282cb, 32'hbf120c33} /* (16, 2, 18) {real, imag} */,
  {32'hbe948e26, 32'h3fe0646f} /* (16, 2, 17) {real, imag} */,
  {32'h3d856b61, 32'hbe5ecb6d} /* (16, 2, 16) {real, imag} */,
  {32'hbf7e096c, 32'hbf30cb2a} /* (16, 2, 15) {real, imag} */,
  {32'hbef9e34a, 32'hbef09ccb} /* (16, 2, 14) {real, imag} */,
  {32'hbf80fd51, 32'hbe6cd2d9} /* (16, 2, 13) {real, imag} */,
  {32'hbd78f5ac, 32'hbf8756a0} /* (16, 2, 12) {real, imag} */,
  {32'h401243cc, 32'h3f72144c} /* (16, 2, 11) {real, imag} */,
  {32'h3fedb83e, 32'h3e8b766b} /* (16, 2, 10) {real, imag} */,
  {32'hbd0fcb66, 32'h3e742233} /* (16, 2, 9) {real, imag} */,
  {32'hbf5d6854, 32'h3f85e826} /* (16, 2, 8) {real, imag} */,
  {32'hbebaca04, 32'h3d818fc8} /* (16, 2, 7) {real, imag} */,
  {32'h3ed49852, 32'h3fb9dd2e} /* (16, 2, 6) {real, imag} */,
  {32'h3fb6a836, 32'hbe811004} /* (16, 2, 5) {real, imag} */,
  {32'hbef0dd36, 32'h3fb30aaf} /* (16, 2, 4) {real, imag} */,
  {32'hbf2b66ba, 32'hbf55954d} /* (16, 2, 3) {real, imag} */,
  {32'hbf04ab9f, 32'h3f30b39f} /* (16, 2, 2) {real, imag} */,
  {32'hbfc6d9e9, 32'h3f12a3af} /* (16, 2, 1) {real, imag} */,
  {32'h3d8ead56, 32'h3e8dc88d} /* (16, 2, 0) {real, imag} */,
  {32'h3f2a469f, 32'h3f9e0196} /* (16, 1, 31) {real, imag} */,
  {32'hbf1b10cc, 32'h3fbd0080} /* (16, 1, 30) {real, imag} */,
  {32'h3ecf393a, 32'h3fb96afd} /* (16, 1, 29) {real, imag} */,
  {32'h3d9816f6, 32'hbd9f17ba} /* (16, 1, 28) {real, imag} */,
  {32'hbe043dbf, 32'hbfadfb23} /* (16, 1, 27) {real, imag} */,
  {32'h3f15915b, 32'h3f75e42e} /* (16, 1, 26) {real, imag} */,
  {32'hbe0e1c56, 32'hbdb79849} /* (16, 1, 25) {real, imag} */,
  {32'hbe50a3a8, 32'hbf81fd71} /* (16, 1, 24) {real, imag} */,
  {32'hbf2da598, 32'hbe7eac86} /* (16, 1, 23) {real, imag} */,
  {32'hbf74bebd, 32'h3f20016f} /* (16, 1, 22) {real, imag} */,
  {32'hbf4e0358, 32'h3e66959a} /* (16, 1, 21) {real, imag} */,
  {32'hc0138540, 32'hbde08795} /* (16, 1, 20) {real, imag} */,
  {32'h3f5416e0, 32'hbf8d26e7} /* (16, 1, 19) {real, imag} */,
  {32'h3f119517, 32'h3f05c3e8} /* (16, 1, 18) {real, imag} */,
  {32'hbdb92454, 32'hbce68a89} /* (16, 1, 17) {real, imag} */,
  {32'h3e00f0fc, 32'h3f9090d9} /* (16, 1, 16) {real, imag} */,
  {32'h3d9616b9, 32'h3be1ba61} /* (16, 1, 15) {real, imag} */,
  {32'hbd4127f2, 32'h3eb2458b} /* (16, 1, 14) {real, imag} */,
  {32'h3eef3160, 32'h3fd9192c} /* (16, 1, 13) {real, imag} */,
  {32'h3e51cb50, 32'hbf6e6ff2} /* (16, 1, 12) {real, imag} */,
  {32'hbeee653d, 32'hc00009f7} /* (16, 1, 11) {real, imag} */,
  {32'hbfeeb48c, 32'h3f16f076} /* (16, 1, 10) {real, imag} */,
  {32'h3f8de299, 32'hbfbcac11} /* (16, 1, 9) {real, imag} */,
  {32'h3dd9cf7f, 32'hbdb04dc8} /* (16, 1, 8) {real, imag} */,
  {32'hbe9f1a5d, 32'hbec72279} /* (16, 1, 7) {real, imag} */,
  {32'h3e8a5470, 32'h3edf3643} /* (16, 1, 6) {real, imag} */,
  {32'h3fad2841, 32'hbec7d2bb} /* (16, 1, 5) {real, imag} */,
  {32'hbfe4a6fe, 32'hbf411c83} /* (16, 1, 4) {real, imag} */,
  {32'hbedb507a, 32'hbf91ea45} /* (16, 1, 3) {real, imag} */,
  {32'hbf525e6a, 32'h3fa5852b} /* (16, 1, 2) {real, imag} */,
  {32'hbe4f5ee5, 32'hbafde438} /* (16, 1, 1) {real, imag} */,
  {32'h3f805e94, 32'hbea769a9} /* (16, 1, 0) {real, imag} */,
  {32'h3f1dec83, 32'h3e771f61} /* (16, 0, 31) {real, imag} */,
  {32'hbd68e28e, 32'hbf257369} /* (16, 0, 30) {real, imag} */,
  {32'h3f61b1ab, 32'h3e0375bb} /* (16, 0, 29) {real, imag} */,
  {32'hbed3bcef, 32'h3eebffd5} /* (16, 0, 28) {real, imag} */,
  {32'hbfbae4d7, 32'hbe88cff7} /* (16, 0, 27) {real, imag} */,
  {32'h3e401683, 32'hbf385c93} /* (16, 0, 26) {real, imag} */,
  {32'hbf366f77, 32'hbfb0063a} /* (16, 0, 25) {real, imag} */,
  {32'h3ea38213, 32'hbf2ed7d5} /* (16, 0, 24) {real, imag} */,
  {32'hc0287cf1, 32'hbf6a1d22} /* (16, 0, 23) {real, imag} */,
  {32'hbf08aea8, 32'hbfca6fea} /* (16, 0, 22) {real, imag} */,
  {32'hbe6089b1, 32'h3f527de2} /* (16, 0, 21) {real, imag} */,
  {32'h3ee9f928, 32'hbf6a0e75} /* (16, 0, 20) {real, imag} */,
  {32'h3de2394e, 32'h3f4fbafd} /* (16, 0, 19) {real, imag} */,
  {32'hbfb26897, 32'hbfcd7b80} /* (16, 0, 18) {real, imag} */,
  {32'h3f276ccd, 32'h3eb1d5e6} /* (16, 0, 17) {real, imag} */,
  {32'hbf6ee06b, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3f276ccd, 32'hbeb1d5e6} /* (16, 0, 15) {real, imag} */,
  {32'hbfb26897, 32'h3fcd7b80} /* (16, 0, 14) {real, imag} */,
  {32'h3de2394e, 32'hbf4fbafd} /* (16, 0, 13) {real, imag} */,
  {32'h3ee9f928, 32'h3f6a0e75} /* (16, 0, 12) {real, imag} */,
  {32'hbe6089b1, 32'hbf527de2} /* (16, 0, 11) {real, imag} */,
  {32'hbf08aea8, 32'h3fca6fea} /* (16, 0, 10) {real, imag} */,
  {32'hc0287cf1, 32'h3f6a1d22} /* (16, 0, 9) {real, imag} */,
  {32'h3ea38213, 32'h3f2ed7d5} /* (16, 0, 8) {real, imag} */,
  {32'hbf366f77, 32'h3fb0063a} /* (16, 0, 7) {real, imag} */,
  {32'h3e401683, 32'h3f385c93} /* (16, 0, 6) {real, imag} */,
  {32'hbfbae4d7, 32'h3e88cff7} /* (16, 0, 5) {real, imag} */,
  {32'hbed3bcef, 32'hbeebffd5} /* (16, 0, 4) {real, imag} */,
  {32'h3f61b1ab, 32'hbe0375bb} /* (16, 0, 3) {real, imag} */,
  {32'hbd68e28e, 32'h3f257369} /* (16, 0, 2) {real, imag} */,
  {32'h3f1dec83, 32'hbe771f61} /* (16, 0, 1) {real, imag} */,
  {32'hbbc48c29, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h3f8ddb01, 32'hbf76c711} /* (15, 31, 31) {real, imag} */,
  {32'hbffb9a3d, 32'h3f68dc30} /* (15, 31, 30) {real, imag} */,
  {32'hbf958e79, 32'h4072430c} /* (15, 31, 29) {real, imag} */,
  {32'h3f3d8caa, 32'h3f731b47} /* (15, 31, 28) {real, imag} */,
  {32'hc037eb6a, 32'h3fd4ba44} /* (15, 31, 27) {real, imag} */,
  {32'hbe388719, 32'h3fcae9d8} /* (15, 31, 26) {real, imag} */,
  {32'h3f741f78, 32'hbf2199f2} /* (15, 31, 25) {real, imag} */,
  {32'hbf86353b, 32'hbea1bd36} /* (15, 31, 24) {real, imag} */,
  {32'hbf52c46a, 32'h3fcfced6} /* (15, 31, 23) {real, imag} */,
  {32'h3f89260e, 32'h3fef1c15} /* (15, 31, 22) {real, imag} */,
  {32'hbe542699, 32'hbfc0363a} /* (15, 31, 21) {real, imag} */,
  {32'h3f666742, 32'hbf72c5a6} /* (15, 31, 20) {real, imag} */,
  {32'hbedaebba, 32'h3fbc585f} /* (15, 31, 19) {real, imag} */,
  {32'hbf8f4a50, 32'hbf43e234} /* (15, 31, 18) {real, imag} */,
  {32'hbf4d1485, 32'h3f9f1b26} /* (15, 31, 17) {real, imag} */,
  {32'h3cdf7016, 32'h3d014a39} /* (15, 31, 16) {real, imag} */,
  {32'h3fe00f12, 32'h3feaac91} /* (15, 31, 15) {real, imag} */,
  {32'hbf2b7ec9, 32'hbe409ea2} /* (15, 31, 14) {real, imag} */,
  {32'h3e8035e9, 32'h3e3163cc} /* (15, 31, 13) {real, imag} */,
  {32'h40580e32, 32'h3e3730f8} /* (15, 31, 12) {real, imag} */,
  {32'h3fb238be, 32'hbec56bc5} /* (15, 31, 11) {real, imag} */,
  {32'h3e00cf5d, 32'h3e4ac89a} /* (15, 31, 10) {real, imag} */,
  {32'h3f84c5ff, 32'hc00aed9e} /* (15, 31, 9) {real, imag} */,
  {32'hbe417e70, 32'hc00d11be} /* (15, 31, 8) {real, imag} */,
  {32'h4018d82f, 32'h3ff9250a} /* (15, 31, 7) {real, imag} */,
  {32'hbf00bcab, 32'h4014775c} /* (15, 31, 6) {real, imag} */,
  {32'h3f903d07, 32'hbfdd53cb} /* (15, 31, 5) {real, imag} */,
  {32'h3d36aaff, 32'h3fa0dd99} /* (15, 31, 4) {real, imag} */,
  {32'h3c82cef3, 32'h3f56007c} /* (15, 31, 3) {real, imag} */,
  {32'hbed99beb, 32'hc00e31dd} /* (15, 31, 2) {real, imag} */,
  {32'h400e6349, 32'h3fd5ef51} /* (15, 31, 1) {real, imag} */,
  {32'h3d06068c, 32'hbf5f05f7} /* (15, 31, 0) {real, imag} */,
  {32'h3d8be3a9, 32'h3f8dfaa4} /* (15, 30, 31) {real, imag} */,
  {32'h402f9dc4, 32'hbfc8d9aa} /* (15, 30, 30) {real, imag} */,
  {32'hbf53af39, 32'hbf33baf4} /* (15, 30, 29) {real, imag} */,
  {32'h3eeeb3be, 32'hbf9b3c8f} /* (15, 30, 28) {real, imag} */,
  {32'hbfb55a5b, 32'hbf040791} /* (15, 30, 27) {real, imag} */,
  {32'h3f078ceb, 32'hbf4321e0} /* (15, 30, 26) {real, imag} */,
  {32'hbfa83419, 32'h3f38f3f2} /* (15, 30, 25) {real, imag} */,
  {32'h3faaba90, 32'hbe75a233} /* (15, 30, 24) {real, imag} */,
  {32'hbf2ab9e5, 32'h3fb36e2b} /* (15, 30, 23) {real, imag} */,
  {32'h3fb18439, 32'h3f1c9b37} /* (15, 30, 22) {real, imag} */,
  {32'h3f57609d, 32'hbf7389f9} /* (15, 30, 21) {real, imag} */,
  {32'h3f362f52, 32'h3f35a23b} /* (15, 30, 20) {real, imag} */,
  {32'hbf07238d, 32'hbe66084d} /* (15, 30, 19) {real, imag} */,
  {32'hbfca0610, 32'h3fa8a7d7} /* (15, 30, 18) {real, imag} */,
  {32'h3f80e86e, 32'hbf664da0} /* (15, 30, 17) {real, imag} */,
  {32'h3f9ec299, 32'hbf54f496} /* (15, 30, 16) {real, imag} */,
  {32'hbf41319e, 32'h3fcfa97d} /* (15, 30, 15) {real, imag} */,
  {32'h3d17cee8, 32'hbf414db0} /* (15, 30, 14) {real, imag} */,
  {32'h3d98e0fb, 32'h3f3a8ce5} /* (15, 30, 13) {real, imag} */,
  {32'h3f37a9cc, 32'h3d96ca50} /* (15, 30, 12) {real, imag} */,
  {32'hc03262a3, 32'h3eca34f2} /* (15, 30, 11) {real, imag} */,
  {32'hbe6a38f4, 32'hbfe9786b} /* (15, 30, 10) {real, imag} */,
  {32'h3d014839, 32'hc03774a2} /* (15, 30, 9) {real, imag} */,
  {32'h3fe3b23a, 32'hbf4fe9fb} /* (15, 30, 8) {real, imag} */,
  {32'hbf497764, 32'h3dc10890} /* (15, 30, 7) {real, imag} */,
  {32'hbe47db9d, 32'hbf4792f0} /* (15, 30, 6) {real, imag} */,
  {32'hbfac4a4e, 32'h3e1c67c8} /* (15, 30, 5) {real, imag} */,
  {32'hbf06f112, 32'hbf18bc6b} /* (15, 30, 4) {real, imag} */,
  {32'h3fa5294a, 32'hbf98404c} /* (15, 30, 3) {real, imag} */,
  {32'h3f41915a, 32'h3d0d90fb} /* (15, 30, 2) {real, imag} */,
  {32'h3d008666, 32'h3fe280bc} /* (15, 30, 1) {real, imag} */,
  {32'hbe96e111, 32'h3f8b6b41} /* (15, 30, 0) {real, imag} */,
  {32'h3f01f624, 32'hbfb85fa7} /* (15, 29, 31) {real, imag} */,
  {32'hbe160cd1, 32'h3f8e1901} /* (15, 29, 30) {real, imag} */,
  {32'hbdb214fb, 32'hbfa5bbca} /* (15, 29, 29) {real, imag} */,
  {32'hbf88b849, 32'h3d4ead9c} /* (15, 29, 28) {real, imag} */,
  {32'h3fb9722c, 32'h3ea04591} /* (15, 29, 27) {real, imag} */,
  {32'hbf466943, 32'hbfc6b178} /* (15, 29, 26) {real, imag} */,
  {32'hbf7200f5, 32'hbfc353d9} /* (15, 29, 25) {real, imag} */,
  {32'h401ffe57, 32'h3f459a64} /* (15, 29, 24) {real, imag} */,
  {32'hbf918a82, 32'h3f56443c} /* (15, 29, 23) {real, imag} */,
  {32'hbfa71b8a, 32'hc00cd184} /* (15, 29, 22) {real, imag} */,
  {32'h3fd73834, 32'h3f233678} /* (15, 29, 21) {real, imag} */,
  {32'hbe4c385f, 32'h401217a0} /* (15, 29, 20) {real, imag} */,
  {32'h3fbf2923, 32'h3e900cd9} /* (15, 29, 19) {real, imag} */,
  {32'hbfebc910, 32'hbf6bff82} /* (15, 29, 18) {real, imag} */,
  {32'hbdbc5097, 32'h3f705e46} /* (15, 29, 17) {real, imag} */,
  {32'h3fc49285, 32'h3ec4a2d9} /* (15, 29, 16) {real, imag} */,
  {32'h3f8905be, 32'hbeb010ba} /* (15, 29, 15) {real, imag} */,
  {32'hbfcc04ae, 32'hbfad75af} /* (15, 29, 14) {real, imag} */,
  {32'h3f6f92a0, 32'h3d452245} /* (15, 29, 13) {real, imag} */,
  {32'hbf0ac1ef, 32'hbfde78db} /* (15, 29, 12) {real, imag} */,
  {32'h3fd2967c, 32'hbfec994f} /* (15, 29, 11) {real, imag} */,
  {32'hbffd21d8, 32'hbefb86be} /* (15, 29, 10) {real, imag} */,
  {32'hbff07a28, 32'h3f8ff85a} /* (15, 29, 9) {real, imag} */,
  {32'h3f204924, 32'hbed41e99} /* (15, 29, 8) {real, imag} */,
  {32'hbf2e4787, 32'h3f5b0ad4} /* (15, 29, 7) {real, imag} */,
  {32'h3f2fd084, 32'hbd944532} /* (15, 29, 6) {real, imag} */,
  {32'hbecf3196, 32'hbf237ec6} /* (15, 29, 5) {real, imag} */,
  {32'hbf3d970a, 32'h3fa28870} /* (15, 29, 4) {real, imag} */,
  {32'hbeed75e2, 32'h3fcc05f0} /* (15, 29, 3) {real, imag} */,
  {32'hbf593557, 32'h3fa9a733} /* (15, 29, 2) {real, imag} */,
  {32'h3f1370bf, 32'h3e7a4608} /* (15, 29, 1) {real, imag} */,
  {32'h3ff86cdd, 32'hbf291748} /* (15, 29, 0) {real, imag} */,
  {32'hbf887e3a, 32'h3f1c928c} /* (15, 28, 31) {real, imag} */,
  {32'h3fd7d5e3, 32'hbf5c0fe5} /* (15, 28, 30) {real, imag} */,
  {32'hbfee8894, 32'hbee65f43} /* (15, 28, 29) {real, imag} */,
  {32'hbcce5924, 32'h40086918} /* (15, 28, 28) {real, imag} */,
  {32'hc04f1b10, 32'h3df5d809} /* (15, 28, 27) {real, imag} */,
  {32'h3efa42ea, 32'h3f4e7310} /* (15, 28, 26) {real, imag} */,
  {32'hbeb60508, 32'hc01c893e} /* (15, 28, 25) {real, imag} */,
  {32'hbef5bbfa, 32'h3f920887} /* (15, 28, 24) {real, imag} */,
  {32'h3e375cc2, 32'hbf8e0b2a} /* (15, 28, 23) {real, imag} */,
  {32'h3f420e3b, 32'h3e1ef4f5} /* (15, 28, 22) {real, imag} */,
  {32'h3f57d638, 32'hbfb5d421} /* (15, 28, 21) {real, imag} */,
  {32'h3fb90d64, 32'hbcdf9e13} /* (15, 28, 20) {real, imag} */,
  {32'h3fd42cc0, 32'h3fc785a5} /* (15, 28, 19) {real, imag} */,
  {32'hbf2c4ad9, 32'h3f989797} /* (15, 28, 18) {real, imag} */,
  {32'hbe3994e5, 32'hbfaf2839} /* (15, 28, 17) {real, imag} */,
  {32'hbdc30125, 32'h3e97691a} /* (15, 28, 16) {real, imag} */,
  {32'h3f11e03d, 32'h3f424b24} /* (15, 28, 15) {real, imag} */,
  {32'h3fbae6bc, 32'h3ce2f6cd} /* (15, 28, 14) {real, imag} */,
  {32'hbe57f9db, 32'h3ebf02dd} /* (15, 28, 13) {real, imag} */,
  {32'hbf457c99, 32'h3ff9f845} /* (15, 28, 12) {real, imag} */,
  {32'hbeb64280, 32'hbd8c646c} /* (15, 28, 11) {real, imag} */,
  {32'hbfc2aab3, 32'hbf40decf} /* (15, 28, 10) {real, imag} */,
  {32'h3f87f9d4, 32'hbd901729} /* (15, 28, 9) {real, imag} */,
  {32'h3ed431f0, 32'h3faf3538} /* (15, 28, 8) {real, imag} */,
  {32'h3f21cc83, 32'hc002087f} /* (15, 28, 7) {real, imag} */,
  {32'h3f49c430, 32'h3f58a704} /* (15, 28, 6) {real, imag} */,
  {32'h3f1a1014, 32'hbf978fde} /* (15, 28, 5) {real, imag} */,
  {32'h3e809714, 32'hc004b35c} /* (15, 28, 4) {real, imag} */,
  {32'h4017a694, 32'h3f40edd3} /* (15, 28, 3) {real, imag} */,
  {32'hbf9863a5, 32'h3fb1c81a} /* (15, 28, 2) {real, imag} */,
  {32'h3df99af2, 32'hbe0264d7} /* (15, 28, 1) {real, imag} */,
  {32'h3f5dfad5, 32'hbf0d5cc3} /* (15, 28, 0) {real, imag} */,
  {32'hbfb50ba0, 32'h402ad701} /* (15, 27, 31) {real, imag} */,
  {32'h40177dd4, 32'hc016be88} /* (15, 27, 30) {real, imag} */,
  {32'h3f1d99de, 32'h3ff7fcdc} /* (15, 27, 29) {real, imag} */,
  {32'hbf6b9ae7, 32'hbf163cfd} /* (15, 27, 28) {real, imag} */,
  {32'h3f73de44, 32'h3fcca47c} /* (15, 27, 27) {real, imag} */,
  {32'hc00cae83, 32'h400cb1eb} /* (15, 27, 26) {real, imag} */,
  {32'hbf6a2747, 32'hbf8fd17a} /* (15, 27, 25) {real, imag} */,
  {32'hbf3e4940, 32'h3f937181} /* (15, 27, 24) {real, imag} */,
  {32'h3f4f7dbf, 32'h3d41ad40} /* (15, 27, 23) {real, imag} */,
  {32'h3f2d5616, 32'hbfc47db8} /* (15, 27, 22) {real, imag} */,
  {32'hc02bc89c, 32'hc03e461a} /* (15, 27, 21) {real, imag} */,
  {32'hbeaddb9d, 32'h3f140586} /* (15, 27, 20) {real, imag} */,
  {32'hbf0c3b70, 32'hbe00a1da} /* (15, 27, 19) {real, imag} */,
  {32'h3fd13e74, 32'h3f71684f} /* (15, 27, 18) {real, imag} */,
  {32'h3fea689f, 32'h3f5dc04a} /* (15, 27, 17) {real, imag} */,
  {32'h3fe0b149, 32'h3f71bfa3} /* (15, 27, 16) {real, imag} */,
  {32'h3e6bf582, 32'h3f4df6ea} /* (15, 27, 15) {real, imag} */,
  {32'h3e08f03b, 32'h3e2e9747} /* (15, 27, 14) {real, imag} */,
  {32'h3e7f7b2c, 32'hbef7a03a} /* (15, 27, 13) {real, imag} */,
  {32'hbf7b4933, 32'hbea1590d} /* (15, 27, 12) {real, imag} */,
  {32'hbf3d4e88, 32'h3e6e40f5} /* (15, 27, 11) {real, imag} */,
  {32'h3f8b239e, 32'h3fff5cee} /* (15, 27, 10) {real, imag} */,
  {32'h3c92b71e, 32'hbe5f2e0f} /* (15, 27, 9) {real, imag} */,
  {32'h3fde42bf, 32'h3f8055f7} /* (15, 27, 8) {real, imag} */,
  {32'hbe039fdb, 32'h400548e2} /* (15, 27, 7) {real, imag} */,
  {32'h3e1e3969, 32'hbfd1784c} /* (15, 27, 6) {real, imag} */,
  {32'hbfaf863a, 32'h3d924427} /* (15, 27, 5) {real, imag} */,
  {32'h3ea972c8, 32'h3fa26716} /* (15, 27, 4) {real, imag} */,
  {32'h3f0c7ed5, 32'hbf2eeb31} /* (15, 27, 3) {real, imag} */,
  {32'h3fa1ad12, 32'h3f8f1a01} /* (15, 27, 2) {real, imag} */,
  {32'hbdb27c76, 32'hbe9dbe6f} /* (15, 27, 1) {real, imag} */,
  {32'h3f562bf3, 32'h3f78089c} /* (15, 27, 0) {real, imag} */,
  {32'h3a9314cd, 32'h3f0fb2aa} /* (15, 26, 31) {real, imag} */,
  {32'hbfb3c8c8, 32'hbfd20771} /* (15, 26, 30) {real, imag} */,
  {32'h3f63f237, 32'hbe41dab4} /* (15, 26, 29) {real, imag} */,
  {32'hc0064ee7, 32'h3ef2384d} /* (15, 26, 28) {real, imag} */,
  {32'hbef49c49, 32'h3e358ec6} /* (15, 26, 27) {real, imag} */,
  {32'h3f2c3123, 32'hbe85da05} /* (15, 26, 26) {real, imag} */,
  {32'hbf89ad43, 32'hbfeb85ae} /* (15, 26, 25) {real, imag} */,
  {32'h3dfeaaf4, 32'hbf9ed0fd} /* (15, 26, 24) {real, imag} */,
  {32'h3ffee693, 32'hbf2e1f8d} /* (15, 26, 23) {real, imag} */,
  {32'hbedeca67, 32'h3dbb6b38} /* (15, 26, 22) {real, imag} */,
  {32'h3f860ee8, 32'hc00b44fa} /* (15, 26, 21) {real, imag} */,
  {32'hbfdffc9c, 32'h3fa23b60} /* (15, 26, 20) {real, imag} */,
  {32'h3e4c4615, 32'hbe51202d} /* (15, 26, 19) {real, imag} */,
  {32'hc0071b0d, 32'h400cab05} /* (15, 26, 18) {real, imag} */,
  {32'hbeb775fe, 32'hbf85b5d2} /* (15, 26, 17) {real, imag} */,
  {32'h3f299518, 32'h3f5c7930} /* (15, 26, 16) {real, imag} */,
  {32'h3f457d4a, 32'hbe9b7e1e} /* (15, 26, 15) {real, imag} */,
  {32'hbf6f4963, 32'h3e6eeda9} /* (15, 26, 14) {real, imag} */,
  {32'hc01fcdea, 32'hbdd8c48e} /* (15, 26, 13) {real, imag} */,
  {32'hc02c86ba, 32'hc0297de4} /* (15, 26, 12) {real, imag} */,
  {32'hbc1abed5, 32'hbe65ad6d} /* (15, 26, 11) {real, imag} */,
  {32'hbfc5deff, 32'hbfcb8d0d} /* (15, 26, 10) {real, imag} */,
  {32'h3e9f063c, 32'h3f8781e3} /* (15, 26, 9) {real, imag} */,
  {32'h3fa01f49, 32'hc0180b19} /* (15, 26, 8) {real, imag} */,
  {32'h3edf6d60, 32'h3f082cea} /* (15, 26, 7) {real, imag} */,
  {32'hbf873945, 32'hbe147957} /* (15, 26, 6) {real, imag} */,
  {32'h3f8e6fa3, 32'hbf0cd824} /* (15, 26, 5) {real, imag} */,
  {32'h3f450f1e, 32'hbe6ad09b} /* (15, 26, 4) {real, imag} */,
  {32'h3fb09952, 32'h3eab757c} /* (15, 26, 3) {real, imag} */,
  {32'h3e826e00, 32'h3f6fe16a} /* (15, 26, 2) {real, imag} */,
  {32'hc04f342d, 32'h3d7ba6c1} /* (15, 26, 1) {real, imag} */,
  {32'hbffb3fbf, 32'hbfda8879} /* (15, 26, 0) {real, imag} */,
  {32'h3ecdbee3, 32'hbecc4608} /* (15, 25, 31) {real, imag} */,
  {32'h3ec6a77b, 32'h3fd2f873} /* (15, 25, 30) {real, imag} */,
  {32'h3fd6b64d, 32'h3e67b80a} /* (15, 25, 29) {real, imag} */,
  {32'hbee82a0d, 32'h3f9b3534} /* (15, 25, 28) {real, imag} */,
  {32'h3e88b9d8, 32'hbf18070f} /* (15, 25, 27) {real, imag} */,
  {32'hbf860526, 32'h3f125c02} /* (15, 25, 26) {real, imag} */,
  {32'h400bc770, 32'hbfb35f9d} /* (15, 25, 25) {real, imag} */,
  {32'h3f92c3f0, 32'h3f4926af} /* (15, 25, 24) {real, imag} */,
  {32'hbf705542, 32'hc02c0172} /* (15, 25, 23) {real, imag} */,
  {32'hc013e3a1, 32'hbdc56fd8} /* (15, 25, 22) {real, imag} */,
  {32'hbfe489dc, 32'h3fd63edf} /* (15, 25, 21) {real, imag} */,
  {32'hbe8ea5ec, 32'hbfcd73c1} /* (15, 25, 20) {real, imag} */,
  {32'h40227c45, 32'hbc258bbe} /* (15, 25, 19) {real, imag} */,
  {32'hbf8bfd5b, 32'h3fadebbc} /* (15, 25, 18) {real, imag} */,
  {32'hbff48f99, 32'h3fc718d5} /* (15, 25, 17) {real, imag} */,
  {32'hbfbc8c91, 32'h40244974} /* (15, 25, 16) {real, imag} */,
  {32'hbf2f476d, 32'hbf2dbada} /* (15, 25, 15) {real, imag} */,
  {32'hc02ceffe, 32'h3fd6cee4} /* (15, 25, 14) {real, imag} */,
  {32'h3ed68818, 32'hbd21fe99} /* (15, 25, 13) {real, imag} */,
  {32'hbeed439e, 32'hbfc737d0} /* (15, 25, 12) {real, imag} */,
  {32'h3f36442e, 32'h40410c2c} /* (15, 25, 11) {real, imag} */,
  {32'h3e8c45a9, 32'hbf22ced2} /* (15, 25, 10) {real, imag} */,
  {32'hbff43708, 32'hbec7e39f} /* (15, 25, 9) {real, imag} */,
  {32'hbe94ef6f, 32'h3f89b8a1} /* (15, 25, 8) {real, imag} */,
  {32'hbfaa790d, 32'hbeba1656} /* (15, 25, 7) {real, imag} */,
  {32'hbfc190f6, 32'hbee2f3ac} /* (15, 25, 6) {real, imag} */,
  {32'hbef94953, 32'h3e6d6bef} /* (15, 25, 5) {real, imag} */,
  {32'h3fb4a9f4, 32'hbbdf28dc} /* (15, 25, 4) {real, imag} */,
  {32'h3ee2f05e, 32'hbf85d651} /* (15, 25, 3) {real, imag} */,
  {32'h3ea1e604, 32'hbf596184} /* (15, 25, 2) {real, imag} */,
  {32'hbfc3204f, 32'hbfa4f957} /* (15, 25, 1) {real, imag} */,
  {32'hc01f6bd4, 32'h3f3b728c} /* (15, 25, 0) {real, imag} */,
  {32'hbf81e573, 32'hbfeb7810} /* (15, 24, 31) {real, imag} */,
  {32'h3dacbfa6, 32'h3f8852b9} /* (15, 24, 30) {real, imag} */,
  {32'h3f997bba, 32'hbf596ac0} /* (15, 24, 29) {real, imag} */,
  {32'h3f9b990c, 32'hbf6c6c7e} /* (15, 24, 28) {real, imag} */,
  {32'hbfc32585, 32'h3fdd94dc} /* (15, 24, 27) {real, imag} */,
  {32'hbda1db43, 32'hbf9cb0d9} /* (15, 24, 26) {real, imag} */,
  {32'h3f44a863, 32'h3ff383c2} /* (15, 24, 25) {real, imag} */,
  {32'hbeb5b6a7, 32'hbe9532b8} /* (15, 24, 24) {real, imag} */,
  {32'hbf46f498, 32'hbf1193a1} /* (15, 24, 23) {real, imag} */,
  {32'h3e6f889f, 32'h3f2a291f} /* (15, 24, 22) {real, imag} */,
  {32'hbf4101d5, 32'h3f481eac} /* (15, 24, 21) {real, imag} */,
  {32'h3faf4c4a, 32'h3f3559b7} /* (15, 24, 20) {real, imag} */,
  {32'hbe81eeea, 32'h3f48b28f} /* (15, 24, 19) {real, imag} */,
  {32'h3eff5ae2, 32'hbf839c58} /* (15, 24, 18) {real, imag} */,
  {32'h3eb31995, 32'h3eec46be} /* (15, 24, 17) {real, imag} */,
  {32'h3f73193c, 32'h400b9326} /* (15, 24, 16) {real, imag} */,
  {32'hbd5881bc, 32'h4031ebc0} /* (15, 24, 15) {real, imag} */,
  {32'hbfcb798f, 32'hbff347e3} /* (15, 24, 14) {real, imag} */,
  {32'h3fcb47d4, 32'hbff0d25a} /* (15, 24, 13) {real, imag} */,
  {32'h3fb0f01d, 32'h3f83f527} /* (15, 24, 12) {real, imag} */,
  {32'h3fd13bf4, 32'h40187536} /* (15, 24, 11) {real, imag} */,
  {32'hbe04462f, 32'h3fadf115} /* (15, 24, 10) {real, imag} */,
  {32'h3e8c9591, 32'hbfd6c6ca} /* (15, 24, 9) {real, imag} */,
  {32'h3ff32954, 32'hbdd79bc1} /* (15, 24, 8) {real, imag} */,
  {32'hbefdaca4, 32'hbd6657a1} /* (15, 24, 7) {real, imag} */,
  {32'h3f106920, 32'hbe5e117a} /* (15, 24, 6) {real, imag} */,
  {32'hbd466ade, 32'h3ffc5edc} /* (15, 24, 5) {real, imag} */,
  {32'hbf993d34, 32'hc0305e31} /* (15, 24, 4) {real, imag} */,
  {32'h3e3545c2, 32'h3ea6c3cf} /* (15, 24, 3) {real, imag} */,
  {32'hbf0de9c1, 32'hbfd67364} /* (15, 24, 2) {real, imag} */,
  {32'hbf04591d, 32'h3f2f1940} /* (15, 24, 1) {real, imag} */,
  {32'h39ae2682, 32'hbf291de5} /* (15, 24, 0) {real, imag} */,
  {32'hbfac91e6, 32'h3e64c335} /* (15, 23, 31) {real, imag} */,
  {32'h400cdf2e, 32'h3f1399e3} /* (15, 23, 30) {real, imag} */,
  {32'hbf954576, 32'h3ffea266} /* (15, 23, 29) {real, imag} */,
  {32'hc01460d2, 32'hbfbd8dae} /* (15, 23, 28) {real, imag} */,
  {32'h3f820ddc, 32'h3f80daea} /* (15, 23, 27) {real, imag} */,
  {32'h3ef9e79a, 32'hbf164b81} /* (15, 23, 26) {real, imag} */,
  {32'hbefbac38, 32'h3f4394c8} /* (15, 23, 25) {real, imag} */,
  {32'h3e2bb564, 32'hbdbbd58a} /* (15, 23, 24) {real, imag} */,
  {32'h3e09f72b, 32'hbf99d682} /* (15, 23, 23) {real, imag} */,
  {32'hbfffc5f9, 32'h3fcf3ab8} /* (15, 23, 22) {real, imag} */,
  {32'hbea0c14d, 32'h3f423fdc} /* (15, 23, 21) {real, imag} */,
  {32'h3f0fbfb2, 32'hbfba5c3e} /* (15, 23, 20) {real, imag} */,
  {32'hbdb273bf, 32'h3f18759b} /* (15, 23, 19) {real, imag} */,
  {32'h3e777e6c, 32'hbf748674} /* (15, 23, 18) {real, imag} */,
  {32'h3ec706df, 32'hbf0e53b4} /* (15, 23, 17) {real, imag} */,
  {32'hbf6f2d32, 32'hbf437a3e} /* (15, 23, 16) {real, imag} */,
  {32'hbf97e7a7, 32'h3e7d59f7} /* (15, 23, 15) {real, imag} */,
  {32'hbf9d1dca, 32'h40036d7d} /* (15, 23, 14) {real, imag} */,
  {32'hc003c96d, 32'hc04c3427} /* (15, 23, 13) {real, imag} */,
  {32'hbe695686, 32'h3fcaef65} /* (15, 23, 12) {real, imag} */,
  {32'h40074aa1, 32'h3dd49621} /* (15, 23, 11) {real, imag} */,
  {32'hbf91a43b, 32'hbf9fb80c} /* (15, 23, 10) {real, imag} */,
  {32'h400eb05f, 32'h400c3925} /* (15, 23, 9) {real, imag} */,
  {32'h3f9a637e, 32'hc0946110} /* (15, 23, 8) {real, imag} */,
  {32'h3fd3698b, 32'hbe330166} /* (15, 23, 7) {real, imag} */,
  {32'hbf3caa6b, 32'hbf03922b} /* (15, 23, 6) {real, imag} */,
  {32'h3e8e58ea, 32'h3f5c1b05} /* (15, 23, 5) {real, imag} */,
  {32'hbfad7319, 32'h3f2fdcdf} /* (15, 23, 4) {real, imag} */,
  {32'hbfd8bf5d, 32'hc011b535} /* (15, 23, 3) {real, imag} */,
  {32'h3e8c05b3, 32'h3f97ac95} /* (15, 23, 2) {real, imag} */,
  {32'hbdc0a9d3, 32'h3f18a91e} /* (15, 23, 1) {real, imag} */,
  {32'hbd975491, 32'hc01e988c} /* (15, 23, 0) {real, imag} */,
  {32'hc0a168a4, 32'hbf883929} /* (15, 22, 31) {real, imag} */,
  {32'hbfa12fd6, 32'h3f31e0db} /* (15, 22, 30) {real, imag} */,
  {32'h3e9ca8c3, 32'hbef02eba} /* (15, 22, 29) {real, imag} */,
  {32'h3f79c698, 32'hc0411eb5} /* (15, 22, 28) {real, imag} */,
  {32'hbf88b499, 32'h3f84538c} /* (15, 22, 27) {real, imag} */,
  {32'h3f0a0bcf, 32'h3faec373} /* (15, 22, 26) {real, imag} */,
  {32'hbf512ff4, 32'hc007ea7c} /* (15, 22, 25) {real, imag} */,
  {32'hbeea3e6a, 32'hbf8348de} /* (15, 22, 24) {real, imag} */,
  {32'hbef600f6, 32'h3fe52368} /* (15, 22, 23) {real, imag} */,
  {32'h3fe99186, 32'h40310435} /* (15, 22, 22) {real, imag} */,
  {32'hbfd4f4f2, 32'hbe2441d1} /* (15, 22, 21) {real, imag} */,
  {32'hbfa12f6c, 32'h4023eabd} /* (15, 22, 20) {real, imag} */,
  {32'h40284891, 32'hbf3b3618} /* (15, 22, 19) {real, imag} */,
  {32'h3f76240d, 32'hbf7f2a24} /* (15, 22, 18) {real, imag} */,
  {32'hbfbfb75f, 32'h3d7629c3} /* (15, 22, 17) {real, imag} */,
  {32'h3fb67368, 32'hbefe9fe5} /* (15, 22, 16) {real, imag} */,
  {32'h4034486e, 32'hbff2f32e} /* (15, 22, 15) {real, imag} */,
  {32'h402b6fcc, 32'h3fa76968} /* (15, 22, 14) {real, imag} */,
  {32'hc021b13a, 32'h3f20677a} /* (15, 22, 13) {real, imag} */,
  {32'hc00a06f4, 32'hbedfdaab} /* (15, 22, 12) {real, imag} */,
  {32'h3fe07b5e, 32'hbe694cd0} /* (15, 22, 11) {real, imag} */,
  {32'h3f667264, 32'hbe9c89c6} /* (15, 22, 10) {real, imag} */,
  {32'hbfb06ad3, 32'h401ca688} /* (15, 22, 9) {real, imag} */,
  {32'hc0047b19, 32'h3f13302a} /* (15, 22, 8) {real, imag} */,
  {32'h3fa12691, 32'h3f58bc30} /* (15, 22, 7) {real, imag} */,
  {32'h3d7f8939, 32'h3e9c8c92} /* (15, 22, 6) {real, imag} */,
  {32'h400e594a, 32'hbfc2a71a} /* (15, 22, 5) {real, imag} */,
  {32'h3fd8f8fd, 32'h3f993279} /* (15, 22, 4) {real, imag} */,
  {32'h3f2cb1a2, 32'h3e6ed326} /* (15, 22, 3) {real, imag} */,
  {32'h3ec884a5, 32'h3fdb3285} /* (15, 22, 2) {real, imag} */,
  {32'h3e52efe2, 32'hbf9f103d} /* (15, 22, 1) {real, imag} */,
  {32'h3ec39a73, 32'hbf9c7423} /* (15, 22, 0) {real, imag} */,
  {32'hbff053de, 32'hbdbb6b1d} /* (15, 21, 31) {real, imag} */,
  {32'hbcaefe83, 32'h3fbf5582} /* (15, 21, 30) {real, imag} */,
  {32'hbf6cc9ab, 32'hbf20759c} /* (15, 21, 29) {real, imag} */,
  {32'h3faf4d94, 32'h401d0233} /* (15, 21, 28) {real, imag} */,
  {32'h3ffb5aa0, 32'hc02f3a40} /* (15, 21, 27) {real, imag} */,
  {32'hbf82b41c, 32'h3f88a972} /* (15, 21, 26) {real, imag} */,
  {32'hbfbe7fb4, 32'h4018b55c} /* (15, 21, 25) {real, imag} */,
  {32'hbee3458c, 32'h3f291b76} /* (15, 21, 24) {real, imag} */,
  {32'h3d626fb6, 32'hbf516278} /* (15, 21, 23) {real, imag} */,
  {32'hbd9d73f1, 32'h3f772093} /* (15, 21, 22) {real, imag} */,
  {32'hc00d74e8, 32'h3f95a725} /* (15, 21, 21) {real, imag} */,
  {32'hbe344454, 32'hc0464e1c} /* (15, 21, 20) {real, imag} */,
  {32'h3fa662f2, 32'h3da87792} /* (15, 21, 19) {real, imag} */,
  {32'h40005e6c, 32'hc001989c} /* (15, 21, 18) {real, imag} */,
  {32'h3fcf0d3f, 32'hbfdb3d56} /* (15, 21, 17) {real, imag} */,
  {32'hbfadd9a6, 32'hbf996283} /* (15, 21, 16) {real, imag} */,
  {32'hbfca2ee8, 32'hbefaaec1} /* (15, 21, 15) {real, imag} */,
  {32'hbe960288, 32'h3eb04bb0} /* (15, 21, 14) {real, imag} */,
  {32'hc02b4862, 32'h3f9c97b6} /* (15, 21, 13) {real, imag} */,
  {32'h4024bbe0, 32'h3f196451} /* (15, 21, 12) {real, imag} */,
  {32'hbf5e095b, 32'hc0021d7a} /* (15, 21, 11) {real, imag} */,
  {32'h3feee609, 32'h3eb97fa9} /* (15, 21, 10) {real, imag} */,
  {32'hbfaab9b3, 32'h40255688} /* (15, 21, 9) {real, imag} */,
  {32'hbe6d41ac, 32'hbf8f7d28} /* (15, 21, 8) {real, imag} */,
  {32'hbf760699, 32'h3f86e425} /* (15, 21, 7) {real, imag} */,
  {32'hc000352a, 32'hbf742695} /* (15, 21, 6) {real, imag} */,
  {32'hbf00384f, 32'hbff7324f} /* (15, 21, 5) {real, imag} */,
  {32'h3f0fa4df, 32'h3f7f3b90} /* (15, 21, 4) {real, imag} */,
  {32'h3ec8204f, 32'hbecde30e} /* (15, 21, 3) {real, imag} */,
  {32'h3f902a0e, 32'hc066eedf} /* (15, 21, 2) {real, imag} */,
  {32'h3ec2ff01, 32'hbf55f42a} /* (15, 21, 1) {real, imag} */,
  {32'h3eda960c, 32'h3f873f38} /* (15, 21, 0) {real, imag} */,
  {32'hbf99ed61, 32'h3f98864c} /* (15, 20, 31) {real, imag} */,
  {32'h3fe4087d, 32'hbf62c8d7} /* (15, 20, 30) {real, imag} */,
  {32'h3f244917, 32'hbef6b977} /* (15, 20, 29) {real, imag} */,
  {32'h3f872a91, 32'hbfdd36c0} /* (15, 20, 28) {real, imag} */,
  {32'hbeb924f8, 32'h3f7d5afe} /* (15, 20, 27) {real, imag} */,
  {32'hbe41c5be, 32'hbf2b4940} /* (15, 20, 26) {real, imag} */,
  {32'hbf4d9027, 32'hbfeeb509} /* (15, 20, 25) {real, imag} */,
  {32'h4039aa56, 32'h4012e219} /* (15, 20, 24) {real, imag} */,
  {32'h3f524c85, 32'h4021691c} /* (15, 20, 23) {real, imag} */,
  {32'h3fc1df46, 32'h3f5ce81d} /* (15, 20, 22) {real, imag} */,
  {32'h3ef3b137, 32'hbdecc12b} /* (15, 20, 21) {real, imag} */,
  {32'h3f25cec0, 32'h402c9f0f} /* (15, 20, 20) {real, imag} */,
  {32'hbee3e42a, 32'hbfee35c6} /* (15, 20, 19) {real, imag} */,
  {32'h401b688c, 32'hbf67637e} /* (15, 20, 18) {real, imag} */,
  {32'h3f6d29ab, 32'hc020eaf2} /* (15, 20, 17) {real, imag} */,
  {32'h3fd2c2d2, 32'hbf8fd482} /* (15, 20, 16) {real, imag} */,
  {32'h3f678ff0, 32'h3f11f83a} /* (15, 20, 15) {real, imag} */,
  {32'h401367d6, 32'h40148b21} /* (15, 20, 14) {real, imag} */,
  {32'h3fbba89b, 32'h3f96882b} /* (15, 20, 13) {real, imag} */,
  {32'hc09b70af, 32'hbfc4ea60} /* (15, 20, 12) {real, imag} */,
  {32'h404004c6, 32'h3f77338f} /* (15, 20, 11) {real, imag} */,
  {32'h3f82d34e, 32'h3fbdf315} /* (15, 20, 10) {real, imag} */,
  {32'hbaa6ac0e, 32'h3fdd4bca} /* (15, 20, 9) {real, imag} */,
  {32'hbfa26b4c, 32'h3db71eac} /* (15, 20, 8) {real, imag} */,
  {32'hbf9e9125, 32'h3e007c84} /* (15, 20, 7) {real, imag} */,
  {32'h3f884501, 32'h3ec3928c} /* (15, 20, 6) {real, imag} */,
  {32'hbfaf3e41, 32'h3fc9a6fb} /* (15, 20, 5) {real, imag} */,
  {32'hbf8ea24e, 32'hbfa8a217} /* (15, 20, 4) {real, imag} */,
  {32'hbf4dd065, 32'h3e640b4e} /* (15, 20, 3) {real, imag} */,
  {32'hbfa3ad86, 32'hbf3a9312} /* (15, 20, 2) {real, imag} */,
  {32'hbf97861c, 32'hbfc345d1} /* (15, 20, 1) {real, imag} */,
  {32'h3f110e34, 32'h3f5674d4} /* (15, 20, 0) {real, imag} */,
  {32'h3fd645f2, 32'hbf658874} /* (15, 19, 31) {real, imag} */,
  {32'h3f2a7329, 32'hbffda5fc} /* (15, 19, 30) {real, imag} */,
  {32'hbeb946f8, 32'hbf90983a} /* (15, 19, 29) {real, imag} */,
  {32'hbc212c0f, 32'h3fb5568d} /* (15, 19, 28) {real, imag} */,
  {32'hbe615c93, 32'h3f7ace13} /* (15, 19, 27) {real, imag} */,
  {32'h3f11e974, 32'h4037adf5} /* (15, 19, 26) {real, imag} */,
  {32'h3f618bce, 32'hbe93d20d} /* (15, 19, 25) {real, imag} */,
  {32'h3feadde4, 32'hbf2775b4} /* (15, 19, 24) {real, imag} */,
  {32'hbfc40de5, 32'hbe4a9699} /* (15, 19, 23) {real, imag} */,
  {32'hbef181ca, 32'h3f7a8113} /* (15, 19, 22) {real, imag} */,
  {32'hbf1ba8e3, 32'h3f76ce27} /* (15, 19, 21) {real, imag} */,
  {32'hbecdef43, 32'h4034e5ce} /* (15, 19, 20) {real, imag} */,
  {32'h3ea27233, 32'hbf70758c} /* (15, 19, 19) {real, imag} */,
  {32'hc0302bfe, 32'h400f83a3} /* (15, 19, 18) {real, imag} */,
  {32'h3fdd5f44, 32'h3fc63948} /* (15, 19, 17) {real, imag} */,
  {32'h3ecafbf8, 32'hbed689cd} /* (15, 19, 16) {real, imag} */,
  {32'hc0322d8d, 32'hbf929f5b} /* (15, 19, 15) {real, imag} */,
  {32'hbfb79ff7, 32'hbf859161} /* (15, 19, 14) {real, imag} */,
  {32'hc02013d6, 32'hc0808730} /* (15, 19, 13) {real, imag} */,
  {32'h3c87dfe1, 32'h3f742cdb} /* (15, 19, 12) {real, imag} */,
  {32'h3fb68174, 32'hbdde077a} /* (15, 19, 11) {real, imag} */,
  {32'h3f1d4e25, 32'h40334e00} /* (15, 19, 10) {real, imag} */,
  {32'h3f8df10b, 32'h3f411431} /* (15, 19, 9) {real, imag} */,
  {32'h3ff7eb60, 32'h3fc2207b} /* (15, 19, 8) {real, imag} */,
  {32'h3f83452d, 32'hbe97e3ec} /* (15, 19, 7) {real, imag} */,
  {32'h3ec8a7af, 32'h3e9cf5de} /* (15, 19, 6) {real, imag} */,
  {32'h3f36ecf8, 32'hbfebc7b1} /* (15, 19, 5) {real, imag} */,
  {32'hbf237542, 32'h3ff80ce8} /* (15, 19, 4) {real, imag} */,
  {32'hbf94c86a, 32'h3f420701} /* (15, 19, 3) {real, imag} */,
  {32'hbf904c04, 32'h3f209d44} /* (15, 19, 2) {real, imag} */,
  {32'h3f36b338, 32'hbec8d049} /* (15, 19, 1) {real, imag} */,
  {32'hbe6591e2, 32'h3eda4732} /* (15, 19, 0) {real, imag} */,
  {32'h3e6e6c19, 32'h3db63b47} /* (15, 18, 31) {real, imag} */,
  {32'h3fc53dac, 32'h3f1a4c90} /* (15, 18, 30) {real, imag} */,
  {32'hbe3af8c6, 32'h3e6921df} /* (15, 18, 29) {real, imag} */,
  {32'h3fc47fbe, 32'h3fc0bbb8} /* (15, 18, 28) {real, imag} */,
  {32'h3eaed351, 32'h3f014ca6} /* (15, 18, 27) {real, imag} */,
  {32'h3fffcd49, 32'h3e9e4032} /* (15, 18, 26) {real, imag} */,
  {32'h4062f1f0, 32'h3d95ce8a} /* (15, 18, 25) {real, imag} */,
  {32'h3f9748d6, 32'hbfb2ae5d} /* (15, 18, 24) {real, imag} */,
  {32'hbf124101, 32'hbe8d2981} /* (15, 18, 23) {real, imag} */,
  {32'hbe855a89, 32'hbfbaf4b0} /* (15, 18, 22) {real, imag} */,
  {32'h400fa60c, 32'h3f5a48e1} /* (15, 18, 21) {real, imag} */,
  {32'hbe45ecf3, 32'h402ba0fe} /* (15, 18, 20) {real, imag} */,
  {32'hc0741b59, 32'h4000ab8b} /* (15, 18, 19) {real, imag} */,
  {32'h3f907ed9, 32'hbed7ad48} /* (15, 18, 18) {real, imag} */,
  {32'hc06d59cb, 32'h3fd94931} /* (15, 18, 17) {real, imag} */,
  {32'hbf9409b4, 32'hbf39c46d} /* (15, 18, 16) {real, imag} */,
  {32'h3f696000, 32'h3f0864bc} /* (15, 18, 15) {real, imag} */,
  {32'hbf8de6d0, 32'h3fb0ec08} /* (15, 18, 14) {real, imag} */,
  {32'hbf14c2d6, 32'h3e3ff145} /* (15, 18, 13) {real, imag} */,
  {32'h3e8cb6a3, 32'hbdef2b7f} /* (15, 18, 12) {real, imag} */,
  {32'h3e5074d9, 32'hc02f2346} /* (15, 18, 11) {real, imag} */,
  {32'h3f266544, 32'hc0147e59} /* (15, 18, 10) {real, imag} */,
  {32'hbf9d7c03, 32'hbfb83bb6} /* (15, 18, 9) {real, imag} */,
  {32'h3dadb7df, 32'hbfaa0d35} /* (15, 18, 8) {real, imag} */,
  {32'h402b5083, 32'hc0018a88} /* (15, 18, 7) {real, imag} */,
  {32'h3f82e67a, 32'hbffe363d} /* (15, 18, 6) {real, imag} */,
  {32'h400f85f1, 32'h3fa916ad} /* (15, 18, 5) {real, imag} */,
  {32'hbdff37b3, 32'hbf858a4c} /* (15, 18, 4) {real, imag} */,
  {32'hbf717369, 32'hbf7ae1fc} /* (15, 18, 3) {real, imag} */,
  {32'h3fce0736, 32'hbf2e3983} /* (15, 18, 2) {real, imag} */,
  {32'h4002fbab, 32'h3f484660} /* (15, 18, 1) {real, imag} */,
  {32'h3c1a3ae0, 32'hbf7a54e1} /* (15, 18, 0) {real, imag} */,
  {32'hbf491c66, 32'h3fa1ebe7} /* (15, 17, 31) {real, imag} */,
  {32'h3f459058, 32'h3e05b820} /* (15, 17, 30) {real, imag} */,
  {32'h3d8fac24, 32'h3f3eedd9} /* (15, 17, 29) {real, imag} */,
  {32'hbc883c33, 32'hbf0a0189} /* (15, 17, 28) {real, imag} */,
  {32'h3d6db068, 32'hbfab368f} /* (15, 17, 27) {real, imag} */,
  {32'h3f013a85, 32'h3f1be958} /* (15, 17, 26) {real, imag} */,
  {32'hbddb760c, 32'h3f8ab28d} /* (15, 17, 25) {real, imag} */,
  {32'h3d5803e5, 32'hbfbca45a} /* (15, 17, 24) {real, imag} */,
  {32'hc018d817, 32'h3e5735ce} /* (15, 17, 23) {real, imag} */,
  {32'hbe2e41db, 32'h4037320c} /* (15, 17, 22) {real, imag} */,
  {32'hbf237865, 32'h3f044da4} /* (15, 17, 21) {real, imag} */,
  {32'hbf6573cd, 32'h3eeab455} /* (15, 17, 20) {real, imag} */,
  {32'hbe503562, 32'hbe9d7e23} /* (15, 17, 19) {real, imag} */,
  {32'hc00fa97e, 32'hbed80984} /* (15, 17, 18) {real, imag} */,
  {32'h3f2d6686, 32'hbf2d2985} /* (15, 17, 17) {real, imag} */,
  {32'h3fbb0b88, 32'hbee515be} /* (15, 17, 16) {real, imag} */,
  {32'h3fd4df10, 32'hbf2b384d} /* (15, 17, 15) {real, imag} */,
  {32'h3fa68fa9, 32'hbe5f0950} /* (15, 17, 14) {real, imag} */,
  {32'h3f88ebbb, 32'h3ffc49ba} /* (15, 17, 13) {real, imag} */,
  {32'h4086ae75, 32'h3fda8d42} /* (15, 17, 12) {real, imag} */,
  {32'hbf7e4f95, 32'hbee499b1} /* (15, 17, 11) {real, imag} */,
  {32'hc01b6603, 32'h3eef8fce} /* (15, 17, 10) {real, imag} */,
  {32'hbf0dbf8e, 32'hbef711fd} /* (15, 17, 9) {real, imag} */,
  {32'hbecd6073, 32'hbed0898d} /* (15, 17, 8) {real, imag} */,
  {32'hc0156461, 32'hbec64132} /* (15, 17, 7) {real, imag} */,
  {32'h3f494566, 32'hbea46778} /* (15, 17, 6) {real, imag} */,
  {32'h3d1c43fe, 32'hbe679f2d} /* (15, 17, 5) {real, imag} */,
  {32'hbe88d8af, 32'h3e113eeb} /* (15, 17, 4) {real, imag} */,
  {32'h3f35ed42, 32'hbd46bcae} /* (15, 17, 3) {real, imag} */,
  {32'hbf0bb2d3, 32'hbe7adb79} /* (15, 17, 2) {real, imag} */,
  {32'h3f3aa1c0, 32'h3fcb3911} /* (15, 17, 1) {real, imag} */,
  {32'hbda5e566, 32'h3f994b53} /* (15, 17, 0) {real, imag} */,
  {32'hbf8fcb91, 32'hbc43f24b} /* (15, 16, 31) {real, imag} */,
  {32'hbe74be81, 32'hbe68f6df} /* (15, 16, 30) {real, imag} */,
  {32'hbf00faed, 32'hbfc9df37} /* (15, 16, 29) {real, imag} */,
  {32'hbfa19092, 32'hbf568133} /* (15, 16, 28) {real, imag} */,
  {32'hbf1f4fad, 32'hbf6c237d} /* (15, 16, 27) {real, imag} */,
  {32'hbf4a970a, 32'h3fa8501c} /* (15, 16, 26) {real, imag} */,
  {32'hbf6fdf5a, 32'h3d5ae745} /* (15, 16, 25) {real, imag} */,
  {32'hbf86259c, 32'hbf7b9aa5} /* (15, 16, 24) {real, imag} */,
  {32'hbd89138b, 32'hc033ee4e} /* (15, 16, 23) {real, imag} */,
  {32'h40679505, 32'hc005af35} /* (15, 16, 22) {real, imag} */,
  {32'hbf00ffed, 32'h3e15344e} /* (15, 16, 21) {real, imag} */,
  {32'h3f548705, 32'h3f7ca1e0} /* (15, 16, 20) {real, imag} */,
  {32'h3fda4479, 32'hbfbdbd4f} /* (15, 16, 19) {real, imag} */,
  {32'hbebd16fc, 32'h3e9a5c26} /* (15, 16, 18) {real, imag} */,
  {32'hbef4b215, 32'h3df0fcee} /* (15, 16, 17) {real, imag} */,
  {32'h3f09eccd, 32'h3e07173b} /* (15, 16, 16) {real, imag} */,
  {32'hbee7db82, 32'hbe0d04b4} /* (15, 16, 15) {real, imag} */,
  {32'hbfcc4354, 32'h3fee2f3d} /* (15, 16, 14) {real, imag} */,
  {32'hbfd0ce89, 32'hbf70d3d8} /* (15, 16, 13) {real, imag} */,
  {32'hbfa5e1f1, 32'hbfc3f12d} /* (15, 16, 12) {real, imag} */,
  {32'h3f032379, 32'hc04a3ec7} /* (15, 16, 11) {real, imag} */,
  {32'h3f2d3b0f, 32'h4048c6ab} /* (15, 16, 10) {real, imag} */,
  {32'hbfabfbf6, 32'h3ed05d3a} /* (15, 16, 9) {real, imag} */,
  {32'h3fd58bd4, 32'hbf0bd83e} /* (15, 16, 8) {real, imag} */,
  {32'hbf01d9b4, 32'hbf4a7a59} /* (15, 16, 7) {real, imag} */,
  {32'h3fada164, 32'hbe84bf07} /* (15, 16, 6) {real, imag} */,
  {32'h3f9cb468, 32'h3fe1f0e2} /* (15, 16, 5) {real, imag} */,
  {32'h3e9960aa, 32'h3f104c73} /* (15, 16, 4) {real, imag} */,
  {32'h3e91331c, 32'hbfbe2009} /* (15, 16, 3) {real, imag} */,
  {32'h3ed4646e, 32'h3f345219} /* (15, 16, 2) {real, imag} */,
  {32'h3ef86493, 32'h3f093b34} /* (15, 16, 1) {real, imag} */,
  {32'h3e87912a, 32'h3f147917} /* (15, 16, 0) {real, imag} */,
  {32'hbe4716d9, 32'hbf28e0ec} /* (15, 15, 31) {real, imag} */,
  {32'hbda808a2, 32'h3e1f295f} /* (15, 15, 30) {real, imag} */,
  {32'h3f1756f2, 32'h3f2ac46d} /* (15, 15, 29) {real, imag} */,
  {32'h3f0438df, 32'hbf53ef1e} /* (15, 15, 28) {real, imag} */,
  {32'h3fb4522b, 32'h3f831669} /* (15, 15, 27) {real, imag} */,
  {32'hbeae9ac4, 32'h3f2cf335} /* (15, 15, 26) {real, imag} */,
  {32'h3fa6b95b, 32'h3feef3d1} /* (15, 15, 25) {real, imag} */,
  {32'h3eb003e1, 32'hbf7b24fd} /* (15, 15, 24) {real, imag} */,
  {32'h3e2e3c78, 32'h3f80eb96} /* (15, 15, 23) {real, imag} */,
  {32'hbf941632, 32'hbec55b8a} /* (15, 15, 22) {real, imag} */,
  {32'hbfca4d88, 32'hbfed7d75} /* (15, 15, 21) {real, imag} */,
  {32'h4006bc8d, 32'hbf1ea21e} /* (15, 15, 20) {real, imag} */,
  {32'h3f0c30c8, 32'h3f662bd1} /* (15, 15, 19) {real, imag} */,
  {32'h3f140607, 32'h40044865} /* (15, 15, 18) {real, imag} */,
  {32'h3f2b9dee, 32'hbf40017d} /* (15, 15, 17) {real, imag} */,
  {32'h3ea87420, 32'hbd54109e} /* (15, 15, 16) {real, imag} */,
  {32'h3f11e700, 32'h4011a27f} /* (15, 15, 15) {real, imag} */,
  {32'h3fc88157, 32'hbf7231e9} /* (15, 15, 14) {real, imag} */,
  {32'h3f44afcf, 32'h3f3e0379} /* (15, 15, 13) {real, imag} */,
  {32'h4007bf40, 32'h40035647} /* (15, 15, 12) {real, imag} */,
  {32'hbfcffed4, 32'h3f9137b2} /* (15, 15, 11) {real, imag} */,
  {32'h40106f63, 32'h3fe84fcc} /* (15, 15, 10) {real, imag} */,
  {32'hbeb936c1, 32'h3f0ecb63} /* (15, 15, 9) {real, imag} */,
  {32'h3e5ddb7c, 32'hbf46e9a3} /* (15, 15, 8) {real, imag} */,
  {32'hbed3772f, 32'hbf13ca60} /* (15, 15, 7) {real, imag} */,
  {32'h3f09ca02, 32'h40200bab} /* (15, 15, 6) {real, imag} */,
  {32'h3f38d8c5, 32'hbfbfb675} /* (15, 15, 5) {real, imag} */,
  {32'h3ee2c9ca, 32'hbb3b4718} /* (15, 15, 4) {real, imag} */,
  {32'hbda79712, 32'hbe2a6a0f} /* (15, 15, 3) {real, imag} */,
  {32'hbf389339, 32'h3f2d2713} /* (15, 15, 2) {real, imag} */,
  {32'hbe88a4af, 32'h3f8a64d6} /* (15, 15, 1) {real, imag} */,
  {32'hbe51b948, 32'hbedb8a09} /* (15, 15, 0) {real, imag} */,
  {32'h3de7c1b5, 32'h3edac20f} /* (15, 14, 31) {real, imag} */,
  {32'hbea865ce, 32'h40111660} /* (15, 14, 30) {real, imag} */,
  {32'h3f4c7450, 32'hbebc7a7e} /* (15, 14, 29) {real, imag} */,
  {32'hbe4b9d03, 32'h3f69fb6c} /* (15, 14, 28) {real, imag} */,
  {32'h3f036c51, 32'hc00c970e} /* (15, 14, 27) {real, imag} */,
  {32'hbf719a57, 32'hbf9e9e2d} /* (15, 14, 26) {real, imag} */,
  {32'hbfbe31a9, 32'hbf8b3d7a} /* (15, 14, 25) {real, imag} */,
  {32'h3c46abe8, 32'h3ff35a72} /* (15, 14, 24) {real, imag} */,
  {32'h3ff00672, 32'hbd11992c} /* (15, 14, 23) {real, imag} */,
  {32'hbea11d23, 32'hbf16ca66} /* (15, 14, 22) {real, imag} */,
  {32'hbea28f52, 32'h3d95a785} /* (15, 14, 21) {real, imag} */,
  {32'hbffa47c4, 32'hbf0cdb72} /* (15, 14, 20) {real, imag} */,
  {32'hbe9e00fd, 32'hbfcfbdfd} /* (15, 14, 19) {real, imag} */,
  {32'hbeabe2d7, 32'h4016cce8} /* (15, 14, 18) {real, imag} */,
  {32'hbf954ea5, 32'hbf33d0e1} /* (15, 14, 17) {real, imag} */,
  {32'hbf9436ec, 32'hc0392c68} /* (15, 14, 16) {real, imag} */,
  {32'h3f838c8a, 32'hbf57b36c} /* (15, 14, 15) {real, imag} */,
  {32'hbf4cc461, 32'h3f51ee42} /* (15, 14, 14) {real, imag} */,
  {32'h3ed97a86, 32'h3fa4f4f8} /* (15, 14, 13) {real, imag} */,
  {32'h3fea7b96, 32'hbf540dc1} /* (15, 14, 12) {real, imag} */,
  {32'hbf91815b, 32'hbf8bdd56} /* (15, 14, 11) {real, imag} */,
  {32'hbf8629b3, 32'h3fbec190} /* (15, 14, 10) {real, imag} */,
  {32'h3fc896dc, 32'h4028e5b1} /* (15, 14, 9) {real, imag} */,
  {32'h3d463271, 32'hbf474438} /* (15, 14, 8) {real, imag} */,
  {32'h3f11f96b, 32'hbf3246fb} /* (15, 14, 7) {real, imag} */,
  {32'hbe442a96, 32'h3ee99ba8} /* (15, 14, 6) {real, imag} */,
  {32'hbf16399e, 32'hc00d0354} /* (15, 14, 5) {real, imag} */,
  {32'h3f64bb65, 32'hbfac4e49} /* (15, 14, 4) {real, imag} */,
  {32'hc00c5f10, 32'hbe457107} /* (15, 14, 3) {real, imag} */,
  {32'hbfd0f96f, 32'h3dcc51f1} /* (15, 14, 2) {real, imag} */,
  {32'h3f1581e5, 32'h3dae8ea7} /* (15, 14, 1) {real, imag} */,
  {32'h3fc3a815, 32'hc008487d} /* (15, 14, 0) {real, imag} */,
  {32'hbfb64e74, 32'h3f3e2124} /* (15, 13, 31) {real, imag} */,
  {32'h3e41a2c5, 32'hbff3efcd} /* (15, 13, 30) {real, imag} */,
  {32'h3ba5ccd3, 32'hbf928a17} /* (15, 13, 29) {real, imag} */,
  {32'h3fe3e333, 32'h3e99ec60} /* (15, 13, 28) {real, imag} */,
  {32'h3ee86266, 32'hbf46e29e} /* (15, 13, 27) {real, imag} */,
  {32'h3f4b3170, 32'hbf399954} /* (15, 13, 26) {real, imag} */,
  {32'hbf84cf29, 32'h3f10bf81} /* (15, 13, 25) {real, imag} */,
  {32'hbe44e2b5, 32'h3fcd620b} /* (15, 13, 24) {real, imag} */,
  {32'hc019f1d1, 32'hbed7653a} /* (15, 13, 23) {real, imag} */,
  {32'h3ecc6795, 32'hbffcf389} /* (15, 13, 22) {real, imag} */,
  {32'hbfb6a79f, 32'hbeba72f3} /* (15, 13, 21) {real, imag} */,
  {32'hbf4df0fa, 32'h3f738c78} /* (15, 13, 20) {real, imag} */,
  {32'hc01f1735, 32'hbf9b2411} /* (15, 13, 19) {real, imag} */,
  {32'hbdbb8691, 32'h4028c3c8} /* (15, 13, 18) {real, imag} */,
  {32'hbf61f115, 32'h3fc7bd4c} /* (15, 13, 17) {real, imag} */,
  {32'h3f40feec, 32'h3de96145} /* (15, 13, 16) {real, imag} */,
  {32'h404cb7dc, 32'hbf9ecc8f} /* (15, 13, 15) {real, imag} */,
  {32'hbf44e223, 32'h40580dc2} /* (15, 13, 14) {real, imag} */,
  {32'hc01f1e0f, 32'h3f99515d} /* (15, 13, 13) {real, imag} */,
  {32'hc02d59b1, 32'h3f7e3321} /* (15, 13, 12) {real, imag} */,
  {32'h3ff5af9c, 32'hbf9a14ce} /* (15, 13, 11) {real, imag} */,
  {32'hbf8ea908, 32'h3ed16994} /* (15, 13, 10) {real, imag} */,
  {32'h400befd9, 32'hc0089207} /* (15, 13, 9) {real, imag} */,
  {32'hbf3d1c68, 32'h3fe9f1f9} /* (15, 13, 8) {real, imag} */,
  {32'hbf0ea01b, 32'hbf1ae39f} /* (15, 13, 7) {real, imag} */,
  {32'h3f761154, 32'hc006c4ee} /* (15, 13, 6) {real, imag} */,
  {32'h3d7396e3, 32'h3f682e73} /* (15, 13, 5) {real, imag} */,
  {32'hbd6e79b0, 32'hbfc34751} /* (15, 13, 4) {real, imag} */,
  {32'h3f504942, 32'hbedc1c8b} /* (15, 13, 3) {real, imag} */,
  {32'hc0642a50, 32'h3ea9d4f0} /* (15, 13, 2) {real, imag} */,
  {32'hbfd38ad5, 32'h3d8d15a6} /* (15, 13, 1) {real, imag} */,
  {32'h3ec059e0, 32'h3f881b32} /* (15, 13, 0) {real, imag} */,
  {32'h40521d81, 32'hbd873841} /* (15, 12, 31) {real, imag} */,
  {32'h3f7a5f6a, 32'hbe671479} /* (15, 12, 30) {real, imag} */,
  {32'hbf0c149f, 32'hbfb5423f} /* (15, 12, 29) {real, imag} */,
  {32'h3f221a34, 32'h3f523211} /* (15, 12, 28) {real, imag} */,
  {32'h4020abf1, 32'h3f3b8e51} /* (15, 12, 27) {real, imag} */,
  {32'h3fab1f41, 32'h3d7b627b} /* (15, 12, 26) {real, imag} */,
  {32'hbf49a285, 32'hbfa0e150} /* (15, 12, 25) {real, imag} */,
  {32'hbed0107a, 32'h3ff67126} /* (15, 12, 24) {real, imag} */,
  {32'h3fa1d28d, 32'hbfc11ce8} /* (15, 12, 23) {real, imag} */,
  {32'h4006c83b, 32'h3f8c32d0} /* (15, 12, 22) {real, imag} */,
  {32'hbf074c66, 32'h3fa35863} /* (15, 12, 21) {real, imag} */,
  {32'h3fa16104, 32'hc040abaa} /* (15, 12, 20) {real, imag} */,
  {32'hbf8ef5b7, 32'h3fb40197} /* (15, 12, 19) {real, imag} */,
  {32'hbfcf3310, 32'hbc531847} /* (15, 12, 18) {real, imag} */,
  {32'h3d4f05d1, 32'h4071c512} /* (15, 12, 17) {real, imag} */,
  {32'hbf39dcd8, 32'h3fb8dbb8} /* (15, 12, 16) {real, imag} */,
  {32'hbe975d36, 32'hbe4c615f} /* (15, 12, 15) {real, imag} */,
  {32'hbfbfa723, 32'h3f45a9ee} /* (15, 12, 14) {real, imag} */,
  {32'h3d8d5b65, 32'hbe2e446f} /* (15, 12, 13) {real, imag} */,
  {32'hbd69df9d, 32'h3f954007} /* (15, 12, 12) {real, imag} */,
  {32'hbe14d744, 32'h3f289cb4} /* (15, 12, 11) {real, imag} */,
  {32'hc003d7fd, 32'hbfa1dc66} /* (15, 12, 10) {real, imag} */,
  {32'hbfa12c67, 32'h3f919de3} /* (15, 12, 9) {real, imag} */,
  {32'h3fe35e09, 32'hbed41abe} /* (15, 12, 8) {real, imag} */,
  {32'hbfad1628, 32'hbf563def} /* (15, 12, 7) {real, imag} */,
  {32'h3f435f1a, 32'h3e8fd109} /* (15, 12, 6) {real, imag} */,
  {32'hbfb278b1, 32'hbf1b6c7f} /* (15, 12, 5) {real, imag} */,
  {32'hbfae3142, 32'hbf3f9018} /* (15, 12, 4) {real, imag} */,
  {32'h3f263f8f, 32'h3d57c749} /* (15, 12, 3) {real, imag} */,
  {32'h3fcea723, 32'hbf8c0494} /* (15, 12, 2) {real, imag} */,
  {32'h3f9002f0, 32'hbec10439} /* (15, 12, 1) {real, imag} */,
  {32'hbfe919db, 32'h3f983312} /* (15, 12, 0) {real, imag} */,
  {32'hbdd07711, 32'h3fb0e1e6} /* (15, 11, 31) {real, imag} */,
  {32'h3e35ec1c, 32'hbf250c5f} /* (15, 11, 30) {real, imag} */,
  {32'h3f9bdd8d, 32'h3fa7c11d} /* (15, 11, 29) {real, imag} */,
  {32'hbfb410d6, 32'hbe5279d4} /* (15, 11, 28) {real, imag} */,
  {32'hbf2f1284, 32'hbc76992c} /* (15, 11, 27) {real, imag} */,
  {32'hbecefc1f, 32'h3d5a3489} /* (15, 11, 26) {real, imag} */,
  {32'h400fd44c, 32'hbf576ab8} /* (15, 11, 25) {real, imag} */,
  {32'hbefbf9dc, 32'h3fd75cf7} /* (15, 11, 24) {real, imag} */,
  {32'hbffa2d4f, 32'h3fa3b680} /* (15, 11, 23) {real, imag} */,
  {32'hc04368b2, 32'hbddba86b} /* (15, 11, 22) {real, imag} */,
  {32'hbfcbe7d6, 32'hbe8c58cc} /* (15, 11, 21) {real, imag} */,
  {32'h3fcf7a34, 32'hbea4ef30} /* (15, 11, 20) {real, imag} */,
  {32'hbf26970b, 32'h404dd0f5} /* (15, 11, 19) {real, imag} */,
  {32'h3f23edac, 32'hbe30ba42} /* (15, 11, 18) {real, imag} */,
  {32'h3e4fb0e9, 32'hbf8bdf5d} /* (15, 11, 17) {real, imag} */,
  {32'h3fd49f9d, 32'hc0204059} /* (15, 11, 16) {real, imag} */,
  {32'h3ed875c3, 32'hbe8f87b9} /* (15, 11, 15) {real, imag} */,
  {32'h3fb9c087, 32'hbca8524b} /* (15, 11, 14) {real, imag} */,
  {32'h3f4e9ca7, 32'hbf3bbb43} /* (15, 11, 13) {real, imag} */,
  {32'hbfbe6dda, 32'h403e2198} /* (15, 11, 12) {real, imag} */,
  {32'hbe9ed564, 32'h3e16bb8e} /* (15, 11, 11) {real, imag} */,
  {32'hbda1fbc0, 32'h3f02ca73} /* (15, 11, 10) {real, imag} */,
  {32'h3fe21964, 32'hbe8631f8} /* (15, 11, 9) {real, imag} */,
  {32'hc01fb69d, 32'hc00bd21d} /* (15, 11, 8) {real, imag} */,
  {32'h3fd7d298, 32'h3e9d646e} /* (15, 11, 7) {real, imag} */,
  {32'h3fed63c3, 32'h3edfd32b} /* (15, 11, 6) {real, imag} */,
  {32'h3ffc03bb, 32'hbf8cb294} /* (15, 11, 5) {real, imag} */,
  {32'hbf8400b5, 32'hc00239cc} /* (15, 11, 4) {real, imag} */,
  {32'hbc32bfd6, 32'hbf452b86} /* (15, 11, 3) {real, imag} */,
  {32'h3e9a2d46, 32'h3e8319df} /* (15, 11, 2) {real, imag} */,
  {32'h3f97baea, 32'h3eff5def} /* (15, 11, 1) {real, imag} */,
  {32'h3f0be871, 32'h3f9c09ac} /* (15, 11, 0) {real, imag} */,
  {32'h3ebe31df, 32'h3f8f7d11} /* (15, 10, 31) {real, imag} */,
  {32'h40000ffc, 32'hbf474254} /* (15, 10, 30) {real, imag} */,
  {32'hbefb5f9a, 32'hbf278ea5} /* (15, 10, 29) {real, imag} */,
  {32'h3e3ef23f, 32'h3f1f0c25} /* (15, 10, 28) {real, imag} */,
  {32'h3ed12325, 32'h3fe4557b} /* (15, 10, 27) {real, imag} */,
  {32'h3ee1d165, 32'h3facec80} /* (15, 10, 26) {real, imag} */,
  {32'hbf814f3a, 32'hc0230f28} /* (15, 10, 25) {real, imag} */,
  {32'hbf4a9c2d, 32'h3f576ce0} /* (15, 10, 24) {real, imag} */,
  {32'h3ff946e7, 32'hc043e999} /* (15, 10, 23) {real, imag} */,
  {32'hc08441c2, 32'hbf99f0f8} /* (15, 10, 22) {real, imag} */,
  {32'h3e37731c, 32'h3e20a966} /* (15, 10, 21) {real, imag} */,
  {32'h3fdc15fc, 32'h3fc618e7} /* (15, 10, 20) {real, imag} */,
  {32'h3f81c1e8, 32'hbe8bb785} /* (15, 10, 19) {real, imag} */,
  {32'hbfc5c551, 32'h3f34f63f} /* (15, 10, 18) {real, imag} */,
  {32'hbfbc2dd2, 32'h3ee4d273} /* (15, 10, 17) {real, imag} */,
  {32'h3f9e5c0c, 32'hbf433aa2} /* (15, 10, 16) {real, imag} */,
  {32'hbf9fb915, 32'hb9f5034f} /* (15, 10, 15) {real, imag} */,
  {32'hbf6aedfc, 32'hbfc7794d} /* (15, 10, 14) {real, imag} */,
  {32'h3fab3c24, 32'hc0301054} /* (15, 10, 13) {real, imag} */,
  {32'hbedfce88, 32'h3ff92f50} /* (15, 10, 12) {real, imag} */,
  {32'hbf3c92eb, 32'h3e854c91} /* (15, 10, 11) {real, imag} */,
  {32'hbe7609b9, 32'h402451c6} /* (15, 10, 10) {real, imag} */,
  {32'h3faa0cdc, 32'hbf1caf45} /* (15, 10, 9) {real, imag} */,
  {32'hbfbf3972, 32'h3f1dc051} /* (15, 10, 8) {real, imag} */,
  {32'hbf6646d9, 32'h3f06d65e} /* (15, 10, 7) {real, imag} */,
  {32'h3faee526, 32'h3fdde08c} /* (15, 10, 6) {real, imag} */,
  {32'h3eae187d, 32'hbf88e980} /* (15, 10, 5) {real, imag} */,
  {32'hbf09cc7c, 32'h4002af5d} /* (15, 10, 4) {real, imag} */,
  {32'h3d0bf12f, 32'hbf0a7b98} /* (15, 10, 3) {real, imag} */,
  {32'h3e35066f, 32'hbf535d62} /* (15, 10, 2) {real, imag} */,
  {32'hbf4780f8, 32'h3f0f4819} /* (15, 10, 1) {real, imag} */,
  {32'hbf877d26, 32'hbd3dd9af} /* (15, 10, 0) {real, imag} */,
  {32'h3dd60c17, 32'h3f80ff19} /* (15, 9, 31) {real, imag} */,
  {32'h3d95bfeb, 32'hbf2df189} /* (15, 9, 30) {real, imag} */,
  {32'hbef92fb9, 32'h3eabf1f7} /* (15, 9, 29) {real, imag} */,
  {32'h3cde9d9e, 32'hbf80cddc} /* (15, 9, 28) {real, imag} */,
  {32'h4010c440, 32'h3f21f712} /* (15, 9, 27) {real, imag} */,
  {32'h3e9179c8, 32'hbf0dfbaf} /* (15, 9, 26) {real, imag} */,
  {32'hbf107692, 32'h3d50c231} /* (15, 9, 25) {real, imag} */,
  {32'hc030d404, 32'h3ff48199} /* (15, 9, 24) {real, imag} */,
  {32'h3f68ef4b, 32'h3fb0ad67} /* (15, 9, 23) {real, imag} */,
  {32'h4035d26f, 32'hc0611c8d} /* (15, 9, 22) {real, imag} */,
  {32'hc066e4b5, 32'h3fdaec09} /* (15, 9, 21) {real, imag} */,
  {32'hbda4c377, 32'h3fd7f5fa} /* (15, 9, 20) {real, imag} */,
  {32'hbe972fbc, 32'h3f4a24d0} /* (15, 9, 19) {real, imag} */,
  {32'h3d7b0c7b, 32'h3f67ce9a} /* (15, 9, 18) {real, imag} */,
  {32'hbf75dfff, 32'hbf3b5ac3} /* (15, 9, 17) {real, imag} */,
  {32'hbf9bccc3, 32'hbf3fb4ef} /* (15, 9, 16) {real, imag} */,
  {32'hbfc57c84, 32'hbfc8cac5} /* (15, 9, 15) {real, imag} */,
  {32'hbfb6ebb5, 32'h40389686} /* (15, 9, 14) {real, imag} */,
  {32'h3f36bde7, 32'h3fbdd018} /* (15, 9, 13) {real, imag} */,
  {32'hc024f651, 32'hbf481bbe} /* (15, 9, 12) {real, imag} */,
  {32'hbfb9c1e1, 32'hbf8f0399} /* (15, 9, 11) {real, imag} */,
  {32'h40a21176, 32'hbfc5fa82} /* (15, 9, 10) {real, imag} */,
  {32'h3fc5e4ea, 32'h4044d7a9} /* (15, 9, 9) {real, imag} */,
  {32'hc030eac2, 32'hbfac0093} /* (15, 9, 8) {real, imag} */,
  {32'h3f9a67c0, 32'hbe86a3f4} /* (15, 9, 7) {real, imag} */,
  {32'h3f5288ae, 32'h4042b90f} /* (15, 9, 6) {real, imag} */,
  {32'h3d99db9a, 32'hbf62b68c} /* (15, 9, 5) {real, imag} */,
  {32'hbeb6f2cc, 32'hbfb8962d} /* (15, 9, 4) {real, imag} */,
  {32'h3f8e3304, 32'hbf6cd11a} /* (15, 9, 3) {real, imag} */,
  {32'h3f08a465, 32'hbfddef9c} /* (15, 9, 2) {real, imag} */,
  {32'h3fad3d25, 32'h3f881d68} /* (15, 9, 1) {real, imag} */,
  {32'h3ebd4a2c, 32'h3d87d0a0} /* (15, 9, 0) {real, imag} */,
  {32'h3ebb9430, 32'hbf01584e} /* (15, 8, 31) {real, imag} */,
  {32'hbc33f99e, 32'hbe405812} /* (15, 8, 30) {real, imag} */,
  {32'h3d90db44, 32'hbfc18cd1} /* (15, 8, 29) {real, imag} */,
  {32'h3fcc16b1, 32'h4024024a} /* (15, 8, 28) {real, imag} */,
  {32'h3f7d36d1, 32'h3f989a90} /* (15, 8, 27) {real, imag} */,
  {32'h3ffdba9d, 32'h3fd24c30} /* (15, 8, 26) {real, imag} */,
  {32'hbf9cd591, 32'hbfba7fe9} /* (15, 8, 25) {real, imag} */,
  {32'hbf7dc052, 32'hbffe8f63} /* (15, 8, 24) {real, imag} */,
  {32'hbf9ba4b9, 32'h400c7eeb} /* (15, 8, 23) {real, imag} */,
  {32'h40283bd5, 32'h3f7ec185} /* (15, 8, 22) {real, imag} */,
  {32'h3f8182ec, 32'h3ee5e11e} /* (15, 8, 21) {real, imag} */,
  {32'h402adb74, 32'h3f804e27} /* (15, 8, 20) {real, imag} */,
  {32'hbe9d191e, 32'h3eb7347f} /* (15, 8, 19) {real, imag} */,
  {32'h3d829e20, 32'hbf58d678} /* (15, 8, 18) {real, imag} */,
  {32'hbf2f0b56, 32'h3e524342} /* (15, 8, 17) {real, imag} */,
  {32'h3fd605cf, 32'h4006c2d5} /* (15, 8, 16) {real, imag} */,
  {32'hbf15b2b9, 32'h3f35e82b} /* (15, 8, 15) {real, imag} */,
  {32'h400eebb5, 32'hbf2d0998} /* (15, 8, 14) {real, imag} */,
  {32'h3f5af744, 32'hbfbd0446} /* (15, 8, 13) {real, imag} */,
  {32'hc002a394, 32'h3fbced59} /* (15, 8, 12) {real, imag} */,
  {32'h3f3ec1e3, 32'hbf9723ba} /* (15, 8, 11) {real, imag} */,
  {32'h3e9490d1, 32'h4023fda5} /* (15, 8, 10) {real, imag} */,
  {32'hbf81034d, 32'h3f995ac0} /* (15, 8, 9) {real, imag} */,
  {32'hbf4102ba, 32'h3fd12a94} /* (15, 8, 8) {real, imag} */,
  {32'hc00aa1d7, 32'h3f3fcdde} /* (15, 8, 7) {real, imag} */,
  {32'hbde93bdd, 32'hbff3ab0d} /* (15, 8, 6) {real, imag} */,
  {32'h3ef07e2a, 32'h3f802760} /* (15, 8, 5) {real, imag} */,
  {32'h40304003, 32'hbfb1ba58} /* (15, 8, 4) {real, imag} */,
  {32'h3f4186ff, 32'h3f09b42f} /* (15, 8, 3) {real, imag} */,
  {32'hbf530dbc, 32'hbf8cd77e} /* (15, 8, 2) {real, imag} */,
  {32'hc0204067, 32'hbef0642c} /* (15, 8, 1) {real, imag} */,
  {32'hc00c5ef2, 32'h3da3951c} /* (15, 8, 0) {real, imag} */,
  {32'hbfb283f5, 32'h40292203} /* (15, 7, 31) {real, imag} */,
  {32'h3fd277ba, 32'h3f8581fe} /* (15, 7, 30) {real, imag} */,
  {32'hbe82d762, 32'hbf884dca} /* (15, 7, 29) {real, imag} */,
  {32'hbf0d6b78, 32'h3ec4e1b4} /* (15, 7, 28) {real, imag} */,
  {32'h3ea7c769, 32'hbd6b12c6} /* (15, 7, 27) {real, imag} */,
  {32'hc031e533, 32'h3eebad37} /* (15, 7, 26) {real, imag} */,
  {32'hbf0ae046, 32'hbfe09af0} /* (15, 7, 25) {real, imag} */,
  {32'hbf113ba3, 32'hbd8de30f} /* (15, 7, 24) {real, imag} */,
  {32'hbf0d0d0c, 32'hbf91be1c} /* (15, 7, 23) {real, imag} */,
  {32'hc02187c4, 32'h3e3d41a7} /* (15, 7, 22) {real, imag} */,
  {32'h3f212b0b, 32'h40148f35} /* (15, 7, 21) {real, imag} */,
  {32'h3fa22f4a, 32'hbf0f3db1} /* (15, 7, 20) {real, imag} */,
  {32'h404cfa0c, 32'h400d9d29} /* (15, 7, 19) {real, imag} */,
  {32'h3f2501dc, 32'h3f63d132} /* (15, 7, 18) {real, imag} */,
  {32'h3e3135da, 32'hbfc7f132} /* (15, 7, 17) {real, imag} */,
  {32'h3e19b40d, 32'h3eedaea8} /* (15, 7, 16) {real, imag} */,
  {32'h3f8a4495, 32'hbee21f1d} /* (15, 7, 15) {real, imag} */,
  {32'hbf413d63, 32'hbf50ec13} /* (15, 7, 14) {real, imag} */,
  {32'hbe940d52, 32'hbe21c7c6} /* (15, 7, 13) {real, imag} */,
  {32'hbf11b708, 32'hbfd07671} /* (15, 7, 12) {real, imag} */,
  {32'h3f1d1d49, 32'h3f92fb41} /* (15, 7, 11) {real, imag} */,
  {32'h3fa8c5f5, 32'hc02d3c02} /* (15, 7, 10) {real, imag} */,
  {32'h4003595f, 32'h3f9c54b7} /* (15, 7, 9) {real, imag} */,
  {32'hbf80c4ae, 32'hbded44e0} /* (15, 7, 8) {real, imag} */,
  {32'h3cd44dd7, 32'h3f91661e} /* (15, 7, 7) {real, imag} */,
  {32'hc01929af, 32'h3dbebd31} /* (15, 7, 6) {real, imag} */,
  {32'h4018f556, 32'h3da79710} /* (15, 7, 5) {real, imag} */,
  {32'h3f60e258, 32'hc00e8f58} /* (15, 7, 4) {real, imag} */,
  {32'h3f1e0f48, 32'hbe162578} /* (15, 7, 3) {real, imag} */,
  {32'h4023cada, 32'h3fa08160} /* (15, 7, 2) {real, imag} */,
  {32'h3ecbd200, 32'h4001bb38} /* (15, 7, 1) {real, imag} */,
  {32'hbcf65638, 32'h3f5ad7c3} /* (15, 7, 0) {real, imag} */,
  {32'hbf359da5, 32'h3eafdd15} /* (15, 6, 31) {real, imag} */,
  {32'h3dd027a7, 32'h3fac0cf6} /* (15, 6, 30) {real, imag} */,
  {32'h3f1ec538, 32'h3e42eb43} /* (15, 6, 29) {real, imag} */,
  {32'h3fa56795, 32'h3edba797} /* (15, 6, 28) {real, imag} */,
  {32'h3f17bd33, 32'hc019fa50} /* (15, 6, 27) {real, imag} */,
  {32'h40466fa3, 32'h3da5294c} /* (15, 6, 26) {real, imag} */,
  {32'hbe9c4273, 32'h3f94626b} /* (15, 6, 25) {real, imag} */,
  {32'hbe704ee7, 32'hbfbc5eb2} /* (15, 6, 24) {real, imag} */,
  {32'hbfaba9db, 32'hbdeed12d} /* (15, 6, 23) {real, imag} */,
  {32'h402426e7, 32'h4010adf9} /* (15, 6, 22) {real, imag} */,
  {32'h3f853853, 32'h3f98b66a} /* (15, 6, 21) {real, imag} */,
  {32'hbeaf73d6, 32'hbf079037} /* (15, 6, 20) {real, imag} */,
  {32'hbbd6bfd5, 32'hbfd39c02} /* (15, 6, 19) {real, imag} */,
  {32'h3fa946af, 32'h3f7b91be} /* (15, 6, 18) {real, imag} */,
  {32'h3d0d74bb, 32'h3fa435bb} /* (15, 6, 17) {real, imag} */,
  {32'hbf07c162, 32'hbf0ff7f9} /* (15, 6, 16) {real, imag} */,
  {32'hbdc91d3c, 32'hbe8a91d2} /* (15, 6, 15) {real, imag} */,
  {32'h402f6297, 32'hc005d2b5} /* (15, 6, 14) {real, imag} */,
  {32'h3f8b7800, 32'h3fb25135} /* (15, 6, 13) {real, imag} */,
  {32'hbfd806e8, 32'h3ea42ecc} /* (15, 6, 12) {real, imag} */,
  {32'h4006314f, 32'h3efc303e} /* (15, 6, 11) {real, imag} */,
  {32'h3d0d58a5, 32'h4030295e} /* (15, 6, 10) {real, imag} */,
  {32'hbeb755e4, 32'hc0255697} /* (15, 6, 9) {real, imag} */,
  {32'hc0958613, 32'hbfea7693} /* (15, 6, 8) {real, imag} */,
  {32'h3eb6842a, 32'hbeb11a1d} /* (15, 6, 7) {real, imag} */,
  {32'hbfb932e6, 32'h3e0a1a79} /* (15, 6, 6) {real, imag} */,
  {32'hbf325478, 32'h3f2c2bf0} /* (15, 6, 5) {real, imag} */,
  {32'h3fe85193, 32'h3e15d9f0} /* (15, 6, 4) {real, imag} */,
  {32'h3f780143, 32'hbf7c6ac7} /* (15, 6, 3) {real, imag} */,
  {32'h3f235d0a, 32'hbf13981d} /* (15, 6, 2) {real, imag} */,
  {32'hbf5cb6f7, 32'h3f86598b} /* (15, 6, 1) {real, imag} */,
  {32'hbf6efa69, 32'hbe672eef} /* (15, 6, 0) {real, imag} */,
  {32'h3fa7d94e, 32'hbdc77e45} /* (15, 5, 31) {real, imag} */,
  {32'h3f15a499, 32'h3f813716} /* (15, 5, 30) {real, imag} */,
  {32'h3de34343, 32'h4031e6f2} /* (15, 5, 29) {real, imag} */,
  {32'h3f92d028, 32'h3eda007b} /* (15, 5, 28) {real, imag} */,
  {32'h3f9ed175, 32'hbdec67df} /* (15, 5, 27) {real, imag} */,
  {32'h4011a322, 32'hc039bcf4} /* (15, 5, 26) {real, imag} */,
  {32'h3f7635ae, 32'h3ff95e66} /* (15, 5, 25) {real, imag} */,
  {32'hbf2c3305, 32'hbec2d032} /* (15, 5, 24) {real, imag} */,
  {32'hbf743c27, 32'h3ff6f2e7} /* (15, 5, 23) {real, imag} */,
  {32'h3d9853c8, 32'h3f59cb93} /* (15, 5, 22) {real, imag} */,
  {32'h3f180f4e, 32'h3ed8df3f} /* (15, 5, 21) {real, imag} */,
  {32'hbf17a806, 32'h3fdefa78} /* (15, 5, 20) {real, imag} */,
  {32'hbf3d5626, 32'h3c9d8f7c} /* (15, 5, 19) {real, imag} */,
  {32'h3e4fdd5e, 32'h3f2734c6} /* (15, 5, 18) {real, imag} */,
  {32'h3ebbbd94, 32'hbf9f8610} /* (15, 5, 17) {real, imag} */,
  {32'hbf2a2ae4, 32'h3e9b5bd7} /* (15, 5, 16) {real, imag} */,
  {32'h3de4579f, 32'h3ee75335} /* (15, 5, 15) {real, imag} */,
  {32'hbf86a1b3, 32'hbfdb1b70} /* (15, 5, 14) {real, imag} */,
  {32'hc00ba6d5, 32'h3f287f53} /* (15, 5, 13) {real, imag} */,
  {32'h3ec3d7f6, 32'hbe97249b} /* (15, 5, 12) {real, imag} */,
  {32'h3fde8c78, 32'h3fbf9953} /* (15, 5, 11) {real, imag} */,
  {32'hbf5e7cf6, 32'h3ea51453} /* (15, 5, 10) {real, imag} */,
  {32'hbeaea8e6, 32'hbf9d38cb} /* (15, 5, 9) {real, imag} */,
  {32'h3f480d4f, 32'hbfc2930a} /* (15, 5, 8) {real, imag} */,
  {32'h3f90dd03, 32'hbf895e91} /* (15, 5, 7) {real, imag} */,
  {32'hbe421711, 32'h3f0a89d7} /* (15, 5, 6) {real, imag} */,
  {32'hbfb4e33f, 32'hbf4affe5} /* (15, 5, 5) {real, imag} */,
  {32'h4032b8c2, 32'hbf9cb962} /* (15, 5, 4) {real, imag} */,
  {32'h3f648615, 32'h3fefecbf} /* (15, 5, 3) {real, imag} */,
  {32'hbf2ff800, 32'h3fd336a5} /* (15, 5, 2) {real, imag} */,
  {32'h40021842, 32'hbed994c6} /* (15, 5, 1) {real, imag} */,
  {32'h3f5d5622, 32'hbfa4903c} /* (15, 5, 0) {real, imag} */,
  {32'h3ec716f6, 32'h3ff6c87c} /* (15, 4, 31) {real, imag} */,
  {32'hbd179372, 32'h3fe2e454} /* (15, 4, 30) {real, imag} */,
  {32'hbe4a0dfb, 32'h3d8cee3b} /* (15, 4, 29) {real, imag} */,
  {32'h3f158a9c, 32'hbfcf734a} /* (15, 4, 28) {real, imag} */,
  {32'h3e680104, 32'hbeb6bc20} /* (15, 4, 27) {real, imag} */,
  {32'hbfad67b7, 32'hbfd3c0ec} /* (15, 4, 26) {real, imag} */,
  {32'h4053fec8, 32'h3fbff6aa} /* (15, 4, 25) {real, imag} */,
  {32'hbd5064eb, 32'hbf7b2505} /* (15, 4, 24) {real, imag} */,
  {32'h3ecbb8d8, 32'hbe666deb} /* (15, 4, 23) {real, imag} */,
  {32'h3fa4c152, 32'hbdc1a8fb} /* (15, 4, 22) {real, imag} */,
  {32'h3d74941e, 32'h3ff4f0fa} /* (15, 4, 21) {real, imag} */,
  {32'h3ec5d48d, 32'hc0063596} /* (15, 4, 20) {real, imag} */,
  {32'hbf8bf166, 32'hbecb6975} /* (15, 4, 19) {real, imag} */,
  {32'h3f35ff73, 32'h3fc751db} /* (15, 4, 18) {real, imag} */,
  {32'h3eeddef8, 32'hc02f0c0e} /* (15, 4, 17) {real, imag} */,
  {32'h3ee9a3a6, 32'h3f5f3902} /* (15, 4, 16) {real, imag} */,
  {32'h3f1c6287, 32'h3f896326} /* (15, 4, 15) {real, imag} */,
  {32'h3f305ce7, 32'hbf09a88e} /* (15, 4, 14) {real, imag} */,
  {32'h3fe1b1a6, 32'hbe62cc86} /* (15, 4, 13) {real, imag} */,
  {32'hbf5b3d42, 32'h402bba8f} /* (15, 4, 12) {real, imag} */,
  {32'h3fe2f5f0, 32'hc00d7554} /* (15, 4, 11) {real, imag} */,
  {32'hc0746db0, 32'hbf03cb88} /* (15, 4, 10) {real, imag} */,
  {32'hbf602572, 32'h3cbc3f54} /* (15, 4, 9) {real, imag} */,
  {32'hbf690a2f, 32'hbece6f1b} /* (15, 4, 8) {real, imag} */,
  {32'hbf8ce9f0, 32'h3f4d43e1} /* (15, 4, 7) {real, imag} */,
  {32'hbd17fbb9, 32'hbfad4d90} /* (15, 4, 6) {real, imag} */,
  {32'h3fb56660, 32'h3ed5127d} /* (15, 4, 5) {real, imag} */,
  {32'h3faa7c7d, 32'h3ff2d255} /* (15, 4, 4) {real, imag} */,
  {32'hbe2830e9, 32'hc0103f78} /* (15, 4, 3) {real, imag} */,
  {32'hbbae8008, 32'hc0004d6a} /* (15, 4, 2) {real, imag} */,
  {32'h3dd68806, 32'hbff57b23} /* (15, 4, 1) {real, imag} */,
  {32'hc02641f7, 32'h3f163fee} /* (15, 4, 0) {real, imag} */,
  {32'h3f634e23, 32'h3e2b3fc6} /* (15, 3, 31) {real, imag} */,
  {32'hbff0bbb3, 32'hc00c67fa} /* (15, 3, 30) {real, imag} */,
  {32'h3cba7973, 32'hbfdc3379} /* (15, 3, 29) {real, imag} */,
  {32'hbe7918cb, 32'hbddb17b2} /* (15, 3, 28) {real, imag} */,
  {32'h40113cc6, 32'h3eabb745} /* (15, 3, 27) {real, imag} */,
  {32'h3f978c70, 32'h3f4dfd64} /* (15, 3, 26) {real, imag} */,
  {32'hbf7c71da, 32'h3fcb9736} /* (15, 3, 25) {real, imag} */,
  {32'hbf6d8b2f, 32'hbf8b2f29} /* (15, 3, 24) {real, imag} */,
  {32'h3eeef134, 32'h3d78a5e0} /* (15, 3, 23) {real, imag} */,
  {32'h3fd5ed76, 32'hbe3798ef} /* (15, 3, 22) {real, imag} */,
  {32'hc05b4c07, 32'h3fb02398} /* (15, 3, 21) {real, imag} */,
  {32'hbfe939ee, 32'h3f3e2ac2} /* (15, 3, 20) {real, imag} */,
  {32'hc025907d, 32'h3e3017eb} /* (15, 3, 19) {real, imag} */,
  {32'h3f266a5e, 32'hbf5a1032} /* (15, 3, 18) {real, imag} */,
  {32'h4012507e, 32'h3fb7a88a} /* (15, 3, 17) {real, imag} */,
  {32'hbee929ae, 32'h3e3e2a38} /* (15, 3, 16) {real, imag} */,
  {32'h3d80f20d, 32'hbf68b90d} /* (15, 3, 15) {real, imag} */,
  {32'hbf900fd1, 32'h3f83d2d9} /* (15, 3, 14) {real, imag} */,
  {32'h3f5f5b7b, 32'h40053bff} /* (15, 3, 13) {real, imag} */,
  {32'h3fc5009b, 32'hbfda6e98} /* (15, 3, 12) {real, imag} */,
  {32'hbf767706, 32'h3f89afb8} /* (15, 3, 11) {real, imag} */,
  {32'hbfec291b, 32'h4034d193} /* (15, 3, 10) {real, imag} */,
  {32'hbf98d5a2, 32'h3d81d472} /* (15, 3, 9) {real, imag} */,
  {32'h3fb4937d, 32'hbf447277} /* (15, 3, 8) {real, imag} */,
  {32'h3e6afeb3, 32'hbf665b6c} /* (15, 3, 7) {real, imag} */,
  {32'h3dd41898, 32'h3f92978c} /* (15, 3, 6) {real, imag} */,
  {32'h3fe5a4c1, 32'hbd85a8e1} /* (15, 3, 5) {real, imag} */,
  {32'h3edeb1b2, 32'h3d821171} /* (15, 3, 4) {real, imag} */,
  {32'h3e8c9b83, 32'h3f841797} /* (15, 3, 3) {real, imag} */,
  {32'hbe6140ac, 32'h3e1dbd86} /* (15, 3, 2) {real, imag} */,
  {32'h3fd08d6d, 32'h3eaf8868} /* (15, 3, 1) {real, imag} */,
  {32'hbfc5f499, 32'h3f2f00af} /* (15, 3, 0) {real, imag} */,
  {32'hbf68f536, 32'hbeb5260c} /* (15, 2, 31) {real, imag} */,
  {32'hbf9a774b, 32'hbe7edf65} /* (15, 2, 30) {real, imag} */,
  {32'h3fa1569a, 32'h3f06214c} /* (15, 2, 29) {real, imag} */,
  {32'hbe86e6d2, 32'hbf78e638} /* (15, 2, 28) {real, imag} */,
  {32'h3ff92aa3, 32'h3f624b3a} /* (15, 2, 27) {real, imag} */,
  {32'h3ed994a0, 32'h403e4912} /* (15, 2, 26) {real, imag} */,
  {32'hbeb9e570, 32'h3fe70d50} /* (15, 2, 25) {real, imag} */,
  {32'hbf24e76a, 32'hbfbf9a3c} /* (15, 2, 24) {real, imag} */,
  {32'hbfd705bc, 32'hc00ce850} /* (15, 2, 23) {real, imag} */,
  {32'h3f235030, 32'hbf64e082} /* (15, 2, 22) {real, imag} */,
  {32'hbe4f5e38, 32'hc05a7516} /* (15, 2, 21) {real, imag} */,
  {32'hbf9305c7, 32'h3d354849} /* (15, 2, 20) {real, imag} */,
  {32'h3f0061ba, 32'h3ff02c3c} /* (15, 2, 19) {real, imag} */,
  {32'h3e626030, 32'hbf1cedc7} /* (15, 2, 18) {real, imag} */,
  {32'h3f5a34e4, 32'hbfda48aa} /* (15, 2, 17) {real, imag} */,
  {32'h3eb5d6c9, 32'hbfda4df2} /* (15, 2, 16) {real, imag} */,
  {32'hbf349d0f, 32'h3ef7123b} /* (15, 2, 15) {real, imag} */,
  {32'hbfcea1e0, 32'hbf171ec0} /* (15, 2, 14) {real, imag} */,
  {32'h3d9298a6, 32'h3ff2d967} /* (15, 2, 13) {real, imag} */,
  {32'h3f8eba1a, 32'hbf869e44} /* (15, 2, 12) {real, imag} */,
  {32'h3e48b437, 32'hbfa59665} /* (15, 2, 11) {real, imag} */,
  {32'hbe615a55, 32'h3f2fe733} /* (15, 2, 10) {real, imag} */,
  {32'h3e215173, 32'h3f5a637e} /* (15, 2, 9) {real, imag} */,
  {32'hbf5a9ebe, 32'h3f0aad17} /* (15, 2, 8) {real, imag} */,
  {32'hbe55d896, 32'hbd0c9f60} /* (15, 2, 7) {real, imag} */,
  {32'hbeba85a6, 32'hc0397ae6} /* (15, 2, 6) {real, imag} */,
  {32'h3f80c55f, 32'hbf2d20a9} /* (15, 2, 5) {real, imag} */,
  {32'hbf3e190d, 32'h3c4eaa38} /* (15, 2, 4) {real, imag} */,
  {32'hc01ef885, 32'h3f71852d} /* (15, 2, 3) {real, imag} */,
  {32'h3f8fbb0c, 32'hbf79cad9} /* (15, 2, 2) {real, imag} */,
  {32'hbfe42a7c, 32'hbfbcff38} /* (15, 2, 1) {real, imag} */,
  {32'h3e95acad, 32'h4027179d} /* (15, 2, 0) {real, imag} */,
  {32'h3fe97c8d, 32'h3ed97682} /* (15, 1, 31) {real, imag} */,
  {32'hbf707c4e, 32'h3f517b55} /* (15, 1, 30) {real, imag} */,
  {32'h3f77752d, 32'h3f1172f4} /* (15, 1, 29) {real, imag} */,
  {32'h3ef53360, 32'hbd1fe423} /* (15, 1, 28) {real, imag} */,
  {32'h3f08202b, 32'hbdd92afe} /* (15, 1, 27) {real, imag} */,
  {32'hbf9956ac, 32'h3e6e1e42} /* (15, 1, 26) {real, imag} */,
  {32'h3f40767d, 32'h3c1c503e} /* (15, 1, 25) {real, imag} */,
  {32'hbec8381a, 32'h3fcf6765} /* (15, 1, 24) {real, imag} */,
  {32'h403b888f, 32'h3f8d85c5} /* (15, 1, 23) {real, imag} */,
  {32'h3e5e0f22, 32'h3f39c547} /* (15, 1, 22) {real, imag} */,
  {32'h3e097fb3, 32'hbf25382a} /* (15, 1, 21) {real, imag} */,
  {32'h3fca1ac8, 32'h3fe84b99} /* (15, 1, 20) {real, imag} */,
  {32'hbf30d1db, 32'hbfaa4b7b} /* (15, 1, 19) {real, imag} */,
  {32'h3ec9f78d, 32'hbf0560de} /* (15, 1, 18) {real, imag} */,
  {32'h3e18dd58, 32'hbf39df0c} /* (15, 1, 17) {real, imag} */,
  {32'hc0034712, 32'hc000e57c} /* (15, 1, 16) {real, imag} */,
  {32'h3f113aa0, 32'hbeb8c647} /* (15, 1, 15) {real, imag} */,
  {32'h3e8491ac, 32'hbfd378a6} /* (15, 1, 14) {real, imag} */,
  {32'h3f779cff, 32'hbf10c976} /* (15, 1, 13) {real, imag} */,
  {32'h3f868d92, 32'hbfd7cc09} /* (15, 1, 12) {real, imag} */,
  {32'h3f7c6cdb, 32'h3fcfefcc} /* (15, 1, 11) {real, imag} */,
  {32'h3f6a5460, 32'hbf81e409} /* (15, 1, 10) {real, imag} */,
  {32'h3fe49559, 32'h3fd22377} /* (15, 1, 9) {real, imag} */,
  {32'hbf8992d8, 32'hbf2f6d9d} /* (15, 1, 8) {real, imag} */,
  {32'h3f2efc71, 32'h3faf30d4} /* (15, 1, 7) {real, imag} */,
  {32'h3e3462e3, 32'h3f198541} /* (15, 1, 6) {real, imag} */,
  {32'hbfe902bc, 32'h3f26e949} /* (15, 1, 5) {real, imag} */,
  {32'h3f5384b5, 32'h3f86d8b1} /* (15, 1, 4) {real, imag} */,
  {32'hbf7b3fb3, 32'hbf0dc7c0} /* (15, 1, 3) {real, imag} */,
  {32'hbff8ee7d, 32'hbff7be5a} /* (15, 1, 2) {real, imag} */,
  {32'h40511ec0, 32'h3f47af05} /* (15, 1, 1) {real, imag} */,
  {32'h3fb21377, 32'h3f8d27de} /* (15, 1, 0) {real, imag} */,
  {32'h3dc8437d, 32'hc010d8a0} /* (15, 0, 31) {real, imag} */,
  {32'h3efb4f57, 32'h3f9ddb2c} /* (15, 0, 30) {real, imag} */,
  {32'hbec0ba3a, 32'hbff1d194} /* (15, 0, 29) {real, imag} */,
  {32'hbfe514ad, 32'hbf81f94e} /* (15, 0, 28) {real, imag} */,
  {32'hbf370a9f, 32'h3f72b8d9} /* (15, 0, 27) {real, imag} */,
  {32'hbf05f859, 32'hbf8625f1} /* (15, 0, 26) {real, imag} */,
  {32'h3f1c58c2, 32'h3e1c26f3} /* (15, 0, 25) {real, imag} */,
  {32'hbfaeed9f, 32'hbc19556c} /* (15, 0, 24) {real, imag} */,
  {32'h3f50deda, 32'h3f473f58} /* (15, 0, 23) {real, imag} */,
  {32'h3f95d059, 32'hbf496e6d} /* (15, 0, 22) {real, imag} */,
  {32'hbf3a5626, 32'h3ee5e02a} /* (15, 0, 21) {real, imag} */,
  {32'h3e90eed7, 32'hbf44e3d5} /* (15, 0, 20) {real, imag} */,
  {32'hbfc42213, 32'h4006f0d2} /* (15, 0, 19) {real, imag} */,
  {32'h4049f3cf, 32'hbf010efb} /* (15, 0, 18) {real, imag} */,
  {32'h3f0ea30c, 32'h3f8a7803} /* (15, 0, 17) {real, imag} */,
  {32'h3f19bb43, 32'h3ead3075} /* (15, 0, 16) {real, imag} */,
  {32'hbd497a38, 32'hbf816bef} /* (15, 0, 15) {real, imag} */,
  {32'hbfb6ad6a, 32'hbf4785bf} /* (15, 0, 14) {real, imag} */,
  {32'h4007e254, 32'h3f26f718} /* (15, 0, 13) {real, imag} */,
  {32'h3f4ba22a, 32'h3e6641f6} /* (15, 0, 12) {real, imag} */,
  {32'hbf81315e, 32'h3fe361d2} /* (15, 0, 11) {real, imag} */,
  {32'hbf26770d, 32'h3f5abacc} /* (15, 0, 10) {real, imag} */,
  {32'h3d8c6d3a, 32'h400e82f2} /* (15, 0, 9) {real, imag} */,
  {32'h404d5e9c, 32'hbf926da6} /* (15, 0, 8) {real, imag} */,
  {32'h3f4446cd, 32'hc01571dc} /* (15, 0, 7) {real, imag} */,
  {32'h3f4d3e85, 32'h3eea1d6e} /* (15, 0, 6) {real, imag} */,
  {32'hbe4c6b6a, 32'hbe69d500} /* (15, 0, 5) {real, imag} */,
  {32'hbfdb7095, 32'hbeb22468} /* (15, 0, 4) {real, imag} */,
  {32'hbfc45292, 32'hbffcfd67} /* (15, 0, 3) {real, imag} */,
  {32'h3c381615, 32'hba300204} /* (15, 0, 2) {real, imag} */,
  {32'hbf754673, 32'hbec821b1} /* (15, 0, 1) {real, imag} */,
  {32'h3f32920e, 32'h3f71358b} /* (15, 0, 0) {real, imag} */,
  {32'hc0b00dcb, 32'h3fa46337} /* (14, 31, 31) {real, imag} */,
  {32'h3f6c3eab, 32'hc055b25b} /* (14, 31, 30) {real, imag} */,
  {32'h3fd0fea4, 32'h3fa9e29c} /* (14, 31, 29) {real, imag} */,
  {32'hbe66489a, 32'h3f6056a8} /* (14, 31, 28) {real, imag} */,
  {32'hbfcefb5c, 32'hbf2668ae} /* (14, 31, 27) {real, imag} */,
  {32'hbf1d7c9e, 32'hbffa526a} /* (14, 31, 26) {real, imag} */,
  {32'hc04c61cc, 32'hbf69af87} /* (14, 31, 25) {real, imag} */,
  {32'h3e0f1b7c, 32'hc01b419d} /* (14, 31, 24) {real, imag} */,
  {32'h3f679673, 32'hbf9fe3ee} /* (14, 31, 23) {real, imag} */,
  {32'h4023710e, 32'h3f87ab50} /* (14, 31, 22) {real, imag} */,
  {32'h400de8a0, 32'hc023fe13} /* (14, 31, 21) {real, imag} */,
  {32'h3f2e963d, 32'h3e88fbb5} /* (14, 31, 20) {real, imag} */,
  {32'h3ef543c7, 32'h3f4a4e3f} /* (14, 31, 19) {real, imag} */,
  {32'h3fb8d597, 32'h3d0a3b4c} /* (14, 31, 18) {real, imag} */,
  {32'hbfb3aeef, 32'hbec25e89} /* (14, 31, 17) {real, imag} */,
  {32'h3ed6632f, 32'hbfe42260} /* (14, 31, 16) {real, imag} */,
  {32'hbf8f8dcd, 32'h3f40516f} /* (14, 31, 15) {real, imag} */,
  {32'h3ed0ca3e, 32'hbf476807} /* (14, 31, 14) {real, imag} */,
  {32'hbff006a7, 32'hbe7881b0} /* (14, 31, 13) {real, imag} */,
  {32'hbf201953, 32'hbc78240c} /* (14, 31, 12) {real, imag} */,
  {32'h404b576b, 32'h3d15e57d} /* (14, 31, 11) {real, imag} */,
  {32'hc03d1811, 32'hbf8a35fd} /* (14, 31, 10) {real, imag} */,
  {32'h3f436756, 32'hbf8c0629} /* (14, 31, 9) {real, imag} */,
  {32'h3e30dc6b, 32'hc007adc3} /* (14, 31, 8) {real, imag} */,
  {32'h3fd9f702, 32'hbf373ca5} /* (14, 31, 7) {real, imag} */,
  {32'hbefa11f4, 32'h4022fd0e} /* (14, 31, 6) {real, imag} */,
  {32'h3fac482e, 32'h3f76e5d0} /* (14, 31, 5) {real, imag} */,
  {32'hbcce9749, 32'h3f6324c3} /* (14, 31, 4) {real, imag} */,
  {32'h3f476487, 32'h3b450ef7} /* (14, 31, 3) {real, imag} */,
  {32'h3fb36a21, 32'hbf6a462c} /* (14, 31, 2) {real, imag} */,
  {32'hc07df3ac, 32'h3f5b45ef} /* (14, 31, 1) {real, imag} */,
  {32'hc03c4dbd, 32'hbe0fb841} /* (14, 31, 0) {real, imag} */,
  {32'h40b0771d, 32'hbec8a1ff} /* (14, 30, 31) {real, imag} */,
  {32'hc060b778, 32'h3f2fdf06} /* (14, 30, 30) {real, imag} */,
  {32'hbe5031b4, 32'h3f2ab9aa} /* (14, 30, 29) {real, imag} */,
  {32'hbde84ad6, 32'h3fec1935} /* (14, 30, 28) {real, imag} */,
  {32'hbfdcf19b, 32'h3fd5e926} /* (14, 30, 27) {real, imag} */,
  {32'hbf8cb089, 32'hbe19b3f1} /* (14, 30, 26) {real, imag} */,
  {32'h3f8ead60, 32'h3fa1f9e5} /* (14, 30, 25) {real, imag} */,
  {32'hc0024e98, 32'hbf331ab1} /* (14, 30, 24) {real, imag} */,
  {32'h3d224423, 32'hbf8a9b3a} /* (14, 30, 23) {real, imag} */,
  {32'h4026d91a, 32'hbec56334} /* (14, 30, 22) {real, imag} */,
  {32'hbe990b5f, 32'h3f7a1821} /* (14, 30, 21) {real, imag} */,
  {32'hbeafa363, 32'h3e9e907c} /* (14, 30, 20) {real, imag} */,
  {32'hc0482179, 32'h3f0d9449} /* (14, 30, 19) {real, imag} */,
  {32'h3f4db245, 32'hbe64d18b} /* (14, 30, 18) {real, imag} */,
  {32'hbe910184, 32'hbeb63d6b} /* (14, 30, 17) {real, imag} */,
  {32'hbfb2644a, 32'hbf1d9c09} /* (14, 30, 16) {real, imag} */,
  {32'hbfeb53cd, 32'h3f4bd02e} /* (14, 30, 15) {real, imag} */,
  {32'hbd463cc2, 32'h4007b646} /* (14, 30, 14) {real, imag} */,
  {32'hbdf12b1b, 32'h3f84ee64} /* (14, 30, 13) {real, imag} */,
  {32'h40088dba, 32'hbf51b19e} /* (14, 30, 12) {real, imag} */,
  {32'hbfa89251, 32'h3f1832e6} /* (14, 30, 11) {real, imag} */,
  {32'h3ff0c7fe, 32'hc00b3000} /* (14, 30, 10) {real, imag} */,
  {32'h40188c17, 32'hbf081b8f} /* (14, 30, 9) {real, imag} */,
  {32'hbfc79a92, 32'h3e10eb83} /* (14, 30, 8) {real, imag} */,
  {32'hbf87826f, 32'h3f5c27e8} /* (14, 30, 7) {real, imag} */,
  {32'h3f3522b6, 32'h3ed24c77} /* (14, 30, 6) {real, imag} */,
  {32'hbf9cfabb, 32'h3f017e05} /* (14, 30, 5) {real, imag} */,
  {32'h400a5bc7, 32'h3f880333} /* (14, 30, 4) {real, imag} */,
  {32'h40023a9d, 32'hbf88360c} /* (14, 30, 3) {real, imag} */,
  {32'hc0684acd, 32'h3e9493c7} /* (14, 30, 2) {real, imag} */,
  {32'h40ab856b, 32'hc006cad8} /* (14, 30, 1) {real, imag} */,
  {32'h4020173e, 32'h3ed7527e} /* (14, 30, 0) {real, imag} */,
  {32'hc01dfb7b, 32'hbd9e1800} /* (14, 29, 31) {real, imag} */,
  {32'h3f83f546, 32'hbf82ec5b} /* (14, 29, 30) {real, imag} */,
  {32'h3f067d33, 32'hc022204b} /* (14, 29, 29) {real, imag} */,
  {32'h3c81a768, 32'hbf622609} /* (14, 29, 28) {real, imag} */,
  {32'hbf9a9446, 32'h3fe0691d} /* (14, 29, 27) {real, imag} */,
  {32'hbe35ec4e, 32'hbe561716} /* (14, 29, 26) {real, imag} */,
  {32'h404cce03, 32'h3fe47ebc} /* (14, 29, 25) {real, imag} */,
  {32'hc030c8a1, 32'hbf2921ba} /* (14, 29, 24) {real, imag} */,
  {32'hbf8ec073, 32'hbfeefb32} /* (14, 29, 23) {real, imag} */,
  {32'h3f9f7818, 32'h3e11af33} /* (14, 29, 22) {real, imag} */,
  {32'hbe4ddbd1, 32'h3fc7373e} /* (14, 29, 21) {real, imag} */,
  {32'hc018fbd3, 32'h3f9c1815} /* (14, 29, 20) {real, imag} */,
  {32'h400496a0, 32'h3f16156f} /* (14, 29, 19) {real, imag} */,
  {32'h3ee47fda, 32'hbf278543} /* (14, 29, 18) {real, imag} */,
  {32'h4028743d, 32'hc019fc20} /* (14, 29, 17) {real, imag} */,
  {32'h3f0ad788, 32'h3f73a11c} /* (14, 29, 16) {real, imag} */,
  {32'hbf9692d2, 32'h3fc21083} /* (14, 29, 15) {real, imag} */,
  {32'h40315954, 32'hbd1d1a0a} /* (14, 29, 14) {real, imag} */,
  {32'h3e9ab749, 32'hbf64ecd2} /* (14, 29, 13) {real, imag} */,
  {32'hbec7bc38, 32'hbf621bff} /* (14, 29, 12) {real, imag} */,
  {32'h3ef1b9ff, 32'h3dbae815} /* (14, 29, 11) {real, imag} */,
  {32'hbfef2446, 32'h3ffe8695} /* (14, 29, 10) {real, imag} */,
  {32'hbf12abe1, 32'h3f2f6847} /* (14, 29, 9) {real, imag} */,
  {32'h3eb5f92f, 32'hbf9759fe} /* (14, 29, 8) {real, imag} */,
  {32'hbf68e8cd, 32'h403ded2c} /* (14, 29, 7) {real, imag} */,
  {32'h4052fea4, 32'h3dfe4a17} /* (14, 29, 6) {real, imag} */,
  {32'h3ebb7cee, 32'h3f3dd477} /* (14, 29, 5) {real, imag} */,
  {32'hbfc55812, 32'h3d8642c5} /* (14, 29, 4) {real, imag} */,
  {32'hc01a0a64, 32'hbfffe960} /* (14, 29, 3) {real, imag} */,
  {32'h3f8f2d41, 32'hbe1041c2} /* (14, 29, 2) {real, imag} */,
  {32'hbeba672a, 32'h3f945ce4} /* (14, 29, 1) {real, imag} */,
  {32'hbfb24d58, 32'h3fbd1608} /* (14, 29, 0) {real, imag} */,
  {32'hbfcb3a94, 32'h407dc960} /* (14, 28, 31) {real, imag} */,
  {32'h4036aba6, 32'h3fbe0d1f} /* (14, 28, 30) {real, imag} */,
  {32'h4017cfb0, 32'h3f11a96b} /* (14, 28, 29) {real, imag} */,
  {32'h3feeb736, 32'h3e0f7d9b} /* (14, 28, 28) {real, imag} */,
  {32'hbe1a1b53, 32'hbfdf00e0} /* (14, 28, 27) {real, imag} */,
  {32'h3f50fe21, 32'hbffa7f29} /* (14, 28, 26) {real, imag} */,
  {32'hc0588763, 32'h3fd78adf} /* (14, 28, 25) {real, imag} */,
  {32'h3fd3b5b2, 32'hc09ea28c} /* (14, 28, 24) {real, imag} */,
  {32'hbed2c60e, 32'h3f125e67} /* (14, 28, 23) {real, imag} */,
  {32'h3de189af, 32'hc031e200} /* (14, 28, 22) {real, imag} */,
  {32'hbff83b33, 32'h3e449646} /* (14, 28, 21) {real, imag} */,
  {32'h3f74d6ff, 32'hbe0fe423} /* (14, 28, 20) {real, imag} */,
  {32'hc023ada2, 32'h3f4380bc} /* (14, 28, 19) {real, imag} */,
  {32'hbf89dbe1, 32'h3e7c4284} /* (14, 28, 18) {real, imag} */,
  {32'h3fe6f0d9, 32'h3f0b4243} /* (14, 28, 17) {real, imag} */,
  {32'hbf2af7e6, 32'h3e8bf860} /* (14, 28, 16) {real, imag} */,
  {32'h3e16c384, 32'h3f4823d2} /* (14, 28, 15) {real, imag} */,
  {32'hc02ee98d, 32'hbfba2b7d} /* (14, 28, 14) {real, imag} */,
  {32'hbf13b6fc, 32'h3df3c73e} /* (14, 28, 13) {real, imag} */,
  {32'hbf9b8738, 32'hbff83c86} /* (14, 28, 12) {real, imag} */,
  {32'hbf865334, 32'h40267db5} /* (14, 28, 11) {real, imag} */,
  {32'hbd68fa29, 32'h3efec91e} /* (14, 28, 10) {real, imag} */,
  {32'hc02aae93, 32'h3e0e95db} /* (14, 28, 9) {real, imag} */,
  {32'h400d5bcb, 32'hbe3252b3} /* (14, 28, 8) {real, imag} */,
  {32'hbf96d50a, 32'hbf78031d} /* (14, 28, 7) {real, imag} */,
  {32'hbe66b9e0, 32'h3e64b950} /* (14, 28, 6) {real, imag} */,
  {32'h405d63dd, 32'hbf8f3f25} /* (14, 28, 5) {real, imag} */,
  {32'hc05bf039, 32'hc02ea756} /* (14, 28, 4) {real, imag} */,
  {32'h40214a95, 32'hbfae1233} /* (14, 28, 3) {real, imag} */,
  {32'hbbfc783c, 32'hbf3dde7b} /* (14, 28, 2) {real, imag} */,
  {32'hc0013e50, 32'h401328f3} /* (14, 28, 1) {real, imag} */,
  {32'hbf932926, 32'hbf2c38bc} /* (14, 28, 0) {real, imag} */,
  {32'h3edce174, 32'h3d99ec12} /* (14, 27, 31) {real, imag} */,
  {32'hbec92072, 32'h40866939} /* (14, 27, 30) {real, imag} */,
  {32'hbfa94193, 32'h3fea7b29} /* (14, 27, 29) {real, imag} */,
  {32'h3e88fba6, 32'h3e7ec093} /* (14, 27, 28) {real, imag} */,
  {32'hbf9597cc, 32'h3f5a12ea} /* (14, 27, 27) {real, imag} */,
  {32'h3fbfe5cc, 32'hbf986996} /* (14, 27, 26) {real, imag} */,
  {32'hbecd4ade, 32'hbfdba501} /* (14, 27, 25) {real, imag} */,
  {32'hbcd5986e, 32'h3ec82817} /* (14, 27, 24) {real, imag} */,
  {32'hc063cc93, 32'hbfc7dae1} /* (14, 27, 23) {real, imag} */,
  {32'hbf44b7ef, 32'hbe91cfe5} /* (14, 27, 22) {real, imag} */,
  {32'hc02175fe, 32'h40416785} /* (14, 27, 21) {real, imag} */,
  {32'hc023a877, 32'hc0150e4c} /* (14, 27, 20) {real, imag} */,
  {32'h3f2ba5d4, 32'hbf1a306a} /* (14, 27, 19) {real, imag} */,
  {32'h3d348ff9, 32'h3f9d91ef} /* (14, 27, 18) {real, imag} */,
  {32'h3f23bb36, 32'hbef7ef0d} /* (14, 27, 17) {real, imag} */,
  {32'h3f6c4b7b, 32'hbe8ee9cd} /* (14, 27, 16) {real, imag} */,
  {32'h401d2be8, 32'hc03f93ae} /* (14, 27, 15) {real, imag} */,
  {32'hbf153ccb, 32'h3f1145ae} /* (14, 27, 14) {real, imag} */,
  {32'hc0192919, 32'hbfa59d4d} /* (14, 27, 13) {real, imag} */,
  {32'hc0260357, 32'hbffe3de8} /* (14, 27, 12) {real, imag} */,
  {32'h3ebf410c, 32'hbf8b2be5} /* (14, 27, 11) {real, imag} */,
  {32'h400ec146, 32'hbf1bd3b0} /* (14, 27, 10) {real, imag} */,
  {32'hbe1bafa2, 32'h3f59826b} /* (14, 27, 9) {real, imag} */,
  {32'h3fac5c80, 32'hc0050aff} /* (14, 27, 8) {real, imag} */,
  {32'h3fac5b9e, 32'hbe5bbf08} /* (14, 27, 7) {real, imag} */,
  {32'hbeb28631, 32'h3fc8d1f0} /* (14, 27, 6) {real, imag} */,
  {32'hbfa2ce58, 32'h401fec49} /* (14, 27, 5) {real, imag} */,
  {32'h40336357, 32'hbf46bb9c} /* (14, 27, 4) {real, imag} */,
  {32'h3f24f4a0, 32'h3e1b9b32} /* (14, 27, 3) {real, imag} */,
  {32'hbfae68d9, 32'h3e92d6fa} /* (14, 27, 2) {real, imag} */,
  {32'h4025f766, 32'hc01d855f} /* (14, 27, 1) {real, imag} */,
  {32'h3fd57dde, 32'h3ff0a8dd} /* (14, 27, 0) {real, imag} */,
  {32'h3f62760e, 32'h3d472edf} /* (14, 26, 31) {real, imag} */,
  {32'h3f96b4d3, 32'h3fb0256e} /* (14, 26, 30) {real, imag} */,
  {32'hbf877797, 32'hbff827db} /* (14, 26, 29) {real, imag} */,
  {32'h3f386fd8, 32'h3f01b69e} /* (14, 26, 28) {real, imag} */,
  {32'hbe324767, 32'h3ea71695} /* (14, 26, 27) {real, imag} */,
  {32'hc03104da, 32'hbe7aed1d} /* (14, 26, 26) {real, imag} */,
  {32'h3f847d62, 32'hc000d662} /* (14, 26, 25) {real, imag} */,
  {32'h3f8430ca, 32'h3ef4e2c4} /* (14, 26, 24) {real, imag} */,
  {32'hbef2d64b, 32'h3f98548b} /* (14, 26, 23) {real, imag} */,
  {32'h40265984, 32'hbfd3c420} /* (14, 26, 22) {real, imag} */,
  {32'h3fcb8713, 32'hbf1f912b} /* (14, 26, 21) {real, imag} */,
  {32'hbf70af3c, 32'h3f5d32b2} /* (14, 26, 20) {real, imag} */,
  {32'hbe1cf528, 32'h3f0a1d55} /* (14, 26, 19) {real, imag} */,
  {32'hbfe71b60, 32'hc049eb27} /* (14, 26, 18) {real, imag} */,
  {32'hbe619acb, 32'hbf59138f} /* (14, 26, 17) {real, imag} */,
  {32'h4016a967, 32'h3f971649} /* (14, 26, 16) {real, imag} */,
  {32'h3f74e743, 32'hbfb60aab} /* (14, 26, 15) {real, imag} */,
  {32'hbf84fc47, 32'h3f8ae316} /* (14, 26, 14) {real, imag} */,
  {32'hbf9dc677, 32'hbdf1b4dd} /* (14, 26, 13) {real, imag} */,
  {32'h3f2425dc, 32'hbf80dfae} /* (14, 26, 12) {real, imag} */,
  {32'hbf3aff73, 32'hbf91dc31} /* (14, 26, 11) {real, imag} */,
  {32'h3fdca29c, 32'h3f6ca5f4} /* (14, 26, 10) {real, imag} */,
  {32'hbeb4e332, 32'hbf9890ef} /* (14, 26, 9) {real, imag} */,
  {32'h3f917095, 32'hbf33f61a} /* (14, 26, 8) {real, imag} */,
  {32'h3f2a98bf, 32'h3e427b53} /* (14, 26, 7) {real, imag} */,
  {32'hbf07ab44, 32'hbe7cbb6b} /* (14, 26, 6) {real, imag} */,
  {32'h3fbc2390, 32'h3d89fc94} /* (14, 26, 5) {real, imag} */,
  {32'hbf9579f1, 32'hbcc46f32} /* (14, 26, 4) {real, imag} */,
  {32'h3eef35cc, 32'h400a4338} /* (14, 26, 3) {real, imag} */,
  {32'hbfe1e314, 32'h3daca3fc} /* (14, 26, 2) {real, imag} */,
  {32'h3ea3bba3, 32'h3fa76f4e} /* (14, 26, 1) {real, imag} */,
  {32'hbffad8dd, 32'h3fc50e77} /* (14, 26, 0) {real, imag} */,
  {32'hc038a073, 32'h3fcaed3f} /* (14, 25, 31) {real, imag} */,
  {32'h3f8883a8, 32'h3ff6e8d6} /* (14, 25, 30) {real, imag} */,
  {32'h3f8af3c5, 32'h3fc2d666} /* (14, 25, 29) {real, imag} */,
  {32'h3eacaa94, 32'hbea63309} /* (14, 25, 28) {real, imag} */,
  {32'h40039643, 32'hc007c89b} /* (14, 25, 27) {real, imag} */,
  {32'hbfc185c1, 32'h3e26deab} /* (14, 25, 26) {real, imag} */,
  {32'h3f159d4d, 32'h3f66c2d9} /* (14, 25, 25) {real, imag} */,
  {32'hbf34ea51, 32'hbebf6193} /* (14, 25, 24) {real, imag} */,
  {32'hbeeceaac, 32'h3fe3fa7d} /* (14, 25, 23) {real, imag} */,
  {32'h40231683, 32'hbed1c766} /* (14, 25, 22) {real, imag} */,
  {32'h3d07c622, 32'h3f095a84} /* (14, 25, 21) {real, imag} */,
  {32'hbf4604d1, 32'hbdb6b968} /* (14, 25, 20) {real, imag} */,
  {32'h3d11e014, 32'hbf8928a4} /* (14, 25, 19) {real, imag} */,
  {32'hbf11a87b, 32'h3fdd4e2d} /* (14, 25, 18) {real, imag} */,
  {32'hbfbac42a, 32'hbfd6539b} /* (14, 25, 17) {real, imag} */,
  {32'h3eef612a, 32'h3f2899c3} /* (14, 25, 16) {real, imag} */,
  {32'hc0030a72, 32'h3f0c2010} /* (14, 25, 15) {real, imag} */,
  {32'hbe6a8938, 32'h3ee5dfc1} /* (14, 25, 14) {real, imag} */,
  {32'h4033bca6, 32'h3f8bf77c} /* (14, 25, 13) {real, imag} */,
  {32'h3ebd1121, 32'h3c90dced} /* (14, 25, 12) {real, imag} */,
  {32'h402ba77e, 32'hbe89c25f} /* (14, 25, 11) {real, imag} */,
  {32'h3f13cbc0, 32'h3e998aa2} /* (14, 25, 10) {real, imag} */,
  {32'h3e30cf5d, 32'h3fd0bd49} /* (14, 25, 9) {real, imag} */,
  {32'hbe7b02df, 32'h3eda3d97} /* (14, 25, 8) {real, imag} */,
  {32'hc0386d1a, 32'hbf6724cd} /* (14, 25, 7) {real, imag} */,
  {32'hbec92e25, 32'hbfcf55ca} /* (14, 25, 6) {real, imag} */,
  {32'hbf4e208f, 32'h3ff06c34} /* (14, 25, 5) {real, imag} */,
  {32'h3e41be8b, 32'hbf93cef1} /* (14, 25, 4) {real, imag} */,
  {32'hc002b561, 32'h3f5bbbed} /* (14, 25, 3) {real, imag} */,
  {32'h40409320, 32'h40312ef3} /* (14, 25, 2) {real, imag} */,
  {32'h3fab096e, 32'h3f3fd247} /* (14, 25, 1) {real, imag} */,
  {32'hbf3d7b39, 32'h3f804248} /* (14, 25, 0) {real, imag} */,
  {32'h3fbeadf6, 32'hbfddcc89} /* (14, 24, 31) {real, imag} */,
  {32'hc036bd04, 32'h3f2ba0bd} /* (14, 24, 30) {real, imag} */,
  {32'hc002bf6a, 32'h3ed4932f} /* (14, 24, 29) {real, imag} */,
  {32'hbf901748, 32'hbfa30fbf} /* (14, 24, 28) {real, imag} */,
  {32'h3ff83570, 32'hbff24b62} /* (14, 24, 27) {real, imag} */,
  {32'h3e74f7a2, 32'hc03cb7de} /* (14, 24, 26) {real, imag} */,
  {32'h3fba3131, 32'hbfbb1e0e} /* (14, 24, 25) {real, imag} */,
  {32'h3ead3312, 32'hc07a2093} /* (14, 24, 24) {real, imag} */,
  {32'h3f69639c, 32'h3f9613db} /* (14, 24, 23) {real, imag} */,
  {32'hc0074c48, 32'h3f415fba} /* (14, 24, 22) {real, imag} */,
  {32'h3e841ee2, 32'h3f9c6f71} /* (14, 24, 21) {real, imag} */,
  {32'hbfb0c84e, 32'h3fc1e514} /* (14, 24, 20) {real, imag} */,
  {32'hc029fd26, 32'h400a84dd} /* (14, 24, 19) {real, imag} */,
  {32'h3e9ab0ae, 32'h3f72b8f4} /* (14, 24, 18) {real, imag} */,
  {32'hbf2e02e2, 32'hbf7ae7af} /* (14, 24, 17) {real, imag} */,
  {32'h3faa471e, 32'h3d8f1b97} /* (14, 24, 16) {real, imag} */,
  {32'hbf62ee12, 32'h3fc440c5} /* (14, 24, 15) {real, imag} */,
  {32'hbf68108e, 32'hbff41a7d} /* (14, 24, 14) {real, imag} */,
  {32'h4094d11c, 32'hc006a223} /* (14, 24, 13) {real, imag} */,
  {32'hbdd2ebe4, 32'h407b4002} /* (14, 24, 12) {real, imag} */,
  {32'h3f20a9a6, 32'h3fa306b3} /* (14, 24, 11) {real, imag} */,
  {32'h3f577dc6, 32'h40011dcc} /* (14, 24, 10) {real, imag} */,
  {32'h3f23e217, 32'h3fc1c5c8} /* (14, 24, 9) {real, imag} */,
  {32'hc03b380e, 32'h3f9442dd} /* (14, 24, 8) {real, imag} */,
  {32'hbf6d3311, 32'h3f1e1c4e} /* (14, 24, 7) {real, imag} */,
  {32'hbf4584a8, 32'hbf57b428} /* (14, 24, 6) {real, imag} */,
  {32'hbfe8ce88, 32'h3f0ee0c9} /* (14, 24, 5) {real, imag} */,
  {32'h3f446d82, 32'h401bd700} /* (14, 24, 4) {real, imag} */,
  {32'h3f27935f, 32'hbe2bdd32} /* (14, 24, 3) {real, imag} */,
  {32'hbf95d973, 32'hbf7bb9e0} /* (14, 24, 2) {real, imag} */,
  {32'h3ec21586, 32'hbfd84a84} /* (14, 24, 1) {real, imag} */,
  {32'h3f1e5721, 32'hbdc88d38} /* (14, 24, 0) {real, imag} */,
  {32'hbf859edc, 32'hbe334be4} /* (14, 23, 31) {real, imag} */,
  {32'hc00095f2, 32'hbf5faf7f} /* (14, 23, 30) {real, imag} */,
  {32'h3fc4da23, 32'h3f19e898} /* (14, 23, 29) {real, imag} */,
  {32'hc05b12fb, 32'hc001a8c8} /* (14, 23, 28) {real, imag} */,
  {32'hc0085920, 32'hbd7f91af} /* (14, 23, 27) {real, imag} */,
  {32'h401c5e5f, 32'h3f8223b5} /* (14, 23, 26) {real, imag} */,
  {32'h3e485989, 32'h3f983d7a} /* (14, 23, 25) {real, imag} */,
  {32'h3f934fff, 32'h3f58e950} /* (14, 23, 24) {real, imag} */,
  {32'hbf4927c7, 32'hbfabd8fd} /* (14, 23, 23) {real, imag} */,
  {32'h3f968033, 32'hc073aeb7} /* (14, 23, 22) {real, imag} */,
  {32'hbf6a85dd, 32'hbfc11ef2} /* (14, 23, 21) {real, imag} */,
  {32'hbf64e0f3, 32'hbf41bff8} /* (14, 23, 20) {real, imag} */,
  {32'h3c3cefc3, 32'hbeb6e0a6} /* (14, 23, 19) {real, imag} */,
  {32'hbee1d024, 32'h3eaa2cb0} /* (14, 23, 18) {real, imag} */,
  {32'h3f41d606, 32'h3e9261e0} /* (14, 23, 17) {real, imag} */,
  {32'hbef4d866, 32'hc0062631} /* (14, 23, 16) {real, imag} */,
  {32'h3fc37955, 32'hbfb6017d} /* (14, 23, 15) {real, imag} */,
  {32'h40027d02, 32'hbf1ded62} /* (14, 23, 14) {real, imag} */,
  {32'h3faec888, 32'hbf23bdba} /* (14, 23, 13) {real, imag} */,
  {32'h3e402d55, 32'hbf8ec9bd} /* (14, 23, 12) {real, imag} */,
  {32'hbfadb98c, 32'h3e273981} /* (14, 23, 11) {real, imag} */,
  {32'hbf622f3e, 32'hbf4148f9} /* (14, 23, 10) {real, imag} */,
  {32'hbf07e7f4, 32'h3f9355d9} /* (14, 23, 9) {real, imag} */,
  {32'h3e2bb97a, 32'h40406c70} /* (14, 23, 8) {real, imag} */,
  {32'h4010e302, 32'hbf83db31} /* (14, 23, 7) {real, imag} */,
  {32'h3f81aee7, 32'h3f006b68} /* (14, 23, 6) {real, imag} */,
  {32'h400efd5e, 32'h3f4a68d3} /* (14, 23, 5) {real, imag} */,
  {32'h400c39a6, 32'h3ea0a593} /* (14, 23, 4) {real, imag} */,
  {32'hc017fd09, 32'h3f8fcc75} /* (14, 23, 3) {real, imag} */,
  {32'hbeb684a2, 32'h40462097} /* (14, 23, 2) {real, imag} */,
  {32'h3f7ece34, 32'h3f5fdade} /* (14, 23, 1) {real, imag} */,
  {32'hbf565ad7, 32'h3fdc73b9} /* (14, 23, 0) {real, imag} */,
  {32'hbe9e16b1, 32'hbe8ce1f2} /* (14, 22, 31) {real, imag} */,
  {32'hbe9b6216, 32'hbe9d8aa6} /* (14, 22, 30) {real, imag} */,
  {32'hbdb80f39, 32'hc0099f5a} /* (14, 22, 29) {real, imag} */,
  {32'hbfa3ebdb, 32'h3faaf527} /* (14, 22, 28) {real, imag} */,
  {32'h3ff7aefd, 32'h3ed7d140} /* (14, 22, 27) {real, imag} */,
  {32'h3f9504e8, 32'h40133d10} /* (14, 22, 26) {real, imag} */,
  {32'hbff7c681, 32'h3fa5dded} /* (14, 22, 25) {real, imag} */,
  {32'h3f37a133, 32'h3ee53a8e} /* (14, 22, 24) {real, imag} */,
  {32'h3f496009, 32'h3f2120b3} /* (14, 22, 23) {real, imag} */,
  {32'h3f99d184, 32'h3f746caa} /* (14, 22, 22) {real, imag} */,
  {32'h3f9cc8cf, 32'h40a08d91} /* (14, 22, 21) {real, imag} */,
  {32'h3f9af22f, 32'h3fb9df1a} /* (14, 22, 20) {real, imag} */,
  {32'h404271b4, 32'hbc58cc69} /* (14, 22, 19) {real, imag} */,
  {32'h3db75319, 32'hbf53073d} /* (14, 22, 18) {real, imag} */,
  {32'hbda68e2c, 32'h3f897884} /* (14, 22, 17) {real, imag} */,
  {32'h3fea7ea9, 32'h3e37e70c} /* (14, 22, 16) {real, imag} */,
  {32'h3f6edf34, 32'hbfaab0d6} /* (14, 22, 15) {real, imag} */,
  {32'h3fb3ac65, 32'hbf46a95e} /* (14, 22, 14) {real, imag} */,
  {32'h3e8eedaa, 32'hbf4806ef} /* (14, 22, 13) {real, imag} */,
  {32'h4058f1e2, 32'h3ebc1501} /* (14, 22, 12) {real, imag} */,
  {32'h3ffa1a8d, 32'hbfa80f6b} /* (14, 22, 11) {real, imag} */,
  {32'hc02367d5, 32'h3faacd54} /* (14, 22, 10) {real, imag} */,
  {32'h3fad402d, 32'hbe8a03cc} /* (14, 22, 9) {real, imag} */,
  {32'hc012b02e, 32'h3de4ec57} /* (14, 22, 8) {real, imag} */,
  {32'h3fbbf9ec, 32'hbfabc9a1} /* (14, 22, 7) {real, imag} */,
  {32'h3e1e1f1a, 32'hbf8c7cd9} /* (14, 22, 6) {real, imag} */,
  {32'hc024e275, 32'h3e9cc57a} /* (14, 22, 5) {real, imag} */,
  {32'hc06cd0d3, 32'h3f1a0655} /* (14, 22, 4) {real, imag} */,
  {32'hbf00cf44, 32'h3e53d251} /* (14, 22, 3) {real, imag} */,
  {32'h400fc1a6, 32'hbfc90fe6} /* (14, 22, 2) {real, imag} */,
  {32'h4024e3e8, 32'h3f6b6b79} /* (14, 22, 1) {real, imag} */,
  {32'h3fbfd123, 32'h3fafaa60} /* (14, 22, 0) {real, imag} */,
  {32'h400ed8a8, 32'h400e393e} /* (14, 21, 31) {real, imag} */,
  {32'hbf67382d, 32'hbe55bf44} /* (14, 21, 30) {real, imag} */,
  {32'h4038de62, 32'hc0162163} /* (14, 21, 29) {real, imag} */,
  {32'h400a6086, 32'h402e1de9} /* (14, 21, 28) {real, imag} */,
  {32'h4058099e, 32'hc014aad3} /* (14, 21, 27) {real, imag} */,
  {32'h3f7edcae, 32'h3e51b83f} /* (14, 21, 26) {real, imag} */,
  {32'h3efb5458, 32'hbfdd6ad6} /* (14, 21, 25) {real, imag} */,
  {32'h406582cc, 32'hbf066a8d} /* (14, 21, 24) {real, imag} */,
  {32'hbf2027f5, 32'h3fcd198f} /* (14, 21, 23) {real, imag} */,
  {32'hc03c613a, 32'h403bc71f} /* (14, 21, 22) {real, imag} */,
  {32'h401d05e5, 32'hbf411d73} /* (14, 21, 21) {real, imag} */,
  {32'hbf01056d, 32'h3d323af9} /* (14, 21, 20) {real, imag} */,
  {32'h3f5564ca, 32'hc01a3ab0} /* (14, 21, 19) {real, imag} */,
  {32'hbfe91475, 32'h40514a68} /* (14, 21, 18) {real, imag} */,
  {32'h40056fa7, 32'hbf667795} /* (14, 21, 17) {real, imag} */,
  {32'h3e11e4ec, 32'hbfd7c304} /* (14, 21, 16) {real, imag} */,
  {32'hc022a286, 32'h3f2ed7d0} /* (14, 21, 15) {real, imag} */,
  {32'h4038e1ad, 32'hbfc6089a} /* (14, 21, 14) {real, imag} */,
  {32'hc00033ed, 32'hc08b6964} /* (14, 21, 13) {real, imag} */,
  {32'h4003f188, 32'h400edd88} /* (14, 21, 12) {real, imag} */,
  {32'hbfd29562, 32'h3e694d6b} /* (14, 21, 11) {real, imag} */,
  {32'h40789ab1, 32'hbf95e2ae} /* (14, 21, 10) {real, imag} */,
  {32'h3e0aa6b4, 32'hbe297a35} /* (14, 21, 9) {real, imag} */,
  {32'hbceffc39, 32'hc007aebb} /* (14, 21, 8) {real, imag} */,
  {32'hbec3225d, 32'h3f54aecd} /* (14, 21, 7) {real, imag} */,
  {32'h3e407d30, 32'hbfbb4752} /* (14, 21, 6) {real, imag} */,
  {32'hbffb0c69, 32'hbea967ef} /* (14, 21, 5) {real, imag} */,
  {32'h3b9cd32e, 32'h3fe17ae7} /* (14, 21, 4) {real, imag} */,
  {32'hbfa14cce, 32'h3e8fd4ad} /* (14, 21, 3) {real, imag} */,
  {32'h3ea7c99e, 32'hc00d4c46} /* (14, 21, 2) {real, imag} */,
  {32'h3fdd552f, 32'hbf4669d4} /* (14, 21, 1) {real, imag} */,
  {32'hbf0464db, 32'hbfb06139} /* (14, 21, 0) {real, imag} */,
  {32'hbf72e530, 32'hbf1a0a2f} /* (14, 20, 31) {real, imag} */,
  {32'h40104f75, 32'hbf85b21b} /* (14, 20, 30) {real, imag} */,
  {32'hbfd8eaec, 32'hbf971fe7} /* (14, 20, 29) {real, imag} */,
  {32'h3ee56289, 32'hbf901cc3} /* (14, 20, 28) {real, imag} */,
  {32'hc070ffa2, 32'h400b03d0} /* (14, 20, 27) {real, imag} */,
  {32'hbf7b8989, 32'h3f0087dd} /* (14, 20, 26) {real, imag} */,
  {32'hc000dc34, 32'h3ef7bc6b} /* (14, 20, 25) {real, imag} */,
  {32'hbfb2d4a4, 32'h3fa1886d} /* (14, 20, 24) {real, imag} */,
  {32'hbf9e5f45, 32'hbe4d765b} /* (14, 20, 23) {real, imag} */,
  {32'h3f79de28, 32'h3fd5495f} /* (14, 20, 22) {real, imag} */,
  {32'hc0bf2a67, 32'hbf724dcc} /* (14, 20, 21) {real, imag} */,
  {32'h3fcd3eb5, 32'hbfac9755} /* (14, 20, 20) {real, imag} */,
  {32'h3f33dbea, 32'hbedfd44d} /* (14, 20, 19) {real, imag} */,
  {32'hbfd9de1e, 32'hbf61a66e} /* (14, 20, 18) {real, imag} */,
  {32'h4048c396, 32'hbf2cf768} /* (14, 20, 17) {real, imag} */,
  {32'hbd524f4d, 32'hbf8092ec} /* (14, 20, 16) {real, imag} */,
  {32'hbed2113c, 32'hbdf1f671} /* (14, 20, 15) {real, imag} */,
  {32'h3e75edd3, 32'h400222fc} /* (14, 20, 14) {real, imag} */,
  {32'h3f20afac, 32'h3e691261} /* (14, 20, 13) {real, imag} */,
  {32'h3fd6c01f, 32'hbfa22fb1} /* (14, 20, 12) {real, imag} */,
  {32'h3f14fed8, 32'h402e5561} /* (14, 20, 11) {real, imag} */,
  {32'hc0517044, 32'h404e6652} /* (14, 20, 10) {real, imag} */,
  {32'h3fb8e4b2, 32'hc00c2a19} /* (14, 20, 9) {real, imag} */,
  {32'h4020b955, 32'h3cc04e8d} /* (14, 20, 8) {real, imag} */,
  {32'h401c04af, 32'h4023f99c} /* (14, 20, 7) {real, imag} */,
  {32'h3e35034a, 32'h3e310f4f} /* (14, 20, 6) {real, imag} */,
  {32'hbfb4bcbf, 32'h401951c4} /* (14, 20, 5) {real, imag} */,
  {32'hc02d08e6, 32'h3fc1468b} /* (14, 20, 4) {real, imag} */,
  {32'h3fc635b0, 32'hbe81655e} /* (14, 20, 3) {real, imag} */,
  {32'hbfc36013, 32'h3f2365a3} /* (14, 20, 2) {real, imag} */,
  {32'h3f33b336, 32'hbf76d34c} /* (14, 20, 1) {real, imag} */,
  {32'h3fb947a7, 32'h3df45269} /* (14, 20, 0) {real, imag} */,
  {32'h3f60f38c, 32'h3f9c2014} /* (14, 19, 31) {real, imag} */,
  {32'hc000f17d, 32'hbcf480f1} /* (14, 19, 30) {real, imag} */,
  {32'hbfec6bfa, 32'hc003b1e2} /* (14, 19, 29) {real, imag} */,
  {32'h3fb27894, 32'hbebc306e} /* (14, 19, 28) {real, imag} */,
  {32'h3f27a967, 32'hbfe0372a} /* (14, 19, 27) {real, imag} */,
  {32'hc023c6e3, 32'hc029bdf6} /* (14, 19, 26) {real, imag} */,
  {32'hbfac1801, 32'hbed99ffb} /* (14, 19, 25) {real, imag} */,
  {32'h400394b3, 32'hc007eecb} /* (14, 19, 24) {real, imag} */,
  {32'h3f007dd5, 32'h3ff27535} /* (14, 19, 23) {real, imag} */,
  {32'h3ee04eb6, 32'hbfea3553} /* (14, 19, 22) {real, imag} */,
  {32'hc00ba7fa, 32'hbf6a5c07} /* (14, 19, 21) {real, imag} */,
  {32'hc03ef542, 32'hc00b5aeb} /* (14, 19, 20) {real, imag} */,
  {32'h400403eb, 32'hbf2c7d69} /* (14, 19, 19) {real, imag} */,
  {32'h4024d21b, 32'hbfadf3f9} /* (14, 19, 18) {real, imag} */,
  {32'h3f8a2e70, 32'h3e414f59} /* (14, 19, 17) {real, imag} */,
  {32'hbfebf84e, 32'h3f82f440} /* (14, 19, 16) {real, imag} */,
  {32'h3f89af47, 32'hbf6b9d69} /* (14, 19, 15) {real, imag} */,
  {32'hbff9a52c, 32'hbebeca9e} /* (14, 19, 14) {real, imag} */,
  {32'hc034ed86, 32'h3efbef07} /* (14, 19, 13) {real, imag} */,
  {32'hbf161f8e, 32'hbdee962e} /* (14, 19, 12) {real, imag} */,
  {32'hbe2f9bbd, 32'h3ff828d2} /* (14, 19, 11) {real, imag} */,
  {32'h3f6ee650, 32'hbd4f1177} /* (14, 19, 10) {real, imag} */,
  {32'h3d8c2b2c, 32'h3f3d9c91} /* (14, 19, 9) {real, imag} */,
  {32'hbf32a31e, 32'h3fc09f08} /* (14, 19, 8) {real, imag} */,
  {32'hbfdd94fb, 32'hbfc638e0} /* (14, 19, 7) {real, imag} */,
  {32'h3fd016fa, 32'h3fda72bc} /* (14, 19, 6) {real, imag} */,
  {32'hbf1f78ca, 32'h3fb118a4} /* (14, 19, 5) {real, imag} */,
  {32'h3e3bd225, 32'h3f9a90f0} /* (14, 19, 4) {real, imag} */,
  {32'h3f805452, 32'hbf395b9d} /* (14, 19, 3) {real, imag} */,
  {32'hbeb32683, 32'h3bddffcc} /* (14, 19, 2) {real, imag} */,
  {32'hbff3d768, 32'hbf2ede0c} /* (14, 19, 1) {real, imag} */,
  {32'hbff547f6, 32'h3fe55025} /* (14, 19, 0) {real, imag} */,
  {32'h3e17d4e6, 32'hbf907715} /* (14, 18, 31) {real, imag} */,
  {32'h3e26f9a2, 32'h3f16b42e} /* (14, 18, 30) {real, imag} */,
  {32'h3e450a0c, 32'h3ff6d351} /* (14, 18, 29) {real, imag} */,
  {32'hbe8d3c34, 32'hbf4a5422} /* (14, 18, 28) {real, imag} */,
  {32'h3e400aa6, 32'h40035be6} /* (14, 18, 27) {real, imag} */,
  {32'h3f4dcd45, 32'hbea6787f} /* (14, 18, 26) {real, imag} */,
  {32'h400e5de7, 32'hbf824f8e} /* (14, 18, 25) {real, imag} */,
  {32'h3f09ddee, 32'hbf296cff} /* (14, 18, 24) {real, imag} */,
  {32'hc07882b6, 32'h402e269a} /* (14, 18, 23) {real, imag} */,
  {32'h4063fc87, 32'h3eadc08b} /* (14, 18, 22) {real, imag} */,
  {32'h400c2994, 32'hbe203568} /* (14, 18, 21) {real, imag} */,
  {32'h3fd1118c, 32'hc02dc919} /* (14, 18, 20) {real, imag} */,
  {32'h3fe19ce5, 32'h402a94a0} /* (14, 18, 19) {real, imag} */,
  {32'h3ef3b773, 32'hbf12afde} /* (14, 18, 18) {real, imag} */,
  {32'h3ef3e47a, 32'hbf811ae3} /* (14, 18, 17) {real, imag} */,
  {32'h3fb6a584, 32'h3e963dc6} /* (14, 18, 16) {real, imag} */,
  {32'h3f5c4240, 32'h3f3f7537} /* (14, 18, 15) {real, imag} */,
  {32'hbfc686a2, 32'h3f6a505e} /* (14, 18, 14) {real, imag} */,
  {32'hc0507069, 32'hc00f9dd8} /* (14, 18, 13) {real, imag} */,
  {32'hc02cfb50, 32'h402518e2} /* (14, 18, 12) {real, imag} */,
  {32'hbf04c868, 32'h402365a1} /* (14, 18, 11) {real, imag} */,
  {32'hc026ade1, 32'h3f09edfb} /* (14, 18, 10) {real, imag} */,
  {32'hbfceb65f, 32'hbe322770} /* (14, 18, 9) {real, imag} */,
  {32'hbe41bcb6, 32'h3f161530} /* (14, 18, 8) {real, imag} */,
  {32'hbfbc2ad3, 32'hbecfe114} /* (14, 18, 7) {real, imag} */,
  {32'hbfc5d1ed, 32'hbf362b77} /* (14, 18, 6) {real, imag} */,
  {32'hbf32a698, 32'h3cfabfb0} /* (14, 18, 5) {real, imag} */,
  {32'h40274549, 32'hbf521645} /* (14, 18, 4) {real, imag} */,
  {32'hbf4260d3, 32'hbf84f40c} /* (14, 18, 3) {real, imag} */,
  {32'h3f8a3318, 32'hbf216cdb} /* (14, 18, 2) {real, imag} */,
  {32'hbde11275, 32'hbfdf079e} /* (14, 18, 1) {real, imag} */,
  {32'hbf01228a, 32'hbf08ae7b} /* (14, 18, 0) {real, imag} */,
  {32'hbfb60dbd, 32'h3e6bf1cf} /* (14, 17, 31) {real, imag} */,
  {32'hbf576529, 32'hbf12a7c3} /* (14, 17, 30) {real, imag} */,
  {32'h3f323739, 32'hbe87fdfd} /* (14, 17, 29) {real, imag} */,
  {32'hbfbbdd4b, 32'hbf5f10ca} /* (14, 17, 28) {real, imag} */,
  {32'h3eea52bb, 32'hbf5677e5} /* (14, 17, 27) {real, imag} */,
  {32'hbf15e6bf, 32'h3d6a4dbb} /* (14, 17, 26) {real, imag} */,
  {32'hbf95d5dd, 32'h3f959a77} /* (14, 17, 25) {real, imag} */,
  {32'h3f47bf98, 32'hbf45cd01} /* (14, 17, 24) {real, imag} */,
  {32'h40246d28, 32'hbfbd039a} /* (14, 17, 23) {real, imag} */,
  {32'h404450bf, 32'hbebd4c3d} /* (14, 17, 22) {real, imag} */,
  {32'hbfe1c515, 32'h3f7c51a8} /* (14, 17, 21) {real, imag} */,
  {32'hbf8d122b, 32'h40a1b7cd} /* (14, 17, 20) {real, imag} */,
  {32'hbfef74ed, 32'hbe534d13} /* (14, 17, 19) {real, imag} */,
  {32'hc0063375, 32'h403ad93e} /* (14, 17, 18) {real, imag} */,
  {32'hc00b7dd9, 32'h3f7eb10b} /* (14, 17, 17) {real, imag} */,
  {32'h3f07586a, 32'h3f82c1fc} /* (14, 17, 16) {real, imag} */,
  {32'hbf177b39, 32'hbfadc64f} /* (14, 17, 15) {real, imag} */,
  {32'h3f5b4391, 32'h3ecc9cce} /* (14, 17, 14) {real, imag} */,
  {32'hbf6c90e4, 32'h4032b94a} /* (14, 17, 13) {real, imag} */,
  {32'hbf8782f4, 32'hbf8d7d00} /* (14, 17, 12) {real, imag} */,
  {32'hbfb0559d, 32'hbd16d2ec} /* (14, 17, 11) {real, imag} */,
  {32'h3fd22c39, 32'hbfb43836} /* (14, 17, 10) {real, imag} */,
  {32'h3f39a58a, 32'h3f960b58} /* (14, 17, 9) {real, imag} */,
  {32'h3f6e60ad, 32'h3fb4ce6b} /* (14, 17, 8) {real, imag} */,
  {32'hbfd7bcaf, 32'h3e5a3b65} /* (14, 17, 7) {real, imag} */,
  {32'h3f84ec83, 32'h40272f75} /* (14, 17, 6) {real, imag} */,
  {32'hbd8e4fd8, 32'h3f1a3193} /* (14, 17, 5) {real, imag} */,
  {32'h3f43b80a, 32'hc0365a70} /* (14, 17, 4) {real, imag} */,
  {32'h3fff0af1, 32'hbe8ca0d1} /* (14, 17, 3) {real, imag} */,
  {32'h3f1cc71a, 32'h3f2926f8} /* (14, 17, 2) {real, imag} */,
  {32'h3ef0f618, 32'hbee8b31d} /* (14, 17, 1) {real, imag} */,
  {32'h3f0541e6, 32'hbe1d72f8} /* (14, 17, 0) {real, imag} */,
  {32'hbf03a6dd, 32'h3dedb29f} /* (14, 16, 31) {real, imag} */,
  {32'hbf072aff, 32'hbf48558c} /* (14, 16, 30) {real, imag} */,
  {32'hbed63e41, 32'hbf3b24c0} /* (14, 16, 29) {real, imag} */,
  {32'h3f5ef34b, 32'h3f88c775} /* (14, 16, 28) {real, imag} */,
  {32'hbec58124, 32'h3f890f4a} /* (14, 16, 27) {real, imag} */,
  {32'hbfb59547, 32'h3fa39ff0} /* (14, 16, 26) {real, imag} */,
  {32'h3f83af5e, 32'hbfb15bb5} /* (14, 16, 25) {real, imag} */,
  {32'hbf426a4b, 32'hbf1eded6} /* (14, 16, 24) {real, imag} */,
  {32'h3f8578be, 32'h3f7c4d6a} /* (14, 16, 23) {real, imag} */,
  {32'h3f6d77bf, 32'hbfa84976} /* (14, 16, 22) {real, imag} */,
  {32'hbd7d0712, 32'hbeb870fe} /* (14, 16, 21) {real, imag} */,
  {32'h3fa9e4c2, 32'h3d9cd32a} /* (14, 16, 20) {real, imag} */,
  {32'h3ff182cd, 32'h40020e37} /* (14, 16, 19) {real, imag} */,
  {32'hbfd37524, 32'h3fa5bf81} /* (14, 16, 18) {real, imag} */,
  {32'hbe6656c2, 32'hbeb6d73c} /* (14, 16, 17) {real, imag} */,
  {32'h3dbbde8d, 32'hbf464312} /* (14, 16, 16) {real, imag} */,
  {32'h3d9fcff8, 32'h3ee6d48a} /* (14, 16, 15) {real, imag} */,
  {32'h3f0d301f, 32'hbef8ead5} /* (14, 16, 14) {real, imag} */,
  {32'hbfb71ac9, 32'hbf5fe7db} /* (14, 16, 13) {real, imag} */,
  {32'h3f4d2559, 32'h3f0b62de} /* (14, 16, 12) {real, imag} */,
  {32'hbef1ac77, 32'hbdadd828} /* (14, 16, 11) {real, imag} */,
  {32'hbe5914c3, 32'hc05901c4} /* (14, 16, 10) {real, imag} */,
  {32'h3eb46a87, 32'hbf72180f} /* (14, 16, 9) {real, imag} */,
  {32'hbedd48f0, 32'h3ee649c6} /* (14, 16, 8) {real, imag} */,
  {32'hbf02412e, 32'hbe9019c9} /* (14, 16, 7) {real, imag} */,
  {32'hbe3e1168, 32'h3f0d9ea1} /* (14, 16, 6) {real, imag} */,
  {32'h3fabfea1, 32'h3f8a90d3} /* (14, 16, 5) {real, imag} */,
  {32'h3f2c963d, 32'h3d69c942} /* (14, 16, 4) {real, imag} */,
  {32'h3f4a98a2, 32'hbf17edab} /* (14, 16, 3) {real, imag} */,
  {32'hbf8e311a, 32'h3fea6114} /* (14, 16, 2) {real, imag} */,
  {32'h3e11f954, 32'hc01a63ef} /* (14, 16, 1) {real, imag} */,
  {32'h3ed49494, 32'h3ea8fb26} /* (14, 16, 0) {real, imag} */,
  {32'hbf5f6e48, 32'hc0082c39} /* (14, 15, 31) {real, imag} */,
  {32'h3caf2f6e, 32'hbe8f3e45} /* (14, 15, 30) {real, imag} */,
  {32'h3fb0f17d, 32'hbf90cc4f} /* (14, 15, 29) {real, imag} */,
  {32'hbfe7146e, 32'h3e107643} /* (14, 15, 28) {real, imag} */,
  {32'h3f6b07e4, 32'hbe6c8fe6} /* (14, 15, 27) {real, imag} */,
  {32'hbfa3fc1c, 32'h3ec698d4} /* (14, 15, 26) {real, imag} */,
  {32'h3f3c2923, 32'h3f54d46f} /* (14, 15, 25) {real, imag} */,
  {32'hbfaf0778, 32'hbf74226b} /* (14, 15, 24) {real, imag} */,
  {32'hbeda0937, 32'h3fb72050} /* (14, 15, 23) {real, imag} */,
  {32'h403214b1, 32'hc00d01a3} /* (14, 15, 22) {real, imag} */,
  {32'h3fed1062, 32'h3fe36b19} /* (14, 15, 21) {real, imag} */,
  {32'h3eac0723, 32'hbf985685} /* (14, 15, 20) {real, imag} */,
  {32'hbfb75ece, 32'h3f4c2615} /* (14, 15, 19) {real, imag} */,
  {32'h3ec7d260, 32'h3e710a51} /* (14, 15, 18) {real, imag} */,
  {32'h3e590001, 32'h3eeb3180} /* (14, 15, 17) {real, imag} */,
  {32'hbe9dbf05, 32'hc00e840d} /* (14, 15, 16) {real, imag} */,
  {32'h3f7490b2, 32'hbfb08eef} /* (14, 15, 15) {real, imag} */,
  {32'h3f6c6a91, 32'hc011188f} /* (14, 15, 14) {real, imag} */,
  {32'hbffc3c23, 32'h402172e6} /* (14, 15, 13) {real, imag} */,
  {32'hbfd4c7b2, 32'hbe4e03be} /* (14, 15, 12) {real, imag} */,
  {32'hbfe788d8, 32'hc02aa2a3} /* (14, 15, 11) {real, imag} */,
  {32'h3fc0d96b, 32'hbe60f8db} /* (14, 15, 10) {real, imag} */,
  {32'h3f58dd14, 32'hbe775b8d} /* (14, 15, 9) {real, imag} */,
  {32'hbeff0a7f, 32'h404fbf86} /* (14, 15, 8) {real, imag} */,
  {32'h3f4bab99, 32'hbd2e1abf} /* (14, 15, 7) {real, imag} */,
  {32'h401466f6, 32'hbff22070} /* (14, 15, 6) {real, imag} */,
  {32'hbebe1fcb, 32'hbe48df82} /* (14, 15, 5) {real, imag} */,
  {32'h3f9e89a6, 32'h3fd7d600} /* (14, 15, 4) {real, imag} */,
  {32'h3f26fd54, 32'h3e679da7} /* (14, 15, 3) {real, imag} */,
  {32'h3e8d252e, 32'h401200c8} /* (14, 15, 2) {real, imag} */,
  {32'h3fa64cee, 32'hbf1982f1} /* (14, 15, 1) {real, imag} */,
  {32'hbfe197d9, 32'hbf486185} /* (14, 15, 0) {real, imag} */,
  {32'h3db4b031, 32'h3f948356} /* (14, 14, 31) {real, imag} */,
  {32'hbef109aa, 32'hbfcfe955} /* (14, 14, 30) {real, imag} */,
  {32'hbe87f262, 32'h3f1a2ac5} /* (14, 14, 29) {real, imag} */,
  {32'h3f2f675f, 32'hbe8b4d10} /* (14, 14, 28) {real, imag} */,
  {32'h4031420c, 32'h4000c7a3} /* (14, 14, 27) {real, imag} */,
  {32'h3ee175be, 32'hbfe12760} /* (14, 14, 26) {real, imag} */,
  {32'hbf078ac4, 32'hbae048cd} /* (14, 14, 25) {real, imag} */,
  {32'h3feec533, 32'hbfa9eeb2} /* (14, 14, 24) {real, imag} */,
  {32'hbfe815fc, 32'hc055a19f} /* (14, 14, 23) {real, imag} */,
  {32'hbf58954a, 32'h3e62f968} /* (14, 14, 22) {real, imag} */,
  {32'h3fc298b1, 32'hbe8ecee2} /* (14, 14, 21) {real, imag} */,
  {32'hbf1c9fb0, 32'hc0011038} /* (14, 14, 20) {real, imag} */,
  {32'h3e133717, 32'h3f4eae4f} /* (14, 14, 19) {real, imag} */,
  {32'h3fe3425d, 32'h3f5f9600} /* (14, 14, 18) {real, imag} */,
  {32'h3f45dd1e, 32'h3f8985d9} /* (14, 14, 17) {real, imag} */,
  {32'hbf27525e, 32'hbff6d98e} /* (14, 14, 16) {real, imag} */,
  {32'h3e8a5624, 32'hbf1cc200} /* (14, 14, 15) {real, imag} */,
  {32'hbe8964a5, 32'hbfc66ce5} /* (14, 14, 14) {real, imag} */,
  {32'h3fa15b45, 32'hc041b9b1} /* (14, 14, 13) {real, imag} */,
  {32'h3f0e3cf2, 32'hbf9130cd} /* (14, 14, 12) {real, imag} */,
  {32'h400a13e5, 32'hbfd17df6} /* (14, 14, 11) {real, imag} */,
  {32'h3e57f7ec, 32'h3f0bb0e9} /* (14, 14, 10) {real, imag} */,
  {32'h3e70a583, 32'h40710eda} /* (14, 14, 9) {real, imag} */,
  {32'hc01f8691, 32'h3f370cf6} /* (14, 14, 8) {real, imag} */,
  {32'hbf3245fd, 32'hbf7a93c0} /* (14, 14, 7) {real, imag} */,
  {32'h403503c6, 32'h3f807330} /* (14, 14, 6) {real, imag} */,
  {32'h3f138d90, 32'hbf84f39a} /* (14, 14, 5) {real, imag} */,
  {32'hbf534bd9, 32'h3fe19a1e} /* (14, 14, 4) {real, imag} */,
  {32'hbf81023a, 32'hbfaadb91} /* (14, 14, 3) {real, imag} */,
  {32'h3f3f5514, 32'h3e8c4fd5} /* (14, 14, 2) {real, imag} */,
  {32'h3f58f2ed, 32'hbf1a8d91} /* (14, 14, 1) {real, imag} */,
  {32'hbd8cf1a1, 32'hbe1e999f} /* (14, 14, 0) {real, imag} */,
  {32'h3f385e0d, 32'hbda42ae1} /* (14, 13, 31) {real, imag} */,
  {32'h3fde86b1, 32'h3ff30754} /* (14, 13, 30) {real, imag} */,
  {32'hbefd8afe, 32'hbdcf3266} /* (14, 13, 29) {real, imag} */,
  {32'h3dfd3612, 32'hbfa82269} /* (14, 13, 28) {real, imag} */,
  {32'h3f6b71e2, 32'h3f0aa162} /* (14, 13, 27) {real, imag} */,
  {32'hbf988220, 32'hc00cb3a7} /* (14, 13, 26) {real, imag} */,
  {32'h3fe89112, 32'hbfb9dda3} /* (14, 13, 25) {real, imag} */,
  {32'hc0202a56, 32'h3db873ef} /* (14, 13, 24) {real, imag} */,
  {32'hbed70a20, 32'h40899333} /* (14, 13, 23) {real, imag} */,
  {32'h406b583a, 32'hbfe019dc} /* (14, 13, 22) {real, imag} */,
  {32'hc0079e30, 32'h3f9549bc} /* (14, 13, 21) {real, imag} */,
  {32'h401ee7c6, 32'hbff23b7f} /* (14, 13, 20) {real, imag} */,
  {32'h3df6b70f, 32'hbf0d42fc} /* (14, 13, 19) {real, imag} */,
  {32'h3e9d2a62, 32'h3f45f0e6} /* (14, 13, 18) {real, imag} */,
  {32'hbf832404, 32'h401c60bc} /* (14, 13, 17) {real, imag} */,
  {32'hbf0ed44d, 32'hbe90eb96} /* (14, 13, 16) {real, imag} */,
  {32'h3ff6fec7, 32'h3f140633} /* (14, 13, 15) {real, imag} */,
  {32'hbfa0edc0, 32'h3f421174} /* (14, 13, 14) {real, imag} */,
  {32'h4010b4e9, 32'hc047921c} /* (14, 13, 13) {real, imag} */,
  {32'h4067c4b5, 32'hbf033f9c} /* (14, 13, 12) {real, imag} */,
  {32'h3f113551, 32'hbfabe13c} /* (14, 13, 11) {real, imag} */,
  {32'hbfbda832, 32'hbe7546aa} /* (14, 13, 10) {real, imag} */,
  {32'hbea17c42, 32'h404f3b60} /* (14, 13, 9) {real, imag} */,
  {32'hbfe70b99, 32'hbf7928fd} /* (14, 13, 8) {real, imag} */,
  {32'hc035c2e4, 32'hbeac0c6c} /* (14, 13, 7) {real, imag} */,
  {32'hbfdcd479, 32'hbf215909} /* (14, 13, 6) {real, imag} */,
  {32'h3fc251ce, 32'hbfa32a23} /* (14, 13, 5) {real, imag} */,
  {32'hbd12dc8e, 32'h3f579859} /* (14, 13, 4) {real, imag} */,
  {32'hbf61fd27, 32'h3f9eb666} /* (14, 13, 3) {real, imag} */,
  {32'hbeb11214, 32'h40148061} /* (14, 13, 2) {real, imag} */,
  {32'h3f094f20, 32'hbd86002c} /* (14, 13, 1) {real, imag} */,
  {32'hc062458e, 32'hbf89a6e8} /* (14, 13, 0) {real, imag} */,
  {32'hbf78086c, 32'hbf9848c1} /* (14, 12, 31) {real, imag} */,
  {32'hbfb3ae27, 32'hbe137bd4} /* (14, 12, 30) {real, imag} */,
  {32'hc0697cac, 32'hbf9580cd} /* (14, 12, 29) {real, imag} */,
  {32'h3fad269d, 32'h40810a9d} /* (14, 12, 28) {real, imag} */,
  {32'h40181399, 32'h3e80898d} /* (14, 12, 27) {real, imag} */,
  {32'hbf95b239, 32'h3feaef01} /* (14, 12, 26) {real, imag} */,
  {32'h3f9951bc, 32'hbd147233} /* (14, 12, 25) {real, imag} */,
  {32'h3f161995, 32'h3f85b3f1} /* (14, 12, 24) {real, imag} */,
  {32'h3f92669a, 32'h4018e40d} /* (14, 12, 23) {real, imag} */,
  {32'h3f5b5715, 32'hc017a4d3} /* (14, 12, 22) {real, imag} */,
  {32'h3f397ab4, 32'hbfd0cfec} /* (14, 12, 21) {real, imag} */,
  {32'hc02418fe, 32'h3fac6c28} /* (14, 12, 20) {real, imag} */,
  {32'hbf4f6896, 32'hbed90862} /* (14, 12, 19) {real, imag} */,
  {32'h3f20de66, 32'hbe8c6c3d} /* (14, 12, 18) {real, imag} */,
  {32'hbe60bcd3, 32'h3e66f59a} /* (14, 12, 17) {real, imag} */,
  {32'hbd66da48, 32'h3fe7ab46} /* (14, 12, 16) {real, imag} */,
  {32'hc026191b, 32'h3fe31f6b} /* (14, 12, 15) {real, imag} */,
  {32'hbf9c5943, 32'hc0969592} /* (14, 12, 14) {real, imag} */,
  {32'hbf9c8e8e, 32'hbe53ee4f} /* (14, 12, 13) {real, imag} */,
  {32'h3f288079, 32'h3f42ae02} /* (14, 12, 12) {real, imag} */,
  {32'hbfc0b2d9, 32'h4010ef99} /* (14, 12, 11) {real, imag} */,
  {32'h40885007, 32'hbf583995} /* (14, 12, 10) {real, imag} */,
  {32'hbf854ce4, 32'h3e2d9eae} /* (14, 12, 9) {real, imag} */,
  {32'hc07eadad, 32'hbf8ef92b} /* (14, 12, 8) {real, imag} */,
  {32'h3fa820a7, 32'hbfd36f33} /* (14, 12, 7) {real, imag} */,
  {32'h3e1c59e6, 32'hbf9eef3c} /* (14, 12, 6) {real, imag} */,
  {32'hc00c0bbf, 32'h3dd1f7ed} /* (14, 12, 5) {real, imag} */,
  {32'h3fef4657, 32'h3def05e5} /* (14, 12, 4) {real, imag} */,
  {32'h3eeb56f8, 32'hbebe1422} /* (14, 12, 3) {real, imag} */,
  {32'hbe69f9cc, 32'hbfb3b7e1} /* (14, 12, 2) {real, imag} */,
  {32'h3f6e5381, 32'hbfc547c2} /* (14, 12, 1) {real, imag} */,
  {32'hbe6051aa, 32'hc053b23b} /* (14, 12, 0) {real, imag} */,
  {32'hbf36f32f, 32'h3f5dc943} /* (14, 11, 31) {real, imag} */,
  {32'hbe65c16c, 32'hbf3b7570} /* (14, 11, 30) {real, imag} */,
  {32'h4009c3d8, 32'h3f6de63c} /* (14, 11, 29) {real, imag} */,
  {32'h3eab734b, 32'hbfb855bf} /* (14, 11, 28) {real, imag} */,
  {32'h3f64db9e, 32'h402edd1b} /* (14, 11, 27) {real, imag} */,
  {32'hbf8c8d7f, 32'hbf29f1bd} /* (14, 11, 26) {real, imag} */,
  {32'hbf2eef27, 32'h3fd47cd1} /* (14, 11, 25) {real, imag} */,
  {32'h3ed40961, 32'h400203f4} /* (14, 11, 24) {real, imag} */,
  {32'hbe034ce1, 32'hbfd90143} /* (14, 11, 23) {real, imag} */,
  {32'h3f2b8ecc, 32'hbec2ccc9} /* (14, 11, 22) {real, imag} */,
  {32'h3fadb7b4, 32'hbfdbe64b} /* (14, 11, 21) {real, imag} */,
  {32'h3f424d8d, 32'h401ad640} /* (14, 11, 20) {real, imag} */,
  {32'hbf353aa5, 32'h40845ef1} /* (14, 11, 19) {real, imag} */,
  {32'h3f657f5c, 32'h40161928} /* (14, 11, 18) {real, imag} */,
  {32'hbf4ab750, 32'hc07aa1d3} /* (14, 11, 17) {real, imag} */,
  {32'hc003979d, 32'h404653c8} /* (14, 11, 16) {real, imag} */,
  {32'hbfce7000, 32'hbf9ff7c2} /* (14, 11, 15) {real, imag} */,
  {32'h3f827e22, 32'hbfe46ab0} /* (14, 11, 14) {real, imag} */,
  {32'h3fb354ff, 32'hc038dc40} /* (14, 11, 13) {real, imag} */,
  {32'h3f2f1b1c, 32'h3f27ecc9} /* (14, 11, 12) {real, imag} */,
  {32'h4086ffd9, 32'hbf79131b} /* (14, 11, 11) {real, imag} */,
  {32'hbe182785, 32'hbedf6d29} /* (14, 11, 10) {real, imag} */,
  {32'hbea51d58, 32'h3f4b51d1} /* (14, 11, 9) {real, imag} */,
  {32'h400931dd, 32'h401c4fb3} /* (14, 11, 8) {real, imag} */,
  {32'h3fbeb044, 32'h3f26e553} /* (14, 11, 7) {real, imag} */,
  {32'h401eda7e, 32'h3eb8cd7a} /* (14, 11, 6) {real, imag} */,
  {32'hbf9df577, 32'hbe43ae0c} /* (14, 11, 5) {real, imag} */,
  {32'hbfa2ba31, 32'hc01ae27f} /* (14, 11, 4) {real, imag} */,
  {32'hbe1f91b3, 32'hbffa2b4d} /* (14, 11, 3) {real, imag} */,
  {32'hbf9eafeb, 32'hc03e80ca} /* (14, 11, 2) {real, imag} */,
  {32'h3d8c16d3, 32'hbcf3e7f6} /* (14, 11, 1) {real, imag} */,
  {32'hbd8a83c6, 32'h3f9a7a33} /* (14, 11, 0) {real, imag} */,
  {32'hbf267017, 32'hbfb14fd8} /* (14, 10, 31) {real, imag} */,
  {32'h402167fa, 32'h3fbd558c} /* (14, 10, 30) {real, imag} */,
  {32'hbf7b3299, 32'hbc982cb9} /* (14, 10, 29) {real, imag} */,
  {32'hbf307d0b, 32'h3f32660e} /* (14, 10, 28) {real, imag} */,
  {32'h3bbaa991, 32'h3f4fd0ab} /* (14, 10, 27) {real, imag} */,
  {32'h4095ff39, 32'h3f06cd2e} /* (14, 10, 26) {real, imag} */,
  {32'h3e81e079, 32'h3e532327} /* (14, 10, 25) {real, imag} */,
  {32'hbe85258e, 32'h3d0d21dc} /* (14, 10, 24) {real, imag} */,
  {32'hbf0190b7, 32'hbf0097c8} /* (14, 10, 23) {real, imag} */,
  {32'hc003228c, 32'hc0458191} /* (14, 10, 22) {real, imag} */,
  {32'hbe17f8f4, 32'hc009e654} /* (14, 10, 21) {real, imag} */,
  {32'h3f2c3df7, 32'h3fbbf155} /* (14, 10, 20) {real, imag} */,
  {32'h404fb919, 32'hbfbd0b17} /* (14, 10, 19) {real, imag} */,
  {32'hbe172c1c, 32'hc0040cf2} /* (14, 10, 18) {real, imag} */,
  {32'hc0423759, 32'h3fb3cc64} /* (14, 10, 17) {real, imag} */,
  {32'hc04c49a8, 32'hbf09c0cd} /* (14, 10, 16) {real, imag} */,
  {32'h3f50a9bb, 32'hbfb8b5f1} /* (14, 10, 15) {real, imag} */,
  {32'hc00a61a0, 32'h403a9329} /* (14, 10, 14) {real, imag} */,
  {32'hbff119ca, 32'hc0a69ace} /* (14, 10, 13) {real, imag} */,
  {32'h3e3dcde6, 32'hbfc0fa02} /* (14, 10, 12) {real, imag} */,
  {32'h3fbcca73, 32'h3f48899d} /* (14, 10, 11) {real, imag} */,
  {32'h407d84bf, 32'h3f18359d} /* (14, 10, 10) {real, imag} */,
  {32'h3e4ec128, 32'hbec861e8} /* (14, 10, 9) {real, imag} */,
  {32'hbfbfe9cd, 32'hbf291346} /* (14, 10, 8) {real, imag} */,
  {32'h4005b5ed, 32'h3f0b3f53} /* (14, 10, 7) {real, imag} */,
  {32'h3fc659a3, 32'hbf5d7cbe} /* (14, 10, 6) {real, imag} */,
  {32'h3f09824c, 32'h3ee1444f} /* (14, 10, 5) {real, imag} */,
  {32'h3e59bef5, 32'hc0085a25} /* (14, 10, 4) {real, imag} */,
  {32'hba614f0d, 32'h3f1981e1} /* (14, 10, 3) {real, imag} */,
  {32'hc0024e07, 32'hbc5bbc6b} /* (14, 10, 2) {real, imag} */,
  {32'hc004c24c, 32'h40381a9d} /* (14, 10, 1) {real, imag} */,
  {32'h401396b3, 32'hbe047c3c} /* (14, 10, 0) {real, imag} */,
  {32'h40019da6, 32'hbf82826b} /* (14, 9, 31) {real, imag} */,
  {32'h3fca9fdf, 32'hbf6dc5b3} /* (14, 9, 30) {real, imag} */,
  {32'hbf6e5df8, 32'h402ef19a} /* (14, 9, 29) {real, imag} */,
  {32'hc08a7887, 32'hbff5f75f} /* (14, 9, 28) {real, imag} */,
  {32'hc05d1e3e, 32'h3fbe6b75} /* (14, 9, 27) {real, imag} */,
  {32'h3fc4fc04, 32'hbf7c3527} /* (14, 9, 26) {real, imag} */,
  {32'h3f2af826, 32'hbe573b91} /* (14, 9, 25) {real, imag} */,
  {32'hbe6ad0ed, 32'hbf9f358d} /* (14, 9, 24) {real, imag} */,
  {32'h3f92f6b9, 32'h3e151908} /* (14, 9, 23) {real, imag} */,
  {32'h4034ac3e, 32'hbfeb6b62} /* (14, 9, 22) {real, imag} */,
  {32'hbfd4ce6e, 32'h3f127c9f} /* (14, 9, 21) {real, imag} */,
  {32'hbf63055a, 32'h3fe82029} /* (14, 9, 20) {real, imag} */,
  {32'h3f37393d, 32'hbfd180d0} /* (14, 9, 19) {real, imag} */,
  {32'hbeb1c269, 32'hbf71d3c5} /* (14, 9, 18) {real, imag} */,
  {32'hbfff5631, 32'h3e8a5e67} /* (14, 9, 17) {real, imag} */,
  {32'h3ffb52fa, 32'hbfec4250} /* (14, 9, 16) {real, imag} */,
  {32'hbe49ed91, 32'hc01d5373} /* (14, 9, 15) {real, imag} */,
  {32'h3fc12456, 32'h40078939} /* (14, 9, 14) {real, imag} */,
  {32'hc016cd8d, 32'hbfeffa74} /* (14, 9, 13) {real, imag} */,
  {32'hbf13aa48, 32'h40393fab} /* (14, 9, 12) {real, imag} */,
  {32'hbe1d8aae, 32'h403fdb17} /* (14, 9, 11) {real, imag} */,
  {32'h400aac15, 32'hbf593572} /* (14, 9, 10) {real, imag} */,
  {32'hbff0ab16, 32'hbf6ae771} /* (14, 9, 9) {real, imag} */,
  {32'h3e14fb4d, 32'h3ffdc5ab} /* (14, 9, 8) {real, imag} */,
  {32'h3f1c3685, 32'hbf83da8d} /* (14, 9, 7) {real, imag} */,
  {32'hbf9a15dc, 32'h3cf48009} /* (14, 9, 6) {real, imag} */,
  {32'h3fac4b67, 32'h3e6bc165} /* (14, 9, 5) {real, imag} */,
  {32'hbfcb4d8f, 32'h3fbe7f6d} /* (14, 9, 4) {real, imag} */,
  {32'hbfc8947d, 32'h3e2ff21b} /* (14, 9, 3) {real, imag} */,
  {32'hbebddb34, 32'hbe027193} /* (14, 9, 2) {real, imag} */,
  {32'hbf4c83f7, 32'hbfbf7f45} /* (14, 9, 1) {real, imag} */,
  {32'h3f7a8384, 32'hbfa368b9} /* (14, 9, 0) {real, imag} */,
  {32'h40263b0e, 32'h403891ed} /* (14, 8, 31) {real, imag} */,
  {32'hbf0b55c6, 32'h3f10120e} /* (14, 8, 30) {real, imag} */,
  {32'hbcf05fdc, 32'hbfe7232d} /* (14, 8, 29) {real, imag} */,
  {32'hbdfca5a7, 32'h3fe29cf3} /* (14, 8, 28) {real, imag} */,
  {32'h3e56062d, 32'hbfcd0117} /* (14, 8, 27) {real, imag} */,
  {32'h3ff9d10f, 32'h3d2e67dd} /* (14, 8, 26) {real, imag} */,
  {32'h3fc808fd, 32'hbff37dfc} /* (14, 8, 25) {real, imag} */,
  {32'h3ee09548, 32'h3ff2f28f} /* (14, 8, 24) {real, imag} */,
  {32'hbf99be02, 32'hc0257be3} /* (14, 8, 23) {real, imag} */,
  {32'hbfde4df7, 32'hbffb9d02} /* (14, 8, 22) {real, imag} */,
  {32'hbed9f408, 32'hbec74ef0} /* (14, 8, 21) {real, imag} */,
  {32'h3ff5c34d, 32'hbffc96f9} /* (14, 8, 20) {real, imag} */,
  {32'hbfcda153, 32'h3ff2eb7c} /* (14, 8, 19) {real, imag} */,
  {32'h40081720, 32'h3d126184} /* (14, 8, 18) {real, imag} */,
  {32'hbe7cbdeb, 32'hbf09d1a6} /* (14, 8, 17) {real, imag} */,
  {32'hc0115996, 32'h3e09ecc3} /* (14, 8, 16) {real, imag} */,
  {32'hbf28e34f, 32'hbf836ae5} /* (14, 8, 15) {real, imag} */,
  {32'hbe999326, 32'h3fd54e71} /* (14, 8, 14) {real, imag} */,
  {32'hbe58597f, 32'h3ffc0592} /* (14, 8, 13) {real, imag} */,
  {32'hbf5fce37, 32'hbfab5030} /* (14, 8, 12) {real, imag} */,
  {32'hc081490a, 32'hbedec9b2} /* (14, 8, 11) {real, imag} */,
  {32'h3f302c78, 32'hbe8becf8} /* (14, 8, 10) {real, imag} */,
  {32'hbfb8972c, 32'hc042cdf6} /* (14, 8, 9) {real, imag} */,
  {32'hc03f4f8d, 32'h3f1887e0} /* (14, 8, 8) {real, imag} */,
  {32'hbf00227d, 32'h3ea79593} /* (14, 8, 7) {real, imag} */,
  {32'hc0099c5a, 32'hbfe98800} /* (14, 8, 6) {real, imag} */,
  {32'hbe688f9c, 32'hbfafe299} /* (14, 8, 5) {real, imag} */,
  {32'hbf8bc52d, 32'hbfa51111} /* (14, 8, 4) {real, imag} */,
  {32'hbe8ee50e, 32'hbf7eb7a4} /* (14, 8, 3) {real, imag} */,
  {32'h3f791b92, 32'h3e1fe80e} /* (14, 8, 2) {real, imag} */,
  {32'h3fd8ea26, 32'hbd14d7d0} /* (14, 8, 1) {real, imag} */,
  {32'hbe232ee2, 32'h3e1e30c9} /* (14, 8, 0) {real, imag} */,
  {32'h3f981c49, 32'hbf43cdfa} /* (14, 7, 31) {real, imag} */,
  {32'hc01f96f7, 32'hbf85d7f5} /* (14, 7, 30) {real, imag} */,
  {32'h3f6a27ad, 32'h3f69266e} /* (14, 7, 29) {real, imag} */,
  {32'h401e4257, 32'hc0664093} /* (14, 7, 28) {real, imag} */,
  {32'hbfc22866, 32'h3fd6fd9f} /* (14, 7, 27) {real, imag} */,
  {32'h3f8ca600, 32'h40265125} /* (14, 7, 26) {real, imag} */,
  {32'hc01a099f, 32'h3f942947} /* (14, 7, 25) {real, imag} */,
  {32'h3f7859d9, 32'hbfd178ab} /* (14, 7, 24) {real, imag} */,
  {32'hbe8f35d0, 32'h3f719118} /* (14, 7, 23) {real, imag} */,
  {32'hbf9e62ff, 32'hc02201af} /* (14, 7, 22) {real, imag} */,
  {32'hbe58e12b, 32'hc019f060} /* (14, 7, 21) {real, imag} */,
  {32'hbf515479, 32'hbf08962a} /* (14, 7, 20) {real, imag} */,
  {32'hbe8e999b, 32'hbe9f4194} /* (14, 7, 19) {real, imag} */,
  {32'h3d62d9ad, 32'h3f6747a7} /* (14, 7, 18) {real, imag} */,
  {32'h3eab22bd, 32'h3dee0b9f} /* (14, 7, 17) {real, imag} */,
  {32'hbe7bf387, 32'hbfb229b4} /* (14, 7, 16) {real, imag} */,
  {32'h3f1a0a51, 32'hbfb776d4} /* (14, 7, 15) {real, imag} */,
  {32'hc024eb87, 32'hbf22a373} /* (14, 7, 14) {real, imag} */,
  {32'h3ffa456b, 32'h3d129cf4} /* (14, 7, 13) {real, imag} */,
  {32'hc0074f6d, 32'h3fbe5848} /* (14, 7, 12) {real, imag} */,
  {32'hbf31474b, 32'hc05f84d6} /* (14, 7, 11) {real, imag} */,
  {32'h40176105, 32'h400d3c1b} /* (14, 7, 10) {real, imag} */,
  {32'hc0008c1e, 32'hbe9cecaf} /* (14, 7, 9) {real, imag} */,
  {32'hbfa7a6c0, 32'hc06b9686} /* (14, 7, 8) {real, imag} */,
  {32'hbee8ee54, 32'hbf0e54c7} /* (14, 7, 7) {real, imag} */,
  {32'h3fab27c1, 32'h3f7b0c5a} /* (14, 7, 6) {real, imag} */,
  {32'h3fb2297c, 32'h3f8d5201} /* (14, 7, 5) {real, imag} */,
  {32'h3f65f31e, 32'h40795d78} /* (14, 7, 4) {real, imag} */,
  {32'h3fb026f3, 32'h3f398413} /* (14, 7, 3) {real, imag} */,
  {32'h3fe26e94, 32'h3fb1032f} /* (14, 7, 2) {real, imag} */,
  {32'hc02ea316, 32'hbfe3709a} /* (14, 7, 1) {real, imag} */,
  {32'hbfa19a10, 32'hbf1b3ac5} /* (14, 7, 0) {real, imag} */,
  {32'h3f741c49, 32'h3f8706b2} /* (14, 6, 31) {real, imag} */,
  {32'h4009e262, 32'h3fc06662} /* (14, 6, 30) {real, imag} */,
  {32'hc05245d6, 32'hbfbf0023} /* (14, 6, 29) {real, imag} */,
  {32'h3f7b0b17, 32'h3f1c3ac1} /* (14, 6, 28) {real, imag} */,
  {32'h3f1f5ea5, 32'h4014e0fc} /* (14, 6, 27) {real, imag} */,
  {32'h3fc1dd15, 32'hbeacc719} /* (14, 6, 26) {real, imag} */,
  {32'hbf44e543, 32'hc004b01f} /* (14, 6, 25) {real, imag} */,
  {32'hbeaa2a60, 32'hbd599590} /* (14, 6, 24) {real, imag} */,
  {32'h3fcfa3c1, 32'h3fcc4791} /* (14, 6, 23) {real, imag} */,
  {32'hbfa54ed6, 32'hc01cc0f3} /* (14, 6, 22) {real, imag} */,
  {32'h3eaa3b2f, 32'h3f873238} /* (14, 6, 21) {real, imag} */,
  {32'h40027723, 32'hbefa3be7} /* (14, 6, 20) {real, imag} */,
  {32'h3f90d80c, 32'hbec66b6c} /* (14, 6, 19) {real, imag} */,
  {32'hbf84d1b8, 32'h3ee5371a} /* (14, 6, 18) {real, imag} */,
  {32'h3f7d36e8, 32'hbebcc1c1} /* (14, 6, 17) {real, imag} */,
  {32'hbfb3f030, 32'hbf6024b3} /* (14, 6, 16) {real, imag} */,
  {32'h3fad3053, 32'h3fdc3ca6} /* (14, 6, 15) {real, imag} */,
  {32'hbf49ec6f, 32'hbf8c59fe} /* (14, 6, 14) {real, imag} */,
  {32'h3e64f96d, 32'h3fdf8c15} /* (14, 6, 13) {real, imag} */,
  {32'hbf6f3bc7, 32'h3ede3510} /* (14, 6, 12) {real, imag} */,
  {32'hbfedc6d1, 32'h3ee60829} /* (14, 6, 11) {real, imag} */,
  {32'h3e578ace, 32'h3f99fd3b} /* (14, 6, 10) {real, imag} */,
  {32'hc0868857, 32'h3fe9ce4a} /* (14, 6, 9) {real, imag} */,
  {32'hbf895ecd, 32'hbfeabf81} /* (14, 6, 8) {real, imag} */,
  {32'h3f80ba74, 32'hbfa6adb4} /* (14, 6, 7) {real, imag} */,
  {32'h3ef066b2, 32'h4000b35b} /* (14, 6, 6) {real, imag} */,
  {32'hbf335dd3, 32'hbf6281e1} /* (14, 6, 5) {real, imag} */,
  {32'h3f98bb4e, 32'hbfad8d0e} /* (14, 6, 4) {real, imag} */,
  {32'h3fa9ec5d, 32'h3fcacd55} /* (14, 6, 3) {real, imag} */,
  {32'hbe29b2c7, 32'h3f351699} /* (14, 6, 2) {real, imag} */,
  {32'h3e0cbb17, 32'hbfd71e07} /* (14, 6, 1) {real, imag} */,
  {32'h400db0fb, 32'hbf8bc8a4} /* (14, 6, 0) {real, imag} */,
  {32'hbf398a48, 32'hbf5753ff} /* (14, 5, 31) {real, imag} */,
  {32'hbdd576a4, 32'hc01ecd31} /* (14, 5, 30) {real, imag} */,
  {32'hbf3935fb, 32'h3faeccb6} /* (14, 5, 29) {real, imag} */,
  {32'h401053be, 32'hbf0e4005} /* (14, 5, 28) {real, imag} */,
  {32'hc001ee96, 32'h3ed00173} /* (14, 5, 27) {real, imag} */,
  {32'hbdbd1019, 32'h3fb269e7} /* (14, 5, 26) {real, imag} */,
  {32'h3fd04142, 32'hbfa75ba4} /* (14, 5, 25) {real, imag} */,
  {32'hbf9e43ae, 32'h40312f5c} /* (14, 5, 24) {real, imag} */,
  {32'h3faeb454, 32'hbf5fe959} /* (14, 5, 23) {real, imag} */,
  {32'hc01155c8, 32'hbfb06b6e} /* (14, 5, 22) {real, imag} */,
  {32'hbfddb845, 32'h3e127d14} /* (14, 5, 21) {real, imag} */,
  {32'hbfce5561, 32'h3f726062} /* (14, 5, 20) {real, imag} */,
  {32'h3fa8bb77, 32'h3fa066ed} /* (14, 5, 19) {real, imag} */,
  {32'hbffa44be, 32'h3fd5886d} /* (14, 5, 18) {real, imag} */,
  {32'hc02eaa38, 32'hbcc67969} /* (14, 5, 17) {real, imag} */,
  {32'h3ff43fd9, 32'h3fb78c2d} /* (14, 5, 16) {real, imag} */,
  {32'hbfa601ac, 32'h3f7f4e4d} /* (14, 5, 15) {real, imag} */,
  {32'h3ff22bc8, 32'h3f8bdef5} /* (14, 5, 14) {real, imag} */,
  {32'h3f9c7e73, 32'hbf571ad8} /* (14, 5, 13) {real, imag} */,
  {32'h3fcaae01, 32'h3f80fb22} /* (14, 5, 12) {real, imag} */,
  {32'h3fb0c9e9, 32'hbe17d07b} /* (14, 5, 11) {real, imag} */,
  {32'hbf084c5f, 32'h3ee7379b} /* (14, 5, 10) {real, imag} */,
  {32'h3fb55b0e, 32'hc08003bb} /* (14, 5, 9) {real, imag} */,
  {32'hbf3641ff, 32'h3fb899c3} /* (14, 5, 8) {real, imag} */,
  {32'hbe3db293, 32'hbf4d5f0b} /* (14, 5, 7) {real, imag} */,
  {32'hbeb3f132, 32'h3f533212} /* (14, 5, 6) {real, imag} */,
  {32'h400d63f3, 32'h3fae1619} /* (14, 5, 5) {real, imag} */,
  {32'h3ee53edb, 32'h40055348} /* (14, 5, 4) {real, imag} */,
  {32'hbd11998d, 32'hbf88a7f4} /* (14, 5, 3) {real, imag} */,
  {32'hbf002a83, 32'hbefc40b1} /* (14, 5, 2) {real, imag} */,
  {32'hbe246ae2, 32'h405fcd2b} /* (14, 5, 1) {real, imag} */,
  {32'h4066416e, 32'h407a28a6} /* (14, 5, 0) {real, imag} */,
  {32'hbffa3342, 32'hc02216a7} /* (14, 4, 31) {real, imag} */,
  {32'h3f6a416a, 32'hbfceb700} /* (14, 4, 30) {real, imag} */,
  {32'h3f4424d7, 32'hc013f8cc} /* (14, 4, 29) {real, imag} */,
  {32'h3e0c2313, 32'h3ee53753} /* (14, 4, 28) {real, imag} */,
  {32'hbf504d70, 32'hbfd1d7b1} /* (14, 4, 27) {real, imag} */,
  {32'h3f366d2f, 32'hbc0cdf0b} /* (14, 4, 26) {real, imag} */,
  {32'h3f35dd3d, 32'hbf8873f9} /* (14, 4, 25) {real, imag} */,
  {32'h3f9e1247, 32'hbf7a0477} /* (14, 4, 24) {real, imag} */,
  {32'h3f5c7975, 32'hbd178f7d} /* (14, 4, 23) {real, imag} */,
  {32'h3d9c102f, 32'h3fbfeb01} /* (14, 4, 22) {real, imag} */,
  {32'hbeb714f1, 32'hbf43af9e} /* (14, 4, 21) {real, imag} */,
  {32'h4027bdd6, 32'h3fcbe0b8} /* (14, 4, 20) {real, imag} */,
  {32'hbf76d3a9, 32'h402e923a} /* (14, 4, 19) {real, imag} */,
  {32'h3f5d1cbf, 32'h3ffba84e} /* (14, 4, 18) {real, imag} */,
  {32'hbda0b828, 32'h3dc47ec7} /* (14, 4, 17) {real, imag} */,
  {32'hbe825e60, 32'hbe2373c4} /* (14, 4, 16) {real, imag} */,
  {32'h3f8b9b26, 32'hbe234d75} /* (14, 4, 15) {real, imag} */,
  {32'hbef3f528, 32'h3ec246ff} /* (14, 4, 14) {real, imag} */,
  {32'hbf178568, 32'h3fabcc16} /* (14, 4, 13) {real, imag} */,
  {32'hbf17b579, 32'h3fb963fd} /* (14, 4, 12) {real, imag} */,
  {32'hc03ab7d1, 32'hbff1d9da} /* (14, 4, 11) {real, imag} */,
  {32'h40068ba9, 32'h3e3e4860} /* (14, 4, 10) {real, imag} */,
  {32'hbf3f9db2, 32'h3e277c17} /* (14, 4, 9) {real, imag} */,
  {32'h3e607231, 32'h3e227bef} /* (14, 4, 8) {real, imag} */,
  {32'hbf8dd23e, 32'h3fa49d12} /* (14, 4, 7) {real, imag} */,
  {32'hbf06c884, 32'hbdaddf93} /* (14, 4, 6) {real, imag} */,
  {32'h3feea5f8, 32'hbfbd4399} /* (14, 4, 5) {real, imag} */,
  {32'h3e65d8dc, 32'hbead1469} /* (14, 4, 4) {real, imag} */,
  {32'h3f1a080e, 32'h3e7a406c} /* (14, 4, 3) {real, imag} */,
  {32'h3f2c2b49, 32'h3f14edf5} /* (14, 4, 2) {real, imag} */,
  {32'hc08ce35d, 32'h4001837a} /* (14, 4, 1) {real, imag} */,
  {32'h3ef877a9, 32'hbf84a29f} /* (14, 4, 0) {real, imag} */,
  {32'h401532fc, 32'hbfeac4e1} /* (14, 3, 31) {real, imag} */,
  {32'h3f98d785, 32'h3ec769d3} /* (14, 3, 30) {real, imag} */,
  {32'hc04cf2cf, 32'h40008afb} /* (14, 3, 29) {real, imag} */,
  {32'hbf44abaf, 32'hbf04f7ae} /* (14, 3, 28) {real, imag} */,
  {32'hbb24c975, 32'hbfeaa16c} /* (14, 3, 27) {real, imag} */,
  {32'hbdbf0c83, 32'hbf7ea94c} /* (14, 3, 26) {real, imag} */,
  {32'h3ee60668, 32'h4035f507} /* (14, 3, 25) {real, imag} */,
  {32'h3f7c54b0, 32'hbe83044d} /* (14, 3, 24) {real, imag} */,
  {32'h3fec21aa, 32'hbf93fc4c} /* (14, 3, 23) {real, imag} */,
  {32'hbf176d5a, 32'h3f7ab9d0} /* (14, 3, 22) {real, imag} */,
  {32'h3fab6233, 32'hbfb117c8} /* (14, 3, 21) {real, imag} */,
  {32'hbd78826d, 32'hbf82945e} /* (14, 3, 20) {real, imag} */,
  {32'h3f38bb48, 32'hbf231307} /* (14, 3, 19) {real, imag} */,
  {32'hbfc60700, 32'h3fe81581} /* (14, 3, 18) {real, imag} */,
  {32'hbfc94eec, 32'hbf63cb04} /* (14, 3, 17) {real, imag} */,
  {32'h3fdd8320, 32'h3db59e46} /* (14, 3, 16) {real, imag} */,
  {32'h402663e2, 32'h3f7417b7} /* (14, 3, 15) {real, imag} */,
  {32'hbf8e51d1, 32'hbec6b439} /* (14, 3, 14) {real, imag} */,
  {32'hbea44045, 32'h3fdd6bb4} /* (14, 3, 13) {real, imag} */,
  {32'hbfcc8eda, 32'h3fb37c17} /* (14, 3, 12) {real, imag} */,
  {32'hbf8745e1, 32'h3ec5af00} /* (14, 3, 11) {real, imag} */,
  {32'hbb72ea3b, 32'hbff3d36b} /* (14, 3, 10) {real, imag} */,
  {32'hbf9a0cab, 32'h3f0985ef} /* (14, 3, 9) {real, imag} */,
  {32'h3f4134d6, 32'h3cc56c8f} /* (14, 3, 8) {real, imag} */,
  {32'h3f149048, 32'hbf62b416} /* (14, 3, 7) {real, imag} */,
  {32'h3ebcbeb1, 32'h3f2f310a} /* (14, 3, 6) {real, imag} */,
  {32'h3ff46435, 32'hbf30b28d} /* (14, 3, 5) {real, imag} */,
  {32'h4016dfe9, 32'hbf95a515} /* (14, 3, 4) {real, imag} */,
  {32'h3dc99dcc, 32'hbfb6f636} /* (14, 3, 3) {real, imag} */,
  {32'hbe23e316, 32'hbde64992} /* (14, 3, 2) {real, imag} */,
  {32'hbf514f08, 32'hbf8b11f1} /* (14, 3, 1) {real, imag} */,
  {32'h3f5221b7, 32'hbebaa896} /* (14, 3, 0) {real, imag} */,
  {32'h40d75171, 32'h3f4b4f32} /* (14, 2, 31) {real, imag} */,
  {32'hc0ac02d5, 32'h40413826} /* (14, 2, 30) {real, imag} */,
  {32'h3f523d10, 32'hc005b64e} /* (14, 2, 29) {real, imag} */,
  {32'h3f6b989a, 32'hbf80336c} /* (14, 2, 28) {real, imag} */,
  {32'h3f2defeb, 32'h4003f152} /* (14, 2, 27) {real, imag} */,
  {32'h400ed288, 32'hbe8b9a71} /* (14, 2, 26) {real, imag} */,
  {32'hbfbb0830, 32'hbedf0d00} /* (14, 2, 25) {real, imag} */,
  {32'hbfb4f19a, 32'h406831e2} /* (14, 2, 24) {real, imag} */,
  {32'h3d20d476, 32'h3f6593ce} /* (14, 2, 23) {real, imag} */,
  {32'h3fec1a75, 32'h3daf978f} /* (14, 2, 22) {real, imag} */,
  {32'hbfb91d08, 32'h3feb14cc} /* (14, 2, 21) {real, imag} */,
  {32'hbe30ea3c, 32'hbd4f678c} /* (14, 2, 20) {real, imag} */,
  {32'h3eb6ffd0, 32'hbefae771} /* (14, 2, 19) {real, imag} */,
  {32'hbf83f2e8, 32'hc01625e0} /* (14, 2, 18) {real, imag} */,
  {32'h3f4f7f4b, 32'hbeba2678} /* (14, 2, 17) {real, imag} */,
  {32'h3f84611e, 32'hbde2e9c2} /* (14, 2, 16) {real, imag} */,
  {32'h3fc4c13e, 32'h3f77421c} /* (14, 2, 15) {real, imag} */,
  {32'hbfb1ad74, 32'hc0158fe9} /* (14, 2, 14) {real, imag} */,
  {32'h3ead31e1, 32'h40499a82} /* (14, 2, 13) {real, imag} */,
  {32'hc03637b0, 32'hbee5ffbb} /* (14, 2, 12) {real, imag} */,
  {32'h3ffde9a3, 32'hc00f5c5b} /* (14, 2, 11) {real, imag} */,
  {32'hc01460fb, 32'h3f81e13a} /* (14, 2, 10) {real, imag} */,
  {32'h3feb97d6, 32'h3f50e2de} /* (14, 2, 9) {real, imag} */,
  {32'h3f921ff6, 32'hbde96992} /* (14, 2, 8) {real, imag} */,
  {32'h3fa8ab10, 32'h3c7200e1} /* (14, 2, 7) {real, imag} */,
  {32'h3f02d062, 32'hbf5e4585} /* (14, 2, 6) {real, imag} */,
  {32'h4043cc49, 32'hbfeae7d8} /* (14, 2, 5) {real, imag} */,
  {32'h3f3b11cf, 32'h3f4000c8} /* (14, 2, 4) {real, imag} */,
  {32'hb980113f, 32'h3fdca0f8} /* (14, 2, 3) {real, imag} */,
  {32'hbf65ca1c, 32'h400343a3} /* (14, 2, 2) {real, imag} */,
  {32'h3fd90ab7, 32'h3e57653d} /* (14, 2, 1) {real, imag} */,
  {32'h40427640, 32'h3f3cb94c} /* (14, 2, 0) {real, imag} */,
  {32'hc09bfa6e, 32'h404d330b} /* (14, 1, 31) {real, imag} */,
  {32'h40558d32, 32'hbf99ed72} /* (14, 1, 30) {real, imag} */,
  {32'h3efe46a8, 32'hbfa8e31e} /* (14, 1, 29) {real, imag} */,
  {32'hbf958401, 32'hbfe1a489} /* (14, 1, 28) {real, imag} */,
  {32'h400d61fa, 32'hc0511bbc} /* (14, 1, 27) {real, imag} */,
  {32'h3f023574, 32'hbd3b0fce} /* (14, 1, 26) {real, imag} */,
  {32'h3f9ebe9e, 32'h3fb81023} /* (14, 1, 25) {real, imag} */,
  {32'hc052b399, 32'h3ffd2a60} /* (14, 1, 24) {real, imag} */,
  {32'h3f55aff0, 32'hbfdc7844} /* (14, 1, 23) {real, imag} */,
  {32'h3f1c49ff, 32'h3f57e0a7} /* (14, 1, 22) {real, imag} */,
  {32'h3fb93fed, 32'h3f962adb} /* (14, 1, 21) {real, imag} */,
  {32'hbfbfd66d, 32'hbf70eed4} /* (14, 1, 20) {real, imag} */,
  {32'h3f07d063, 32'hbe9e3b29} /* (14, 1, 19) {real, imag} */,
  {32'h3edbc00d, 32'hbd99c303} /* (14, 1, 18) {real, imag} */,
  {32'h3e7c95c3, 32'hc01a0c57} /* (14, 1, 17) {real, imag} */,
  {32'h3d386da8, 32'hbdbf91e9} /* (14, 1, 16) {real, imag} */,
  {32'hbfdc3ef5, 32'hc0004dc3} /* (14, 1, 15) {real, imag} */,
  {32'hbfbeef32, 32'h3fc99d5b} /* (14, 1, 14) {real, imag} */,
  {32'h3fee71a8, 32'hbf610b67} /* (14, 1, 13) {real, imag} */,
  {32'hbd1623d0, 32'hbf2b703f} /* (14, 1, 12) {real, imag} */,
  {32'h3f8f9e27, 32'hbf5348fb} /* (14, 1, 11) {real, imag} */,
  {32'h3f8a64eb, 32'h40272f91} /* (14, 1, 10) {real, imag} */,
  {32'h40361ac9, 32'h3eec06b1} /* (14, 1, 9) {real, imag} */,
  {32'hbf01db57, 32'hbf3b1b7a} /* (14, 1, 8) {real, imag} */,
  {32'h3f80bc36, 32'h3baf7bdd} /* (14, 1, 7) {real, imag} */,
  {32'hbf0e2a67, 32'hbfcb2a48} /* (14, 1, 6) {real, imag} */,
  {32'hbe854b3d, 32'h3e857007} /* (14, 1, 5) {real, imag} */,
  {32'hbfabcfbf, 32'h400f47ad} /* (14, 1, 4) {real, imag} */,
  {32'hbeead71e, 32'h3f0af515} /* (14, 1, 3) {real, imag} */,
  {32'h40898cca, 32'h3e787ee6} /* (14, 1, 2) {real, imag} */,
  {32'hc0d3b970, 32'hc044ea7d} /* (14, 1, 1) {real, imag} */,
  {32'hc08991b1, 32'h3f03be47} /* (14, 1, 0) {real, imag} */,
  {32'hbf7935ec, 32'h3fd9163a} /* (14, 0, 31) {real, imag} */,
  {32'h3f14056c, 32'h3f81543c} /* (14, 0, 30) {real, imag} */,
  {32'h3f52be18, 32'hbfe637ab} /* (14, 0, 29) {real, imag} */,
  {32'h401bf50c, 32'hbec09f4b} /* (14, 0, 28) {real, imag} */,
  {32'h3ff37a52, 32'hbd2e893b} /* (14, 0, 27) {real, imag} */,
  {32'hc0112a53, 32'h403b0452} /* (14, 0, 26) {real, imag} */,
  {32'h3ffe8523, 32'h4047c1f0} /* (14, 0, 25) {real, imag} */,
  {32'hbfed6d0e, 32'hbf784581} /* (14, 0, 24) {real, imag} */,
  {32'h40167802, 32'hbfd38a71} /* (14, 0, 23) {real, imag} */,
  {32'h3e5294f0, 32'h3f3d4601} /* (14, 0, 22) {real, imag} */,
  {32'h3f77379d, 32'hbee38d3e} /* (14, 0, 21) {real, imag} */,
  {32'hbca740b3, 32'h3dfab48c} /* (14, 0, 20) {real, imag} */,
  {32'h3d8271dd, 32'h3fa0f6a5} /* (14, 0, 19) {real, imag} */,
  {32'hbf84f327, 32'hbead51c1} /* (14, 0, 18) {real, imag} */,
  {32'h3ee40a0c, 32'h3dc55b19} /* (14, 0, 17) {real, imag} */,
  {32'hbfa6ba06, 32'hbf8bbece} /* (14, 0, 16) {real, imag} */,
  {32'h3f69a5ca, 32'h402e482e} /* (14, 0, 15) {real, imag} */,
  {32'h3f1982f7, 32'h3f2dbcbf} /* (14, 0, 14) {real, imag} */,
  {32'hbf93ec11, 32'h3f4ed9bb} /* (14, 0, 13) {real, imag} */,
  {32'h3f626239, 32'h3d306639} /* (14, 0, 12) {real, imag} */,
  {32'h3e98ef32, 32'h3fe0571e} /* (14, 0, 11) {real, imag} */,
  {32'hbf7fec6a, 32'h3ff87ce1} /* (14, 0, 10) {real, imag} */,
  {32'h3f9e5b2a, 32'hc0863a11} /* (14, 0, 9) {real, imag} */,
  {32'hbfca1147, 32'h3e7184b8} /* (14, 0, 8) {real, imag} */,
  {32'hbfec47c9, 32'hbdb15c6b} /* (14, 0, 7) {real, imag} */,
  {32'hbf8473bd, 32'hbf3366be} /* (14, 0, 6) {real, imag} */,
  {32'h3d5f5beb, 32'h3e3d9de2} /* (14, 0, 5) {real, imag} */,
  {32'hbf97ba16, 32'h3d3ebf79} /* (14, 0, 4) {real, imag} */,
  {32'hc013d3bb, 32'hbefd7ea7} /* (14, 0, 3) {real, imag} */,
  {32'h403a7e8a, 32'h3f541e48} /* (14, 0, 2) {real, imag} */,
  {32'hbfc2025c, 32'hc05bc53f} /* (14, 0, 1) {real, imag} */,
  {32'hbff4f8bc, 32'h3fd9fdda} /* (14, 0, 0) {real, imag} */,
  {32'hbea0a70e, 32'hbfa972ed} /* (13, 31, 31) {real, imag} */,
  {32'hbf4ad4a2, 32'hbdf1b2d4} /* (13, 31, 30) {real, imag} */,
  {32'hbf0573fd, 32'h3f86df1e} /* (13, 31, 29) {real, imag} */,
  {32'h40148d9e, 32'hbef5a9ba} /* (13, 31, 28) {real, imag} */,
  {32'hc028e4ec, 32'h3f833175} /* (13, 31, 27) {real, imag} */,
  {32'h3cd2a8b6, 32'hbfbdd617} /* (13, 31, 26) {real, imag} */,
  {32'hbfbb2c7a, 32'h3e9f72b6} /* (13, 31, 25) {real, imag} */,
  {32'h3fff4c8f, 32'hbfd48c05} /* (13, 31, 24) {real, imag} */,
  {32'hbfb197d5, 32'hbf8473dc} /* (13, 31, 23) {real, imag} */,
  {32'h3f5b1b7c, 32'hc009d831} /* (13, 31, 22) {real, imag} */,
  {32'h3f1e5676, 32'h4079fe77} /* (13, 31, 21) {real, imag} */,
  {32'hbf2ec150, 32'h3fc13e4b} /* (13, 31, 20) {real, imag} */,
  {32'hc012248d, 32'h3f828752} /* (13, 31, 19) {real, imag} */,
  {32'hbd839fd4, 32'hbfbc7c48} /* (13, 31, 18) {real, imag} */,
  {32'h3f6e564c, 32'h3e539b0b} /* (13, 31, 17) {real, imag} */,
  {32'hbe6262a8, 32'hbf2f44b7} /* (13, 31, 16) {real, imag} */,
  {32'h3fa4da85, 32'hbf11d487} /* (13, 31, 15) {real, imag} */,
  {32'h3e2fb7e5, 32'h3f4cd226} /* (13, 31, 14) {real, imag} */,
  {32'hbd169314, 32'hbe8fdd21} /* (13, 31, 13) {real, imag} */,
  {32'h3ff1c961, 32'hbff1d33a} /* (13, 31, 12) {real, imag} */,
  {32'hbfb5ecaf, 32'hbfcde70d} /* (13, 31, 11) {real, imag} */,
  {32'h3d967cb9, 32'h401ed1ce} /* (13, 31, 10) {real, imag} */,
  {32'hbef8bb2f, 32'h4064a2e2} /* (13, 31, 9) {real, imag} */,
  {32'hbdb9545b, 32'h3ed0e0b9} /* (13, 31, 8) {real, imag} */,
  {32'hbfa0271c, 32'h3e642e89} /* (13, 31, 7) {real, imag} */,
  {32'h3f444f7d, 32'hc05a95d1} /* (13, 31, 6) {real, imag} */,
  {32'h3f9d75a7, 32'hc0487447} /* (13, 31, 5) {real, imag} */,
  {32'h3e35aae4, 32'hbf401dbd} /* (13, 31, 4) {real, imag} */,
  {32'hc01ed3c0, 32'h3faa5300} /* (13, 31, 3) {real, imag} */,
  {32'h3ff71f03, 32'hbe8d60e0} /* (13, 31, 2) {real, imag} */,
  {32'h3f2ef35a, 32'hbee2f513} /* (13, 31, 1) {real, imag} */,
  {32'h3f41c080, 32'h3f286788} /* (13, 31, 0) {real, imag} */,
  {32'hbf8f1f45, 32'hc0056b4b} /* (13, 30, 31) {real, imag} */,
  {32'h3f81e39c, 32'h3fb4e074} /* (13, 30, 30) {real, imag} */,
  {32'hbf909032, 32'hbd099eba} /* (13, 30, 29) {real, imag} */,
  {32'h3ed1fe4e, 32'hbf5f6810} /* (13, 30, 28) {real, imag} */,
  {32'h3f3e3fac, 32'h3dd35f49} /* (13, 30, 27) {real, imag} */,
  {32'hbeca0764, 32'h4000fbff} /* (13, 30, 26) {real, imag} */,
  {32'h3e2714a9, 32'hc0089e36} /* (13, 30, 25) {real, imag} */,
  {32'hbe67bafb, 32'h3dbb9ccc} /* (13, 30, 24) {real, imag} */,
  {32'h3f5f9e4f, 32'hbf84548b} /* (13, 30, 23) {real, imag} */,
  {32'h400bd7db, 32'h3fb60958} /* (13, 30, 22) {real, imag} */,
  {32'hbeff58d7, 32'h3ea01119} /* (13, 30, 21) {real, imag} */,
  {32'h4019f84e, 32'h3f53bb8f} /* (13, 30, 20) {real, imag} */,
  {32'h3d353410, 32'h3fc6aec9} /* (13, 30, 19) {real, imag} */,
  {32'hbf782684, 32'h3fa983b4} /* (13, 30, 18) {real, imag} */,
  {32'h3f118474, 32'hbef1a3c3} /* (13, 30, 17) {real, imag} */,
  {32'hbfa35fda, 32'h3ffefc0a} /* (13, 30, 16) {real, imag} */,
  {32'h3f07d194, 32'h3e7ea1dc} /* (13, 30, 15) {real, imag} */,
  {32'h3e5facd3, 32'h3ebc6d4a} /* (13, 30, 14) {real, imag} */,
  {32'hbfc68e8e, 32'hbf648dd5} /* (13, 30, 13) {real, imag} */,
  {32'hbf027857, 32'hbf914281} /* (13, 30, 12) {real, imag} */,
  {32'h4039c234, 32'h3fcf5390} /* (13, 30, 11) {real, imag} */,
  {32'h401cbddf, 32'h3e502065} /* (13, 30, 10) {real, imag} */,
  {32'hbf86fa20, 32'h4013f16c} /* (13, 30, 9) {real, imag} */,
  {32'h40068fc2, 32'h3ff514ce} /* (13, 30, 8) {real, imag} */,
  {32'hbfa05bbc, 32'hc05b2b21} /* (13, 30, 7) {real, imag} */,
  {32'hc05f7d8a, 32'hbe7e3163} /* (13, 30, 6) {real, imag} */,
  {32'hbfe7c642, 32'h3fd80312} /* (13, 30, 5) {real, imag} */,
  {32'hbf6b0955, 32'h3fd613d4} /* (13, 30, 4) {real, imag} */,
  {32'h3f43bfc4, 32'h3fefc689} /* (13, 30, 3) {real, imag} */,
  {32'h3f3315c4, 32'hc053ea2b} /* (13, 30, 2) {real, imag} */,
  {32'h3effd838, 32'hbf722086} /* (13, 30, 1) {real, imag} */,
  {32'hbfc4e39d, 32'hbf34589e} /* (13, 30, 0) {real, imag} */,
  {32'h3fdd4bdd, 32'h3f96ae68} /* (13, 29, 31) {real, imag} */,
  {32'hbff0673c, 32'hbf38f065} /* (13, 29, 30) {real, imag} */,
  {32'hbfa5244d, 32'hbd204964} /* (13, 29, 29) {real, imag} */,
  {32'hbffe29a0, 32'hbfe6db48} /* (13, 29, 28) {real, imag} */,
  {32'h3dad3d8d, 32'hbeacd4e5} /* (13, 29, 27) {real, imag} */,
  {32'h40896e94, 32'h3f6ba95c} /* (13, 29, 26) {real, imag} */,
  {32'hbf4fc6a7, 32'h3f4cf577} /* (13, 29, 25) {real, imag} */,
  {32'h400e1d7c, 32'hc00dabf9} /* (13, 29, 24) {real, imag} */,
  {32'h3ea9e1b3, 32'h3ec27f2b} /* (13, 29, 23) {real, imag} */,
  {32'h3fec9a34, 32'h3ed9f288} /* (13, 29, 22) {real, imag} */,
  {32'hc011b8f8, 32'hbf025f71} /* (13, 29, 21) {real, imag} */,
  {32'h4022aba4, 32'h40288f1f} /* (13, 29, 20) {real, imag} */,
  {32'h3f964bb4, 32'hc0362592} /* (13, 29, 19) {real, imag} */,
  {32'hbe46fcfe, 32'h4044965f} /* (13, 29, 18) {real, imag} */,
  {32'h3d885361, 32'h3fd6fbcd} /* (13, 29, 17) {real, imag} */,
  {32'hbfb99bf3, 32'h3fdcad23} /* (13, 29, 16) {real, imag} */,
  {32'hbf655a0f, 32'h3fcbdd9d} /* (13, 29, 15) {real, imag} */,
  {32'hbf556262, 32'hbfaa388c} /* (13, 29, 14) {real, imag} */,
  {32'hbf159321, 32'hbffe0073} /* (13, 29, 13) {real, imag} */,
  {32'h3e015286, 32'h3f95955c} /* (13, 29, 12) {real, imag} */,
  {32'hc02b195f, 32'hbff37214} /* (13, 29, 11) {real, imag} */,
  {32'hc002fe60, 32'hc006de93} /* (13, 29, 10) {real, imag} */,
  {32'h3f1a1a52, 32'hbf807460} /* (13, 29, 9) {real, imag} */,
  {32'hbfb5a16e, 32'hbf1d85a9} /* (13, 29, 8) {real, imag} */,
  {32'h3f924d37, 32'hbfa337b1} /* (13, 29, 7) {real, imag} */,
  {32'h3f23adfe, 32'hbf813d8b} /* (13, 29, 6) {real, imag} */,
  {32'hbfcf71f7, 32'hbf6981eb} /* (13, 29, 5) {real, imag} */,
  {32'h3e9a6d24, 32'h4004c063} /* (13, 29, 4) {real, imag} */,
  {32'hbdda91ce, 32'h4020b40d} /* (13, 29, 3) {real, imag} */,
  {32'h3f2c8bc4, 32'hc01bbeb5} /* (13, 29, 2) {real, imag} */,
  {32'hbd872f9c, 32'h3fffecc2} /* (13, 29, 1) {real, imag} */,
  {32'h3ebf3eb5, 32'h3f88494d} /* (13, 29, 0) {real, imag} */,
  {32'hbd099138, 32'hc0667871} /* (13, 28, 31) {real, imag} */,
  {32'h3fca7b9d, 32'h4069ce15} /* (13, 28, 30) {real, imag} */,
  {32'hbfb8d0a2, 32'hbfbbb737} /* (13, 28, 29) {real, imag} */,
  {32'h3f2ea902, 32'h3fc69aea} /* (13, 28, 28) {real, imag} */,
  {32'hbf5154d4, 32'hbf67840a} /* (13, 28, 27) {real, imag} */,
  {32'hbfb6cd7a, 32'h3f449f0a} /* (13, 28, 26) {real, imag} */,
  {32'h3e64e239, 32'hbf47f661} /* (13, 28, 25) {real, imag} */,
  {32'h3f104bf6, 32'hbf2649ec} /* (13, 28, 24) {real, imag} */,
  {32'hbd8fe2cc, 32'h400a7694} /* (13, 28, 23) {real, imag} */,
  {32'h3fa52772, 32'h3e8e6396} /* (13, 28, 22) {real, imag} */,
  {32'hc01c0ebb, 32'hc0155bd6} /* (13, 28, 21) {real, imag} */,
  {32'hbf9b5818, 32'hc0192717} /* (13, 28, 20) {real, imag} */,
  {32'hbe07d7d4, 32'hbfa6a208} /* (13, 28, 19) {real, imag} */,
  {32'h3facf103, 32'hbf7c5f50} /* (13, 28, 18) {real, imag} */,
  {32'hbfd08462, 32'hbffccd6f} /* (13, 28, 17) {real, imag} */,
  {32'h3f42487b, 32'hbf5c9da4} /* (13, 28, 16) {real, imag} */,
  {32'h3f5c8079, 32'h3f7098ed} /* (13, 28, 15) {real, imag} */,
  {32'hbf91c6db, 32'hc02a2d8f} /* (13, 28, 14) {real, imag} */,
  {32'hc043e36e, 32'hc014e6ae} /* (13, 28, 13) {real, imag} */,
  {32'hc067cf31, 32'hbe06a32d} /* (13, 28, 12) {real, imag} */,
  {32'h3fc06290, 32'h3fd8dabb} /* (13, 28, 11) {real, imag} */,
  {32'h402a6c2f, 32'h40145b6b} /* (13, 28, 10) {real, imag} */,
  {32'hc009defe, 32'h3f0cd779} /* (13, 28, 9) {real, imag} */,
  {32'h3fcbc0c5, 32'h40199400} /* (13, 28, 8) {real, imag} */,
  {32'h404ab81f, 32'h3fb115c8} /* (13, 28, 7) {real, imag} */,
  {32'hbf860d01, 32'hc00d7c88} /* (13, 28, 6) {real, imag} */,
  {32'h3e0fefe6, 32'hbdca351d} /* (13, 28, 5) {real, imag} */,
  {32'h3f853523, 32'hbe1b1393} /* (13, 28, 4) {real, imag} */,
  {32'h3d855dac, 32'hbf87f1a6} /* (13, 28, 3) {real, imag} */,
  {32'hc05e57e2, 32'hc000dff6} /* (13, 28, 2) {real, imag} */,
  {32'h3f318107, 32'h3f95acbe} /* (13, 28, 1) {real, imag} */,
  {32'hc00d0987, 32'h3dfa706b} /* (13, 28, 0) {real, imag} */,
  {32'h3f1b382c, 32'hc0261133} /* (13, 27, 31) {real, imag} */,
  {32'h3e932ddc, 32'h3d8f60d4} /* (13, 27, 30) {real, imag} */,
  {32'h4023c5c4, 32'h3f76e7a8} /* (13, 27, 29) {real, imag} */,
  {32'hbff9c7a0, 32'hbf675c9c} /* (13, 27, 28) {real, imag} */,
  {32'h40285685, 32'hbffbe71c} /* (13, 27, 27) {real, imag} */,
  {32'h3ea68e7a, 32'h4015b32a} /* (13, 27, 26) {real, imag} */,
  {32'hc043d8d1, 32'hbe293f47} /* (13, 27, 25) {real, imag} */,
  {32'hc07d655a, 32'hbf651364} /* (13, 27, 24) {real, imag} */,
  {32'h402825c3, 32'hbd9c62f7} /* (13, 27, 23) {real, imag} */,
  {32'h4042520b, 32'h3f9a84ec} /* (13, 27, 22) {real, imag} */,
  {32'h3f02861d, 32'h3f99397f} /* (13, 27, 21) {real, imag} */,
  {32'h3ed2e465, 32'h3f753ccd} /* (13, 27, 20) {real, imag} */,
  {32'h3eb96862, 32'hbfb164b1} /* (13, 27, 19) {real, imag} */,
  {32'hc00a1b70, 32'hbf2310a5} /* (13, 27, 18) {real, imag} */,
  {32'hbf1c64e0, 32'hbee30bfb} /* (13, 27, 17) {real, imag} */,
  {32'h3ee9bb01, 32'h3fad1683} /* (13, 27, 16) {real, imag} */,
  {32'h3f3c61a8, 32'h402c0fc2} /* (13, 27, 15) {real, imag} */,
  {32'hc01721c4, 32'h404bd86b} /* (13, 27, 14) {real, imag} */,
  {32'hbf178001, 32'h3ef75b5b} /* (13, 27, 13) {real, imag} */,
  {32'hbeccf355, 32'h3fbbc49b} /* (13, 27, 12) {real, imag} */,
  {32'h4047f8fa, 32'h3c9d0982} /* (13, 27, 11) {real, imag} */,
  {32'h3e037307, 32'h402c6d53} /* (13, 27, 10) {real, imag} */,
  {32'hc0330aec, 32'hbf20edec} /* (13, 27, 9) {real, imag} */,
  {32'hc0066bd6, 32'hbfd1692a} /* (13, 27, 8) {real, imag} */,
  {32'hbfd81ef2, 32'hbecc1bfe} /* (13, 27, 7) {real, imag} */,
  {32'h4003822a, 32'h3f3c5e2a} /* (13, 27, 6) {real, imag} */,
  {32'hc013d293, 32'hbfa1503a} /* (13, 27, 5) {real, imag} */,
  {32'hbd27e359, 32'hc068b32c} /* (13, 27, 4) {real, imag} */,
  {32'hbe9cc80f, 32'h3f4ff48a} /* (13, 27, 3) {real, imag} */,
  {32'hbfc4fdb8, 32'h3f4eaf14} /* (13, 27, 2) {real, imag} */,
  {32'h3f237f33, 32'h3fdda81e} /* (13, 27, 1) {real, imag} */,
  {32'hbfeb117c, 32'hbf9dc393} /* (13, 27, 0) {real, imag} */,
  {32'h400ca8ea, 32'h4044238f} /* (13, 26, 31) {real, imag} */,
  {32'hbfd33b26, 32'h3f95cfb5} /* (13, 26, 30) {real, imag} */,
  {32'hbfadf627, 32'h3fbb1a00} /* (13, 26, 29) {real, imag} */,
  {32'h3f986231, 32'h3ee17696} /* (13, 26, 28) {real, imag} */,
  {32'h3f85bd92, 32'h3fe73392} /* (13, 26, 27) {real, imag} */,
  {32'hc0191ea7, 32'hbe2a0e17} /* (13, 26, 26) {real, imag} */,
  {32'hc0383d42, 32'h3f2b3fce} /* (13, 26, 25) {real, imag} */,
  {32'hbe9c5a90, 32'hbf82febe} /* (13, 26, 24) {real, imag} */,
  {32'hc060d929, 32'h3fe27258} /* (13, 26, 23) {real, imag} */,
  {32'hbf14c43a, 32'h3f183dc8} /* (13, 26, 22) {real, imag} */,
  {32'h3fcb16e6, 32'hc0090d79} /* (13, 26, 21) {real, imag} */,
  {32'h3fd8fd13, 32'hbf832d61} /* (13, 26, 20) {real, imag} */,
  {32'h3f06c96f, 32'hbf823e39} /* (13, 26, 19) {real, imag} */,
  {32'hc0857c87, 32'hc01ccdcb} /* (13, 26, 18) {real, imag} */,
  {32'hbf8d5abf, 32'h3fd6e089} /* (13, 26, 17) {real, imag} */,
  {32'h3f06ff5b, 32'hc0050ebe} /* (13, 26, 16) {real, imag} */,
  {32'h3f29d381, 32'hc0030d48} /* (13, 26, 15) {real, imag} */,
  {32'h3f6cf7d0, 32'hbfce541a} /* (13, 26, 14) {real, imag} */,
  {32'hbf6d6404, 32'h3f43d20c} /* (13, 26, 13) {real, imag} */,
  {32'h3f43f133, 32'h3d9b5cf1} /* (13, 26, 12) {real, imag} */,
  {32'h3fbc9430, 32'hbf411cd4} /* (13, 26, 11) {real, imag} */,
  {32'hc02c05b5, 32'hbeb293af} /* (13, 26, 10) {real, imag} */,
  {32'h3fc3d318, 32'hbfd502c8} /* (13, 26, 9) {real, imag} */,
  {32'h3d883b3c, 32'h402038fb} /* (13, 26, 8) {real, imag} */,
  {32'h3f652444, 32'hc0210e59} /* (13, 26, 7) {real, imag} */,
  {32'hbfb8c8b7, 32'h3f8ec327} /* (13, 26, 6) {real, imag} */,
  {32'h3ebc335f, 32'hbf0a3dd8} /* (13, 26, 5) {real, imag} */,
  {32'hbf304605, 32'hbf916529} /* (13, 26, 4) {real, imag} */,
  {32'h40036281, 32'h3faafc99} /* (13, 26, 3) {real, imag} */,
  {32'h3f2cbe54, 32'h3f38c539} /* (13, 26, 2) {real, imag} */,
  {32'h403217d7, 32'h40336ce9} /* (13, 26, 1) {real, imag} */,
  {32'h3d53f41a, 32'hc003807d} /* (13, 26, 0) {real, imag} */,
  {32'hbf881d0d, 32'h3f1203ba} /* (13, 25, 31) {real, imag} */,
  {32'hc0926d36, 32'hbf8da410} /* (13, 25, 30) {real, imag} */,
  {32'hbfa2c4f9, 32'h3ee35204} /* (13, 25, 29) {real, imag} */,
  {32'h3f37e1a9, 32'hbfbf5c5e} /* (13, 25, 28) {real, imag} */,
  {32'hc020f95d, 32'h3e4b289e} /* (13, 25, 27) {real, imag} */,
  {32'hbf6d6bbe, 32'h4046944d} /* (13, 25, 26) {real, imag} */,
  {32'hc0085214, 32'hbf092a69} /* (13, 25, 25) {real, imag} */,
  {32'h3e864f1a, 32'h3ed9412e} /* (13, 25, 24) {real, imag} */,
  {32'h3fa8c0b6, 32'h3f8ecb1a} /* (13, 25, 23) {real, imag} */,
  {32'h3ffcb52e, 32'h3f2b87ee} /* (13, 25, 22) {real, imag} */,
  {32'h3f039d20, 32'hbf90e26a} /* (13, 25, 21) {real, imag} */,
  {32'h40108c00, 32'hc01db4a6} /* (13, 25, 20) {real, imag} */,
  {32'h3f85fa31, 32'h3ea8f0f6} /* (13, 25, 19) {real, imag} */,
  {32'hbf2d21bf, 32'hbfb2ae55} /* (13, 25, 18) {real, imag} */,
  {32'h3f318348, 32'h3dd1115b} /* (13, 25, 17) {real, imag} */,
  {32'h3f241a50, 32'hbf225f1f} /* (13, 25, 16) {real, imag} */,
  {32'hbf855535, 32'h3e93177b} /* (13, 25, 15) {real, imag} */,
  {32'h3f3a0807, 32'hbee11498} /* (13, 25, 14) {real, imag} */,
  {32'h3fa8d75e, 32'h40383439} /* (13, 25, 13) {real, imag} */,
  {32'h3ef6a463, 32'h400a68ba} /* (13, 25, 12) {real, imag} */,
  {32'h3fe48ff9, 32'h3fda3c1c} /* (13, 25, 11) {real, imag} */,
  {32'h406b60bc, 32'h3f3059ce} /* (13, 25, 10) {real, imag} */,
  {32'h3d3cf253, 32'hbeb8ee35} /* (13, 25, 9) {real, imag} */,
  {32'hbff4463c, 32'hbfd276fd} /* (13, 25, 8) {real, imag} */,
  {32'h4042ea35, 32'hc00601f6} /* (13, 25, 7) {real, imag} */,
  {32'hbebb8dd3, 32'hbfb921b2} /* (13, 25, 6) {real, imag} */,
  {32'hbfc9c89f, 32'h4065e5bc} /* (13, 25, 5) {real, imag} */,
  {32'hbdcbc391, 32'hbe874311} /* (13, 25, 4) {real, imag} */,
  {32'hbe9b615e, 32'hc04e9027} /* (13, 25, 3) {real, imag} */,
  {32'h3deb1db7, 32'h4047a9b4} /* (13, 25, 2) {real, imag} */,
  {32'hbf9debd9, 32'h3f134d54} /* (13, 25, 1) {real, imag} */,
  {32'h3f5bccdf, 32'hbf1bec7e} /* (13, 25, 0) {real, imag} */,
  {32'hbf2657a0, 32'h3d52db8b} /* (13, 24, 31) {real, imag} */,
  {32'hc0014a6f, 32'hbfd347b6} /* (13, 24, 30) {real, imag} */,
  {32'hbfa9e043, 32'h3ec79c04} /* (13, 24, 29) {real, imag} */,
  {32'hbe910c86, 32'h3f79ab2a} /* (13, 24, 28) {real, imag} */,
  {32'hbd997626, 32'hbffac31f} /* (13, 24, 27) {real, imag} */,
  {32'hbfbd4312, 32'h3ffe50aa} /* (13, 24, 26) {real, imag} */,
  {32'h3e70104b, 32'hbec3b6bc} /* (13, 24, 25) {real, imag} */,
  {32'h40939bbc, 32'hbee6e0e1} /* (13, 24, 24) {real, imag} */,
  {32'hbf563b5d, 32'hbf29db63} /* (13, 24, 23) {real, imag} */,
  {32'h3ee00def, 32'hbfa3a700} /* (13, 24, 22) {real, imag} */,
  {32'h403a1f72, 32'hc00f910b} /* (13, 24, 21) {real, imag} */,
  {32'hbfccb8d9, 32'hbdf5e3ee} /* (13, 24, 20) {real, imag} */,
  {32'hbfa37834, 32'hbfb93a0e} /* (13, 24, 19) {real, imag} */,
  {32'h3ec5ae7e, 32'h4038d761} /* (13, 24, 18) {real, imag} */,
  {32'hc010b464, 32'h3e2c432e} /* (13, 24, 17) {real, imag} */,
  {32'hbdeb2d30, 32'h3f4d63b2} /* (13, 24, 16) {real, imag} */,
  {32'h3f38eb89, 32'h3f58a271} /* (13, 24, 15) {real, imag} */,
  {32'h3e98394b, 32'h3fad6dea} /* (13, 24, 14) {real, imag} */,
  {32'h3ffb3670, 32'hc08e5b74} /* (13, 24, 13) {real, imag} */,
  {32'hbf4c54c0, 32'h3fab6e09} /* (13, 24, 12) {real, imag} */,
  {32'h3ed56f74, 32'h3f173496} /* (13, 24, 11) {real, imag} */,
  {32'hbf8fd421, 32'h3f12fe5c} /* (13, 24, 10) {real, imag} */,
  {32'h3f76234b, 32'h3f0b3a56} /* (13, 24, 9) {real, imag} */,
  {32'h3f66824c, 32'hbff82c36} /* (13, 24, 8) {real, imag} */,
  {32'hbf772111, 32'hc00c2330} /* (13, 24, 7) {real, imag} */,
  {32'h3f090b7b, 32'h3f8725da} /* (13, 24, 6) {real, imag} */,
  {32'hbf7a2724, 32'h3f5b6795} /* (13, 24, 5) {real, imag} */,
  {32'h4005a25b, 32'h4008bb97} /* (13, 24, 4) {real, imag} */,
  {32'hbe84368d, 32'hbe930abd} /* (13, 24, 3) {real, imag} */,
  {32'h3f85b4db, 32'hbfb0119f} /* (13, 24, 2) {real, imag} */,
  {32'hbede5528, 32'hc003af7d} /* (13, 24, 1) {real, imag} */,
  {32'h3f0293ba, 32'hbf2a190b} /* (13, 24, 0) {real, imag} */,
  {32'hc001e325, 32'h40381a1a} /* (13, 23, 31) {real, imag} */,
  {32'h3ed2a0c2, 32'h400803b9} /* (13, 23, 30) {real, imag} */,
  {32'h3f9d368a, 32'h3e38b741} /* (13, 23, 29) {real, imag} */,
  {32'h3f046593, 32'hbf5cd0f7} /* (13, 23, 28) {real, imag} */,
  {32'hbfeb414e, 32'h3da934ca} /* (13, 23, 27) {real, imag} */,
  {32'h3f109a31, 32'hc070cbe1} /* (13, 23, 26) {real, imag} */,
  {32'hbf3c60e7, 32'hbf5555ec} /* (13, 23, 25) {real, imag} */,
  {32'h3f94855e, 32'hc08d5266} /* (13, 23, 24) {real, imag} */,
  {32'hbf1da512, 32'h402c41df} /* (13, 23, 23) {real, imag} */,
  {32'h3d7f093e, 32'h3e0c4140} /* (13, 23, 22) {real, imag} */,
  {32'h3f7d83f7, 32'h3f0f2889} /* (13, 23, 21) {real, imag} */,
  {32'h3ccb8c60, 32'hc03502ad} /* (13, 23, 20) {real, imag} */,
  {32'h3f126178, 32'h3bbb8de3} /* (13, 23, 19) {real, imag} */,
  {32'h3f98aabf, 32'h3f0890ea} /* (13, 23, 18) {real, imag} */,
  {32'hbfc85edf, 32'hbec91a28} /* (13, 23, 17) {real, imag} */,
  {32'hbfa5a0a6, 32'hbfb2159f} /* (13, 23, 16) {real, imag} */,
  {32'hc0190014, 32'hbeaa8ee8} /* (13, 23, 15) {real, imag} */,
  {32'hc0208e79, 32'h4083fc26} /* (13, 23, 14) {real, imag} */,
  {32'h408cb313, 32'h3fbecbfb} /* (13, 23, 13) {real, imag} */,
  {32'h3e407775, 32'hbf2655b5} /* (13, 23, 12) {real, imag} */,
  {32'h400aadde, 32'hc07f6599} /* (13, 23, 11) {real, imag} */,
  {32'hbf11fd85, 32'hc010011a} /* (13, 23, 10) {real, imag} */,
  {32'hc0040494, 32'hbffd8222} /* (13, 23, 9) {real, imag} */,
  {32'hbe86cbb3, 32'h401429cc} /* (13, 23, 8) {real, imag} */,
  {32'h3f4de0ca, 32'h3fc8b86c} /* (13, 23, 7) {real, imag} */,
  {32'hbf5badd3, 32'hc0734be4} /* (13, 23, 6) {real, imag} */,
  {32'h400abcee, 32'h3f997643} /* (13, 23, 5) {real, imag} */,
  {32'h3e27a190, 32'h3d09ee74} /* (13, 23, 4) {real, imag} */,
  {32'hbe5a34fb, 32'hbf4aabec} /* (13, 23, 3) {real, imag} */,
  {32'h4031b6a8, 32'hbfcef66e} /* (13, 23, 2) {real, imag} */,
  {32'h3f835112, 32'h402e41ff} /* (13, 23, 1) {real, imag} */,
  {32'hbefef943, 32'h3fad98f3} /* (13, 23, 0) {real, imag} */,
  {32'hbf1d459e, 32'h400abd72} /* (13, 22, 31) {real, imag} */,
  {32'hbf7054c5, 32'hbf0553fe} /* (13, 22, 30) {real, imag} */,
  {32'h3ff9f9c6, 32'hbfcf8540} /* (13, 22, 29) {real, imag} */,
  {32'h3e914bd5, 32'hbfbda0d5} /* (13, 22, 28) {real, imag} */,
  {32'hbf548591, 32'h3f6d566b} /* (13, 22, 27) {real, imag} */,
  {32'hbf028ee2, 32'h3f5cd0f4} /* (13, 22, 26) {real, imag} */,
  {32'hbfcd0069, 32'hbf24714c} /* (13, 22, 25) {real, imag} */,
  {32'h401c4b6d, 32'hbf022060} /* (13, 22, 24) {real, imag} */,
  {32'h3f138e67, 32'hc051795f} /* (13, 22, 23) {real, imag} */,
  {32'hc051a0cf, 32'hbfe78265} /* (13, 22, 22) {real, imag} */,
  {32'hc0a0d07c, 32'h3ef33680} /* (13, 22, 21) {real, imag} */,
  {32'h3f055f30, 32'h404b430a} /* (13, 22, 20) {real, imag} */,
  {32'h3fe57acc, 32'h3f0f9460} /* (13, 22, 19) {real, imag} */,
  {32'h3e987bed, 32'h408cc98a} /* (13, 22, 18) {real, imag} */,
  {32'hbf1fd9f1, 32'h3d8d74ec} /* (13, 22, 17) {real, imag} */,
  {32'hbf19dfc3, 32'h3c14cedd} /* (13, 22, 16) {real, imag} */,
  {32'hc013758b, 32'hbf66260d} /* (13, 22, 15) {real, imag} */,
  {32'h3f8b574d, 32'hc02a823e} /* (13, 22, 14) {real, imag} */,
  {32'hbff96347, 32'hbec92b28} /* (13, 22, 13) {real, imag} */,
  {32'h3f2abf6c, 32'h3f637970} /* (13, 22, 12) {real, imag} */,
  {32'hc00e9055, 32'h400542fe} /* (13, 22, 11) {real, imag} */,
  {32'h3fc90a29, 32'h3e5ec26c} /* (13, 22, 10) {real, imag} */,
  {32'h3fae7ec8, 32'h3e10b62f} /* (13, 22, 9) {real, imag} */,
  {32'h3f12f01b, 32'h3ed22d13} /* (13, 22, 8) {real, imag} */,
  {32'h3f54260a, 32'h3ff48446} /* (13, 22, 7) {real, imag} */,
  {32'hc049f214, 32'h40153c08} /* (13, 22, 6) {real, imag} */,
  {32'h3ffece93, 32'h400419e8} /* (13, 22, 5) {real, imag} */,
  {32'h3fa25a21, 32'hbfcb312f} /* (13, 22, 4) {real, imag} */,
  {32'h3fc4ac77, 32'hbd899b15} /* (13, 22, 3) {real, imag} */,
  {32'hbfb65988, 32'hbd563b9e} /* (13, 22, 2) {real, imag} */,
  {32'hc000eb2c, 32'hbf81c1c7} /* (13, 22, 1) {real, imag} */,
  {32'h3feada62, 32'hbffabfb5} /* (13, 22, 0) {real, imag} */,
  {32'hbdebf633, 32'h3f58659c} /* (13, 21, 31) {real, imag} */,
  {32'hbf69f417, 32'h4068d311} /* (13, 21, 30) {real, imag} */,
  {32'h40758a6b, 32'h407559be} /* (13, 21, 29) {real, imag} */,
  {32'h3ed98103, 32'hbccde61f} /* (13, 21, 28) {real, imag} */,
  {32'hbef2aab1, 32'hc02e53fe} /* (13, 21, 27) {real, imag} */,
  {32'hc00bacc7, 32'h3f3bb078} /* (13, 21, 26) {real, imag} */,
  {32'h4055da5c, 32'h3dceffa3} /* (13, 21, 25) {real, imag} */,
  {32'hbf80530a, 32'h40022742} /* (13, 21, 24) {real, imag} */,
  {32'hbdfc744a, 32'hbdddf18c} /* (13, 21, 23) {real, imag} */,
  {32'hbeee8998, 32'hbec57de0} /* (13, 21, 22) {real, imag} */,
  {32'h4053cdca, 32'hbfacda74} /* (13, 21, 21) {real, imag} */,
  {32'h3e8223c6, 32'hc007a0a8} /* (13, 21, 20) {real, imag} */,
  {32'hc01c3ed8, 32'h3f1c3af7} /* (13, 21, 19) {real, imag} */,
  {32'h3f09b1d8, 32'h3f984ce3} /* (13, 21, 18) {real, imag} */,
  {32'h3da40425, 32'hbed55bb5} /* (13, 21, 17) {real, imag} */,
  {32'hbeb1b03a, 32'h3f84b4f9} /* (13, 21, 16) {real, imag} */,
  {32'hbfe0ce3e, 32'hc0013f04} /* (13, 21, 15) {real, imag} */,
  {32'hbe8f7c1f, 32'hbf952d6c} /* (13, 21, 14) {real, imag} */,
  {32'h406ac0f3, 32'h3efecb1a} /* (13, 21, 13) {real, imag} */,
  {32'h3ff4ce83, 32'h3f262235} /* (13, 21, 12) {real, imag} */,
  {32'h3f1c8841, 32'h406bca9d} /* (13, 21, 11) {real, imag} */,
  {32'hbf2f59f9, 32'h3f81a9e0} /* (13, 21, 10) {real, imag} */,
  {32'h3fba2f74, 32'hc00ab74c} /* (13, 21, 9) {real, imag} */,
  {32'h400ed26e, 32'hbfcd03d9} /* (13, 21, 8) {real, imag} */,
  {32'hc0350b4f, 32'h3ddc3fed} /* (13, 21, 7) {real, imag} */,
  {32'h3f882ee1, 32'hc0abe9ec} /* (13, 21, 6) {real, imag} */,
  {32'hbf2f0dfa, 32'h3f8350bc} /* (13, 21, 5) {real, imag} */,
  {32'h3d1b1c2c, 32'h3fa765fe} /* (13, 21, 4) {real, imag} */,
  {32'h3f81bcbe, 32'h3d955671} /* (13, 21, 3) {real, imag} */,
  {32'h3fe52ec4, 32'hbe675589} /* (13, 21, 2) {real, imag} */,
  {32'h3d75cc5b, 32'hbef4c4d9} /* (13, 21, 1) {real, imag} */,
  {32'hbe90bead, 32'hbe0ba29d} /* (13, 21, 0) {real, imag} */,
  {32'hbf88a583, 32'hbea655b4} /* (13, 20, 31) {real, imag} */,
  {32'hbfbb940c, 32'hbed885b8} /* (13, 20, 30) {real, imag} */,
  {32'h3ff41e99, 32'h3f48c0eb} /* (13, 20, 29) {real, imag} */,
  {32'hbfeba1f5, 32'hbe116c39} /* (13, 20, 28) {real, imag} */,
  {32'h3f93d534, 32'hbe561239} /* (13, 20, 27) {real, imag} */,
  {32'hbfabc57c, 32'h3cea22f9} /* (13, 20, 26) {real, imag} */,
  {32'h3fac4d7e, 32'hc083f835} /* (13, 20, 25) {real, imag} */,
  {32'hbf71328d, 32'h3f2ddcfe} /* (13, 20, 24) {real, imag} */,
  {32'h3fc24ae2, 32'h3f8537eb} /* (13, 20, 23) {real, imag} */,
  {32'h4039039c, 32'hbfa7869b} /* (13, 20, 22) {real, imag} */,
  {32'hbf5eaa59, 32'h3fd92540} /* (13, 20, 21) {real, imag} */,
  {32'hbf0cd96b, 32'hbe906ea9} /* (13, 20, 20) {real, imag} */,
  {32'h3f6e77b4, 32'hbfb30f0c} /* (13, 20, 19) {real, imag} */,
  {32'hbe2ecb74, 32'h400e015b} /* (13, 20, 18) {real, imag} */,
  {32'h3f01d1d2, 32'hbf9f6df6} /* (13, 20, 17) {real, imag} */,
  {32'h3f576731, 32'hbf2bdbb2} /* (13, 20, 16) {real, imag} */,
  {32'h3fe10d94, 32'hbfa26324} /* (13, 20, 15) {real, imag} */,
  {32'h3f96b06c, 32'hbf154edc} /* (13, 20, 14) {real, imag} */,
  {32'h3e4b886d, 32'h3f7068fd} /* (13, 20, 13) {real, imag} */,
  {32'h3fe20a7f, 32'h3e78b6e6} /* (13, 20, 12) {real, imag} */,
  {32'hbfc29bd1, 32'h4050b69e} /* (13, 20, 11) {real, imag} */,
  {32'hbfce5e24, 32'h3f9bc9ed} /* (13, 20, 10) {real, imag} */,
  {32'hbf011c04, 32'hbfae3da3} /* (13, 20, 9) {real, imag} */,
  {32'h3fd0a68a, 32'hbf93aee0} /* (13, 20, 8) {real, imag} */,
  {32'hbe64c248, 32'h3f8469b5} /* (13, 20, 7) {real, imag} */,
  {32'h40636ecf, 32'h3ee31699} /* (13, 20, 6) {real, imag} */,
  {32'hc01eef89, 32'hbf97d24e} /* (13, 20, 5) {real, imag} */,
  {32'hbf0419d9, 32'h3f64e045} /* (13, 20, 4) {real, imag} */,
  {32'h402ae09a, 32'hbdd7c69a} /* (13, 20, 3) {real, imag} */,
  {32'hbf52eb1b, 32'h3fe3473c} /* (13, 20, 2) {real, imag} */,
  {32'hbf5c55e2, 32'hbf7635b9} /* (13, 20, 1) {real, imag} */,
  {32'hbf23a953, 32'h3f8b44af} /* (13, 20, 0) {real, imag} */,
  {32'hbdfcfd58, 32'hbfac982b} /* (13, 19, 31) {real, imag} */,
  {32'hbe33bd2b, 32'hbe957a55} /* (13, 19, 30) {real, imag} */,
  {32'h3ed8166b, 32'h3f1e9bf1} /* (13, 19, 29) {real, imag} */,
  {32'h3f4f0c68, 32'hbeec9da3} /* (13, 19, 28) {real, imag} */,
  {32'hc02436ac, 32'hbfa53524} /* (13, 19, 27) {real, imag} */,
  {32'h3fc66bc3, 32'h3f7a1418} /* (13, 19, 26) {real, imag} */,
  {32'hc02a591a, 32'hbfa44010} /* (13, 19, 25) {real, imag} */,
  {32'h3f3696b9, 32'hbf6cb34b} /* (13, 19, 24) {real, imag} */,
  {32'h3ee05e4d, 32'h3fd9e257} /* (13, 19, 23) {real, imag} */,
  {32'hbf3ae4b2, 32'h3f11c999} /* (13, 19, 22) {real, imag} */,
  {32'hc00bf900, 32'h3dd36021} /* (13, 19, 21) {real, imag} */,
  {32'hbea6095b, 32'h3c938828} /* (13, 19, 20) {real, imag} */,
  {32'h3f2c5fc4, 32'hbc7e2968} /* (13, 19, 19) {real, imag} */,
  {32'hbfc3db61, 32'hc01218c3} /* (13, 19, 18) {real, imag} */,
  {32'h40515ae3, 32'hbf52bc0a} /* (13, 19, 17) {real, imag} */,
  {32'hbf5af67e, 32'h3f8a2583} /* (13, 19, 16) {real, imag} */,
  {32'hbed70870, 32'hbe95b68d} /* (13, 19, 15) {real, imag} */,
  {32'hc012e86d, 32'h3eddab12} /* (13, 19, 14) {real, imag} */,
  {32'hbde17dc0, 32'hbfe687e9} /* (13, 19, 13) {real, imag} */,
  {32'hbf78f7fd, 32'h3f9cb760} /* (13, 19, 12) {real, imag} */,
  {32'h3fc67818, 32'h404494d1} /* (13, 19, 11) {real, imag} */,
  {32'hbdcf7ad6, 32'hc0123641} /* (13, 19, 10) {real, imag} */,
  {32'h3fa9c1a6, 32'hbfae7845} /* (13, 19, 9) {real, imag} */,
  {32'hbec5755b, 32'hc01ae52c} /* (13, 19, 8) {real, imag} */,
  {32'h3e98a113, 32'h4026248a} /* (13, 19, 7) {real, imag} */,
  {32'h3eb36d49, 32'hbdceed45} /* (13, 19, 6) {real, imag} */,
  {32'hbf0985d8, 32'hbe9675c6} /* (13, 19, 5) {real, imag} */,
  {32'hc00e3b89, 32'hbf4bd277} /* (13, 19, 4) {real, imag} */,
  {32'hc040e9a1, 32'hbf82214a} /* (13, 19, 3) {real, imag} */,
  {32'h3f3d35d2, 32'h3f2532f0} /* (13, 19, 2) {real, imag} */,
  {32'h3f45979b, 32'hbff3b7ea} /* (13, 19, 1) {real, imag} */,
  {32'hbf933048, 32'hbfae7eac} /* (13, 19, 0) {real, imag} */,
  {32'hbe73f42e, 32'hbfb3014b} /* (13, 18, 31) {real, imag} */,
  {32'h3ee9ad22, 32'hbfa87307} /* (13, 18, 30) {real, imag} */,
  {32'hbfe30497, 32'hbf026881} /* (13, 18, 29) {real, imag} */,
  {32'h3ea38a97, 32'h3f438e22} /* (13, 18, 28) {real, imag} */,
  {32'hbf68b3e3, 32'hc0173fd6} /* (13, 18, 27) {real, imag} */,
  {32'h3ffad4e1, 32'hbec8396b} /* (13, 18, 26) {real, imag} */,
  {32'h401d00c6, 32'hc02c482e} /* (13, 18, 25) {real, imag} */,
  {32'h40193025, 32'hc014f584} /* (13, 18, 24) {real, imag} */,
  {32'h3f8a0fe2, 32'h401b58e3} /* (13, 18, 23) {real, imag} */,
  {32'hc0bbd7bc, 32'h3f1d7e9a} /* (13, 18, 22) {real, imag} */,
  {32'h3e29de31, 32'hbed90493} /* (13, 18, 21) {real, imag} */,
  {32'hbfcd16fe, 32'hbf439c14} /* (13, 18, 20) {real, imag} */,
  {32'hbfa5fef5, 32'h3fa32849} /* (13, 18, 19) {real, imag} */,
  {32'hbe50b200, 32'hbfa7be6e} /* (13, 18, 18) {real, imag} */,
  {32'h3f07807c, 32'h3dc11487} /* (13, 18, 17) {real, imag} */,
  {32'h3fdbcfac, 32'h400b32b7} /* (13, 18, 16) {real, imag} */,
  {32'h3f46cc17, 32'h3fab0647} /* (13, 18, 15) {real, imag} */,
  {32'hc0138fbd, 32'hbfec5fc5} /* (13, 18, 14) {real, imag} */,
  {32'h3f238c42, 32'hbfad1cae} /* (13, 18, 13) {real, imag} */,
  {32'hbfc3b41c, 32'hbfab2d64} /* (13, 18, 12) {real, imag} */,
  {32'hc05e0a65, 32'h40179fcf} /* (13, 18, 11) {real, imag} */,
  {32'h3f40cac3, 32'h401ebcb2} /* (13, 18, 10) {real, imag} */,
  {32'hbfcbe129, 32'hbf948145} /* (13, 18, 9) {real, imag} */,
  {32'hbf2f9ebb, 32'hc0086762} /* (13, 18, 8) {real, imag} */,
  {32'hbe4445f8, 32'h401c3efa} /* (13, 18, 7) {real, imag} */,
  {32'h3ea233de, 32'h400452e2} /* (13, 18, 6) {real, imag} */,
  {32'h3f835aa0, 32'hbf8fecc5} /* (13, 18, 5) {real, imag} */,
  {32'h3fca4a76, 32'h3da439fc} /* (13, 18, 4) {real, imag} */,
  {32'hc013810f, 32'h40031a23} /* (13, 18, 3) {real, imag} */,
  {32'hc02b976e, 32'h3f138f63} /* (13, 18, 2) {real, imag} */,
  {32'h3d2d682d, 32'hbf000194} /* (13, 18, 1) {real, imag} */,
  {32'hbeae6f2f, 32'hbf949a4a} /* (13, 18, 0) {real, imag} */,
  {32'hbf237886, 32'h3e552452} /* (13, 17, 31) {real, imag} */,
  {32'h3f57503a, 32'hbfe04e83} /* (13, 17, 30) {real, imag} */,
  {32'h3efe6433, 32'h4062a024} /* (13, 17, 29) {real, imag} */,
  {32'h3f8ec325, 32'h3ef06e27} /* (13, 17, 28) {real, imag} */,
  {32'hbe44ea1e, 32'h3fc5c89f} /* (13, 17, 27) {real, imag} */,
  {32'hbf4032f7, 32'hbf1af2f5} /* (13, 17, 26) {real, imag} */,
  {32'hbf40c055, 32'h3f45da1a} /* (13, 17, 25) {real, imag} */,
  {32'h3e8852d8, 32'hbfa6c178} /* (13, 17, 24) {real, imag} */,
  {32'hbf2a19ec, 32'h3f4ff088} /* (13, 17, 23) {real, imag} */,
  {32'h3f845b5c, 32'hbdc495dc} /* (13, 17, 22) {real, imag} */,
  {32'h3f0a4dc9, 32'hbd9d5ccf} /* (13, 17, 21) {real, imag} */,
  {32'hbf6b3b1c, 32'hbeac2688} /* (13, 17, 20) {real, imag} */,
  {32'h3fbf2634, 32'hbfd189df} /* (13, 17, 19) {real, imag} */,
  {32'h401351d7, 32'h3e0d49af} /* (13, 17, 18) {real, imag} */,
  {32'h3ec5152c, 32'h3e74e783} /* (13, 17, 17) {real, imag} */,
  {32'hbf857067, 32'h3f94f879} /* (13, 17, 16) {real, imag} */,
  {32'hc036d731, 32'hbd1ea616} /* (13, 17, 15) {real, imag} */,
  {32'hbf80a0de, 32'hbc70b1e5} /* (13, 17, 14) {real, imag} */,
  {32'hbec48254, 32'hbd1b9b56} /* (13, 17, 13) {real, imag} */,
  {32'h3e6ceb2a, 32'hbf98cae2} /* (13, 17, 12) {real, imag} */,
  {32'h3fda5035, 32'hbda43e5a} /* (13, 17, 11) {real, imag} */,
  {32'h3fb01ac3, 32'hbd78c2c4} /* (13, 17, 10) {real, imag} */,
  {32'h3f2434da, 32'hbf47abd7} /* (13, 17, 9) {real, imag} */,
  {32'h3f16db45, 32'h3fa48eaa} /* (13, 17, 8) {real, imag} */,
  {32'h3fdd05be, 32'h3f0575fe} /* (13, 17, 7) {real, imag} */,
  {32'hbf83a557, 32'hbe5e8b25} /* (13, 17, 6) {real, imag} */,
  {32'hbf07d166, 32'h3e9c7114} /* (13, 17, 5) {real, imag} */,
  {32'hbf7a70fa, 32'hbf96271c} /* (13, 17, 4) {real, imag} */,
  {32'hc0268ab0, 32'h3f186a94} /* (13, 17, 3) {real, imag} */,
  {32'hbd0c06b6, 32'h3ec8438b} /* (13, 17, 2) {real, imag} */,
  {32'hbe3dcdf9, 32'h3faf6cf6} /* (13, 17, 1) {real, imag} */,
  {32'h3f46ced1, 32'hbe41b3c8} /* (13, 17, 0) {real, imag} */,
  {32'h3f0ff3c9, 32'h3d189fa1} /* (13, 16, 31) {real, imag} */,
  {32'h3fcaa806, 32'h3fe73e4a} /* (13, 16, 30) {real, imag} */,
  {32'hbf9680d5, 32'h3f071950} /* (13, 16, 29) {real, imag} */,
  {32'h3cf3009b, 32'h3f9cacf9} /* (13, 16, 28) {real, imag} */,
  {32'h3fc94ff9, 32'h400c07e5} /* (13, 16, 27) {real, imag} */,
  {32'h3f86ebaa, 32'h3e4b0fec} /* (13, 16, 26) {real, imag} */,
  {32'hbedbf7b9, 32'h40313432} /* (13, 16, 25) {real, imag} */,
  {32'hbf2f73c0, 32'hbf5c451e} /* (13, 16, 24) {real, imag} */,
  {32'hbf7434f2, 32'h40316357} /* (13, 16, 23) {real, imag} */,
  {32'hbfc34321, 32'hc00f59ac} /* (13, 16, 22) {real, imag} */,
  {32'h4008460d, 32'hbf31ba2e} /* (13, 16, 21) {real, imag} */,
  {32'h3ee3fb54, 32'h3e5af1d4} /* (13, 16, 20) {real, imag} */,
  {32'h40085193, 32'h3f7956e4} /* (13, 16, 19) {real, imag} */,
  {32'hbc253161, 32'h40577551} /* (13, 16, 18) {real, imag} */,
  {32'hbe0791e9, 32'hbf1b8bd0} /* (13, 16, 17) {real, imag} */,
  {32'hbf20bb1f, 32'hbf9a96fe} /* (13, 16, 16) {real, imag} */,
  {32'h3f1b60f5, 32'hbf166301} /* (13, 16, 15) {real, imag} */,
  {32'hbf8d6e5a, 32'h3efe03c4} /* (13, 16, 14) {real, imag} */,
  {32'hbfce3366, 32'h3d3ee92f} /* (13, 16, 13) {real, imag} */,
  {32'hc010e3fb, 32'h3dd69703} /* (13, 16, 12) {real, imag} */,
  {32'hbee026f1, 32'hc0029e39} /* (13, 16, 11) {real, imag} */,
  {32'hbf0d57c0, 32'hbf76732d} /* (13, 16, 10) {real, imag} */,
  {32'h4020162c, 32'h3f914218} /* (13, 16, 9) {real, imag} */,
  {32'hbe8447c4, 32'h3ec05fd9} /* (13, 16, 8) {real, imag} */,
  {32'hbf1c8f39, 32'h3ff7e58f} /* (13, 16, 7) {real, imag} */,
  {32'h3f1dd661, 32'hbfb7864f} /* (13, 16, 6) {real, imag} */,
  {32'h3d9fa8f6, 32'hbfd47da6} /* (13, 16, 5) {real, imag} */,
  {32'hbe3ddd05, 32'hbf8b9da8} /* (13, 16, 4) {real, imag} */,
  {32'h3e554fb9, 32'hbf42fe85} /* (13, 16, 3) {real, imag} */,
  {32'h4003dc6c, 32'hbfc2f38c} /* (13, 16, 2) {real, imag} */,
  {32'hbf6ff833, 32'h3eecdc92} /* (13, 16, 1) {real, imag} */,
  {32'h3f3885e1, 32'hbf780bfb} /* (13, 16, 0) {real, imag} */,
  {32'hbf9854c8, 32'hbf43a710} /* (13, 15, 31) {real, imag} */,
  {32'h3da8a69a, 32'hbdf73aaa} /* (13, 15, 30) {real, imag} */,
  {32'h3f58ed2a, 32'h3efaddba} /* (13, 15, 29) {real, imag} */,
  {32'h400a8685, 32'hbe01a3e7} /* (13, 15, 28) {real, imag} */,
  {32'h3f7eb95d, 32'h3ee6d227} /* (13, 15, 27) {real, imag} */,
  {32'hbf18a1de, 32'hbf3dcf7e} /* (13, 15, 26) {real, imag} */,
  {32'hbef0a80a, 32'h3f871cea} /* (13, 15, 25) {real, imag} */,
  {32'h3f5465dc, 32'h3f231496} /* (13, 15, 24) {real, imag} */,
  {32'hbca6ca54, 32'h3dc7d157} /* (13, 15, 23) {real, imag} */,
  {32'hbfb6bf5e, 32'h3e7b4f0e} /* (13, 15, 22) {real, imag} */,
  {32'h3f6c1846, 32'h3f8e3129} /* (13, 15, 21) {real, imag} */,
  {32'hc008e09c, 32'h3fb9ae5a} /* (13, 15, 20) {real, imag} */,
  {32'h3ee6e1e4, 32'h3fb0f647} /* (13, 15, 19) {real, imag} */,
  {32'hbf5c2129, 32'h3e649832} /* (13, 15, 18) {real, imag} */,
  {32'h3f028724, 32'h3fb1db63} /* (13, 15, 17) {real, imag} */,
  {32'h3fbd2dce, 32'hbf4f5cbc} /* (13, 15, 16) {real, imag} */,
  {32'hbf94466c, 32'hc0263210} /* (13, 15, 15) {real, imag} */,
  {32'h3fac567d, 32'hbf2e8b4a} /* (13, 15, 14) {real, imag} */,
  {32'hbedf579c, 32'h3fba6c64} /* (13, 15, 13) {real, imag} */,
  {32'h3f874344, 32'h3f885b96} /* (13, 15, 12) {real, imag} */,
  {32'h3fa0f7f3, 32'h40305a14} /* (13, 15, 11) {real, imag} */,
  {32'h3ff0f5ba, 32'h3f1d9928} /* (13, 15, 10) {real, imag} */,
  {32'hc037dd7f, 32'hbf56c9bd} /* (13, 15, 9) {real, imag} */,
  {32'h3e89d2f3, 32'h3da0d87f} /* (13, 15, 8) {real, imag} */,
  {32'hbfcac17a, 32'hbfc1bb31} /* (13, 15, 7) {real, imag} */,
  {32'hbfa6db22, 32'h3f880834} /* (13, 15, 6) {real, imag} */,
  {32'h3fc2c4ee, 32'hbf9d03ff} /* (13, 15, 5) {real, imag} */,
  {32'h3fd022c6, 32'h3f39e560} /* (13, 15, 4) {real, imag} */,
  {32'hbfd27acd, 32'h3fe5f0c9} /* (13, 15, 3) {real, imag} */,
  {32'hbdbeca8f, 32'hbfc103fd} /* (13, 15, 2) {real, imag} */,
  {32'hbf80db8b, 32'hbf4745ab} /* (13, 15, 1) {real, imag} */,
  {32'h3ffc6568, 32'hbebaed0b} /* (13, 15, 0) {real, imag} */,
  {32'hbff3e427, 32'h3e947c78} /* (13, 14, 31) {real, imag} */,
  {32'h3f6353d8, 32'hc01740c0} /* (13, 14, 30) {real, imag} */,
  {32'h3fff4a89, 32'h3fb42bb6} /* (13, 14, 29) {real, imag} */,
  {32'hbf963353, 32'hbd54ea70} /* (13, 14, 28) {real, imag} */,
  {32'hbf9fd329, 32'hbd54d256} /* (13, 14, 27) {real, imag} */,
  {32'hbe09f012, 32'h3ff0a386} /* (13, 14, 26) {real, imag} */,
  {32'hbd5bf6e9, 32'hbfcc26c5} /* (13, 14, 25) {real, imag} */,
  {32'hbe35a9ac, 32'h3eafb979} /* (13, 14, 24) {real, imag} */,
  {32'h400901e3, 32'h3fc06b3b} /* (13, 14, 23) {real, imag} */,
  {32'h3fbd116e, 32'hbeebf94a} /* (13, 14, 22) {real, imag} */,
  {32'h3fac868e, 32'hc017b78d} /* (13, 14, 21) {real, imag} */,
  {32'h3f9a852d, 32'hbfc5c3a6} /* (13, 14, 20) {real, imag} */,
  {32'hc02677ae, 32'hbf312a25} /* (13, 14, 19) {real, imag} */,
  {32'hbd8637b3, 32'h3d72a82e} /* (13, 14, 18) {real, imag} */,
  {32'h3ea8f39e, 32'hbf5c4203} /* (13, 14, 17) {real, imag} */,
  {32'h3f56e660, 32'h3ff3598d} /* (13, 14, 16) {real, imag} */,
  {32'hbdf5c81d, 32'hbf49a37f} /* (13, 14, 15) {real, imag} */,
  {32'h3f1ea056, 32'h3fd4be8c} /* (13, 14, 14) {real, imag} */,
  {32'hbe3d624e, 32'hc013b136} /* (13, 14, 13) {real, imag} */,
  {32'h3ecec165, 32'hbfa2ea9a} /* (13, 14, 12) {real, imag} */,
  {32'h3feb6b28, 32'h3fafd231} /* (13, 14, 11) {real, imag} */,
  {32'hbfe6239c, 32'hbf43f5ce} /* (13, 14, 10) {real, imag} */,
  {32'hbf59376c, 32'h3f3626dd} /* (13, 14, 9) {real, imag} */,
  {32'h3ff87ec6, 32'hbfe8c47a} /* (13, 14, 8) {real, imag} */,
  {32'h3f2baa71, 32'hbf813474} /* (13, 14, 7) {real, imag} */,
  {32'h3efc260b, 32'hbf2293b1} /* (13, 14, 6) {real, imag} */,
  {32'h3f883a57, 32'hbeadb709} /* (13, 14, 5) {real, imag} */,
  {32'hbf882183, 32'hbf449f52} /* (13, 14, 4) {real, imag} */,
  {32'h3f3f06af, 32'hbf498a12} /* (13, 14, 3) {real, imag} */,
  {32'hbf7b1a8c, 32'h3e88a067} /* (13, 14, 2) {real, imag} */,
  {32'hbd977fe2, 32'h3fba3804} /* (13, 14, 1) {real, imag} */,
  {32'h3fe2d336, 32'hbfd7f5dd} /* (13, 14, 0) {real, imag} */,
  {32'hbfe1c129, 32'h3fbf4de9} /* (13, 13, 31) {real, imag} */,
  {32'h401f3a67, 32'h3e862cb9} /* (13, 13, 30) {real, imag} */,
  {32'hc033113e, 32'hc02b0751} /* (13, 13, 29) {real, imag} */,
  {32'hbfd9f33b, 32'hbf9e772f} /* (13, 13, 28) {real, imag} */,
  {32'h3dde66eb, 32'hc04ace5c} /* (13, 13, 27) {real, imag} */,
  {32'h3f4a93e5, 32'h40315689} /* (13, 13, 26) {real, imag} */,
  {32'hbf553842, 32'hbfbb4369} /* (13, 13, 25) {real, imag} */,
  {32'h4024f532, 32'h3fe2133d} /* (13, 13, 24) {real, imag} */,
  {32'hc0467609, 32'hbfc82641} /* (13, 13, 23) {real, imag} */,
  {32'hbfa31857, 32'h400e8f7d} /* (13, 13, 22) {real, imag} */,
  {32'hbfa314b3, 32'h400993b6} /* (13, 13, 21) {real, imag} */,
  {32'h3f50847b, 32'hc001b31c} /* (13, 13, 20) {real, imag} */,
  {32'hbfde6fce, 32'hbf90b982} /* (13, 13, 19) {real, imag} */,
  {32'hbf2d29af, 32'hbf601dec} /* (13, 13, 18) {real, imag} */,
  {32'hbed82108, 32'hbe749a28} /* (13, 13, 17) {real, imag} */,
  {32'h3fa10963, 32'hbfedd0f6} /* (13, 13, 16) {real, imag} */,
  {32'hbfb9a974, 32'h400c8f15} /* (13, 13, 15) {real, imag} */,
  {32'hbfb03540, 32'hbffe24bb} /* (13, 13, 14) {real, imag} */,
  {32'h4065a4eb, 32'hbdc3b4ed} /* (13, 13, 13) {real, imag} */,
  {32'hbea4e538, 32'h3f96091e} /* (13, 13, 12) {real, imag} */,
  {32'hc0164bf9, 32'hbe80efa1} /* (13, 13, 11) {real, imag} */,
  {32'h3f936d78, 32'hbf048822} /* (13, 13, 10) {real, imag} */,
  {32'hbfe8f661, 32'hbddeffdc} /* (13, 13, 9) {real, imag} */,
  {32'hc03df95f, 32'hbfae26e4} /* (13, 13, 8) {real, imag} */,
  {32'h3f602965, 32'h4003fb9f} /* (13, 13, 7) {real, imag} */,
  {32'h4074bc1c, 32'hc00d7979} /* (13, 13, 6) {real, imag} */,
  {32'h3fb4a374, 32'h3fc436bc} /* (13, 13, 5) {real, imag} */,
  {32'h3e9e5014, 32'hbfb84e8d} /* (13, 13, 4) {real, imag} */,
  {32'h3f80efc8, 32'h3f0dcac4} /* (13, 13, 3) {real, imag} */,
  {32'h3fadc6f4, 32'hbfc7b3ec} /* (13, 13, 2) {real, imag} */,
  {32'h3fd97e4e, 32'h3e08820d} /* (13, 13, 1) {real, imag} */,
  {32'hc0074a2b, 32'hbfac5356} /* (13, 13, 0) {real, imag} */,
  {32'h3df9ce5f, 32'hbecef558} /* (13, 12, 31) {real, imag} */,
  {32'hbfe8bc01, 32'h3f736ed4} /* (13, 12, 30) {real, imag} */,
  {32'h3e3a74c8, 32'hbf15cbe3} /* (13, 12, 29) {real, imag} */,
  {32'h3f71683f, 32'hbf1a72a3} /* (13, 12, 28) {real, imag} */,
  {32'h3f751ad7, 32'h3ffa035f} /* (13, 12, 27) {real, imag} */,
  {32'hc049b980, 32'h3e84cbdb} /* (13, 12, 26) {real, imag} */,
  {32'h408bc49c, 32'hbe6e3f76} /* (13, 12, 25) {real, imag} */,
  {32'hbfe53bdd, 32'hbde56009} /* (13, 12, 24) {real, imag} */,
  {32'h3fef5214, 32'h3c081609} /* (13, 12, 23) {real, imag} */,
  {32'h3ffad3c9, 32'h3e59c2a9} /* (13, 12, 22) {real, imag} */,
  {32'h402ca14e, 32'hc0115f64} /* (13, 12, 21) {real, imag} */,
  {32'h3fb0b3ef, 32'h3f470bda} /* (13, 12, 20) {real, imag} */,
  {32'hbea9a16c, 32'hbfdeeb59} /* (13, 12, 19) {real, imag} */,
  {32'hbfdb175d, 32'h3fa34eea} /* (13, 12, 18) {real, imag} */,
  {32'h3f7b5c52, 32'h3ff01bca} /* (13, 12, 17) {real, imag} */,
  {32'hbf00a307, 32'h3f762eb9} /* (13, 12, 16) {real, imag} */,
  {32'h3f8bf1b8, 32'hc06eea54} /* (13, 12, 15) {real, imag} */,
  {32'h3f8d457d, 32'h3e09753e} /* (13, 12, 14) {real, imag} */,
  {32'hbfa76d94, 32'hbf4e547a} /* (13, 12, 13) {real, imag} */,
  {32'h40552f89, 32'h3f487b8e} /* (13, 12, 12) {real, imag} */,
  {32'h404c7f5b, 32'hbf13a5e0} /* (13, 12, 11) {real, imag} */,
  {32'hbedaa8e8, 32'h3ea37902} /* (13, 12, 10) {real, imag} */,
  {32'hbe583f65, 32'h3e4a2231} /* (13, 12, 9) {real, imag} */,
  {32'hbee2a07b, 32'hbfff0568} /* (13, 12, 8) {real, imag} */,
  {32'h3fae155b, 32'h3e8e1909} /* (13, 12, 7) {real, imag} */,
  {32'hbeb0fa30, 32'h3ea41465} /* (13, 12, 6) {real, imag} */,
  {32'hbf84deee, 32'h3e229aa6} /* (13, 12, 5) {real, imag} */,
  {32'hc0623927, 32'h3f570449} /* (13, 12, 4) {real, imag} */,
  {32'h3e9df65a, 32'hc0760909} /* (13, 12, 3) {real, imag} */,
  {32'h3fc927fa, 32'hbf2fe65a} /* (13, 12, 2) {real, imag} */,
  {32'h401b7dfa, 32'h3fadb0ef} /* (13, 12, 1) {real, imag} */,
  {32'hbfbfe181, 32'h3f969a3a} /* (13, 12, 0) {real, imag} */,
  {32'h3ee19ea7, 32'h3ec691a5} /* (13, 11, 31) {real, imag} */,
  {32'h3f2db778, 32'hbf64d3fe} /* (13, 11, 30) {real, imag} */,
  {32'hbf489c71, 32'h3f234598} /* (13, 11, 29) {real, imag} */,
  {32'h3f281d7f, 32'hbf0795e9} /* (13, 11, 28) {real, imag} */,
  {32'h3f704311, 32'h3c9ccfcd} /* (13, 11, 27) {real, imag} */,
  {32'h3f2fde4e, 32'h3f6815b6} /* (13, 11, 26) {real, imag} */,
  {32'hc00225d9, 32'hc0040c5b} /* (13, 11, 25) {real, imag} */,
  {32'hbf7c3765, 32'h3e875ea7} /* (13, 11, 24) {real, imag} */,
  {32'hc0bb86a6, 32'h3ebf3d3e} /* (13, 11, 23) {real, imag} */,
  {32'hc01b1335, 32'hbfccee60} /* (13, 11, 22) {real, imag} */,
  {32'hc0259ab9, 32'hbe8dbd41} /* (13, 11, 21) {real, imag} */,
  {32'h404645ec, 32'h3dcf8046} /* (13, 11, 20) {real, imag} */,
  {32'h3de559ad, 32'h3fb158e9} /* (13, 11, 19) {real, imag} */,
  {32'h402a3b6d, 32'h3f86985a} /* (13, 11, 18) {real, imag} */,
  {32'h3fe6c289, 32'hbfcf8b69} /* (13, 11, 17) {real, imag} */,
  {32'hbf85087e, 32'h3f252377} /* (13, 11, 16) {real, imag} */,
  {32'hbf737054, 32'hbf816476} /* (13, 11, 15) {real, imag} */,
  {32'h3f0d85b0, 32'h3f0b2515} /* (13, 11, 14) {real, imag} */,
  {32'h3fd50e94, 32'h3ebc220e} /* (13, 11, 13) {real, imag} */,
  {32'h3fa7d286, 32'h402703d1} /* (13, 11, 12) {real, imag} */,
  {32'h40235a64, 32'hc070dcb5} /* (13, 11, 11) {real, imag} */,
  {32'hbe672b65, 32'h3fc046f8} /* (13, 11, 10) {real, imag} */,
  {32'hbf9f0cb6, 32'h402819d8} /* (13, 11, 9) {real, imag} */,
  {32'hbfcc70b4, 32'hc03c162c} /* (13, 11, 8) {real, imag} */,
  {32'h3d4dafc1, 32'h3f4a0d2a} /* (13, 11, 7) {real, imag} */,
  {32'hc0946d3b, 32'h3ed970a0} /* (13, 11, 6) {real, imag} */,
  {32'hc08e8da5, 32'h3f68d3a1} /* (13, 11, 5) {real, imag} */,
  {32'hbf043c7b, 32'h3e640b7a} /* (13, 11, 4) {real, imag} */,
  {32'h4028502b, 32'hc015a05c} /* (13, 11, 3) {real, imag} */,
  {32'h3f61d6c5, 32'h3f860ac2} /* (13, 11, 2) {real, imag} */,
  {32'hbe7d1e0c, 32'hc030e11e} /* (13, 11, 1) {real, imag} */,
  {32'hbf2b8aae, 32'h3f9fe013} /* (13, 11, 0) {real, imag} */,
  {32'h3fd5df99, 32'h3fd7784c} /* (13, 10, 31) {real, imag} */,
  {32'hc00f549b, 32'h3e180029} /* (13, 10, 30) {real, imag} */,
  {32'hc00193c1, 32'hbec1d886} /* (13, 10, 29) {real, imag} */,
  {32'hc0997d10, 32'hbfeaccb9} /* (13, 10, 28) {real, imag} */,
  {32'h408d6831, 32'hbf26396e} /* (13, 10, 27) {real, imag} */,
  {32'h3e3925a8, 32'h3f940af7} /* (13, 10, 26) {real, imag} */,
  {32'h3fff0210, 32'h3f4df922} /* (13, 10, 25) {real, imag} */,
  {32'h3f1d94f2, 32'hc03549df} /* (13, 10, 24) {real, imag} */,
  {32'h3f53728b, 32'hc00ca96d} /* (13, 10, 23) {real, imag} */,
  {32'hbf53e341, 32'hc02a7d53} /* (13, 10, 22) {real, imag} */,
  {32'h3fc85fa8, 32'h4094cd68} /* (13, 10, 21) {real, imag} */,
  {32'h3f1f362d, 32'h40562599} /* (13, 10, 20) {real, imag} */,
  {32'h3ffb0c36, 32'hc03de546} /* (13, 10, 19) {real, imag} */,
  {32'hbf4660ce, 32'h400c9df1} /* (13, 10, 18) {real, imag} */,
  {32'hbea42b22, 32'hc021c2ee} /* (13, 10, 17) {real, imag} */,
  {32'h400d7380, 32'hbf24fc67} /* (13, 10, 16) {real, imag} */,
  {32'hbeef3738, 32'h3ebefdfd} /* (13, 10, 15) {real, imag} */,
  {32'hbfcd52ce, 32'hbe4b3c1e} /* (13, 10, 14) {real, imag} */,
  {32'h404d7484, 32'hbfcf4732} /* (13, 10, 13) {real, imag} */,
  {32'hc06f36cd, 32'hbf699f52} /* (13, 10, 12) {real, imag} */,
  {32'h3fc231a1, 32'hbde19939} /* (13, 10, 11) {real, imag} */,
  {32'h3e2bfcdd, 32'hbf5f0040} /* (13, 10, 10) {real, imag} */,
  {32'hbffc29a3, 32'hbffebd03} /* (13, 10, 9) {real, imag} */,
  {32'h3fec8ba9, 32'h3f922d42} /* (13, 10, 8) {real, imag} */,
  {32'h3fcdbe99, 32'hbf8a217a} /* (13, 10, 7) {real, imag} */,
  {32'hbf54e5a4, 32'h404a9e3c} /* (13, 10, 6) {real, imag} */,
  {32'hbea43f6b, 32'h40633d74} /* (13, 10, 5) {real, imag} */,
  {32'hbf95b8e1, 32'hc07d2e5e} /* (13, 10, 4) {real, imag} */,
  {32'h3fbd2040, 32'hbcdea7cc} /* (13, 10, 3) {real, imag} */,
  {32'hbfbf7c0d, 32'h3fd81d65} /* (13, 10, 2) {real, imag} */,
  {32'hbf4af6e6, 32'hbf59c725} /* (13, 10, 1) {real, imag} */,
  {32'h3fb4f637, 32'hc04e2337} /* (13, 10, 0) {real, imag} */,
  {32'hc0060f5b, 32'hc0704b5c} /* (13, 9, 31) {real, imag} */,
  {32'h3ebb4c94, 32'hbfddb6fe} /* (13, 9, 30) {real, imag} */,
  {32'hbe1f37ed, 32'h40982a76} /* (13, 9, 29) {real, imag} */,
  {32'hbfc0f4d0, 32'h3fa459cc} /* (13, 9, 28) {real, imag} */,
  {32'h3e3b2643, 32'h40054ae6} /* (13, 9, 27) {real, imag} */,
  {32'hc05e5538, 32'h3fe94258} /* (13, 9, 26) {real, imag} */,
  {32'hbf621b8d, 32'hbfda0bbb} /* (13, 9, 25) {real, imag} */,
  {32'h3f031fe9, 32'hc0820a6e} /* (13, 9, 24) {real, imag} */,
  {32'h3fe4ece5, 32'hc0512c40} /* (13, 9, 23) {real, imag} */,
  {32'h3fd48a44, 32'h403af0ea} /* (13, 9, 22) {real, imag} */,
  {32'h4089b701, 32'hbf847c62} /* (13, 9, 21) {real, imag} */,
  {32'h3f3b4ada, 32'hc0b97782} /* (13, 9, 20) {real, imag} */,
  {32'hbf1a9bd0, 32'h3f10eb1a} /* (13, 9, 19) {real, imag} */,
  {32'hc0347085, 32'h3eb69091} /* (13, 9, 18) {real, imag} */,
  {32'hbf00d6e3, 32'h3fe70ca6} /* (13, 9, 17) {real, imag} */,
  {32'h3f1c2661, 32'hbf678fd9} /* (13, 9, 16) {real, imag} */,
  {32'h3fad855a, 32'h4000a674} /* (13, 9, 15) {real, imag} */,
  {32'hbfbd9904, 32'hbf878673} /* (13, 9, 14) {real, imag} */,
  {32'hbe5e3601, 32'hbeb5a0eb} /* (13, 9, 13) {real, imag} */,
  {32'hbd36ed29, 32'hc00cdf11} /* (13, 9, 12) {real, imag} */,
  {32'h3f24d7bc, 32'hbee65785} /* (13, 9, 11) {real, imag} */,
  {32'hc02b8a45, 32'h3d91c9d6} /* (13, 9, 10) {real, imag} */,
  {32'h40451674, 32'hbdfd8d80} /* (13, 9, 9) {real, imag} */,
  {32'h40339858, 32'h3f92f4c2} /* (13, 9, 8) {real, imag} */,
  {32'hbf8a5d6a, 32'h3f22cfaf} /* (13, 9, 7) {real, imag} */,
  {32'hc00cd02f, 32'h3f9c877f} /* (13, 9, 6) {real, imag} */,
  {32'hc044201a, 32'h400f5374} /* (13, 9, 5) {real, imag} */,
  {32'h3eb3cbdc, 32'hbf5c279b} /* (13, 9, 4) {real, imag} */,
  {32'hbfe72e27, 32'hbfb88718} /* (13, 9, 3) {real, imag} */,
  {32'hc0258bf0, 32'hbeb08897} /* (13, 9, 2) {real, imag} */,
  {32'h402ae57e, 32'hbed2c271} /* (13, 9, 1) {real, imag} */,
  {32'hbfaa57ec, 32'h3e88b47a} /* (13, 9, 0) {real, imag} */,
  {32'h40022526, 32'hbf0b90c0} /* (13, 8, 31) {real, imag} */,
  {32'hc02afbc6, 32'h3f95d4ea} /* (13, 8, 30) {real, imag} */,
  {32'h403c77c9, 32'hc0207ec1} /* (13, 8, 29) {real, imag} */,
  {32'h400d5161, 32'hc0021caf} /* (13, 8, 28) {real, imag} */,
  {32'h3f62a1fd, 32'h3ee5f01d} /* (13, 8, 27) {real, imag} */,
  {32'h4032897b, 32'hbf9f025d} /* (13, 8, 26) {real, imag} */,
  {32'hbf85a304, 32'h3f507ae3} /* (13, 8, 25) {real, imag} */,
  {32'h3f05ab6a, 32'hbea51bca} /* (13, 8, 24) {real, imag} */,
  {32'h3f0b8017, 32'hc06bbd88} /* (13, 8, 23) {real, imag} */,
  {32'h3f744da6, 32'h3fa25abe} /* (13, 8, 22) {real, imag} */,
  {32'hc05d2f68, 32'h3f46b1e7} /* (13, 8, 21) {real, imag} */,
  {32'h3de33229, 32'h40112e18} /* (13, 8, 20) {real, imag} */,
  {32'hbfcaae43, 32'hc02671da} /* (13, 8, 19) {real, imag} */,
  {32'h3e910145, 32'h3e9953bb} /* (13, 8, 18) {real, imag} */,
  {32'hbe998c83, 32'hbfa9ea8d} /* (13, 8, 17) {real, imag} */,
  {32'h3c80a0fb, 32'h3cc4e8c1} /* (13, 8, 16) {real, imag} */,
  {32'h3f31f6e7, 32'h3f30bda6} /* (13, 8, 15) {real, imag} */,
  {32'hbff649b4, 32'hbfa755e2} /* (13, 8, 14) {real, imag} */,
  {32'hbfa386d9, 32'h40158260} /* (13, 8, 13) {real, imag} */,
  {32'h3ec371d0, 32'h40152cab} /* (13, 8, 12) {real, imag} */,
  {32'hbe9bbfee, 32'hc02c6f11} /* (13, 8, 11) {real, imag} */,
  {32'h402c9384, 32'hc05734ca} /* (13, 8, 10) {real, imag} */,
  {32'hbfc4cc84, 32'h3fe75624} /* (13, 8, 9) {real, imag} */,
  {32'h3d884931, 32'hbfdbb3f4} /* (13, 8, 8) {real, imag} */,
  {32'hbec28b77, 32'hbe539820} /* (13, 8, 7) {real, imag} */,
  {32'hbfacf580, 32'hbf78c3cc} /* (13, 8, 6) {real, imag} */,
  {32'hbfba8927, 32'h3fe2b499} /* (13, 8, 5) {real, imag} */,
  {32'hbbb96907, 32'h401a7133} /* (13, 8, 4) {real, imag} */,
  {32'hc04fa65d, 32'h3f612851} /* (13, 8, 3) {real, imag} */,
  {32'h3e6c0c4a, 32'hc0059c9b} /* (13, 8, 2) {real, imag} */,
  {32'h3eabf47a, 32'hbd95bdd2} /* (13, 8, 1) {real, imag} */,
  {32'h40254c0a, 32'hbf9adad2} /* (13, 8, 0) {real, imag} */,
  {32'h3f9a0939, 32'hbf6796dc} /* (13, 7, 31) {real, imag} */,
  {32'hbed2b684, 32'hbf99179d} /* (13, 7, 30) {real, imag} */,
  {32'hbf3d6d43, 32'hbdaa6315} /* (13, 7, 29) {real, imag} */,
  {32'h3f22ca7a, 32'hbf44dbfb} /* (13, 7, 28) {real, imag} */,
  {32'hbfeb69ae, 32'hbf78da98} /* (13, 7, 27) {real, imag} */,
  {32'hbc13e87f, 32'hbfe4dba6} /* (13, 7, 26) {real, imag} */,
  {32'hbfedbb0d, 32'h3f3c2eb9} /* (13, 7, 25) {real, imag} */,
  {32'hbdd8dcdf, 32'h3f1f21ba} /* (13, 7, 24) {real, imag} */,
  {32'hbf125002, 32'hbfac41c1} /* (13, 7, 23) {real, imag} */,
  {32'h3f89e65d, 32'hbf98b75d} /* (13, 7, 22) {real, imag} */,
  {32'h4038e56c, 32'h400e3212} /* (13, 7, 21) {real, imag} */,
  {32'hc000da1a, 32'h3e83a415} /* (13, 7, 20) {real, imag} */,
  {32'hc043bc1e, 32'hbdbdb9da} /* (13, 7, 19) {real, imag} */,
  {32'h3fb052eb, 32'hbf81482b} /* (13, 7, 18) {real, imag} */,
  {32'hbe0e2f76, 32'hbca7175c} /* (13, 7, 17) {real, imag} */,
  {32'h40021f9d, 32'h3fa05372} /* (13, 7, 16) {real, imag} */,
  {32'h3eaf7b10, 32'h3ef59fcb} /* (13, 7, 15) {real, imag} */,
  {32'h3f13cd23, 32'hc016f46f} /* (13, 7, 14) {real, imag} */,
  {32'h3e4c8573, 32'h3ee9d413} /* (13, 7, 13) {real, imag} */,
  {32'h3f8ac1fd, 32'h3f94f8e2} /* (13, 7, 12) {real, imag} */,
  {32'hbfa43007, 32'hc0347249} /* (13, 7, 11) {real, imag} */,
  {32'hbf29e6fb, 32'h40016ce5} /* (13, 7, 10) {real, imag} */,
  {32'hbd9345c3, 32'h4081cc57} /* (13, 7, 9) {real, imag} */,
  {32'hbe8bfc60, 32'hbfe4aef6} /* (13, 7, 8) {real, imag} */,
  {32'h405845a3, 32'hc08696dc} /* (13, 7, 7) {real, imag} */,
  {32'h3f13642a, 32'h3f93ec52} /* (13, 7, 6) {real, imag} */,
  {32'hbe7a7918, 32'h402f817a} /* (13, 7, 5) {real, imag} */,
  {32'h3f19002d, 32'hbed8e2b8} /* (13, 7, 4) {real, imag} */,
  {32'hbf2931b7, 32'h3ea7d3be} /* (13, 7, 3) {real, imag} */,
  {32'hc05606da, 32'h3f906d0e} /* (13, 7, 2) {real, imag} */,
  {32'h400a54cf, 32'h3f4f8662} /* (13, 7, 1) {real, imag} */,
  {32'hc018a51c, 32'hbf7eb79b} /* (13, 7, 0) {real, imag} */,
  {32'hc00d90d1, 32'h3f2fa8e4} /* (13, 6, 31) {real, imag} */,
  {32'hbfb8e03a, 32'h401a8681} /* (13, 6, 30) {real, imag} */,
  {32'h3f285495, 32'hbf879f68} /* (13, 6, 29) {real, imag} */,
  {32'hbf447f03, 32'h3fe5a1b6} /* (13, 6, 28) {real, imag} */,
  {32'h3f4a48bb, 32'hbfeca2cc} /* (13, 6, 27) {real, imag} */,
  {32'hbfb1ac2d, 32'hc0252143} /* (13, 6, 26) {real, imag} */,
  {32'hbedb604c, 32'h3fb0d238} /* (13, 6, 25) {real, imag} */,
  {32'hc02cadfe, 32'hc0b56797} /* (13, 6, 24) {real, imag} */,
  {32'h401ac73a, 32'hc01786f6} /* (13, 6, 23) {real, imag} */,
  {32'hbf504b96, 32'h3d9e6e5c} /* (13, 6, 22) {real, imag} */,
  {32'h3f129ffd, 32'h3f24134a} /* (13, 6, 21) {real, imag} */,
  {32'hbe5bf036, 32'hbe4ae801} /* (13, 6, 20) {real, imag} */,
  {32'h4007ab9c, 32'h408b60be} /* (13, 6, 19) {real, imag} */,
  {32'h3fd44997, 32'hbfcf8dc3} /* (13, 6, 18) {real, imag} */,
  {32'hbff1f211, 32'h3e946595} /* (13, 6, 17) {real, imag} */,
  {32'hbf27fd27, 32'h3ebc62a3} /* (13, 6, 16) {real, imag} */,
  {32'hc00b16b2, 32'hc04346ca} /* (13, 6, 15) {real, imag} */,
  {32'h4002352a, 32'h3de82ff1} /* (13, 6, 14) {real, imag} */,
  {32'h3f95c385, 32'h3f2d2c32} /* (13, 6, 13) {real, imag} */,
  {32'h3f2f94bc, 32'hbf5df98c} /* (13, 6, 12) {real, imag} */,
  {32'hbfe25e40, 32'h401477e1} /* (13, 6, 11) {real, imag} */,
  {32'hbf62d741, 32'hc0056fbd} /* (13, 6, 10) {real, imag} */,
  {32'h3fec594e, 32'hbfd68576} /* (13, 6, 9) {real, imag} */,
  {32'hc0123c29, 32'hbf8ca6dc} /* (13, 6, 8) {real, imag} */,
  {32'hbf1b1131, 32'h3ff58259} /* (13, 6, 7) {real, imag} */,
  {32'h3fb16526, 32'h4042d155} /* (13, 6, 6) {real, imag} */,
  {32'h402dd21b, 32'h3eb99221} /* (13, 6, 5) {real, imag} */,
  {32'hbfc0af12, 32'hbee594c9} /* (13, 6, 4) {real, imag} */,
  {32'hbfcf8705, 32'hbe4bf5e2} /* (13, 6, 3) {real, imag} */,
  {32'h4048ba89, 32'hbfcf02d7} /* (13, 6, 2) {real, imag} */,
  {32'h3dd11308, 32'hbef2c552} /* (13, 6, 1) {real, imag} */,
  {32'h3f972bce, 32'h3f977ee5} /* (13, 6, 0) {real, imag} */,
  {32'h3e9df34d, 32'hbfc79c9a} /* (13, 5, 31) {real, imag} */,
  {32'h3fc425dd, 32'hc000a02c} /* (13, 5, 30) {real, imag} */,
  {32'hbf5ed454, 32'hbfe24350} /* (13, 5, 29) {real, imag} */,
  {32'hbf8b7d65, 32'h3fba37ed} /* (13, 5, 28) {real, imag} */,
  {32'hbf827f03, 32'h3ddc344f} /* (13, 5, 27) {real, imag} */,
  {32'h3db14a91, 32'h3f4bc184} /* (13, 5, 26) {real, imag} */,
  {32'hbfd8ad18, 32'hbf6db43e} /* (13, 5, 25) {real, imag} */,
  {32'hc00c1fa3, 32'h3febe8ea} /* (13, 5, 24) {real, imag} */,
  {32'h3d411437, 32'h3f45ea5e} /* (13, 5, 23) {real, imag} */,
  {32'hc06e59a6, 32'hc03cff64} /* (13, 5, 22) {real, imag} */,
  {32'hc073f807, 32'h400a7406} /* (13, 5, 21) {real, imag} */,
  {32'hbeff8c18, 32'hbfa49b34} /* (13, 5, 20) {real, imag} */,
  {32'hc0085a9a, 32'hbf201f61} /* (13, 5, 19) {real, imag} */,
  {32'hbeea2f3e, 32'hbee9ae43} /* (13, 5, 18) {real, imag} */,
  {32'hbf991ebf, 32'h3f3a9619} /* (13, 5, 17) {real, imag} */,
  {32'h3fe8e2ab, 32'h3f18c676} /* (13, 5, 16) {real, imag} */,
  {32'h3e5f6051, 32'h3f9f9914} /* (13, 5, 15) {real, imag} */,
  {32'h40025853, 32'hbd92e46e} /* (13, 5, 14) {real, imag} */,
  {32'h3f03c398, 32'hbf30870d} /* (13, 5, 13) {real, imag} */,
  {32'hbfbd67a4, 32'hbfe0064d} /* (13, 5, 12) {real, imag} */,
  {32'hc0714c9d, 32'hbfc55bfe} /* (13, 5, 11) {real, imag} */,
  {32'hbf7aa3bb, 32'hbec8e78b} /* (13, 5, 10) {real, imag} */,
  {32'hbfd8c696, 32'h3e8904c4} /* (13, 5, 9) {real, imag} */,
  {32'h40301ed7, 32'hbf8d2f6d} /* (13, 5, 8) {real, imag} */,
  {32'hc08cda59, 32'hc0188e12} /* (13, 5, 7) {real, imag} */,
  {32'h40b0332c, 32'h3e1601a8} /* (13, 5, 6) {real, imag} */,
  {32'h3e2fa555, 32'h3ada68e1} /* (13, 5, 5) {real, imag} */,
  {32'h3f57beca, 32'h3e086c00} /* (13, 5, 4) {real, imag} */,
  {32'h40709f2f, 32'h3ecbe447} /* (13, 5, 3) {real, imag} */,
  {32'h3e35d7e1, 32'h40277c61} /* (13, 5, 2) {real, imag} */,
  {32'hbfab5413, 32'h3fee8417} /* (13, 5, 1) {real, imag} */,
  {32'h401307d8, 32'hbf28c4b8} /* (13, 5, 0) {real, imag} */,
  {32'h3f26cdf2, 32'hbfdce42d} /* (13, 4, 31) {real, imag} */,
  {32'hbfaa2afd, 32'h40145d43} /* (13, 4, 30) {real, imag} */,
  {32'h3f8bcae2, 32'h3eeff98f} /* (13, 4, 29) {real, imag} */,
  {32'h3fce1d81, 32'hbfd79b52} /* (13, 4, 28) {real, imag} */,
  {32'hbfd19c68, 32'hbff28d11} /* (13, 4, 27) {real, imag} */,
  {32'hbe122b31, 32'h3face116} /* (13, 4, 26) {real, imag} */,
  {32'h3f389705, 32'hbf4f9e41} /* (13, 4, 25) {real, imag} */,
  {32'h3f690ed0, 32'hbf516cb9} /* (13, 4, 24) {real, imag} */,
  {32'h3f544f22, 32'hbfe04af2} /* (13, 4, 23) {real, imag} */,
  {32'h3f237385, 32'hbe9b9326} /* (13, 4, 22) {real, imag} */,
  {32'h3eec4060, 32'h3f1a2f4b} /* (13, 4, 21) {real, imag} */,
  {32'hbfbb29a3, 32'hbf4b5269} /* (13, 4, 20) {real, imag} */,
  {32'h3f68ad1c, 32'hbf3098dc} /* (13, 4, 19) {real, imag} */,
  {32'h3e09e542, 32'hc039ad84} /* (13, 4, 18) {real, imag} */,
  {32'hbf91525f, 32'h3f796df4} /* (13, 4, 17) {real, imag} */,
  {32'h3f6e1cd1, 32'h3e9e2942} /* (13, 4, 16) {real, imag} */,
  {32'hbe5f330f, 32'h3ec80b1b} /* (13, 4, 15) {real, imag} */,
  {32'h3ec0d176, 32'h3f289496} /* (13, 4, 14) {real, imag} */,
  {32'h400554bb, 32'h3fcb21d8} /* (13, 4, 13) {real, imag} */,
  {32'hbd5cfd2f, 32'hbfa0f563} /* (13, 4, 12) {real, imag} */,
  {32'h3e87c2f0, 32'hbfa45970} /* (13, 4, 11) {real, imag} */,
  {32'hbf918ada, 32'h3fedf3f0} /* (13, 4, 10) {real, imag} */,
  {32'h3f298d74, 32'hbc9b8c57} /* (13, 4, 9) {real, imag} */,
  {32'hbc8c022f, 32'hc0268f1a} /* (13, 4, 8) {real, imag} */,
  {32'h3f7984fb, 32'hbf4ab943} /* (13, 4, 7) {real, imag} */,
  {32'hbe50513b, 32'hbf3eefc3} /* (13, 4, 6) {real, imag} */,
  {32'h3de7b84e, 32'hc00550d2} /* (13, 4, 5) {real, imag} */,
  {32'hc00166fa, 32'h408efde1} /* (13, 4, 4) {real, imag} */,
  {32'hbe2104a1, 32'h3fb6598e} /* (13, 4, 3) {real, imag} */,
  {32'h3fb1c3c0, 32'hbded8590} /* (13, 4, 2) {real, imag} */,
  {32'h3f2d201d, 32'h3fcacd2e} /* (13, 4, 1) {real, imag} */,
  {32'h3f57d80a, 32'hc01c6833} /* (13, 4, 0) {real, imag} */,
  {32'hbf1a7842, 32'h3f097b7d} /* (13, 3, 31) {real, imag} */,
  {32'hbfa1a81d, 32'hbfa79b23} /* (13, 3, 30) {real, imag} */,
  {32'hbf0c03d6, 32'hc02efc89} /* (13, 3, 29) {real, imag} */,
  {32'h3f5c925f, 32'hbeee4fb1} /* (13, 3, 28) {real, imag} */,
  {32'hbdcd6359, 32'hbf381db6} /* (13, 3, 27) {real, imag} */,
  {32'hbe5d0b71, 32'h40316017} /* (13, 3, 26) {real, imag} */,
  {32'h3fd9c80c, 32'h3e1b9f5b} /* (13, 3, 25) {real, imag} */,
  {32'hbf36c356, 32'h3c70c214} /* (13, 3, 24) {real, imag} */,
  {32'h3eea9f93, 32'hbd94841a} /* (13, 3, 23) {real, imag} */,
  {32'h3f38a998, 32'hc016f5e4} /* (13, 3, 22) {real, imag} */,
  {32'hbe9e3a90, 32'hbe82d19d} /* (13, 3, 21) {real, imag} */,
  {32'hbfd0fd63, 32'h3f537382} /* (13, 3, 20) {real, imag} */,
  {32'hbd383792, 32'h3ffe2f27} /* (13, 3, 19) {real, imag} */,
  {32'hbe9de14b, 32'h3fcbe46f} /* (13, 3, 18) {real, imag} */,
  {32'hbf7842bd, 32'h3dfa5757} /* (13, 3, 17) {real, imag} */,
  {32'hbf79d807, 32'hbebc6559} /* (13, 3, 16) {real, imag} */,
  {32'h3f0e0ac2, 32'hbf1ec444} /* (13, 3, 15) {real, imag} */,
  {32'hc0415085, 32'hbf381f3b} /* (13, 3, 14) {real, imag} */,
  {32'h3f033ab8, 32'h400c9ee2} /* (13, 3, 13) {real, imag} */,
  {32'h3f11e9a7, 32'h3f28ed63} /* (13, 3, 12) {real, imag} */,
  {32'hbff34ae9, 32'h3eb75671} /* (13, 3, 11) {real, imag} */,
  {32'h3e802b7e, 32'h3fd75631} /* (13, 3, 10) {real, imag} */,
  {32'h3ff0ead8, 32'hbf27882d} /* (13, 3, 9) {real, imag} */,
  {32'hbf27904f, 32'h40666253} /* (13, 3, 8) {real, imag} */,
  {32'h3ecb1292, 32'h3fd99de1} /* (13, 3, 7) {real, imag} */,
  {32'hbf0792bd, 32'h3efc7d7f} /* (13, 3, 6) {real, imag} */,
  {32'hbf229048, 32'h3f997c0d} /* (13, 3, 5) {real, imag} */,
  {32'h3fdc208d, 32'h3f916241} /* (13, 3, 4) {real, imag} */,
  {32'hbf74c1cf, 32'hbe0d785c} /* (13, 3, 3) {real, imag} */,
  {32'hbfb73a16, 32'h3f16494f} /* (13, 3, 2) {real, imag} */,
  {32'hbf91de9e, 32'hbf880cc7} /* (13, 3, 1) {real, imag} */,
  {32'hbfd84f38, 32'hbc2452e7} /* (13, 3, 0) {real, imag} */,
  {32'hbf83cb0c, 32'h3f982026} /* (13, 2, 31) {real, imag} */,
  {32'h40189c0d, 32'h404bf6ac} /* (13, 2, 30) {real, imag} */,
  {32'h40654440, 32'hbf91b5bd} /* (13, 2, 29) {real, imag} */,
  {32'h40213ab3, 32'h3f731676} /* (13, 2, 28) {real, imag} */,
  {32'hc025c19d, 32'h3e4812f8} /* (13, 2, 27) {real, imag} */,
  {32'hbea50518, 32'hc05c286e} /* (13, 2, 26) {real, imag} */,
  {32'h3fd767eb, 32'hbf3ff10e} /* (13, 2, 25) {real, imag} */,
  {32'hc00d9236, 32'hc012484c} /* (13, 2, 24) {real, imag} */,
  {32'h3f887a21, 32'h40227a14} /* (13, 2, 23) {real, imag} */,
  {32'hc0174af6, 32'hbf2ed9f9} /* (13, 2, 22) {real, imag} */,
  {32'hc0224b80, 32'h3f7695e8} /* (13, 2, 21) {real, imag} */,
  {32'hbece1432, 32'h3f58010f} /* (13, 2, 20) {real, imag} */,
  {32'hbf7dc12e, 32'h3f42e472} /* (13, 2, 19) {real, imag} */,
  {32'h400245d6, 32'h3fd3a507} /* (13, 2, 18) {real, imag} */,
  {32'hbe82d4d9, 32'hbf3ee339} /* (13, 2, 17) {real, imag} */,
  {32'h3f275e41, 32'h3e1abbdf} /* (13, 2, 16) {real, imag} */,
  {32'h3fe548b6, 32'hbf9f1b56} /* (13, 2, 15) {real, imag} */,
  {32'h3f92baef, 32'h401e400c} /* (13, 2, 14) {real, imag} */,
  {32'hbe2669e4, 32'hbffd7e34} /* (13, 2, 13) {real, imag} */,
  {32'hc000e0cb, 32'hc0129e02} /* (13, 2, 12) {real, imag} */,
  {32'h3e112ffd, 32'h3fcb6f41} /* (13, 2, 11) {real, imag} */,
  {32'hbf332ffd, 32'h3e9f697f} /* (13, 2, 10) {real, imag} */,
  {32'hbfd22f14, 32'hbf441fbb} /* (13, 2, 9) {real, imag} */,
  {32'hc051c68a, 32'h4003112c} /* (13, 2, 8) {real, imag} */,
  {32'hbf7b5cac, 32'hbfd5f7cb} /* (13, 2, 7) {real, imag} */,
  {32'hc0123416, 32'hbfbfd488} /* (13, 2, 6) {real, imag} */,
  {32'hbf87ebb6, 32'hc02cfb89} /* (13, 2, 5) {real, imag} */,
  {32'h3ebfce07, 32'h4035740e} /* (13, 2, 4) {real, imag} */,
  {32'h3f834024, 32'hbeac8c61} /* (13, 2, 3) {real, imag} */,
  {32'hbf92ac44, 32'h4013ea78} /* (13, 2, 2) {real, imag} */,
  {32'h3fb7d2ab, 32'hc074c0c2} /* (13, 2, 1) {real, imag} */,
  {32'h40248d38, 32'h3f15ce9b} /* (13, 2, 0) {real, imag} */,
  {32'h402262d6, 32'h3f40a034} /* (13, 1, 31) {real, imag} */,
  {32'h3fc2ecdc, 32'h3f8d7499} /* (13, 1, 30) {real, imag} */,
  {32'h407ed389, 32'h3ed0b449} /* (13, 1, 29) {real, imag} */,
  {32'h3f459bc3, 32'hbe0ca201} /* (13, 1, 28) {real, imag} */,
  {32'hbf4e480e, 32'h401dff43} /* (13, 1, 27) {real, imag} */,
  {32'h3f641856, 32'h3e3c644f} /* (13, 1, 26) {real, imag} */,
  {32'h3f25fdee, 32'h3fbc35c2} /* (13, 1, 25) {real, imag} */,
  {32'h400a21f2, 32'h4025278e} /* (13, 1, 24) {real, imag} */,
  {32'h3f3fd089, 32'h400a1f28} /* (13, 1, 23) {real, imag} */,
  {32'h3f97d99d, 32'h3eb031ef} /* (13, 1, 22) {real, imag} */,
  {32'hbfb4f54c, 32'h3f0a6624} /* (13, 1, 21) {real, imag} */,
  {32'hc066d15e, 32'h3ee91c83} /* (13, 1, 20) {real, imag} */,
  {32'h3f8753c5, 32'h3df1dee6} /* (13, 1, 19) {real, imag} */,
  {32'h3eb2d486, 32'h3f7549cb} /* (13, 1, 18) {real, imag} */,
  {32'hbfd8a9eb, 32'hbe48fc8e} /* (13, 1, 17) {real, imag} */,
  {32'h4007f799, 32'hc05c7144} /* (13, 1, 16) {real, imag} */,
  {32'hbed44af6, 32'h3f75638a} /* (13, 1, 15) {real, imag} */,
  {32'h3e9c93a4, 32'hbfcbcb22} /* (13, 1, 14) {real, imag} */,
  {32'h3f1c7ead, 32'hbea37ae2} /* (13, 1, 13) {real, imag} */,
  {32'hbf69a8ef, 32'hbf62ade9} /* (13, 1, 12) {real, imag} */,
  {32'h4090042d, 32'hbe57b685} /* (13, 1, 11) {real, imag} */,
  {32'h3f8b99b8, 32'h3f1c411d} /* (13, 1, 10) {real, imag} */,
  {32'hbfb90cb1, 32'hc0a2682e} /* (13, 1, 9) {real, imag} */,
  {32'hbf4a644a, 32'h3e261d30} /* (13, 1, 8) {real, imag} */,
  {32'hbfd7d06a, 32'hbea6a295} /* (13, 1, 7) {real, imag} */,
  {32'h3fcf8fd5, 32'h3e9a1776} /* (13, 1, 6) {real, imag} */,
  {32'hbf68337f, 32'h3eb4016f} /* (13, 1, 5) {real, imag} */,
  {32'hbef04e4b, 32'h3fda43ac} /* (13, 1, 4) {real, imag} */,
  {32'h3f34f383, 32'hbfa6a455} /* (13, 1, 3) {real, imag} */,
  {32'hbf22766c, 32'h401bd976} /* (13, 1, 2) {real, imag} */,
  {32'hc02f143b, 32'hbe4f21ec} /* (13, 1, 1) {real, imag} */,
  {32'h3fe7ff12, 32'h3f4ef287} /* (13, 1, 0) {real, imag} */,
  {32'hbff1a0c9, 32'h3ee70613} /* (13, 0, 31) {real, imag} */,
  {32'h40023ce4, 32'h3fd673ce} /* (13, 0, 30) {real, imag} */,
  {32'h3ecdea9b, 32'hc04a69d5} /* (13, 0, 29) {real, imag} */,
  {32'h3ec7640b, 32'h4013245d} /* (13, 0, 28) {real, imag} */,
  {32'hbfb6217e, 32'hbe8caa03} /* (13, 0, 27) {real, imag} */,
  {32'hbf9868eb, 32'hbf915ec2} /* (13, 0, 26) {real, imag} */,
  {32'hbfd7437a, 32'hbe964c45} /* (13, 0, 25) {real, imag} */,
  {32'hc003ad94, 32'h401e3624} /* (13, 0, 24) {real, imag} */,
  {32'h4060cd5d, 32'hbe989d7a} /* (13, 0, 23) {real, imag} */,
  {32'hbfa1de18, 32'h40394282} /* (13, 0, 22) {real, imag} */,
  {32'h4085d3b0, 32'hbfc6840e} /* (13, 0, 21) {real, imag} */,
  {32'hbfd0895a, 32'h3ef1c6e8} /* (13, 0, 20) {real, imag} */,
  {32'hbffedce4, 32'h3f7d5a94} /* (13, 0, 19) {real, imag} */,
  {32'h3e7112b4, 32'h3f3008c5} /* (13, 0, 18) {real, imag} */,
  {32'h3fea22f4, 32'hbf1b8138} /* (13, 0, 17) {real, imag} */,
  {32'hc0101cdb, 32'h400d34d1} /* (13, 0, 16) {real, imag} */,
  {32'hbe702583, 32'hbe83d7cf} /* (13, 0, 15) {real, imag} */,
  {32'h3d26f8f6, 32'h3e0acad4} /* (13, 0, 14) {real, imag} */,
  {32'h3f0eb28f, 32'h3ee95a10} /* (13, 0, 13) {real, imag} */,
  {32'h3f130ef1, 32'hbef3fef0} /* (13, 0, 12) {real, imag} */,
  {32'h3f61efb8, 32'h3f71d034} /* (13, 0, 11) {real, imag} */,
  {32'hc0077c1f, 32'hbfaaa56f} /* (13, 0, 10) {real, imag} */,
  {32'h3d9a6281, 32'hbf86ff59} /* (13, 0, 9) {real, imag} */,
  {32'hbfb158f0, 32'h3e69df8a} /* (13, 0, 8) {real, imag} */,
  {32'hbf2e55e9, 32'h3fb0cd75} /* (13, 0, 7) {real, imag} */,
  {32'hc0160973, 32'hbfacb501} /* (13, 0, 6) {real, imag} */,
  {32'h3dc7bdbf, 32'hbf8ee409} /* (13, 0, 5) {real, imag} */,
  {32'h3f9407a7, 32'hc01e3167} /* (13, 0, 4) {real, imag} */,
  {32'h3fdce0fe, 32'hbfb5c528} /* (13, 0, 3) {real, imag} */,
  {32'hbe97d10c, 32'hbfb1fa94} /* (13, 0, 2) {real, imag} */,
  {32'h3f459184, 32'hc03aceef} /* (13, 0, 1) {real, imag} */,
  {32'hbe7ff58c, 32'hbd3ae56e} /* (13, 0, 0) {real, imag} */,
  {32'hc0353655, 32'h3f6c2883} /* (12, 31, 31) {real, imag} */,
  {32'hc047278d, 32'h3e8a880b} /* (12, 31, 30) {real, imag} */,
  {32'hbfb617dd, 32'hbf846d04} /* (12, 31, 29) {real, imag} */,
  {32'h3dd25a15, 32'hc01dddca} /* (12, 31, 28) {real, imag} */,
  {32'hbf0796c6, 32'h3f2104a0} /* (12, 31, 27) {real, imag} */,
  {32'hc0475e0b, 32'hbda474d5} /* (12, 31, 26) {real, imag} */,
  {32'h3ff28215, 32'h40608b89} /* (12, 31, 25) {real, imag} */,
  {32'hbfdda269, 32'h3f1da6f0} /* (12, 31, 24) {real, imag} */,
  {32'hbee9764b, 32'h3f28ee77} /* (12, 31, 23) {real, imag} */,
  {32'hc00c2906, 32'hbf6995d6} /* (12, 31, 22) {real, imag} */,
  {32'h40602b63, 32'hbf724f7e} /* (12, 31, 21) {real, imag} */,
  {32'h3e295be1, 32'hbeec99ab} /* (12, 31, 20) {real, imag} */,
  {32'h3eeb5468, 32'h3ffaadee} /* (12, 31, 19) {real, imag} */,
  {32'h401bda2d, 32'h3f541e5c} /* (12, 31, 18) {real, imag} */,
  {32'hbf6cbdac, 32'h3ec5a969} /* (12, 31, 17) {real, imag} */,
  {32'hbb65d508, 32'hbf83f9c5} /* (12, 31, 16) {real, imag} */,
  {32'hc016d070, 32'h40024d60} /* (12, 31, 15) {real, imag} */,
  {32'h3d12c71d, 32'h3d8cb836} /* (12, 31, 14) {real, imag} */,
  {32'h3fe647d7, 32'h40536300} /* (12, 31, 13) {real, imag} */,
  {32'h3f325091, 32'hbf06b9ea} /* (12, 31, 12) {real, imag} */,
  {32'hbfaf7141, 32'h408d86cf} /* (12, 31, 11) {real, imag} */,
  {32'h402fe66c, 32'hbf0babba} /* (12, 31, 10) {real, imag} */,
  {32'h4030353e, 32'h3e429bb6} /* (12, 31, 9) {real, imag} */,
  {32'h3fd00779, 32'h3eee4179} /* (12, 31, 8) {real, imag} */,
  {32'hbf613532, 32'h3f473900} /* (12, 31, 7) {real, imag} */,
  {32'h3f4f2ae7, 32'h3fd11fd7} /* (12, 31, 6) {real, imag} */,
  {32'h400d385f, 32'hbfbb7db6} /* (12, 31, 5) {real, imag} */,
  {32'hbfa003cf, 32'hbe85d632} /* (12, 31, 4) {real, imag} */,
  {32'h3fa398ab, 32'h3f110027} /* (12, 31, 3) {real, imag} */,
  {32'hbe1389bb, 32'h3f434144} /* (12, 31, 2) {real, imag} */,
  {32'hbfb7e887, 32'hbebda4ea} /* (12, 31, 1) {real, imag} */,
  {32'h3fd3f4f3, 32'h3fb0827a} /* (12, 31, 0) {real, imag} */,
  {32'hbf5a4b5f, 32'hbef661fc} /* (12, 30, 31) {real, imag} */,
  {32'hc01323ab, 32'h3f4a1eb7} /* (12, 30, 30) {real, imag} */,
  {32'h3fd7b40f, 32'h3faf0664} /* (12, 30, 29) {real, imag} */,
  {32'h3eb73e12, 32'hbf42c140} /* (12, 30, 28) {real, imag} */,
  {32'h3fc443dd, 32'hbf70d5df} /* (12, 30, 27) {real, imag} */,
  {32'h3f7c7eeb, 32'hbe22ae1c} /* (12, 30, 26) {real, imag} */,
  {32'h3fe4549b, 32'h4014a118} /* (12, 30, 25) {real, imag} */,
  {32'h3fa39cd9, 32'h3ed54fe1} /* (12, 30, 24) {real, imag} */,
  {32'h3fe0d7fe, 32'h3ee4fd5a} /* (12, 30, 23) {real, imag} */,
  {32'hbf062f74, 32'h3e63489f} /* (12, 30, 22) {real, imag} */,
  {32'hc0054e60, 32'h3ed60041} /* (12, 30, 21) {real, imag} */,
  {32'h4058abb9, 32'h4018998c} /* (12, 30, 20) {real, imag} */,
  {32'hbf4822bf, 32'hbefdb01f} /* (12, 30, 19) {real, imag} */,
  {32'hbfef57c9, 32'h3f8144ab} /* (12, 30, 18) {real, imag} */,
  {32'hbf852081, 32'h3eb23713} /* (12, 30, 17) {real, imag} */,
  {32'hbf7590ba, 32'hbf9e4966} /* (12, 30, 16) {real, imag} */,
  {32'h3f8619d6, 32'hbfa17f75} /* (12, 30, 15) {real, imag} */,
  {32'h3fc2849b, 32'hbfaae9f2} /* (12, 30, 14) {real, imag} */,
  {32'hbf6ff8ce, 32'h3e5ada41} /* (12, 30, 13) {real, imag} */,
  {32'h3f21f1a8, 32'hbe3e4814} /* (12, 30, 12) {real, imag} */,
  {32'hbdec559b, 32'h3f8b4a9f} /* (12, 30, 11) {real, imag} */,
  {32'hbdaf0a77, 32'h3ec9862f} /* (12, 30, 10) {real, imag} */,
  {32'hbf32a676, 32'h3fab55cd} /* (12, 30, 9) {real, imag} */,
  {32'hbebfd46c, 32'hbe1c3ae9} /* (12, 30, 8) {real, imag} */,
  {32'h4084d19e, 32'hbf5df565} /* (12, 30, 7) {real, imag} */,
  {32'h3fb94a0b, 32'h3f75cf09} /* (12, 30, 6) {real, imag} */,
  {32'h3fb54a8e, 32'hbf800d31} /* (12, 30, 5) {real, imag} */,
  {32'h3d70608b, 32'hc01003d9} /* (12, 30, 4) {real, imag} */,
  {32'h40432d51, 32'hc0052cc1} /* (12, 30, 3) {real, imag} */,
  {32'hbf748537, 32'h3dc3fb60} /* (12, 30, 2) {real, imag} */,
  {32'h3fdc1830, 32'h40a31230} /* (12, 30, 1) {real, imag} */,
  {32'h3f0907e4, 32'hbfcb7206} /* (12, 30, 0) {real, imag} */,
  {32'h3ef3b9c0, 32'h40a34614} /* (12, 29, 31) {real, imag} */,
  {32'h4005eaf3, 32'hbf4da739} /* (12, 29, 30) {real, imag} */,
  {32'h3ffe5b77, 32'hc00c60db} /* (12, 29, 29) {real, imag} */,
  {32'h3fe60eac, 32'hbfc606c1} /* (12, 29, 28) {real, imag} */,
  {32'h3e8b88d1, 32'h3f2251c8} /* (12, 29, 27) {real, imag} */,
  {32'hbe24f9a9, 32'h3e0fff0d} /* (12, 29, 26) {real, imag} */,
  {32'hbe7cabf5, 32'hbf99d7b7} /* (12, 29, 25) {real, imag} */,
  {32'h40063d5c, 32'h3fbec654} /* (12, 29, 24) {real, imag} */,
  {32'h3fc0b84c, 32'hbf9b510e} /* (12, 29, 23) {real, imag} */,
  {32'hbecaa01b, 32'h405fdafd} /* (12, 29, 22) {real, imag} */,
  {32'hbee0aa15, 32'h3e5ecaca} /* (12, 29, 21) {real, imag} */,
  {32'hbf2128fe, 32'hc0237b9b} /* (12, 29, 20) {real, imag} */,
  {32'hc0386609, 32'h3f8be949} /* (12, 29, 19) {real, imag} */,
  {32'h3ed6ee6f, 32'h3e8de53e} /* (12, 29, 18) {real, imag} */,
  {32'hc00e9726, 32'h40202454} /* (12, 29, 17) {real, imag} */,
  {32'h3ea72d25, 32'h3f17c891} /* (12, 29, 16) {real, imag} */,
  {32'hbdf17ff5, 32'hbf153b8a} /* (12, 29, 15) {real, imag} */,
  {32'hbf58b9a7, 32'hbfda278c} /* (12, 29, 14) {real, imag} */,
  {32'hbf47c8f3, 32'hbf75001f} /* (12, 29, 13) {real, imag} */,
  {32'h3fd54999, 32'hbf1ecb03} /* (12, 29, 12) {real, imag} */,
  {32'h3adb17d8, 32'hbf40f567} /* (12, 29, 11) {real, imag} */,
  {32'hc0309cc5, 32'h3fa4ec57} /* (12, 29, 10) {real, imag} */,
  {32'hbee8be94, 32'h3d3ce824} /* (12, 29, 9) {real, imag} */,
  {32'hbfda5028, 32'hbed1a5d8} /* (12, 29, 8) {real, imag} */,
  {32'h3f945b3c, 32'hc05ab407} /* (12, 29, 7) {real, imag} */,
  {32'h3e8c103a, 32'hbfc6d3da} /* (12, 29, 6) {real, imag} */,
  {32'hbf97b651, 32'hbea891ad} /* (12, 29, 5) {real, imag} */,
  {32'h3fd24078, 32'h402db80c} /* (12, 29, 4) {real, imag} */,
  {32'hbf35df50, 32'hc099ecdc} /* (12, 29, 3) {real, imag} */,
  {32'h3f926d01, 32'h3f468f35} /* (12, 29, 2) {real, imag} */,
  {32'h3f3a4129, 32'hc030a671} /* (12, 29, 1) {real, imag} */,
  {32'h3eed901c, 32'hbe7dfc2e} /* (12, 29, 0) {real, imag} */,
  {32'hbf200783, 32'h3f6ad6d3} /* (12, 28, 31) {real, imag} */,
  {32'hc0008d7d, 32'h3f8f8212} /* (12, 28, 30) {real, imag} */,
  {32'hbf034a98, 32'hbffe966c} /* (12, 28, 29) {real, imag} */,
  {32'h3ede4271, 32'h3f967aff} /* (12, 28, 28) {real, imag} */,
  {32'hc016ef47, 32'hbe7c64f9} /* (12, 28, 27) {real, imag} */,
  {32'hbdfab129, 32'h3f6f6817} /* (12, 28, 26) {real, imag} */,
  {32'h3ee1d115, 32'hc0000a1b} /* (12, 28, 25) {real, imag} */,
  {32'hbfbf8a65, 32'hbf6ccd61} /* (12, 28, 24) {real, imag} */,
  {32'h3ef01ccf, 32'hc059acc6} /* (12, 28, 23) {real, imag} */,
  {32'hc06cd84e, 32'h3ff78efc} /* (12, 28, 22) {real, imag} */,
  {32'hbe93e3f6, 32'h3f4b3618} /* (12, 28, 21) {real, imag} */,
  {32'h3fa49e7a, 32'hbe522390} /* (12, 28, 20) {real, imag} */,
  {32'hbfd69bc0, 32'h3fc8c46d} /* (12, 28, 19) {real, imag} */,
  {32'h3fa40293, 32'h3e9ad510} /* (12, 28, 18) {real, imag} */,
  {32'h3f67a946, 32'h3f2b57f6} /* (12, 28, 17) {real, imag} */,
  {32'hbec1b1cb, 32'hbef51fca} /* (12, 28, 16) {real, imag} */,
  {32'h3f574873, 32'h3faaabe1} /* (12, 28, 15) {real, imag} */,
  {32'h3f1f0c2c, 32'hc0306c07} /* (12, 28, 14) {real, imag} */,
  {32'h3f2c3640, 32'h3e2ed077} /* (12, 28, 13) {real, imag} */,
  {32'hbfbf9734, 32'hbf12524b} /* (12, 28, 12) {real, imag} */,
  {32'hc066fa13, 32'h3f712fe4} /* (12, 28, 11) {real, imag} */,
  {32'h3fbfb096, 32'h3fed7e91} /* (12, 28, 10) {real, imag} */,
  {32'h40104a83, 32'h3f8863ec} /* (12, 28, 9) {real, imag} */,
  {32'hc023f797, 32'h4024cfea} /* (12, 28, 8) {real, imag} */,
  {32'h3f1eb2dd, 32'hbe9880d0} /* (12, 28, 7) {real, imag} */,
  {32'h4015ed4f, 32'hbf95b10c} /* (12, 28, 6) {real, imag} */,
  {32'h3cd26528, 32'hc05c09a1} /* (12, 28, 5) {real, imag} */,
  {32'hbf5765d8, 32'h3eea82cb} /* (12, 28, 4) {real, imag} */,
  {32'hc01bcc4a, 32'hbe52d956} /* (12, 28, 3) {real, imag} */,
  {32'h3fc0fdfe, 32'h3fa65a87} /* (12, 28, 2) {real, imag} */,
  {32'h3f69dc05, 32'h3eab84dd} /* (12, 28, 1) {real, imag} */,
  {32'h3f1f386a, 32'h40008e0b} /* (12, 28, 0) {real, imag} */,
  {32'h3f93b6cf, 32'hc00f80a2} /* (12, 27, 31) {real, imag} */,
  {32'hbfbeab12, 32'h3ba6dcf5} /* (12, 27, 30) {real, imag} */,
  {32'hbf81a7b6, 32'h3eeed2a6} /* (12, 27, 29) {real, imag} */,
  {32'hbf01f52e, 32'hc01149bf} /* (12, 27, 28) {real, imag} */,
  {32'hbfe2c7af, 32'hc01e6a55} /* (12, 27, 27) {real, imag} */,
  {32'hbfe9aff0, 32'hbfade756} /* (12, 27, 26) {real, imag} */,
  {32'h400f9332, 32'h3fffac1e} /* (12, 27, 25) {real, imag} */,
  {32'hbe2966ec, 32'h4057ac12} /* (12, 27, 24) {real, imag} */,
  {32'hc006e7ce, 32'hbfc88063} /* (12, 27, 23) {real, imag} */,
  {32'hbfb8f875, 32'h3effda43} /* (12, 27, 22) {real, imag} */,
  {32'h40154bfe, 32'hbf03113c} /* (12, 27, 21) {real, imag} */,
  {32'hbe197aa5, 32'h3f829bd8} /* (12, 27, 20) {real, imag} */,
  {32'h3e5df4a1, 32'hbfb1194c} /* (12, 27, 19) {real, imag} */,
  {32'h3e06f591, 32'hbf52e916} /* (12, 27, 18) {real, imag} */,
  {32'hbe65ee37, 32'hbfc20f72} /* (12, 27, 17) {real, imag} */,
  {32'hbfdd5939, 32'hbeacf1d8} /* (12, 27, 16) {real, imag} */,
  {32'h3f34d7bc, 32'hbde3fee8} /* (12, 27, 15) {real, imag} */,
  {32'hbfb33a99, 32'hbf1b57d3} /* (12, 27, 14) {real, imag} */,
  {32'h3f3b69fd, 32'h3f3d08b9} /* (12, 27, 13) {real, imag} */,
  {32'hbeb81324, 32'hc0054147} /* (12, 27, 12) {real, imag} */,
  {32'hc004d13c, 32'h4073f2b1} /* (12, 27, 11) {real, imag} */,
  {32'hbf6c48d1, 32'h3ebaf89f} /* (12, 27, 10) {real, imag} */,
  {32'h40077c28, 32'hc0533c57} /* (12, 27, 9) {real, imag} */,
  {32'hc056dcea, 32'h3f790597} /* (12, 27, 8) {real, imag} */,
  {32'hbf634473, 32'hbee745a0} /* (12, 27, 7) {real, imag} */,
  {32'hbf14720f, 32'hc0344ea8} /* (12, 27, 6) {real, imag} */,
  {32'h3f5f9e9f, 32'hbfd03172} /* (12, 27, 5) {real, imag} */,
  {32'hbf80f8b2, 32'hbe3998f5} /* (12, 27, 4) {real, imag} */,
  {32'hc033ce62, 32'h3fdf6244} /* (12, 27, 3) {real, imag} */,
  {32'h3e063e45, 32'h3f1031cf} /* (12, 27, 2) {real, imag} */,
  {32'h3f918d6d, 32'h3d5e6d0d} /* (12, 27, 1) {real, imag} */,
  {32'h3f9e5285, 32'hbf2a5b82} /* (12, 27, 0) {real, imag} */,
  {32'hbfac2b45, 32'h402f1c1f} /* (12, 26, 31) {real, imag} */,
  {32'h3f9d136c, 32'h3d28bd1f} /* (12, 26, 30) {real, imag} */,
  {32'h40329c15, 32'h3f910e56} /* (12, 26, 29) {real, imag} */,
  {32'hbf2ca3dc, 32'hc073154d} /* (12, 26, 28) {real, imag} */,
  {32'h3e778a0c, 32'h3f878b64} /* (12, 26, 27) {real, imag} */,
  {32'h3e3b2f4a, 32'hbf989242} /* (12, 26, 26) {real, imag} */,
  {32'h405ab3bf, 32'hbdbbf1a9} /* (12, 26, 25) {real, imag} */,
  {32'hbfe39220, 32'h3f92be5c} /* (12, 26, 24) {real, imag} */,
  {32'hbfe11ebe, 32'h3f9803f9} /* (12, 26, 23) {real, imag} */,
  {32'h3f1a7cc2, 32'hbed3e339} /* (12, 26, 22) {real, imag} */,
  {32'hbf61b187, 32'hbe823514} /* (12, 26, 21) {real, imag} */,
  {32'h3fe41644, 32'h3f9b9bad} /* (12, 26, 20) {real, imag} */,
  {32'h3f52a280, 32'hbf65b811} /* (12, 26, 19) {real, imag} */,
  {32'h3fefdd36, 32'h3d8c7160} /* (12, 26, 18) {real, imag} */,
  {32'hbfbe24e8, 32'h3fd1966a} /* (12, 26, 17) {real, imag} */,
  {32'hbd8b7b59, 32'hbf59cc7b} /* (12, 26, 16) {real, imag} */,
  {32'h3fc33686, 32'hbf78fa83} /* (12, 26, 15) {real, imag} */,
  {32'h3ee4fefb, 32'h4012ec89} /* (12, 26, 14) {real, imag} */,
  {32'h4032dacb, 32'hbe1545dd} /* (12, 26, 13) {real, imag} */,
  {32'hbf7053ca, 32'h4024ce4c} /* (12, 26, 12) {real, imag} */,
  {32'hbf3c901a, 32'hbfa7f6aa} /* (12, 26, 11) {real, imag} */,
  {32'h3ee79523, 32'hbfff9486} /* (12, 26, 10) {real, imag} */,
  {32'hbfa5eee3, 32'h3f887ab3} /* (12, 26, 9) {real, imag} */,
  {32'h4031dd4c, 32'h3f8b70fb} /* (12, 26, 8) {real, imag} */,
  {32'h3f4ff034, 32'hbf57148b} /* (12, 26, 7) {real, imag} */,
  {32'hc084394e, 32'hbf56be4d} /* (12, 26, 6) {real, imag} */,
  {32'h401d5eef, 32'hbf318257} /* (12, 26, 5) {real, imag} */,
  {32'h3fc8ce81, 32'hbefa17f0} /* (12, 26, 4) {real, imag} */,
  {32'h3f8e87d6, 32'h4020817b} /* (12, 26, 3) {real, imag} */,
  {32'hc0756c00, 32'h3f947e50} /* (12, 26, 2) {real, imag} */,
  {32'hbfaa0cbb, 32'hbf08cde2} /* (12, 26, 1) {real, imag} */,
  {32'hbec6219a, 32'h3e959412} /* (12, 26, 0) {real, imag} */,
  {32'h3fa32e66, 32'h3fdbdaf3} /* (12, 25, 31) {real, imag} */,
  {32'h402476d2, 32'h3f092fe3} /* (12, 25, 30) {real, imag} */,
  {32'hbeca7ea4, 32'h3f4d4516} /* (12, 25, 29) {real, imag} */,
  {32'hbf97acf1, 32'h3f8a011c} /* (12, 25, 28) {real, imag} */,
  {32'hc023a366, 32'h3fded2a8} /* (12, 25, 27) {real, imag} */,
  {32'h40278247, 32'h3fd119a7} /* (12, 25, 26) {real, imag} */,
  {32'h3f1c3181, 32'h3f2695f8} /* (12, 25, 25) {real, imag} */,
  {32'hbfe21c87, 32'hc071f08b} /* (12, 25, 24) {real, imag} */,
  {32'h401e0b23, 32'hbfb27d6e} /* (12, 25, 23) {real, imag} */,
  {32'hbfec8db3, 32'hc006af4b} /* (12, 25, 22) {real, imag} */,
  {32'h3ec433b9, 32'hbf175f86} /* (12, 25, 21) {real, imag} */,
  {32'hbfac9207, 32'h3f37ee51} /* (12, 25, 20) {real, imag} */,
  {32'hbe91cade, 32'hc0250f97} /* (12, 25, 19) {real, imag} */,
  {32'h401d5de9, 32'hbf7fd037} /* (12, 25, 18) {real, imag} */,
  {32'hbf8dfd73, 32'hbfabaae1} /* (12, 25, 17) {real, imag} */,
  {32'hc017cc6c, 32'hbdf61074} /* (12, 25, 16) {real, imag} */,
  {32'hbfb15f30, 32'h3ed60e27} /* (12, 25, 15) {real, imag} */,
  {32'h400e8f0b, 32'hbe73b03b} /* (12, 25, 14) {real, imag} */,
  {32'hbeb0f837, 32'h3e4e6461} /* (12, 25, 13) {real, imag} */,
  {32'h3ef015f5, 32'h3f1c3a04} /* (12, 25, 12) {real, imag} */,
  {32'h3e8010d2, 32'hbfc7c573} /* (12, 25, 11) {real, imag} */,
  {32'h3fd4fc8a, 32'hbff71eb0} /* (12, 25, 10) {real, imag} */,
  {32'hbfddafae, 32'hbf72d25e} /* (12, 25, 9) {real, imag} */,
  {32'h3f0b2098, 32'hbf41343c} /* (12, 25, 8) {real, imag} */,
  {32'h3f8b47be, 32'hbfdfacb5} /* (12, 25, 7) {real, imag} */,
  {32'h3fea54c7, 32'h406e6f20} /* (12, 25, 6) {real, imag} */,
  {32'h3d8ac1c2, 32'hbf838d28} /* (12, 25, 5) {real, imag} */,
  {32'hbe756771, 32'h3f9c6da0} /* (12, 25, 4) {real, imag} */,
  {32'hc0006f24, 32'hc06ff3e6} /* (12, 25, 3) {real, imag} */,
  {32'hbf2427b1, 32'h3e85bc84} /* (12, 25, 2) {real, imag} */,
  {32'h3f0a9506, 32'hc03da33f} /* (12, 25, 1) {real, imag} */,
  {32'hbfd58b62, 32'h3fb5f782} /* (12, 25, 0) {real, imag} */,
  {32'h3f1b54f4, 32'hbf804f9b} /* (12, 24, 31) {real, imag} */,
  {32'hbf8dd066, 32'h3f42f672} /* (12, 24, 30) {real, imag} */,
  {32'h3f8e558e, 32'h40871654} /* (12, 24, 29) {real, imag} */,
  {32'hc002eac2, 32'h3fcdac38} /* (12, 24, 28) {real, imag} */,
  {32'hbf3c0d97, 32'hc06f8b0c} /* (12, 24, 27) {real, imag} */,
  {32'h3f7741c3, 32'h4073b581} /* (12, 24, 26) {real, imag} */,
  {32'hc0536a38, 32'hbe1607db} /* (12, 24, 25) {real, imag} */,
  {32'hbb6b258f, 32'h402333b4} /* (12, 24, 24) {real, imag} */,
  {32'hbcb75507, 32'h3fab7943} /* (12, 24, 23) {real, imag} */,
  {32'hc09071da, 32'h4064fafa} /* (12, 24, 22) {real, imag} */,
  {32'hbf2c155d, 32'hbff6a43c} /* (12, 24, 21) {real, imag} */,
  {32'h40557013, 32'h4081590c} /* (12, 24, 20) {real, imag} */,
  {32'h40962234, 32'h3f08ec1b} /* (12, 24, 19) {real, imag} */,
  {32'hc0181875, 32'hc018b43e} /* (12, 24, 18) {real, imag} */,
  {32'h3f1bfc9a, 32'h3f42b4fe} /* (12, 24, 17) {real, imag} */,
  {32'h3f3c0c17, 32'hbf329603} /* (12, 24, 16) {real, imag} */,
  {32'hbf004c7f, 32'hbed08236} /* (12, 24, 15) {real, imag} */,
  {32'h3e4cb5ae, 32'h3fc9c3e3} /* (12, 24, 14) {real, imag} */,
  {32'h3ee6965f, 32'h3e9671e5} /* (12, 24, 13) {real, imag} */,
  {32'h3e66aeef, 32'h3f959640} /* (12, 24, 12) {real, imag} */,
  {32'h3f4d703f, 32'hc031fcbb} /* (12, 24, 11) {real, imag} */,
  {32'h3eee08ff, 32'h40359582} /* (12, 24, 10) {real, imag} */,
  {32'h3fac76a8, 32'hbfbc7409} /* (12, 24, 9) {real, imag} */,
  {32'hbf0b017d, 32'h405c489e} /* (12, 24, 8) {real, imag} */,
  {32'hbf759b33, 32'hbf87ee7e} /* (12, 24, 7) {real, imag} */,
  {32'h3dc46363, 32'hbebf2758} /* (12, 24, 6) {real, imag} */,
  {32'h3f1a445b, 32'h3f47c0d9} /* (12, 24, 5) {real, imag} */,
  {32'h3fbf35cf, 32'h3f4392da} /* (12, 24, 4) {real, imag} */,
  {32'hc0201642, 32'hbe98109a} /* (12, 24, 3) {real, imag} */,
  {32'hbfb5873d, 32'h3fd1831b} /* (12, 24, 2) {real, imag} */,
  {32'hbf8e8727, 32'h3e1b72bd} /* (12, 24, 1) {real, imag} */,
  {32'h406ebcf4, 32'h3e25a5e2} /* (12, 24, 0) {real, imag} */,
  {32'hbf12e421, 32'hc080a40b} /* (12, 23, 31) {real, imag} */,
  {32'hbf7bc307, 32'hbd9a20ae} /* (12, 23, 30) {real, imag} */,
  {32'h3fa79f4b, 32'h3fe1e93a} /* (12, 23, 29) {real, imag} */,
  {32'hc00fc45b, 32'hbfa5729d} /* (12, 23, 28) {real, imag} */,
  {32'h4075b5ab, 32'hbfc2accf} /* (12, 23, 27) {real, imag} */,
  {32'h3e839b7b, 32'h4041fb1d} /* (12, 23, 26) {real, imag} */,
  {32'h3f1bbde3, 32'h3f352d3e} /* (12, 23, 25) {real, imag} */,
  {32'hbff2e9b5, 32'hbfc4ae6b} /* (12, 23, 24) {real, imag} */,
  {32'hbfdfd3cf, 32'hbf9bc7b6} /* (12, 23, 23) {real, imag} */,
  {32'hbf8111a1, 32'hbfc83b35} /* (12, 23, 22) {real, imag} */,
  {32'h400b6520, 32'hbf8dff7b} /* (12, 23, 21) {real, imag} */,
  {32'h4067ea49, 32'hbfce8079} /* (12, 23, 20) {real, imag} */,
  {32'hbeea3c64, 32'h40824a3c} /* (12, 23, 19) {real, imag} */,
  {32'h3f8ca945, 32'hc0408828} /* (12, 23, 18) {real, imag} */,
  {32'hbf031162, 32'hbfb53561} /* (12, 23, 17) {real, imag} */,
  {32'h3e6c1117, 32'h3fbef189} /* (12, 23, 16) {real, imag} */,
  {32'hbf21fc06, 32'hbeac4071} /* (12, 23, 15) {real, imag} */,
  {32'h3f2085de, 32'hbfeb3b71} /* (12, 23, 14) {real, imag} */,
  {32'h4037df22, 32'h4011a829} /* (12, 23, 13) {real, imag} */,
  {32'hbf490462, 32'hc07f7605} /* (12, 23, 12) {real, imag} */,
  {32'hbf2779bb, 32'hbf8490eb} /* (12, 23, 11) {real, imag} */,
  {32'h3ed11ffa, 32'h3c3d4c60} /* (12, 23, 10) {real, imag} */,
  {32'h3f280a6b, 32'hbf77728c} /* (12, 23, 9) {real, imag} */,
  {32'hbe1ff9b9, 32'h3f079d47} /* (12, 23, 8) {real, imag} */,
  {32'h3fae62f5, 32'hbf25ea80} /* (12, 23, 7) {real, imag} */,
  {32'hbf15812e, 32'h400bbd13} /* (12, 23, 6) {real, imag} */,
  {32'hbd9007c4, 32'h401f188c} /* (12, 23, 5) {real, imag} */,
  {32'hbf6e051b, 32'h4014a646} /* (12, 23, 4) {real, imag} */,
  {32'hbe757597, 32'h3ea71633} /* (12, 23, 3) {real, imag} */,
  {32'h3fcfff49, 32'hbf707ef2} /* (12, 23, 2) {real, imag} */,
  {32'hbffc706a, 32'h3f29ba2e} /* (12, 23, 1) {real, imag} */,
  {32'hc002456d, 32'h4001a142} /* (12, 23, 0) {real, imag} */,
  {32'hc02d40f7, 32'h3de06018} /* (12, 22, 31) {real, imag} */,
  {32'h401dc9b2, 32'hbca9325e} /* (12, 22, 30) {real, imag} */,
  {32'hc0a8f58e, 32'hbf27790f} /* (12, 22, 29) {real, imag} */,
  {32'h3fcf89fe, 32'hbf9de663} /* (12, 22, 28) {real, imag} */,
  {32'h3f601b2f, 32'hc05cfd22} /* (12, 22, 27) {real, imag} */,
  {32'hbe395746, 32'h3f896ce0} /* (12, 22, 26) {real, imag} */,
  {32'h400a20dd, 32'h4012d7b1} /* (12, 22, 25) {real, imag} */,
  {32'h3fd42b4c, 32'hbfa5469c} /* (12, 22, 24) {real, imag} */,
  {32'hbc1a73fe, 32'hbf10ce72} /* (12, 22, 23) {real, imag} */,
  {32'h40246315, 32'h4068c343} /* (12, 22, 22) {real, imag} */,
  {32'h3ff9fd79, 32'hbd565956} /* (12, 22, 21) {real, imag} */,
  {32'h3f042e83, 32'h3f0e1aaf} /* (12, 22, 20) {real, imag} */,
  {32'hbec58dbe, 32'hbf22b557} /* (12, 22, 19) {real, imag} */,
  {32'hc0042e7e, 32'h3f604428} /* (12, 22, 18) {real, imag} */,
  {32'hbf19d1e3, 32'hbe1972fc} /* (12, 22, 17) {real, imag} */,
  {32'h3ff5a745, 32'h406101d0} /* (12, 22, 16) {real, imag} */,
  {32'h3fa3808d, 32'hbffa907d} /* (12, 22, 15) {real, imag} */,
  {32'h3e430285, 32'h3f8cc265} /* (12, 22, 14) {real, imag} */,
  {32'hbf4304b2, 32'h3ed97482} /* (12, 22, 13) {real, imag} */,
  {32'hc0240904, 32'hbf66da9d} /* (12, 22, 12) {real, imag} */,
  {32'hbfbbe448, 32'h400d613e} /* (12, 22, 11) {real, imag} */,
  {32'hbfc56a2f, 32'h3f3396de} /* (12, 22, 10) {real, imag} */,
  {32'h3f456b61, 32'h3dee141e} /* (12, 22, 9) {real, imag} */,
  {32'hc00728ff, 32'hbebf3568} /* (12, 22, 8) {real, imag} */,
  {32'hbf896959, 32'hbfa5ba82} /* (12, 22, 7) {real, imag} */,
  {32'h3fd35737, 32'hc05b7784} /* (12, 22, 6) {real, imag} */,
  {32'h3fe6b7ab, 32'h3f111498} /* (12, 22, 5) {real, imag} */,
  {32'hbe10e74c, 32'hbfdaed98} /* (12, 22, 4) {real, imag} */,
  {32'h40474c6c, 32'hbfa57442} /* (12, 22, 3) {real, imag} */,
  {32'h40317ff4, 32'h3e3c16b3} /* (12, 22, 2) {real, imag} */,
  {32'hbeafe728, 32'h40518868} /* (12, 22, 1) {real, imag} */,
  {32'hbe402dbb, 32'h402677c2} /* (12, 22, 0) {real, imag} */,
  {32'h3f1a279d, 32'h3fa536c2} /* (12, 21, 31) {real, imag} */,
  {32'h3fa2b3fa, 32'hbef87f0b} /* (12, 21, 30) {real, imag} */,
  {32'hbf9f638d, 32'hbfc09dfa} /* (12, 21, 29) {real, imag} */,
  {32'h3fe95e1c, 32'hbf0df359} /* (12, 21, 28) {real, imag} */,
  {32'hc0192ce6, 32'h3fa13f2d} /* (12, 21, 27) {real, imag} */,
  {32'hbe0801d2, 32'hbf0ddcf6} /* (12, 21, 26) {real, imag} */,
  {32'hc03c3087, 32'hbf50c036} /* (12, 21, 25) {real, imag} */,
  {32'h400ff4dc, 32'h3fbef08c} /* (12, 21, 24) {real, imag} */,
  {32'h402c37e0, 32'h4015b7d2} /* (12, 21, 23) {real, imag} */,
  {32'hbdd6d806, 32'h3fe41515} /* (12, 21, 22) {real, imag} */,
  {32'h400c89d4, 32'h4070fbd3} /* (12, 21, 21) {real, imag} */,
  {32'hc02e0748, 32'hc01d143f} /* (12, 21, 20) {real, imag} */,
  {32'hc03a52ab, 32'hc04851ce} /* (12, 21, 19) {real, imag} */,
  {32'h3e5012f7, 32'hc001c318} /* (12, 21, 18) {real, imag} */,
  {32'hbfc2ac5f, 32'hbd677150} /* (12, 21, 17) {real, imag} */,
  {32'h3d539b9c, 32'hbf161b55} /* (12, 21, 16) {real, imag} */,
  {32'h3f0e5e18, 32'h3f5ff3c3} /* (12, 21, 15) {real, imag} */,
  {32'hbdcffaf0, 32'h3f8bb87a} /* (12, 21, 14) {real, imag} */,
  {32'h3fcf0d43, 32'h3f553332} /* (12, 21, 13) {real, imag} */,
  {32'h3fc5bcdb, 32'hbfc745ba} /* (12, 21, 12) {real, imag} */,
  {32'hbfd7059a, 32'hbf304f91} /* (12, 21, 11) {real, imag} */,
  {32'hc040b3fb, 32'h4079b743} /* (12, 21, 10) {real, imag} */,
  {32'h3f90abcf, 32'hbfd914e9} /* (12, 21, 9) {real, imag} */,
  {32'hbfe75fdd, 32'h3eee877c} /* (12, 21, 8) {real, imag} */,
  {32'h4045b4e8, 32'hbfe5f36b} /* (12, 21, 7) {real, imag} */,
  {32'hc017fbdd, 32'h3fc055f7} /* (12, 21, 6) {real, imag} */,
  {32'h4033f85c, 32'hbfa83b92} /* (12, 21, 5) {real, imag} */,
  {32'h3f80b937, 32'hc0589461} /* (12, 21, 4) {real, imag} */,
  {32'hbcb44756, 32'h3ff59807} /* (12, 21, 3) {real, imag} */,
  {32'h3fd3816e, 32'hc0132395} /* (12, 21, 2) {real, imag} */,
  {32'h3fa85bcb, 32'h3fc7a285} /* (12, 21, 1) {real, imag} */,
  {32'h3ee6b147, 32'hbf0fdb89} /* (12, 21, 0) {real, imag} */,
  {32'h3fbd0add, 32'hbfa5a5aa} /* (12, 20, 31) {real, imag} */,
  {32'hbf162136, 32'hc0908909} /* (12, 20, 30) {real, imag} */,
  {32'h3fcb420b, 32'hc0048403} /* (12, 20, 29) {real, imag} */,
  {32'hbfd8071a, 32'h3e045b21} /* (12, 20, 28) {real, imag} */,
  {32'h3fcddf16, 32'h3f1b6258} /* (12, 20, 27) {real, imag} */,
  {32'h3fc89cf1, 32'hbec18edf} /* (12, 20, 26) {real, imag} */,
  {32'hbecba4a3, 32'hbfcb954a} /* (12, 20, 25) {real, imag} */,
  {32'hc08107bc, 32'h3e1adae1} /* (12, 20, 24) {real, imag} */,
  {32'h3fcc84b5, 32'h3f813d2a} /* (12, 20, 23) {real, imag} */,
  {32'h3e620893, 32'hbec95777} /* (12, 20, 22) {real, imag} */,
  {32'hc042d8b7, 32'h3fb44acb} /* (12, 20, 21) {real, imag} */,
  {32'h404e570b, 32'h3fa46307} /* (12, 20, 20) {real, imag} */,
  {32'h3fe079d6, 32'h3f7a8fc4} /* (12, 20, 19) {real, imag} */,
  {32'hbfe791f2, 32'h3fe64d6e} /* (12, 20, 18) {real, imag} */,
  {32'h3fb2ca3e, 32'h4004b91c} /* (12, 20, 17) {real, imag} */,
  {32'hbf45ec5e, 32'h3ec178e2} /* (12, 20, 16) {real, imag} */,
  {32'hbfa7af62, 32'hbf329bab} /* (12, 20, 15) {real, imag} */,
  {32'h3dbb61f5, 32'h3fd58787} /* (12, 20, 14) {real, imag} */,
  {32'h40000c0e, 32'h3f060037} /* (12, 20, 13) {real, imag} */,
  {32'h3f31460a, 32'h409e2580} /* (12, 20, 12) {real, imag} */,
  {32'h402456f2, 32'h3dc683b1} /* (12, 20, 11) {real, imag} */,
  {32'hbfbf6323, 32'hc0d92c77} /* (12, 20, 10) {real, imag} */,
  {32'hc02d4b37, 32'hbeb49ea0} /* (12, 20, 9) {real, imag} */,
  {32'hbf91079a, 32'hc02a2a73} /* (12, 20, 8) {real, imag} */,
  {32'h3fa380b4, 32'h40513992} /* (12, 20, 7) {real, imag} */,
  {32'hbf492fae, 32'h3e674648} /* (12, 20, 6) {real, imag} */,
  {32'hc0a25162, 32'h3e299506} /* (12, 20, 5) {real, imag} */,
  {32'h3f9fa606, 32'h403c9b4f} /* (12, 20, 4) {real, imag} */,
  {32'h3fd51dd9, 32'h3f67d6d7} /* (12, 20, 3) {real, imag} */,
  {32'h3ecbbda3, 32'h3e9e8a03} /* (12, 20, 2) {real, imag} */,
  {32'h3fed8861, 32'hbf7f460e} /* (12, 20, 1) {real, imag} */,
  {32'hbe128460, 32'h3f598984} /* (12, 20, 0) {real, imag} */,
  {32'h3f11e5bb, 32'hbef9d52e} /* (12, 19, 31) {real, imag} */,
  {32'hbe9a21e5, 32'h4014432a} /* (12, 19, 30) {real, imag} */,
  {32'h3fc6c438, 32'hbff4bbac} /* (12, 19, 29) {real, imag} */,
  {32'h3fe80a22, 32'h4036ff78} /* (12, 19, 28) {real, imag} */,
  {32'h3d3b97bb, 32'h406d5839} /* (12, 19, 27) {real, imag} */,
  {32'h3f9235a4, 32'hc08c313a} /* (12, 19, 26) {real, imag} */,
  {32'hbf313b96, 32'hbfd47a8a} /* (12, 19, 25) {real, imag} */,
  {32'hbf201674, 32'hbc9e6b9e} /* (12, 19, 24) {real, imag} */,
  {32'hc046523c, 32'h3d1e0cee} /* (12, 19, 23) {real, imag} */,
  {32'h40a47bd1, 32'hc06c24b8} /* (12, 19, 22) {real, imag} */,
  {32'h3e55ccd1, 32'h40000efe} /* (12, 19, 21) {real, imag} */,
  {32'h3f24a0ad, 32'hbfa8144a} /* (12, 19, 20) {real, imag} */,
  {32'h3d360781, 32'h40222e50} /* (12, 19, 19) {real, imag} */,
  {32'h3f83989e, 32'h3f4b0909} /* (12, 19, 18) {real, imag} */,
  {32'h3fef02c6, 32'hbe89ffbd} /* (12, 19, 17) {real, imag} */,
  {32'hbf725cdc, 32'hbf023a15} /* (12, 19, 16) {real, imag} */,
  {32'hbfcb475d, 32'hbf02999c} /* (12, 19, 15) {real, imag} */,
  {32'h3f5463bc, 32'h3fb147c8} /* (12, 19, 14) {real, imag} */,
  {32'h3fccc05a, 32'hbdf8a4ef} /* (12, 19, 13) {real, imag} */,
  {32'h4053ad46, 32'h3f93df98} /* (12, 19, 12) {real, imag} */,
  {32'hbfd450e1, 32'hbf23fb04} /* (12, 19, 11) {real, imag} */,
  {32'hbd86df7b, 32'h3ed5eb44} /* (12, 19, 10) {real, imag} */,
  {32'hbf90f216, 32'h3e3a9aa3} /* (12, 19, 9) {real, imag} */,
  {32'hc01fd145, 32'h40555d0c} /* (12, 19, 8) {real, imag} */,
  {32'hbebb1cdc, 32'hbeb51690} /* (12, 19, 7) {real, imag} */,
  {32'hc009e29c, 32'hc03b30f5} /* (12, 19, 6) {real, imag} */,
  {32'hbf8829ee, 32'hbfc38690} /* (12, 19, 5) {real, imag} */,
  {32'h3efb1933, 32'hbeb9e83f} /* (12, 19, 4) {real, imag} */,
  {32'hbd0bc284, 32'hbff87f30} /* (12, 19, 3) {real, imag} */,
  {32'h40225349, 32'h3fcc53ec} /* (12, 19, 2) {real, imag} */,
  {32'h3faf2de7, 32'h40008c9c} /* (12, 19, 1) {real, imag} */,
  {32'hbe01ab71, 32'hc0321a55} /* (12, 19, 0) {real, imag} */,
  {32'h3f22f672, 32'h3f6c16c9} /* (12, 18, 31) {real, imag} */,
  {32'hbfb1008c, 32'hbc21e5d3} /* (12, 18, 30) {real, imag} */,
  {32'h403ffe8b, 32'hbf8e1c9d} /* (12, 18, 29) {real, imag} */,
  {32'h3f804535, 32'hbf8bec81} /* (12, 18, 28) {real, imag} */,
  {32'hbf4c9cc6, 32'h3fd6fffa} /* (12, 18, 27) {real, imag} */,
  {32'h3d60cd61, 32'h3e993f72} /* (12, 18, 26) {real, imag} */,
  {32'h3f6be1d4, 32'hbeb706c8} /* (12, 18, 25) {real, imag} */,
  {32'hbe4e8f41, 32'hbf01555d} /* (12, 18, 24) {real, imag} */,
  {32'h3f1ea82c, 32'h40192d24} /* (12, 18, 23) {real, imag} */,
  {32'hc06136d6, 32'hc02912dd} /* (12, 18, 22) {real, imag} */,
  {32'h3ffa9d8f, 32'h3ffb2d37} /* (12, 18, 21) {real, imag} */,
  {32'hbfedbbff, 32'hbe94e180} /* (12, 18, 20) {real, imag} */,
  {32'h3f1c9412, 32'h4003dbec} /* (12, 18, 19) {real, imag} */,
  {32'hbfd45b3d, 32'hc087fbd8} /* (12, 18, 18) {real, imag} */,
  {32'hbe0c09eb, 32'hbfac2e4c} /* (12, 18, 17) {real, imag} */,
  {32'hc0281794, 32'hbf009579} /* (12, 18, 16) {real, imag} */,
  {32'hc048af3c, 32'hbf760916} /* (12, 18, 15) {real, imag} */,
  {32'hbf54f018, 32'hc08ab0d7} /* (12, 18, 14) {real, imag} */,
  {32'h4028c5f0, 32'h4041dd30} /* (12, 18, 13) {real, imag} */,
  {32'hc042034d, 32'h3efd7aff} /* (12, 18, 12) {real, imag} */,
  {32'hc0157be1, 32'hbfd08331} /* (12, 18, 11) {real, imag} */,
  {32'h403f7356, 32'h405c7be4} /* (12, 18, 10) {real, imag} */,
  {32'h405e2676, 32'hbf481baf} /* (12, 18, 9) {real, imag} */,
  {32'hbf12ee71, 32'hbfa09f3a} /* (12, 18, 8) {real, imag} */,
  {32'h3f9b2fe5, 32'h3f1f8e88} /* (12, 18, 7) {real, imag} */,
  {32'hbeda4206, 32'hc06ca04a} /* (12, 18, 6) {real, imag} */,
  {32'h3f852203, 32'h3f906fe2} /* (12, 18, 5) {real, imag} */,
  {32'h3de36833, 32'hbfe38b7b} /* (12, 18, 4) {real, imag} */,
  {32'hbf631cfa, 32'h3f24b9b6} /* (12, 18, 3) {real, imag} */,
  {32'hbf68a7ac, 32'h403768e5} /* (12, 18, 2) {real, imag} */,
  {32'h4001f8cb, 32'hbe1995f4} /* (12, 18, 1) {real, imag} */,
  {32'h3f8d035b, 32'h3feccbf7} /* (12, 18, 0) {real, imag} */,
  {32'hbdd82d2e, 32'hbea95ddf} /* (12, 17, 31) {real, imag} */,
  {32'h40102cde, 32'hbf0abc52} /* (12, 17, 30) {real, imag} */,
  {32'hbf922855, 32'hbe21dc96} /* (12, 17, 29) {real, imag} */,
  {32'h3fba5641, 32'h40371b7d} /* (12, 17, 28) {real, imag} */,
  {32'h3f1076bc, 32'h3f1ad45c} /* (12, 17, 27) {real, imag} */,
  {32'h3e2e31c5, 32'h40508e94} /* (12, 17, 26) {real, imag} */,
  {32'hbfd2625e, 32'hc00e196c} /* (12, 17, 25) {real, imag} */,
  {32'hbf0e07ca, 32'h3f27c2f8} /* (12, 17, 24) {real, imag} */,
  {32'hc04ac0f5, 32'hc00c18c4} /* (12, 17, 23) {real, imag} */,
  {32'h4017b767, 32'h402d21dd} /* (12, 17, 22) {real, imag} */,
  {32'h3f4b36d3, 32'hbf93a560} /* (12, 17, 21) {real, imag} */,
  {32'h3fa42bd7, 32'h3f864ae4} /* (12, 17, 20) {real, imag} */,
  {32'h3f84a4b7, 32'h3edafa6e} /* (12, 17, 19) {real, imag} */,
  {32'hbf04ba9e, 32'h3f2af483} /* (12, 17, 18) {real, imag} */,
  {32'hbe25b574, 32'hbeb8c881} /* (12, 17, 17) {real, imag} */,
  {32'hbe3398f9, 32'h3d9fdcd7} /* (12, 17, 16) {real, imag} */,
  {32'h3fc38680, 32'hbf68160a} /* (12, 17, 15) {real, imag} */,
  {32'h403dc201, 32'h3fa53030} /* (12, 17, 14) {real, imag} */,
  {32'hbf6fe58c, 32'h3fa705cb} /* (12, 17, 13) {real, imag} */,
  {32'hbe450c16, 32'h3f4e608e} /* (12, 17, 12) {real, imag} */,
  {32'hbf289f01, 32'h3f27fb2e} /* (12, 17, 11) {real, imag} */,
  {32'hbf7e69a2, 32'h3f48d81c} /* (12, 17, 10) {real, imag} */,
  {32'hbf99d544, 32'h4014febb} /* (12, 17, 9) {real, imag} */,
  {32'h3c9a6d5a, 32'hc058a489} /* (12, 17, 8) {real, imag} */,
  {32'h4014e15a, 32'hbf0d8a31} /* (12, 17, 7) {real, imag} */,
  {32'h409965a7, 32'hbf82d5bf} /* (12, 17, 6) {real, imag} */,
  {32'hbfb00ee9, 32'h40098dda} /* (12, 17, 5) {real, imag} */,
  {32'hbed1794e, 32'h3c51137b} /* (12, 17, 4) {real, imag} */,
  {32'h3f8cb042, 32'hbf711a82} /* (12, 17, 3) {real, imag} */,
  {32'h3f0b78c5, 32'h3f09d159} /* (12, 17, 2) {real, imag} */,
  {32'hbf265b59, 32'hc03d077e} /* (12, 17, 1) {real, imag} */,
  {32'hbe98e0ce, 32'hbfdfebaf} /* (12, 17, 0) {real, imag} */,
  {32'h3f2bd5ba, 32'hbfc505db} /* (12, 16, 31) {real, imag} */,
  {32'h3ff2a6f4, 32'h401452a9} /* (12, 16, 30) {real, imag} */,
  {32'hbf8c45bb, 32'h3fa365ac} /* (12, 16, 29) {real, imag} */,
  {32'hc0045fd3, 32'hbf52b3ed} /* (12, 16, 28) {real, imag} */,
  {32'h3e43e027, 32'h4005f5d8} /* (12, 16, 27) {real, imag} */,
  {32'hbf1618e0, 32'hbf7c7489} /* (12, 16, 26) {real, imag} */,
  {32'h3f090236, 32'h3f65c0c7} /* (12, 16, 25) {real, imag} */,
  {32'hbfe8aa4f, 32'hbf807358} /* (12, 16, 24) {real, imag} */,
  {32'h3f830de3, 32'h3ec1d4e7} /* (12, 16, 23) {real, imag} */,
  {32'hbe502012, 32'hbfafdf01} /* (12, 16, 22) {real, imag} */,
  {32'h402bbc3a, 32'hbf5edddb} /* (12, 16, 21) {real, imag} */,
  {32'h40323e11, 32'hbd9dbb6e} /* (12, 16, 20) {real, imag} */,
  {32'hc03fa6da, 32'h40209f0e} /* (12, 16, 19) {real, imag} */,
  {32'h3f51f7f0, 32'hbf4c1a65} /* (12, 16, 18) {real, imag} */,
  {32'h3f8111e2, 32'h3fef683a} /* (12, 16, 17) {real, imag} */,
  {32'hbfc1df6b, 32'h3e4c9cc8} /* (12, 16, 16) {real, imag} */,
  {32'hbfe3a9ad, 32'h40095252} /* (12, 16, 15) {real, imag} */,
  {32'hbfc52942, 32'h3f3aa457} /* (12, 16, 14) {real, imag} */,
  {32'hc02bdce6, 32'h40042b6c} /* (12, 16, 13) {real, imag} */,
  {32'hbfef3e28, 32'hbf1cde93} /* (12, 16, 12) {real, imag} */,
  {32'h3e3ef911, 32'h3c910b05} /* (12, 16, 11) {real, imag} */,
  {32'hbf8238a3, 32'h3ed6269f} /* (12, 16, 10) {real, imag} */,
  {32'h3fc23be7, 32'h3ff3cfe6} /* (12, 16, 9) {real, imag} */,
  {32'hbe514099, 32'hbfeaf68d} /* (12, 16, 8) {real, imag} */,
  {32'h3ea90121, 32'hbfe0c467} /* (12, 16, 7) {real, imag} */,
  {32'hc00ebe0b, 32'hbfb71fcf} /* (12, 16, 6) {real, imag} */,
  {32'h3c3080e3, 32'h3f681d90} /* (12, 16, 5) {real, imag} */,
  {32'hbce569f3, 32'h3f94e02c} /* (12, 16, 4) {real, imag} */,
  {32'hbfdd63c1, 32'hbea39bad} /* (12, 16, 3) {real, imag} */,
  {32'hbe8b5bee, 32'h3f3dd707} /* (12, 16, 2) {real, imag} */,
  {32'h3f2529cf, 32'hbd00e017} /* (12, 16, 1) {real, imag} */,
  {32'h3f0abea4, 32'hbe3f69e3} /* (12, 16, 0) {real, imag} */,
  {32'h3f82bc03, 32'hbf2e4b04} /* (12, 15, 31) {real, imag} */,
  {32'h3f4e47c1, 32'h3f807a16} /* (12, 15, 30) {real, imag} */,
  {32'h3fb908cc, 32'hbea86160} /* (12, 15, 29) {real, imag} */,
  {32'h3f67a170, 32'h3eb16c01} /* (12, 15, 28) {real, imag} */,
  {32'hbf54a706, 32'h3ed843fe} /* (12, 15, 27) {real, imag} */,
  {32'hbf27d347, 32'h3fde5093} /* (12, 15, 26) {real, imag} */,
  {32'hbf59509b, 32'h3f9b4496} /* (12, 15, 25) {real, imag} */,
  {32'h401950fc, 32'h3f74ed77} /* (12, 15, 24) {real, imag} */,
  {32'h407dc0f5, 32'hbe4a5996} /* (12, 15, 23) {real, imag} */,
  {32'h3dd5e219, 32'hbf449978} /* (12, 15, 22) {real, imag} */,
  {32'hbfdd7160, 32'h3f8c6fee} /* (12, 15, 21) {real, imag} */,
  {32'hc0b07864, 32'h3ee245ee} /* (12, 15, 20) {real, imag} */,
  {32'h3ed0b70f, 32'h3ea1700d} /* (12, 15, 19) {real, imag} */,
  {32'h3f8f7b45, 32'hbf5ecf11} /* (12, 15, 18) {real, imag} */,
  {32'h3fe08baa, 32'h40379828} /* (12, 15, 17) {real, imag} */,
  {32'hbe56fdb3, 32'h3f526464} /* (12, 15, 16) {real, imag} */,
  {32'hbf048156, 32'hbfa07be2} /* (12, 15, 15) {real, imag} */,
  {32'hbf1767a6, 32'h3eb7ab6e} /* (12, 15, 14) {real, imag} */,
  {32'h40229a95, 32'hbfe83aca} /* (12, 15, 13) {real, imag} */,
  {32'h3f5f9209, 32'hc074ee95} /* (12, 15, 12) {real, imag} */,
  {32'h3f130728, 32'h400dac11} /* (12, 15, 11) {real, imag} */,
  {32'hc01e0c5c, 32'hbe727fde} /* (12, 15, 10) {real, imag} */,
  {32'hbe22222d, 32'h3f15f434} /* (12, 15, 9) {real, imag} */,
  {32'h3f1bfad5, 32'hc01d043f} /* (12, 15, 8) {real, imag} */,
  {32'h3e96f053, 32'h3fb53dbd} /* (12, 15, 7) {real, imag} */,
  {32'h3e9845de, 32'hc04c058e} /* (12, 15, 6) {real, imag} */,
  {32'hbf7dabd1, 32'h3fc179bb} /* (12, 15, 5) {real, imag} */,
  {32'hbff63321, 32'hc00ba828} /* (12, 15, 4) {real, imag} */,
  {32'hbf429e0a, 32'h3d813a4b} /* (12, 15, 3) {real, imag} */,
  {32'h3de3f83b, 32'h3e945530} /* (12, 15, 2) {real, imag} */,
  {32'h3e8fb452, 32'h3f54503a} /* (12, 15, 1) {real, imag} */,
  {32'h3fe05b1b, 32'h3d1a311e} /* (12, 15, 0) {real, imag} */,
  {32'hbfcaa632, 32'hbf863b1a} /* (12, 14, 31) {real, imag} */,
  {32'hbfbf4465, 32'h3fc080c5} /* (12, 14, 30) {real, imag} */,
  {32'h3e9d1181, 32'h3e8afa69} /* (12, 14, 29) {real, imag} */,
  {32'h404845f9, 32'hbd5ba71e} /* (12, 14, 28) {real, imag} */,
  {32'h3dbaa385, 32'hbffc648a} /* (12, 14, 27) {real, imag} */,
  {32'hc03fef6a, 32'h3f99230d} /* (12, 14, 26) {real, imag} */,
  {32'hbfa17348, 32'h3ebaa10f} /* (12, 14, 25) {real, imag} */,
  {32'hbe3d98f6, 32'h3f46d18f} /* (12, 14, 24) {real, imag} */,
  {32'hc01ad171, 32'h3f7d4db5} /* (12, 14, 23) {real, imag} */,
  {32'hc0821b83, 32'h3e161651} /* (12, 14, 22) {real, imag} */,
  {32'h4059893c, 32'hbfef379b} /* (12, 14, 21) {real, imag} */,
  {32'h40267253, 32'hbf83e160} /* (12, 14, 20) {real, imag} */,
  {32'h4014d0bb, 32'hc0007a47} /* (12, 14, 19) {real, imag} */,
  {32'h3e83a305, 32'h3e384be8} /* (12, 14, 18) {real, imag} */,
  {32'hbf307fc3, 32'h3f5a5ff6} /* (12, 14, 17) {real, imag} */,
  {32'hbf119345, 32'hc0116ef4} /* (12, 14, 16) {real, imag} */,
  {32'h4091ce37, 32'hc041802a} /* (12, 14, 15) {real, imag} */,
  {32'h3fd90387, 32'hc06eb69a} /* (12, 14, 14) {real, imag} */,
  {32'h3fe9b6b2, 32'h3febe771} /* (12, 14, 13) {real, imag} */,
  {32'h3e728038, 32'h3f960282} /* (12, 14, 12) {real, imag} */,
  {32'h3fb8e01a, 32'h3f97ef20} /* (12, 14, 11) {real, imag} */,
  {32'hbf81819c, 32'h3f8fa31e} /* (12, 14, 10) {real, imag} */,
  {32'hc02a1c2b, 32'h3fb91066} /* (12, 14, 9) {real, imag} */,
  {32'h3f5f3b1c, 32'h3dfd3135} /* (12, 14, 8) {real, imag} */,
  {32'hc0826b3d, 32'hbde5b106} /* (12, 14, 7) {real, imag} */,
  {32'hbf87da4f, 32'hc002a569} /* (12, 14, 6) {real, imag} */,
  {32'hbf973665, 32'hc0934b76} /* (12, 14, 5) {real, imag} */,
  {32'hc01d59f0, 32'h3fe76d2b} /* (12, 14, 4) {real, imag} */,
  {32'hbfbaf525, 32'hbdada517} /* (12, 14, 3) {real, imag} */,
  {32'h3faa6259, 32'hbf7c4ec0} /* (12, 14, 2) {real, imag} */,
  {32'h3eca8ee3, 32'hbe8b0c63} /* (12, 14, 1) {real, imag} */,
  {32'hbe86f147, 32'h3f8e6d70} /* (12, 14, 0) {real, imag} */,
  {32'hc02c0579, 32'hbf25da9e} /* (12, 13, 31) {real, imag} */,
  {32'h3fd72be4, 32'h3f515754} /* (12, 13, 30) {real, imag} */,
  {32'hc03e3e7d, 32'h40428389} /* (12, 13, 29) {real, imag} */,
  {32'hbf41d0e6, 32'hbe25b63d} /* (12, 13, 28) {real, imag} */,
  {32'hc0160970, 32'h4033612d} /* (12, 13, 27) {real, imag} */,
  {32'hbf9715b7, 32'h40444c45} /* (12, 13, 26) {real, imag} */,
  {32'h3e7d3b45, 32'h3eee89c6} /* (12, 13, 25) {real, imag} */,
  {32'h3fc686c5, 32'h3d9753e2} /* (12, 13, 24) {real, imag} */,
  {32'h3faf5f47, 32'hbf628b0f} /* (12, 13, 23) {real, imag} */,
  {32'h3e64195b, 32'h3ebcb788} /* (12, 13, 22) {real, imag} */,
  {32'h406d3527, 32'h3e810a5f} /* (12, 13, 21) {real, imag} */,
  {32'hbebf6773, 32'h4046b167} /* (12, 13, 20) {real, imag} */,
  {32'hbfdf40fa, 32'h3f7903a5} /* (12, 13, 19) {real, imag} */,
  {32'hc01f549f, 32'h401827df} /* (12, 13, 18) {real, imag} */,
  {32'hbf89d200, 32'hbfae348d} /* (12, 13, 17) {real, imag} */,
  {32'hc02a11ba, 32'h3f0a21d0} /* (12, 13, 16) {real, imag} */,
  {32'hbf9421d9, 32'h3f974416} /* (12, 13, 15) {real, imag} */,
  {32'hbf771f1f, 32'hbeb87b44} /* (12, 13, 14) {real, imag} */,
  {32'hbe76b5e8, 32'h3ec06895} /* (12, 13, 13) {real, imag} */,
  {32'hbe848ae0, 32'hbfe0170e} /* (12, 13, 12) {real, imag} */,
  {32'h40252f6f, 32'h40061470} /* (12, 13, 11) {real, imag} */,
  {32'h3f23eedb, 32'hbfd4214c} /* (12, 13, 10) {real, imag} */,
  {32'h401e23ca, 32'h3e2abb57} /* (12, 13, 9) {real, imag} */,
  {32'h4008858a, 32'hbd892e22} /* (12, 13, 8) {real, imag} */,
  {32'h3fb49727, 32'hbf818ab4} /* (12, 13, 7) {real, imag} */,
  {32'h3e88a4f6, 32'h3ea70d50} /* (12, 13, 6) {real, imag} */,
  {32'h4096f567, 32'hbf16e7b9} /* (12, 13, 5) {real, imag} */,
  {32'hbfa00a1c, 32'hc0441b7e} /* (12, 13, 4) {real, imag} */,
  {32'h3e945014, 32'hbffaf401} /* (12, 13, 3) {real, imag} */,
  {32'hbee45358, 32'hbf1221ba} /* (12, 13, 2) {real, imag} */,
  {32'hbf95fe39, 32'h400f57db} /* (12, 13, 1) {real, imag} */,
  {32'h400cec7f, 32'h3e503136} /* (12, 13, 0) {real, imag} */,
  {32'hbf9cf633, 32'h40063484} /* (12, 12, 31) {real, imag} */,
  {32'h3e80b3c2, 32'hbf70fa74} /* (12, 12, 30) {real, imag} */,
  {32'h4004ecaa, 32'h40055d11} /* (12, 12, 29) {real, imag} */,
  {32'hc00cb56f, 32'h3f4ee717} /* (12, 12, 28) {real, imag} */,
  {32'hbf1adf75, 32'hbf915cad} /* (12, 12, 27) {real, imag} */,
  {32'h3f0197a2, 32'hbfd411f5} /* (12, 12, 26) {real, imag} */,
  {32'hbeaab354, 32'hbfefa64f} /* (12, 12, 25) {real, imag} */,
  {32'h3f4c6b67, 32'hbfc53b3e} /* (12, 12, 24) {real, imag} */,
  {32'hbfc4ea4f, 32'hbfdf2169} /* (12, 12, 23) {real, imag} */,
  {32'h3fb10c91, 32'hbfffb21b} /* (12, 12, 22) {real, imag} */,
  {32'h3cb41ef0, 32'h3cf222ea} /* (12, 12, 21) {real, imag} */,
  {32'h3eb11e9f, 32'h3fe56224} /* (12, 12, 20) {real, imag} */,
  {32'hbfbaf1f2, 32'hc0077ac1} /* (12, 12, 19) {real, imag} */,
  {32'hc030fa65, 32'h3f172d66} /* (12, 12, 18) {real, imag} */,
  {32'hbfbe876d, 32'hbe49bcef} /* (12, 12, 17) {real, imag} */,
  {32'h401cbca5, 32'h3f921c15} /* (12, 12, 16) {real, imag} */,
  {32'h3fa55409, 32'hbfaa9d65} /* (12, 12, 15) {real, imag} */,
  {32'hc0019e27, 32'hc00c02c3} /* (12, 12, 14) {real, imag} */,
  {32'hc01ce977, 32'hbe1a3e83} /* (12, 12, 13) {real, imag} */,
  {32'hc06ea7c4, 32'hbfc5f4f4} /* (12, 12, 12) {real, imag} */,
  {32'hbdc39445, 32'hbff18ca1} /* (12, 12, 11) {real, imag} */,
  {32'hc00f083d, 32'h405bc8eb} /* (12, 12, 10) {real, imag} */,
  {32'h409d855e, 32'hc03a521b} /* (12, 12, 9) {real, imag} */,
  {32'hbf74fbef, 32'h3e54f0e2} /* (12, 12, 8) {real, imag} */,
  {32'hbee031be, 32'h3f0534c1} /* (12, 12, 7) {real, imag} */,
  {32'hbec050b8, 32'hc0769b75} /* (12, 12, 6) {real, imag} */,
  {32'h40060571, 32'hbfa338aa} /* (12, 12, 5) {real, imag} */,
  {32'hbf35fc58, 32'hbe98941d} /* (12, 12, 4) {real, imag} */,
  {32'h4041e546, 32'h401919cf} /* (12, 12, 3) {real, imag} */,
  {32'hbec8c877, 32'hbfe1330d} /* (12, 12, 2) {real, imag} */,
  {32'hbf373c8c, 32'hbf6b6c7b} /* (12, 12, 1) {real, imag} */,
  {32'h40295a6f, 32'h408729c3} /* (12, 12, 0) {real, imag} */,
  {32'h3f09371e, 32'hc00a3a31} /* (12, 11, 31) {real, imag} */,
  {32'hc02a587e, 32'hbf99edf4} /* (12, 11, 30) {real, imag} */,
  {32'h3fd68f45, 32'hbf7790a9} /* (12, 11, 29) {real, imag} */,
  {32'hbfef6cea, 32'h3f023bce} /* (12, 11, 28) {real, imag} */,
  {32'h3f094f89, 32'h3fcbc111} /* (12, 11, 27) {real, imag} */,
  {32'h3f784c89, 32'hbe315bfa} /* (12, 11, 26) {real, imag} */,
  {32'h408108bf, 32'hbea2bf5f} /* (12, 11, 25) {real, imag} */,
  {32'h3f126521, 32'hc01a5a9f} /* (12, 11, 24) {real, imag} */,
  {32'hbf81d346, 32'h3ef56ef7} /* (12, 11, 23) {real, imag} */,
  {32'h4046791b, 32'h3f923cc3} /* (12, 11, 22) {real, imag} */,
  {32'h400fce49, 32'hc00c240c} /* (12, 11, 21) {real, imag} */,
  {32'h4070927a, 32'h40394cbf} /* (12, 11, 20) {real, imag} */,
  {32'hbe81fc22, 32'h405efddf} /* (12, 11, 19) {real, imag} */,
  {32'h3fddada8, 32'hbeed6f10} /* (12, 11, 18) {real, imag} */,
  {32'hbe4d47fc, 32'hbf839b31} /* (12, 11, 17) {real, imag} */,
  {32'h3e941d7c, 32'h3fc02c9e} /* (12, 11, 16) {real, imag} */,
  {32'hbf70ac81, 32'hc00daaa9} /* (12, 11, 15) {real, imag} */,
  {32'h3fb5b406, 32'h3fcb0163} /* (12, 11, 14) {real, imag} */,
  {32'hbfc4bf51, 32'hbe894e1f} /* (12, 11, 13) {real, imag} */,
  {32'h402d8c4f, 32'hbf272085} /* (12, 11, 12) {real, imag} */,
  {32'h3f2283c0, 32'h3f947792} /* (12, 11, 11) {real, imag} */,
  {32'hc03af8fb, 32'hbf3b3951} /* (12, 11, 10) {real, imag} */,
  {32'h4095d4ae, 32'h40866ad3} /* (12, 11, 9) {real, imag} */,
  {32'h4020d5c3, 32'h3fba3023} /* (12, 11, 8) {real, imag} */,
  {32'hc0040cf5, 32'h3fd63479} /* (12, 11, 7) {real, imag} */,
  {32'hc067109f, 32'h3df94e45} /* (12, 11, 6) {real, imag} */,
  {32'h3ef71dde, 32'h3f91d6db} /* (12, 11, 5) {real, imag} */,
  {32'h3e1259b6, 32'hbf69a7b1} /* (12, 11, 4) {real, imag} */,
  {32'h403a6a17, 32'h3fcb26af} /* (12, 11, 3) {real, imag} */,
  {32'h401a659c, 32'h3fc4d913} /* (12, 11, 2) {real, imag} */,
  {32'hbe5ba1c6, 32'hbf38645d} /* (12, 11, 1) {real, imag} */,
  {32'hbf0ae548, 32'hc032bcf6} /* (12, 11, 0) {real, imag} */,
  {32'hc00214f3, 32'h3ec91c52} /* (12, 10, 31) {real, imag} */,
  {32'hbedecf38, 32'h3f559ddd} /* (12, 10, 30) {real, imag} */,
  {32'hbebd3cf4, 32'hbf99591a} /* (12, 10, 29) {real, imag} */,
  {32'h3f16ee62, 32'hbef316a6} /* (12, 10, 28) {real, imag} */,
  {32'hbf330825, 32'h407a452f} /* (12, 10, 27) {real, imag} */,
  {32'hc014f1cb, 32'hbe6b2ecf} /* (12, 10, 26) {real, imag} */,
  {32'h3e583a26, 32'hbf70fa4b} /* (12, 10, 25) {real, imag} */,
  {32'hbfab611f, 32'hc0086432} /* (12, 10, 24) {real, imag} */,
  {32'h3e7f4eb1, 32'hbfce8f31} /* (12, 10, 23) {real, imag} */,
  {32'h3f7a0a57, 32'hbe6f257e} /* (12, 10, 22) {real, imag} */,
  {32'h3fd026b8, 32'h3dcd44bf} /* (12, 10, 21) {real, imag} */,
  {32'h3f308b5f, 32'hbf611dd4} /* (12, 10, 20) {real, imag} */,
  {32'h400eed35, 32'h3fc53f1e} /* (12, 10, 19) {real, imag} */,
  {32'hc0244066, 32'hbfd542b2} /* (12, 10, 18) {real, imag} */,
  {32'hbedd057b, 32'hbbaf5c9b} /* (12, 10, 17) {real, imag} */,
  {32'hbfb0d33f, 32'h3e37b6e0} /* (12, 10, 16) {real, imag} */,
  {32'h4049b8b8, 32'h404fe67b} /* (12, 10, 15) {real, imag} */,
  {32'h40a7542e, 32'hbfb605a4} /* (12, 10, 14) {real, imag} */,
  {32'hbfafe83f, 32'h3d4598f5} /* (12, 10, 13) {real, imag} */,
  {32'hc01f32d1, 32'h40538daa} /* (12, 10, 12) {real, imag} */,
  {32'hbf272fa6, 32'hbd36a3b2} /* (12, 10, 11) {real, imag} */,
  {32'hbedf6e4c, 32'h3f226fd3} /* (12, 10, 10) {real, imag} */,
  {32'hc0153672, 32'hbe2850a5} /* (12, 10, 9) {real, imag} */,
  {32'hbe83165e, 32'hbf8e2eee} /* (12, 10, 8) {real, imag} */,
  {32'hbf7ac57b, 32'hbfa73ee8} /* (12, 10, 7) {real, imag} */,
  {32'hc081171b, 32'hbf541278} /* (12, 10, 6) {real, imag} */,
  {32'hbfc4dbe6, 32'h3fc01e74} /* (12, 10, 5) {real, imag} */,
  {32'h401ab7ad, 32'hbf40ed81} /* (12, 10, 4) {real, imag} */,
  {32'hc03b388c, 32'hbf9115ef} /* (12, 10, 3) {real, imag} */,
  {32'h3fc092fb, 32'h3f74c236} /* (12, 10, 2) {real, imag} */,
  {32'hbfa54dcd, 32'hc01de49d} /* (12, 10, 1) {real, imag} */,
  {32'hbf314444, 32'hbf172a66} /* (12, 10, 0) {real, imag} */,
  {32'hbfb67aef, 32'h3f9490d7} /* (12, 9, 31) {real, imag} */,
  {32'h3e00e999, 32'h408e209e} /* (12, 9, 30) {real, imag} */,
  {32'h3f5439a7, 32'h3fb7285f} /* (12, 9, 29) {real, imag} */,
  {32'h3de961e0, 32'h3f5bcbb7} /* (12, 9, 28) {real, imag} */,
  {32'hbe1e6095, 32'h3f8c3d84} /* (12, 9, 27) {real, imag} */,
  {32'hbe459573, 32'h3df7a872} /* (12, 9, 26) {real, imag} */,
  {32'hbf1e55b5, 32'hc03f2222} /* (12, 9, 25) {real, imag} */,
  {32'h3facef0c, 32'h3f524124} /* (12, 9, 24) {real, imag} */,
  {32'hc0850b75, 32'h4001dd52} /* (12, 9, 23) {real, imag} */,
  {32'hbef2cef3, 32'hbedd8b62} /* (12, 9, 22) {real, imag} */,
  {32'hbe37c96d, 32'hbea351d0} /* (12, 9, 21) {real, imag} */,
  {32'hbf31ad54, 32'hbfbeaac0} /* (12, 9, 20) {real, imag} */,
  {32'h40367ecd, 32'hbf8e503e} /* (12, 9, 19) {real, imag} */,
  {32'h3e9a4dcf, 32'hbf01acf4} /* (12, 9, 18) {real, imag} */,
  {32'h3e346baf, 32'hbff90358} /* (12, 9, 17) {real, imag} */,
  {32'h3ec67b46, 32'h3f57eb2c} /* (12, 9, 16) {real, imag} */,
  {32'hbf906f97, 32'h3f1ecf79} /* (12, 9, 15) {real, imag} */,
  {32'hbf9ab209, 32'h40488f7a} /* (12, 9, 14) {real, imag} */,
  {32'hc017dfbd, 32'h3fbb1acc} /* (12, 9, 13) {real, imag} */,
  {32'hbfbb50c9, 32'hbf1f9274} /* (12, 9, 12) {real, imag} */,
  {32'h3f5d7720, 32'h40603f07} /* (12, 9, 11) {real, imag} */,
  {32'hc01986bb, 32'h3fd3bf31} /* (12, 9, 10) {real, imag} */,
  {32'hbfb0e3b9, 32'hbf7a8c1f} /* (12, 9, 9) {real, imag} */,
  {32'hbfba0627, 32'hbe93b85f} /* (12, 9, 8) {real, imag} */,
  {32'hbfc6fdba, 32'hbec6e3ed} /* (12, 9, 7) {real, imag} */,
  {32'h3fdb3324, 32'hbf160293} /* (12, 9, 6) {real, imag} */,
  {32'h405839de, 32'hbfd6a5bf} /* (12, 9, 5) {real, imag} */,
  {32'hbfd0767e, 32'h3f80ef85} /* (12, 9, 4) {real, imag} */,
  {32'hbfab0b3d, 32'hc04e546a} /* (12, 9, 3) {real, imag} */,
  {32'hbf0a5037, 32'hbee44d2c} /* (12, 9, 2) {real, imag} */,
  {32'hc0708f0d, 32'hbfd19d44} /* (12, 9, 1) {real, imag} */,
  {32'h3ef3b4b2, 32'hbfdbebc3} /* (12, 9, 0) {real, imag} */,
  {32'hbf5a1dda, 32'h3feade83} /* (12, 8, 31) {real, imag} */,
  {32'hbff070a9, 32'hc004c3b4} /* (12, 8, 30) {real, imag} */,
  {32'hbf8e2801, 32'h3f7db5c9} /* (12, 8, 29) {real, imag} */,
  {32'h3faa8367, 32'h3f588590} /* (12, 8, 28) {real, imag} */,
  {32'hc00a6fef, 32'h3e8643ab} /* (12, 8, 27) {real, imag} */,
  {32'h3ee98aff, 32'h3fe825bc} /* (12, 8, 26) {real, imag} */,
  {32'h3faacda1, 32'hbec7b355} /* (12, 8, 25) {real, imag} */,
  {32'hbef13d6f, 32'h40244269} /* (12, 8, 24) {real, imag} */,
  {32'h3dc3e983, 32'h3f937a11} /* (12, 8, 23) {real, imag} */,
  {32'hbff9a9d2, 32'hbef48c00} /* (12, 8, 22) {real, imag} */,
  {32'h3e104349, 32'h3dfabeb7} /* (12, 8, 21) {real, imag} */,
  {32'h3e722b6e, 32'h3df55a55} /* (12, 8, 20) {real, imag} */,
  {32'hbf7b35fe, 32'hbecc875c} /* (12, 8, 19) {real, imag} */,
  {32'h3f1ee021, 32'hbf0a6607} /* (12, 8, 18) {real, imag} */,
  {32'h3f6ec3b8, 32'h3f83b9f4} /* (12, 8, 17) {real, imag} */,
  {32'hbf4aeadb, 32'h4011d567} /* (12, 8, 16) {real, imag} */,
  {32'hbeb8073d, 32'h3fa83e56} /* (12, 8, 15) {real, imag} */,
  {32'hbf9d6d81, 32'h40114813} /* (12, 8, 14) {real, imag} */,
  {32'h3fadd750, 32'hbf33c075} /* (12, 8, 13) {real, imag} */,
  {32'h40266fad, 32'hbf7cda85} /* (12, 8, 12) {real, imag} */,
  {32'h3f234298, 32'h3dd98936} /* (12, 8, 11) {real, imag} */,
  {32'hbfa75b11, 32'hbf11d415} /* (12, 8, 10) {real, imag} */,
  {32'hc02c5c66, 32'hbf9b4ec9} /* (12, 8, 9) {real, imag} */,
  {32'hbecd896e, 32'h3fb52feb} /* (12, 8, 8) {real, imag} */,
  {32'h400e24ab, 32'h3f7ab8ac} /* (12, 8, 7) {real, imag} */,
  {32'h40069077, 32'h3e7774dc} /* (12, 8, 6) {real, imag} */,
  {32'h3f378914, 32'h3fb4bb25} /* (12, 8, 5) {real, imag} */,
  {32'h402a4d3b, 32'hbf8b125e} /* (12, 8, 4) {real, imag} */,
  {32'h4035c874, 32'h3fa39a89} /* (12, 8, 3) {real, imag} */,
  {32'h405db04f, 32'hc00e60a2} /* (12, 8, 2) {real, imag} */,
  {32'h3e12cb44, 32'hbf1c58c9} /* (12, 8, 1) {real, imag} */,
  {32'h3f034000, 32'hbd8ec137} /* (12, 8, 0) {real, imag} */,
  {32'h3fb6676d, 32'h3f76033b} /* (12, 7, 31) {real, imag} */,
  {32'hbe1edd95, 32'hbf3bff19} /* (12, 7, 30) {real, imag} */,
  {32'h3f263049, 32'hbfbb7dae} /* (12, 7, 29) {real, imag} */,
  {32'h3f93fd5f, 32'h3fa44649} /* (12, 7, 28) {real, imag} */,
  {32'h3fb0d042, 32'h403a4232} /* (12, 7, 27) {real, imag} */,
  {32'hc0135c0f, 32'hbf3dbabe} /* (12, 7, 26) {real, imag} */,
  {32'hbfc3bca9, 32'hbff76edc} /* (12, 7, 25) {real, imag} */,
  {32'hbffa4101, 32'h4045bf51} /* (12, 7, 24) {real, imag} */,
  {32'h40842474, 32'h3e298107} /* (12, 7, 23) {real, imag} */,
  {32'h3f2b94b6, 32'hbf9d819d} /* (12, 7, 22) {real, imag} */,
  {32'h3f21ec92, 32'hc006cf7c} /* (12, 7, 21) {real, imag} */,
  {32'hbf5a15f1, 32'h3fb91a42} /* (12, 7, 20) {real, imag} */,
  {32'h3f621fed, 32'h3d09c997} /* (12, 7, 19) {real, imag} */,
  {32'hc06974c7, 32'hbec64aaa} /* (12, 7, 18) {real, imag} */,
  {32'hbf018ddd, 32'hbfbfa66d} /* (12, 7, 17) {real, imag} */,
  {32'h4005ed5a, 32'hc03eef9a} /* (12, 7, 16) {real, imag} */,
  {32'h3f9b4b43, 32'h3fc30ed3} /* (12, 7, 15) {real, imag} */,
  {32'h3fd3fa65, 32'hbfc83961} /* (12, 7, 14) {real, imag} */,
  {32'hbe355215, 32'hbfea9572} /* (12, 7, 13) {real, imag} */,
  {32'h4052830c, 32'h3f5d9140} /* (12, 7, 12) {real, imag} */,
  {32'hc02107df, 32'h3e9a164e} /* (12, 7, 11) {real, imag} */,
  {32'hbfc0db66, 32'h3f9d9670} /* (12, 7, 10) {real, imag} */,
  {32'hbfbf57a3, 32'hbe3668f4} /* (12, 7, 9) {real, imag} */,
  {32'h401fbe62, 32'hbf194b0b} /* (12, 7, 8) {real, imag} */,
  {32'hbf936138, 32'hbf9c0509} /* (12, 7, 7) {real, imag} */,
  {32'hbfe3fccb, 32'h3f6ec713} /* (12, 7, 6) {real, imag} */,
  {32'h3f5ca7fa, 32'hbe4bb56e} /* (12, 7, 5) {real, imag} */,
  {32'h3ed77ac6, 32'hbfee76ff} /* (12, 7, 4) {real, imag} */,
  {32'h3fd56dd6, 32'hbff3eaf3} /* (12, 7, 3) {real, imag} */,
  {32'hc007d201, 32'h40118c4a} /* (12, 7, 2) {real, imag} */,
  {32'hc00d10f4, 32'h3ffc5d0c} /* (12, 7, 1) {real, imag} */,
  {32'h3fd8faaa, 32'hc04fed1c} /* (12, 7, 0) {real, imag} */,
  {32'h3fa1c29f, 32'hc01d5b98} /* (12, 6, 31) {real, imag} */,
  {32'h3f68096a, 32'h3ff84dca} /* (12, 6, 30) {real, imag} */,
  {32'hc0092a5c, 32'hbeed1535} /* (12, 6, 29) {real, imag} */,
  {32'hbf68e345, 32'hbf86f7f6} /* (12, 6, 28) {real, imag} */,
  {32'h3f8340e3, 32'hbfd22f6d} /* (12, 6, 27) {real, imag} */,
  {32'h3fbfefe9, 32'hc03593e1} /* (12, 6, 26) {real, imag} */,
  {32'h3d12ce04, 32'h3fe74235} /* (12, 6, 25) {real, imag} */,
  {32'hc03cc10c, 32'hc01825a2} /* (12, 6, 24) {real, imag} */,
  {32'h3f25dfda, 32'h3fcd5946} /* (12, 6, 23) {real, imag} */,
  {32'h3fcf2a29, 32'h3e1f7fdb} /* (12, 6, 22) {real, imag} */,
  {32'h3f7becd5, 32'h3fd74261} /* (12, 6, 21) {real, imag} */,
  {32'hbf6b37be, 32'hbfd968f5} /* (12, 6, 20) {real, imag} */,
  {32'h3f9361d1, 32'h40003763} /* (12, 6, 19) {real, imag} */,
  {32'h3f59feb2, 32'hbf93ffbf} /* (12, 6, 18) {real, imag} */,
  {32'hbfe15c8d, 32'h3e3809fb} /* (12, 6, 17) {real, imag} */,
  {32'hbf1cbb02, 32'h3f00fd46} /* (12, 6, 16) {real, imag} */,
  {32'h3eea9c46, 32'hbe0c2d9e} /* (12, 6, 15) {real, imag} */,
  {32'h3f22720e, 32'h4035c5a3} /* (12, 6, 14) {real, imag} */,
  {32'h3f98e002, 32'h3e4a63ce} /* (12, 6, 13) {real, imag} */,
  {32'hbf2ec99c, 32'hbf6f0b45} /* (12, 6, 12) {real, imag} */,
  {32'hc03a5a4b, 32'hbd119ab4} /* (12, 6, 11) {real, imag} */,
  {32'h3fafd7d7, 32'h3e514aa9} /* (12, 6, 10) {real, imag} */,
  {32'h3f269043, 32'h3f7f986c} /* (12, 6, 9) {real, imag} */,
  {32'h3f10724e, 32'h3f9bf8ad} /* (12, 6, 8) {real, imag} */,
  {32'hc01c909c, 32'h3f1ecd9f} /* (12, 6, 7) {real, imag} */,
  {32'h4018619a, 32'hbf169bf2} /* (12, 6, 6) {real, imag} */,
  {32'hc061b7e0, 32'hbf04e562} /* (12, 6, 5) {real, imag} */,
  {32'h3f14f106, 32'hbdc3c8dd} /* (12, 6, 4) {real, imag} */,
  {32'h3ede7837, 32'h3e944ad3} /* (12, 6, 3) {real, imag} */,
  {32'h3fec6c83, 32'h3ffc75d5} /* (12, 6, 2) {real, imag} */,
  {32'hc0010780, 32'hbffc2d41} /* (12, 6, 1) {real, imag} */,
  {32'hbfddf40e, 32'h3ff7b456} /* (12, 6, 0) {real, imag} */,
  {32'h40008b5a, 32'hc019bd99} /* (12, 5, 31) {real, imag} */,
  {32'h3fcc72ca, 32'h3eba528a} /* (12, 5, 30) {real, imag} */,
  {32'h3ed4a938, 32'h406dc03d} /* (12, 5, 29) {real, imag} */,
  {32'h3f907caa, 32'h400a0833} /* (12, 5, 28) {real, imag} */,
  {32'hbfa2bf12, 32'hbf531cf2} /* (12, 5, 27) {real, imag} */,
  {32'h4010b6bd, 32'h3fa15a67} /* (12, 5, 26) {real, imag} */,
  {32'h3eed4340, 32'hc01570ff} /* (12, 5, 25) {real, imag} */,
  {32'hbe93a6bd, 32'hc03aa7ff} /* (12, 5, 24) {real, imag} */,
  {32'hc0927f5b, 32'h3fec55e8} /* (12, 5, 23) {real, imag} */,
  {32'h3ff6409e, 32'h40af30d0} /* (12, 5, 22) {real, imag} */,
  {32'hbfb5ebca, 32'hbfb16615} /* (12, 5, 21) {real, imag} */,
  {32'hc073d7e6, 32'hbf28e908} /* (12, 5, 20) {real, imag} */,
  {32'h3e3c747e, 32'hbf6c55cc} /* (12, 5, 19) {real, imag} */,
  {32'hbe5c12b3, 32'hc0124dd9} /* (12, 5, 18) {real, imag} */,
  {32'h401e10b9, 32'h3f900563} /* (12, 5, 17) {real, imag} */,
  {32'h3e5fbe59, 32'h3ef76083} /* (12, 5, 16) {real, imag} */,
  {32'hbff2867e, 32'hbffad4ce} /* (12, 5, 15) {real, imag} */,
  {32'h3fb74b8c, 32'hbfd73a7e} /* (12, 5, 14) {real, imag} */,
  {32'hbed16b71, 32'hc00ec0b8} /* (12, 5, 13) {real, imag} */,
  {32'h4035c874, 32'h3ff11c40} /* (12, 5, 12) {real, imag} */,
  {32'h401c046c, 32'hbf320a98} /* (12, 5, 11) {real, imag} */,
  {32'h3f1919eb, 32'hbe656db9} /* (12, 5, 10) {real, imag} */,
  {32'hbf6affcf, 32'h3f91e0c0} /* (12, 5, 9) {real, imag} */,
  {32'hbf8903ba, 32'h401bd864} /* (12, 5, 8) {real, imag} */,
  {32'h4039fb0c, 32'h3f08fa03} /* (12, 5, 7) {real, imag} */,
  {32'hc09c61dc, 32'hbeca85bd} /* (12, 5, 6) {real, imag} */,
  {32'hbfe149bf, 32'h3f6afc48} /* (12, 5, 5) {real, imag} */,
  {32'hbf267282, 32'hbf215094} /* (12, 5, 4) {real, imag} */,
  {32'hbf16b030, 32'h4072983e} /* (12, 5, 3) {real, imag} */,
  {32'hc064e193, 32'hc05a58ea} /* (12, 5, 2) {real, imag} */,
  {32'h3fc48926, 32'hc032e290} /* (12, 5, 1) {real, imag} */,
  {32'hbf6d011d, 32'hbf8266de} /* (12, 5, 0) {real, imag} */,
  {32'h3e989e6a, 32'hbf0f8922} /* (12, 4, 31) {real, imag} */,
  {32'h3f406762, 32'hc02ad6c4} /* (12, 4, 30) {real, imag} */,
  {32'hc039f364, 32'h3febf440} /* (12, 4, 29) {real, imag} */,
  {32'hc0184694, 32'h4067c80f} /* (12, 4, 28) {real, imag} */,
  {32'h3fb6d2dd, 32'hbf59475f} /* (12, 4, 27) {real, imag} */,
  {32'h3f462836, 32'hbf0b4c6d} /* (12, 4, 26) {real, imag} */,
  {32'hbf3ca5a8, 32'h3e42904a} /* (12, 4, 25) {real, imag} */,
  {32'h3f4d8bca, 32'h3f67341e} /* (12, 4, 24) {real, imag} */,
  {32'h4017c7fd, 32'hbf322b80} /* (12, 4, 23) {real, imag} */,
  {32'hbf8999eb, 32'h3f8e79c7} /* (12, 4, 22) {real, imag} */,
  {32'h406186b9, 32'hbeb21419} /* (12, 4, 21) {real, imag} */,
  {32'hc0286788, 32'h3fa20209} /* (12, 4, 20) {real, imag} */,
  {32'hc011a5e3, 32'h3f7f8585} /* (12, 4, 19) {real, imag} */,
  {32'hbeefc9e4, 32'hc071ce35} /* (12, 4, 18) {real, imag} */,
  {32'hbbd4998d, 32'h3df796a5} /* (12, 4, 17) {real, imag} */,
  {32'h3e2a3758, 32'hbf479526} /* (12, 4, 16) {real, imag} */,
  {32'h3e986cca, 32'hc00154b4} /* (12, 4, 15) {real, imag} */,
  {32'h3de92f93, 32'h3e8b04f3} /* (12, 4, 14) {real, imag} */,
  {32'h3c8d087b, 32'hbec7c17c} /* (12, 4, 13) {real, imag} */,
  {32'h3db989a1, 32'h3ef9e80f} /* (12, 4, 12) {real, imag} */,
  {32'h3f103b26, 32'h404b2eac} /* (12, 4, 11) {real, imag} */,
  {32'h3fc1b747, 32'h3f8fca49} /* (12, 4, 10) {real, imag} */,
  {32'h3fa2da65, 32'hbf9a52e4} /* (12, 4, 9) {real, imag} */,
  {32'h404c08f7, 32'h3f42f251} /* (12, 4, 8) {real, imag} */,
  {32'hbdd8e6b2, 32'hbfa00466} /* (12, 4, 7) {real, imag} */,
  {32'h3f66ef2f, 32'hbf9168e2} /* (12, 4, 6) {real, imag} */,
  {32'hbf3c1074, 32'h4053928b} /* (12, 4, 5) {real, imag} */,
  {32'hbf90a112, 32'hbf032f17} /* (12, 4, 4) {real, imag} */,
  {32'h3fe8ee78, 32'h3f84aa7b} /* (12, 4, 3) {real, imag} */,
  {32'h3e7c9985, 32'h401d3901} /* (12, 4, 2) {real, imag} */,
  {32'h3fd33fe9, 32'h3ce466d0} /* (12, 4, 1) {real, imag} */,
  {32'hc022a435, 32'hbfa3dc1e} /* (12, 4, 0) {real, imag} */,
  {32'h404a734b, 32'hbf823454} /* (12, 3, 31) {real, imag} */,
  {32'hbfe19be8, 32'h3ee7a972} /* (12, 3, 30) {real, imag} */,
  {32'h3fb9425c, 32'hbf90bad8} /* (12, 3, 29) {real, imag} */,
  {32'hbfb1a083, 32'h4040b8a8} /* (12, 3, 28) {real, imag} */,
  {32'hbfadd8de, 32'hbf2ae5da} /* (12, 3, 27) {real, imag} */,
  {32'h3f81dd1e, 32'hbedcd278} /* (12, 3, 26) {real, imag} */,
  {32'hbee9a6c1, 32'hbf978a46} /* (12, 3, 25) {real, imag} */,
  {32'h3f40cdf3, 32'hbf03564f} /* (12, 3, 24) {real, imag} */,
  {32'h3e4225a4, 32'h3ee559da} /* (12, 3, 23) {real, imag} */,
  {32'h3f9423d2, 32'hbe7c1963} /* (12, 3, 22) {real, imag} */,
  {32'h40525502, 32'h4017bf80} /* (12, 3, 21) {real, imag} */,
  {32'h3f5a8c4d, 32'hbf6d0ac6} /* (12, 3, 20) {real, imag} */,
  {32'h3fba5958, 32'h3f1ac303} /* (12, 3, 19) {real, imag} */,
  {32'h3fd2c13f, 32'h3ea08ccb} /* (12, 3, 18) {real, imag} */,
  {32'hbf7dc35d, 32'h3fb9b6de} /* (12, 3, 17) {real, imag} */,
  {32'h3d92112d, 32'h3fc99ff7} /* (12, 3, 16) {real, imag} */,
  {32'h3ffc3e31, 32'h4029b8d6} /* (12, 3, 15) {real, imag} */,
  {32'hbfdb2a4d, 32'hbdd59ae7} /* (12, 3, 14) {real, imag} */,
  {32'h3e4ee5e9, 32'h3e152e94} /* (12, 3, 13) {real, imag} */,
  {32'hbe02e0d2, 32'hbee312ae} /* (12, 3, 12) {real, imag} */,
  {32'h403664d5, 32'hbcadfcb6} /* (12, 3, 11) {real, imag} */,
  {32'h3dc00796, 32'h3faac7be} /* (12, 3, 10) {real, imag} */,
  {32'hbd4b455a, 32'hc0384f3a} /* (12, 3, 9) {real, imag} */,
  {32'h3f9db46a, 32'h3e78340e} /* (12, 3, 8) {real, imag} */,
  {32'hbfb038de, 32'hbf981aa7} /* (12, 3, 7) {real, imag} */,
  {32'hbf1f20bc, 32'hc049b5e3} /* (12, 3, 6) {real, imag} */,
  {32'h3e81ca2d, 32'h400419c6} /* (12, 3, 5) {real, imag} */,
  {32'h3f2d2d22, 32'hbe57bbae} /* (12, 3, 4) {real, imag} */,
  {32'hc061cab9, 32'h3fec3c28} /* (12, 3, 3) {real, imag} */,
  {32'h402b599a, 32'hbf0c9970} /* (12, 3, 2) {real, imag} */,
  {32'hbf72485c, 32'hbfa9fd36} /* (12, 3, 1) {real, imag} */,
  {32'h3fc8f89a, 32'h3cdcd572} /* (12, 3, 0) {real, imag} */,
  {32'h3dac474e, 32'hc02c9139} /* (12, 2, 31) {real, imag} */,
  {32'hbf61fcec, 32'h3f7bd3ef} /* (12, 2, 30) {real, imag} */,
  {32'hbfcf12e3, 32'h3fe50ac9} /* (12, 2, 29) {real, imag} */,
  {32'h3fbfb0da, 32'hbf92548e} /* (12, 2, 28) {real, imag} */,
  {32'h40034cc7, 32'h3eb9a7d2} /* (12, 2, 27) {real, imag} */,
  {32'hc0874c12, 32'hbf822b0d} /* (12, 2, 26) {real, imag} */,
  {32'h3e8abad0, 32'hbf088b96} /* (12, 2, 25) {real, imag} */,
  {32'h3f76ec04, 32'h400df0a4} /* (12, 2, 24) {real, imag} */,
  {32'hbfff5adf, 32'hbe710394} /* (12, 2, 23) {real, imag} */,
  {32'hc00799a9, 32'hc00abb6d} /* (12, 2, 22) {real, imag} */,
  {32'h3eca87d9, 32'h40709cda} /* (12, 2, 21) {real, imag} */,
  {32'h3d8b3bf5, 32'hbfd84507} /* (12, 2, 20) {real, imag} */,
  {32'hbf7f723d, 32'hbf966ca6} /* (12, 2, 19) {real, imag} */,
  {32'hc00b70fe, 32'h4010620f} /* (12, 2, 18) {real, imag} */,
  {32'h401f878f, 32'h3f9510de} /* (12, 2, 17) {real, imag} */,
  {32'h3ea94a27, 32'hbe6f35e8} /* (12, 2, 16) {real, imag} */,
  {32'hbf228023, 32'hbf270d47} /* (12, 2, 15) {real, imag} */,
  {32'h3f713faf, 32'hc0408275} /* (12, 2, 14) {real, imag} */,
  {32'h3fb49cbd, 32'hbe9eb972} /* (12, 2, 13) {real, imag} */,
  {32'hc0347969, 32'h3fa65353} /* (12, 2, 12) {real, imag} */,
  {32'h3f2d9c3d, 32'hbf4be5bf} /* (12, 2, 11) {real, imag} */,
  {32'hbfc8fe2f, 32'hbfa60e4c} /* (12, 2, 10) {real, imag} */,
  {32'h3de329d9, 32'hc00ae267} /* (12, 2, 9) {real, imag} */,
  {32'hc0037745, 32'hc0419849} /* (12, 2, 8) {real, imag} */,
  {32'h3ef95b07, 32'hc07444ba} /* (12, 2, 7) {real, imag} */,
  {32'h403d5a6e, 32'h4014f162} /* (12, 2, 6) {real, imag} */,
  {32'hbf79b789, 32'h3f92019c} /* (12, 2, 5) {real, imag} */,
  {32'hbe4edb86, 32'hc014c007} /* (12, 2, 4) {real, imag} */,
  {32'h3f7ada9b, 32'hbfe4b5a6} /* (12, 2, 3) {real, imag} */,
  {32'hbf78a9c6, 32'h401e8d08} /* (12, 2, 2) {real, imag} */,
  {32'h3fce5582, 32'h4039435c} /* (12, 2, 1) {real, imag} */,
  {32'hbf424646, 32'h3f14e922} /* (12, 2, 0) {real, imag} */,
  {32'hbfab8a9f, 32'hbc382ecc} /* (12, 1, 31) {real, imag} */,
  {32'h402a2e88, 32'hbf175360} /* (12, 1, 30) {real, imag} */,
  {32'h3e9c6fa6, 32'h3d415fe3} /* (12, 1, 29) {real, imag} */,
  {32'hc05721c9, 32'h3fd63ebf} /* (12, 1, 28) {real, imag} */,
  {32'hc04352a0, 32'hbf3839c0} /* (12, 1, 27) {real, imag} */,
  {32'hbff79a61, 32'hbfa77511} /* (12, 1, 26) {real, imag} */,
  {32'h3f4e3952, 32'h3eec5c11} /* (12, 1, 25) {real, imag} */,
  {32'hbf65f51f, 32'h3fbe32a7} /* (12, 1, 24) {real, imag} */,
  {32'h3f499a36, 32'hbf1cb28c} /* (12, 1, 23) {real, imag} */,
  {32'hbf50bbd2, 32'h3ffe8608} /* (12, 1, 22) {real, imag} */,
  {32'h3f3c4f9c, 32'h3f70a06c} /* (12, 1, 21) {real, imag} */,
  {32'hc0022e3a, 32'hc00676a3} /* (12, 1, 20) {real, imag} */,
  {32'h3d8a8ca6, 32'hbfc86757} /* (12, 1, 19) {real, imag} */,
  {32'hbf4d1c74, 32'hbe984437} /* (12, 1, 18) {real, imag} */,
  {32'h3fabb085, 32'hbf02bdd9} /* (12, 1, 17) {real, imag} */,
  {32'h3fa9a920, 32'h3eccb87b} /* (12, 1, 16) {real, imag} */,
  {32'h3ec65d0e, 32'h3f5e8d3d} /* (12, 1, 15) {real, imag} */,
  {32'h3e10b2bf, 32'hbe795db6} /* (12, 1, 14) {real, imag} */,
  {32'h3fd84387, 32'hbf30dd3f} /* (12, 1, 13) {real, imag} */,
  {32'hbfe05357, 32'h3fc58625} /* (12, 1, 12) {real, imag} */,
  {32'h3fc50994, 32'hc00c6ed7} /* (12, 1, 11) {real, imag} */,
  {32'hbf327edf, 32'hbfc2277d} /* (12, 1, 10) {real, imag} */,
  {32'hbf9ed500, 32'h3f81ce74} /* (12, 1, 9) {real, imag} */,
  {32'h40302fff, 32'h3fc78066} /* (12, 1, 8) {real, imag} */,
  {32'hbf1a5f26, 32'h3fc5e4ac} /* (12, 1, 7) {real, imag} */,
  {32'hbe9b6a59, 32'h401a6eac} /* (12, 1, 6) {real, imag} */,
  {32'hbeb041a4, 32'h40281ea9} /* (12, 1, 5) {real, imag} */,
  {32'hc06959f4, 32'h3f2b9f14} /* (12, 1, 4) {real, imag} */,
  {32'h3fc8b5a5, 32'h3fb1eb00} /* (12, 1, 3) {real, imag} */,
  {32'h400d5587, 32'hbfcc1124} /* (12, 1, 2) {real, imag} */,
  {32'h3f88e6e3, 32'h3c7f6f40} /* (12, 1, 1) {real, imag} */,
  {32'h4008c1e6, 32'h3e0dbdf0} /* (12, 1, 0) {real, imag} */,
  {32'hbe8bf94f, 32'h3e16ccc1} /* (12, 0, 31) {real, imag} */,
  {32'hbffc9831, 32'hbf503040} /* (12, 0, 30) {real, imag} */,
  {32'h3ef90143, 32'hbeac0c34} /* (12, 0, 29) {real, imag} */,
  {32'h3c306939, 32'h3f97cb17} /* (12, 0, 28) {real, imag} */,
  {32'h404e8951, 32'hc07b4beb} /* (12, 0, 27) {real, imag} */,
  {32'h3fbfebcd, 32'hbfeafe26} /* (12, 0, 26) {real, imag} */,
  {32'hbe913aee, 32'h3fe87782} /* (12, 0, 25) {real, imag} */,
  {32'h406225d9, 32'h40027d4a} /* (12, 0, 24) {real, imag} */,
  {32'hbf8f6c2b, 32'h3fa3ec82} /* (12, 0, 23) {real, imag} */,
  {32'h3f8ef3e4, 32'hbe78263b} /* (12, 0, 22) {real, imag} */,
  {32'hc037ffef, 32'h3e1d6dbe} /* (12, 0, 21) {real, imag} */,
  {32'h3f0215d5, 32'hbfa7046b} /* (12, 0, 20) {real, imag} */,
  {32'h3f2a932c, 32'hc057eda3} /* (12, 0, 19) {real, imag} */,
  {32'h3de21874, 32'h4024b3b3} /* (12, 0, 18) {real, imag} */,
  {32'hbeeb5e17, 32'hbf269a52} /* (12, 0, 17) {real, imag} */,
  {32'hbe435355, 32'hbee851c1} /* (12, 0, 16) {real, imag} */,
  {32'h3eb858e2, 32'h3fe1bb52} /* (12, 0, 15) {real, imag} */,
  {32'h3fafb135, 32'hbf2da643} /* (12, 0, 14) {real, imag} */,
  {32'hbef7d602, 32'hbf833efe} /* (12, 0, 13) {real, imag} */,
  {32'hbff2f38e, 32'hbfebb336} /* (12, 0, 12) {real, imag} */,
  {32'h3f045e72, 32'hbfb5ac5e} /* (12, 0, 11) {real, imag} */,
  {32'h3f4d741b, 32'hc00667d6} /* (12, 0, 10) {real, imag} */,
  {32'h40528817, 32'hc0443fd5} /* (12, 0, 9) {real, imag} */,
  {32'h3fcb0c0a, 32'hbea4cb91} /* (12, 0, 8) {real, imag} */,
  {32'hbf1e5af9, 32'hbe4613f1} /* (12, 0, 7) {real, imag} */,
  {32'h4093aa2b, 32'h400bc0a3} /* (12, 0, 6) {real, imag} */,
  {32'hc0106c4f, 32'hbeca04a9} /* (12, 0, 5) {real, imag} */,
  {32'h3fad0d11, 32'hbf5f9cba} /* (12, 0, 4) {real, imag} */,
  {32'hc019341b, 32'h3ed24ddb} /* (12, 0, 3) {real, imag} */,
  {32'hbf80ea4a, 32'h4010e22c} /* (12, 0, 2) {real, imag} */,
  {32'h3ed627e2, 32'hbfd78dc6} /* (12, 0, 1) {real, imag} */,
  {32'hbfa13490, 32'hbfeb4004} /* (12, 0, 0) {real, imag} */,
  {32'h40a48cfd, 32'hc0babc42} /* (11, 31, 31) {real, imag} */,
  {32'hc0224b97, 32'h41112e0f} /* (11, 31, 30) {real, imag} */,
  {32'hbe3879a0, 32'h3faa4256} /* (11, 31, 29) {real, imag} */,
  {32'hc06d7c55, 32'hc086522e} /* (11, 31, 28) {real, imag} */,
  {32'hbf9bdb95, 32'hbf524e95} /* (11, 31, 27) {real, imag} */,
  {32'h3fff5d0f, 32'h3f605648} /* (11, 31, 26) {real, imag} */,
  {32'h40478fc3, 32'hc00295ad} /* (11, 31, 25) {real, imag} */,
  {32'h3fb2f58c, 32'h3f1f4fc9} /* (11, 31, 24) {real, imag} */,
  {32'hc0152c14, 32'hbfb848c1} /* (11, 31, 23) {real, imag} */,
  {32'hc02fa291, 32'h3ff3ec37} /* (11, 31, 22) {real, imag} */,
  {32'h3f1ac058, 32'h4051e020} /* (11, 31, 21) {real, imag} */,
  {32'hbd8f2125, 32'h3f05d54f} /* (11, 31, 20) {real, imag} */,
  {32'h4019a6a4, 32'h3f9c9810} /* (11, 31, 19) {real, imag} */,
  {32'hbefb475a, 32'h4043df99} /* (11, 31, 18) {real, imag} */,
  {32'h3f5b8332, 32'h3fe1e5d1} /* (11, 31, 17) {real, imag} */,
  {32'h3f1ebaee, 32'h3f3088d2} /* (11, 31, 16) {real, imag} */,
  {32'h3fceaf83, 32'hbfab20e7} /* (11, 31, 15) {real, imag} */,
  {32'hc02ad555, 32'h3d35ae47} /* (11, 31, 14) {real, imag} */,
  {32'h3f8aeb02, 32'hc01e6750} /* (11, 31, 13) {real, imag} */,
  {32'hc0225ee3, 32'h3f04801f} /* (11, 31, 12) {real, imag} */,
  {32'hc020162f, 32'hbfd3e53b} /* (11, 31, 11) {real, imag} */,
  {32'h3f94d4c4, 32'hc02cef25} /* (11, 31, 10) {real, imag} */,
  {32'h40346c75, 32'h403f3a4f} /* (11, 31, 9) {real, imag} */,
  {32'hbfe09173, 32'hbd2d9d22} /* (11, 31, 8) {real, imag} */,
  {32'h3f2a2d00, 32'hbfbe33af} /* (11, 31, 7) {real, imag} */,
  {32'h401ddf82, 32'h3fca6630} /* (11, 31, 6) {real, imag} */,
  {32'hbf267b66, 32'h4084381d} /* (11, 31, 5) {real, imag} */,
  {32'h3a089aef, 32'hc04ec705} /* (11, 31, 4) {real, imag} */,
  {32'h4001c368, 32'hc01509b6} /* (11, 31, 3) {real, imag} */,
  {32'h3fb0dd0e, 32'h40985605} /* (11, 31, 2) {real, imag} */,
  {32'h402ddff7, 32'hbf9d6480} /* (11, 31, 1) {real, imag} */,
  {32'h409c9c9d, 32'hc0fb8d1d} /* (11, 31, 0) {real, imag} */,
  {32'hc017d342, 32'h402f2403} /* (11, 30, 31) {real, imag} */,
  {32'h408cb9d4, 32'hbe767f08} /* (11, 30, 30) {real, imag} */,
  {32'hbfadb355, 32'hc014893c} /* (11, 30, 29) {real, imag} */,
  {32'h405c2168, 32'h3fe952fb} /* (11, 30, 28) {real, imag} */,
  {32'hbf8ca14a, 32'hbf81892f} /* (11, 30, 27) {real, imag} */,
  {32'h3f876722, 32'hc09ab441} /* (11, 30, 26) {real, imag} */,
  {32'h3f3875f0, 32'hbff3d1ad} /* (11, 30, 25) {real, imag} */,
  {32'h3fb713c1, 32'hbfd51014} /* (11, 30, 24) {real, imag} */,
  {32'h400011e6, 32'hbf531346} /* (11, 30, 23) {real, imag} */,
  {32'h4067aea7, 32'h3fd7793e} /* (11, 30, 22) {real, imag} */,
  {32'hbf015a47, 32'hc0143a9c} /* (11, 30, 21) {real, imag} */,
  {32'h3f3bef51, 32'hbf755526} /* (11, 30, 20) {real, imag} */,
  {32'h3f99dbcd, 32'h400d20bf} /* (11, 30, 19) {real, imag} */,
  {32'h3f8ab6ef, 32'hc00cb573} /* (11, 30, 18) {real, imag} */,
  {32'h3ffe40fe, 32'h3fc9ceaf} /* (11, 30, 17) {real, imag} */,
  {32'h3e396810, 32'h3f5f404f} /* (11, 30, 16) {real, imag} */,
  {32'h3dfc6892, 32'hbfc34112} /* (11, 30, 15) {real, imag} */,
  {32'h3e465f8f, 32'h3f19c5c5} /* (11, 30, 14) {real, imag} */,
  {32'h3fe9605b, 32'h3f17097e} /* (11, 30, 13) {real, imag} */,
  {32'hc07a3c42, 32'h3f40a828} /* (11, 30, 12) {real, imag} */,
  {32'hbf29312b, 32'hbfcc6859} /* (11, 30, 11) {real, imag} */,
  {32'h3e13c68c, 32'hbf60b813} /* (11, 30, 10) {real, imag} */,
  {32'hc008b163, 32'h3e664720} /* (11, 30, 9) {real, imag} */,
  {32'h3ff0e6cf, 32'hbf361612} /* (11, 30, 8) {real, imag} */,
  {32'h401ea008, 32'h3e98dcf5} /* (11, 30, 7) {real, imag} */,
  {32'hbfe53fd2, 32'h3eb2b38f} /* (11, 30, 6) {real, imag} */,
  {32'h3ca342ec, 32'hbf173b72} /* (11, 30, 5) {real, imag} */,
  {32'hbfd7a324, 32'hbfeba21c} /* (11, 30, 4) {real, imag} */,
  {32'hc0531f70, 32'h3f89e528} /* (11, 30, 3) {real, imag} */,
  {32'h40ce527a, 32'hc0570112} /* (11, 30, 2) {real, imag} */,
  {32'hc0e5e651, 32'h40385c2b} /* (11, 30, 1) {real, imag} */,
  {32'hbf9aa279, 32'h40821432} /* (11, 30, 0) {real, imag} */,
  {32'h3f23713e, 32'hc0663582} /* (11, 29, 31) {real, imag} */,
  {32'h4006b267, 32'h4082c047} /* (11, 29, 30) {real, imag} */,
  {32'hbf7c124b, 32'hbede4d2d} /* (11, 29, 29) {real, imag} */,
  {32'h3ea4c835, 32'hbff31295} /* (11, 29, 28) {real, imag} */,
  {32'h40505f52, 32'hc001d162} /* (11, 29, 27) {real, imag} */,
  {32'h3fa2e90c, 32'hbecc368e} /* (11, 29, 26) {real, imag} */,
  {32'hbe3bdabf, 32'h3fa4b883} /* (11, 29, 25) {real, imag} */,
  {32'hbf8762d6, 32'h403c14cc} /* (11, 29, 24) {real, imag} */,
  {32'hbe2c7502, 32'hbfcca917} /* (11, 29, 23) {real, imag} */,
  {32'h3fb56989, 32'h3d0cad65} /* (11, 29, 22) {real, imag} */,
  {32'hbfa51f87, 32'hbe92572b} /* (11, 29, 21) {real, imag} */,
  {32'hbfef3af6, 32'hc02160c9} /* (11, 29, 20) {real, imag} */,
  {32'h3f6191b7, 32'h3f7e3f42} /* (11, 29, 19) {real, imag} */,
  {32'h3f0204b1, 32'hbde6bd76} /* (11, 29, 18) {real, imag} */,
  {32'hbfdb0a9e, 32'hbfdb2446} /* (11, 29, 17) {real, imag} */,
  {32'h40099b8e, 32'hc0683d14} /* (11, 29, 16) {real, imag} */,
  {32'h3f60e435, 32'hbefd576f} /* (11, 29, 15) {real, imag} */,
  {32'hc01d6236, 32'h3ef5cca6} /* (11, 29, 14) {real, imag} */,
  {32'h40494c70, 32'hbf5409d6} /* (11, 29, 13) {real, imag} */,
  {32'h3ea1ee2a, 32'hbeb25c1d} /* (11, 29, 12) {real, imag} */,
  {32'hbf099d38, 32'hbf1c3599} /* (11, 29, 11) {real, imag} */,
  {32'h4053f38d, 32'h3e3b7bc2} /* (11, 29, 10) {real, imag} */,
  {32'hc03aff3b, 32'h3f1c1796} /* (11, 29, 9) {real, imag} */,
  {32'hbf9d3e5b, 32'h3f8899cd} /* (11, 29, 8) {real, imag} */,
  {32'h3efcc359, 32'h40801f8d} /* (11, 29, 7) {real, imag} */,
  {32'hbfade4da, 32'hbff2a325} /* (11, 29, 6) {real, imag} */,
  {32'h3fa85e94, 32'hbfbe2077} /* (11, 29, 5) {real, imag} */,
  {32'h3f00c68d, 32'hbf8740e5} /* (11, 29, 4) {real, imag} */,
  {32'h3f83957a, 32'h3f2a578b} /* (11, 29, 3) {real, imag} */,
  {32'hbf173548, 32'h40a27ce9} /* (11, 29, 2) {real, imag} */,
  {32'hbfa6026e, 32'hbfabbd61} /* (11, 29, 1) {real, imag} */,
  {32'h3f42c461, 32'h3fd6417d} /* (11, 29, 0) {real, imag} */,
  {32'h40251210, 32'h3e89a83f} /* (11, 28, 31) {real, imag} */,
  {32'h4080b98a, 32'hbfa2c832} /* (11, 28, 30) {real, imag} */,
  {32'hbf168378, 32'hc00dfd6e} /* (11, 28, 29) {real, imag} */,
  {32'hbf6e99b9, 32'hbf17f5ea} /* (11, 28, 28) {real, imag} */,
  {32'h3f179caf, 32'hbfe5291f} /* (11, 28, 27) {real, imag} */,
  {32'h40310f3c, 32'hbff3be31} /* (11, 28, 26) {real, imag} */,
  {32'hbea9d152, 32'hbebd99b6} /* (11, 28, 25) {real, imag} */,
  {32'hc02a1d49, 32'h4010fbe4} /* (11, 28, 24) {real, imag} */,
  {32'h3f74b8d5, 32'hbfc9bbe3} /* (11, 28, 23) {real, imag} */,
  {32'h3fdcb2db, 32'hc0149bb1} /* (11, 28, 22) {real, imag} */,
  {32'hbe219331, 32'hbece53c7} /* (11, 28, 21) {real, imag} */,
  {32'hbf7c08f7, 32'h3d3beb02} /* (11, 28, 20) {real, imag} */,
  {32'h3fc53a46, 32'hbe87f9be} /* (11, 28, 19) {real, imag} */,
  {32'h3e6c4241, 32'h4014ad45} /* (11, 28, 18) {real, imag} */,
  {32'hbfb336a1, 32'hbf6819f9} /* (11, 28, 17) {real, imag} */,
  {32'h3fc65444, 32'h401d21b7} /* (11, 28, 16) {real, imag} */,
  {32'hbdb639d4, 32'hbf1baa11} /* (11, 28, 15) {real, imag} */,
  {32'hbff51eac, 32'hbef3a6fb} /* (11, 28, 14) {real, imag} */,
  {32'hbff91a98, 32'h400dec83} /* (11, 28, 13) {real, imag} */,
  {32'h3f9c17eb, 32'hbcd9a37d} /* (11, 28, 12) {real, imag} */,
  {32'h3f952543, 32'hbf21c53a} /* (11, 28, 11) {real, imag} */,
  {32'hbf1b7678, 32'hbeaf19ad} /* (11, 28, 10) {real, imag} */,
  {32'hc0380ff5, 32'hbd9a7091} /* (11, 28, 9) {real, imag} */,
  {32'hc00916d9, 32'h3f40303d} /* (11, 28, 8) {real, imag} */,
  {32'h3f9393b5, 32'hc024a071} /* (11, 28, 7) {real, imag} */,
  {32'hbef32d36, 32'hbfb03a64} /* (11, 28, 6) {real, imag} */,
  {32'h3f47aa35, 32'h3f83aab5} /* (11, 28, 5) {real, imag} */,
  {32'hbe92b84b, 32'hbeb1e73a} /* (11, 28, 4) {real, imag} */,
  {32'h40215f82, 32'hc0c8eaad} /* (11, 28, 3) {real, imag} */,
  {32'hc038a00a, 32'h3fbab1a2} /* (11, 28, 2) {real, imag} */,
  {32'hbeaaae75, 32'h3f8c4df0} /* (11, 28, 1) {real, imag} */,
  {32'h3dd1aaa8, 32'hbce1bf18} /* (11, 28, 0) {real, imag} */,
  {32'hbf78dcca, 32'h405e1db4} /* (11, 27, 31) {real, imag} */,
  {32'hc0205958, 32'hbf8f8026} /* (11, 27, 30) {real, imag} */,
  {32'hbf833dcd, 32'hbfe8ff2d} /* (11, 27, 29) {real, imag} */,
  {32'h3f46c7bb, 32'hbb2d54c4} /* (11, 27, 28) {real, imag} */,
  {32'h409e58d0, 32'h3cc8abc0} /* (11, 27, 27) {real, imag} */,
  {32'hc009dd13, 32'h3f483e96} /* (11, 27, 26) {real, imag} */,
  {32'hbf721d35, 32'hc073ab55} /* (11, 27, 25) {real, imag} */,
  {32'h403c8678, 32'h400ba7ba} /* (11, 27, 24) {real, imag} */,
  {32'h3fc19e79, 32'h3f1c8a02} /* (11, 27, 23) {real, imag} */,
  {32'h3f12ed63, 32'hc02a7645} /* (11, 27, 22) {real, imag} */,
  {32'h3e22f85c, 32'h3fcf3278} /* (11, 27, 21) {real, imag} */,
  {32'hbf6fda95, 32'h3f8e8fd7} /* (11, 27, 20) {real, imag} */,
  {32'h3f0982a6, 32'hbf74a8dc} /* (11, 27, 19) {real, imag} */,
  {32'h3f07d474, 32'h3fa816ed} /* (11, 27, 18) {real, imag} */,
  {32'h4022bf37, 32'h4032b069} /* (11, 27, 17) {real, imag} */,
  {32'h3f8de73f, 32'h3e31052b} /* (11, 27, 16) {real, imag} */,
  {32'hbf81989c, 32'h3dc697ef} /* (11, 27, 15) {real, imag} */,
  {32'hbeb4563d, 32'hbd2ee610} /* (11, 27, 14) {real, imag} */,
  {32'h3fa7cc68, 32'hbf264d32} /* (11, 27, 13) {real, imag} */,
  {32'h3f896299, 32'hbe494646} /* (11, 27, 12) {real, imag} */,
  {32'hbf501f22, 32'h3f8e129c} /* (11, 27, 11) {real, imag} */,
  {32'hbfc8f11c, 32'hbfbef702} /* (11, 27, 10) {real, imag} */,
  {32'h3fb1239d, 32'h3efca579} /* (11, 27, 9) {real, imag} */,
  {32'h4010b269, 32'hbf726876} /* (11, 27, 8) {real, imag} */,
  {32'hbf81058c, 32'h400541ce} /* (11, 27, 7) {real, imag} */,
  {32'hbec2dffb, 32'h40388d54} /* (11, 27, 6) {real, imag} */,
  {32'hbf2d5ede, 32'hc02688e7} /* (11, 27, 5) {real, imag} */,
  {32'hbf9ae26f, 32'hbf88c8f0} /* (11, 27, 4) {real, imag} */,
  {32'h3ecaa699, 32'h3f27117f} /* (11, 27, 3) {real, imag} */,
  {32'h3f5bfd40, 32'hc0c81473} /* (11, 27, 2) {real, imag} */,
  {32'hbfa278ea, 32'h3e6ec5bf} /* (11, 27, 1) {real, imag} */,
  {32'hc00bf33f, 32'h407bab26} /* (11, 27, 0) {real, imag} */,
  {32'h3f13ffe0, 32'hc0115396} /* (11, 26, 31) {real, imag} */,
  {32'hc0424c84, 32'hc0814888} /* (11, 26, 30) {real, imag} */,
  {32'hbfc437fe, 32'h40212fd7} /* (11, 26, 29) {real, imag} */,
  {32'h401ea4b3, 32'h40183878} /* (11, 26, 28) {real, imag} */,
  {32'h3f7e8e95, 32'hbe032cc2} /* (11, 26, 27) {real, imag} */,
  {32'h3f8ba47b, 32'hbf3ad1c9} /* (11, 26, 26) {real, imag} */,
  {32'h401e4945, 32'hbff17769} /* (11, 26, 25) {real, imag} */,
  {32'hbf31d009, 32'h3f054ec7} /* (11, 26, 24) {real, imag} */,
  {32'hbed45004, 32'hbfcade5b} /* (11, 26, 23) {real, imag} */,
  {32'h3eb9e07c, 32'hbe89484b} /* (11, 26, 22) {real, imag} */,
  {32'h401fde3a, 32'h402834bb} /* (11, 26, 21) {real, imag} */,
  {32'hbfe9e36a, 32'h3f805d12} /* (11, 26, 20) {real, imag} */,
  {32'hbfb65090, 32'h3fa330b8} /* (11, 26, 19) {real, imag} */,
  {32'hbfd7acbd, 32'hc04459eb} /* (11, 26, 18) {real, imag} */,
  {32'h3fce4aec, 32'h3fb7972f} /* (11, 26, 17) {real, imag} */,
  {32'hbf83ed89, 32'h3f1abcc5} /* (11, 26, 16) {real, imag} */,
  {32'hc0105395, 32'hbdee13bd} /* (11, 26, 15) {real, imag} */,
  {32'h3f7266ca, 32'hc033b1f9} /* (11, 26, 14) {real, imag} */,
  {32'h3f974f0b, 32'h3fc6dc76} /* (11, 26, 13) {real, imag} */,
  {32'h3faa35f3, 32'hbf0d7a07} /* (11, 26, 12) {real, imag} */,
  {32'hbfa04c97, 32'h3f8d7eb7} /* (11, 26, 11) {real, imag} */,
  {32'hbe83a1d5, 32'h3ffe6399} /* (11, 26, 10) {real, imag} */,
  {32'h408e64c6, 32'h40170aae} /* (11, 26, 9) {real, imag} */,
  {32'h3fd04e4b, 32'hc0258abc} /* (11, 26, 8) {real, imag} */,
  {32'hbe8970be, 32'h3e48885a} /* (11, 26, 7) {real, imag} */,
  {32'h3ff3c7da, 32'hbf6f921f} /* (11, 26, 6) {real, imag} */,
  {32'hc01fdad9, 32'hbfe06dd5} /* (11, 26, 5) {real, imag} */,
  {32'hbf489226, 32'hbf8b891a} /* (11, 26, 4) {real, imag} */,
  {32'hbfc1f9f6, 32'h3f73f99b} /* (11, 26, 3) {real, imag} */,
  {32'hbf39d5e2, 32'hbfbfce76} /* (11, 26, 2) {real, imag} */,
  {32'hbf4ee889, 32'h3f83b6d5} /* (11, 26, 1) {real, imag} */,
  {32'h3fe89fa9, 32'h3ffe36d9} /* (11, 26, 0) {real, imag} */,
  {32'h3faee9a2, 32'h3eab8811} /* (11, 25, 31) {real, imag} */,
  {32'hbd57cdce, 32'hbf3d7d17} /* (11, 25, 30) {real, imag} */,
  {32'hbf7d5297, 32'h3fdb692b} /* (11, 25, 29) {real, imag} */,
  {32'hbe1911d6, 32'hbf1e1283} /* (11, 25, 28) {real, imag} */,
  {32'hbf69233d, 32'hbf95f1f6} /* (11, 25, 27) {real, imag} */,
  {32'hc019c08e, 32'h3f82fcc0} /* (11, 25, 26) {real, imag} */,
  {32'hbf801648, 32'h3f8c1dc2} /* (11, 25, 25) {real, imag} */,
  {32'h3f62445d, 32'h3fd50788} /* (11, 25, 24) {real, imag} */,
  {32'hbf88ca4b, 32'hbfd8de9a} /* (11, 25, 23) {real, imag} */,
  {32'hbf8dba55, 32'h3fcac671} /* (11, 25, 22) {real, imag} */,
  {32'hbe970d7a, 32'hbf664686} /* (11, 25, 21) {real, imag} */,
  {32'h3ff9f5e6, 32'hc0343801} /* (11, 25, 20) {real, imag} */,
  {32'h3fc4e97c, 32'h3e96f887} /* (11, 25, 19) {real, imag} */,
  {32'hc027e368, 32'hbfe8397b} /* (11, 25, 18) {real, imag} */,
  {32'h3fc48983, 32'h3fd0e187} /* (11, 25, 17) {real, imag} */,
  {32'h3c1b5c3e, 32'h3e2e4d97} /* (11, 25, 16) {real, imag} */,
  {32'hbfa87da8, 32'h405b0ad6} /* (11, 25, 15) {real, imag} */,
  {32'hbf542ffe, 32'h3e840576} /* (11, 25, 14) {real, imag} */,
  {32'hbe305aa2, 32'hbf285b46} /* (11, 25, 13) {real, imag} */,
  {32'hbc402298, 32'h40148868} /* (11, 25, 12) {real, imag} */,
  {32'h3e93e995, 32'h3f927bd0} /* (11, 25, 11) {real, imag} */,
  {32'h400b4ff4, 32'hc010af1f} /* (11, 25, 10) {real, imag} */,
  {32'hbfca6c59, 32'hbf6ff27d} /* (11, 25, 9) {real, imag} */,
  {32'h40093f74, 32'hbfa333b4} /* (11, 25, 8) {real, imag} */,
  {32'h3c77e64d, 32'h3fbaafa0} /* (11, 25, 7) {real, imag} */,
  {32'hbff55492, 32'hc0607e35} /* (11, 25, 6) {real, imag} */,
  {32'h3faa0a14, 32'hc050b501} /* (11, 25, 5) {real, imag} */,
  {32'h3fbc1b6f, 32'h3f7b4082} /* (11, 25, 4) {real, imag} */,
  {32'hbeb10af1, 32'h3f05de76} /* (11, 25, 3) {real, imag} */,
  {32'h3ebd8765, 32'hc00d4bd3} /* (11, 25, 2) {real, imag} */,
  {32'hbfcf234a, 32'h3e3ceaf1} /* (11, 25, 1) {real, imag} */,
  {32'h402da826, 32'h3f9d155c} /* (11, 25, 0) {real, imag} */,
  {32'hbf8a53dd, 32'hbe8b5795} /* (11, 24, 31) {real, imag} */,
  {32'hc0352fbf, 32'h3f8d7557} /* (11, 24, 30) {real, imag} */,
  {32'h3fed146a, 32'hbfe78c4c} /* (11, 24, 29) {real, imag} */,
  {32'h3ec1d27c, 32'h402607da} /* (11, 24, 28) {real, imag} */,
  {32'h4020c6ab, 32'hc005f7bf} /* (11, 24, 27) {real, imag} */,
  {32'hc01f6497, 32'hbe304998} /* (11, 24, 26) {real, imag} */,
  {32'hbfee4717, 32'hc04a005a} /* (11, 24, 25) {real, imag} */,
  {32'hc02e0f36, 32'hbf8d5f38} /* (11, 24, 24) {real, imag} */,
  {32'hbf291fbf, 32'h3f3b2c57} /* (11, 24, 23) {real, imag} */,
  {32'h3fe28a2e, 32'h3f79a4cd} /* (11, 24, 22) {real, imag} */,
  {32'hbf277434, 32'h3ec13ac8} /* (11, 24, 21) {real, imag} */,
  {32'hbfd5d893, 32'hbed85da3} /* (11, 24, 20) {real, imag} */,
  {32'h3f9d2f63, 32'hc034ca8a} /* (11, 24, 19) {real, imag} */,
  {32'hbfc7af11, 32'hbfa9ebf1} /* (11, 24, 18) {real, imag} */,
  {32'hbef6bbde, 32'hbea7f38c} /* (11, 24, 17) {real, imag} */,
  {32'h3ffbc800, 32'h400379a4} /* (11, 24, 16) {real, imag} */,
  {32'h3f7f651e, 32'hbeec671b} /* (11, 24, 15) {real, imag} */,
  {32'hbc72ff3e, 32'hbd7fead0} /* (11, 24, 14) {real, imag} */,
  {32'h400dd31e, 32'hbf264dc6} /* (11, 24, 13) {real, imag} */,
  {32'hbf16c34c, 32'hbfa015a9} /* (11, 24, 12) {real, imag} */,
  {32'hc0064ff7, 32'hbee5eed4} /* (11, 24, 11) {real, imag} */,
  {32'hbf8c29a8, 32'h401dccc4} /* (11, 24, 10) {real, imag} */,
  {32'hc071b6ce, 32'h3fcb1f17} /* (11, 24, 9) {real, imag} */,
  {32'h3f5c39d6, 32'hbfe60143} /* (11, 24, 8) {real, imag} */,
  {32'h3fea5f36, 32'h403b3f77} /* (11, 24, 7) {real, imag} */,
  {32'h4092ace4, 32'hbf299312} /* (11, 24, 6) {real, imag} */,
  {32'hbd9ec6ae, 32'h3f0ec493} /* (11, 24, 5) {real, imag} */,
  {32'h3feba00a, 32'hbf82c415} /* (11, 24, 4) {real, imag} */,
  {32'h3f293640, 32'hbdf639e2} /* (11, 24, 3) {real, imag} */,
  {32'h4039fa80, 32'h4015f877} /* (11, 24, 2) {real, imag} */,
  {32'hbfe77675, 32'h40313b07} /* (11, 24, 1) {real, imag} */,
  {32'hc028da7b, 32'h40781ce6} /* (11, 24, 0) {real, imag} */,
  {32'hbea189e9, 32'h3f3aa165} /* (11, 23, 31) {real, imag} */,
  {32'hc089a4a9, 32'h4038df42} /* (11, 23, 30) {real, imag} */,
  {32'h3ff9e434, 32'hbf50bcd7} /* (11, 23, 29) {real, imag} */,
  {32'hbfad79be, 32'hbf4c5cb3} /* (11, 23, 28) {real, imag} */,
  {32'hbfff847f, 32'hbf50157f} /* (11, 23, 27) {real, imag} */,
  {32'h4012de66, 32'hc00bb805} /* (11, 23, 26) {real, imag} */,
  {32'hc040e8cf, 32'h3fa6f180} /* (11, 23, 25) {real, imag} */,
  {32'h3fb1157f, 32'h3f9ada10} /* (11, 23, 24) {real, imag} */,
  {32'h3ff2ceaa, 32'hbf95ce5f} /* (11, 23, 23) {real, imag} */,
  {32'h40679e88, 32'hbfbaa108} /* (11, 23, 22) {real, imag} */,
  {32'hc00ed613, 32'h3fe2d323} /* (11, 23, 21) {real, imag} */,
  {32'h3f2fd20a, 32'h3eec2c46} /* (11, 23, 20) {real, imag} */,
  {32'hbff844ac, 32'hbf6b3a49} /* (11, 23, 19) {real, imag} */,
  {32'hc017b1c5, 32'h3e779884} /* (11, 23, 18) {real, imag} */,
  {32'h3f40eb31, 32'hbf27ee3d} /* (11, 23, 17) {real, imag} */,
  {32'h3f9fa886, 32'h3f8adfe5} /* (11, 23, 16) {real, imag} */,
  {32'hbfa0b9d1, 32'h3f8b70a6} /* (11, 23, 15) {real, imag} */,
  {32'h3ed69248, 32'h3e88f270} /* (11, 23, 14) {real, imag} */,
  {32'h3e8a601e, 32'h3edf405f} /* (11, 23, 13) {real, imag} */,
  {32'hbe487a3c, 32'hbf899311} /* (11, 23, 12) {real, imag} */,
  {32'h3f424f2f, 32'hc01499be} /* (11, 23, 11) {real, imag} */,
  {32'h3e9f364a, 32'h3fc54be8} /* (11, 23, 10) {real, imag} */,
  {32'h403251e5, 32'h3d8bfb28} /* (11, 23, 9) {real, imag} */,
  {32'h402aad4a, 32'h400ca745} /* (11, 23, 8) {real, imag} */,
  {32'h3f5bc071, 32'h3f9d0564} /* (11, 23, 7) {real, imag} */,
  {32'h3fb89bb5, 32'h3f76f4e5} /* (11, 23, 6) {real, imag} */,
  {32'hc007dfb1, 32'hc024a849} /* (11, 23, 5) {real, imag} */,
  {32'hbf1cd483, 32'hbf8cb578} /* (11, 23, 4) {real, imag} */,
  {32'hbf010d53, 32'h402ad08a} /* (11, 23, 3) {real, imag} */,
  {32'hbfd62560, 32'h3ed7b142} /* (11, 23, 2) {real, imag} */,
  {32'hbfc19b09, 32'h3f9a80ec} /* (11, 23, 1) {real, imag} */,
  {32'h3f5030f3, 32'hbf59839d} /* (11, 23, 0) {real, imag} */,
  {32'h3e037d99, 32'hc0508ad0} /* (11, 22, 31) {real, imag} */,
  {32'h3e67205a, 32'hbfa1b924} /* (11, 22, 30) {real, imag} */,
  {32'hbf3bc425, 32'h3f82b209} /* (11, 22, 29) {real, imag} */,
  {32'hc05d51f3, 32'h3f88c92e} /* (11, 22, 28) {real, imag} */,
  {32'h4016321d, 32'h400c3fe2} /* (11, 22, 27) {real, imag} */,
  {32'h400168e9, 32'h3fde995a} /* (11, 22, 26) {real, imag} */,
  {32'h40123e14, 32'h3e8b0d30} /* (11, 22, 25) {real, imag} */,
  {32'h406c8806, 32'h3ef488bf} /* (11, 22, 24) {real, imag} */,
  {32'hbf919346, 32'h40a6873f} /* (11, 22, 23) {real, imag} */,
  {32'hc011c1ed, 32'hbea6cf04} /* (11, 22, 22) {real, imag} */,
  {32'hbea4bb34, 32'hc0682d15} /* (11, 22, 21) {real, imag} */,
  {32'hbfd25fcf, 32'hbf515bc3} /* (11, 22, 20) {real, imag} */,
  {32'hbfc6462f, 32'h3f391e10} /* (11, 22, 19) {real, imag} */,
  {32'h40d7ca0c, 32'hc00cbd9c} /* (11, 22, 18) {real, imag} */,
  {32'hbf8f23ab, 32'h3c2d3de3} /* (11, 22, 17) {real, imag} */,
  {32'hbfd695ae, 32'hbe90e20d} /* (11, 22, 16) {real, imag} */,
  {32'hbdeadb31, 32'h40386358} /* (11, 22, 15) {real, imag} */,
  {32'hbfd1dadb, 32'h4079542e} /* (11, 22, 14) {real, imag} */,
  {32'h3bec1200, 32'h404707d4} /* (11, 22, 13) {real, imag} */,
  {32'hc01919cf, 32'hbd92ef76} /* (11, 22, 12) {real, imag} */,
  {32'h4051a0fe, 32'hbde223a4} /* (11, 22, 11) {real, imag} */,
  {32'h400fb9a2, 32'h3b4c04ca} /* (11, 22, 10) {real, imag} */,
  {32'hbfbd60a1, 32'hc0853799} /* (11, 22, 9) {real, imag} */,
  {32'h4025fe29, 32'h4018bd47} /* (11, 22, 8) {real, imag} */,
  {32'h3fc6ee77, 32'hbe224946} /* (11, 22, 7) {real, imag} */,
  {32'h4019d641, 32'h3fbc5da6} /* (11, 22, 6) {real, imag} */,
  {32'hc015b03d, 32'hbf6d8f64} /* (11, 22, 5) {real, imag} */,
  {32'hbf9ea46b, 32'hbde9000b} /* (11, 22, 4) {real, imag} */,
  {32'h3f54e69d, 32'hbd4e4934} /* (11, 22, 3) {real, imag} */,
  {32'hbe42963b, 32'hbedf0e8e} /* (11, 22, 2) {real, imag} */,
  {32'hbdc51524, 32'hbf1dd81e} /* (11, 22, 1) {real, imag} */,
  {32'h3e6ddb65, 32'h3f4af8b7} /* (11, 22, 0) {real, imag} */,
  {32'hbfede088, 32'h4072fd80} /* (11, 21, 31) {real, imag} */,
  {32'h3e8a59f4, 32'hbf335ea3} /* (11, 21, 30) {real, imag} */,
  {32'h3f90de44, 32'hc082a857} /* (11, 21, 29) {real, imag} */,
  {32'hc00fe600, 32'h3e00fc6d} /* (11, 21, 28) {real, imag} */,
  {32'hbf233742, 32'h3f5ca0ad} /* (11, 21, 27) {real, imag} */,
  {32'h4019be4d, 32'h3f6d2101} /* (11, 21, 26) {real, imag} */,
  {32'h3fda0558, 32'hc08c08d7} /* (11, 21, 25) {real, imag} */,
  {32'hc082256a, 32'hbfdc2df1} /* (11, 21, 24) {real, imag} */,
  {32'h3f52848a, 32'h4041d91b} /* (11, 21, 23) {real, imag} */,
  {32'h3c43e698, 32'h3f559711} /* (11, 21, 22) {real, imag} */,
  {32'h3f3ae74f, 32'h3cd4d463} /* (11, 21, 21) {real, imag} */,
  {32'h3ea04607, 32'h3f7f5c0d} /* (11, 21, 20) {real, imag} */,
  {32'h3f952d5f, 32'hbf80119b} /* (11, 21, 19) {real, imag} */,
  {32'h3f238cc9, 32'h40412045} /* (11, 21, 18) {real, imag} */,
  {32'hbfac4646, 32'hbe893628} /* (11, 21, 17) {real, imag} */,
  {32'hc03988b0, 32'h3f2bad5a} /* (11, 21, 16) {real, imag} */,
  {32'h3f91a4ee, 32'hbfaa22f9} /* (11, 21, 15) {real, imag} */,
  {32'hbf4b492c, 32'hbe8394ef} /* (11, 21, 14) {real, imag} */,
  {32'h3f98cfe1, 32'hbf8d67a8} /* (11, 21, 13) {real, imag} */,
  {32'hbf5cfb27, 32'h4055817a} /* (11, 21, 12) {real, imag} */,
  {32'hbfce288d, 32'hbf2a85cb} /* (11, 21, 11) {real, imag} */,
  {32'hbf9e8b02, 32'hbf89fa6c} /* (11, 21, 10) {real, imag} */,
  {32'h4001af55, 32'hbba7c68a} /* (11, 21, 9) {real, imag} */,
  {32'hbf599f70, 32'hbd9279fc} /* (11, 21, 8) {real, imag} */,
  {32'h4009cd1d, 32'hbd659cad} /* (11, 21, 7) {real, imag} */,
  {32'hbfe48e3d, 32'hbfcee5ef} /* (11, 21, 6) {real, imag} */,
  {32'h3f0fca19, 32'h3fd74209} /* (11, 21, 5) {real, imag} */,
  {32'h3fa51fad, 32'h3fe7fa96} /* (11, 21, 4) {real, imag} */,
  {32'hc032076d, 32'hbfacecee} /* (11, 21, 3) {real, imag} */,
  {32'h3fdb5ea8, 32'hbf4cac77} /* (11, 21, 2) {real, imag} */,
  {32'h3fdd0e7f, 32'h40211964} /* (11, 21, 1) {real, imag} */,
  {32'hc05451b4, 32'h3dd798fc} /* (11, 21, 0) {real, imag} */,
  {32'h3de8f94c, 32'h3ed8affa} /* (11, 20, 31) {real, imag} */,
  {32'h3faf6842, 32'h3ea717d5} /* (11, 20, 30) {real, imag} */,
  {32'hbddc7645, 32'h3fa1ee35} /* (11, 20, 29) {real, imag} */,
  {32'hbfa3adac, 32'hbf3c18d8} /* (11, 20, 28) {real, imag} */,
  {32'h401749b4, 32'hbf4d1069} /* (11, 20, 27) {real, imag} */,
  {32'hc04b56ff, 32'hbfb37cd2} /* (11, 20, 26) {real, imag} */,
  {32'h3eebeb70, 32'h3ee2327e} /* (11, 20, 25) {real, imag} */,
  {32'h3f06a0b3, 32'h3ff006fe} /* (11, 20, 24) {real, imag} */,
  {32'hc0796a4d, 32'hbf8ee1e7} /* (11, 20, 23) {real, imag} */,
  {32'hc0920035, 32'h401ddb73} /* (11, 20, 22) {real, imag} */,
  {32'h3fb7b7ec, 32'h3e7aced1} /* (11, 20, 21) {real, imag} */,
  {32'hbf9b9a82, 32'hc03e0a63} /* (11, 20, 20) {real, imag} */,
  {32'h401a9545, 32'h3fba1465} /* (11, 20, 19) {real, imag} */,
  {32'hbff2f56e, 32'h3e39efd0} /* (11, 20, 18) {real, imag} */,
  {32'h3f922667, 32'h3fc6d972} /* (11, 20, 17) {real, imag} */,
  {32'hbfbb8585, 32'hbf6aa5f0} /* (11, 20, 16) {real, imag} */,
  {32'hbfd33ba7, 32'hc00d1e7c} /* (11, 20, 15) {real, imag} */,
  {32'h402dbf7a, 32'hc0232a07} /* (11, 20, 14) {real, imag} */,
  {32'h3fc08735, 32'hc03bd07a} /* (11, 20, 13) {real, imag} */,
  {32'h40175c1e, 32'hc003963d} /* (11, 20, 12) {real, imag} */,
  {32'hbfaf077a, 32'hbf050232} /* (11, 20, 11) {real, imag} */,
  {32'hbf6b6393, 32'h40a5c8a5} /* (11, 20, 10) {real, imag} */,
  {32'hbd0d1265, 32'h3f4ac2de} /* (11, 20, 9) {real, imag} */,
  {32'hc00e0bb7, 32'h3fbe3eca} /* (11, 20, 8) {real, imag} */,
  {32'h3fb4e413, 32'hbff927c1} /* (11, 20, 7) {real, imag} */,
  {32'h3f1705d8, 32'h3f8dd5c5} /* (11, 20, 6) {real, imag} */,
  {32'hbf9d017e, 32'h404b14ce} /* (11, 20, 5) {real, imag} */,
  {32'hbdccf729, 32'h3f4d46a2} /* (11, 20, 4) {real, imag} */,
  {32'h401c666a, 32'hbe18105e} /* (11, 20, 3) {real, imag} */,
  {32'hbfa329b7, 32'h3f9e6d31} /* (11, 20, 2) {real, imag} */,
  {32'hbef7271a, 32'hbf9c0bf0} /* (11, 20, 1) {real, imag} */,
  {32'hc007e07f, 32'hbfbdb675} /* (11, 20, 0) {real, imag} */,
  {32'h40361a10, 32'hbfdc8ab8} /* (11, 19, 31) {real, imag} */,
  {32'h3fe925e8, 32'h3e647b7f} /* (11, 19, 30) {real, imag} */,
  {32'h4008cd23, 32'h402bc49e} /* (11, 19, 29) {real, imag} */,
  {32'h404fc5fb, 32'hbfe31ff4} /* (11, 19, 28) {real, imag} */,
  {32'h3f69923f, 32'hbfe8f297} /* (11, 19, 27) {real, imag} */,
  {32'hbf5fd561, 32'h4055f229} /* (11, 19, 26) {real, imag} */,
  {32'hb9ebebf3, 32'hbfadb042} /* (11, 19, 25) {real, imag} */,
  {32'h3fb7f9a9, 32'hbf21dfc9} /* (11, 19, 24) {real, imag} */,
  {32'hc0909243, 32'h3fd73ba9} /* (11, 19, 23) {real, imag} */,
  {32'h3f541ca5, 32'h403b55ff} /* (11, 19, 22) {real, imag} */,
  {32'hc0786e46, 32'hbfad36bc} /* (11, 19, 21) {real, imag} */,
  {32'hbd61f916, 32'h403774d1} /* (11, 19, 20) {real, imag} */,
  {32'h3ea940ae, 32'hbeb9fe44} /* (11, 19, 19) {real, imag} */,
  {32'h3fc27f5a, 32'h3f0e149f} /* (11, 19, 18) {real, imag} */,
  {32'hbf201932, 32'hc02adee0} /* (11, 19, 17) {real, imag} */,
  {32'h3ea521dc, 32'hbfde8fa9} /* (11, 19, 16) {real, imag} */,
  {32'h4005a8e9, 32'hbfa91469} /* (11, 19, 15) {real, imag} */,
  {32'hc0053662, 32'hbee2d883} /* (11, 19, 14) {real, imag} */,
  {32'h3ef7abe2, 32'hbfc24426} /* (11, 19, 13) {real, imag} */,
  {32'hbcb670a4, 32'h3f0bbcd9} /* (11, 19, 12) {real, imag} */,
  {32'hbf7cdf05, 32'h3e90d767} /* (11, 19, 11) {real, imag} */,
  {32'hbf659b07, 32'hbf9b9983} /* (11, 19, 10) {real, imag} */,
  {32'h404fc16d, 32'hc0039138} /* (11, 19, 9) {real, imag} */,
  {32'hbf04f19e, 32'hbfbe28b5} /* (11, 19, 8) {real, imag} */,
  {32'hbf72a1c6, 32'h4022ad7e} /* (11, 19, 7) {real, imag} */,
  {32'h3fa95e3d, 32'h3fcf1a00} /* (11, 19, 6) {real, imag} */,
  {32'h3e8f61ea, 32'h3fba80fc} /* (11, 19, 5) {real, imag} */,
  {32'h3f722936, 32'h3f755e9c} /* (11, 19, 4) {real, imag} */,
  {32'hbedea681, 32'hbfe721d6} /* (11, 19, 3) {real, imag} */,
  {32'hbcea39a2, 32'hbf509738} /* (11, 19, 2) {real, imag} */,
  {32'hbf5ed44d, 32'hbf056ac8} /* (11, 19, 1) {real, imag} */,
  {32'hbd9e6f6f, 32'hbf6db5ef} /* (11, 19, 0) {real, imag} */,
  {32'h3fa14081, 32'h3fee188e} /* (11, 18, 31) {real, imag} */,
  {32'h3ff5ba49, 32'h402f7018} /* (11, 18, 30) {real, imag} */,
  {32'hbeefb87e, 32'hbf0b0a65} /* (11, 18, 29) {real, imag} */,
  {32'h3e6af56a, 32'hbf3b216c} /* (11, 18, 28) {real, imag} */,
  {32'hbf8c399f, 32'h3fe8b884} /* (11, 18, 27) {real, imag} */,
  {32'h3dd4d6d9, 32'hbf6d03e4} /* (11, 18, 26) {real, imag} */,
  {32'h400c07ce, 32'hbe879bd9} /* (11, 18, 25) {real, imag} */,
  {32'hbffe0675, 32'h3f896687} /* (11, 18, 24) {real, imag} */,
  {32'h3df4b129, 32'h406a31e8} /* (11, 18, 23) {real, imag} */,
  {32'h3f604be6, 32'h40580caa} /* (11, 18, 22) {real, imag} */,
  {32'hbf9fa6c1, 32'hbe84fd47} /* (11, 18, 21) {real, imag} */,
  {32'hbfd3ac4e, 32'hbf35ac5c} /* (11, 18, 20) {real, imag} */,
  {32'h3f93eedf, 32'h403797e0} /* (11, 18, 19) {real, imag} */,
  {32'h3f69a875, 32'h40232c3a} /* (11, 18, 18) {real, imag} */,
  {32'hbe35e345, 32'h3e99e265} /* (11, 18, 17) {real, imag} */,
  {32'h401ab647, 32'hbf45ca7d} /* (11, 18, 16) {real, imag} */,
  {32'h4005d873, 32'h400bca01} /* (11, 18, 15) {real, imag} */,
  {32'h406895cf, 32'h3ee41431} /* (11, 18, 14) {real, imag} */,
  {32'hbfbd5ccf, 32'hbf65a586} /* (11, 18, 13) {real, imag} */,
  {32'h3fe988f5, 32'hc0223ddb} /* (11, 18, 12) {real, imag} */,
  {32'hbedcea16, 32'h406094eb} /* (11, 18, 11) {real, imag} */,
  {32'h3ecf63b7, 32'h3feea4ea} /* (11, 18, 10) {real, imag} */,
  {32'h4032844e, 32'hbfd4d877} /* (11, 18, 9) {real, imag} */,
  {32'h3f5894b3, 32'hbf875ac3} /* (11, 18, 8) {real, imag} */,
  {32'hbf754a9a, 32'hbfb36279} /* (11, 18, 7) {real, imag} */,
  {32'hbf585c2d, 32'h3d4145e2} /* (11, 18, 6) {real, imag} */,
  {32'hbfd6bef4, 32'h3e07d195} /* (11, 18, 5) {real, imag} */,
  {32'h3de2f9b4, 32'h3ee6cb95} /* (11, 18, 4) {real, imag} */,
  {32'h3ea9cad5, 32'hbff005c0} /* (11, 18, 3) {real, imag} */,
  {32'hbe891f0e, 32'h3f5f3577} /* (11, 18, 2) {real, imag} */,
  {32'h3f2e5186, 32'hbe61ce19} /* (11, 18, 1) {real, imag} */,
  {32'h3f9ba926, 32'hbe9ecfd7} /* (11, 18, 0) {real, imag} */,
  {32'h3f8751f7, 32'hbef0c56d} /* (11, 17, 31) {real, imag} */,
  {32'h3f8fb071, 32'h3f3f3881} /* (11, 17, 30) {real, imag} */,
  {32'hbe50bf7b, 32'h402e992f} /* (11, 17, 29) {real, imag} */,
  {32'hbe1cd454, 32'hbfa206b1} /* (11, 17, 28) {real, imag} */,
  {32'hbf9a243a, 32'hbf4e6674} /* (11, 17, 27) {real, imag} */,
  {32'h3eaa4c75, 32'hbf86789c} /* (11, 17, 26) {real, imag} */,
  {32'h3f5b8e18, 32'h3fa9cf24} /* (11, 17, 25) {real, imag} */,
  {32'hbff54931, 32'h3eacce54} /* (11, 17, 24) {real, imag} */,
  {32'hbf951a84, 32'hbff40730} /* (11, 17, 23) {real, imag} */,
  {32'h3f2b951f, 32'hbc3f7b20} /* (11, 17, 22) {real, imag} */,
  {32'hc02b0e64, 32'hc06de636} /* (11, 17, 21) {real, imag} */,
  {32'hbef82465, 32'hbf7ac534} /* (11, 17, 20) {real, imag} */,
  {32'h3d613245, 32'hbe5bd4d9} /* (11, 17, 19) {real, imag} */,
  {32'h3fb65747, 32'h3dbf90bb} /* (11, 17, 18) {real, imag} */,
  {32'hbff3e997, 32'hbdce3df3} /* (11, 17, 17) {real, imag} */,
  {32'hbfb5c8c1, 32'h3fc88451} /* (11, 17, 16) {real, imag} */,
  {32'hbff262fd, 32'h3f46d9ed} /* (11, 17, 15) {real, imag} */,
  {32'h3e406efe, 32'h3fa6f738} /* (11, 17, 14) {real, imag} */,
  {32'hc028aada, 32'hbf8f113c} /* (11, 17, 13) {real, imag} */,
  {32'h3e5550c3, 32'h3fb2df6c} /* (11, 17, 12) {real, imag} */,
  {32'hc00ecb50, 32'h4021d7fa} /* (11, 17, 11) {real, imag} */,
  {32'h3f04260e, 32'hbf67fd93} /* (11, 17, 10) {real, imag} */,
  {32'hbff6992e, 32'hbfc0f88d} /* (11, 17, 9) {real, imag} */,
  {32'hbd8de0ac, 32'h3e86b1b5} /* (11, 17, 8) {real, imag} */,
  {32'hc025e906, 32'hbecb032e} /* (11, 17, 7) {real, imag} */,
  {32'hbfefbc2c, 32'h3fd9e60d} /* (11, 17, 6) {real, imag} */,
  {32'h3f93d410, 32'hbf8a6b85} /* (11, 17, 5) {real, imag} */,
  {32'h3e6c8c2e, 32'hbf8bdb90} /* (11, 17, 4) {real, imag} */,
  {32'h3f51abe4, 32'hbfa3463a} /* (11, 17, 3) {real, imag} */,
  {32'h408a33fb, 32'h3e764095} /* (11, 17, 2) {real, imag} */,
  {32'hbf80985e, 32'h3db739f2} /* (11, 17, 1) {real, imag} */,
  {32'hbf2fd553, 32'hbf8ae94e} /* (11, 17, 0) {real, imag} */,
  {32'hbda28af3, 32'h3f44160d} /* (11, 16, 31) {real, imag} */,
  {32'hbd22a7b8, 32'h3dba06b4} /* (11, 16, 30) {real, imag} */,
  {32'hbf4e9d25, 32'hbef05a6e} /* (11, 16, 29) {real, imag} */,
  {32'hbf590ea9, 32'h3de99a01} /* (11, 16, 28) {real, imag} */,
  {32'h3d330c01, 32'h40062225} /* (11, 16, 27) {real, imag} */,
  {32'hbf9215d0, 32'hbf47f623} /* (11, 16, 26) {real, imag} */,
  {32'hbeed29e2, 32'h3e7604cf} /* (11, 16, 25) {real, imag} */,
  {32'h3f965d9a, 32'hbf12eec1} /* (11, 16, 24) {real, imag} */,
  {32'h408a8007, 32'h3ef721a4} /* (11, 16, 23) {real, imag} */,
  {32'hbed09cf9, 32'h3ede6055} /* (11, 16, 22) {real, imag} */,
  {32'hbf8b0ec5, 32'h3fed9f24} /* (11, 16, 21) {real, imag} */,
  {32'hbf9d8f2b, 32'hbf901518} /* (11, 16, 20) {real, imag} */,
  {32'hbf8af5e9, 32'h3f993f2d} /* (11, 16, 19) {real, imag} */,
  {32'h3f038e8d, 32'h3ef68f3b} /* (11, 16, 18) {real, imag} */,
  {32'h3f9c52cd, 32'hbe1dc05d} /* (11, 16, 17) {real, imag} */,
  {32'h3ed1fee4, 32'h3da47fe8} /* (11, 16, 16) {real, imag} */,
  {32'hbf70c087, 32'hbf9f13fc} /* (11, 16, 15) {real, imag} */,
  {32'h3cebd6e3, 32'hbec80168} /* (11, 16, 14) {real, imag} */,
  {32'h4038fab3, 32'hbf86f750} /* (11, 16, 13) {real, imag} */,
  {32'h3f26b087, 32'h3fa4ea3c} /* (11, 16, 12) {real, imag} */,
  {32'h3f507182, 32'hbfcc6e45} /* (11, 16, 11) {real, imag} */,
  {32'hbf3eb191, 32'hbf7f54e8} /* (11, 16, 10) {real, imag} */,
  {32'hbd427509, 32'hc03c4802} /* (11, 16, 9) {real, imag} */,
  {32'h3f8ae2be, 32'hbff10e60} /* (11, 16, 8) {real, imag} */,
  {32'h3fa0a7f5, 32'hc0111045} /* (11, 16, 7) {real, imag} */,
  {32'h3e25e021, 32'h3fc8d1d6} /* (11, 16, 6) {real, imag} */,
  {32'hbfc45bd9, 32'h3f1e2642} /* (11, 16, 5) {real, imag} */,
  {32'h3f6241c5, 32'hbdd33b76} /* (11, 16, 4) {real, imag} */,
  {32'h3f9d3176, 32'hbdc30b37} /* (11, 16, 3) {real, imag} */,
  {32'h3eee991c, 32'h3f5973d2} /* (11, 16, 2) {real, imag} */,
  {32'hbf2cbdb0, 32'hbf1ff262} /* (11, 16, 1) {real, imag} */,
  {32'h3ff417fc, 32'h3ecbf637} /* (11, 16, 0) {real, imag} */,
  {32'h3fdf9015, 32'hbf6e6a00} /* (11, 15, 31) {real, imag} */,
  {32'hbfac40cf, 32'h3e695ff6} /* (11, 15, 30) {real, imag} */,
  {32'hbfa793e7, 32'h3f9b3b06} /* (11, 15, 29) {real, imag} */,
  {32'hbebd155b, 32'hbdf2455a} /* (11, 15, 28) {real, imag} */,
  {32'hbe97dd9b, 32'h4005605f} /* (11, 15, 27) {real, imag} */,
  {32'h3e0b101b, 32'hbf0e77a5} /* (11, 15, 26) {real, imag} */,
  {32'h3ed6efd4, 32'hbf339d59} /* (11, 15, 25) {real, imag} */,
  {32'hc0423654, 32'h401146c2} /* (11, 15, 24) {real, imag} */,
  {32'hbfb44c35, 32'hbefa7885} /* (11, 15, 23) {real, imag} */,
  {32'h3e85ffad, 32'h3f26d2b7} /* (11, 15, 22) {real, imag} */,
  {32'h3fd8e01e, 32'h40080fbd} /* (11, 15, 21) {real, imag} */,
  {32'hbfbe72de, 32'hbf769fba} /* (11, 15, 20) {real, imag} */,
  {32'h3f1aa5de, 32'hc01aafb7} /* (11, 15, 19) {real, imag} */,
  {32'h3f074e39, 32'hbff48117} /* (11, 15, 18) {real, imag} */,
  {32'h3dd7a7e7, 32'hbef75ce6} /* (11, 15, 17) {real, imag} */,
  {32'hbfb9c564, 32'h3f085960} /* (11, 15, 16) {real, imag} */,
  {32'hbf6a1370, 32'hbecba7e8} /* (11, 15, 15) {real, imag} */,
  {32'h3ecb01ac, 32'h3f739c94} /* (11, 15, 14) {real, imag} */,
  {32'hc02934b5, 32'hbf19289d} /* (11, 15, 13) {real, imag} */,
  {32'h3f2ba702, 32'hbec76247} /* (11, 15, 12) {real, imag} */,
  {32'h4038899b, 32'hc037a75d} /* (11, 15, 11) {real, imag} */,
  {32'h3f81478b, 32'hbf869a87} /* (11, 15, 10) {real, imag} */,
  {32'hbf879099, 32'h3e0476ed} /* (11, 15, 9) {real, imag} */,
  {32'hbe0ba70c, 32'h3fec050c} /* (11, 15, 8) {real, imag} */,
  {32'h3f83afa5, 32'hbf5a5759} /* (11, 15, 7) {real, imag} */,
  {32'hbf5293d7, 32'h3fa47fbb} /* (11, 15, 6) {real, imag} */,
  {32'h3fc14131, 32'h3f9df864} /* (11, 15, 5) {real, imag} */,
  {32'h3e85f17e, 32'hbfd8735d} /* (11, 15, 4) {real, imag} */,
  {32'hbd08861f, 32'h3fe8ee6d} /* (11, 15, 3) {real, imag} */,
  {32'h3e2cf09b, 32'hbccbbb12} /* (11, 15, 2) {real, imag} */,
  {32'h3f6a26c8, 32'h3f36886b} /* (11, 15, 1) {real, imag} */,
  {32'h3f4180e1, 32'hbe0b031a} /* (11, 15, 0) {real, imag} */,
  {32'hbe5b2e85, 32'hbfee0be7} /* (11, 14, 31) {real, imag} */,
  {32'hbfa4a4b6, 32'h3fadd63e} /* (11, 14, 30) {real, imag} */,
  {32'h3f6b8ffb, 32'hbfe6232f} /* (11, 14, 29) {real, imag} */,
  {32'hbf5a6aa6, 32'h3f74bd3e} /* (11, 14, 28) {real, imag} */,
  {32'h3eed0bdc, 32'hbd197b12} /* (11, 14, 27) {real, imag} */,
  {32'hbf5a5cdb, 32'h3e20b4c7} /* (11, 14, 26) {real, imag} */,
  {32'hbd6dfbd0, 32'h3de8ab52} /* (11, 14, 25) {real, imag} */,
  {32'hbfd53c65, 32'hc021b1db} /* (11, 14, 24) {real, imag} */,
  {32'h3ff96ca6, 32'h3f9a19f7} /* (11, 14, 23) {real, imag} */,
  {32'hc0914c44, 32'h3de65791} /* (11, 14, 22) {real, imag} */,
  {32'hbe290387, 32'h3e4d06b4} /* (11, 14, 21) {real, imag} */,
  {32'hbe7cb05f, 32'hbdc2f9a1} /* (11, 14, 20) {real, imag} */,
  {32'h3f9dec76, 32'hbfdd4322} /* (11, 14, 19) {real, imag} */,
  {32'h405095d3, 32'h3fdac6ef} /* (11, 14, 18) {real, imag} */,
  {32'h3efdc52b, 32'h3f559def} /* (11, 14, 17) {real, imag} */,
  {32'h40062259, 32'hc035ab7e} /* (11, 14, 16) {real, imag} */,
  {32'hbf7c3d50, 32'h3f98f5be} /* (11, 14, 15) {real, imag} */,
  {32'h3f482d1b, 32'hbf555a70} /* (11, 14, 14) {real, imag} */,
  {32'h40107f40, 32'h3f8c8bda} /* (11, 14, 13) {real, imag} */,
  {32'h3e3f1539, 32'hbf8cc537} /* (11, 14, 12) {real, imag} */,
  {32'hbe4b932c, 32'h4007b41e} /* (11, 14, 11) {real, imag} */,
  {32'hbfb489fa, 32'h3ea8867e} /* (11, 14, 10) {real, imag} */,
  {32'hbf6afd8e, 32'hbeec0126} /* (11, 14, 9) {real, imag} */,
  {32'h3e147c1c, 32'hbf56d275} /* (11, 14, 8) {real, imag} */,
  {32'hbfcc91b5, 32'hbe792c11} /* (11, 14, 7) {real, imag} */,
  {32'hbd072152, 32'hbf597190} /* (11, 14, 6) {real, imag} */,
  {32'h3e3d7d6d, 32'h400f49e9} /* (11, 14, 5) {real, imag} */,
  {32'h3dec5466, 32'hbea1f45a} /* (11, 14, 4) {real, imag} */,
  {32'h3e0f7cf0, 32'hbfcbac0f} /* (11, 14, 3) {real, imag} */,
  {32'h3f8ad87e, 32'h3ed13814} /* (11, 14, 2) {real, imag} */,
  {32'hbfdbaaf2, 32'h401a1f97} /* (11, 14, 1) {real, imag} */,
  {32'hbeec714b, 32'hbfe007ad} /* (11, 14, 0) {real, imag} */,
  {32'h3f5700f0, 32'hbfc52460} /* (11, 13, 31) {real, imag} */,
  {32'h3f3adde9, 32'h400e84c0} /* (11, 13, 30) {real, imag} */,
  {32'h3f28789d, 32'h3fd74b47} /* (11, 13, 29) {real, imag} */,
  {32'hbf0d2e7d, 32'hbd3d19a4} /* (11, 13, 28) {real, imag} */,
  {32'hbf95621c, 32'h3fc7b2b2} /* (11, 13, 27) {real, imag} */,
  {32'h3fa020e1, 32'h3f012953} /* (11, 13, 26) {real, imag} */,
  {32'h4025bcc5, 32'hbf84ac4d} /* (11, 13, 25) {real, imag} */,
  {32'h3f282fb8, 32'h3e3f43c3} /* (11, 13, 24) {real, imag} */,
  {32'h402e75ab, 32'h40024a31} /* (11, 13, 23) {real, imag} */,
  {32'h40008981, 32'hc0484377} /* (11, 13, 22) {real, imag} */,
  {32'hbe05366e, 32'hbed3608b} /* (11, 13, 21) {real, imag} */,
  {32'h3f794910, 32'h400ac292} /* (11, 13, 20) {real, imag} */,
  {32'hbf13554d, 32'hbfc077d3} /* (11, 13, 19) {real, imag} */,
  {32'h3d156ef7, 32'h4057c6fd} /* (11, 13, 18) {real, imag} */,
  {32'hbfe52b87, 32'h3ef296b2} /* (11, 13, 17) {real, imag} */,
  {32'hbf49c893, 32'hbf30cc1f} /* (11, 13, 16) {real, imag} */,
  {32'hbf55dc86, 32'hbf968568} /* (11, 13, 15) {real, imag} */,
  {32'h3f2cc80f, 32'hbf312d81} /* (11, 13, 14) {real, imag} */,
  {32'hbebe8561, 32'hbfc42530} /* (11, 13, 13) {real, imag} */,
  {32'h3fbb5c65, 32'hbfb0b2ed} /* (11, 13, 12) {real, imag} */,
  {32'h3fa4fde9, 32'hc020a02a} /* (11, 13, 11) {real, imag} */,
  {32'h3f09376d, 32'h3f540168} /* (11, 13, 10) {real, imag} */,
  {32'hbf49af94, 32'hbfe1b5e7} /* (11, 13, 9) {real, imag} */,
  {32'h3fba3564, 32'hbf4655e0} /* (11, 13, 8) {real, imag} */,
  {32'hbe43d348, 32'h3f19ddae} /* (11, 13, 7) {real, imag} */,
  {32'h3ff5350c, 32'h3d17fdc0} /* (11, 13, 6) {real, imag} */,
  {32'h3ebf280a, 32'hc0181ddc} /* (11, 13, 5) {real, imag} */,
  {32'h3f8928ba, 32'h3f840c4e} /* (11, 13, 4) {real, imag} */,
  {32'hc0004306, 32'hbe31e30f} /* (11, 13, 3) {real, imag} */,
  {32'hbf55d0ef, 32'h3fbd31e3} /* (11, 13, 2) {real, imag} */,
  {32'hbf825772, 32'h3eb837a7} /* (11, 13, 1) {real, imag} */,
  {32'h3fee56d4, 32'h3f8fe7b6} /* (11, 13, 0) {real, imag} */,
  {32'h3fc64aa1, 32'h40085727} /* (11, 12, 31) {real, imag} */,
  {32'hc0316679, 32'hbe65f308} /* (11, 12, 30) {real, imag} */,
  {32'hbd0d7db0, 32'h3e25b892} /* (11, 12, 29) {real, imag} */,
  {32'h3fdc02a4, 32'h3ebf34b8} /* (11, 12, 28) {real, imag} */,
  {32'h3fafa3d5, 32'hbfb5aa56} /* (11, 12, 27) {real, imag} */,
  {32'hc0008776, 32'h4050f2bb} /* (11, 12, 26) {real, imag} */,
  {32'hbfece681, 32'h3fd5c6be} /* (11, 12, 25) {real, imag} */,
  {32'h3ef58bbd, 32'h4042b3f5} /* (11, 12, 24) {real, imag} */,
  {32'hbf80fbdb, 32'hbf812fe6} /* (11, 12, 23) {real, imag} */,
  {32'hc00792a8, 32'hc03299ed} /* (11, 12, 22) {real, imag} */,
  {32'h3ec6f48f, 32'hc05374ad} /* (11, 12, 21) {real, imag} */,
  {32'hbeedfdab, 32'hc06fe19f} /* (11, 12, 20) {real, imag} */,
  {32'hc0132842, 32'h403393c0} /* (11, 12, 19) {real, imag} */,
  {32'h4037db7a, 32'hc07d2c5e} /* (11, 12, 18) {real, imag} */,
  {32'hbfa0335c, 32'hc02d6f02} /* (11, 12, 17) {real, imag} */,
  {32'hbef4b74e, 32'hbddbb3dd} /* (11, 12, 16) {real, imag} */,
  {32'hbf6242e5, 32'hc01b14d2} /* (11, 12, 15) {real, imag} */,
  {32'h3e19084f, 32'h3fb9b5d4} /* (11, 12, 14) {real, imag} */,
  {32'h3f8887d2, 32'hc06a0afc} /* (11, 12, 13) {real, imag} */,
  {32'hbd17b16f, 32'hbf66aa35} /* (11, 12, 12) {real, imag} */,
  {32'hbf870c26, 32'hbf59269d} /* (11, 12, 11) {real, imag} */,
  {32'h3f5c98c9, 32'h3d828133} /* (11, 12, 10) {real, imag} */,
  {32'h3f07ad0d, 32'h3f29e3ad} /* (11, 12, 9) {real, imag} */,
  {32'hbfdb9d08, 32'hbfc244b1} /* (11, 12, 8) {real, imag} */,
  {32'h40335867, 32'hbeea0727} /* (11, 12, 7) {real, imag} */,
  {32'h3f253058, 32'hbe6b0dc7} /* (11, 12, 6) {real, imag} */,
  {32'hbf8850bc, 32'hc0067273} /* (11, 12, 5) {real, imag} */,
  {32'h3f05724a, 32'h3e67668f} /* (11, 12, 4) {real, imag} */,
  {32'hbfa66bdd, 32'h3f23df64} /* (11, 12, 3) {real, imag} */,
  {32'hc0093ae7, 32'h401bef47} /* (11, 12, 2) {real, imag} */,
  {32'hc012b468, 32'hc000ce3b} /* (11, 12, 1) {real, imag} */,
  {32'h3e6f1eb1, 32'hbfca36ed} /* (11, 12, 0) {real, imag} */,
  {32'hc08906a2, 32'h3f7e6603} /* (11, 11, 31) {real, imag} */,
  {32'hbfef6388, 32'h407fc043} /* (11, 11, 30) {real, imag} */,
  {32'hc00babd5, 32'h3f34306d} /* (11, 11, 29) {real, imag} */,
  {32'hbee45db7, 32'hbef5b72e} /* (11, 11, 28) {real, imag} */,
  {32'hbf3a6105, 32'hbfd70572} /* (11, 11, 27) {real, imag} */,
  {32'h3fb78b0b, 32'hc01cc3d4} /* (11, 11, 26) {real, imag} */,
  {32'hc017e1f5, 32'hbfa09256} /* (11, 11, 25) {real, imag} */,
  {32'h40078cb1, 32'hbff3131c} /* (11, 11, 24) {real, imag} */,
  {32'hbf31fd9a, 32'hbe3bd98a} /* (11, 11, 23) {real, imag} */,
  {32'h40054836, 32'hbfa7b376} /* (11, 11, 22) {real, imag} */,
  {32'h3f5ded65, 32'hbfb4694f} /* (11, 11, 21) {real, imag} */,
  {32'hbfaf74c9, 32'hc08ca1de} /* (11, 11, 20) {real, imag} */,
  {32'hbfbf0b3c, 32'hbf9356cf} /* (11, 11, 19) {real, imag} */,
  {32'hc0661975, 32'hc02a01ef} /* (11, 11, 18) {real, imag} */,
  {32'hbf099bde, 32'h402c1c24} /* (11, 11, 17) {real, imag} */,
  {32'hbf4fa3c0, 32'hbf7ae806} /* (11, 11, 16) {real, imag} */,
  {32'h3eb9e2f6, 32'h3f9050b9} /* (11, 11, 15) {real, imag} */,
  {32'hbf71d263, 32'hc018e844} /* (11, 11, 14) {real, imag} */,
  {32'hbf70072f, 32'hbf48b902} /* (11, 11, 13) {real, imag} */,
  {32'h4000173e, 32'h3f65af6c} /* (11, 11, 12) {real, imag} */,
  {32'hbdef3216, 32'h406e0b4b} /* (11, 11, 11) {real, imag} */,
  {32'h3f14663d, 32'hbfcc6b3e} /* (11, 11, 10) {real, imag} */,
  {32'hbfdb6f59, 32'hbf87204e} /* (11, 11, 9) {real, imag} */,
  {32'h3eeea5fd, 32'h3f7f4d99} /* (11, 11, 8) {real, imag} */,
  {32'hbdc6f15d, 32'hbeb5bfc6} /* (11, 11, 7) {real, imag} */,
  {32'hbf2538d6, 32'hbfef03a3} /* (11, 11, 6) {real, imag} */,
  {32'hbecd51ff, 32'hbef3a6d9} /* (11, 11, 5) {real, imag} */,
  {32'hc06dd8a1, 32'h4074044f} /* (11, 11, 4) {real, imag} */,
  {32'hc0447e9c, 32'h3f023503} /* (11, 11, 3) {real, imag} */,
  {32'hbf80046f, 32'h3de5c42a} /* (11, 11, 2) {real, imag} */,
  {32'hbda77b81, 32'hbf535290} /* (11, 11, 1) {real, imag} */,
  {32'hbf924a23, 32'hc015a117} /* (11, 11, 0) {real, imag} */,
  {32'hbee5d1c0, 32'h3e129e3a} /* (11, 10, 31) {real, imag} */,
  {32'hbf5549a4, 32'hbf154948} /* (11, 10, 30) {real, imag} */,
  {32'h40121e3a, 32'hbfbc74fa} /* (11, 10, 29) {real, imag} */,
  {32'h3ef1d154, 32'h40099466} /* (11, 10, 28) {real, imag} */,
  {32'h400c206d, 32'hbf795a1f} /* (11, 10, 27) {real, imag} */,
  {32'hbf49ebbb, 32'hc01c821d} /* (11, 10, 26) {real, imag} */,
  {32'hbe266f6a, 32'h409e0088} /* (11, 10, 25) {real, imag} */,
  {32'h40be212d, 32'hc09c66d9} /* (11, 10, 24) {real, imag} */,
  {32'hc096f2ba, 32'h401f8404} /* (11, 10, 23) {real, imag} */,
  {32'hbfd0e7f0, 32'hbd4c5904} /* (11, 10, 22) {real, imag} */,
  {32'h3f98169f, 32'h3f0b38c1} /* (11, 10, 21) {real, imag} */,
  {32'hc0275ea1, 32'h3f84c2c8} /* (11, 10, 20) {real, imag} */,
  {32'h3f3961a8, 32'hbf7618a4} /* (11, 10, 19) {real, imag} */,
  {32'hc0096c94, 32'h400cbd35} /* (11, 10, 18) {real, imag} */,
  {32'h3fb6049a, 32'hbe51f497} /* (11, 10, 17) {real, imag} */,
  {32'hbe252814, 32'hbfa667e4} /* (11, 10, 16) {real, imag} */,
  {32'hbe0d85c0, 32'h3ef15fa1} /* (11, 10, 15) {real, imag} */,
  {32'h405d3c32, 32'h3faceb75} /* (11, 10, 14) {real, imag} */,
  {32'hc055514a, 32'hbfbc1784} /* (11, 10, 13) {real, imag} */,
  {32'h405506f2, 32'h3f2b473b} /* (11, 10, 12) {real, imag} */,
  {32'h3f30d726, 32'hbea651d6} /* (11, 10, 11) {real, imag} */,
  {32'h3fcf626b, 32'h4043db4d} /* (11, 10, 10) {real, imag} */,
  {32'hc02e5550, 32'hc09b5cc6} /* (11, 10, 9) {real, imag} */,
  {32'h3fbe059d, 32'hc03622a6} /* (11, 10, 8) {real, imag} */,
  {32'h3f3a3e76, 32'hbdcaaa59} /* (11, 10, 7) {real, imag} */,
  {32'h3f59b8bb, 32'hbf585b72} /* (11, 10, 6) {real, imag} */,
  {32'hbf8e5fda, 32'hbfb40ea8} /* (11, 10, 5) {real, imag} */,
  {32'hbf9b5e9c, 32'h3fac0757} /* (11, 10, 4) {real, imag} */,
  {32'hbf56ce19, 32'h40095724} /* (11, 10, 3) {real, imag} */,
  {32'hbfe6014d, 32'hbf3efff2} /* (11, 10, 2) {real, imag} */,
  {32'hc067df18, 32'h4014797a} /* (11, 10, 1) {real, imag} */,
  {32'hbf56ea16, 32'h408a1edd} /* (11, 10, 0) {real, imag} */,
  {32'hc00a72e8, 32'hbeee4b1e} /* (11, 9, 31) {real, imag} */,
  {32'h40096e6b, 32'h4002ca42} /* (11, 9, 30) {real, imag} */,
  {32'hc0028fab, 32'h3e601c48} /* (11, 9, 29) {real, imag} */,
  {32'hc04ef84a, 32'h3f009ef8} /* (11, 9, 28) {real, imag} */,
  {32'hbfdfb7ad, 32'h400102ff} /* (11, 9, 27) {real, imag} */,
  {32'hbdc8c7ff, 32'hbf0979ce} /* (11, 9, 26) {real, imag} */,
  {32'h3ffe2e18, 32'h402c0a1b} /* (11, 9, 25) {real, imag} */,
  {32'hc037efbf, 32'h401b890d} /* (11, 9, 24) {real, imag} */,
  {32'hc02025c9, 32'h3fe131c9} /* (11, 9, 23) {real, imag} */,
  {32'hc07690a9, 32'hc040391e} /* (11, 9, 22) {real, imag} */,
  {32'h3fa21831, 32'hbf9534e8} /* (11, 9, 21) {real, imag} */,
  {32'hbf46dc88, 32'hbf8eef93} /* (11, 9, 20) {real, imag} */,
  {32'h3f88574a, 32'h3f9752bf} /* (11, 9, 19) {real, imag} */,
  {32'hbf558cc9, 32'h3e84ba23} /* (11, 9, 18) {real, imag} */,
  {32'hbf8a61b0, 32'hc087af4e} /* (11, 9, 17) {real, imag} */,
  {32'h3f6745cb, 32'hbfd96933} /* (11, 9, 16) {real, imag} */,
  {32'hbfbf33a8, 32'hbeced4bb} /* (11, 9, 15) {real, imag} */,
  {32'hbfeba8f5, 32'h3f2b5c9e} /* (11, 9, 14) {real, imag} */,
  {32'h3f41b52b, 32'h400800ab} /* (11, 9, 13) {real, imag} */,
  {32'h3fbdd610, 32'h40222ac7} /* (11, 9, 12) {real, imag} */,
  {32'hc01f1de0, 32'h3f281372} /* (11, 9, 11) {real, imag} */,
  {32'hbffa931a, 32'hbe06bb8f} /* (11, 9, 10) {real, imag} */,
  {32'hc0072b9d, 32'hbe8200ef} /* (11, 9, 9) {real, imag} */,
  {32'h401b2b48, 32'h3f02a021} /* (11, 9, 8) {real, imag} */,
  {32'hbe4e6550, 32'h3f2c67eb} /* (11, 9, 7) {real, imag} */,
  {32'h3f1d6da6, 32'h400a6c5d} /* (11, 9, 6) {real, imag} */,
  {32'h3feb19a6, 32'hbf7067ee} /* (11, 9, 5) {real, imag} */,
  {32'hbd8c66a2, 32'h3fb154fb} /* (11, 9, 4) {real, imag} */,
  {32'h3e96484e, 32'hc0280bd1} /* (11, 9, 3) {real, imag} */,
  {32'hbdb8f85c, 32'hc0161168} /* (11, 9, 2) {real, imag} */,
  {32'h409f3251, 32'h3ec3ef9c} /* (11, 9, 1) {real, imag} */,
  {32'h40325ad0, 32'hc0437eda} /* (11, 9, 0) {real, imag} */,
  {32'hbed1e88a, 32'hbfc50d44} /* (11, 8, 31) {real, imag} */,
  {32'hbfc34675, 32'h3f5f60e6} /* (11, 8, 30) {real, imag} */,
  {32'hbf8e72b2, 32'h3f5bcc39} /* (11, 8, 29) {real, imag} */,
  {32'h3ff040ca, 32'hc0041b37} /* (11, 8, 28) {real, imag} */,
  {32'h3e27e788, 32'hbffd182f} /* (11, 8, 27) {real, imag} */,
  {32'h3f0dd042, 32'hbf0156e2} /* (11, 8, 26) {real, imag} */,
  {32'hc093e57d, 32'hbfc3597e} /* (11, 8, 25) {real, imag} */,
  {32'hbfd1c85e, 32'hbfee92b7} /* (11, 8, 24) {real, imag} */,
  {32'hbef17046, 32'h400a2e36} /* (11, 8, 23) {real, imag} */,
  {32'h40856658, 32'h4006b1ad} /* (11, 8, 22) {real, imag} */,
  {32'h4092bf08, 32'h3e06f85e} /* (11, 8, 21) {real, imag} */,
  {32'hbe880eef, 32'hbfca28d2} /* (11, 8, 20) {real, imag} */,
  {32'hbe024d93, 32'h3f06fcf7} /* (11, 8, 19) {real, imag} */,
  {32'h400e1da0, 32'hbff064b9} /* (11, 8, 18) {real, imag} */,
  {32'hbfa79d1e, 32'hbf9c2503} /* (11, 8, 17) {real, imag} */,
  {32'h3f6347a5, 32'hbd188e42} /* (11, 8, 16) {real, imag} */,
  {32'hbfa7be59, 32'h3f2c8133} /* (11, 8, 15) {real, imag} */,
  {32'hbf931733, 32'h3f18fe43} /* (11, 8, 14) {real, imag} */,
  {32'h3fc959ef, 32'h40a0b63d} /* (11, 8, 13) {real, imag} */,
  {32'hbedd36b4, 32'h3fc21ab2} /* (11, 8, 12) {real, imag} */,
  {32'hbed7b49b, 32'hbffe4493} /* (11, 8, 11) {real, imag} */,
  {32'hbfff125c, 32'hbfbf64f1} /* (11, 8, 10) {real, imag} */,
  {32'hbfc7fda6, 32'hbf2fde58} /* (11, 8, 9) {real, imag} */,
  {32'h4051e72e, 32'hbe7dab3e} /* (11, 8, 8) {real, imag} */,
  {32'h40434d19, 32'h3e353c20} /* (11, 8, 7) {real, imag} */,
  {32'hc061918a, 32'h3fdf0f92} /* (11, 8, 6) {real, imag} */,
  {32'hbfa9bbd2, 32'h4012cb4c} /* (11, 8, 5) {real, imag} */,
  {32'hc00a5606, 32'h3feb09ea} /* (11, 8, 4) {real, imag} */,
  {32'h3f943f0d, 32'h3d27080e} /* (11, 8, 3) {real, imag} */,
  {32'hbfb92b4e, 32'h3c5ac838} /* (11, 8, 2) {real, imag} */,
  {32'h3d948aa4, 32'hbf89e71d} /* (11, 8, 1) {real, imag} */,
  {32'h3f533ab1, 32'h3f762b7d} /* (11, 8, 0) {real, imag} */,
  {32'h4074ca4d, 32'hbf7e1b77} /* (11, 7, 31) {real, imag} */,
  {32'hc00639c0, 32'hbe4b436b} /* (11, 7, 30) {real, imag} */,
  {32'h402bd3ad, 32'h40745c28} /* (11, 7, 29) {real, imag} */,
  {32'h3d5bb6f3, 32'hbf9cb73c} /* (11, 7, 28) {real, imag} */,
  {32'hc04c0859, 32'h3f3ee9e8} /* (11, 7, 27) {real, imag} */,
  {32'hbfb2dd6a, 32'hbf990f96} /* (11, 7, 26) {real, imag} */,
  {32'hbedfac49, 32'hbf7124f4} /* (11, 7, 25) {real, imag} */,
  {32'h400e1184, 32'hbed003d6} /* (11, 7, 24) {real, imag} */,
  {32'hc038c07f, 32'hbf99dc3e} /* (11, 7, 23) {real, imag} */,
  {32'h3e797008, 32'h407db43f} /* (11, 7, 22) {real, imag} */,
  {32'hc02e825a, 32'hbe64a38e} /* (11, 7, 21) {real, imag} */,
  {32'h4096dfa8, 32'h3fd4b642} /* (11, 7, 20) {real, imag} */,
  {32'hbf890f46, 32'h406052bf} /* (11, 7, 19) {real, imag} */,
  {32'hbec1c3a0, 32'hbf81cad2} /* (11, 7, 18) {real, imag} */,
  {32'h3f21e498, 32'h3f0188ee} /* (11, 7, 17) {real, imag} */,
  {32'hc001d7be, 32'hbe465af5} /* (11, 7, 16) {real, imag} */,
  {32'hbfb5b28b, 32'h4005233a} /* (11, 7, 15) {real, imag} */,
  {32'h3f464e0a, 32'hbfbac320} /* (11, 7, 14) {real, imag} */,
  {32'hc001a47d, 32'hc02d0695} /* (11, 7, 13) {real, imag} */,
  {32'hbe76afc3, 32'hbd8d39c2} /* (11, 7, 12) {real, imag} */,
  {32'h403a1907, 32'h4008e4a2} /* (11, 7, 11) {real, imag} */,
  {32'hbf23d677, 32'hbf910cac} /* (11, 7, 10) {real, imag} */,
  {32'h3f6f70cf, 32'hb97e78f8} /* (11, 7, 9) {real, imag} */,
  {32'h4031f627, 32'h3f434b65} /* (11, 7, 8) {real, imag} */,
  {32'h3fb06c72, 32'h403d3d64} /* (11, 7, 7) {real, imag} */,
  {32'h4085617d, 32'hbdeec9da} /* (11, 7, 6) {real, imag} */,
  {32'hc00272df, 32'hc08f6688} /* (11, 7, 5) {real, imag} */,
  {32'h3fe79009, 32'h3f77b9d6} /* (11, 7, 4) {real, imag} */,
  {32'hbfa28867, 32'hc06e4237} /* (11, 7, 3) {real, imag} */,
  {32'hbcdd89a7, 32'h3e91ebe6} /* (11, 7, 2) {real, imag} */,
  {32'h40896800, 32'hbf8c6d8f} /* (11, 7, 1) {real, imag} */,
  {32'hc0523611, 32'h3faa0fd6} /* (11, 7, 0) {real, imag} */,
  {32'h40b78efd, 32'h3ff6ba9a} /* (11, 6, 31) {real, imag} */,
  {32'hbe795c78, 32'h3fb3d539} /* (11, 6, 30) {real, imag} */,
  {32'hc02a9bbe, 32'hc010b18f} /* (11, 6, 29) {real, imag} */,
  {32'h3fd8d137, 32'hbf53f608} /* (11, 6, 28) {real, imag} */,
  {32'hc01ac7c0, 32'h3f84e087} /* (11, 6, 27) {real, imag} */,
  {32'hbfff8755, 32'hbf8621a6} /* (11, 6, 26) {real, imag} */,
  {32'hbee5fda1, 32'hbf9a3f49} /* (11, 6, 25) {real, imag} */,
  {32'hc065a4b5, 32'h40205e9f} /* (11, 6, 24) {real, imag} */,
  {32'h3f57e807, 32'hbee172d2} /* (11, 6, 23) {real, imag} */,
  {32'h3e5e30d2, 32'hc02b1332} /* (11, 6, 22) {real, imag} */,
  {32'hbf4e8969, 32'h3fb94286} /* (11, 6, 21) {real, imag} */,
  {32'h3ff2b7b4, 32'h404b0aaf} /* (11, 6, 20) {real, imag} */,
  {32'hbfe7eee8, 32'hbff8cdc7} /* (11, 6, 19) {real, imag} */,
  {32'h3ffbf315, 32'h3fd2c8e3} /* (11, 6, 18) {real, imag} */,
  {32'h3f970194, 32'hbff52ec9} /* (11, 6, 17) {real, imag} */,
  {32'h3fc83131, 32'h3fde0c38} /* (11, 6, 16) {real, imag} */,
  {32'h3f0ce067, 32'hbf67a811} /* (11, 6, 15) {real, imag} */,
  {32'hbf353a97, 32'h3f75ba74} /* (11, 6, 14) {real, imag} */,
  {32'hbf67447c, 32'h3efd710f} /* (11, 6, 13) {real, imag} */,
  {32'hbdbc56de, 32'h40146082} /* (11, 6, 12) {real, imag} */,
  {32'h3f3f4eef, 32'h401f13f8} /* (11, 6, 11) {real, imag} */,
  {32'hbe1c32cb, 32'h409c1725} /* (11, 6, 10) {real, imag} */,
  {32'h4039d466, 32'h40056b0b} /* (11, 6, 9) {real, imag} */,
  {32'hc01f57df, 32'hbea311cf} /* (11, 6, 8) {real, imag} */,
  {32'hbff5512b, 32'hbf814a29} /* (11, 6, 7) {real, imag} */,
  {32'hbff13e56, 32'h401cdf96} /* (11, 6, 6) {real, imag} */,
  {32'h3fe23ff5, 32'hbf574563} /* (11, 6, 5) {real, imag} */,
  {32'h401e9db7, 32'hbff7aba0} /* (11, 6, 4) {real, imag} */,
  {32'h3fd91974, 32'h3ec68958} /* (11, 6, 3) {real, imag} */,
  {32'hbe9c760a, 32'h3fdfb3d4} /* (11, 6, 2) {real, imag} */,
  {32'h4001f84b, 32'h3f52d613} /* (11, 6, 1) {real, imag} */,
  {32'hc070d5c4, 32'hbf2bb91e} /* (11, 6, 0) {real, imag} */,
  {32'hc020077c, 32'h405e5d75} /* (11, 5, 31) {real, imag} */,
  {32'h3fd9d152, 32'h401108c9} /* (11, 5, 30) {real, imag} */,
  {32'h3e9c1be3, 32'h3d30678c} /* (11, 5, 29) {real, imag} */,
  {32'h3f845a37, 32'hc039cc84} /* (11, 5, 28) {real, imag} */,
  {32'h3fec4949, 32'hbf960986} /* (11, 5, 27) {real, imag} */,
  {32'hbf1c9fde, 32'h3f0fed86} /* (11, 5, 26) {real, imag} */,
  {32'hbfa37a0d, 32'h400b2349} /* (11, 5, 25) {real, imag} */,
  {32'h3eeea292, 32'h3ed7490a} /* (11, 5, 24) {real, imag} */,
  {32'h3d97b5d8, 32'hbfe4c1ed} /* (11, 5, 23) {real, imag} */,
  {32'hc022c9f7, 32'h3ed8b16e} /* (11, 5, 22) {real, imag} */,
  {32'h3fa2bee0, 32'hbff3523a} /* (11, 5, 21) {real, imag} */,
  {32'h3f82ce52, 32'h3f912def} /* (11, 5, 20) {real, imag} */,
  {32'hbf32ece2, 32'h404b9f53} /* (11, 5, 19) {real, imag} */,
  {32'hbf839e61, 32'hbf4db962} /* (11, 5, 18) {real, imag} */,
  {32'hbe3d883a, 32'h3ea8509f} /* (11, 5, 17) {real, imag} */,
  {32'h3fea6f47, 32'hbdad585e} /* (11, 5, 16) {real, imag} */,
  {32'h4016bccf, 32'hbf52a3fb} /* (11, 5, 15) {real, imag} */,
  {32'hbfd45e1d, 32'h3ec041ca} /* (11, 5, 14) {real, imag} */,
  {32'hc017a706, 32'h3f9ebc3e} /* (11, 5, 13) {real, imag} */,
  {32'hc0598c76, 32'hbe9864dc} /* (11, 5, 12) {real, imag} */,
  {32'h3ff3ff47, 32'h4037d502} /* (11, 5, 11) {real, imag} */,
  {32'hbeb16946, 32'h3ff1242b} /* (11, 5, 10) {real, imag} */,
  {32'h3fae60cf, 32'hc03b7957} /* (11, 5, 9) {real, imag} */,
  {32'h4030f941, 32'h3f7ac793} /* (11, 5, 8) {real, imag} */,
  {32'hc0128b94, 32'hbffbde9e} /* (11, 5, 7) {real, imag} */,
  {32'hbf686a81, 32'hbf4e5870} /* (11, 5, 6) {real, imag} */,
  {32'h3f506413, 32'h403d684a} /* (11, 5, 5) {real, imag} */,
  {32'hbf0db96f, 32'hc031cc62} /* (11, 5, 4) {real, imag} */,
  {32'hbe020cc0, 32'hc011495a} /* (11, 5, 3) {real, imag} */,
  {32'h400eab21, 32'hbf7e72b1} /* (11, 5, 2) {real, imag} */,
  {32'hc0cfde39, 32'hc00ec508} /* (11, 5, 1) {real, imag} */,
  {32'hc0142e01, 32'h3f69279a} /* (11, 5, 0) {real, imag} */,
  {32'h3ef2fb35, 32'h3f622a32} /* (11, 4, 31) {real, imag} */,
  {32'h3da6de0a, 32'hc040c515} /* (11, 4, 30) {real, imag} */,
  {32'hbe82165c, 32'h3fe6a094} /* (11, 4, 29) {real, imag} */,
  {32'h3f02e598, 32'hbff0b2f2} /* (11, 4, 28) {real, imag} */,
  {32'hc08fdc85, 32'h400d36ac} /* (11, 4, 27) {real, imag} */,
  {32'h4004b748, 32'hbfbabcaa} /* (11, 4, 26) {real, imag} */,
  {32'hbf14df6d, 32'h408f7186} /* (11, 4, 25) {real, imag} */,
  {32'h3ed8eb17, 32'h3f12b04d} /* (11, 4, 24) {real, imag} */,
  {32'hbfd33170, 32'hbf77805f} /* (11, 4, 23) {real, imag} */,
  {32'hc0540cab, 32'h3e498505} /* (11, 4, 22) {real, imag} */,
  {32'hbd980a98, 32'h3f9a61d0} /* (11, 4, 21) {real, imag} */,
  {32'h3fd2d8da, 32'h3ff70c57} /* (11, 4, 20) {real, imag} */,
  {32'h3fd95fd4, 32'hbf8571df} /* (11, 4, 19) {real, imag} */,
  {32'h3e2b20ce, 32'hbfea8d65} /* (11, 4, 18) {real, imag} */,
  {32'hbc413bbe, 32'hc01a0724} /* (11, 4, 17) {real, imag} */,
  {32'hbe939bb3, 32'h3feddea6} /* (11, 4, 16) {real, imag} */,
  {32'h3fefc660, 32'h3e61125a} /* (11, 4, 15) {real, imag} */,
  {32'hbe4d77dd, 32'h3fb8a10e} /* (11, 4, 14) {real, imag} */,
  {32'hc03d5931, 32'hbeed9433} /* (11, 4, 13) {real, imag} */,
  {32'hc02e7302, 32'h400ed925} /* (11, 4, 12) {real, imag} */,
  {32'hc0205b87, 32'h3ef9842c} /* (11, 4, 11) {real, imag} */,
  {32'h3e2832d7, 32'hc00cc0fd} /* (11, 4, 10) {real, imag} */,
  {32'hbe150668, 32'hc0655e30} /* (11, 4, 9) {real, imag} */,
  {32'hbea0b66d, 32'hbf87dece} /* (11, 4, 8) {real, imag} */,
  {32'h40862ecc, 32'hc019cad0} /* (11, 4, 7) {real, imag} */,
  {32'hc066ff14, 32'h4017c864} /* (11, 4, 6) {real, imag} */,
  {32'hc01e8834, 32'h3fa777b0} /* (11, 4, 5) {real, imag} */,
  {32'h3f43eb6a, 32'h3ff3cc68} /* (11, 4, 4) {real, imag} */,
  {32'h405abfbf, 32'hbf9e813b} /* (11, 4, 3) {real, imag} */,
  {32'hc064cefb, 32'hc0972fb3} /* (11, 4, 2) {real, imag} */,
  {32'h4098d628, 32'h3d8ca88c} /* (11, 4, 1) {real, imag} */,
  {32'h3fbca97c, 32'hbf1c5702} /* (11, 4, 0) {real, imag} */,
  {32'h3fb54741, 32'h407c8032} /* (11, 3, 31) {real, imag} */,
  {32'hbf558be6, 32'hc0905791} /* (11, 3, 30) {real, imag} */,
  {32'h400a63c3, 32'h3fc65da5} /* (11, 3, 29) {real, imag} */,
  {32'h3ff69c34, 32'hbfa54b53} /* (11, 3, 28) {real, imag} */,
  {32'h3f9f362b, 32'hc0909ae0} /* (11, 3, 27) {real, imag} */,
  {32'hc0042671, 32'h4013c982} /* (11, 3, 26) {real, imag} */,
  {32'hbfedf34a, 32'hc05bd519} /* (11, 3, 25) {real, imag} */,
  {32'hbe8ea97c, 32'hbffe52ea} /* (11, 3, 24) {real, imag} */,
  {32'h403063af, 32'hbfcbc745} /* (11, 3, 23) {real, imag} */,
  {32'hc002f4ef, 32'hbf6397eb} /* (11, 3, 22) {real, imag} */,
  {32'hc03c1de5, 32'hbf42eb9e} /* (11, 3, 21) {real, imag} */,
  {32'hbfa057bd, 32'h40857f6b} /* (11, 3, 20) {real, imag} */,
  {32'hbfa3834d, 32'hbebfe63a} /* (11, 3, 19) {real, imag} */,
  {32'hbfadb0b0, 32'h3f937ceb} /* (11, 3, 18) {real, imag} */,
  {32'h3f092744, 32'h3fab6932} /* (11, 3, 17) {real, imag} */,
  {32'hc01192f5, 32'hbf0e3d21} /* (11, 3, 16) {real, imag} */,
  {32'hbf73b350, 32'hbf86d639} /* (11, 3, 15) {real, imag} */,
  {32'h3ff6f097, 32'h3fb01e9f} /* (11, 3, 14) {real, imag} */,
  {32'h3fa11eb7, 32'hbf480516} /* (11, 3, 13) {real, imag} */,
  {32'hbfad19d0, 32'h4014b63f} /* (11, 3, 12) {real, imag} */,
  {32'h3ff24116, 32'h4012f167} /* (11, 3, 11) {real, imag} */,
  {32'hbff439ea, 32'hbe8d5878} /* (11, 3, 10) {real, imag} */,
  {32'h4060cba1, 32'hbf3e06b3} /* (11, 3, 9) {real, imag} */,
  {32'hbf8a6b1b, 32'h402b442e} /* (11, 3, 8) {real, imag} */,
  {32'h3f904625, 32'h3e1476d5} /* (11, 3, 7) {real, imag} */,
  {32'h3f6d054c, 32'hbf90c87e} /* (11, 3, 6) {real, imag} */,
  {32'hbf3589ff, 32'hbf629589} /* (11, 3, 5) {real, imag} */,
  {32'hbf909028, 32'h3f83286b} /* (11, 3, 4) {real, imag} */,
  {32'hc04d6430, 32'hbfd8c081} /* (11, 3, 3) {real, imag} */,
  {32'hc07d042f, 32'hbe05ac81} /* (11, 3, 2) {real, imag} */,
  {32'hbf7ca812, 32'h3fe1b321} /* (11, 3, 1) {real, imag} */,
  {32'h405f37f9, 32'h3fc8fa33} /* (11, 3, 0) {real, imag} */,
  {32'hc0dde7e2, 32'h40774c7a} /* (11, 2, 31) {real, imag} */,
  {32'h40cfdbd2, 32'hbeb9a1f9} /* (11, 2, 30) {real, imag} */,
  {32'h3e8db507, 32'hbd133e04} /* (11, 2, 29) {real, imag} */,
  {32'h3f127a9c, 32'hbe51d806} /* (11, 2, 28) {real, imag} */,
  {32'hbe3b92bd, 32'h3f3c4d6c} /* (11, 2, 27) {real, imag} */,
  {32'h3f351b61, 32'h40057ebe} /* (11, 2, 26) {real, imag} */,
  {32'hc03127cb, 32'h409558ca} /* (11, 2, 25) {real, imag} */,
  {32'h3f07fbcc, 32'hc0684a1d} /* (11, 2, 24) {real, imag} */,
  {32'h403cda25, 32'h3e546a10} /* (11, 2, 23) {real, imag} */,
  {32'h3ed6a724, 32'h3f9c9315} /* (11, 2, 22) {real, imag} */,
  {32'h3e82da76, 32'hbf86a30c} /* (11, 2, 21) {real, imag} */,
  {32'hbf9e6b0e, 32'h400775bd} /* (11, 2, 20) {real, imag} */,
  {32'h3fe3ffd1, 32'h3ef5a885} /* (11, 2, 19) {real, imag} */,
  {32'hbf67c6ef, 32'h3e7738a4} /* (11, 2, 18) {real, imag} */,
  {32'hbec11458, 32'h40140693} /* (11, 2, 17) {real, imag} */,
  {32'h3b35d331, 32'h3f507b76} /* (11, 2, 16) {real, imag} */,
  {32'h3f587d0c, 32'hc0399f35} /* (11, 2, 15) {real, imag} */,
  {32'hbff81028, 32'hbeb58d4c} /* (11, 2, 14) {real, imag} */,
  {32'hbfdea654, 32'hbf1a3f8d} /* (11, 2, 13) {real, imag} */,
  {32'h40932071, 32'h3e508b69} /* (11, 2, 12) {real, imag} */,
  {32'h4000917d, 32'h40453c17} /* (11, 2, 11) {real, imag} */,
  {32'hc09f8aaf, 32'hbf031d29} /* (11, 2, 10) {real, imag} */,
  {32'hc0068ea7, 32'hc02902c6} /* (11, 2, 9) {real, imag} */,
  {32'hbf97f716, 32'h4066934f} /* (11, 2, 8) {real, imag} */,
  {32'h3fa78bfe, 32'h3fa8204b} /* (11, 2, 7) {real, imag} */,
  {32'h3f6ed9a5, 32'hbfffe64e} /* (11, 2, 6) {real, imag} */,
  {32'h40123ea6, 32'h3f065393} /* (11, 2, 5) {real, imag} */,
  {32'hc002089d, 32'hbfbaa0e6} /* (11, 2, 4) {real, imag} */,
  {32'hbf7e50f4, 32'hbd42d83d} /* (11, 2, 3) {real, imag} */,
  {32'h3f2fffd1, 32'hc0a8d90f} /* (11, 2, 2) {real, imag} */,
  {32'hbfd1a6c7, 32'h3f93fad1} /* (11, 2, 1) {real, imag} */,
  {32'hc064d99f, 32'h3e60e8f7} /* (11, 2, 0) {real, imag} */,
  {32'h3fab1fcf, 32'hc0545e40} /* (11, 1, 31) {real, imag} */,
  {32'hc088c9c8, 32'hbed34f0a} /* (11, 1, 30) {real, imag} */,
  {32'hbec2c814, 32'h3fe25dd3} /* (11, 1, 29) {real, imag} */,
  {32'h4000925a, 32'h409c0f50} /* (11, 1, 28) {real, imag} */,
  {32'hc0a27ac4, 32'h4014f00f} /* (11, 1, 27) {real, imag} */,
  {32'hc01862f6, 32'h3f18e742} /* (11, 1, 26) {real, imag} */,
  {32'hbf53e957, 32'hc0161357} /* (11, 1, 25) {real, imag} */,
  {32'h3fad385e, 32'hc0970be0} /* (11, 1, 24) {real, imag} */,
  {32'hbe8a4378, 32'hbf5afe45} /* (11, 1, 23) {real, imag} */,
  {32'hbf040ed4, 32'hbffda74e} /* (11, 1, 22) {real, imag} */,
  {32'hbef461d7, 32'hbf100575} /* (11, 1, 21) {real, imag} */,
  {32'h3f5475ea, 32'h4053aaa0} /* (11, 1, 20) {real, imag} */,
  {32'h3f295fbb, 32'hc02911ac} /* (11, 1, 19) {real, imag} */,
  {32'hbe3a74ac, 32'hbe58d53e} /* (11, 1, 18) {real, imag} */,
  {32'h4036ae06, 32'hc007aae6} /* (11, 1, 17) {real, imag} */,
  {32'hbee7ce01, 32'hbf847826} /* (11, 1, 16) {real, imag} */,
  {32'hbe59249e, 32'h3ff5abbf} /* (11, 1, 15) {real, imag} */,
  {32'h4088fc43, 32'hbfe744ed} /* (11, 1, 14) {real, imag} */,
  {32'h3fbd872e, 32'hbf39e714} /* (11, 1, 13) {real, imag} */,
  {32'hbe924442, 32'h3fc1bf1c} /* (11, 1, 12) {real, imag} */,
  {32'hbfc61399, 32'hbe4aa935} /* (11, 1, 11) {real, imag} */,
  {32'hbd811423, 32'h3f35fce1} /* (11, 1, 10) {real, imag} */,
  {32'h4028900f, 32'hbf9fb47f} /* (11, 1, 9) {real, imag} */,
  {32'hc082ae66, 32'h3ffd345c} /* (11, 1, 8) {real, imag} */,
  {32'hbfcb21e5, 32'hbf9db62c} /* (11, 1, 7) {real, imag} */,
  {32'h403aeecb, 32'hbf314612} /* (11, 1, 6) {real, imag} */,
  {32'hc03890c4, 32'h3fa3ab52} /* (11, 1, 5) {real, imag} */,
  {32'h3fad4cf9, 32'h3fd64ac0} /* (11, 1, 4) {real, imag} */,
  {32'h40181de8, 32'h3f53cb6b} /* (11, 1, 3) {real, imag} */,
  {32'hc0e4c1a5, 32'hc007de89} /* (11, 1, 2) {real, imag} */,
  {32'h41206b4f, 32'h3f84d39a} /* (11, 1, 1) {real, imag} */,
  {32'h40cae1a2, 32'hbfa40baf} /* (11, 1, 0) {real, imag} */,
  {32'h403b2e35, 32'hc0a67a93} /* (11, 0, 31) {real, imag} */,
  {32'h408e33fc, 32'h3ed6407a} /* (11, 0, 30) {real, imag} */,
  {32'h3fb14fca, 32'h4088222d} /* (11, 0, 29) {real, imag} */,
  {32'h3f28e0fe, 32'hbf213ad3} /* (11, 0, 28) {real, imag} */,
  {32'hc0375c99, 32'hc00cbb08} /* (11, 0, 27) {real, imag} */,
  {32'h3f8cfe43, 32'hbecb5782} /* (11, 0, 26) {real, imag} */,
  {32'hbf125de9, 32'h3ed12ea8} /* (11, 0, 25) {real, imag} */,
  {32'h408d1cc1, 32'h40d7b5e2} /* (11, 0, 24) {real, imag} */,
  {32'hc037921e, 32'h4075a332} /* (11, 0, 23) {real, imag} */,
  {32'hbf53d1b6, 32'h3fde753f} /* (11, 0, 22) {real, imag} */,
  {32'h3f5786da, 32'h3fede211} /* (11, 0, 21) {real, imag} */,
  {32'h3f6b7c4a, 32'hbf0d8289} /* (11, 0, 20) {real, imag} */,
  {32'hbf74d1a2, 32'hbec3865f} /* (11, 0, 19) {real, imag} */,
  {32'h3f5a4a53, 32'hbebedea8} /* (11, 0, 18) {real, imag} */,
  {32'hbf59dc98, 32'hbfdb4f82} /* (11, 0, 17) {real, imag} */,
  {32'h3f5d8d92, 32'hbf973574} /* (11, 0, 16) {real, imag} */,
  {32'hbf6294db, 32'h3f1e354e} /* (11, 0, 15) {real, imag} */,
  {32'h3d8dd622, 32'hc06ba86e} /* (11, 0, 14) {real, imag} */,
  {32'hc01543e0, 32'hbff8fd3d} /* (11, 0, 13) {real, imag} */,
  {32'h3f0fac48, 32'hbfc0e668} /* (11, 0, 12) {real, imag} */,
  {32'hbee0a41d, 32'hbf86f5d9} /* (11, 0, 11) {real, imag} */,
  {32'hbf6d346d, 32'hbf0aa7b9} /* (11, 0, 10) {real, imag} */,
  {32'hbfc8817d, 32'hbfdfc8f6} /* (11, 0, 9) {real, imag} */,
  {32'hbfb26c67, 32'h3f63d9a4} /* (11, 0, 8) {real, imag} */,
  {32'h3fc91117, 32'hc026aa7a} /* (11, 0, 7) {real, imag} */,
  {32'hbf9636ae, 32'hbeae3df9} /* (11, 0, 6) {real, imag} */,
  {32'h3fa88b87, 32'h3fda968b} /* (11, 0, 5) {real, imag} */,
  {32'h40390405, 32'hbf022669} /* (11, 0, 4) {real, imag} */,
  {32'h3fa9a847, 32'hbda83f92} /* (11, 0, 3) {real, imag} */,
  {32'hbf91f44e, 32'hc09baedb} /* (11, 0, 2) {real, imag} */,
  {32'h40a302b6, 32'hc02ec925} /* (11, 0, 1) {real, imag} */,
  {32'h4094392b, 32'hc02b81b0} /* (11, 0, 0) {real, imag} */,
  {32'hc013519c, 32'h409d3234} /* (10, 31, 31) {real, imag} */,
  {32'h3f905a44, 32'hc0568bca} /* (10, 31, 30) {real, imag} */,
  {32'h40a1adbe, 32'hbc738e87} /* (10, 31, 29) {real, imag} */,
  {32'hbfcc9ff5, 32'h3f1cd8cb} /* (10, 31, 28) {real, imag} */,
  {32'h40af2bc6, 32'hbfdcc56d} /* (10, 31, 27) {real, imag} */,
  {32'h3fcf82f2, 32'hbfa7ebfa} /* (10, 31, 26) {real, imag} */,
  {32'h3eaa8ff9, 32'h408c971f} /* (10, 31, 25) {real, imag} */,
  {32'hbf6a9a19, 32'h3fb404c2} /* (10, 31, 24) {real, imag} */,
  {32'hc06080df, 32'h3f9d9471} /* (10, 31, 23) {real, imag} */,
  {32'h3ef81ffa, 32'hbfd93b90} /* (10, 31, 22) {real, imag} */,
  {32'h3f04dc08, 32'h3fe5ee1f} /* (10, 31, 21) {real, imag} */,
  {32'hbfa9e635, 32'h3dde5f4b} /* (10, 31, 20) {real, imag} */,
  {32'hbf2fbc7e, 32'h3edd5b5f} /* (10, 31, 19) {real, imag} */,
  {32'hbf9bd7c2, 32'h3f5d377f} /* (10, 31, 18) {real, imag} */,
  {32'h3f8a9f7a, 32'hbf60c0bf} /* (10, 31, 17) {real, imag} */,
  {32'h3f14caa0, 32'hbe1a9b5a} /* (10, 31, 16) {real, imag} */,
  {32'hbf6814f4, 32'h3fdf62da} /* (10, 31, 15) {real, imag} */,
  {32'hbf14df8e, 32'h3f2dc6c0} /* (10, 31, 14) {real, imag} */,
  {32'h4012fa9e, 32'hc0447a5b} /* (10, 31, 13) {real, imag} */,
  {32'h3e05a053, 32'hbf0b269a} /* (10, 31, 12) {real, imag} */,
  {32'h3f18caf5, 32'h3f0d0c41} /* (10, 31, 11) {real, imag} */,
  {32'h3fcebf8d, 32'hbfa89fce} /* (10, 31, 10) {real, imag} */,
  {32'h3f4eb966, 32'h3ec22ad4} /* (10, 31, 9) {real, imag} */,
  {32'hbec60bcd, 32'hc02f71d8} /* (10, 31, 8) {real, imag} */,
  {32'hbf8e2b40, 32'h3fd1edb7} /* (10, 31, 7) {real, imag} */,
  {32'hbf633628, 32'hbff832b8} /* (10, 31, 6) {real, imag} */,
  {32'hbf6fb7af, 32'hc0c83fdd} /* (10, 31, 5) {real, imag} */,
  {32'hbfc19935, 32'h3cda9c06} /* (10, 31, 4) {real, imag} */,
  {32'h3f85465d, 32'h4066cbb6} /* (10, 31, 3) {real, imag} */,
  {32'h4027ba79, 32'hc07333e0} /* (10, 31, 2) {real, imag} */,
  {32'hc0583de1, 32'h3fc3d800} /* (10, 31, 1) {real, imag} */,
  {32'h4011481f, 32'h40aff7c3} /* (10, 31, 0) {real, imag} */,
  {32'h3f9ae4e7, 32'h40323dc3} /* (10, 30, 31) {real, imag} */,
  {32'hc0bfd73a, 32'hbe831296} /* (10, 30, 30) {real, imag} */,
  {32'hbefd11a0, 32'hc057060c} /* (10, 30, 29) {real, imag} */,
  {32'h3eb77618, 32'hc011790c} /* (10, 30, 28) {real, imag} */,
  {32'hc04b0a80, 32'h3fdb78e7} /* (10, 30, 27) {real, imag} */,
  {32'h3ea11706, 32'h3f815475} /* (10, 30, 26) {real, imag} */,
  {32'h3ea4010a, 32'hc039901d} /* (10, 30, 25) {real, imag} */,
  {32'hc0077c8d, 32'h408af7c0} /* (10, 30, 24) {real, imag} */,
  {32'hbfb45ca7, 32'h3f8587dd} /* (10, 30, 23) {real, imag} */,
  {32'hbf73b0fa, 32'hc0178c83} /* (10, 30, 22) {real, imag} */,
  {32'hbe078c0c, 32'hbf88ba3f} /* (10, 30, 21) {real, imag} */,
  {32'hbfc51771, 32'h3ff47655} /* (10, 30, 20) {real, imag} */,
  {32'h3f1bc4a8, 32'h40169f12} /* (10, 30, 19) {real, imag} */,
  {32'h4036106b, 32'h400bcfd9} /* (10, 30, 18) {real, imag} */,
  {32'h3e9b55a8, 32'hbf2c35de} /* (10, 30, 17) {real, imag} */,
  {32'h3edb7423, 32'h3c9fcb79} /* (10, 30, 16) {real, imag} */,
  {32'hbf72d12c, 32'hbeeebef3} /* (10, 30, 15) {real, imag} */,
  {32'h3f9cc296, 32'hc0221db0} /* (10, 30, 14) {real, imag} */,
  {32'h3f30f373, 32'hbf936f36} /* (10, 30, 13) {real, imag} */,
  {32'hbfd395ae, 32'hc02dd145} /* (10, 30, 12) {real, imag} */,
  {32'hbee5f106, 32'hbe72ec1b} /* (10, 30, 11) {real, imag} */,
  {32'h3e8c3f7f, 32'h3ee8ec53} /* (10, 30, 10) {real, imag} */,
  {32'hbfe32c25, 32'hbe0de28a} /* (10, 30, 9) {real, imag} */,
  {32'hc03e9bbc, 32'h3fae29da} /* (10, 30, 8) {real, imag} */,
  {32'hbed8a7a5, 32'h3febd391} /* (10, 30, 7) {real, imag} */,
  {32'h3faf83a3, 32'hbfdcdee8} /* (10, 30, 6) {real, imag} */,
  {32'hbe534921, 32'h401d1651} /* (10, 30, 5) {real, imag} */,
  {32'h3f26aca7, 32'h40e30dec} /* (10, 30, 4) {real, imag} */,
  {32'h407fe443, 32'hbe68f325} /* (10, 30, 3) {real, imag} */,
  {32'hbeb20184, 32'hbf023292} /* (10, 30, 2) {real, imag} */,
  {32'h40190bd2, 32'hc05497a5} /* (10, 30, 1) {real, imag} */,
  {32'h40acaeb1, 32'hbf8fbba7} /* (10, 30, 0) {real, imag} */,
  {32'hc0265a76, 32'hc0100153} /* (10, 29, 31) {real, imag} */,
  {32'hbf3bb982, 32'hbffbd3dd} /* (10, 29, 30) {real, imag} */,
  {32'hc0008451, 32'hbe31621a} /* (10, 29, 29) {real, imag} */,
  {32'hbf548813, 32'h3ebcd1f8} /* (10, 29, 28) {real, imag} */,
  {32'hbfb327da, 32'h40619aef} /* (10, 29, 27) {real, imag} */,
  {32'h3f3b97f5, 32'h407cdf92} /* (10, 29, 26) {real, imag} */,
  {32'hbfbfffda, 32'hbf48f322} /* (10, 29, 25) {real, imag} */,
  {32'hbf82d697, 32'hbf033314} /* (10, 29, 24) {real, imag} */,
  {32'h3fba1fd4, 32'h3fa70a26} /* (10, 29, 23) {real, imag} */,
  {32'hbe336dc2, 32'hbf73b12c} /* (10, 29, 22) {real, imag} */,
  {32'hbfb826c0, 32'hbf13d9c4} /* (10, 29, 21) {real, imag} */,
  {32'h40491993, 32'hbec9e3a5} /* (10, 29, 20) {real, imag} */,
  {32'hbfabe1bf, 32'hbf1dfbd2} /* (10, 29, 19) {real, imag} */,
  {32'hbf82c2a6, 32'hc0255835} /* (10, 29, 18) {real, imag} */,
  {32'h3f497730, 32'h3f0c3f0c} /* (10, 29, 17) {real, imag} */,
  {32'h3fce048d, 32'hbfae0ffa} /* (10, 29, 16) {real, imag} */,
  {32'h3cc754c5, 32'hbf85e220} /* (10, 29, 15) {real, imag} */,
  {32'hbf690c39, 32'h40428a0a} /* (10, 29, 14) {real, imag} */,
  {32'hbf1f313d, 32'h3f985513} /* (10, 29, 13) {real, imag} */,
  {32'h3f27e388, 32'h40314a14} /* (10, 29, 12) {real, imag} */,
  {32'hbfafb3d4, 32'h3f2317e7} /* (10, 29, 11) {real, imag} */,
  {32'hc0770bcf, 32'h3fc7273e} /* (10, 29, 10) {real, imag} */,
  {32'h3fba375b, 32'h3e4f4b7f} /* (10, 29, 9) {real, imag} */,
  {32'h3eb4d0cb, 32'h40940932} /* (10, 29, 8) {real, imag} */,
  {32'hbeca9f7f, 32'h3f616e66} /* (10, 29, 7) {real, imag} */,
  {32'h3e92e248, 32'h3f87c10c} /* (10, 29, 6) {real, imag} */,
  {32'h3fb19bb3, 32'hbffd024c} /* (10, 29, 5) {real, imag} */,
  {32'h3fc6018c, 32'hbf8030fb} /* (10, 29, 4) {real, imag} */,
  {32'hbe850959, 32'h3f550c50} /* (10, 29, 3) {real, imag} */,
  {32'hbf9ccab7, 32'hc06b367b} /* (10, 29, 2) {real, imag} */,
  {32'hc07375bd, 32'hc0082344} /* (10, 29, 1) {real, imag} */,
  {32'hc0203052, 32'hc0630c80} /* (10, 29, 0) {real, imag} */,
  {32'h3f62f05e, 32'h4001cebd} /* (10, 28, 31) {real, imag} */,
  {32'hbff0782d, 32'hc035e3dd} /* (10, 28, 30) {real, imag} */,
  {32'h3d37a4be, 32'h3f6e666d} /* (10, 28, 29) {real, imag} */,
  {32'hc0cd905f, 32'h3dc77034} /* (10, 28, 28) {real, imag} */,
  {32'h3e60aeea, 32'hc00442e0} /* (10, 28, 27) {real, imag} */,
  {32'hbd2d543b, 32'hbde1cfec} /* (10, 28, 26) {real, imag} */,
  {32'h3ff293fa, 32'h4002a851} /* (10, 28, 25) {real, imag} */,
  {32'h40088c8e, 32'h3f9ed6e7} /* (10, 28, 24) {real, imag} */,
  {32'h3d995478, 32'hbfe9edd7} /* (10, 28, 23) {real, imag} */,
  {32'h3cb0e54b, 32'hc0013807} /* (10, 28, 22) {real, imag} */,
  {32'h3ed525d2, 32'h3f87e1d2} /* (10, 28, 21) {real, imag} */,
  {32'hbfafed0e, 32'hbf6a6340} /* (10, 28, 20) {real, imag} */,
  {32'h3f788fef, 32'h3f472f31} /* (10, 28, 19) {real, imag} */,
  {32'hbfe636c9, 32'h3f946642} /* (10, 28, 18) {real, imag} */,
  {32'h3f58589e, 32'hbeb491c0} /* (10, 28, 17) {real, imag} */,
  {32'hbf6fd324, 32'hbf0d8995} /* (10, 28, 16) {real, imag} */,
  {32'h3f84c619, 32'h3fc3cf03} /* (10, 28, 15) {real, imag} */,
  {32'hbfbf7357, 32'h3f88dfd4} /* (10, 28, 14) {real, imag} */,
  {32'h3fb5ec17, 32'h3e6cdbf6} /* (10, 28, 13) {real, imag} */,
  {32'hc0b7a8dd, 32'h4042cf8c} /* (10, 28, 12) {real, imag} */,
  {32'h40858f03, 32'hbea27e98} /* (10, 28, 11) {real, imag} */,
  {32'hbe4e324a, 32'hc02d3aa5} /* (10, 28, 10) {real, imag} */,
  {32'hc016f291, 32'hbf341bee} /* (10, 28, 9) {real, imag} */,
  {32'h3fa9a75f, 32'hbe326ae0} /* (10, 28, 8) {real, imag} */,
  {32'h3fc2bacc, 32'h3fbcd10c} /* (10, 28, 7) {real, imag} */,
  {32'hc05fd663, 32'h4075e57b} /* (10, 28, 6) {real, imag} */,
  {32'hbf9fadd5, 32'hbf407440} /* (10, 28, 5) {real, imag} */,
  {32'h3e1d061d, 32'h404c3cc1} /* (10, 28, 4) {real, imag} */,
  {32'hc00ff585, 32'hc026c586} /* (10, 28, 3) {real, imag} */,
  {32'h3e7a1e6e, 32'hc01b86c2} /* (10, 28, 2) {real, imag} */,
  {32'h3fb931e5, 32'hbf5e7b61} /* (10, 28, 1) {real, imag} */,
  {32'hbf016d31, 32'h3fd061ae} /* (10, 28, 0) {real, imag} */,
  {32'hbffc1429, 32'hbead76cd} /* (10, 27, 31) {real, imag} */,
  {32'hbfc08945, 32'h3eb651a0} /* (10, 27, 30) {real, imag} */,
  {32'hc02d98e7, 32'hbfe97d78} /* (10, 27, 29) {real, imag} */,
  {32'h400d5673, 32'hc026498f} /* (10, 27, 28) {real, imag} */,
  {32'h3edfb491, 32'h400ea6f3} /* (10, 27, 27) {real, imag} */,
  {32'hbfb910e7, 32'hc0022ac0} /* (10, 27, 26) {real, imag} */,
  {32'hbecd0a1f, 32'h3fd1c069} /* (10, 27, 25) {real, imag} */,
  {32'hbdb5f954, 32'hbeca823a} /* (10, 27, 24) {real, imag} */,
  {32'h3fa8a679, 32'hbfd5c8b7} /* (10, 27, 23) {real, imag} */,
  {32'hc0306c38, 32'h3eae15ec} /* (10, 27, 22) {real, imag} */,
  {32'h400a9e51, 32'hbf579f57} /* (10, 27, 21) {real, imag} */,
  {32'h3eec3a8f, 32'h3f79a45c} /* (10, 27, 20) {real, imag} */,
  {32'hbe62d1f7, 32'h3f2eb232} /* (10, 27, 19) {real, imag} */,
  {32'h3f5d7d9d, 32'h3f8e4841} /* (10, 27, 18) {real, imag} */,
  {32'hbe4abd5c, 32'h3f0acda9} /* (10, 27, 17) {real, imag} */,
  {32'hc0176176, 32'h3f308956} /* (10, 27, 16) {real, imag} */,
  {32'h3eef720e, 32'hbc6c98f0} /* (10, 27, 15) {real, imag} */,
  {32'h402f1d55, 32'hbe4c1d49} /* (10, 27, 14) {real, imag} */,
  {32'h3ef8fda0, 32'h3ea71679} /* (10, 27, 13) {real, imag} */,
  {32'hbf041381, 32'hbfef5042} /* (10, 27, 12) {real, imag} */,
  {32'h3f46c98e, 32'hbfb33a22} /* (10, 27, 11) {real, imag} */,
  {32'h3f5fea57, 32'hc060811a} /* (10, 27, 10) {real, imag} */,
  {32'hbe5bb8a6, 32'h3f9e3d20} /* (10, 27, 9) {real, imag} */,
  {32'hbfe06e81, 32'h3f236fdd} /* (10, 27, 8) {real, imag} */,
  {32'h3f40a913, 32'h3f9d8f26} /* (10, 27, 7) {real, imag} */,
  {32'h3fbe3b76, 32'h403f312f} /* (10, 27, 6) {real, imag} */,
  {32'h405acb1e, 32'hbf811965} /* (10, 27, 5) {real, imag} */,
  {32'hc088d3e0, 32'hbf177fd7} /* (10, 27, 4) {real, imag} */,
  {32'h3f410bf0, 32'hc016ba7c} /* (10, 27, 3) {real, imag} */,
  {32'h3d77b14c, 32'hbf80008a} /* (10, 27, 2) {real, imag} */,
  {32'h3f6b758b, 32'h4015c892} /* (10, 27, 1) {real, imag} */,
  {32'h3fec85d7, 32'h3fd20dd2} /* (10, 27, 0) {real, imag} */,
  {32'h3dd4c029, 32'h3f6085f6} /* (10, 26, 31) {real, imag} */,
  {32'hc0491000, 32'hbfe08a85} /* (10, 26, 30) {real, imag} */,
  {32'hbe8f7632, 32'h401ed2b9} /* (10, 26, 29) {real, imag} */,
  {32'hbeb791e9, 32'h3f608e00} /* (10, 26, 28) {real, imag} */,
  {32'hc064ec50, 32'hbe858e74} /* (10, 26, 27) {real, imag} */,
  {32'h4000f523, 32'h3fce24c7} /* (10, 26, 26) {real, imag} */,
  {32'h3f3ac312, 32'hbecc5d64} /* (10, 26, 25) {real, imag} */,
  {32'h401e7779, 32'h3e68400f} /* (10, 26, 24) {real, imag} */,
  {32'hbe9ee226, 32'hbefa82b8} /* (10, 26, 23) {real, imag} */,
  {32'h3fb162ef, 32'h3fd827b6} /* (10, 26, 22) {real, imag} */,
  {32'h3f1a5631, 32'hc030481a} /* (10, 26, 21) {real, imag} */,
  {32'h3f6d067b, 32'hc083e350} /* (10, 26, 20) {real, imag} */,
  {32'h408819d9, 32'hbfd8b7eb} /* (10, 26, 19) {real, imag} */,
  {32'hbf98adf0, 32'h3f15c33d} /* (10, 26, 18) {real, imag} */,
  {32'h3fe58188, 32'h3ee165db} /* (10, 26, 17) {real, imag} */,
  {32'hbeb235c6, 32'hbe8aa72a} /* (10, 26, 16) {real, imag} */,
  {32'hbf98bd38, 32'hbdaa34ae} /* (10, 26, 15) {real, imag} */,
  {32'hbee644fc, 32'hbfc059df} /* (10, 26, 14) {real, imag} */,
  {32'h3f948627, 32'h3ec4f340} /* (10, 26, 13) {real, imag} */,
  {32'h3ff88123, 32'h3ea57da1} /* (10, 26, 12) {real, imag} */,
  {32'hbdf84f71, 32'h40350a25} /* (10, 26, 11) {real, imag} */,
  {32'h3f5f7e72, 32'h3fdb357d} /* (10, 26, 10) {real, imag} */,
  {32'hbe51b4d0, 32'h3e9d6422} /* (10, 26, 9) {real, imag} */,
  {32'hbf1db47a, 32'h3f6e34b1} /* (10, 26, 8) {real, imag} */,
  {32'h406fd052, 32'hc002e2ed} /* (10, 26, 7) {real, imag} */,
  {32'h3e0bd1a6, 32'h3d88fc34} /* (10, 26, 6) {real, imag} */,
  {32'hc02373ee, 32'hc06148fa} /* (10, 26, 5) {real, imag} */,
  {32'hc06f6833, 32'h3f348c79} /* (10, 26, 4) {real, imag} */,
  {32'h40698d26, 32'h3f0c8199} /* (10, 26, 3) {real, imag} */,
  {32'h3f071d4b, 32'hbe25a469} /* (10, 26, 2) {real, imag} */,
  {32'h3f397361, 32'hbeb409fe} /* (10, 26, 1) {real, imag} */,
  {32'h4013fb5f, 32'hc008aeaf} /* (10, 26, 0) {real, imag} */,
  {32'h40326d7c, 32'hc02f6d2a} /* (10, 25, 31) {real, imag} */,
  {32'h3f8cd5a2, 32'h3f49a274} /* (10, 25, 30) {real, imag} */,
  {32'h402cf930, 32'hbf51a532} /* (10, 25, 29) {real, imag} */,
  {32'h3e9aaa1e, 32'h3fa61775} /* (10, 25, 28) {real, imag} */,
  {32'h404ca5d4, 32'h3f9a0104} /* (10, 25, 27) {real, imag} */,
  {32'h40508566, 32'hc04623a7} /* (10, 25, 26) {real, imag} */,
  {32'h3e081cab, 32'h404b11d2} /* (10, 25, 25) {real, imag} */,
  {32'hbfc030dc, 32'hbf000bf6} /* (10, 25, 24) {real, imag} */,
  {32'hbd31ef64, 32'hc0503571} /* (10, 25, 23) {real, imag} */,
  {32'hc02f1a34, 32'h4028bc69} /* (10, 25, 22) {real, imag} */,
  {32'hbfbbb7e7, 32'h3fb41dd4} /* (10, 25, 21) {real, imag} */,
  {32'h3f828bb5, 32'h3f9b66d6} /* (10, 25, 20) {real, imag} */,
  {32'hbfaec064, 32'h3fa5d27c} /* (10, 25, 19) {real, imag} */,
  {32'h3e6a7dbe, 32'h4013e6a7} /* (10, 25, 18) {real, imag} */,
  {32'h3f096ec4, 32'hc016bc4a} /* (10, 25, 17) {real, imag} */,
  {32'hbf95f7c6, 32'hbf45dfa7} /* (10, 25, 16) {real, imag} */,
  {32'hbea2ce89, 32'h3d50dd05} /* (10, 25, 15) {real, imag} */,
  {32'h3f38b9b1, 32'h3ebca950} /* (10, 25, 14) {real, imag} */,
  {32'hc05a0d57, 32'hbf1bc88e} /* (10, 25, 13) {real, imag} */,
  {32'hbfb7f22f, 32'hbec4f9d1} /* (10, 25, 12) {real, imag} */,
  {32'hbf85dbf5, 32'h40057ce3} /* (10, 25, 11) {real, imag} */,
  {32'h3f8360ed, 32'hc037b693} /* (10, 25, 10) {real, imag} */,
  {32'hbeacb4da, 32'h3f413873} /* (10, 25, 9) {real, imag} */,
  {32'h3f6cfc47, 32'hbf0f2e5f} /* (10, 25, 8) {real, imag} */,
  {32'hbf9dc9b7, 32'h402a6680} /* (10, 25, 7) {real, imag} */,
  {32'hc05bac33, 32'hbf49cacb} /* (10, 25, 6) {real, imag} */,
  {32'h4025c10b, 32'hc04cf3ee} /* (10, 25, 5) {real, imag} */,
  {32'h3f9ba783, 32'hbdd45c8e} /* (10, 25, 4) {real, imag} */,
  {32'hc0357fb4, 32'hc02a2611} /* (10, 25, 3) {real, imag} */,
  {32'hbfb12df1, 32'hc03e8797} /* (10, 25, 2) {real, imag} */,
  {32'hbf8a3253, 32'h3f817a42} /* (10, 25, 1) {real, imag} */,
  {32'hbf8d1d77, 32'h3fb3b0c9} /* (10, 25, 0) {real, imag} */,
  {32'h40065e6c, 32'h3f32f4f8} /* (10, 24, 31) {real, imag} */,
  {32'hbfb9213d, 32'h3ff40c55} /* (10, 24, 30) {real, imag} */,
  {32'h3f74ec4f, 32'hc0588202} /* (10, 24, 29) {real, imag} */,
  {32'hbf0b399e, 32'h4004a878} /* (10, 24, 28) {real, imag} */,
  {32'h4080d1b7, 32'h4051590c} /* (10, 24, 27) {real, imag} */,
  {32'hc09d8db0, 32'hbe4bc4b2} /* (10, 24, 26) {real, imag} */,
  {32'hc00a948e, 32'hc03d4cf7} /* (10, 24, 25) {real, imag} */,
  {32'hbf506504, 32'h3d3cf415} /* (10, 24, 24) {real, imag} */,
  {32'h3f387817, 32'h3fa8c50c} /* (10, 24, 23) {real, imag} */,
  {32'hbfaa4a90, 32'h401d2aa9} /* (10, 24, 22) {real, imag} */,
  {32'hbf04c1c0, 32'hbfcbcfb1} /* (10, 24, 21) {real, imag} */,
  {32'h3ffecc15, 32'hc0446c0c} /* (10, 24, 20) {real, imag} */,
  {32'hbf048374, 32'hbfc1ad14} /* (10, 24, 19) {real, imag} */,
  {32'h3f9c2e17, 32'hbf37798e} /* (10, 24, 18) {real, imag} */,
  {32'h409c6375, 32'h3f66a685} /* (10, 24, 17) {real, imag} */,
  {32'h3eabfcf1, 32'h3e113f5e} /* (10, 24, 16) {real, imag} */,
  {32'hc08740be, 32'hbcd6e610} /* (10, 24, 15) {real, imag} */,
  {32'h3f9379ac, 32'h3e892cd5} /* (10, 24, 14) {real, imag} */,
  {32'hbfb8bdf0, 32'h3f08d211} /* (10, 24, 13) {real, imag} */,
  {32'hc0900306, 32'h3f8a4afa} /* (10, 24, 12) {real, imag} */,
  {32'h3e9effdb, 32'h3e6d104e} /* (10, 24, 11) {real, imag} */,
  {32'hbf2c8826, 32'hbf548123} /* (10, 24, 10) {real, imag} */,
  {32'h3ef3ec91, 32'h3f8489f2} /* (10, 24, 9) {real, imag} */,
  {32'h3f2d9fcb, 32'hbe585b32} /* (10, 24, 8) {real, imag} */,
  {32'h3c64bf5c, 32'h3f26692d} /* (10, 24, 7) {real, imag} */,
  {32'hc0468d62, 32'h400d91d5} /* (10, 24, 6) {real, imag} */,
  {32'hbf7960b7, 32'hc015995c} /* (10, 24, 5) {real, imag} */,
  {32'h3ec7651c, 32'hc00e0e19} /* (10, 24, 4) {real, imag} */,
  {32'h3f5945bb, 32'h4048c49a} /* (10, 24, 3) {real, imag} */,
  {32'h3efcf2a7, 32'h3f9ff7ac} /* (10, 24, 2) {real, imag} */,
  {32'hbdb00ea5, 32'hbfd8c730} /* (10, 24, 1) {real, imag} */,
  {32'hbe4daabc, 32'h3f1550c8} /* (10, 24, 0) {real, imag} */,
  {32'h3e8da07c, 32'h402dc880} /* (10, 23, 31) {real, imag} */,
  {32'hc00c5e34, 32'h3f55ac02} /* (10, 23, 30) {real, imag} */,
  {32'h3f8f0003, 32'h3f9fd23d} /* (10, 23, 29) {real, imag} */,
  {32'hbfd83886, 32'hbfc4f66b} /* (10, 23, 28) {real, imag} */,
  {32'hbfb78c08, 32'hc0056b7a} /* (10, 23, 27) {real, imag} */,
  {32'h403ebf20, 32'hbea05656} /* (10, 23, 26) {real, imag} */,
  {32'h3f6f1d77, 32'hbffab64e} /* (10, 23, 25) {real, imag} */,
  {32'hbed54421, 32'h3f425120} /* (10, 23, 24) {real, imag} */,
  {32'hc098fc29, 32'h3c984f8d} /* (10, 23, 23) {real, imag} */,
  {32'h3fab9a44, 32'h403400c9} /* (10, 23, 22) {real, imag} */,
  {32'h406342ba, 32'hbe39049e} /* (10, 23, 21) {real, imag} */,
  {32'h3fa0d68d, 32'hc099973f} /* (10, 23, 20) {real, imag} */,
  {32'hbf12ccb4, 32'h3e1f9681} /* (10, 23, 19) {real, imag} */,
  {32'h40527cca, 32'hbdb99568} /* (10, 23, 18) {real, imag} */,
  {32'h3fde932e, 32'h3f9aacc3} /* (10, 23, 17) {real, imag} */,
  {32'h3f909ec4, 32'h3fb196e3} /* (10, 23, 16) {real, imag} */,
  {32'h3f71cc1d, 32'hbf9ba667} /* (10, 23, 15) {real, imag} */,
  {32'hbf86b1df, 32'hbf3f27f9} /* (10, 23, 14) {real, imag} */,
  {32'h3fe9f564, 32'hc06a2feb} /* (10, 23, 13) {real, imag} */,
  {32'h40627641, 32'hbf073753} /* (10, 23, 12) {real, imag} */,
  {32'hc00e7109, 32'h40128e3d} /* (10, 23, 11) {real, imag} */,
  {32'hc02be764, 32'hbf3d098f} /* (10, 23, 10) {real, imag} */,
  {32'h401db943, 32'hbf4b79a5} /* (10, 23, 9) {real, imag} */,
  {32'h3ec6ecbf, 32'hbfe72567} /* (10, 23, 8) {real, imag} */,
  {32'hc038d2a0, 32'h3fc19686} /* (10, 23, 7) {real, imag} */,
  {32'hbfd9d52f, 32'hc0216461} /* (10, 23, 6) {real, imag} */,
  {32'hbf4e52bc, 32'h3fdece17} /* (10, 23, 5) {real, imag} */,
  {32'h4032cc08, 32'hbe3adfa5} /* (10, 23, 4) {real, imag} */,
  {32'h3e6f3c23, 32'h40057e98} /* (10, 23, 3) {real, imag} */,
  {32'h40049cdd, 32'hc0281c63} /* (10, 23, 2) {real, imag} */,
  {32'h3fbc5356, 32'hbf3fbf18} /* (10, 23, 1) {real, imag} */,
  {32'hbdc5d7b9, 32'hbf21c875} /* (10, 23, 0) {real, imag} */,
  {32'hbf9b5e24, 32'h3f857338} /* (10, 22, 31) {real, imag} */,
  {32'h3f7f7917, 32'hbfae51b5} /* (10, 22, 30) {real, imag} */,
  {32'hbfce7db2, 32'h3e3409f7} /* (10, 22, 29) {real, imag} */,
  {32'h3f27ca0b, 32'h3ff4a8cc} /* (10, 22, 28) {real, imag} */,
  {32'h3ecacabb, 32'hc07770ce} /* (10, 22, 27) {real, imag} */,
  {32'hbfffbaee, 32'hc0717755} /* (10, 22, 26) {real, imag} */,
  {32'h3f659cb2, 32'h40136d25} /* (10, 22, 25) {real, imag} */,
  {32'hbfb721df, 32'hc020f597} /* (10, 22, 24) {real, imag} */,
  {32'hbfd638d1, 32'h3e060543} /* (10, 22, 23) {real, imag} */,
  {32'h3f6cee8a, 32'hc0431901} /* (10, 22, 22) {real, imag} */,
  {32'h3e6a0c74, 32'hbf165948} /* (10, 22, 21) {real, imag} */,
  {32'hc0280541, 32'hbe8d4310} /* (10, 22, 20) {real, imag} */,
  {32'hc0574f0c, 32'h3f13622e} /* (10, 22, 19) {real, imag} */,
  {32'h3ffa4b8b, 32'hbf5d6290} /* (10, 22, 18) {real, imag} */,
  {32'h3e75c05d, 32'h40091486} /* (10, 22, 17) {real, imag} */,
  {32'hbed74ce8, 32'hbf6f29e2} /* (10, 22, 16) {real, imag} */,
  {32'hbf5824ad, 32'hbf93c94c} /* (10, 22, 15) {real, imag} */,
  {32'hbfad264a, 32'hbf3f5147} /* (10, 22, 14) {real, imag} */,
  {32'hc0184234, 32'hc0840420} /* (10, 22, 13) {real, imag} */,
  {32'h3eeaf063, 32'hbe6b4b8e} /* (10, 22, 12) {real, imag} */,
  {32'hc03341ba, 32'hbe846ef4} /* (10, 22, 11) {real, imag} */,
  {32'h3fafd3d6, 32'hbf36d014} /* (10, 22, 10) {real, imag} */,
  {32'h3f589ca3, 32'hbddef880} /* (10, 22, 9) {real, imag} */,
  {32'h3e8dcb9c, 32'hbfb82b5f} /* (10, 22, 8) {real, imag} */,
  {32'h3e9ef75f, 32'h3eaab9e9} /* (10, 22, 7) {real, imag} */,
  {32'hbf1554d7, 32'hbeb1ed69} /* (10, 22, 6) {real, imag} */,
  {32'h3fb7b64b, 32'hbd4cfbce} /* (10, 22, 5) {real, imag} */,
  {32'h3f9e172f, 32'h3e4de288} /* (10, 22, 4) {real, imag} */,
  {32'hbfcf910b, 32'h3fa7517f} /* (10, 22, 3) {real, imag} */,
  {32'hbfbc8167, 32'h4001126b} /* (10, 22, 2) {real, imag} */,
  {32'h3f1446b3, 32'h3e6f2783} /* (10, 22, 1) {real, imag} */,
  {32'h3f63ceb4, 32'hc01deaee} /* (10, 22, 0) {real, imag} */,
  {32'h3e289649, 32'hbf7daa8b} /* (10, 21, 31) {real, imag} */,
  {32'hbffa4807, 32'hbe18c390} /* (10, 21, 30) {real, imag} */,
  {32'h3f1dcf16, 32'h404c7f11} /* (10, 21, 29) {real, imag} */,
  {32'h3f064acc, 32'hbf73ed4e} /* (10, 21, 28) {real, imag} */,
  {32'h3f7983ee, 32'h407b681e} /* (10, 21, 27) {real, imag} */,
  {32'hc04aef3a, 32'hbfb034f2} /* (10, 21, 26) {real, imag} */,
  {32'hc02e3672, 32'hc009c9a5} /* (10, 21, 25) {real, imag} */,
  {32'hbf2795db, 32'hbf5691b3} /* (10, 21, 24) {real, imag} */,
  {32'hbf5cce10, 32'hbf0ed739} /* (10, 21, 23) {real, imag} */,
  {32'hbf7a2442, 32'h4018a46f} /* (10, 21, 22) {real, imag} */,
  {32'h3fb50009, 32'h3e9320f3} /* (10, 21, 21) {real, imag} */,
  {32'h3fcd9d13, 32'hbf82ff70} /* (10, 21, 20) {real, imag} */,
  {32'h3fdc4e16, 32'hbfeb5bbc} /* (10, 21, 19) {real, imag} */,
  {32'hbfdf5837, 32'h3fb088f3} /* (10, 21, 18) {real, imag} */,
  {32'hbe36401c, 32'hbfd21a20} /* (10, 21, 17) {real, imag} */,
  {32'h4004f973, 32'h3fe1ad41} /* (10, 21, 16) {real, imag} */,
  {32'h3f62d08e, 32'h3e0b9ab5} /* (10, 21, 15) {real, imag} */,
  {32'hc04fc2c5, 32'hbf0b5642} /* (10, 21, 14) {real, imag} */,
  {32'hbd8abfd0, 32'h405fd6dc} /* (10, 21, 13) {real, imag} */,
  {32'hc0089143, 32'h3f472ad5} /* (10, 21, 12) {real, imag} */,
  {32'h40486c1f, 32'h401e8334} /* (10, 21, 11) {real, imag} */,
  {32'hbf467d89, 32'h3d508127} /* (10, 21, 10) {real, imag} */,
  {32'h40783885, 32'hc0437a7f} /* (10, 21, 9) {real, imag} */,
  {32'hbf462883, 32'h40729b1f} /* (10, 21, 8) {real, imag} */,
  {32'h3e186e77, 32'hbf57ab68} /* (10, 21, 7) {real, imag} */,
  {32'h402f8977, 32'h406d6c58} /* (10, 21, 6) {real, imag} */,
  {32'hbfcc823a, 32'h3fecc789} /* (10, 21, 5) {real, imag} */,
  {32'hbed2ac37, 32'h3f3bc01f} /* (10, 21, 4) {real, imag} */,
  {32'h3f4bf169, 32'hbdb14f8f} /* (10, 21, 3) {real, imag} */,
  {32'h3f8551c2, 32'hbf6ed28f} /* (10, 21, 2) {real, imag} */,
  {32'hc02c6858, 32'h3fac2bb7} /* (10, 21, 1) {real, imag} */,
  {32'h40284cf8, 32'hbf9a95d5} /* (10, 21, 0) {real, imag} */,
  {32'h3fba1edb, 32'h3ecb8926} /* (10, 20, 31) {real, imag} */,
  {32'h3e0931c2, 32'hbfaddf58} /* (10, 20, 30) {real, imag} */,
  {32'hc02e109b, 32'hbfad6aba} /* (10, 20, 29) {real, imag} */,
  {32'h40118b8e, 32'hbeb41913} /* (10, 20, 28) {real, imag} */,
  {32'hbe14772a, 32'hbe31e63b} /* (10, 20, 27) {real, imag} */,
  {32'hbffb135b, 32'hbfc9daa2} /* (10, 20, 26) {real, imag} */,
  {32'h3fe97042, 32'hc039a65c} /* (10, 20, 25) {real, imag} */,
  {32'h3f825e25, 32'hbf5f90ac} /* (10, 20, 24) {real, imag} */,
  {32'h3f23c5af, 32'h3fad035c} /* (10, 20, 23) {real, imag} */,
  {32'h3f393125, 32'hbf985e93} /* (10, 20, 22) {real, imag} */,
  {32'h3f8b8680, 32'hbfac079f} /* (10, 20, 21) {real, imag} */,
  {32'hbffd0adc, 32'h3fd53e06} /* (10, 20, 20) {real, imag} */,
  {32'h3e399146, 32'h3fd4d31f} /* (10, 20, 19) {real, imag} */,
  {32'hbfb63731, 32'hbf070cfd} /* (10, 20, 18) {real, imag} */,
  {32'hbecfc8a7, 32'h3dec02d6} /* (10, 20, 17) {real, imag} */,
  {32'h40855895, 32'h3e93e847} /* (10, 20, 16) {real, imag} */,
  {32'hbf698aa2, 32'h40004dc4} /* (10, 20, 15) {real, imag} */,
  {32'h405938c7, 32'hc0524923} /* (10, 20, 14) {real, imag} */,
  {32'h3fc617bd, 32'hbe6e0644} /* (10, 20, 13) {real, imag} */,
  {32'hc0355e83, 32'h40214ae4} /* (10, 20, 12) {real, imag} */,
  {32'hbff1654a, 32'hbe1dc369} /* (10, 20, 11) {real, imag} */,
  {32'hc03ae12a, 32'h3c3674b0} /* (10, 20, 10) {real, imag} */,
  {32'hbffed559, 32'h3fcc9a1b} /* (10, 20, 9) {real, imag} */,
  {32'hbf032cec, 32'h3ff44ad0} /* (10, 20, 8) {real, imag} */,
  {32'hbfe83156, 32'h401fa420} /* (10, 20, 7) {real, imag} */,
  {32'h40411f5d, 32'hc0499e5d} /* (10, 20, 6) {real, imag} */,
  {32'h3e2be6a5, 32'hbccb9f0a} /* (10, 20, 5) {real, imag} */,
  {32'hbff22ec3, 32'hc0192e0b} /* (10, 20, 4) {real, imag} */,
  {32'hc01e2492, 32'hbe6bcfd4} /* (10, 20, 3) {real, imag} */,
  {32'h3f60f55b, 32'h3e5fdb76} /* (10, 20, 2) {real, imag} */,
  {32'hbeb1cf46, 32'h4016486b} /* (10, 20, 1) {real, imag} */,
  {32'h3f2f33c9, 32'h40013f34} /* (10, 20, 0) {real, imag} */,
  {32'hbee198f9, 32'h3f2fad6a} /* (10, 19, 31) {real, imag} */,
  {32'hbfecc115, 32'h3fc27318} /* (10, 19, 30) {real, imag} */,
  {32'h3fa878ec, 32'hbf6af79f} /* (10, 19, 29) {real, imag} */,
  {32'h405def47, 32'hbe2613cd} /* (10, 19, 28) {real, imag} */,
  {32'hc0278752, 32'h400f7318} /* (10, 19, 27) {real, imag} */,
  {32'h3fc0f12a, 32'h3eff020a} /* (10, 19, 26) {real, imag} */,
  {32'hc005b1f1, 32'h3fcd42e5} /* (10, 19, 25) {real, imag} */,
  {32'h3ed36c62, 32'h3fbc96ce} /* (10, 19, 24) {real, imag} */,
  {32'hc00fa76b, 32'hc04b008d} /* (10, 19, 23) {real, imag} */,
  {32'h4004efad, 32'hc035b7ac} /* (10, 19, 22) {real, imag} */,
  {32'h3da8b993, 32'hc063cb5f} /* (10, 19, 21) {real, imag} */,
  {32'h3f085158, 32'h3f4d4aad} /* (10, 19, 20) {real, imag} */,
  {32'hc0076683, 32'h3fb9619c} /* (10, 19, 19) {real, imag} */,
  {32'h3f65ca62, 32'h401a6031} /* (10, 19, 18) {real, imag} */,
  {32'h4032cb52, 32'hc03ede15} /* (10, 19, 17) {real, imag} */,
  {32'h40279950, 32'hbfd2ad2d} /* (10, 19, 16) {real, imag} */,
  {32'h3f7d290f, 32'h3fb4187e} /* (10, 19, 15) {real, imag} */,
  {32'h3e9fbf49, 32'h40956c56} /* (10, 19, 14) {real, imag} */,
  {32'h4002d379, 32'h402cc9c2} /* (10, 19, 13) {real, imag} */,
  {32'hbfc6d23b, 32'hbfe8bbfa} /* (10, 19, 12) {real, imag} */,
  {32'hbfc58670, 32'hbf9a3360} /* (10, 19, 11) {real, imag} */,
  {32'h3f97348e, 32'h4041c30b} /* (10, 19, 10) {real, imag} */,
  {32'hc038a006, 32'hbf5dc0fa} /* (10, 19, 9) {real, imag} */,
  {32'hbf7f9ad7, 32'h3ebec6a3} /* (10, 19, 8) {real, imag} */,
  {32'h3fa9aebd, 32'hbfc24924} /* (10, 19, 7) {real, imag} */,
  {32'h40c7f964, 32'hc017dc00} /* (10, 19, 6) {real, imag} */,
  {32'h3eb633ef, 32'h3c24c657} /* (10, 19, 5) {real, imag} */,
  {32'hbfb5b003, 32'hbf7c3998} /* (10, 19, 4) {real, imag} */,
  {32'hc01679a6, 32'h3d8613ca} /* (10, 19, 3) {real, imag} */,
  {32'h4004b533, 32'h3f8c9bfb} /* (10, 19, 2) {real, imag} */,
  {32'h3fd1b436, 32'hbbad47d0} /* (10, 19, 1) {real, imag} */,
  {32'hbf41e102, 32'hbeb281e8} /* (10, 19, 0) {real, imag} */,
  {32'hbcefd0ca, 32'hbf159e07} /* (10, 18, 31) {real, imag} */,
  {32'h3e8f5dd1, 32'h402041b4} /* (10, 18, 30) {real, imag} */,
  {32'h3cd74114, 32'hbf29f410} /* (10, 18, 29) {real, imag} */,
  {32'h3ffd8dd0, 32'hbf8059fb} /* (10, 18, 28) {real, imag} */,
  {32'h3f971738, 32'h3fa0da58} /* (10, 18, 27) {real, imag} */,
  {32'hbf83cb1f, 32'hbee828d4} /* (10, 18, 26) {real, imag} */,
  {32'h3f9f5090, 32'h3f5426e3} /* (10, 18, 25) {real, imag} */,
  {32'hbd9bead9, 32'h3f700863} /* (10, 18, 24) {real, imag} */,
  {32'h4030ee3e, 32'h3f9f7395} /* (10, 18, 23) {real, imag} */,
  {32'h3fe92726, 32'h404c156c} /* (10, 18, 22) {real, imag} */,
  {32'hbfcb1c0e, 32'hbf4871ed} /* (10, 18, 21) {real, imag} */,
  {32'hc0264530, 32'h3ff712ef} /* (10, 18, 20) {real, imag} */,
  {32'h3eaf401c, 32'h3f866adf} /* (10, 18, 19) {real, imag} */,
  {32'hc04fc6c7, 32'h3f208e8b} /* (10, 18, 18) {real, imag} */,
  {32'h3f5d6ced, 32'h3f8e23a4} /* (10, 18, 17) {real, imag} */,
  {32'hbed0f266, 32'h3f27bf67} /* (10, 18, 16) {real, imag} */,
  {32'hbf93cb52, 32'hbf534a9b} /* (10, 18, 15) {real, imag} */,
  {32'h3f89d71b, 32'h3fba489e} /* (10, 18, 14) {real, imag} */,
  {32'hbff0555c, 32'h3fa97618} /* (10, 18, 13) {real, imag} */,
  {32'h4053d01f, 32'hc0dfbb88} /* (10, 18, 12) {real, imag} */,
  {32'hbe375c40, 32'hbfac9751} /* (10, 18, 11) {real, imag} */,
  {32'h3fb965c9, 32'h403f5dd6} /* (10, 18, 10) {real, imag} */,
  {32'hbfd1e03f, 32'hbf969ed3} /* (10, 18, 9) {real, imag} */,
  {32'h3f96414a, 32'hbf479230} /* (10, 18, 8) {real, imag} */,
  {32'h3e58fddd, 32'hbf778d12} /* (10, 18, 7) {real, imag} */,
  {32'hbf66100a, 32'h3f8d6b06} /* (10, 18, 6) {real, imag} */,
  {32'h403ce435, 32'hbf9cd3d1} /* (10, 18, 5) {real, imag} */,
  {32'h3f14825b, 32'h3f73b947} /* (10, 18, 4) {real, imag} */,
  {32'h3f293cc5, 32'hbfb7be48} /* (10, 18, 3) {real, imag} */,
  {32'h3d18b048, 32'h3fdfc853} /* (10, 18, 2) {real, imag} */,
  {32'h4049e850, 32'h3e70ca74} /* (10, 18, 1) {real, imag} */,
  {32'hbf581eb2, 32'hbfff58e1} /* (10, 18, 0) {real, imag} */,
  {32'hbf3b55b7, 32'h3f3382b4} /* (10, 17, 31) {real, imag} */,
  {32'h3f1a3ee2, 32'hc0214eb4} /* (10, 17, 30) {real, imag} */,
  {32'hbe8f1427, 32'hbf87f69d} /* (10, 17, 29) {real, imag} */,
  {32'h3ee18ec0, 32'h3ec94b8d} /* (10, 17, 28) {real, imag} */,
  {32'hbf878d5d, 32'hbf62c8c4} /* (10, 17, 27) {real, imag} */,
  {32'h3ee1cddb, 32'h3f5803b9} /* (10, 17, 26) {real, imag} */,
  {32'h3f1858a7, 32'h3fbcc9cd} /* (10, 17, 25) {real, imag} */,
  {32'h3fa0af5b, 32'h3fba05b7} /* (10, 17, 24) {real, imag} */,
  {32'h4082d8bc, 32'h3906addc} /* (10, 17, 23) {real, imag} */,
  {32'hc019c248, 32'hbf35008c} /* (10, 17, 22) {real, imag} */,
  {32'hbea924a2, 32'h3e7e72c5} /* (10, 17, 21) {real, imag} */,
  {32'h3da87f80, 32'h40300052} /* (10, 17, 20) {real, imag} */,
  {32'h3fc1d80d, 32'hc0109f03} /* (10, 17, 19) {real, imag} */,
  {32'h3f6313b5, 32'hbfe84148} /* (10, 17, 18) {real, imag} */,
  {32'hbb404c97, 32'h3e1167b8} /* (10, 17, 17) {real, imag} */,
  {32'hbe40db98, 32'hbd7e20d5} /* (10, 17, 16) {real, imag} */,
  {32'h3fc7d358, 32'h3c023cf1} /* (10, 17, 15) {real, imag} */,
  {32'h403a783e, 32'hbedebe5f} /* (10, 17, 14) {real, imag} */,
  {32'h3f3499b6, 32'h3fbcdd9c} /* (10, 17, 13) {real, imag} */,
  {32'hbfa194d4, 32'hbeddd8bb} /* (10, 17, 12) {real, imag} */,
  {32'h3f480a64, 32'h3fbc894f} /* (10, 17, 11) {real, imag} */,
  {32'hc00df91a, 32'h3f9579cc} /* (10, 17, 10) {real, imag} */,
  {32'h3e81b543, 32'h3fa6cad3} /* (10, 17, 9) {real, imag} */,
  {32'hbe30a7ab, 32'hc0191dac} /* (10, 17, 8) {real, imag} */,
  {32'h3ea4589e, 32'hbf16616e} /* (10, 17, 7) {real, imag} */,
  {32'hbef5ba00, 32'hbfdb33ff} /* (10, 17, 6) {real, imag} */,
  {32'h3e92f5aa, 32'hbf716df4} /* (10, 17, 5) {real, imag} */,
  {32'hc006cc0f, 32'h403b7f18} /* (10, 17, 4) {real, imag} */,
  {32'h3ec9b51b, 32'h3f72936a} /* (10, 17, 3) {real, imag} */,
  {32'h3d9271fe, 32'hbff65b52} /* (10, 17, 2) {real, imag} */,
  {32'h3e29cc4c, 32'hbdbf4c01} /* (10, 17, 1) {real, imag} */,
  {32'h3f7396ff, 32'hbe778b79} /* (10, 17, 0) {real, imag} */,
  {32'hbfc66b06, 32'hbecf27fe} /* (10, 16, 31) {real, imag} */,
  {32'h3e2a41c9, 32'hbed262e0} /* (10, 16, 30) {real, imag} */,
  {32'hbfe257d7, 32'hbedccd64} /* (10, 16, 29) {real, imag} */,
  {32'hc017c86f, 32'hbf042e72} /* (10, 16, 28) {real, imag} */,
  {32'hbf5c280b, 32'h3fabe971} /* (10, 16, 27) {real, imag} */,
  {32'h3f8f04f7, 32'hbf6922a3} /* (10, 16, 26) {real, imag} */,
  {32'h3ecba60c, 32'h407d8069} /* (10, 16, 25) {real, imag} */,
  {32'hbf5fe327, 32'hbea943df} /* (10, 16, 24) {real, imag} */,
  {32'h401d9812, 32'hbfaa01e4} /* (10, 16, 23) {real, imag} */,
  {32'hbf567a52, 32'h3d126c80} /* (10, 16, 22) {real, imag} */,
  {32'hbffac8b5, 32'hbd1d1d02} /* (10, 16, 21) {real, imag} */,
  {32'hc0215c85, 32'h3fbe96e7} /* (10, 16, 20) {real, imag} */,
  {32'h3f6c57f6, 32'h3fa7cf1b} /* (10, 16, 19) {real, imag} */,
  {32'h3f96061f, 32'hbfad1c8a} /* (10, 16, 18) {real, imag} */,
  {32'h3f7b244a, 32'h3fdb58d2} /* (10, 16, 17) {real, imag} */,
  {32'hbf059ea7, 32'hbecdd518} /* (10, 16, 16) {real, imag} */,
  {32'h3f81560f, 32'hbfd36cf0} /* (10, 16, 15) {real, imag} */,
  {32'h3fcef83d, 32'h3fd9e69c} /* (10, 16, 14) {real, imag} */,
  {32'hbfea9ca7, 32'h3ef921a2} /* (10, 16, 13) {real, imag} */,
  {32'h3df04954, 32'h3f76c7f0} /* (10, 16, 12) {real, imag} */,
  {32'h3df1ad81, 32'h3fd37660} /* (10, 16, 11) {real, imag} */,
  {32'h3ebe931c, 32'h3bcdf030} /* (10, 16, 10) {real, imag} */,
  {32'h3f1f29db, 32'hbf402675} /* (10, 16, 9) {real, imag} */,
  {32'hbfbe304e, 32'h3fab2491} /* (10, 16, 8) {real, imag} */,
  {32'hbd066b41, 32'hbe524078} /* (10, 16, 7) {real, imag} */,
  {32'hbf1cfdd1, 32'h3f4ca268} /* (10, 16, 6) {real, imag} */,
  {32'h3f1182e9, 32'hbfa22bca} /* (10, 16, 5) {real, imag} */,
  {32'h3ff7d1b9, 32'h3f5db462} /* (10, 16, 4) {real, imag} */,
  {32'h4000fac2, 32'h3fa8919b} /* (10, 16, 3) {real, imag} */,
  {32'h3fb262c7, 32'hbf3047d8} /* (10, 16, 2) {real, imag} */,
  {32'h3fe54e1c, 32'h3f1b29c8} /* (10, 16, 1) {real, imag} */,
  {32'h3fa6465c, 32'h3e7ebe3b} /* (10, 16, 0) {real, imag} */,
  {32'hbe68475a, 32'h3f6808c5} /* (10, 15, 31) {real, imag} */,
  {32'h3f9beb90, 32'h3f588d7e} /* (10, 15, 30) {real, imag} */,
  {32'h3f9889cc, 32'h3fd7119b} /* (10, 15, 29) {real, imag} */,
  {32'hbf34e70e, 32'hbe4abf96} /* (10, 15, 28) {real, imag} */,
  {32'hbfb8e0f7, 32'hbbbb7337} /* (10, 15, 27) {real, imag} */,
  {32'hbf3f3df8, 32'hbf028c5f} /* (10, 15, 26) {real, imag} */,
  {32'h4047d1f5, 32'hc08fc273} /* (10, 15, 25) {real, imag} */,
  {32'hbdd7bc96, 32'h4035ad65} /* (10, 15, 24) {real, imag} */,
  {32'hc049fddc, 32'h3fe02144} /* (10, 15, 23) {real, imag} */,
  {32'h4046b427, 32'h3ed5f439} /* (10, 15, 22) {real, imag} */,
  {32'hbf11971e, 32'h3fa7fec8} /* (10, 15, 21) {real, imag} */,
  {32'hbd9d5b7e, 32'hc018c0f2} /* (10, 15, 20) {real, imag} */,
  {32'h3fb148d5, 32'h4099b764} /* (10, 15, 19) {real, imag} */,
  {32'h3f751aea, 32'hbfbe066c} /* (10, 15, 18) {real, imag} */,
  {32'hbea7915a, 32'hbf31af4d} /* (10, 15, 17) {real, imag} */,
  {32'h3f6d7c14, 32'h3f07fc11} /* (10, 15, 16) {real, imag} */,
  {32'hbed59b0a, 32'hbf86666b} /* (10, 15, 15) {real, imag} */,
  {32'hbfea0d2b, 32'h40771734} /* (10, 15, 14) {real, imag} */,
  {32'hbf03eee4, 32'hc05e153d} /* (10, 15, 13) {real, imag} */,
  {32'hbefa1ef7, 32'h3fb72782} /* (10, 15, 12) {real, imag} */,
  {32'h3fb457b1, 32'hc03af092} /* (10, 15, 11) {real, imag} */,
  {32'hbf4524f2, 32'h3f960b0e} /* (10, 15, 10) {real, imag} */,
  {32'h3ed865ff, 32'hc032919b} /* (10, 15, 9) {real, imag} */,
  {32'h3ea6f73c, 32'h3df9a6b5} /* (10, 15, 8) {real, imag} */,
  {32'h3f73cc44, 32'h401d1b80} /* (10, 15, 7) {real, imag} */,
  {32'hbeaa63c2, 32'h3e93182f} /* (10, 15, 6) {real, imag} */,
  {32'h4036649c, 32'h3e36b818} /* (10, 15, 5) {real, imag} */,
  {32'h3f5ade3d, 32'h3db7e922} /* (10, 15, 4) {real, imag} */,
  {32'h3e977207, 32'hbea4b5b0} /* (10, 15, 3) {real, imag} */,
  {32'h3e72fa52, 32'h3ed9ea05} /* (10, 15, 2) {real, imag} */,
  {32'hbe832cb5, 32'hbf093f3b} /* (10, 15, 1) {real, imag} */,
  {32'h3dd8349d, 32'h400dc4f1} /* (10, 15, 0) {real, imag} */,
  {32'h3e22d61d, 32'h3e9f2dcf} /* (10, 14, 31) {real, imag} */,
  {32'h3ff32c9a, 32'h3e62015e} /* (10, 14, 30) {real, imag} */,
  {32'hbfc7a4de, 32'hbf818954} /* (10, 14, 29) {real, imag} */,
  {32'h3fdb30d5, 32'h3e44ea03} /* (10, 14, 28) {real, imag} */,
  {32'h3d58adf9, 32'h400a2a74} /* (10, 14, 27) {real, imag} */,
  {32'h3f8e73bb, 32'hbfebb425} /* (10, 14, 26) {real, imag} */,
  {32'hbf8cb4c5, 32'hbfbff869} /* (10, 14, 25) {real, imag} */,
  {32'h3f08c5d7, 32'hbf2ea662} /* (10, 14, 24) {real, imag} */,
  {32'h3fc3b4fc, 32'hc02546e2} /* (10, 14, 23) {real, imag} */,
  {32'h403200da, 32'h3ed919f3} /* (10, 14, 22) {real, imag} */,
  {32'h401a7f2e, 32'h3fa4e089} /* (10, 14, 21) {real, imag} */,
  {32'h4066227c, 32'h3f8f48e3} /* (10, 14, 20) {real, imag} */,
  {32'hc00c2ab0, 32'hbe8503a9} /* (10, 14, 19) {real, imag} */,
  {32'hc00b1884, 32'hbe475150} /* (10, 14, 18) {real, imag} */,
  {32'hbf95c28d, 32'hc08676fb} /* (10, 14, 17) {real, imag} */,
  {32'h3f82cb96, 32'hbe5cde0f} /* (10, 14, 16) {real, imag} */,
  {32'hbfb1b9e4, 32'h4011b52f} /* (10, 14, 15) {real, imag} */,
  {32'hbed78420, 32'h40273fda} /* (10, 14, 14) {real, imag} */,
  {32'hbde23a87, 32'h3e8885ba} /* (10, 14, 13) {real, imag} */,
  {32'h3fff33e0, 32'h3fd8bfbd} /* (10, 14, 12) {real, imag} */,
  {32'hc01f290e, 32'hbf56e59b} /* (10, 14, 11) {real, imag} */,
  {32'h3ee19e3a, 32'hc086bf73} /* (10, 14, 10) {real, imag} */,
  {32'hc03e3c34, 32'hbf832e1c} /* (10, 14, 9) {real, imag} */,
  {32'hbe5116ca, 32'hbf6f805b} /* (10, 14, 8) {real, imag} */,
  {32'h3f130675, 32'hc00257d1} /* (10, 14, 7) {real, imag} */,
  {32'hbf0b2246, 32'hc01d9800} /* (10, 14, 6) {real, imag} */,
  {32'hbfb75ff1, 32'hbfba43eb} /* (10, 14, 5) {real, imag} */,
  {32'h3e4c821b, 32'h402ea5ae} /* (10, 14, 4) {real, imag} */,
  {32'h3fd37897, 32'hbdfe3d42} /* (10, 14, 3) {real, imag} */,
  {32'hbf9daf8a, 32'hbd0a0ddc} /* (10, 14, 2) {real, imag} */,
  {32'hc0329400, 32'h405a3e43} /* (10, 14, 1) {real, imag} */,
  {32'hbf97d98e, 32'h3fab4e52} /* (10, 14, 0) {real, imag} */,
  {32'h4004ae51, 32'hbf3f9be7} /* (10, 13, 31) {real, imag} */,
  {32'h3fd3af73, 32'hbefd121f} /* (10, 13, 30) {real, imag} */,
  {32'hc02d110b, 32'hbf6d1e9b} /* (10, 13, 29) {real, imag} */,
  {32'hbfc78914, 32'hbfe5c1af} /* (10, 13, 28) {real, imag} */,
  {32'h4000282a, 32'h3e74c5d6} /* (10, 13, 27) {real, imag} */,
  {32'h3f72e428, 32'h3fb7df88} /* (10, 13, 26) {real, imag} */,
  {32'h3fa1a393, 32'hbedba50f} /* (10, 13, 25) {real, imag} */,
  {32'hbfda1776, 32'hbb853030} /* (10, 13, 24) {real, imag} */,
  {32'h3fea6268, 32'hbf4e3788} /* (10, 13, 23) {real, imag} */,
  {32'h3e857859, 32'h3f32e44d} /* (10, 13, 22) {real, imag} */,
  {32'hbd285919, 32'hbe8a9ca0} /* (10, 13, 21) {real, imag} */,
  {32'hc03b1880, 32'h408a98a6} /* (10, 13, 20) {real, imag} */,
  {32'h400364a7, 32'h4008e64a} /* (10, 13, 19) {real, imag} */,
  {32'hc006e442, 32'h40849903} /* (10, 13, 18) {real, imag} */,
  {32'hbf1423d3, 32'h3f2e36a8} /* (10, 13, 17) {real, imag} */,
  {32'hbf8fbbb2, 32'hc07e9809} /* (10, 13, 16) {real, imag} */,
  {32'h3dce66c4, 32'h40336e9a} /* (10, 13, 15) {real, imag} */,
  {32'hbfb6f36c, 32'hbf9664ec} /* (10, 13, 14) {real, imag} */,
  {32'hbfffad27, 32'hbff7bbd1} /* (10, 13, 13) {real, imag} */,
  {32'h401876e5, 32'hbea2d722} /* (10, 13, 12) {real, imag} */,
  {32'hbf91cbe6, 32'h3fc3572c} /* (10, 13, 11) {real, imag} */,
  {32'h4049cc4a, 32'hbdbd38be} /* (10, 13, 10) {real, imag} */,
  {32'h3e8346f2, 32'h402410a2} /* (10, 13, 9) {real, imag} */,
  {32'h3f76ad13, 32'hbf0f9137} /* (10, 13, 8) {real, imag} */,
  {32'h3fbce31b, 32'h3e6e6708} /* (10, 13, 7) {real, imag} */,
  {32'h3e98da25, 32'hbd4e2d80} /* (10, 13, 6) {real, imag} */,
  {32'h3fe41b62, 32'h3fb3712c} /* (10, 13, 5) {real, imag} */,
  {32'hbf79e366, 32'h3ea8d56e} /* (10, 13, 4) {real, imag} */,
  {32'h3f1661ec, 32'h3f265447} /* (10, 13, 3) {real, imag} */,
  {32'h3f76e24d, 32'hbe885eb0} /* (10, 13, 2) {real, imag} */,
  {32'hbf4488c1, 32'hbfcd7066} /* (10, 13, 1) {real, imag} */,
  {32'h3f4a081d, 32'h403edc98} /* (10, 13, 0) {real, imag} */,
  {32'h3e988290, 32'h401f4aa8} /* (10, 12, 31) {real, imag} */,
  {32'h4024b266, 32'h3f3c231b} /* (10, 12, 30) {real, imag} */,
  {32'h3ff4b707, 32'h3f4da56b} /* (10, 12, 29) {real, imag} */,
  {32'h403e9f15, 32'hbe2d73fd} /* (10, 12, 28) {real, imag} */,
  {32'hbfcad4eb, 32'h407d7550} /* (10, 12, 27) {real, imag} */,
  {32'h3f99b4fe, 32'hbf769837} /* (10, 12, 26) {real, imag} */,
  {32'hc002d927, 32'h3c0b90af} /* (10, 12, 25) {real, imag} */,
  {32'hc03a0465, 32'hc07a8e8c} /* (10, 12, 24) {real, imag} */,
  {32'h3fb59e63, 32'h3f4618ed} /* (10, 12, 23) {real, imag} */,
  {32'hc027ac65, 32'hbe09d0d4} /* (10, 12, 22) {real, imag} */,
  {32'hc029d234, 32'h3fae9ee3} /* (10, 12, 21) {real, imag} */,
  {32'hbd861c0b, 32'h3fae976a} /* (10, 12, 20) {real, imag} */,
  {32'h4042156f, 32'hc019b692} /* (10, 12, 19) {real, imag} */,
  {32'h3fa1830c, 32'h3cb46037} /* (10, 12, 18) {real, imag} */,
  {32'h3e02a4a1, 32'hbfaaf340} /* (10, 12, 17) {real, imag} */,
  {32'hc01c6be1, 32'hbdb65edf} /* (10, 12, 16) {real, imag} */,
  {32'h3e2350f7, 32'h405df816} /* (10, 12, 15) {real, imag} */,
  {32'h40502467, 32'hbee6c891} /* (10, 12, 14) {real, imag} */,
  {32'h4028cadb, 32'hbfc4ec04} /* (10, 12, 13) {real, imag} */,
  {32'h3fa77b0e, 32'h3e231724} /* (10, 12, 12) {real, imag} */,
  {32'h3fe67047, 32'hbf317b3b} /* (10, 12, 11) {real, imag} */,
  {32'h3f0b4b5d, 32'h405cc0fc} /* (10, 12, 10) {real, imag} */,
  {32'h3ff6cbac, 32'h40485842} /* (10, 12, 9) {real, imag} */,
  {32'h3f90b405, 32'hc07e5f85} /* (10, 12, 8) {real, imag} */,
  {32'h4036ec43, 32'hc02b280a} /* (10, 12, 7) {real, imag} */,
  {32'hbfac7f26, 32'h3f148a2a} /* (10, 12, 6) {real, imag} */,
  {32'hc09d721f, 32'h40030c53} /* (10, 12, 5) {real, imag} */,
  {32'hbf62c5eb, 32'hbad7ed99} /* (10, 12, 4) {real, imag} */,
  {32'hbeaeb71e, 32'h3f25b61a} /* (10, 12, 3) {real, imag} */,
  {32'h4017bfcd, 32'hbf3c9eb6} /* (10, 12, 2) {real, imag} */,
  {32'h3e44c6bc, 32'hc0240cb1} /* (10, 12, 1) {real, imag} */,
  {32'hc046768a, 32'h3c6f38ed} /* (10, 12, 0) {real, imag} */,
  {32'hbb0215f2, 32'hc020c9c5} /* (10, 11, 31) {real, imag} */,
  {32'h3debd6a2, 32'hc0779052} /* (10, 11, 30) {real, imag} */,
  {32'h40591187, 32'h3f9b622f} /* (10, 11, 29) {real, imag} */,
  {32'h3e1fcb00, 32'hc07fa7d4} /* (10, 11, 28) {real, imag} */,
  {32'hbfc0621f, 32'hbf8df519} /* (10, 11, 27) {real, imag} */,
  {32'hbf3b14d2, 32'h4029fb7f} /* (10, 11, 26) {real, imag} */,
  {32'h3f945bcc, 32'h3ee5a884} /* (10, 11, 25) {real, imag} */,
  {32'hbff53f37, 32'h4091605e} /* (10, 11, 24) {real, imag} */,
  {32'hc01c4248, 32'h3fc7078e} /* (10, 11, 23) {real, imag} */,
  {32'hc08b41e1, 32'h406104c8} /* (10, 11, 22) {real, imag} */,
  {32'hc05fd1d6, 32'hc0377047} /* (10, 11, 21) {real, imag} */,
  {32'h3ec2faea, 32'hc04ad4c1} /* (10, 11, 20) {real, imag} */,
  {32'h3fc94751, 32'hbf6787e0} /* (10, 11, 19) {real, imag} */,
  {32'hbfb31bd0, 32'h4028e9c7} /* (10, 11, 18) {real, imag} */,
  {32'h3fb5f98c, 32'h3f803581} /* (10, 11, 17) {real, imag} */,
  {32'hbf88d3ca, 32'hc0107fa5} /* (10, 11, 16) {real, imag} */,
  {32'h3efcd476, 32'hbebb8e05} /* (10, 11, 15) {real, imag} */,
  {32'hbfb10537, 32'h3c18c3a8} /* (10, 11, 14) {real, imag} */,
  {32'h401603d0, 32'hbe6ea323} /* (10, 11, 13) {real, imag} */,
  {32'h3f1f14ee, 32'h3f14731a} /* (10, 11, 12) {real, imag} */,
  {32'hc024a0c0, 32'h401d568e} /* (10, 11, 11) {real, imag} */,
  {32'hbfbba844, 32'h3f094c9a} /* (10, 11, 10) {real, imag} */,
  {32'hbff12934, 32'h3fa8ec29} /* (10, 11, 9) {real, imag} */,
  {32'hbf0a94f4, 32'h40cf6629} /* (10, 11, 8) {real, imag} */,
  {32'hbec71054, 32'hc05183a3} /* (10, 11, 7) {real, imag} */,
  {32'h3e7d50c2, 32'hc00d7e3e} /* (10, 11, 6) {real, imag} */,
  {32'hbe30b894, 32'h405afa83} /* (10, 11, 5) {real, imag} */,
  {32'hc097ebbc, 32'hbe49f4a2} /* (10, 11, 4) {real, imag} */,
  {32'hc0648e19, 32'h3eb1ee73} /* (10, 11, 3) {real, imag} */,
  {32'h3db6850e, 32'h3e049052} /* (10, 11, 2) {real, imag} */,
  {32'hbe0a8627, 32'hc01513fa} /* (10, 11, 1) {real, imag} */,
  {32'hbfeea6fa, 32'h3f1d1e02} /* (10, 11, 0) {real, imag} */,
  {32'h3ff134e3, 32'h3fa80605} /* (10, 10, 31) {real, imag} */,
  {32'h3f847530, 32'hbe6810df} /* (10, 10, 30) {real, imag} */,
  {32'h3fa6c51c, 32'h3f85a963} /* (10, 10, 29) {real, imag} */,
  {32'hbfbbe794, 32'h3fef80c1} /* (10, 10, 28) {real, imag} */,
  {32'h3f3fec26, 32'hc0005c04} /* (10, 10, 27) {real, imag} */,
  {32'hbf8b9d5e, 32'hbf1dcdcf} /* (10, 10, 26) {real, imag} */,
  {32'h3ee7358f, 32'h3f06d111} /* (10, 10, 25) {real, imag} */,
  {32'h401e5587, 32'hbef46446} /* (10, 10, 24) {real, imag} */,
  {32'h403cf4e5, 32'hc048bf4b} /* (10, 10, 23) {real, imag} */,
  {32'h3ebd19e4, 32'h407cf4c1} /* (10, 10, 22) {real, imag} */,
  {32'h405b5f49, 32'h3d8ae73a} /* (10, 10, 21) {real, imag} */,
  {32'h3fb00f53, 32'hbff0defe} /* (10, 10, 20) {real, imag} */,
  {32'h403513c0, 32'h3fae2b69} /* (10, 10, 19) {real, imag} */,
  {32'hbf2842ca, 32'h402ecad7} /* (10, 10, 18) {real, imag} */,
  {32'h3f026efb, 32'hbfa53952} /* (10, 10, 17) {real, imag} */,
  {32'hbfbf8ccd, 32'hbe5f92c9} /* (10, 10, 16) {real, imag} */,
  {32'h402e0ac2, 32'hbf131343} /* (10, 10, 15) {real, imag} */,
  {32'h3e914caa, 32'h40349833} /* (10, 10, 14) {real, imag} */,
  {32'h3e270f30, 32'hbfc1124f} /* (10, 10, 13) {real, imag} */,
  {32'h3dd41362, 32'hbfd50f0e} /* (10, 10, 12) {real, imag} */,
  {32'h40571001, 32'hc0053009} /* (10, 10, 11) {real, imag} */,
  {32'hc054ff42, 32'hbf2bb2f5} /* (10, 10, 10) {real, imag} */,
  {32'hc029bf98, 32'hbfb9313f} /* (10, 10, 9) {real, imag} */,
  {32'hbe7dd266, 32'h3ff8d187} /* (10, 10, 8) {real, imag} */,
  {32'hbfbba98d, 32'hbf7c069e} /* (10, 10, 7) {real, imag} */,
  {32'h3fe84b95, 32'h40508d57} /* (10, 10, 6) {real, imag} */,
  {32'hbebea6cc, 32'hbf06e482} /* (10, 10, 5) {real, imag} */,
  {32'hc0122404, 32'hc06b0370} /* (10, 10, 4) {real, imag} */,
  {32'h3fd26bad, 32'h3e7154fd} /* (10, 10, 3) {real, imag} */,
  {32'h3f9e3991, 32'hbfb4eb7b} /* (10, 10, 2) {real, imag} */,
  {32'h403851c9, 32'hbfdfd941} /* (10, 10, 1) {real, imag} */,
  {32'hbf5dec20, 32'h3d30a3d1} /* (10, 10, 0) {real, imag} */,
  {32'h3f53e147, 32'h3f664910} /* (10, 9, 31) {real, imag} */,
  {32'hbff380a4, 32'h3f9df8ff} /* (10, 9, 30) {real, imag} */,
  {32'h3efc3426, 32'h40052a97} /* (10, 9, 29) {real, imag} */,
  {32'hbf1c00ec, 32'h3f3f3be7} /* (10, 9, 28) {real, imag} */,
  {32'h3febc31d, 32'h40131c6c} /* (10, 9, 27) {real, imag} */,
  {32'hbda418cb, 32'hc00bd930} /* (10, 9, 26) {real, imag} */,
  {32'h3ef0acf2, 32'hbf083041} /* (10, 9, 25) {real, imag} */,
  {32'h3f5710e3, 32'hbc89197f} /* (10, 9, 24) {real, imag} */,
  {32'hbf886543, 32'h401bb668} /* (10, 9, 23) {real, imag} */,
  {32'hbfbd7f34, 32'h406ace24} /* (10, 9, 22) {real, imag} */,
  {32'hc000c1af, 32'hbf70abb3} /* (10, 9, 21) {real, imag} */,
  {32'hc03b82f1, 32'hbf8aaff8} /* (10, 9, 20) {real, imag} */,
  {32'hbf918c27, 32'h3e8cba51} /* (10, 9, 19) {real, imag} */,
  {32'hbfd0b506, 32'h3f08f070} /* (10, 9, 18) {real, imag} */,
  {32'hbde6d90d, 32'h3fc1d743} /* (10, 9, 17) {real, imag} */,
  {32'hbe1a1bca, 32'h3fd90bd4} /* (10, 9, 16) {real, imag} */,
  {32'h3f83ac21, 32'hbdd5618e} /* (10, 9, 15) {real, imag} */,
  {32'hbf340c7a, 32'h3e390c02} /* (10, 9, 14) {real, imag} */,
  {32'hc04eebcb, 32'h3ee49202} /* (10, 9, 13) {real, imag} */,
  {32'h3f8dfe67, 32'h3df2d8e7} /* (10, 9, 12) {real, imag} */,
  {32'h3f7ce782, 32'hbfe662ad} /* (10, 9, 11) {real, imag} */,
  {32'h3f99a054, 32'hc03f56ab} /* (10, 9, 10) {real, imag} */,
  {32'h3e768ae4, 32'h4032e8b6} /* (10, 9, 9) {real, imag} */,
  {32'h40860e1a, 32'h3df5774a} /* (10, 9, 8) {real, imag} */,
  {32'h403d7fff, 32'h4063ac1d} /* (10, 9, 7) {real, imag} */,
  {32'h3f22b18a, 32'hbf8bfb21} /* (10, 9, 6) {real, imag} */,
  {32'hbeef6455, 32'h3f32a9ae} /* (10, 9, 5) {real, imag} */,
  {32'h3fb15e18, 32'h3f9d64e3} /* (10, 9, 4) {real, imag} */,
  {32'h40175395, 32'h3fd3448b} /* (10, 9, 3) {real, imag} */,
  {32'hbe822e96, 32'h40945261} /* (10, 9, 2) {real, imag} */,
  {32'hbfee8b15, 32'h4009cbf3} /* (10, 9, 1) {real, imag} */,
  {32'h3dc20707, 32'hc01e9c6c} /* (10, 9, 0) {real, imag} */,
  {32'hbec90470, 32'h3f1f56ef} /* (10, 8, 31) {real, imag} */,
  {32'hbf6f5b67, 32'h3fc883a1} /* (10, 8, 30) {real, imag} */,
  {32'hc0046efc, 32'h3f7ca0b3} /* (10, 8, 29) {real, imag} */,
  {32'hbfcd77a8, 32'hc0060ea8} /* (10, 8, 28) {real, imag} */,
  {32'h4000d970, 32'hbee01724} /* (10, 8, 27) {real, imag} */,
  {32'hc0583d9e, 32'hbf88dd28} /* (10, 8, 26) {real, imag} */,
  {32'hc039ec5d, 32'h3ecfeaaa} /* (10, 8, 25) {real, imag} */,
  {32'h3fbac5c4, 32'h3e75a383} /* (10, 8, 24) {real, imag} */,
  {32'hbe37e526, 32'h3f3b8d25} /* (10, 8, 23) {real, imag} */,
  {32'hbf96ea19, 32'hbf07baca} /* (10, 8, 22) {real, imag} */,
  {32'h3dbe2885, 32'h3fa81ef7} /* (10, 8, 21) {real, imag} */,
  {32'hc023cc80, 32'h3ff856b7} /* (10, 8, 20) {real, imag} */,
  {32'h3e39256d, 32'hbfad19be} /* (10, 8, 19) {real, imag} */,
  {32'h3fc17d9c, 32'hbf3be9d0} /* (10, 8, 18) {real, imag} */,
  {32'h3e1f6444, 32'hbfe8fba1} /* (10, 8, 17) {real, imag} */,
  {32'h3fd6669f, 32'h3fbb08fc} /* (10, 8, 16) {real, imag} */,
  {32'h3e42c791, 32'h3f989bf3} /* (10, 8, 15) {real, imag} */,
  {32'h40017313, 32'hc016d908} /* (10, 8, 14) {real, imag} */,
  {32'h3fab53d0, 32'h3fad830f} /* (10, 8, 13) {real, imag} */,
  {32'hc05b2368, 32'h3fcd1334} /* (10, 8, 12) {real, imag} */,
  {32'h4044fe80, 32'hbeae749f} /* (10, 8, 11) {real, imag} */,
  {32'hbdc9859a, 32'hbed3c894} /* (10, 8, 10) {real, imag} */,
  {32'hc01ddfe9, 32'hbfab8e98} /* (10, 8, 9) {real, imag} */,
  {32'hbed79700, 32'h405acbd7} /* (10, 8, 8) {real, imag} */,
  {32'h408bc487, 32'hbe6ea931} /* (10, 8, 7) {real, imag} */,
  {32'h404ff133, 32'h3fc06ccc} /* (10, 8, 6) {real, imag} */,
  {32'h3faaf357, 32'hc0010822} /* (10, 8, 5) {real, imag} */,
  {32'h3f3539fb, 32'h402b6639} /* (10, 8, 4) {real, imag} */,
  {32'h40459ec3, 32'hbf9926bc} /* (10, 8, 3) {real, imag} */,
  {32'hc0302b1b, 32'hbfe5a293} /* (10, 8, 2) {real, imag} */,
  {32'hbf6210f0, 32'h3fa19aa5} /* (10, 8, 1) {real, imag} */,
  {32'h407c9133, 32'hbfba31ee} /* (10, 8, 0) {real, imag} */,
  {32'hbfdfdbc3, 32'h402090f5} /* (10, 7, 31) {real, imag} */,
  {32'h3f140983, 32'h403d14ac} /* (10, 7, 30) {real, imag} */,
  {32'hbfc60fce, 32'h3f09ea20} /* (10, 7, 29) {real, imag} */,
  {32'h40332444, 32'h400bfc07} /* (10, 7, 28) {real, imag} */,
  {32'h3ff52553, 32'h401f03c3} /* (10, 7, 27) {real, imag} */,
  {32'h3f400b58, 32'hbf2ca8bc} /* (10, 7, 26) {real, imag} */,
  {32'h402b2d59, 32'hbfba38b3} /* (10, 7, 25) {real, imag} */,
  {32'h3f61500b, 32'hc086844f} /* (10, 7, 24) {real, imag} */,
  {32'h3fc5ff16, 32'hc00dce63} /* (10, 7, 23) {real, imag} */,
  {32'h3e2cc0ed, 32'hbfd1b4af} /* (10, 7, 22) {real, imag} */,
  {32'hbedbe6cd, 32'hc00b4ec1} /* (10, 7, 21) {real, imag} */,
  {32'hbf06d25b, 32'hbf4aeb29} /* (10, 7, 20) {real, imag} */,
  {32'hbf4fde3b, 32'hc0349082} /* (10, 7, 19) {real, imag} */,
  {32'h3f11209b, 32'hbe94030b} /* (10, 7, 18) {real, imag} */,
  {32'hbf27cda2, 32'h404110df} /* (10, 7, 17) {real, imag} */,
  {32'hbec8173a, 32'hc04c4e20} /* (10, 7, 16) {real, imag} */,
  {32'hc0019500, 32'h3f8a02b7} /* (10, 7, 15) {real, imag} */,
  {32'h3ec2efa4, 32'hbf84f9c9} /* (10, 7, 14) {real, imag} */,
  {32'h404475d6, 32'hbc3a4bc3} /* (10, 7, 13) {real, imag} */,
  {32'hbfac5c3a, 32'h3f791f2f} /* (10, 7, 12) {real, imag} */,
  {32'h3fabb16a, 32'h3f7e9b6f} /* (10, 7, 11) {real, imag} */,
  {32'hc00bc91e, 32'hc08307b8} /* (10, 7, 10) {real, imag} */,
  {32'h3ffdaec4, 32'hc02c0bd2} /* (10, 7, 9) {real, imag} */,
  {32'hbf8ce558, 32'hbf0e7af9} /* (10, 7, 8) {real, imag} */,
  {32'hbf536a2b, 32'h3edbca99} /* (10, 7, 7) {real, imag} */,
  {32'h3f7a8153, 32'hc03145ee} /* (10, 7, 6) {real, imag} */,
  {32'h3f4e94c5, 32'hc001bac3} /* (10, 7, 5) {real, imag} */,
  {32'h3eb7338a, 32'hbfa79e44} /* (10, 7, 4) {real, imag} */,
  {32'hbf1a48da, 32'h3fae5256} /* (10, 7, 3) {real, imag} */,
  {32'hbfc94de0, 32'hc06578ca} /* (10, 7, 2) {real, imag} */,
  {32'h3ec4bbc5, 32'hc04dbded} /* (10, 7, 1) {real, imag} */,
  {32'h3fe552dd, 32'hc000af49} /* (10, 7, 0) {real, imag} */,
  {32'h3fd36b9b, 32'hbfa1ea66} /* (10, 6, 31) {real, imag} */,
  {32'h3e1a7411, 32'h3fa01c07} /* (10, 6, 30) {real, imag} */,
  {32'hc091fbb4, 32'hbd1ba9bc} /* (10, 6, 29) {real, imag} */,
  {32'h405845be, 32'h3e13b4c9} /* (10, 6, 28) {real, imag} */,
  {32'hbeb9180f, 32'hc0476c33} /* (10, 6, 27) {real, imag} */,
  {32'hbe20dfb3, 32'hbee16a7b} /* (10, 6, 26) {real, imag} */,
  {32'h3e7a7bc1, 32'hbf0690ac} /* (10, 6, 25) {real, imag} */,
  {32'h3ea67c83, 32'h3f6df1ce} /* (10, 6, 24) {real, imag} */,
  {32'h40402f5c, 32'hc01a24c5} /* (10, 6, 23) {real, imag} */,
  {32'hbf6269f7, 32'h4095a3ca} /* (10, 6, 22) {real, imag} */,
  {32'hbdc4499d, 32'hbf021626} /* (10, 6, 21) {real, imag} */,
  {32'h3ff485bd, 32'hbdd5fe71} /* (10, 6, 20) {real, imag} */,
  {32'hbe178999, 32'h4005569d} /* (10, 6, 19) {real, imag} */,
  {32'h3d24f8b4, 32'hc04c4ad0} /* (10, 6, 18) {real, imag} */,
  {32'hbf565831, 32'h3f068e6d} /* (10, 6, 17) {real, imag} */,
  {32'hbfb81417, 32'h3e91219d} /* (10, 6, 16) {real, imag} */,
  {32'hc01d659a, 32'h400713ee} /* (10, 6, 15) {real, imag} */,
  {32'h3e1710c9, 32'h3fddae66} /* (10, 6, 14) {real, imag} */,
  {32'h3f3f5d85, 32'hc014e0af} /* (10, 6, 13) {real, imag} */,
  {32'hbe2c5411, 32'h3fe0b90b} /* (10, 6, 12) {real, imag} */,
  {32'hbd4f4668, 32'h406f1b51} /* (10, 6, 11) {real, imag} */,
  {32'hc0674205, 32'hbff88a96} /* (10, 6, 10) {real, imag} */,
  {32'hbfbd2a2d, 32'h3dd2fa33} /* (10, 6, 9) {real, imag} */,
  {32'h408aa356, 32'h3fd67756} /* (10, 6, 8) {real, imag} */,
  {32'h3f845d82, 32'hc03b74a2} /* (10, 6, 7) {real, imag} */,
  {32'h3eb3fba7, 32'h3fe28c2f} /* (10, 6, 6) {real, imag} */,
  {32'hbf8d310e, 32'hbf9b9fec} /* (10, 6, 5) {real, imag} */,
  {32'h3dd39a64, 32'h3f4cc599} /* (10, 6, 4) {real, imag} */,
  {32'h4002e242, 32'h3fa3869b} /* (10, 6, 3) {real, imag} */,
  {32'hc06ff9db, 32'hbfc66f5f} /* (10, 6, 2) {real, imag} */,
  {32'h3f4d6435, 32'h40537bfa} /* (10, 6, 1) {real, imag} */,
  {32'hc0291434, 32'hbfc0168f} /* (10, 6, 0) {real, imag} */,
  {32'hc003262f, 32'hc0a801b3} /* (10, 5, 31) {real, imag} */,
  {32'hbf29d46e, 32'h4012d480} /* (10, 5, 30) {real, imag} */,
  {32'h3ffb724c, 32'h3d1f73dd} /* (10, 5, 29) {real, imag} */,
  {32'hbf21496b, 32'hbf9af39e} /* (10, 5, 28) {real, imag} */,
  {32'hc0335a35, 32'hbf157e4c} /* (10, 5, 27) {real, imag} */,
  {32'h3ffba6f1, 32'h4017c68b} /* (10, 5, 26) {real, imag} */,
  {32'hbdadd4d1, 32'hbf074483} /* (10, 5, 25) {real, imag} */,
  {32'hbfca9484, 32'hbfc37305} /* (10, 5, 24) {real, imag} */,
  {32'h3bbd4e62, 32'h3fba76d5} /* (10, 5, 23) {real, imag} */,
  {32'hbfc9d177, 32'h40acab65} /* (10, 5, 22) {real, imag} */,
  {32'h3fa86a19, 32'hbf7b5156} /* (10, 5, 21) {real, imag} */,
  {32'hbc29e98c, 32'h3f9c3510} /* (10, 5, 20) {real, imag} */,
  {32'hbef6121f, 32'hbfcaaa27} /* (10, 5, 19) {real, imag} */,
  {32'hbef69b1d, 32'hbfd78ca4} /* (10, 5, 18) {real, imag} */,
  {32'h3fedaaa1, 32'hbe77a1f4} /* (10, 5, 17) {real, imag} */,
  {32'hbf93a3ee, 32'hbe8a5f2c} /* (10, 5, 16) {real, imag} */,
  {32'hbfc67d3d, 32'h3f7aec49} /* (10, 5, 15) {real, imag} */,
  {32'h40270950, 32'hbfaa3e2e} /* (10, 5, 14) {real, imag} */,
  {32'hc00796da, 32'hc00f4e61} /* (10, 5, 13) {real, imag} */,
  {32'h3f6551d8, 32'h3d42f0d0} /* (10, 5, 12) {real, imag} */,
  {32'hbf512710, 32'h40277dfd} /* (10, 5, 11) {real, imag} */,
  {32'hbfce1b3f, 32'hc0153e95} /* (10, 5, 10) {real, imag} */,
  {32'h3fbb4cba, 32'hbd6183bd} /* (10, 5, 9) {real, imag} */,
  {32'hbe82b86d, 32'hbfc80b81} /* (10, 5, 8) {real, imag} */,
  {32'h4074b05b, 32'h3e702a62} /* (10, 5, 7) {real, imag} */,
  {32'hbffac1ce, 32'h4025ab2e} /* (10, 5, 6) {real, imag} */,
  {32'hc034f1d3, 32'h3fe9f1c2} /* (10, 5, 5) {real, imag} */,
  {32'h3fdd0b8d, 32'hbfd65f7b} /* (10, 5, 4) {real, imag} */,
  {32'h3f34cee9, 32'hbf5e10f0} /* (10, 5, 3) {real, imag} */,
  {32'h3de1832d, 32'hbf94d869} /* (10, 5, 2) {real, imag} */,
  {32'h400aa003, 32'h405a5646} /* (10, 5, 1) {real, imag} */,
  {32'h40168054, 32'hc04c39a3} /* (10, 5, 0) {real, imag} */,
  {32'h3eeaa31d, 32'hbe416681} /* (10, 4, 31) {real, imag} */,
  {32'h405bb3d5, 32'hbdd7b80f} /* (10, 4, 30) {real, imag} */,
  {32'hc05b4105, 32'h4059fd8b} /* (10, 4, 29) {real, imag} */,
  {32'h408e6ce8, 32'h3f34f7fb} /* (10, 4, 28) {real, imag} */,
  {32'h3f750961, 32'h3fafb6f3} /* (10, 4, 27) {real, imag} */,
  {32'hbfdbff57, 32'h4001ca60} /* (10, 4, 26) {real, imag} */,
  {32'h3faaa25c, 32'h3f5ecd1e} /* (10, 4, 25) {real, imag} */,
  {32'hbf2f34a2, 32'hc093e56a} /* (10, 4, 24) {real, imag} */,
  {32'hbff391fb, 32'hc01f3d1e} /* (10, 4, 23) {real, imag} */,
  {32'hbfdb7c71, 32'hc07163c1} /* (10, 4, 22) {real, imag} */,
  {32'hbe1b9f31, 32'hbf37245d} /* (10, 4, 21) {real, imag} */,
  {32'hbf83f56f, 32'h400098c5} /* (10, 4, 20) {real, imag} */,
  {32'h3f3ddda8, 32'hc0ae73b3} /* (10, 4, 19) {real, imag} */,
  {32'h3f884887, 32'h401b23f1} /* (10, 4, 18) {real, imag} */,
  {32'h3e960f90, 32'hbe5c2d37} /* (10, 4, 17) {real, imag} */,
  {32'h3e39cf40, 32'hbea3f13c} /* (10, 4, 16) {real, imag} */,
  {32'hc019dd9c, 32'h3f4d921f} /* (10, 4, 15) {real, imag} */,
  {32'h3dc9a35f, 32'h4022921d} /* (10, 4, 14) {real, imag} */,
  {32'h3f9f9aa4, 32'hbe66976f} /* (10, 4, 13) {real, imag} */,
  {32'hbeb8f922, 32'h3fc5db16} /* (10, 4, 12) {real, imag} */,
  {32'hc0040c3e, 32'h3edccd16} /* (10, 4, 11) {real, imag} */,
  {32'h3f60b1b0, 32'h3f9f26b7} /* (10, 4, 10) {real, imag} */,
  {32'hbe5f1607, 32'hc04aa0cb} /* (10, 4, 9) {real, imag} */,
  {32'hbf8faacf, 32'hbf95eae2} /* (10, 4, 8) {real, imag} */,
  {32'hc08624e3, 32'hbffffa36} /* (10, 4, 7) {real, imag} */,
  {32'hbfcd4867, 32'h3e85733f} /* (10, 4, 6) {real, imag} */,
  {32'hbed0378e, 32'hbfd756d7} /* (10, 4, 5) {real, imag} */,
  {32'hbd80e380, 32'hc02672cf} /* (10, 4, 4) {real, imag} */,
  {32'hc029b529, 32'h402fd856} /* (10, 4, 3) {real, imag} */,
  {32'h40469f43, 32'h3fd7642a} /* (10, 4, 2) {real, imag} */,
  {32'hbf8ed19a, 32'hc09b5e6f} /* (10, 4, 1) {real, imag} */,
  {32'hc0538784, 32'hbf73d7e0} /* (10, 4, 0) {real, imag} */,
  {32'h40000009, 32'h400e55aa} /* (10, 3, 31) {real, imag} */,
  {32'h40af9652, 32'hbc97124a} /* (10, 3, 30) {real, imag} */,
  {32'h3f1a79ca, 32'hc0406fc1} /* (10, 3, 29) {real, imag} */,
  {32'h3dc65705, 32'h3fb14634} /* (10, 3, 28) {real, imag} */,
  {32'h4028e837, 32'hc0117534} /* (10, 3, 27) {real, imag} */,
  {32'hbfce0fb8, 32'h402d170c} /* (10, 3, 26) {real, imag} */,
  {32'h3f3ad48a, 32'hbe486953} /* (10, 3, 25) {real, imag} */,
  {32'h40238516, 32'h407c3593} /* (10, 3, 24) {real, imag} */,
  {32'hbf9aa05f, 32'h4034a5cc} /* (10, 3, 23) {real, imag} */,
  {32'hbfc7a916, 32'hbf04d7d8} /* (10, 3, 22) {real, imag} */,
  {32'h3f05b7de, 32'h3e1b4bab} /* (10, 3, 21) {real, imag} */,
  {32'hc05324ba, 32'h3f42dfed} /* (10, 3, 20) {real, imag} */,
  {32'h3f9d58a3, 32'h4032c67e} /* (10, 3, 19) {real, imag} */,
  {32'h3f35904d, 32'h4017409f} /* (10, 3, 18) {real, imag} */,
  {32'hbf051afc, 32'h3e179a26} /* (10, 3, 17) {real, imag} */,
  {32'hbe8ee991, 32'hbf818b18} /* (10, 3, 16) {real, imag} */,
  {32'h3e2ba2b6, 32'hbf37f8da} /* (10, 3, 15) {real, imag} */,
  {32'hbe787dfe, 32'h3f11ca2b} /* (10, 3, 14) {real, imag} */,
  {32'hbf9e48dc, 32'hbf97340c} /* (10, 3, 13) {real, imag} */,
  {32'h3ee79ed2, 32'hbf44b069} /* (10, 3, 12) {real, imag} */,
  {32'h3f922476, 32'hc0275a31} /* (10, 3, 11) {real, imag} */,
  {32'hbfbcba60, 32'h3f1bf204} /* (10, 3, 10) {real, imag} */,
  {32'hbf6c1703, 32'hbff9498d} /* (10, 3, 9) {real, imag} */,
  {32'h3f851839, 32'hbfced198} /* (10, 3, 8) {real, imag} */,
  {32'hbe342cd2, 32'hbf2859d1} /* (10, 3, 7) {real, imag} */,
  {32'h3e9ddc3a, 32'hbfe5dbbc} /* (10, 3, 6) {real, imag} */,
  {32'h3ee42af1, 32'h3baa31c3} /* (10, 3, 5) {real, imag} */,
  {32'h3f8645c3, 32'hbfcf8dbf} /* (10, 3, 4) {real, imag} */,
  {32'hbfa96f00, 32'hc02d30c0} /* (10, 3, 3) {real, imag} */,
  {32'h40738009, 32'h400f20eb} /* (10, 3, 2) {real, imag} */,
  {32'h3f0f3155, 32'h400b471e} /* (10, 3, 1) {real, imag} */,
  {32'hbf6fde3f, 32'hbeb2a3d7} /* (10, 3, 0) {real, imag} */,
  {32'h40915925, 32'h3ef604b4} /* (10, 2, 31) {real, imag} */,
  {32'hc0b49156, 32'hbea2a22d} /* (10, 2, 30) {real, imag} */,
  {32'hc01f9bef, 32'hc058b26c} /* (10, 2, 29) {real, imag} */,
  {32'h40071ddf, 32'hbffafc0c} /* (10, 2, 28) {real, imag} */,
  {32'hbf73ae5d, 32'h3ca28444} /* (10, 2, 27) {real, imag} */,
  {32'hbf2994bc, 32'hbfe0ad3e} /* (10, 2, 26) {real, imag} */,
  {32'hbe6144e5, 32'hbe8d28a0} /* (10, 2, 25) {real, imag} */,
  {32'h40ba3aa8, 32'hc00e4500} /* (10, 2, 24) {real, imag} */,
  {32'hc00242f5, 32'hbf213c4a} /* (10, 2, 23) {real, imag} */,
  {32'h40827059, 32'h401bf96a} /* (10, 2, 22) {real, imag} */,
  {32'hbd443505, 32'hbf03fc25} /* (10, 2, 21) {real, imag} */,
  {32'hbffff781, 32'h3f923027} /* (10, 2, 20) {real, imag} */,
  {32'hc01ad820, 32'h4014a858} /* (10, 2, 19) {real, imag} */,
  {32'h3fc34ac9, 32'hbf9be0c6} /* (10, 2, 18) {real, imag} */,
  {32'hc043fcb6, 32'hbe8cc3f2} /* (10, 2, 17) {real, imag} */,
  {32'h3ff26f0b, 32'hbe350b2b} /* (10, 2, 16) {real, imag} */,
  {32'h403c0e32, 32'hc00d6e43} /* (10, 2, 15) {real, imag} */,
  {32'hc048d2a2, 32'h3fae1f35} /* (10, 2, 14) {real, imag} */,
  {32'hbf1b01d4, 32'h4063094b} /* (10, 2, 13) {real, imag} */,
  {32'hbf676d5a, 32'hbf0290b1} /* (10, 2, 12) {real, imag} */,
  {32'h4009742f, 32'hc02b42d1} /* (10, 2, 11) {real, imag} */,
  {32'h3f80f979, 32'h3f612bbd} /* (10, 2, 10) {real, imag} */,
  {32'hbfc59f61, 32'hbf990dad} /* (10, 2, 9) {real, imag} */,
  {32'hbfff0db0, 32'h404a85f1} /* (10, 2, 8) {real, imag} */,
  {32'h402587cd, 32'hbfda8676} /* (10, 2, 7) {real, imag} */,
  {32'h400e869e, 32'hbf066719} /* (10, 2, 6) {real, imag} */,
  {32'hc029807c, 32'h3ed96395} /* (10, 2, 5) {real, imag} */,
  {32'h3dd03329, 32'hc03bac2a} /* (10, 2, 4) {real, imag} */,
  {32'hbfcd3a82, 32'h3ffbbccf} /* (10, 2, 3) {real, imag} */,
  {32'hc079d3ab, 32'hbd817b95} /* (10, 2, 2) {real, imag} */,
  {32'h4034da8f, 32'hbe3ca191} /* (10, 2, 1) {real, imag} */,
  {32'h3fc99a19, 32'hbeef91fa} /* (10, 2, 0) {real, imag} */,
  {32'hc0802796, 32'h4013f0bd} /* (10, 1, 31) {real, imag} */,
  {32'h403e6834, 32'h3f39062d} /* (10, 1, 30) {real, imag} */,
  {32'h3f817d9d, 32'hbff3b824} /* (10, 1, 29) {real, imag} */,
  {32'hbf889eab, 32'h4093c751} /* (10, 1, 28) {real, imag} */,
  {32'h405855a2, 32'hbffbda73} /* (10, 1, 27) {real, imag} */,
  {32'h4084dd57, 32'h407c1fac} /* (10, 1, 26) {real, imag} */,
  {32'h3f063af6, 32'hbf53f031} /* (10, 1, 25) {real, imag} */,
  {32'h3e194e06, 32'hbebb746a} /* (10, 1, 24) {real, imag} */,
  {32'hbe99f76b, 32'h3fd98705} /* (10, 1, 23) {real, imag} */,
  {32'hc033cd48, 32'h3fb0319b} /* (10, 1, 22) {real, imag} */,
  {32'h40493d46, 32'hbf2361d2} /* (10, 1, 21) {real, imag} */,
  {32'h3f99424a, 32'h3fb00233} /* (10, 1, 20) {real, imag} */,
  {32'h3fa80ee0, 32'hbddbf6c1} /* (10, 1, 19) {real, imag} */,
  {32'hbe35c250, 32'hbed4c88d} /* (10, 1, 18) {real, imag} */,
  {32'hc0026a9a, 32'hbe6843ca} /* (10, 1, 17) {real, imag} */,
  {32'hbfcedf37, 32'h3feeaf51} /* (10, 1, 16) {real, imag} */,
  {32'h3d2b31ae, 32'hc00e2cb3} /* (10, 1, 15) {real, imag} */,
  {32'h3ec112da, 32'h406d9826} /* (10, 1, 14) {real, imag} */,
  {32'hbf473146, 32'h3c998392} /* (10, 1, 13) {real, imag} */,
  {32'hbfa944f9, 32'h3e475b76} /* (10, 1, 12) {real, imag} */,
  {32'h3fe457d7, 32'h404cb76c} /* (10, 1, 11) {real, imag} */,
  {32'h3d4f296c, 32'h3ec3919a} /* (10, 1, 10) {real, imag} */,
  {32'h40091df0, 32'h3f7fc3a1} /* (10, 1, 9) {real, imag} */,
  {32'hbfdaf627, 32'h3e34f5df} /* (10, 1, 8) {real, imag} */,
  {32'h3fad3868, 32'h3f623d4c} /* (10, 1, 7) {real, imag} */,
  {32'h3fa9356a, 32'h3fdc50e6} /* (10, 1, 6) {real, imag} */,
  {32'h3ed04664, 32'hbf3cd501} /* (10, 1, 5) {real, imag} */,
  {32'hbfa75200, 32'h3fab561f} /* (10, 1, 4) {real, imag} */,
  {32'h3fff5fcc, 32'h403ae37e} /* (10, 1, 3) {real, imag} */,
  {32'h3f99d0bf, 32'hc017ac5f} /* (10, 1, 2) {real, imag} */,
  {32'hc0c6f1ad, 32'hbffb317d} /* (10, 1, 1) {real, imag} */,
  {32'hc0112cf1, 32'h3fdbcdff} /* (10, 1, 0) {real, imag} */,
  {32'hbfbcbd1b, 32'h3f806b45} /* (10, 0, 31) {real, imag} */,
  {32'hbe5d3967, 32'hbf70e9d7} /* (10, 0, 30) {real, imag} */,
  {32'hc03437b5, 32'hbff36dd0} /* (10, 0, 29) {real, imag} */,
  {32'h4063d4b2, 32'hc085e23c} /* (10, 0, 28) {real, imag} */,
  {32'h40d4245e, 32'hc02a3fa4} /* (10, 0, 27) {real, imag} */,
  {32'hc0149a7a, 32'hc09bd375} /* (10, 0, 26) {real, imag} */,
  {32'h3f8ef49a, 32'hbf4fe837} /* (10, 0, 25) {real, imag} */,
  {32'hbf3dda03, 32'h3f72551b} /* (10, 0, 24) {real, imag} */,
  {32'h40997dc7, 32'hbf1999ef} /* (10, 0, 23) {real, imag} */,
  {32'hbf575956, 32'h3fd5904c} /* (10, 0, 22) {real, imag} */,
  {32'h40051461, 32'hbfb514d9} /* (10, 0, 21) {real, imag} */,
  {32'h401b723c, 32'h3eee5e66} /* (10, 0, 20) {real, imag} */,
  {32'hbfd6e878, 32'hc00ad271} /* (10, 0, 19) {real, imag} */,
  {32'hbf33dc51, 32'hbea843ae} /* (10, 0, 18) {real, imag} */,
  {32'h3f07571a, 32'hbfe5bd17} /* (10, 0, 17) {real, imag} */,
  {32'h3fc00d36, 32'h4044a113} /* (10, 0, 16) {real, imag} */,
  {32'h3f678b61, 32'h3f5e8391} /* (10, 0, 15) {real, imag} */,
  {32'hbf1740a7, 32'hbfbdc252} /* (10, 0, 14) {real, imag} */,
  {32'h3eae4200, 32'h402339b0} /* (10, 0, 13) {real, imag} */,
  {32'h3e9c74e4, 32'hbfaf3677} /* (10, 0, 12) {real, imag} */,
  {32'hbe40b3cb, 32'hc03ad638} /* (10, 0, 11) {real, imag} */,
  {32'hbea95f87, 32'h3edb4452} /* (10, 0, 10) {real, imag} */,
  {32'h404915c8, 32'h403db2fe} /* (10, 0, 9) {real, imag} */,
  {32'hc06e9456, 32'h3ffc3910} /* (10, 0, 8) {real, imag} */,
  {32'hc0020cfb, 32'h406247bd} /* (10, 0, 7) {real, imag} */,
  {32'h3eeb14b2, 32'h3e30681d} /* (10, 0, 6) {real, imag} */,
  {32'hbf76bfa4, 32'h4022768b} /* (10, 0, 5) {real, imag} */,
  {32'hbec3296a, 32'h3cdea6b0} /* (10, 0, 4) {real, imag} */,
  {32'hc0a20d8b, 32'hbe95d545} /* (10, 0, 3) {real, imag} */,
  {32'h3fe19ba9, 32'hc041b0e9} /* (10, 0, 2) {real, imag} */,
  {32'hc06c4dbd, 32'hc0690ed4} /* (10, 0, 1) {real, imag} */,
  {32'hbfa85644, 32'hbfa639ca} /* (10, 0, 0) {real, imag} */,
  {32'hc0531de6, 32'h40d21818} /* (9, 31, 31) {real, imag} */,
  {32'hbf4e8aea, 32'hc08cc193} /* (9, 31, 30) {real, imag} */,
  {32'hbfbc6c65, 32'h3ea5f303} /* (9, 31, 29) {real, imag} */,
  {32'hbf3046d0, 32'h402de475} /* (9, 31, 28) {real, imag} */,
  {32'h3fd653dd, 32'h3f267a08} /* (9, 31, 27) {real, imag} */,
  {32'hbf9d96ac, 32'h3f208883} /* (9, 31, 26) {real, imag} */,
  {32'h400728c1, 32'hbf5392f9} /* (9, 31, 25) {real, imag} */,
  {32'hbf955d41, 32'hc0774128} /* (9, 31, 24) {real, imag} */,
  {32'hbf2dfccb, 32'h40599e8a} /* (9, 31, 23) {real, imag} */,
  {32'hbf6ac2d7, 32'h3fed6f8f} /* (9, 31, 22) {real, imag} */,
  {32'h4015d8fd, 32'hc006ea8c} /* (9, 31, 21) {real, imag} */,
  {32'h3f28e0d2, 32'hc000a2bd} /* (9, 31, 20) {real, imag} */,
  {32'hbf590bab, 32'h3f2b8d53} /* (9, 31, 19) {real, imag} */,
  {32'hc02cc534, 32'hbfdb6b0c} /* (9, 31, 18) {real, imag} */,
  {32'hbcba9dde, 32'hbef7415e} /* (9, 31, 17) {real, imag} */,
  {32'h40072a6f, 32'h3fb77283} /* (9, 31, 16) {real, imag} */,
  {32'h3ff247b3, 32'hc00469b1} /* (9, 31, 15) {real, imag} */,
  {32'h3fa4b829, 32'hbf7a87c1} /* (9, 31, 14) {real, imag} */,
  {32'hbfd90c67, 32'hbfbf1f68} /* (9, 31, 13) {real, imag} */,
  {32'h401ef282, 32'h3eac95e9} /* (9, 31, 12) {real, imag} */,
  {32'h405c0c4a, 32'h3f86dbe6} /* (9, 31, 11) {real, imag} */,
  {32'h3f1bbd10, 32'h3e770cb3} /* (9, 31, 10) {real, imag} */,
  {32'h3f81418c, 32'hbfff66be} /* (9, 31, 9) {real, imag} */,
  {32'hbf9d6ecb, 32'hbfaeb2e4} /* (9, 31, 8) {real, imag} */,
  {32'h3fc8e050, 32'h3fe14e42} /* (9, 31, 7) {real, imag} */,
  {32'h3f08902e, 32'hbdbeb6aa} /* (9, 31, 6) {real, imag} */,
  {32'h3fa9ecda, 32'hbfcadf11} /* (9, 31, 5) {real, imag} */,
  {32'hbfde0a13, 32'h3fbca16b} /* (9, 31, 4) {real, imag} */,
  {32'h402ca188, 32'h4019ac45} /* (9, 31, 3) {real, imag} */,
  {32'hbee0795d, 32'h3f853feb} /* (9, 31, 2) {real, imag} */,
  {32'hc02ed7e0, 32'h40750b3d} /* (9, 31, 1) {real, imag} */,
  {32'hc093381e, 32'h4099176f} /* (9, 31, 0) {real, imag} */,
  {32'h408ad91b, 32'h40197944} /* (9, 30, 31) {real, imag} */,
  {32'hbfee7678, 32'h40bc1e31} /* (9, 30, 30) {real, imag} */,
  {32'h3fa5be0e, 32'hc05bbdbd} /* (9, 30, 29) {real, imag} */,
  {32'hbff79f84, 32'hbfe1747a} /* (9, 30, 28) {real, imag} */,
  {32'hbe2fd68f, 32'hc04735e4} /* (9, 30, 27) {real, imag} */,
  {32'hbf58da36, 32'hbfa7ab98} /* (9, 30, 26) {real, imag} */,
  {32'h402c6be5, 32'hbf931256} /* (9, 30, 25) {real, imag} */,
  {32'h3fbef27b, 32'h409bd6bb} /* (9, 30, 24) {real, imag} */,
  {32'h3fd2fb1f, 32'h3faa02f2} /* (9, 30, 23) {real, imag} */,
  {32'hbfedcadc, 32'h40001d24} /* (9, 30, 22) {real, imag} */,
  {32'h3f434c88, 32'h403e2f77} /* (9, 30, 21) {real, imag} */,
  {32'h3e487ff3, 32'h3fed3350} /* (9, 30, 20) {real, imag} */,
  {32'hbfe4052e, 32'hc00a3a2b} /* (9, 30, 19) {real, imag} */,
  {32'hbf2b0188, 32'hbf22503b} /* (9, 30, 18) {real, imag} */,
  {32'h3f654553, 32'h3f0d3a26} /* (9, 30, 17) {real, imag} */,
  {32'hbf5fb73e, 32'hbe3162d7} /* (9, 30, 16) {real, imag} */,
  {32'h3e6e4797, 32'hbfc307e8} /* (9, 30, 15) {real, imag} */,
  {32'hbef59f1d, 32'hc018d31e} /* (9, 30, 14) {real, imag} */,
  {32'h4015b910, 32'h3e3cba08} /* (9, 30, 13) {real, imag} */,
  {32'hbe3487a6, 32'h402bae58} /* (9, 30, 12) {real, imag} */,
  {32'hbf1bad4e, 32'h40845108} /* (9, 30, 11) {real, imag} */,
  {32'h3fc2cf91, 32'hc0425139} /* (9, 30, 10) {real, imag} */,
  {32'h3f0c1eb8, 32'h3fb22a83} /* (9, 30, 9) {real, imag} */,
  {32'hbfdaa068, 32'hc01bf77f} /* (9, 30, 8) {real, imag} */,
  {32'h3e94fbfb, 32'hc07d0d32} /* (9, 30, 7) {real, imag} */,
  {32'hc097bbd2, 32'h400ea312} /* (9, 30, 6) {real, imag} */,
  {32'hbee34bb2, 32'hbfd7287d} /* (9, 30, 5) {real, imag} */,
  {32'h403edb13, 32'h3ce35992} /* (9, 30, 4) {real, imag} */,
  {32'hc09df5cb, 32'h400d7d4f} /* (9, 30, 3) {real, imag} */,
  {32'hc06140ec, 32'h404f6867} /* (9, 30, 2) {real, imag} */,
  {32'h408f90bc, 32'hc02b0af6} /* (9, 30, 1) {real, imag} */,
  {32'hbdd16f89, 32'hc013ae42} /* (9, 30, 0) {real, imag} */,
  {32'hbec1e0fc, 32'h405dfdc6} /* (9, 29, 31) {real, imag} */,
  {32'hc09e6758, 32'hc09d48f0} /* (9, 29, 30) {real, imag} */,
  {32'h403ccb35, 32'h40249750} /* (9, 29, 29) {real, imag} */,
  {32'h3de40bdd, 32'h3fcbf35c} /* (9, 29, 28) {real, imag} */,
  {32'h3f96a2ce, 32'h402493ed} /* (9, 29, 27) {real, imag} */,
  {32'hbf7f1795, 32'h3f84befc} /* (9, 29, 26) {real, imag} */,
  {32'h3fa62fdd, 32'h3f852626} /* (9, 29, 25) {real, imag} */,
  {32'hbc6f985d, 32'h40136166} /* (9, 29, 24) {real, imag} */,
  {32'h3f97ff0b, 32'h3fbce95a} /* (9, 29, 23) {real, imag} */,
  {32'h4008887d, 32'hbfe2fdb6} /* (9, 29, 22) {real, imag} */,
  {32'hbfee4223, 32'h401d67cf} /* (9, 29, 21) {real, imag} */,
  {32'hc0078891, 32'hc07b7b3d} /* (9, 29, 20) {real, imag} */,
  {32'hbfbc172f, 32'hbfb2a52c} /* (9, 29, 19) {real, imag} */,
  {32'h3f309dfa, 32'h3fa4ffff} /* (9, 29, 18) {real, imag} */,
  {32'hbec1a5c6, 32'h3f3ddf20} /* (9, 29, 17) {real, imag} */,
  {32'hbf1d80fc, 32'hbe65b04e} /* (9, 29, 16) {real, imag} */,
  {32'hc0077093, 32'hbf8889e3} /* (9, 29, 15) {real, imag} */,
  {32'h3f8274b4, 32'h3ef21d7b} /* (9, 29, 14) {real, imag} */,
  {32'h3f28be6b, 32'h4018d869} /* (9, 29, 13) {real, imag} */,
  {32'h3fcdc884, 32'hc007cfd5} /* (9, 29, 12) {real, imag} */,
  {32'hbf89d165, 32'h3e3b2e3c} /* (9, 29, 11) {real, imag} */,
  {32'h4058a784, 32'h3f254ad2} /* (9, 29, 10) {real, imag} */,
  {32'hbf24d7d3, 32'hbf85b729} /* (9, 29, 9) {real, imag} */,
  {32'h400bf5e6, 32'hc0194128} /* (9, 29, 8) {real, imag} */,
  {32'hbf46b213, 32'h3f817bbd} /* (9, 29, 7) {real, imag} */,
  {32'h3eda0eaf, 32'h3fcc3e98} /* (9, 29, 6) {real, imag} */,
  {32'h404344ef, 32'h40167f9a} /* (9, 29, 5) {real, imag} */,
  {32'hc030707e, 32'h3f73d795} /* (9, 29, 4) {real, imag} */,
  {32'hbe0b221e, 32'h3f727172} /* (9, 29, 3) {real, imag} */,
  {32'hc09f517d, 32'hc0453953} /* (9, 29, 2) {real, imag} */,
  {32'hbce755bc, 32'hc094a05e} /* (9, 29, 1) {real, imag} */,
  {32'hbdb38734, 32'h40193730} /* (9, 29, 0) {real, imag} */,
  {32'h3f9efcdf, 32'hbfe404c9} /* (9, 28, 31) {real, imag} */,
  {32'hbfd258e9, 32'h3f8d221d} /* (9, 28, 30) {real, imag} */,
  {32'hbf05f2ae, 32'h401c08ec} /* (9, 28, 29) {real, imag} */,
  {32'h400956fc, 32'hbe624fd6} /* (9, 28, 28) {real, imag} */,
  {32'h4020bb48, 32'hc01d47e5} /* (9, 28, 27) {real, imag} */,
  {32'h4042c4d5, 32'hc060c04e} /* (9, 28, 26) {real, imag} */,
  {32'hbf46b170, 32'hbffc6676} /* (9, 28, 25) {real, imag} */,
  {32'h405b6b6c, 32'hc0012418} /* (9, 28, 24) {real, imag} */,
  {32'h3fd440ce, 32'h3fd15940} /* (9, 28, 23) {real, imag} */,
  {32'h3fef7dc5, 32'h3ee6c5dd} /* (9, 28, 22) {real, imag} */,
  {32'h3e08f994, 32'hbfb637be} /* (9, 28, 21) {real, imag} */,
  {32'h404b34b5, 32'h40185780} /* (9, 28, 20) {real, imag} */,
  {32'hbfde4275, 32'h3ff40104} /* (9, 28, 19) {real, imag} */,
  {32'hbf773e55, 32'h40090f2e} /* (9, 28, 18) {real, imag} */,
  {32'hbfa3929b, 32'hbe513591} /* (9, 28, 17) {real, imag} */,
  {32'h3fb58293, 32'h3fc95495} /* (9, 28, 16) {real, imag} */,
  {32'h3ea556e7, 32'hbfbbf704} /* (9, 28, 15) {real, imag} */,
  {32'h3fe4e549, 32'h40512365} /* (9, 28, 14) {real, imag} */,
  {32'hbfb8d9d0, 32'hbfdce455} /* (9, 28, 13) {real, imag} */,
  {32'hbeb72828, 32'hbf0a0cbf} /* (9, 28, 12) {real, imag} */,
  {32'hbf683337, 32'h3f9d763e} /* (9, 28, 11) {real, imag} */,
  {32'hbf8c48f6, 32'hbfe888de} /* (9, 28, 10) {real, imag} */,
  {32'hbfe34b7d, 32'h3f4054e2} /* (9, 28, 9) {real, imag} */,
  {32'hc0c66462, 32'hbfe44d79} /* (9, 28, 8) {real, imag} */,
  {32'h3f5e2984, 32'hbfbf2f29} /* (9, 28, 7) {real, imag} */,
  {32'h3fb1680f, 32'h3f6e504b} /* (9, 28, 6) {real, imag} */,
  {32'hbf9cbc63, 32'hbffc5bbb} /* (9, 28, 5) {real, imag} */,
  {32'hbfac0f31, 32'h3eb87404} /* (9, 28, 4) {real, imag} */,
  {32'hc00fbf40, 32'h40152154} /* (9, 28, 3) {real, imag} */,
  {32'hbfd64f74, 32'hc04acf98} /* (9, 28, 2) {real, imag} */,
  {32'h3ff9d852, 32'h405b0d7a} /* (9, 28, 1) {real, imag} */,
  {32'h3f7446d4, 32'hc05a4495} /* (9, 28, 0) {real, imag} */,
  {32'h4014e92a, 32'hc083a0a6} /* (9, 27, 31) {real, imag} */,
  {32'hc0134480, 32'h3ff8d91e} /* (9, 27, 30) {real, imag} */,
  {32'h4028f603, 32'hbf87f3bc} /* (9, 27, 29) {real, imag} */,
  {32'h3f2f2128, 32'hbfd9c576} /* (9, 27, 28) {real, imag} */,
  {32'h3f911d87, 32'h3e87af9a} /* (9, 27, 27) {real, imag} */,
  {32'hc00d0095, 32'h404e5e9a} /* (9, 27, 26) {real, imag} */,
  {32'h400dce51, 32'hc083d6fc} /* (9, 27, 25) {real, imag} */,
  {32'hbf73bd75, 32'hc030d6dd} /* (9, 27, 24) {real, imag} */,
  {32'hbfbbcb26, 32'h40747a1f} /* (9, 27, 23) {real, imag} */,
  {32'h3d6dd515, 32'h40879e88} /* (9, 27, 22) {real, imag} */,
  {32'h3e9905ed, 32'h401b70c5} /* (9, 27, 21) {real, imag} */,
  {32'hc07eacf1, 32'hbd8144e1} /* (9, 27, 20) {real, imag} */,
  {32'h3dcbfa2b, 32'h3f82425d} /* (9, 27, 19) {real, imag} */,
  {32'h3e18e900, 32'hbf70cfa7} /* (9, 27, 18) {real, imag} */,
  {32'h3f8410d5, 32'hbfd8356c} /* (9, 27, 17) {real, imag} */,
  {32'hbfa470bf, 32'h3f9b8a6f} /* (9, 27, 16) {real, imag} */,
  {32'hbd938016, 32'h3e36bf1d} /* (9, 27, 15) {real, imag} */,
  {32'hbff3e4c3, 32'hc0130e1d} /* (9, 27, 14) {real, imag} */,
  {32'hbf1195b1, 32'hbf98c398} /* (9, 27, 13) {real, imag} */,
  {32'h3f8f2c34, 32'hbedcf1bb} /* (9, 27, 12) {real, imag} */,
  {32'hbff186a7, 32'hbf0e3c3b} /* (9, 27, 11) {real, imag} */,
  {32'h3fd5d054, 32'hc07bde98} /* (9, 27, 10) {real, imag} */,
  {32'h4035f7bb, 32'h40540a45} /* (9, 27, 9) {real, imag} */,
  {32'h4053f79e, 32'h403ffdea} /* (9, 27, 8) {real, imag} */,
  {32'h4014d275, 32'h3e31bc41} /* (9, 27, 7) {real, imag} */,
  {32'hbfc12cd1, 32'h40442ec8} /* (9, 27, 6) {real, imag} */,
  {32'h3cd5fa22, 32'h401bbe9c} /* (9, 27, 5) {real, imag} */,
  {32'hbec02ca0, 32'hbf4dc756} /* (9, 27, 4) {real, imag} */,
  {32'hc048f778, 32'h3fc94b3c} /* (9, 27, 3) {real, imag} */,
  {32'h3ffa48b2, 32'h40035df3} /* (9, 27, 2) {real, imag} */,
  {32'hbf9de27b, 32'hbfc31c7a} /* (9, 27, 1) {real, imag} */,
  {32'h3f676323, 32'h3faf8a11} /* (9, 27, 0) {real, imag} */,
  {32'hc02a1e1a, 32'hc03d1472} /* (9, 26, 31) {real, imag} */,
  {32'h3fee28c9, 32'hbf557e14} /* (9, 26, 30) {real, imag} */,
  {32'h400d0a80, 32'hc0d78fc9} /* (9, 26, 29) {real, imag} */,
  {32'h401a6caa, 32'h3e4f9e07} /* (9, 26, 28) {real, imag} */,
  {32'hbfb7a40d, 32'h3f28a956} /* (9, 26, 27) {real, imag} */,
  {32'h3f08b514, 32'hbf919d0d} /* (9, 26, 26) {real, imag} */,
  {32'h3f9ca35a, 32'hbd0752c0} /* (9, 26, 25) {real, imag} */,
  {32'hbece8a1b, 32'h3fba09f3} /* (9, 26, 24) {real, imag} */,
  {32'h402e7d63, 32'h3ff530fd} /* (9, 26, 23) {real, imag} */,
  {32'hbdf9e090, 32'hc00dadb4} /* (9, 26, 22) {real, imag} */,
  {32'h3e97a5bf, 32'h4081cc98} /* (9, 26, 21) {real, imag} */,
  {32'hbfda9ead, 32'hc044332f} /* (9, 26, 20) {real, imag} */,
  {32'hbf48a343, 32'hbf583406} /* (9, 26, 19) {real, imag} */,
  {32'hc02de3dd, 32'hc0105eb9} /* (9, 26, 18) {real, imag} */,
  {32'hbfe40a5c, 32'h3e51ebab} /* (9, 26, 17) {real, imag} */,
  {32'hbf92ae04, 32'hbfd1604a} /* (9, 26, 16) {real, imag} */,
  {32'h40819090, 32'hbfdd5e2b} /* (9, 26, 15) {real, imag} */,
  {32'hbeb1b596, 32'hbf5c1aaa} /* (9, 26, 14) {real, imag} */,
  {32'hbf0e2e2d, 32'h3e5ac6fa} /* (9, 26, 13) {real, imag} */,
  {32'h3fbaceb2, 32'h3f9ddd93} /* (9, 26, 12) {real, imag} */,
  {32'h3f3f7223, 32'h400d4ab6} /* (9, 26, 11) {real, imag} */,
  {32'hc06d250d, 32'hc0a3f5cb} /* (9, 26, 10) {real, imag} */,
  {32'h3fb77d9a, 32'h3c5744c2} /* (9, 26, 9) {real, imag} */,
  {32'hbf16c3fa, 32'hc032b249} /* (9, 26, 8) {real, imag} */,
  {32'h3f100527, 32'h40105218} /* (9, 26, 7) {real, imag} */,
  {32'hc00de6a8, 32'h40131a71} /* (9, 26, 6) {real, imag} */,
  {32'hc06a8daa, 32'h3f1cbdf5} /* (9, 26, 5) {real, imag} */,
  {32'h3fffae94, 32'h4042ea0d} /* (9, 26, 4) {real, imag} */,
  {32'hc0463b53, 32'hbea7aff5} /* (9, 26, 3) {real, imag} */,
  {32'hbf834d4a, 32'h3ea9387b} /* (9, 26, 2) {real, imag} */,
  {32'h403f89fc, 32'h3f29586e} /* (9, 26, 1) {real, imag} */,
  {32'hc0098b8a, 32'hbebb9601} /* (9, 26, 0) {real, imag} */,
  {32'h3fed628e, 32'hbf9bba7c} /* (9, 25, 31) {real, imag} */,
  {32'h3e6e2442, 32'hc0589349} /* (9, 25, 30) {real, imag} */,
  {32'hbd97f52c, 32'h3e541a1f} /* (9, 25, 29) {real, imag} */,
  {32'h3f742777, 32'h3f87ed14} /* (9, 25, 28) {real, imag} */,
  {32'hbfaf3161, 32'h4035d11a} /* (9, 25, 27) {real, imag} */,
  {32'hc041fd3a, 32'h3fa65901} /* (9, 25, 26) {real, imag} */,
  {32'hbf662aa7, 32'h3f24eb19} /* (9, 25, 25) {real, imag} */,
  {32'h3fe3a70e, 32'hbf4a54fd} /* (9, 25, 24) {real, imag} */,
  {32'hc001eeb9, 32'h3eadd4fd} /* (9, 25, 23) {real, imag} */,
  {32'hc02bcd7e, 32'h4049a94a} /* (9, 25, 22) {real, imag} */,
  {32'hc0188327, 32'hc02ad367} /* (9, 25, 21) {real, imag} */,
  {32'hbc8f7591, 32'h3decb28e} /* (9, 25, 20) {real, imag} */,
  {32'hbfc67561, 32'hc03834b8} /* (9, 25, 19) {real, imag} */,
  {32'h3fd79863, 32'h3f22c321} /* (9, 25, 18) {real, imag} */,
  {32'h4006f098, 32'h3fc29936} /* (9, 25, 17) {real, imag} */,
  {32'h3f707ebb, 32'hbface86e} /* (9, 25, 16) {real, imag} */,
  {32'hbf874103, 32'h3ebafe79} /* (9, 25, 15) {real, imag} */,
  {32'h3efae09f, 32'hbfb4ea30} /* (9, 25, 14) {real, imag} */,
  {32'h3ec82e1b, 32'hbfca3be6} /* (9, 25, 13) {real, imag} */,
  {32'hbf5205ad, 32'hbf27ec5b} /* (9, 25, 12) {real, imag} */,
  {32'hbff649d3, 32'hbedd740f} /* (9, 25, 11) {real, imag} */,
  {32'hc05aca0d, 32'h400f3a38} /* (9, 25, 10) {real, imag} */,
  {32'hbfe84857, 32'h3fd512fc} /* (9, 25, 9) {real, imag} */,
  {32'h400853da, 32'h3ff04667} /* (9, 25, 8) {real, imag} */,
  {32'h3f528d4f, 32'h3fc15caa} /* (9, 25, 7) {real, imag} */,
  {32'hc03d0d7f, 32'h3e1b07a4} /* (9, 25, 6) {real, imag} */,
  {32'h40908d43, 32'hc0c27e3e} /* (9, 25, 5) {real, imag} */,
  {32'h3f9e123a, 32'hbf923749} /* (9, 25, 4) {real, imag} */,
  {32'h3fd8e17f, 32'hbfe8727b} /* (9, 25, 3) {real, imag} */,
  {32'h3f0877c1, 32'hbfb91dd1} /* (9, 25, 2) {real, imag} */,
  {32'h3fb713a0, 32'h40a1ee17} /* (9, 25, 1) {real, imag} */,
  {32'h3f6e7c90, 32'hbf16876e} /* (9, 25, 0) {real, imag} */,
  {32'h3dd85674, 32'h4029c27e} /* (9, 24, 31) {real, imag} */,
  {32'hbfe24b2f, 32'h3fac7aef} /* (9, 24, 30) {real, imag} */,
  {32'hbf7f2d6f, 32'hbf9094ee} /* (9, 24, 29) {real, imag} */,
  {32'hbf84fdaa, 32'h3fe8a16f} /* (9, 24, 28) {real, imag} */,
  {32'h3fd11c06, 32'hc076648b} /* (9, 24, 27) {real, imag} */,
  {32'hbfea674e, 32'hbffceb00} /* (9, 24, 26) {real, imag} */,
  {32'hbfd68c5a, 32'h4019493f} /* (9, 24, 25) {real, imag} */,
  {32'h40367a95, 32'hbf1f855b} /* (9, 24, 24) {real, imag} */,
  {32'hbf85efbb, 32'hbf49239d} /* (9, 24, 23) {real, imag} */,
  {32'h3ed70fd4, 32'hc01856b6} /* (9, 24, 22) {real, imag} */,
  {32'h3e1c3da9, 32'hbf1fa28c} /* (9, 24, 21) {real, imag} */,
  {32'hbe5bb8cd, 32'h403d69b2} /* (9, 24, 20) {real, imag} */,
  {32'h3f8b7dfb, 32'h3f948bee} /* (9, 24, 19) {real, imag} */,
  {32'h4048f626, 32'hbf05f913} /* (9, 24, 18) {real, imag} */,
  {32'hbf295758, 32'hbca484f6} /* (9, 24, 17) {real, imag} */,
  {32'hbf1b962a, 32'h4016872c} /* (9, 24, 16) {real, imag} */,
  {32'hbf42a106, 32'hc01b22cc} /* (9, 24, 15) {real, imag} */,
  {32'h3fd88c23, 32'h3f6bb7b5} /* (9, 24, 14) {real, imag} */,
  {32'h3fe0590e, 32'h4082850f} /* (9, 24, 13) {real, imag} */,
  {32'hbd220ae9, 32'hc0574af5} /* (9, 24, 12) {real, imag} */,
  {32'hbd3efb09, 32'hc062cbbe} /* (9, 24, 11) {real, imag} */,
  {32'h40437c57, 32'hbec45884} /* (9, 24, 10) {real, imag} */,
  {32'h3fab9d3e, 32'h3fd96774} /* (9, 24, 9) {real, imag} */,
  {32'hbfcdc65f, 32'h401712b5} /* (9, 24, 8) {real, imag} */,
  {32'hbe9e522a, 32'h3f91292e} /* (9, 24, 7) {real, imag} */,
  {32'hbe9cd8b4, 32'h3e7cd07b} /* (9, 24, 6) {real, imag} */,
  {32'h3ec28791, 32'h404089b7} /* (9, 24, 5) {real, imag} */,
  {32'h405d6cd9, 32'hbf55921d} /* (9, 24, 4) {real, imag} */,
  {32'hbf0b37d3, 32'hbf30f12f} /* (9, 24, 3) {real, imag} */,
  {32'hbeea31c8, 32'h401c2275} /* (9, 24, 2) {real, imag} */,
  {32'h3f5aea9f, 32'hbed4987a} /* (9, 24, 1) {real, imag} */,
  {32'hbf7a4474, 32'hc040d217} /* (9, 24, 0) {real, imag} */,
  {32'hc041209f, 32'hc09ff4f2} /* (9, 23, 31) {real, imag} */,
  {32'h3f8096cb, 32'hbeee0c02} /* (9, 23, 30) {real, imag} */,
  {32'hbe89b1f7, 32'hbf74f951} /* (9, 23, 29) {real, imag} */,
  {32'h3f987b94, 32'h3f8a100d} /* (9, 23, 28) {real, imag} */,
  {32'hbf9f90e4, 32'hbcdecbab} /* (9, 23, 27) {real, imag} */,
  {32'h3f8874ee, 32'h4021311a} /* (9, 23, 26) {real, imag} */,
  {32'hbffbe287, 32'h3fb7d9cc} /* (9, 23, 25) {real, imag} */,
  {32'hbf42aa57, 32'hbf2d7bd5} /* (9, 23, 24) {real, imag} */,
  {32'hbfb905eb, 32'h3de0cb43} /* (9, 23, 23) {real, imag} */,
  {32'hbf8d7c44, 32'hbf93dc16} /* (9, 23, 22) {real, imag} */,
  {32'hc0149c67, 32'h3f61386c} /* (9, 23, 21) {real, imag} */,
  {32'h3fc52a9f, 32'hbfe047e4} /* (9, 23, 20) {real, imag} */,
  {32'hc00fc5a7, 32'h3f95cb6f} /* (9, 23, 19) {real, imag} */,
  {32'hbfb2f7ec, 32'h3ef99571} /* (9, 23, 18) {real, imag} */,
  {32'h4004fea7, 32'hbeba27b7} /* (9, 23, 17) {real, imag} */,
  {32'h3ee325a7, 32'h3eb4b580} /* (9, 23, 16) {real, imag} */,
  {32'hbf5e7444, 32'hbf1a9683} /* (9, 23, 15) {real, imag} */,
  {32'hbfb921ce, 32'h3ef22b73} /* (9, 23, 14) {real, imag} */,
  {32'h40135703, 32'hbf99433a} /* (9, 23, 13) {real, imag} */,
  {32'hbffc20e7, 32'h3e80ae7c} /* (9, 23, 12) {real, imag} */,
  {32'hbfbb8e34, 32'h3f8b1ffb} /* (9, 23, 11) {real, imag} */,
  {32'hbfeb0828, 32'h3ff9a610} /* (9, 23, 10) {real, imag} */,
  {32'hc0145a95, 32'h3ee591cc} /* (9, 23, 9) {real, imag} */,
  {32'h40c6b775, 32'hbf490c65} /* (9, 23, 8) {real, imag} */,
  {32'h3e1b6633, 32'hbf736339} /* (9, 23, 7) {real, imag} */,
  {32'h40058b56, 32'h3f3bcbb7} /* (9, 23, 6) {real, imag} */,
  {32'h3ff9a90c, 32'h3fa7a63a} /* (9, 23, 5) {real, imag} */,
  {32'hbfb22c5c, 32'h4089fff7} /* (9, 23, 4) {real, imag} */,
  {32'h3eab0d76, 32'hbf73ccd0} /* (9, 23, 3) {real, imag} */,
  {32'hbf42dd17, 32'hbf00dd19} /* (9, 23, 2) {real, imag} */,
  {32'h3f4cea85, 32'h40262cfa} /* (9, 23, 1) {real, imag} */,
  {32'h3f1eb59a, 32'h3ef9f15d} /* (9, 23, 0) {real, imag} */,
  {32'hbfdeccc6, 32'h4038f664} /* (9, 22, 31) {real, imag} */,
  {32'hbe8de840, 32'hc08188e9} /* (9, 22, 30) {real, imag} */,
  {32'hbfa03846, 32'h3f3dd51a} /* (9, 22, 29) {real, imag} */,
  {32'h3e8e1b11, 32'h402c7ebc} /* (9, 22, 28) {real, imag} */,
  {32'h3f0fed89, 32'h3fba361f} /* (9, 22, 27) {real, imag} */,
  {32'h401d3484, 32'hbe06a0d9} /* (9, 22, 26) {real, imag} */,
  {32'hc08a9ffe, 32'h3ffc41a8} /* (9, 22, 25) {real, imag} */,
  {32'hc0022602, 32'h3fc0e573} /* (9, 22, 24) {real, imag} */,
  {32'h3f3cd5f9, 32'hc00120f6} /* (9, 22, 23) {real, imag} */,
  {32'h3f68c817, 32'hbf5f94a3} /* (9, 22, 22) {real, imag} */,
  {32'hbf8e7b29, 32'hbe04e27b} /* (9, 22, 21) {real, imag} */,
  {32'h4078ad70, 32'hbffa8b84} /* (9, 22, 20) {real, imag} */,
  {32'hbe7adc2d, 32'hc01870e0} /* (9, 22, 19) {real, imag} */,
  {32'hbf798d14, 32'h3ec39c5c} /* (9, 22, 18) {real, imag} */,
  {32'h3ca755d4, 32'hbc2800b5} /* (9, 22, 17) {real, imag} */,
  {32'h3c477ec5, 32'h4004ce44} /* (9, 22, 16) {real, imag} */,
  {32'hbf0d57ab, 32'h3f07832b} /* (9, 22, 15) {real, imag} */,
  {32'h3db96266, 32'hbf9485e6} /* (9, 22, 14) {real, imag} */,
  {32'hbf8f1d62, 32'hc085cb11} /* (9, 22, 13) {real, imag} */,
  {32'h3fe71f2f, 32'hbfa9801f} /* (9, 22, 12) {real, imag} */,
  {32'h40295632, 32'h3fec0842} /* (9, 22, 11) {real, imag} */,
  {32'h3eff2056, 32'hc00bdfe1} /* (9, 22, 10) {real, imag} */,
  {32'h3f181b4b, 32'h4025618a} /* (9, 22, 9) {real, imag} */,
  {32'hbf7ea01c, 32'hbec1c92f} /* (9, 22, 8) {real, imag} */,
  {32'h3f917b22, 32'hbea27a04} /* (9, 22, 7) {real, imag} */,
  {32'h3f513ac4, 32'h4051335a} /* (9, 22, 6) {real, imag} */,
  {32'h3e2db7ad, 32'h3fa151f6} /* (9, 22, 5) {real, imag} */,
  {32'h3f021bcb, 32'hc0886396} /* (9, 22, 4) {real, imag} */,
  {32'h3ffb056d, 32'hbd508c0e} /* (9, 22, 3) {real, imag} */,
  {32'h3e864133, 32'h3e8eacca} /* (9, 22, 2) {real, imag} */,
  {32'h3fd115e8, 32'hbfca4872} /* (9, 22, 1) {real, imag} */,
  {32'h3f3049e5, 32'h3e1f653b} /* (9, 22, 0) {real, imag} */,
  {32'hbfb7d2c6, 32'h3f61331a} /* (9, 21, 31) {real, imag} */,
  {32'h3f982105, 32'hc0139c1b} /* (9, 21, 30) {real, imag} */,
  {32'hbf288060, 32'h40156c57} /* (9, 21, 29) {real, imag} */,
  {32'hbf47b9d8, 32'hc03567a6} /* (9, 21, 28) {real, imag} */,
  {32'hbf47814f, 32'h4003c81d} /* (9, 21, 27) {real, imag} */,
  {32'h4085a8d5, 32'hc01e89a9} /* (9, 21, 26) {real, imag} */,
  {32'h404167fa, 32'h3f9fd417} /* (9, 21, 25) {real, imag} */,
  {32'h3c9b4b9a, 32'h3f8e54c1} /* (9, 21, 24) {real, imag} */,
  {32'hbf06c4af, 32'hbedfd13b} /* (9, 21, 23) {real, imag} */,
  {32'hbd507cf4, 32'h3fce7ebb} /* (9, 21, 22) {real, imag} */,
  {32'hbf8aa64e, 32'h3f3ccea3} /* (9, 21, 21) {real, imag} */,
  {32'hbfcc4ba3, 32'h3f0f1d18} /* (9, 21, 20) {real, imag} */,
  {32'hbf75b414, 32'h4039e9a6} /* (9, 21, 19) {real, imag} */,
  {32'h4060fdfe, 32'hbf7af6bf} /* (9, 21, 18) {real, imag} */,
  {32'h3f4de953, 32'h3fa953b5} /* (9, 21, 17) {real, imag} */,
  {32'h3cf91bcf, 32'hbeea490b} /* (9, 21, 16) {real, imag} */,
  {32'h3cb48e7b, 32'hbf4a7ee3} /* (9, 21, 15) {real, imag} */,
  {32'hbf6f4f54, 32'hbe50d0e5} /* (9, 21, 14) {real, imag} */,
  {32'hbf1a87e2, 32'h3e217027} /* (9, 21, 13) {real, imag} */,
  {32'h3fe65ba9, 32'h3f6d6edc} /* (9, 21, 12) {real, imag} */,
  {32'h40123b9e, 32'h3fd244bf} /* (9, 21, 11) {real, imag} */,
  {32'hbf86dd36, 32'h3ffc5d92} /* (9, 21, 10) {real, imag} */,
  {32'hc0929feb, 32'h3e85deec} /* (9, 21, 9) {real, imag} */,
  {32'h3eeb6b80, 32'h3fc6f8a8} /* (9, 21, 8) {real, imag} */,
  {32'h3f1fb6e4, 32'hbf7b9aa6} /* (9, 21, 7) {real, imag} */,
  {32'h3f054095, 32'hc057c841} /* (9, 21, 6) {real, imag} */,
  {32'h405d7357, 32'h3eef0dd5} /* (9, 21, 5) {real, imag} */,
  {32'hc02c7a66, 32'hc001918a} /* (9, 21, 4) {real, imag} */,
  {32'hbdb7f06d, 32'hbf0dc19f} /* (9, 21, 3) {real, imag} */,
  {32'h3f922314, 32'h3fcc5df7} /* (9, 21, 2) {real, imag} */,
  {32'h3f056e42, 32'hbebc14bd} /* (9, 21, 1) {real, imag} */,
  {32'h3f8249bb, 32'h3faf3e72} /* (9, 21, 0) {real, imag} */,
  {32'h3f21df2b, 32'h3eb6a106} /* (9, 20, 31) {real, imag} */,
  {32'h3fba32ae, 32'h3f46b4c0} /* (9, 20, 30) {real, imag} */,
  {32'h3fb802c1, 32'hbf5f5761} /* (9, 20, 29) {real, imag} */,
  {32'h3f9727c1, 32'h3f7f8688} /* (9, 20, 28) {real, imag} */,
  {32'hc0081d20, 32'hbe909158} /* (9, 20, 27) {real, imag} */,
  {32'h3ebb17a8, 32'hbed15870} /* (9, 20, 26) {real, imag} */,
  {32'h3f276018, 32'h40802e2a} /* (9, 20, 25) {real, imag} */,
  {32'hbfef1bee, 32'hbe46e92e} /* (9, 20, 24) {real, imag} */,
  {32'hc0862b8b, 32'h3ed3e5ae} /* (9, 20, 23) {real, imag} */,
  {32'hbf3b770d, 32'h3f3f78f0} /* (9, 20, 22) {real, imag} */,
  {32'hbff39a91, 32'hbc98e734} /* (9, 20, 21) {real, imag} */,
  {32'h3fe533ea, 32'hc0a84dfd} /* (9, 20, 20) {real, imag} */,
  {32'h3f6047ea, 32'h40474382} /* (9, 20, 19) {real, imag} */,
  {32'h3f8bcc7d, 32'hbffc23e2} /* (9, 20, 18) {real, imag} */,
  {32'h3f134d5c, 32'h3f43d92b} /* (9, 20, 17) {real, imag} */,
  {32'hbed6c996, 32'h3f9e0d4d} /* (9, 20, 16) {real, imag} */,
  {32'hbf486a46, 32'h3f3efdff} /* (9, 20, 15) {real, imag} */,
  {32'hbf345e53, 32'h40154866} /* (9, 20, 14) {real, imag} */,
  {32'h3fe50a2b, 32'h3ea716ba} /* (9, 20, 13) {real, imag} */,
  {32'hbf1f698b, 32'h3fb6c1b5} /* (9, 20, 12) {real, imag} */,
  {32'hc02e219a, 32'h4043f163} /* (9, 20, 11) {real, imag} */,
  {32'h3ff6e304, 32'hbfba437b} /* (9, 20, 10) {real, imag} */,
  {32'hc005c47b, 32'hbfbfb2e8} /* (9, 20, 9) {real, imag} */,
  {32'h3ffd944f, 32'hbfa33b5c} /* (9, 20, 8) {real, imag} */,
  {32'hbfd736b5, 32'hbf2f0edd} /* (9, 20, 7) {real, imag} */,
  {32'h3fad766c, 32'hc02c1507} /* (9, 20, 6) {real, imag} */,
  {32'h3ec15963, 32'h3d831297} /* (9, 20, 5) {real, imag} */,
  {32'h3f70f6f9, 32'h3f9e492c} /* (9, 20, 4) {real, imag} */,
  {32'hc00d3275, 32'hc014762b} /* (9, 20, 3) {real, imag} */,
  {32'hbfcf89f2, 32'hbf62c604} /* (9, 20, 2) {real, imag} */,
  {32'h3eb53e03, 32'hbfdb28fc} /* (9, 20, 1) {real, imag} */,
  {32'h3fb3e015, 32'h3e73b4d7} /* (9, 20, 0) {real, imag} */,
  {32'hbc5d6502, 32'hbf104937} /* (9, 19, 31) {real, imag} */,
  {32'hbf60613b, 32'h3e8714a0} /* (9, 19, 30) {real, imag} */,
  {32'h3f634d83, 32'hbf871686} /* (9, 19, 29) {real, imag} */,
  {32'hc001f283, 32'h3ed7e745} /* (9, 19, 28) {real, imag} */,
  {32'h3f770f94, 32'h40179f45} /* (9, 19, 27) {real, imag} */,
  {32'hbd8a024c, 32'h3f35734a} /* (9, 19, 26) {real, imag} */,
  {32'h3fc0f1fd, 32'h3f3ae3da} /* (9, 19, 25) {real, imag} */,
  {32'h4049783f, 32'h3fc8bc3c} /* (9, 19, 24) {real, imag} */,
  {32'hbf150990, 32'hbf8eba21} /* (9, 19, 23) {real, imag} */,
  {32'hc0085bfa, 32'h3eccc82d} /* (9, 19, 22) {real, imag} */,
  {32'hc0226f8d, 32'h3ec361e5} /* (9, 19, 21) {real, imag} */,
  {32'h3fd1425c, 32'hc0486079} /* (9, 19, 20) {real, imag} */,
  {32'h3f9da7a6, 32'hc0053a7f} /* (9, 19, 19) {real, imag} */,
  {32'h3ff1c125, 32'hbf8a7348} /* (9, 19, 18) {real, imag} */,
  {32'hc001794c, 32'hbfe2599e} /* (9, 19, 17) {real, imag} */,
  {32'h3e069dbe, 32'hbe8dd6f8} /* (9, 19, 16) {real, imag} */,
  {32'h3f9cd22c, 32'h40541a71} /* (9, 19, 15) {real, imag} */,
  {32'h3f7350ee, 32'h3fdc2476} /* (9, 19, 14) {real, imag} */,
  {32'h401201de, 32'h3e01d939} /* (9, 19, 13) {real, imag} */,
  {32'hbf37adef, 32'h3f2c45e3} /* (9, 19, 12) {real, imag} */,
  {32'hbf4dc1ee, 32'hc04839fd} /* (9, 19, 11) {real, imag} */,
  {32'hc06a8826, 32'h3e95dff8} /* (9, 19, 10) {real, imag} */,
  {32'h3f5d6560, 32'hbf10ce59} /* (9, 19, 9) {real, imag} */,
  {32'hbe495688, 32'hbf342a06} /* (9, 19, 8) {real, imag} */,
  {32'hbebd1eb5, 32'h3dffdf45} /* (9, 19, 7) {real, imag} */,
  {32'hbffc42e8, 32'hbe8a6e4d} /* (9, 19, 6) {real, imag} */,
  {32'hbef31227, 32'h3fc6c667} /* (9, 19, 5) {real, imag} */,
  {32'hbfa2ea40, 32'hc062c51a} /* (9, 19, 4) {real, imag} */,
  {32'h3f770754, 32'h3ff55952} /* (9, 19, 3) {real, imag} */,
  {32'hbe847887, 32'hbf658aa3} /* (9, 19, 2) {real, imag} */,
  {32'h3f1135f0, 32'hbff3f4ca} /* (9, 19, 1) {real, imag} */,
  {32'hc01293d0, 32'hc08bfbc8} /* (9, 19, 0) {real, imag} */,
  {32'h3ef629c7, 32'h3fcced10} /* (9, 18, 31) {real, imag} */,
  {32'h3f8b08eb, 32'hc00f0ab3} /* (9, 18, 30) {real, imag} */,
  {32'hbe81080f, 32'h3f6613e6} /* (9, 18, 29) {real, imag} */,
  {32'hbf7853aa, 32'hbfad3737} /* (9, 18, 28) {real, imag} */,
  {32'hbff0cf1b, 32'hbe4709bd} /* (9, 18, 27) {real, imag} */,
  {32'h3eff622e, 32'hbf8b55ed} /* (9, 18, 26) {real, imag} */,
  {32'h3f3d0be8, 32'h3f50db64} /* (9, 18, 25) {real, imag} */,
  {32'hbe29b724, 32'h3ee9d7ce} /* (9, 18, 24) {real, imag} */,
  {32'h3ee6e345, 32'hbe18691d} /* (9, 18, 23) {real, imag} */,
  {32'h402e474a, 32'h3f4517de} /* (9, 18, 22) {real, imag} */,
  {32'h3cfcac86, 32'hc018e331} /* (9, 18, 21) {real, imag} */,
  {32'h401c4953, 32'h4091bef0} /* (9, 18, 20) {real, imag} */,
  {32'hbf3ac754, 32'hbf6ae710} /* (9, 18, 19) {real, imag} */,
  {32'h3fa39bd7, 32'hbe85394b} /* (9, 18, 18) {real, imag} */,
  {32'hbfd805fa, 32'h3f7535be} /* (9, 18, 17) {real, imag} */,
  {32'hbf112645, 32'hbf5982c2} /* (9, 18, 16) {real, imag} */,
  {32'h3f52fbda, 32'hbfb913d5} /* (9, 18, 15) {real, imag} */,
  {32'h3f7c2137, 32'h3f8a409f} /* (9, 18, 14) {real, imag} */,
  {32'h3f94a5bb, 32'hbfd103f5} /* (9, 18, 13) {real, imag} */,
  {32'h3fdc6f6c, 32'h3e74bb0d} /* (9, 18, 12) {real, imag} */,
  {32'hbdf01ea6, 32'hbfe0ec05} /* (9, 18, 11) {real, imag} */,
  {32'h3fdaaeca, 32'hbfa3ab88} /* (9, 18, 10) {real, imag} */,
  {32'hbf20ab09, 32'hbfe0f14c} /* (9, 18, 9) {real, imag} */,
  {32'hc037dded, 32'hc0107b4e} /* (9, 18, 8) {real, imag} */,
  {32'hc00d55ee, 32'h3df1184d} /* (9, 18, 7) {real, imag} */,
  {32'h3fc2e92a, 32'h3f241456} /* (9, 18, 6) {real, imag} */,
  {32'h3fa0e388, 32'h4042c7fa} /* (9, 18, 5) {real, imag} */,
  {32'hbf9817fe, 32'h3f99e51b} /* (9, 18, 4) {real, imag} */,
  {32'h3fbc3c51, 32'h3fa3a288} /* (9, 18, 3) {real, imag} */,
  {32'hbf8b290b, 32'hbfd752bd} /* (9, 18, 2) {real, imag} */,
  {32'hbf01e355, 32'h3f5aaeb5} /* (9, 18, 1) {real, imag} */,
  {32'h3e965097, 32'hbf293d1e} /* (9, 18, 0) {real, imag} */,
  {32'hbf82982b, 32'h3f94f5c4} /* (9, 17, 31) {real, imag} */,
  {32'h3e4bcf0f, 32'hc0052852} /* (9, 17, 30) {real, imag} */,
  {32'h3f9d04c0, 32'h3f2e8a4b} /* (9, 17, 29) {real, imag} */,
  {32'hbfd8d04c, 32'hbe0d5d9a} /* (9, 17, 28) {real, imag} */,
  {32'h3eeeb2e6, 32'h40199b7d} /* (9, 17, 27) {real, imag} */,
  {32'hbfef754c, 32'hbfef14f8} /* (9, 17, 26) {real, imag} */,
  {32'h3dcefd24, 32'h3f81fb34} /* (9, 17, 25) {real, imag} */,
  {32'h408fb545, 32'h3fee17ad} /* (9, 17, 24) {real, imag} */,
  {32'h40192aa4, 32'h3f812629} /* (9, 17, 23) {real, imag} */,
  {32'h3f2b557c, 32'h3ee73a98} /* (9, 17, 22) {real, imag} */,
  {32'hbf875c67, 32'h3da1e611} /* (9, 17, 21) {real, imag} */,
  {32'h3f831d43, 32'h3f8d19e9} /* (9, 17, 20) {real, imag} */,
  {32'h3fa77384, 32'h3f71f340} /* (9, 17, 19) {real, imag} */,
  {32'h3e936cb1, 32'h3f81db40} /* (9, 17, 18) {real, imag} */,
  {32'hbfa152d3, 32'hbff477ba} /* (9, 17, 17) {real, imag} */,
  {32'hbfefcebf, 32'h3dc4afe3} /* (9, 17, 16) {real, imag} */,
  {32'hbf67ea5f, 32'h3f0bb671} /* (9, 17, 15) {real, imag} */,
  {32'hbec6ee28, 32'hbf3379fb} /* (9, 17, 14) {real, imag} */,
  {32'hbe458612, 32'hbff312ae} /* (9, 17, 13) {real, imag} */,
  {32'h3f66f9a3, 32'h400ad2e1} /* (9, 17, 12) {real, imag} */,
  {32'hbfa241dd, 32'hc06ba6ea} /* (9, 17, 11) {real, imag} */,
  {32'h3ee53a32, 32'h3fdc70e7} /* (9, 17, 10) {real, imag} */,
  {32'h402d5388, 32'h3f014b09} /* (9, 17, 9) {real, imag} */,
  {32'hbe853cba, 32'h3f8e1c7a} /* (9, 17, 8) {real, imag} */,
  {32'hbf106048, 32'h3f844713} /* (9, 17, 7) {real, imag} */,
  {32'hbf90f2d4, 32'hc01dd175} /* (9, 17, 6) {real, imag} */,
  {32'hbed00341, 32'hbe08ccb8} /* (9, 17, 5) {real, imag} */,
  {32'h3fc2bc36, 32'hbf9c5e63} /* (9, 17, 4) {real, imag} */,
  {32'hbe83da49, 32'h3f677a2a} /* (9, 17, 3) {real, imag} */,
  {32'hbb7b9626, 32'hbfe9c1c9} /* (9, 17, 2) {real, imag} */,
  {32'h3f933411, 32'hbf35f179} /* (9, 17, 1) {real, imag} */,
  {32'h3ff80c0c, 32'hbe38f19e} /* (9, 17, 0) {real, imag} */,
  {32'hbefd2ba3, 32'h3f2bd271} /* (9, 16, 31) {real, imag} */,
  {32'h3f4fb198, 32'hbe82b21e} /* (9, 16, 30) {real, imag} */,
  {32'h3f131eca, 32'hbf533f3e} /* (9, 16, 29) {real, imag} */,
  {32'h3e936e1d, 32'h3f96bc94} /* (9, 16, 28) {real, imag} */,
  {32'h3e897f5d, 32'h3ecf734f} /* (9, 16, 27) {real, imag} */,
  {32'h3f87abd4, 32'h3f83d20a} /* (9, 16, 26) {real, imag} */,
  {32'hbe83bd65, 32'hbf3843c9} /* (9, 16, 25) {real, imag} */,
  {32'hbf48aa8c, 32'hbf3bc06f} /* (9, 16, 24) {real, imag} */,
  {32'h3f897879, 32'h3f8360ee} /* (9, 16, 23) {real, imag} */,
  {32'h3ed390b1, 32'h3fc008ed} /* (9, 16, 22) {real, imag} */,
  {32'hbe39e4f3, 32'hbfbdf706} /* (9, 16, 21) {real, imag} */,
  {32'hbfc307e4, 32'h40663ee8} /* (9, 16, 20) {real, imag} */,
  {32'h3f9f6a95, 32'hbe2a7b91} /* (9, 16, 19) {real, imag} */,
  {32'h3ee035d6, 32'hbe4e0af1} /* (9, 16, 18) {real, imag} */,
  {32'hbfc15ce8, 32'hbffa315a} /* (9, 16, 17) {real, imag} */,
  {32'hbf4a02a2, 32'hc00f3871} /* (9, 16, 16) {real, imag} */,
  {32'h3fbb722c, 32'hbf288735} /* (9, 16, 15) {real, imag} */,
  {32'hbff91166, 32'hbeb0384f} /* (9, 16, 14) {real, imag} */,
  {32'hc023e0af, 32'hbf91a5a2} /* (9, 16, 13) {real, imag} */,
  {32'hbf91d25c, 32'hbfd003be} /* (9, 16, 12) {real, imag} */,
  {32'h3f049f35, 32'h400f124e} /* (9, 16, 11) {real, imag} */,
  {32'h3ebe0ca1, 32'h3f26beae} /* (9, 16, 10) {real, imag} */,
  {32'h3d17ecfb, 32'hbf650485} /* (9, 16, 9) {real, imag} */,
  {32'h3f333cf4, 32'h3fe189e1} /* (9, 16, 8) {real, imag} */,
  {32'h3f61a49f, 32'h3fbadf7b} /* (9, 16, 7) {real, imag} */,
  {32'h3e1347be, 32'h3fe69eca} /* (9, 16, 6) {real, imag} */,
  {32'h3ff6c504, 32'hbfa62a73} /* (9, 16, 5) {real, imag} */,
  {32'h3f20ecd3, 32'hbfed8738} /* (9, 16, 4) {real, imag} */,
  {32'hbf145187, 32'h3f12e541} /* (9, 16, 3) {real, imag} */,
  {32'hbf0747ed, 32'hbe050f39} /* (9, 16, 2) {real, imag} */,
  {32'h3f9baa43, 32'h3fae4b03} /* (9, 16, 1) {real, imag} */,
  {32'h3f2c2349, 32'hc0003d48} /* (9, 16, 0) {real, imag} */,
  {32'hbea9dc68, 32'hbce411b3} /* (9, 15, 31) {real, imag} */,
  {32'h3e8353dc, 32'h3f8b1737} /* (9, 15, 30) {real, imag} */,
  {32'h3fe81a1d, 32'h3ff2e3a1} /* (9, 15, 29) {real, imag} */,
  {32'hbf85d4e2, 32'hbf633958} /* (9, 15, 28) {real, imag} */,
  {32'h3f1cd9c8, 32'h400f7abc} /* (9, 15, 27) {real, imag} */,
  {32'h3f0e0cf8, 32'h3e77aa3e} /* (9, 15, 26) {real, imag} */,
  {32'hbfd99d06, 32'hbf86d7d7} /* (9, 15, 25) {real, imag} */,
  {32'hbf5f69fa, 32'hbf380d28} /* (9, 15, 24) {real, imag} */,
  {32'hbf6a77d2, 32'hbeef68d5} /* (9, 15, 23) {real, imag} */,
  {32'hc0127789, 32'hbf899f10} /* (9, 15, 22) {real, imag} */,
  {32'hbe727dd1, 32'h3f9afdb2} /* (9, 15, 21) {real, imag} */,
  {32'hbee06e9d, 32'hbfe197c5} /* (9, 15, 20) {real, imag} */,
  {32'h3fb841ed, 32'h40081b81} /* (9, 15, 19) {real, imag} */,
  {32'h3e720c25, 32'h3ed06f19} /* (9, 15, 18) {real, imag} */,
  {32'h3f448e39, 32'hbefc8c3e} /* (9, 15, 17) {real, imag} */,
  {32'hbf34e185, 32'hbf58dbee} /* (9, 15, 16) {real, imag} */,
  {32'h4037670e, 32'h3f9a7dd8} /* (9, 15, 15) {real, imag} */,
  {32'h3ff6e5fc, 32'hbfe29496} /* (9, 15, 14) {real, imag} */,
  {32'h403347ec, 32'hbef96fa0} /* (9, 15, 13) {real, imag} */,
  {32'hbf99db31, 32'hbfc0fc84} /* (9, 15, 12) {real, imag} */,
  {32'hbffdbccf, 32'h3f812175} /* (9, 15, 11) {real, imag} */,
  {32'h3fd34d31, 32'h4016a1d8} /* (9, 15, 10) {real, imag} */,
  {32'hbeef2bc2, 32'hbf1d48c7} /* (9, 15, 9) {real, imag} */,
  {32'h402337ff, 32'hbedf8d05} /* (9, 15, 8) {real, imag} */,
  {32'h3f26afb9, 32'hbf823536} /* (9, 15, 7) {real, imag} */,
  {32'hc0060ed0, 32'h3f350f69} /* (9, 15, 6) {real, imag} */,
  {32'hbf7fb184, 32'hbede322b} /* (9, 15, 5) {real, imag} */,
  {32'hbfe4bef2, 32'hbdd12ada} /* (9, 15, 4) {real, imag} */,
  {32'h3e8dd83a, 32'hbf12e251} /* (9, 15, 3) {real, imag} */,
  {32'hbd89ec92, 32'h3f8f5892} /* (9, 15, 2) {real, imag} */,
  {32'hbfe283d9, 32'h3fc875c0} /* (9, 15, 1) {real, imag} */,
  {32'h3f4fd711, 32'hbf0eb377} /* (9, 15, 0) {real, imag} */,
  {32'h3f741555, 32'h3f0be4ff} /* (9, 14, 31) {real, imag} */,
  {32'hc011a5e8, 32'hbf245269} /* (9, 14, 30) {real, imag} */,
  {32'hc012a127, 32'h3eadb345} /* (9, 14, 29) {real, imag} */,
  {32'h3fb6bef6, 32'h4064f356} /* (9, 14, 28) {real, imag} */,
  {32'hbd1603d0, 32'hc013fe01} /* (9, 14, 27) {real, imag} */,
  {32'hbfa3646a, 32'hbee8d012} /* (9, 14, 26) {real, imag} */,
  {32'hc01c6af1, 32'hbfa4cff8} /* (9, 14, 25) {real, imag} */,
  {32'hbf650c94, 32'hbde37e46} /* (9, 14, 24) {real, imag} */,
  {32'h3d99cb12, 32'hbfe8f128} /* (9, 14, 23) {real, imag} */,
  {32'h3e8ebf59, 32'hbfe287ad} /* (9, 14, 22) {real, imag} */,
  {32'hbfa6d6da, 32'hbfce79da} /* (9, 14, 21) {real, imag} */,
  {32'hbf64e02a, 32'h3fbfef1e} /* (9, 14, 20) {real, imag} */,
  {32'hbfce3d25, 32'hc00a1228} /* (9, 14, 19) {real, imag} */,
  {32'hbc007ed6, 32'h3ec4ae78} /* (9, 14, 18) {real, imag} */,
  {32'h3ef34559, 32'hbfe6f128} /* (9, 14, 17) {real, imag} */,
  {32'hbf1f3fcf, 32'h3f06afcf} /* (9, 14, 16) {real, imag} */,
  {32'hbf136f93, 32'hbd97011a} /* (9, 14, 15) {real, imag} */,
  {32'hbf2b9b10, 32'hbf578d83} /* (9, 14, 14) {real, imag} */,
  {32'h3c93484b, 32'h3ee580ee} /* (9, 14, 13) {real, imag} */,
  {32'hbf518f8e, 32'hbd92d2bb} /* (9, 14, 12) {real, imag} */,
  {32'h3f972402, 32'h3fb86e1a} /* (9, 14, 11) {real, imag} */,
  {32'hbf03f4e7, 32'h403a84e0} /* (9, 14, 10) {real, imag} */,
  {32'hbfc97631, 32'h3f9a1d9a} /* (9, 14, 9) {real, imag} */,
  {32'h3fd76763, 32'hbff32086} /* (9, 14, 8) {real, imag} */,
  {32'hc094ad49, 32'hbf9d8b69} /* (9, 14, 7) {real, imag} */,
  {32'h3dda5bb8, 32'h3e38beae} /* (9, 14, 6) {real, imag} */,
  {32'h3f942711, 32'h3e9e4618} /* (9, 14, 5) {real, imag} */,
  {32'h4034a3e6, 32'h405475cc} /* (9, 14, 4) {real, imag} */,
  {32'h3f15e2fb, 32'h3fe0098b} /* (9, 14, 3) {real, imag} */,
  {32'hbfbc4d46, 32'h3dcb897b} /* (9, 14, 2) {real, imag} */,
  {32'hbf82d915, 32'h3feec0ae} /* (9, 14, 1) {real, imag} */,
  {32'hbeea9cf2, 32'h4004fed9} /* (9, 14, 0) {real, imag} */,
  {32'hbede8263, 32'hbfc6f924} /* (9, 13, 31) {real, imag} */,
  {32'h400e6d33, 32'hbea534e0} /* (9, 13, 30) {real, imag} */,
  {32'h3e165320, 32'h3fc80033} /* (9, 13, 29) {real, imag} */,
  {32'h3f177e7a, 32'hc04d31bb} /* (9, 13, 28) {real, imag} */,
  {32'h3ef800ec, 32'hbf4a9435} /* (9, 13, 27) {real, imag} */,
  {32'hbfd6ac68, 32'hbf72be00} /* (9, 13, 26) {real, imag} */,
  {32'h3efe313e, 32'h3f295541} /* (9, 13, 25) {real, imag} */,
  {32'h3f8a1812, 32'hc042a340} /* (9, 13, 24) {real, imag} */,
  {32'h3ef3d317, 32'hbf960a41} /* (9, 13, 23) {real, imag} */,
  {32'h3fa3129c, 32'hbfc945ac} /* (9, 13, 22) {real, imag} */,
  {32'h3e8c453d, 32'h3f29fe08} /* (9, 13, 21) {real, imag} */,
  {32'hbe543ce2, 32'hc0296ab6} /* (9, 13, 20) {real, imag} */,
  {32'h3f1e4111, 32'h40609a50} /* (9, 13, 19) {real, imag} */,
  {32'h3ed59c9b, 32'hbe175254} /* (9, 13, 18) {real, imag} */,
  {32'h3faaa389, 32'h3fb35754} /* (9, 13, 17) {real, imag} */,
  {32'hbe3d89c6, 32'h3de0ea18} /* (9, 13, 16) {real, imag} */,
  {32'hbf780e0f, 32'hbef8c572} /* (9, 13, 15) {real, imag} */,
  {32'h3e1beadf, 32'h3f254493} /* (9, 13, 14) {real, imag} */,
  {32'h3f9365a1, 32'h3ff651fd} /* (9, 13, 13) {real, imag} */,
  {32'hbec284bc, 32'h404f7c50} /* (9, 13, 12) {real, imag} */,
  {32'h407b2778, 32'hbfe09245} /* (9, 13, 11) {real, imag} */,
  {32'hc0257d2d, 32'h3fd948df} /* (9, 13, 10) {real, imag} */,
  {32'hc033a6be, 32'h4003ad44} /* (9, 13, 9) {real, imag} */,
  {32'hbfda96f6, 32'hbf84e225} /* (9, 13, 8) {real, imag} */,
  {32'hbd0e830a, 32'hbd149e4e} /* (9, 13, 7) {real, imag} */,
  {32'h3d742bc8, 32'h3f93f0b4} /* (9, 13, 6) {real, imag} */,
  {32'hc05657e9, 32'h3fbe896f} /* (9, 13, 5) {real, imag} */,
  {32'h40587ba0, 32'h3f59d3fc} /* (9, 13, 4) {real, imag} */,
  {32'hbf31c132, 32'hc0240681} /* (9, 13, 3) {real, imag} */,
  {32'hbf5b566c, 32'hbfcfa0ce} /* (9, 13, 2) {real, imag} */,
  {32'hc023ccc4, 32'hbf4a415c} /* (9, 13, 1) {real, imag} */,
  {32'hbe37d244, 32'hbefd3603} /* (9, 13, 0) {real, imag} */,
  {32'h3fecb699, 32'h40280949} /* (9, 12, 31) {real, imag} */,
  {32'hbf2e980a, 32'h3ed33c99} /* (9, 12, 30) {real, imag} */,
  {32'hc01edcfa, 32'h3eb3473e} /* (9, 12, 29) {real, imag} */,
  {32'hbe6e5ac1, 32'h3fe48789} /* (9, 12, 28) {real, imag} */,
  {32'hbf604ae0, 32'hc0102067} /* (9, 12, 27) {real, imag} */,
  {32'hc04741f7, 32'h4030b850} /* (9, 12, 26) {real, imag} */,
  {32'hbf2d23b1, 32'hbffd2219} /* (9, 12, 25) {real, imag} */,
  {32'h3fd551d4, 32'h3fb19888} /* (9, 12, 24) {real, imag} */,
  {32'hbf9d983e, 32'h4050a318} /* (9, 12, 23) {real, imag} */,
  {32'hbfc13925, 32'hbfaa2699} /* (9, 12, 22) {real, imag} */,
  {32'h3fe6190d, 32'h408970c6} /* (9, 12, 21) {real, imag} */,
  {32'h3eb82e41, 32'h3dbab44f} /* (9, 12, 20) {real, imag} */,
  {32'h400f5ef9, 32'hbf0047e6} /* (9, 12, 19) {real, imag} */,
  {32'h406b1ad3, 32'h3ef1a48a} /* (9, 12, 18) {real, imag} */,
  {32'h4022c8f8, 32'h3f34fc0b} /* (9, 12, 17) {real, imag} */,
  {32'hc019fb8b, 32'hbf5aaa89} /* (9, 12, 16) {real, imag} */,
  {32'hbeabe509, 32'hbf6b7d0d} /* (9, 12, 15) {real, imag} */,
  {32'h3f0a0db5, 32'hbf7bd7ab} /* (9, 12, 14) {real, imag} */,
  {32'h3ff4eceb, 32'h3fe84b38} /* (9, 12, 13) {real, imag} */,
  {32'h3fa5325f, 32'hbe1b4b1f} /* (9, 12, 12) {real, imag} */,
  {32'h3fe2fa5f, 32'hbf66522c} /* (9, 12, 11) {real, imag} */,
  {32'hbf79577f, 32'h3ff68c1e} /* (9, 12, 10) {real, imag} */,
  {32'h3c27b10d, 32'hc0226588} /* (9, 12, 9) {real, imag} */,
  {32'hbd6b0d36, 32'h4009f749} /* (9, 12, 8) {real, imag} */,
  {32'h3fe38429, 32'h3ebbb3bf} /* (9, 12, 7) {real, imag} */,
  {32'h3f3f1d99, 32'h3f656beb} /* (9, 12, 6) {real, imag} */,
  {32'h3fa04d8f, 32'hbff1573b} /* (9, 12, 5) {real, imag} */,
  {32'h3f19756f, 32'h3eb8ad75} /* (9, 12, 4) {real, imag} */,
  {32'hbfbcf93e, 32'h3d2d99ee} /* (9, 12, 3) {real, imag} */,
  {32'h401145ff, 32'h3f024809} /* (9, 12, 2) {real, imag} */,
  {32'h4017e819, 32'hbfbc6fae} /* (9, 12, 1) {real, imag} */,
  {32'hbfc99c3d, 32'h3f0acaaf} /* (9, 12, 0) {real, imag} */,
  {32'hbf320b7f, 32'hbf4afcc1} /* (9, 11, 31) {real, imag} */,
  {32'hbe96f736, 32'hc00be92c} /* (9, 11, 30) {real, imag} */,
  {32'hc026f07a, 32'hbf66638d} /* (9, 11, 29) {real, imag} */,
  {32'hbfc40310, 32'hbeeb4664} /* (9, 11, 28) {real, imag} */,
  {32'hc082594b, 32'h3fa77802} /* (9, 11, 27) {real, imag} */,
  {32'h3fa9c588, 32'h40104b74} /* (9, 11, 26) {real, imag} */,
  {32'h40854ae2, 32'h401599a9} /* (9, 11, 25) {real, imag} */,
  {32'h405e1900, 32'hbe7874ee} /* (9, 11, 24) {real, imag} */,
  {32'hc08272bb, 32'hbef36b3c} /* (9, 11, 23) {real, imag} */,
  {32'hbda72796, 32'h3fee1654} /* (9, 11, 22) {real, imag} */,
  {32'hc03faa41, 32'hc042deae} /* (9, 11, 21) {real, imag} */,
  {32'h3f906ecc, 32'hc00a6f88} /* (9, 11, 20) {real, imag} */,
  {32'h3ffada80, 32'hbf87f42a} /* (9, 11, 19) {real, imag} */,
  {32'hbe72262c, 32'h3fefe00b} /* (9, 11, 18) {real, imag} */,
  {32'h3fa536c5, 32'hc02775c0} /* (9, 11, 17) {real, imag} */,
  {32'hbe9d34e6, 32'hbf8e0200} /* (9, 11, 16) {real, imag} */,
  {32'hbfe3a2be, 32'h3fbd23aa} /* (9, 11, 15) {real, imag} */,
  {32'h3fe73e75, 32'h3f293f4d} /* (9, 11, 14) {real, imag} */,
  {32'h3e6412cd, 32'h3fec2fdb} /* (9, 11, 13) {real, imag} */,
  {32'h3fbad6dc, 32'h3fa1eaf9} /* (9, 11, 12) {real, imag} */,
  {32'hc02ea8b1, 32'hbe5fc7da} /* (9, 11, 11) {real, imag} */,
  {32'h3fe16bfc, 32'h40812dca} /* (9, 11, 10) {real, imag} */,
  {32'h405c94b1, 32'hbe1478a1} /* (9, 11, 9) {real, imag} */,
  {32'h40063b05, 32'h3fd48214} /* (9, 11, 8) {real, imag} */,
  {32'h40175d68, 32'h3fdadbae} /* (9, 11, 7) {real, imag} */,
  {32'h3f7beeaa, 32'h401129d5} /* (9, 11, 6) {real, imag} */,
  {32'h40436bc9, 32'h40652a47} /* (9, 11, 5) {real, imag} */,
  {32'h3fce272b, 32'hbfa4a288} /* (9, 11, 4) {real, imag} */,
  {32'hbff20695, 32'h4080ddd9} /* (9, 11, 3) {real, imag} */,
  {32'hbe6d371b, 32'h3fc73765} /* (9, 11, 2) {real, imag} */,
  {32'h4020f36d, 32'h3f1e9735} /* (9, 11, 1) {real, imag} */,
  {32'hc029d401, 32'h3f886829} /* (9, 11, 0) {real, imag} */,
  {32'h3f79a495, 32'hbfa0fe17} /* (9, 10, 31) {real, imag} */,
  {32'hc0284e2c, 32'hbf2622fa} /* (9, 10, 30) {real, imag} */,
  {32'h3eceae8f, 32'hbf89dc8b} /* (9, 10, 29) {real, imag} */,
  {32'h3e38411e, 32'h3f13cea0} /* (9, 10, 28) {real, imag} */,
  {32'h40511454, 32'hbfcbe563} /* (9, 10, 27) {real, imag} */,
  {32'h3fa69518, 32'h401e8f20} /* (9, 10, 26) {real, imag} */,
  {32'h40098d08, 32'h3a9aecbf} /* (9, 10, 25) {real, imag} */,
  {32'hbf5cdaae, 32'h401619c8} /* (9, 10, 24) {real, imag} */,
  {32'h402b5225, 32'h4010a382} /* (9, 10, 23) {real, imag} */,
  {32'hbf629766, 32'h3fd02024} /* (9, 10, 22) {real, imag} */,
  {32'h4023837e, 32'h3eb47964} /* (9, 10, 21) {real, imag} */,
  {32'hbe81cfcb, 32'hc08ee777} /* (9, 10, 20) {real, imag} */,
  {32'hc08a4673, 32'hc0097116} /* (9, 10, 19) {real, imag} */,
  {32'h3f9d2c70, 32'hc03753e7} /* (9, 10, 18) {real, imag} */,
  {32'h3fc6e694, 32'hbf203fea} /* (9, 10, 17) {real, imag} */,
  {32'h3fc05df6, 32'h40211ae2} /* (9, 10, 16) {real, imag} */,
  {32'hc002f9bb, 32'hc0068384} /* (9, 10, 15) {real, imag} */,
  {32'hbea6b2ea, 32'hc03552e2} /* (9, 10, 14) {real, imag} */,
  {32'hbee0a02b, 32'hbfbbbd7c} /* (9, 10, 13) {real, imag} */,
  {32'h3fbc4052, 32'hbfbc6e45} /* (9, 10, 12) {real, imag} */,
  {32'h402ca666, 32'h3d85e7fb} /* (9, 10, 11) {real, imag} */,
  {32'hbee21476, 32'hbffd04ae} /* (9, 10, 10) {real, imag} */,
  {32'h3f6dbd98, 32'h3f82a51e} /* (9, 10, 9) {real, imag} */,
  {32'h3f4ae95b, 32'hbfacb308} /* (9, 10, 8) {real, imag} */,
  {32'hbff9ce8c, 32'hbf50f466} /* (9, 10, 7) {real, imag} */,
  {32'hbe6f66f4, 32'hbf5b8c4a} /* (9, 10, 6) {real, imag} */,
  {32'h3f3fc053, 32'h3faef594} /* (9, 10, 5) {real, imag} */,
  {32'h3cda1e06, 32'h3f90d47f} /* (9, 10, 4) {real, imag} */,
  {32'hc028c3a6, 32'h40372761} /* (9, 10, 3) {real, imag} */,
  {32'h409cbffb, 32'h3eab053d} /* (9, 10, 2) {real, imag} */,
  {32'hbeff9441, 32'hbcab2acb} /* (9, 10, 1) {real, imag} */,
  {32'hbfae5fff, 32'h3f7779ee} /* (9, 10, 0) {real, imag} */,
  {32'hc022111f, 32'h3fd6d9a6} /* (9, 9, 31) {real, imag} */,
  {32'h401988ff, 32'hbfebee37} /* (9, 9, 30) {real, imag} */,
  {32'h3f327902, 32'h3f06937a} /* (9, 9, 29) {real, imag} */,
  {32'h3fce36f8, 32'h3fbcb4e5} /* (9, 9, 28) {real, imag} */,
  {32'hbf5a2846, 32'hbeea76a3} /* (9, 9, 27) {real, imag} */,
  {32'hc03b030c, 32'hc01181c5} /* (9, 9, 26) {real, imag} */,
  {32'hc02f73ac, 32'h4005a414} /* (9, 9, 25) {real, imag} */,
  {32'h3ddfaf54, 32'h3e6f1be3} /* (9, 9, 24) {real, imag} */,
  {32'hbe0c3a69, 32'h3e5bdd8b} /* (9, 9, 23) {real, imag} */,
  {32'h3e0ce500, 32'hc088bf68} /* (9, 9, 22) {real, imag} */,
  {32'h400284d4, 32'hbf2c123c} /* (9, 9, 21) {real, imag} */,
  {32'h3fe827ef, 32'h3fdfdbd4} /* (9, 9, 20) {real, imag} */,
  {32'h402c9d8a, 32'hc0339f9d} /* (9, 9, 19) {real, imag} */,
  {32'h3bc98101, 32'h3e5a2630} /* (9, 9, 18) {real, imag} */,
  {32'hbf39f8f1, 32'hbfcefdfd} /* (9, 9, 17) {real, imag} */,
  {32'h3e0e76dc, 32'hbff7a879} /* (9, 9, 16) {real, imag} */,
  {32'hbef9ae05, 32'hbf1aded0} /* (9, 9, 15) {real, imag} */,
  {32'hbf8471f5, 32'h3fecf7d0} /* (9, 9, 14) {real, imag} */,
  {32'hbed9019c, 32'h3ea0ee6f} /* (9, 9, 13) {real, imag} */,
  {32'hc0229e00, 32'hc06ddd51} /* (9, 9, 12) {real, imag} */,
  {32'hc00dda31, 32'h3fda676c} /* (9, 9, 11) {real, imag} */,
  {32'h3ff8e9b5, 32'h406cee5d} /* (9, 9, 10) {real, imag} */,
  {32'hc00264eb, 32'hbfe4575b} /* (9, 9, 9) {real, imag} */,
  {32'hc019e2bc, 32'hbfa82735} /* (9, 9, 8) {real, imag} */,
  {32'hc05cd6c3, 32'hbfc3f7eb} /* (9, 9, 7) {real, imag} */,
  {32'h3f3d8c92, 32'hc00ecceb} /* (9, 9, 6) {real, imag} */,
  {32'h4009c474, 32'h3df85654} /* (9, 9, 5) {real, imag} */,
  {32'h3f4b679d, 32'hc0254adf} /* (9, 9, 4) {real, imag} */,
  {32'h3fbe2006, 32'h3d8736b3} /* (9, 9, 3) {real, imag} */,
  {32'h3fe67506, 32'h3fb106da} /* (9, 9, 2) {real, imag} */,
  {32'hbfcb7f9c, 32'hbfb97542} /* (9, 9, 1) {real, imag} */,
  {32'hbfb6e826, 32'h4065a94e} /* (9, 9, 0) {real, imag} */,
  {32'hc07b5bd9, 32'hbfb9f17b} /* (9, 8, 31) {real, imag} */,
  {32'hbff96900, 32'h3fc8e5be} /* (9, 8, 30) {real, imag} */,
  {32'h3f36a20e, 32'h3fc9acf7} /* (9, 8, 29) {real, imag} */,
  {32'hbf1cb02e, 32'hc0050079} /* (9, 8, 28) {real, imag} */,
  {32'h3eb6036f, 32'hbf3087dd} /* (9, 8, 27) {real, imag} */,
  {32'h40b0e5f6, 32'hbf2bf2e6} /* (9, 8, 26) {real, imag} */,
  {32'hbea6aa0b, 32'hbe67cb85} /* (9, 8, 25) {real, imag} */,
  {32'hbf910e8a, 32'hc0033889} /* (9, 8, 24) {real, imag} */,
  {32'h3d4dd413, 32'h3d636c87} /* (9, 8, 23) {real, imag} */,
  {32'h3f804f97, 32'hbf8ff5c4} /* (9, 8, 22) {real, imag} */,
  {32'hc02dff8a, 32'h3fb8c80d} /* (9, 8, 21) {real, imag} */,
  {32'hbeb0af6e, 32'h3f060d19} /* (9, 8, 20) {real, imag} */,
  {32'hbdaf4aaf, 32'h40549abb} /* (9, 8, 19) {real, imag} */,
  {32'h3e93df68, 32'hbf4b01fc} /* (9, 8, 18) {real, imag} */,
  {32'hc037dbc4, 32'h3e9aa30e} /* (9, 8, 17) {real, imag} */,
  {32'hbf745773, 32'hbfd1e5e2} /* (9, 8, 16) {real, imag} */,
  {32'hbf7e410d, 32'hc00661c5} /* (9, 8, 15) {real, imag} */,
  {32'h40192b43, 32'h3e87386a} /* (9, 8, 14) {real, imag} */,
  {32'hbfef0b3d, 32'h3e05fc50} /* (9, 8, 13) {real, imag} */,
  {32'hbfa94c56, 32'h40097a58} /* (9, 8, 12) {real, imag} */,
  {32'h3fcfd71f, 32'h3f844d17} /* (9, 8, 11) {real, imag} */,
  {32'h3ed5e31a, 32'hc0731855} /* (9, 8, 10) {real, imag} */,
  {32'hbece7c44, 32'hc08b5067} /* (9, 8, 9) {real, imag} */,
  {32'hbf4f03b3, 32'h3fb9c8d7} /* (9, 8, 8) {real, imag} */,
  {32'hbf6668d7, 32'hbf9ca17b} /* (9, 8, 7) {real, imag} */,
  {32'hbfe8e60d, 32'h3ef38d90} /* (9, 8, 6) {real, imag} */,
  {32'hc0984ad0, 32'h3fc0987c} /* (9, 8, 5) {real, imag} */,
  {32'h3fa90101, 32'h407ce36d} /* (9, 8, 4) {real, imag} */,
  {32'h3f550148, 32'hbfe3c3f3} /* (9, 8, 3) {real, imag} */,
  {32'h3e0d8906, 32'h3ea2361d} /* (9, 8, 2) {real, imag} */,
  {32'h4058c030, 32'hbf97c090} /* (9, 8, 1) {real, imag} */,
  {32'h40d79b1a, 32'hbf198ed6} /* (9, 8, 0) {real, imag} */,
  {32'hbf3df1dc, 32'h3e87bf23} /* (9, 7, 31) {real, imag} */,
  {32'h4005c648, 32'h404d1323} /* (9, 7, 30) {real, imag} */,
  {32'hc009f2f7, 32'hbfba51ff} /* (9, 7, 29) {real, imag} */,
  {32'h409df532, 32'h3ee83376} /* (9, 7, 28) {real, imag} */,
  {32'h3f376268, 32'hc02a42fd} /* (9, 7, 27) {real, imag} */,
  {32'hbee46497, 32'hc07dfc36} /* (9, 7, 26) {real, imag} */,
  {32'hbf63a57c, 32'hbecbf20c} /* (9, 7, 25) {real, imag} */,
  {32'hc0dd9195, 32'h3c93c59e} /* (9, 7, 24) {real, imag} */,
  {32'h40022acd, 32'hbf34b0f9} /* (9, 7, 23) {real, imag} */,
  {32'hbf8c040f, 32'h3e3961a9} /* (9, 7, 22) {real, imag} */,
  {32'hbea8fa71, 32'hbf76212e} /* (9, 7, 21) {real, imag} */,
  {32'h402a3d88, 32'hc089d349} /* (9, 7, 20) {real, imag} */,
  {32'hbfcca234, 32'h4017d3fc} /* (9, 7, 19) {real, imag} */,
  {32'h3fd8ae0d, 32'hbfd4ef6c} /* (9, 7, 18) {real, imag} */,
  {32'hbfb15951, 32'h3f280180} /* (9, 7, 17) {real, imag} */,
  {32'hbfc5a2ef, 32'h3ef36fae} /* (9, 7, 16) {real, imag} */,
  {32'hbfdb9301, 32'h3f12c45c} /* (9, 7, 15) {real, imag} */,
  {32'h3f7001ec, 32'h3f718d8e} /* (9, 7, 14) {real, imag} */,
  {32'hbf1e3a27, 32'h40a4a81d} /* (9, 7, 13) {real, imag} */,
  {32'hc00bce92, 32'h402f9a16} /* (9, 7, 12) {real, imag} */,
  {32'h3f9d9882, 32'h3f2f6a5d} /* (9, 7, 11) {real, imag} */,
  {32'hbfed6608, 32'hbfb94a08} /* (9, 7, 10) {real, imag} */,
  {32'hc003262e, 32'h3f81e0e7} /* (9, 7, 9) {real, imag} */,
  {32'hbfe6e0cc, 32'hc0991d2c} /* (9, 7, 8) {real, imag} */,
  {32'hbfe6374c, 32'h3f7db322} /* (9, 7, 7) {real, imag} */,
  {32'h3f556517, 32'h3f33b8fa} /* (9, 7, 6) {real, imag} */,
  {32'h3e7a5752, 32'hbfb1cadf} /* (9, 7, 5) {real, imag} */,
  {32'hc02fe68e, 32'h3eaf2795} /* (9, 7, 4) {real, imag} */,
  {32'hbf8afb51, 32'h40186e39} /* (9, 7, 3) {real, imag} */,
  {32'hc056a3a7, 32'hbf45057f} /* (9, 7, 2) {real, imag} */,
  {32'hbf625f1d, 32'hc08ace93} /* (9, 7, 1) {real, imag} */,
  {32'hc0225ccb, 32'h400c7df1} /* (9, 7, 0) {real, imag} */,
  {32'h403ca14f, 32'hbf569625} /* (9, 6, 31) {real, imag} */,
  {32'h402f741c, 32'h4004b847} /* (9, 6, 30) {real, imag} */,
  {32'h3e9dd5a8, 32'h3eddd2a6} /* (9, 6, 29) {real, imag} */,
  {32'hbfbd5c16, 32'hbfb51d7e} /* (9, 6, 28) {real, imag} */,
  {32'h3ecef923, 32'hbf41e415} /* (9, 6, 27) {real, imag} */,
  {32'h3fe628f7, 32'h40a179ce} /* (9, 6, 26) {real, imag} */,
  {32'h3f2db2ff, 32'hbee63088} /* (9, 6, 25) {real, imag} */,
  {32'h3f96f40d, 32'h3f4b4d0e} /* (9, 6, 24) {real, imag} */,
  {32'h4072ffd5, 32'h3f8a8c5d} /* (9, 6, 23) {real, imag} */,
  {32'h3ec369d7, 32'hbd802423} /* (9, 6, 22) {real, imag} */,
  {32'h3ed1990d, 32'hbf04e1c5} /* (9, 6, 21) {real, imag} */,
  {32'hbfd34540, 32'h403fb550} /* (9, 6, 20) {real, imag} */,
  {32'h3eb91dcd, 32'h3f1e5d0b} /* (9, 6, 19) {real, imag} */,
  {32'hc00425e6, 32'h40037391} /* (9, 6, 18) {real, imag} */,
  {32'hbda15e16, 32'hbedb142b} /* (9, 6, 17) {real, imag} */,
  {32'h3fd39da0, 32'hbf50e2be} /* (9, 6, 16) {real, imag} */,
  {32'h3f1a7ebd, 32'h3f7fa184} /* (9, 6, 15) {real, imag} */,
  {32'hbfc108f7, 32'h400be29f} /* (9, 6, 14) {real, imag} */,
  {32'h3fd32a1f, 32'hbf895a10} /* (9, 6, 13) {real, imag} */,
  {32'h407ee619, 32'h3e70f368} /* (9, 6, 12) {real, imag} */,
  {32'hbf3ca313, 32'hc071c129} /* (9, 6, 11) {real, imag} */,
  {32'h3fba306f, 32'hbf188372} /* (9, 6, 10) {real, imag} */,
  {32'h3f3896c3, 32'h3ee328ca} /* (9, 6, 9) {real, imag} */,
  {32'h40021d0f, 32'hbf8d7ee4} /* (9, 6, 8) {real, imag} */,
  {32'h3fd834b4, 32'hbfb39f1a} /* (9, 6, 7) {real, imag} */,
  {32'hbfb9fccc, 32'hc022f7a1} /* (9, 6, 6) {real, imag} */,
  {32'hc023d39b, 32'h3f19a6e6} /* (9, 6, 5) {real, imag} */,
  {32'hc01d2098, 32'hc03cd6fc} /* (9, 6, 4) {real, imag} */,
  {32'h3f36c393, 32'h3eaddc1d} /* (9, 6, 3) {real, imag} */,
  {32'h3f9989d2, 32'h40a0dfbe} /* (9, 6, 2) {real, imag} */,
  {32'h403c063b, 32'hbf669e22} /* (9, 6, 1) {real, imag} */,
  {32'hc076aa4f, 32'h3ec47798} /* (9, 6, 0) {real, imag} */,
  {32'hbe6f2eba, 32'hc002c889} /* (9, 5, 31) {real, imag} */,
  {32'hc04bac71, 32'h400075f2} /* (9, 5, 30) {real, imag} */,
  {32'hc012c316, 32'hc05094f8} /* (9, 5, 29) {real, imag} */,
  {32'h3ff02108, 32'hbfba0b79} /* (9, 5, 28) {real, imag} */,
  {32'h3ed14f0b, 32'h4006b1ed} /* (9, 5, 27) {real, imag} */,
  {32'h3fbf5924, 32'hbe61f20b} /* (9, 5, 26) {real, imag} */,
  {32'h3e129b63, 32'h400106e8} /* (9, 5, 25) {real, imag} */,
  {32'hbfcd482e, 32'hc0a0859f} /* (9, 5, 24) {real, imag} */,
  {32'hbfc3ffad, 32'hc03bff91} /* (9, 5, 23) {real, imag} */,
  {32'h3fe82b0c, 32'hbe09f7dd} /* (9, 5, 22) {real, imag} */,
  {32'hbfdb40b8, 32'h3f37eb17} /* (9, 5, 21) {real, imag} */,
  {32'hbce4a788, 32'h3fe2e1ac} /* (9, 5, 20) {real, imag} */,
  {32'h40a0aef1, 32'hc0165597} /* (9, 5, 19) {real, imag} */,
  {32'h4002498d, 32'hbe8e77f6} /* (9, 5, 18) {real, imag} */,
  {32'h3f1c9598, 32'hbf3427d8} /* (9, 5, 17) {real, imag} */,
  {32'hbeac56ea, 32'hbea25177} /* (9, 5, 16) {real, imag} */,
  {32'h3fb8b85d, 32'hc0550381} /* (9, 5, 15) {real, imag} */,
  {32'hbea96874, 32'h3f51a117} /* (9, 5, 14) {real, imag} */,
  {32'h40102ddb, 32'hbf993dde} /* (9, 5, 13) {real, imag} */,
  {32'h3fd949df, 32'h3f4478ea} /* (9, 5, 12) {real, imag} */,
  {32'hc0283eec, 32'hc0b13eea} /* (9, 5, 11) {real, imag} */,
  {32'hbe8b0948, 32'h3ea871da} /* (9, 5, 10) {real, imag} */,
  {32'h403293e9, 32'hc008045d} /* (9, 5, 9) {real, imag} */,
  {32'h3e2dbcb3, 32'hbf6d4a2b} /* (9, 5, 8) {real, imag} */,
  {32'h403e23d5, 32'hbe47d633} /* (9, 5, 7) {real, imag} */,
  {32'hc06c66a5, 32'hbe7aac49} /* (9, 5, 6) {real, imag} */,
  {32'h4014c1e1, 32'hbddab100} /* (9, 5, 5) {real, imag} */,
  {32'hbfc096d6, 32'h401b6a1b} /* (9, 5, 4) {real, imag} */,
  {32'hc04ab467, 32'hbec9c2c0} /* (9, 5, 3) {real, imag} */,
  {32'h3fb3450d, 32'hc01838b8} /* (9, 5, 2) {real, imag} */,
  {32'h3fddb791, 32'hbf3754df} /* (9, 5, 1) {real, imag} */,
  {32'h4029aef4, 32'hc03d7f3b} /* (9, 5, 0) {real, imag} */,
  {32'h3ff0ade2, 32'h3f894f97} /* (9, 4, 31) {real, imag} */,
  {32'h3fd7c9d6, 32'hbfeec363} /* (9, 4, 30) {real, imag} */,
  {32'h3f23121f, 32'h408ab943} /* (9, 4, 29) {real, imag} */,
  {32'h40007c0c, 32'hbef1241d} /* (9, 4, 28) {real, imag} */,
  {32'hc072ed4d, 32'h4099880e} /* (9, 4, 27) {real, imag} */,
  {32'h3f513d3a, 32'h402c195a} /* (9, 4, 26) {real, imag} */,
  {32'h40b9470c, 32'h3f8e863e} /* (9, 4, 25) {real, imag} */,
  {32'hc014912e, 32'h3fcf76cc} /* (9, 4, 24) {real, imag} */,
  {32'hbff022d4, 32'hbfc33b4a} /* (9, 4, 23) {real, imag} */,
  {32'hc0600d20, 32'hc00f678d} /* (9, 4, 22) {real, imag} */,
  {32'h3f363454, 32'hbfe2c579} /* (9, 4, 21) {real, imag} */,
  {32'h3f21fea5, 32'h4014fb1d} /* (9, 4, 20) {real, imag} */,
  {32'h3d95979c, 32'h4021d9e9} /* (9, 4, 19) {real, imag} */,
  {32'h3f9c1a1b, 32'h3f8f23d5} /* (9, 4, 18) {real, imag} */,
  {32'hbfce91d2, 32'h3f351988} /* (9, 4, 17) {real, imag} */,
  {32'hbf09c9f0, 32'h3f443f13} /* (9, 4, 16) {real, imag} */,
  {32'hc01a2f13, 32'h3f91cf40} /* (9, 4, 15) {real, imag} */,
  {32'h3f492bfb, 32'hbf7e170f} /* (9, 4, 14) {real, imag} */,
  {32'h3fba47ef, 32'h3fc6594d} /* (9, 4, 13) {real, imag} */,
  {32'hbef2e2dd, 32'hbfebfb49} /* (9, 4, 12) {real, imag} */,
  {32'h408531b1, 32'hbfbb0f39} /* (9, 4, 11) {real, imag} */,
  {32'h3fad266e, 32'hc005ebd4} /* (9, 4, 10) {real, imag} */,
  {32'h3fda0671, 32'h40292900} /* (9, 4, 9) {real, imag} */,
  {32'hbf998bae, 32'hbf920c4f} /* (9, 4, 8) {real, imag} */,
  {32'h3f59c70c, 32'hbfccdbdc} /* (9, 4, 7) {real, imag} */,
  {32'hc0784cf0, 32'h401fade9} /* (9, 4, 6) {real, imag} */,
  {32'hbf82a5df, 32'hbf3a1b57} /* (9, 4, 5) {real, imag} */,
  {32'hbf747114, 32'h3f8a411f} /* (9, 4, 4) {real, imag} */,
  {32'h4083391c, 32'h3e5633e7} /* (9, 4, 3) {real, imag} */,
  {32'hbd6f8a91, 32'h3f654a3d} /* (9, 4, 2) {real, imag} */,
  {32'hbe443d65, 32'h3fb28a2a} /* (9, 4, 1) {real, imag} */,
  {32'h3e3e2208, 32'h3f032feb} /* (9, 4, 0) {real, imag} */,
  {32'hbdea6b3b, 32'h3e225eab} /* (9, 3, 31) {real, imag} */,
  {32'hbea7d01e, 32'h3f9979e6} /* (9, 3, 30) {real, imag} */,
  {32'h406d8087, 32'h3efe7171} /* (9, 3, 29) {real, imag} */,
  {32'hbdac85c4, 32'h3f7f6ce6} /* (9, 3, 28) {real, imag} */,
  {32'h3f5302ff, 32'h3f8134fb} /* (9, 3, 27) {real, imag} */,
  {32'h3f881e1f, 32'hc0236057} /* (9, 3, 26) {real, imag} */,
  {32'h3fd6c827, 32'h3ff7427a} /* (9, 3, 25) {real, imag} */,
  {32'hbbe86860, 32'h3f0e52b9} /* (9, 3, 24) {real, imag} */,
  {32'hbfaaa029, 32'hc07008b7} /* (9, 3, 23) {real, imag} */,
  {32'hc03c504f, 32'h3db1a6bb} /* (9, 3, 22) {real, imag} */,
  {32'h3f0bf89d, 32'hbf926f3a} /* (9, 3, 21) {real, imag} */,
  {32'h3e2141a4, 32'h3fa4d060} /* (9, 3, 20) {real, imag} */,
  {32'h4022bbf5, 32'hbe5c62a2} /* (9, 3, 19) {real, imag} */,
  {32'hc01c6b5a, 32'h3e2bd09e} /* (9, 3, 18) {real, imag} */,
  {32'h400a3db8, 32'hbf0e127a} /* (9, 3, 17) {real, imag} */,
  {32'hbea4cca3, 32'h3f44a1b1} /* (9, 3, 16) {real, imag} */,
  {32'hbf33b5b9, 32'h400846ad} /* (9, 3, 15) {real, imag} */,
  {32'hc033db19, 32'h3f7a9d28} /* (9, 3, 14) {real, imag} */,
  {32'h3f191754, 32'hc0a7dea3} /* (9, 3, 13) {real, imag} */,
  {32'h3ff64458, 32'hbfa251ae} /* (9, 3, 12) {real, imag} */,
  {32'hbf3b7e87, 32'h40670d4c} /* (9, 3, 11) {real, imag} */,
  {32'hbe3e2f17, 32'h3e986382} /* (9, 3, 10) {real, imag} */,
  {32'hbf361f91, 32'hbd75c4b8} /* (9, 3, 9) {real, imag} */,
  {32'h3ffc95c5, 32'h3f08baad} /* (9, 3, 8) {real, imag} */,
  {32'hc005189a, 32'h3ff818b5} /* (9, 3, 7) {real, imag} */,
  {32'h40196575, 32'hc088867a} /* (9, 3, 6) {real, imag} */,
  {32'h40334283, 32'h3ea5eeda} /* (9, 3, 5) {real, imag} */,
  {32'hbed41e36, 32'h40581431} /* (9, 3, 4) {real, imag} */,
  {32'h404a9674, 32'hbf853b92} /* (9, 3, 3) {real, imag} */,
  {32'hc053c5ba, 32'hc0bd31c7} /* (9, 3, 2) {real, imag} */,
  {32'hbe8bf30d, 32'hbfb4151d} /* (9, 3, 1) {real, imag} */,
  {32'h4045de60, 32'hbeef567a} /* (9, 3, 0) {real, imag} */,
  {32'h3f93fb79, 32'hc05db407} /* (9, 2, 31) {real, imag} */,
  {32'hbfb882e9, 32'h40be8d4b} /* (9, 2, 30) {real, imag} */,
  {32'hc0a5d16b, 32'h3b7376c4} /* (9, 2, 29) {real, imag} */,
  {32'hc03396bf, 32'hc0850785} /* (9, 2, 28) {real, imag} */,
  {32'h3d92a698, 32'h3f83ffb5} /* (9, 2, 27) {real, imag} */,
  {32'h3fbe06ef, 32'h40424e9b} /* (9, 2, 26) {real, imag} */,
  {32'h3f2c78b1, 32'h4009e451} /* (9, 2, 25) {real, imag} */,
  {32'hbfa14203, 32'hbf30b40a} /* (9, 2, 24) {real, imag} */,
  {32'hbf7f47e2, 32'hbf6c0d50} /* (9, 2, 23) {real, imag} */,
  {32'h405d11a7, 32'h3fa82d3f} /* (9, 2, 22) {real, imag} */,
  {32'h3fdbb9c1, 32'h3f524e41} /* (9, 2, 21) {real, imag} */,
  {32'h3eae206b, 32'hc0182c87} /* (9, 2, 20) {real, imag} */,
  {32'hc04e2125, 32'h3fb61fc7} /* (9, 2, 19) {real, imag} */,
  {32'h3f9da7fa, 32'h4029cd58} /* (9, 2, 18) {real, imag} */,
  {32'hbf0cad44, 32'h3e9ed13d} /* (9, 2, 17) {real, imag} */,
  {32'h3fa7fd29, 32'hbe8b7be0} /* (9, 2, 16) {real, imag} */,
  {32'h403496e8, 32'h40148395} /* (9, 2, 15) {real, imag} */,
  {32'h401d89c3, 32'hbf065fde} /* (9, 2, 14) {real, imag} */,
  {32'hbf581265, 32'hbf90145d} /* (9, 2, 13) {real, imag} */,
  {32'h3f94f51a, 32'hbf10310a} /* (9, 2, 12) {real, imag} */,
  {32'hc04393b3, 32'hbfbce410} /* (9, 2, 11) {real, imag} */,
  {32'h402b98b8, 32'h401af434} /* (9, 2, 10) {real, imag} */,
  {32'hbda36622, 32'hbfc1b402} /* (9, 2, 9) {real, imag} */,
  {32'hc05ada4d, 32'h3f8eeda7} /* (9, 2, 8) {real, imag} */,
  {32'h408789f5, 32'hbf6d32a2} /* (9, 2, 7) {real, imag} */,
  {32'h40226ac5, 32'h3f9ff0c2} /* (9, 2, 6) {real, imag} */,
  {32'hc02b3f91, 32'hbf8f3f1f} /* (9, 2, 5) {real, imag} */,
  {32'h3ff2b67b, 32'hc08f2e1b} /* (9, 2, 4) {real, imag} */,
  {32'hc00e4f6d, 32'h4071f8f4} /* (9, 2, 3) {real, imag} */,
  {32'h3fe1a416, 32'h40ee9c4a} /* (9, 2, 2) {real, imag} */,
  {32'h406c017c, 32'hc0820344} /* (9, 2, 1) {real, imag} */,
  {32'h3f53835d, 32'hc0840c4a} /* (9, 2, 0) {real, imag} */,
  {32'hbf94afa2, 32'h40891c5a} /* (9, 1, 31) {real, imag} */,
  {32'h4022aa49, 32'hc05c953f} /* (9, 1, 30) {real, imag} */,
  {32'h3e3f5e91, 32'hbda627d4} /* (9, 1, 29) {real, imag} */,
  {32'hbc9e394e, 32'h3fb4ca3b} /* (9, 1, 28) {real, imag} */,
  {32'h3f6715bf, 32'h3fc85114} /* (9, 1, 27) {real, imag} */,
  {32'hc0812aa1, 32'h403a4fc4} /* (9, 1, 26) {real, imag} */,
  {32'hc02c0a97, 32'h3f99fb0c} /* (9, 1, 25) {real, imag} */,
  {32'h3f3b8934, 32'hbfa29869} /* (9, 1, 24) {real, imag} */,
  {32'h3ea061f3, 32'hbfbeebf1} /* (9, 1, 23) {real, imag} */,
  {32'h401a184a, 32'hbfac0cde} /* (9, 1, 22) {real, imag} */,
  {32'h3fe0c154, 32'h3f082c7c} /* (9, 1, 21) {real, imag} */,
  {32'hc0491cbc, 32'hbf334756} /* (9, 1, 20) {real, imag} */,
  {32'h3fc952e5, 32'hbfdfeb82} /* (9, 1, 19) {real, imag} */,
  {32'h3f63549e, 32'hbf683da2} /* (9, 1, 18) {real, imag} */,
  {32'h3f2339fb, 32'h3fae282e} /* (9, 1, 17) {real, imag} */,
  {32'h3f2cd194, 32'hbfebdbbf} /* (9, 1, 16) {real, imag} */,
  {32'h3f2d60eb, 32'hbdb55d04} /* (9, 1, 15) {real, imag} */,
  {32'hbfbeeee5, 32'hbf3a040e} /* (9, 1, 14) {real, imag} */,
  {32'hbebbb032, 32'hc03796ca} /* (9, 1, 13) {real, imag} */,
  {32'hbf999226, 32'h3eeb1789} /* (9, 1, 12) {real, imag} */,
  {32'hbfbcb05e, 32'hbcfb0928} /* (9, 1, 11) {real, imag} */,
  {32'hbfca08bf, 32'h3fe70597} /* (9, 1, 10) {real, imag} */,
  {32'h3fae36fe, 32'h403b26a2} /* (9, 1, 9) {real, imag} */,
  {32'hc03fd469, 32'h40be2e36} /* (9, 1, 8) {real, imag} */,
  {32'h3ff9993d, 32'h3fd39f1b} /* (9, 1, 7) {real, imag} */,
  {32'h3fd5afbc, 32'hbfc8f943} /* (9, 1, 6) {real, imag} */,
  {32'h402a5695, 32'hbefb70a5} /* (9, 1, 5) {real, imag} */,
  {32'hbf1c9d85, 32'h4017bdc4} /* (9, 1, 4) {real, imag} */,
  {32'h3ed4e7bd, 32'hc10f0324} /* (9, 1, 3) {real, imag} */,
  {32'h40ab1cac, 32'hc078dc3d} /* (9, 1, 2) {real, imag} */,
  {32'hc0b610c6, 32'hbed07cdb} /* (9, 1, 1) {real, imag} */,
  {32'hc0a72a0d, 32'hc017e4c4} /* (9, 1, 0) {real, imag} */,
  {32'hc00ee180, 32'h40837ce9} /* (9, 0, 31) {real, imag} */,
  {32'h3f8ecfa0, 32'hbf6f1d6f} /* (9, 0, 30) {real, imag} */,
  {32'hc032302b, 32'h3f1e4a15} /* (9, 0, 29) {real, imag} */,
  {32'h3fee085d, 32'h3eb5ab91} /* (9, 0, 28) {real, imag} */,
  {32'h3fede971, 32'hbe9e9138} /* (9, 0, 27) {real, imag} */,
  {32'hc02adc2c, 32'h3f1dc253} /* (9, 0, 26) {real, imag} */,
  {32'h3f1efe38, 32'h3fa86126} /* (9, 0, 25) {real, imag} */,
  {32'hc0503152, 32'hc068e117} /* (9, 0, 24) {real, imag} */,
  {32'h3f751e28, 32'hc03b4a7d} /* (9, 0, 23) {real, imag} */,
  {32'h409895ca, 32'hbf66736f} /* (9, 0, 22) {real, imag} */,
  {32'hbf8fa1fc, 32'h3e2b4619} /* (9, 0, 21) {real, imag} */,
  {32'h3e2b9282, 32'hbd2f7457} /* (9, 0, 20) {real, imag} */,
  {32'h40262e93, 32'hbf25c551} /* (9, 0, 19) {real, imag} */,
  {32'hbfb2dcd6, 32'hbf84ccad} /* (9, 0, 18) {real, imag} */,
  {32'hbf131872, 32'h3f10de1b} /* (9, 0, 17) {real, imag} */,
  {32'h3ef93f34, 32'hbfc5475c} /* (9, 0, 16) {real, imag} */,
  {32'hbe852b95, 32'hbf3727cc} /* (9, 0, 15) {real, imag} */,
  {32'h3fae65eb, 32'h3fef1c08} /* (9, 0, 14) {real, imag} */,
  {32'hbffb400d, 32'h3f303189} /* (9, 0, 13) {real, imag} */,
  {32'h3ec04596, 32'h3f8b6c48} /* (9, 0, 12) {real, imag} */,
  {32'hbf54bb1b, 32'hc01e43ac} /* (9, 0, 11) {real, imag} */,
  {32'hbfc46b08, 32'h4007097f} /* (9, 0, 10) {real, imag} */,
  {32'h3fae1b9e, 32'hbe91d2c3} /* (9, 0, 9) {real, imag} */,
  {32'h40654fa5, 32'h40be5f0e} /* (9, 0, 8) {real, imag} */,
  {32'hbfe691ea, 32'h400263d2} /* (9, 0, 7) {real, imag} */,
  {32'hbf1b0960, 32'hc02e1c5c} /* (9, 0, 6) {real, imag} */,
  {32'h401bd1ef, 32'hbfcb4204} /* (9, 0, 5) {real, imag} */,
  {32'hc02c8495, 32'h40153e38} /* (9, 0, 4) {real, imag} */,
  {32'h40afc7ae, 32'hbf06c377} /* (9, 0, 3) {real, imag} */,
  {32'hc0021e29, 32'hbf03f796} /* (9, 0, 2) {real, imag} */,
  {32'hc09a5d46, 32'hc015fe48} /* (9, 0, 1) {real, imag} */,
  {32'hbf3cbe3f, 32'h40daa393} /* (9, 0, 0) {real, imag} */,
  {32'hc0b68caa, 32'h41dcba48} /* (8, 31, 31) {real, imag} */,
  {32'hc0017c6b, 32'hc191019a} /* (8, 31, 30) {real, imag} */,
  {32'hbe699550, 32'h3f353691} /* (8, 31, 29) {real, imag} */,
  {32'h4057a30f, 32'hc02a42f5} /* (8, 31, 28) {real, imag} */,
  {32'h3f68f5d2, 32'hc0971572} /* (8, 31, 27) {real, imag} */,
  {32'hbee83711, 32'h3e61a2ea} /* (8, 31, 26) {real, imag} */,
  {32'hbfa9ab52, 32'h3e77cb01} /* (8, 31, 25) {real, imag} */,
  {32'hc054765d, 32'hc08f18a2} /* (8, 31, 24) {real, imag} */,
  {32'hc05525c1, 32'hbf89d94f} /* (8, 31, 23) {real, imag} */,
  {32'h405be2bd, 32'h402bd702} /* (8, 31, 22) {real, imag} */,
  {32'h3e8b4a9d, 32'hc07772c6} /* (8, 31, 21) {real, imag} */,
  {32'hc01fc3b8, 32'hbe750a29} /* (8, 31, 20) {real, imag} */,
  {32'hbe5599f4, 32'h3faff77f} /* (8, 31, 19) {real, imag} */,
  {32'hbf7e1054, 32'h3c924251} /* (8, 31, 18) {real, imag} */,
  {32'h409cca41, 32'hbdba117c} /* (8, 31, 17) {real, imag} */,
  {32'hbf927fe3, 32'h3f96aff4} /* (8, 31, 16) {real, imag} */,
  {32'hbf5f97ad, 32'hbf733048} /* (8, 31, 15) {real, imag} */,
  {32'h3f7d2d34, 32'h407dab9e} /* (8, 31, 14) {real, imag} */,
  {32'h3e14c8ed, 32'hbfd4ac8c} /* (8, 31, 13) {real, imag} */,
  {32'h3e945379, 32'h3fa1aab1} /* (8, 31, 12) {real, imag} */,
  {32'hbf8aa415, 32'h3fb737a3} /* (8, 31, 11) {real, imag} */,
  {32'hbe7f9e17, 32'h3dbb3276} /* (8, 31, 10) {real, imag} */,
  {32'h3f3cb06d, 32'hc087c4d2} /* (8, 31, 9) {real, imag} */,
  {32'h3f1ac76e, 32'h3fd8a2a9} /* (8, 31, 8) {real, imag} */,
  {32'h4042a95d, 32'h3f0a3d47} /* (8, 31, 7) {real, imag} */,
  {32'hc012d13f, 32'hbf29efec} /* (8, 31, 6) {real, imag} */,
  {32'h4020d0b0, 32'hc0d14ab4} /* (8, 31, 5) {real, imag} */,
  {32'h3fb3eba7, 32'h40750f12} /* (8, 31, 4) {real, imag} */,
  {32'h3f5fb74e, 32'hbf53c37e} /* (8, 31, 3) {real, imag} */,
  {32'h40fa8ebe, 32'hc0b3c9b3} /* (8, 31, 2) {real, imag} */,
  {32'hc127fe79, 32'h4130aa59} /* (8, 31, 1) {real, imag} */,
  {32'hc10d65e9, 32'h4186824f} /* (8, 31, 0) {real, imag} */,
  {32'h413ad087, 32'hbf9e23e5} /* (8, 30, 31) {real, imag} */,
  {32'hc136d204, 32'h41632eec} /* (8, 30, 30) {real, imag} */,
  {32'h407bf02d, 32'h3faf7adc} /* (8, 30, 29) {real, imag} */,
  {32'h4086965f, 32'hbff0e715} /* (8, 30, 28) {real, imag} */,
  {32'h40183e01, 32'h40e08e3a} /* (8, 30, 27) {real, imag} */,
  {32'h3e4d7df5, 32'h3f186f2a} /* (8, 30, 26) {real, imag} */,
  {32'hbfb69288, 32'h402da91c} /* (8, 30, 25) {real, imag} */,
  {32'hbf015189, 32'h40883606} /* (8, 30, 24) {real, imag} */,
  {32'hbdac4e0e, 32'hbf832ec8} /* (8, 30, 23) {real, imag} */,
  {32'hbfd7ba62, 32'h3f06cfc8} /* (8, 30, 22) {real, imag} */,
  {32'h3f8b0811, 32'h3eecbb8c} /* (8, 30, 21) {real, imag} */,
  {32'h402c2b10, 32'hc02f0620} /* (8, 30, 20) {real, imag} */,
  {32'h3f1a376c, 32'hbd506f5f} /* (8, 30, 19) {real, imag} */,
  {32'hbea0f244, 32'hbeb811ff} /* (8, 30, 18) {real, imag} */,
  {32'hbf2dc6a5, 32'h3e99ca75} /* (8, 30, 17) {real, imag} */,
  {32'h3f5a4ab6, 32'hbf90c299} /* (8, 30, 16) {real, imag} */,
  {32'hbec70f61, 32'h3ca71186} /* (8, 30, 15) {real, imag} */,
  {32'h3f597afe, 32'h3fdd4f33} /* (8, 30, 14) {real, imag} */,
  {32'h402549c6, 32'h3fe737f8} /* (8, 30, 13) {real, imag} */,
  {32'hbf4b64ec, 32'h4086130c} /* (8, 30, 12) {real, imag} */,
  {32'h3f80d480, 32'hbf7d7657} /* (8, 30, 11) {real, imag} */,
  {32'h3f977384, 32'h3fa257db} /* (8, 30, 10) {real, imag} */,
  {32'hbfa4da82, 32'hbf8d4278} /* (8, 30, 9) {real, imag} */,
  {32'hc0e5cc89, 32'h3f8b7909} /* (8, 30, 8) {real, imag} */,
  {32'h3f3991d9, 32'hbe6eb536} /* (8, 30, 7) {real, imag} */,
  {32'h403be27b, 32'hc094c0e4} /* (8, 30, 6) {real, imag} */,
  {32'hc0cadcfa, 32'h3f560c02} /* (8, 30, 5) {real, imag} */,
  {32'h3fe0ca6b, 32'h3fee1a85} /* (8, 30, 4) {real, imag} */,
  {32'h404192d0, 32'hbfe30827} /* (8, 30, 3) {real, imag} */,
  {32'hc11771e0, 32'h4052697c} /* (8, 30, 2) {real, imag} */,
  {32'h411fc6b6, 32'hc18ec8ab} /* (8, 30, 1) {real, imag} */,
  {32'h4093fb62, 32'hc12332ec} /* (8, 30, 0) {real, imag} */,
  {32'hbfaac526, 32'h4027b645} /* (8, 29, 31) {real, imag} */,
  {32'hc018f632, 32'hbfcf4d99} /* (8, 29, 30) {real, imag} */,
  {32'h4079923f, 32'hc06f860d} /* (8, 29, 29) {real, imag} */,
  {32'h4016551b, 32'hc0162b3a} /* (8, 29, 28) {real, imag} */,
  {32'h3f0b88a5, 32'h40286c7b} /* (8, 29, 27) {real, imag} */,
  {32'hbffd03ab, 32'hbe830eb3} /* (8, 29, 26) {real, imag} */,
  {32'hc000cfd4, 32'h3e84f345} /* (8, 29, 25) {real, imag} */,
  {32'h3fe5b1a9, 32'hbe073605} /* (8, 29, 24) {real, imag} */,
  {32'h3ef48cd2, 32'h3d93712c} /* (8, 29, 23) {real, imag} */,
  {32'h3ed63b64, 32'h3f260a6f} /* (8, 29, 22) {real, imag} */,
  {32'hbf131d2c, 32'h3f5f2302} /* (8, 29, 21) {real, imag} */,
  {32'hc0083636, 32'hc04d6ff2} /* (8, 29, 20) {real, imag} */,
  {32'hc02e29b4, 32'hbfb82e6a} /* (8, 29, 19) {real, imag} */,
  {32'h3e8ed735, 32'h40375bfc} /* (8, 29, 18) {real, imag} */,
  {32'h3fa0c5ea, 32'hc02d8c78} /* (8, 29, 17) {real, imag} */,
  {32'hbf6b8482, 32'hbf22fe9a} /* (8, 29, 16) {real, imag} */,
  {32'h3e08aa62, 32'hbfa10f13} /* (8, 29, 15) {real, imag} */,
  {32'hc03943a1, 32'h40053c07} /* (8, 29, 14) {real, imag} */,
  {32'hbfd11528, 32'h3f38adf6} /* (8, 29, 13) {real, imag} */,
  {32'hbe4d225d, 32'hbffa59c6} /* (8, 29, 12) {real, imag} */,
  {32'hc0391be9, 32'h400bbea3} /* (8, 29, 11) {real, imag} */,
  {32'h405fc0b6, 32'hbd8d4602} /* (8, 29, 10) {real, imag} */,
  {32'h3f71f7fc, 32'hc023b259} /* (8, 29, 9) {real, imag} */,
  {32'hbfe76184, 32'hc0534954} /* (8, 29, 8) {real, imag} */,
  {32'hbfe6131c, 32'hbf5d336f} /* (8, 29, 7) {real, imag} */,
  {32'h4079c33d, 32'h403ed1e7} /* (8, 29, 6) {real, imag} */,
  {32'h4027ca12, 32'h3d252fcd} /* (8, 29, 5) {real, imag} */,
  {32'h3fbc2c84, 32'h40d97ae1} /* (8, 29, 4) {real, imag} */,
  {32'hc04080a8, 32'hc0e52a61} /* (8, 29, 3) {real, imag} */,
  {32'hc00b38b9, 32'h3ffc2f8c} /* (8, 29, 2) {real, imag} */,
  {32'h40a71ba9, 32'h3f3618d6} /* (8, 29, 1) {real, imag} */,
  {32'h401b26a6, 32'h3f8d57a3} /* (8, 29, 0) {real, imag} */,
  {32'hbffbbe2b, 32'h40fd4999} /* (8, 28, 31) {real, imag} */,
  {32'hc015f9c4, 32'hc0cc05c6} /* (8, 28, 30) {real, imag} */,
  {32'hbf963530, 32'h40a48062} /* (8, 28, 29) {real, imag} */,
  {32'h405c0091, 32'h408a42c9} /* (8, 28, 28) {real, imag} */,
  {32'h3fa91cf5, 32'hbe969e2d} /* (8, 28, 27) {real, imag} */,
  {32'h3f0b96f1, 32'h3f0c9868} /* (8, 28, 26) {real, imag} */,
  {32'h3f492778, 32'h40a98ea8} /* (8, 28, 25) {real, imag} */,
  {32'h3eb959ad, 32'hbe54f482} /* (8, 28, 24) {real, imag} */,
  {32'hc0a1fa89, 32'hbfff493b} /* (8, 28, 23) {real, imag} */,
  {32'h3fd24613, 32'hbf125cb5} /* (8, 28, 22) {real, imag} */,
  {32'hc06b04b5, 32'hc08aec72} /* (8, 28, 21) {real, imag} */,
  {32'hbf863f88, 32'h3f9d01c7} /* (8, 28, 20) {real, imag} */,
  {32'h3f9f49c8, 32'h3fd8b267} /* (8, 28, 19) {real, imag} */,
  {32'hbe534efd, 32'hc024f027} /* (8, 28, 18) {real, imag} */,
  {32'h3ed9593c, 32'hbf0483d6} /* (8, 28, 17) {real, imag} */,
  {32'h3e917385, 32'h3f458cb4} /* (8, 28, 16) {real, imag} */,
  {32'hbf2e9fe5, 32'hbfd5aa5a} /* (8, 28, 15) {real, imag} */,
  {32'hbfc913db, 32'hc0040dfc} /* (8, 28, 14) {real, imag} */,
  {32'h3f3cc48b, 32'h3f7bda8a} /* (8, 28, 13) {real, imag} */,
  {32'hbf1ada8e, 32'hbfa8e3fb} /* (8, 28, 12) {real, imag} */,
  {32'hbf52552a, 32'h3f19328c} /* (8, 28, 11) {real, imag} */,
  {32'h3ec827b4, 32'h4007e35f} /* (8, 28, 10) {real, imag} */,
  {32'h3f94da11, 32'h3f70f248} /* (8, 28, 9) {real, imag} */,
  {32'h401bf96d, 32'h3f89a9db} /* (8, 28, 8) {real, imag} */,
  {32'h3fad5868, 32'hbde11b4e} /* (8, 28, 7) {real, imag} */,
  {32'h3f88c44f, 32'hbf1395d3} /* (8, 28, 6) {real, imag} */,
  {32'h3eb1cf76, 32'h40d8b883} /* (8, 28, 5) {real, imag} */,
  {32'hbffa6fef, 32'h3d93ebfb} /* (8, 28, 4) {real, imag} */,
  {32'h3fac6465, 32'h40a7c524} /* (8, 28, 3) {real, imag} */,
  {32'h3fa71b21, 32'hc0ca7a8e} /* (8, 28, 2) {real, imag} */,
  {32'hbdc8299f, 32'h402be5ae} /* (8, 28, 1) {real, imag} */,
  {32'hbe22dbef, 32'h3f7523e4} /* (8, 28, 0) {real, imag} */,
  {32'hbfe92936, 32'hbf763e7c} /* (8, 27, 31) {real, imag} */,
  {32'h3f936aeb, 32'h405a7ffa} /* (8, 27, 30) {real, imag} */,
  {32'h3e3cd7b7, 32'hbca2fab1} /* (8, 27, 29) {real, imag} */,
  {32'h4040f972, 32'h406c2ede} /* (8, 27, 28) {real, imag} */,
  {32'h3f9fd05c, 32'hbdf9f9d8} /* (8, 27, 27) {real, imag} */,
  {32'h3f6e7bdb, 32'hbe4937ee} /* (8, 27, 26) {real, imag} */,
  {32'hc03df135, 32'hbfbe2a06} /* (8, 27, 25) {real, imag} */,
  {32'h4032c488, 32'h4001635a} /* (8, 27, 24) {real, imag} */,
  {32'h3f37444a, 32'hbf556545} /* (8, 27, 23) {real, imag} */,
  {32'hbf20c1d9, 32'h3c7a2994} /* (8, 27, 22) {real, imag} */,
  {32'h3fa5441f, 32'h3eee09e5} /* (8, 27, 21) {real, imag} */,
  {32'h404c7ec2, 32'hbec7c731} /* (8, 27, 20) {real, imag} */,
  {32'hc0977cd8, 32'h3ecf434f} /* (8, 27, 19) {real, imag} */,
  {32'hbfaa2d50, 32'hbfc4cfb2} /* (8, 27, 18) {real, imag} */,
  {32'hbf0f88a0, 32'h3fff02f3} /* (8, 27, 17) {real, imag} */,
  {32'h3fdb15c3, 32'hc06f5f64} /* (8, 27, 16) {real, imag} */,
  {32'hbf13e13b, 32'h3f47d754} /* (8, 27, 15) {real, imag} */,
  {32'hbfb7beac, 32'hbfcadea2} /* (8, 27, 14) {real, imag} */,
  {32'hbeb22f7a, 32'h3f348d97} /* (8, 27, 13) {real, imag} */,
  {32'hbfc28a58, 32'hbf0ee336} /* (8, 27, 12) {real, imag} */,
  {32'h3f1e0b19, 32'hc02db0c7} /* (8, 27, 11) {real, imag} */,
  {32'hbd595f00, 32'h3e65444e} /* (8, 27, 10) {real, imag} */,
  {32'h3f1c34c9, 32'h3dc1d931} /* (8, 27, 9) {real, imag} */,
  {32'hbf9ea7a0, 32'h3f8aac5f} /* (8, 27, 8) {real, imag} */,
  {32'h4021b97e, 32'hbf83ad38} /* (8, 27, 7) {real, imag} */,
  {32'hbf95c49b, 32'hbf96c37e} /* (8, 27, 6) {real, imag} */,
  {32'hc0287bfe, 32'hbfa2f215} /* (8, 27, 5) {real, imag} */,
  {32'h3ff07814, 32'h3ee0116d} /* (8, 27, 4) {real, imag} */,
  {32'h3f505465, 32'hbec1bb26} /* (8, 27, 3) {real, imag} */,
  {32'hbff5c55a, 32'h404f2798} /* (8, 27, 2) {real, imag} */,
  {32'h4006fdba, 32'hc0534277} /* (8, 27, 1) {real, imag} */,
  {32'h3f5fd3f5, 32'hc0296de4} /* (8, 27, 0) {real, imag} */,
  {32'h3f39593f, 32'h404780cd} /* (8, 26, 31) {real, imag} */,
  {32'h3f5886f8, 32'hbedfa4fd} /* (8, 26, 30) {real, imag} */,
  {32'h403abadd, 32'h3f8695c7} /* (8, 26, 29) {real, imag} */,
  {32'h4019a69b, 32'hbf3147fd} /* (8, 26, 28) {real, imag} */,
  {32'h3ea36240, 32'h4086f02b} /* (8, 26, 27) {real, imag} */,
  {32'h3f897e95, 32'h3fd39486} /* (8, 26, 26) {real, imag} */,
  {32'hbd449725, 32'hc07d8057} /* (8, 26, 25) {real, imag} */,
  {32'hbf63154e, 32'hbdffbaf6} /* (8, 26, 24) {real, imag} */,
  {32'h3e7372f4, 32'hbf4964f9} /* (8, 26, 23) {real, imag} */,
  {32'hc0203493, 32'hc04d0d31} /* (8, 26, 22) {real, imag} */,
  {32'hc08be198, 32'hbfab74bc} /* (8, 26, 21) {real, imag} */,
  {32'h3f89f65b, 32'hbf9c2a54} /* (8, 26, 20) {real, imag} */,
  {32'h3fece129, 32'h3e346570} /* (8, 26, 19) {real, imag} */,
  {32'h3f939c85, 32'h3d33ce51} /* (8, 26, 18) {real, imag} */,
  {32'h3f45e901, 32'h3fe6adc9} /* (8, 26, 17) {real, imag} */,
  {32'hbe390bc5, 32'h3eb1752a} /* (8, 26, 16) {real, imag} */,
  {32'h3f60e330, 32'hbecd52c1} /* (8, 26, 15) {real, imag} */,
  {32'hc021c5c7, 32'h3fc00ce7} /* (8, 26, 14) {real, imag} */,
  {32'h4083f2bd, 32'hc04581ef} /* (8, 26, 13) {real, imag} */,
  {32'hbf047bc4, 32'h40015670} /* (8, 26, 12) {real, imag} */,
  {32'h3f46178b, 32'h3f7ad896} /* (8, 26, 11) {real, imag} */,
  {32'hbf5cf2d6, 32'h40245e9d} /* (8, 26, 10) {real, imag} */,
  {32'hbfcec06a, 32'h3f93432f} /* (8, 26, 9) {real, imag} */,
  {32'hc02b0991, 32'h3fe19dda} /* (8, 26, 8) {real, imag} */,
  {32'hbf5d393c, 32'hc04a1e7d} /* (8, 26, 7) {real, imag} */,
  {32'hc04abc21, 32'hbf6403bc} /* (8, 26, 6) {real, imag} */,
  {32'h408c3e11, 32'hbf986466} /* (8, 26, 5) {real, imag} */,
  {32'h406c1d8e, 32'hc09b4062} /* (8, 26, 4) {real, imag} */,
  {32'h4002383b, 32'h3f8a7e1d} /* (8, 26, 3) {real, imag} */,
  {32'hbcdba04a, 32'hc0a10d38} /* (8, 26, 2) {real, imag} */,
  {32'hc076475d, 32'h3faac55a} /* (8, 26, 1) {real, imag} */,
  {32'hc02525c3, 32'h3ea5dace} /* (8, 26, 0) {real, imag} */,
  {32'h3fc944ed, 32'hbda8c5b1} /* (8, 25, 31) {real, imag} */,
  {32'hbf65e14e, 32'h3f590af0} /* (8, 25, 30) {real, imag} */,
  {32'hc07ff1bb, 32'hbe9cbd5f} /* (8, 25, 29) {real, imag} */,
  {32'h3f3f6969, 32'hbf55a413} /* (8, 25, 28) {real, imag} */,
  {32'h3fe00cd7, 32'hc076fb7d} /* (8, 25, 27) {real, imag} */,
  {32'hc088387d, 32'h3ffbec55} /* (8, 25, 26) {real, imag} */,
  {32'h3f9b9b50, 32'h3e7678bd} /* (8, 25, 25) {real, imag} */,
  {32'hbf7d8090, 32'hbfe8ec30} /* (8, 25, 24) {real, imag} */,
  {32'hbfaa8660, 32'hbebda981} /* (8, 25, 23) {real, imag} */,
  {32'h403c563c, 32'h3ff1fa6b} /* (8, 25, 22) {real, imag} */,
  {32'h3f1ee1a5, 32'h3fbf5105} /* (8, 25, 21) {real, imag} */,
  {32'hbefd470c, 32'hbf7a4b57} /* (8, 25, 20) {real, imag} */,
  {32'hbf921a0e, 32'h40115ae8} /* (8, 25, 19) {real, imag} */,
  {32'h40117946, 32'h3fca6058} /* (8, 25, 18) {real, imag} */,
  {32'hbf02f168, 32'h3efbabf3} /* (8, 25, 17) {real, imag} */,
  {32'h3d667af6, 32'h3ff1743a} /* (8, 25, 16) {real, imag} */,
  {32'hbf8d970d, 32'hbf53d23b} /* (8, 25, 15) {real, imag} */,
  {32'hbf03d28f, 32'hbede2452} /* (8, 25, 14) {real, imag} */,
  {32'h3f835075, 32'h3ec7acc7} /* (8, 25, 13) {real, imag} */,
  {32'hc00f1c4c, 32'hc07550b5} /* (8, 25, 12) {real, imag} */,
  {32'hbf97e8b1, 32'h3f3152cb} /* (8, 25, 11) {real, imag} */,
  {32'hbf304d03, 32'h4055df68} /* (8, 25, 10) {real, imag} */,
  {32'h402ec423, 32'h3fa59977} /* (8, 25, 9) {real, imag} */,
  {32'h40622b4c, 32'hbfae6536} /* (8, 25, 8) {real, imag} */,
  {32'h403c31fe, 32'hc04634a8} /* (8, 25, 7) {real, imag} */,
  {32'h3f6a943f, 32'h40712c61} /* (8, 25, 6) {real, imag} */,
  {32'hbeedda40, 32'h406f5cbc} /* (8, 25, 5) {real, imag} */,
  {32'hc00eb141, 32'h403628da} /* (8, 25, 4) {real, imag} */,
  {32'h401687b1, 32'h3fb48a0f} /* (8, 25, 3) {real, imag} */,
  {32'h3fecccdb, 32'hc0907925} /* (8, 25, 2) {real, imag} */,
  {32'hbfe83aac, 32'hbf593256} /* (8, 25, 1) {real, imag} */,
  {32'hbfe1bc8d, 32'h4093c6b7} /* (8, 25, 0) {real, imag} */,
  {32'h4022beb3, 32'hc0c9f02f} /* (8, 24, 31) {real, imag} */,
  {32'hbec2af62, 32'h4038e26c} /* (8, 24, 30) {real, imag} */,
  {32'hc07f9759, 32'hbfd5ea30} /* (8, 24, 29) {real, imag} */,
  {32'h3ff6a202, 32'h3f4cfafe} /* (8, 24, 28) {real, imag} */,
  {32'h3e70b571, 32'h4064645d} /* (8, 24, 27) {real, imag} */,
  {32'h3e8bc5c5, 32'h40006fe4} /* (8, 24, 26) {real, imag} */,
  {32'hc08d0146, 32'hbe9cb98a} /* (8, 24, 25) {real, imag} */,
  {32'h3ff216df, 32'hbf2693ce} /* (8, 24, 24) {real, imag} */,
  {32'hbfb29a42, 32'hc0403ea2} /* (8, 24, 23) {real, imag} */,
  {32'h3f852361, 32'h3f916a17} /* (8, 24, 22) {real, imag} */,
  {32'h3f20a758, 32'hbfd77344} /* (8, 24, 21) {real, imag} */,
  {32'h3f309b1a, 32'hbf8f63cf} /* (8, 24, 20) {real, imag} */,
  {32'h400d6860, 32'hc03ea852} /* (8, 24, 19) {real, imag} */,
  {32'h3f896f09, 32'hbff87b18} /* (8, 24, 18) {real, imag} */,
  {32'hbed00231, 32'hbfd488b5} /* (8, 24, 17) {real, imag} */,
  {32'hbd018bf5, 32'h3fc9bac7} /* (8, 24, 16) {real, imag} */,
  {32'h3f935d0c, 32'hbe554049} /* (8, 24, 15) {real, imag} */,
  {32'h3f853d01, 32'hbebbe18d} /* (8, 24, 14) {real, imag} */,
  {32'hbf897d97, 32'h3fc87b9b} /* (8, 24, 13) {real, imag} */,
  {32'h3fdf954e, 32'h3f601ba9} /* (8, 24, 12) {real, imag} */,
  {32'hbecbe5fa, 32'hbec6fbe8} /* (8, 24, 11) {real, imag} */,
  {32'hbfb82030, 32'hbf8297f7} /* (8, 24, 10) {real, imag} */,
  {32'h3f50a3d8, 32'h3cb43b3b} /* (8, 24, 9) {real, imag} */,
  {32'hc09ac38c, 32'hbdeec6fa} /* (8, 24, 8) {real, imag} */,
  {32'hc04cc6ef, 32'hbf211cda} /* (8, 24, 7) {real, imag} */,
  {32'h3ff6da26, 32'h3e454a84} /* (8, 24, 6) {real, imag} */,
  {32'hbfd50256, 32'h3fd0bb3d} /* (8, 24, 5) {real, imag} */,
  {32'h3ff2d67a, 32'h40a08055} /* (8, 24, 4) {real, imag} */,
  {32'h403d89a0, 32'hc062c656} /* (8, 24, 3) {real, imag} */,
  {32'hc0856f3e, 32'h40c2d127} /* (8, 24, 2) {real, imag} */,
  {32'h3db0e881, 32'hc0d8e539} /* (8, 24, 1) {real, imag} */,
  {32'h402dc63a, 32'hbf963580} /* (8, 24, 0) {real, imag} */,
  {32'hbf8fec25, 32'hc06e37af} /* (8, 23, 31) {real, imag} */,
  {32'hbf855394, 32'hc05b7306} /* (8, 23, 30) {real, imag} */,
  {32'h3f0b3487, 32'h40148b21} /* (8, 23, 29) {real, imag} */,
  {32'h40012b8e, 32'h3e4c1eeb} /* (8, 23, 28) {real, imag} */,
  {32'h3e4e190b, 32'hbf236e39} /* (8, 23, 27) {real, imag} */,
  {32'h3f54a110, 32'hbf23aa15} /* (8, 23, 26) {real, imag} */,
  {32'h3febd5ce, 32'hbfaac166} /* (8, 23, 25) {real, imag} */,
  {32'hbf1421fe, 32'hbf09bdf4} /* (8, 23, 24) {real, imag} */,
  {32'h3ef6a47b, 32'hc006a36e} /* (8, 23, 23) {real, imag} */,
  {32'hbf8a6c01, 32'h3fa31f54} /* (8, 23, 22) {real, imag} */,
  {32'h3ef46629, 32'h40585d9b} /* (8, 23, 21) {real, imag} */,
  {32'h3f5d0d42, 32'h401a702a} /* (8, 23, 20) {real, imag} */,
  {32'hc0bd2bc7, 32'h3fafbfb6} /* (8, 23, 19) {real, imag} */,
  {32'h40264227, 32'h3f12b357} /* (8, 23, 18) {real, imag} */,
  {32'hbe1a4712, 32'h3fae2abf} /* (8, 23, 17) {real, imag} */,
  {32'hbfc8d6dd, 32'h3e990e8f} /* (8, 23, 16) {real, imag} */,
  {32'hbea4cb1e, 32'h40698207} /* (8, 23, 15) {real, imag} */,
  {32'hc0303eb8, 32'hc0d50226} /* (8, 23, 14) {real, imag} */,
  {32'hc0167e9c, 32'h3fa08064} /* (8, 23, 13) {real, imag} */,
  {32'h402ed0b9, 32'h3ff7a508} /* (8, 23, 12) {real, imag} */,
  {32'h3f528af8, 32'h402b985a} /* (8, 23, 11) {real, imag} */,
  {32'hbed9f97e, 32'h3f961a0c} /* (8, 23, 10) {real, imag} */,
  {32'hc00f0240, 32'hbf8c0798} /* (8, 23, 9) {real, imag} */,
  {32'hbfe6b0cb, 32'hbfe258cf} /* (8, 23, 8) {real, imag} */,
  {32'h3f15a46d, 32'h401faf55} /* (8, 23, 7) {real, imag} */,
  {32'hbf61fc77, 32'hbf65b504} /* (8, 23, 6) {real, imag} */,
  {32'hc009bc3f, 32'hc008f0be} /* (8, 23, 5) {real, imag} */,
  {32'h3e88bc2b, 32'h400dd446} /* (8, 23, 4) {real, imag} */,
  {32'hbf8fb1a9, 32'h40034005} /* (8, 23, 3) {real, imag} */,
  {32'h3f8c9b05, 32'h408583e8} /* (8, 23, 2) {real, imag} */,
  {32'h3cde947c, 32'hbfc5d969} /* (8, 23, 1) {real, imag} */,
  {32'hbe84d13e, 32'h40845dcb} /* (8, 23, 0) {real, imag} */,
  {32'hbf970ef7, 32'hbf5adeac} /* (8, 22, 31) {real, imag} */,
  {32'h3ffd5a5f, 32'h3e4c7b92} /* (8, 22, 30) {real, imag} */,
  {32'h3fd1e116, 32'h3e9eb1df} /* (8, 22, 29) {real, imag} */,
  {32'h405c4543, 32'h3f3f6e94} /* (8, 22, 28) {real, imag} */,
  {32'hbe52f120, 32'h40aca82a} /* (8, 22, 27) {real, imag} */,
  {32'hbf86a598, 32'hbf696ae2} /* (8, 22, 26) {real, imag} */,
  {32'hbf8edb33, 32'hbfe3598c} /* (8, 22, 25) {real, imag} */,
  {32'hbf96b30c, 32'hbeddb02c} /* (8, 22, 24) {real, imag} */,
  {32'h3f9362a8, 32'hbf54be83} /* (8, 22, 23) {real, imag} */,
  {32'h3fb82880, 32'h3ff49547} /* (8, 22, 22) {real, imag} */,
  {32'hbd222105, 32'hbf2fe9d7} /* (8, 22, 21) {real, imag} */,
  {32'h3fd4ee42, 32'h404889c5} /* (8, 22, 20) {real, imag} */,
  {32'h3f5a3b46, 32'h3f81bacf} /* (8, 22, 19) {real, imag} */,
  {32'hc002e8c3, 32'h3ea7725d} /* (8, 22, 18) {real, imag} */,
  {32'h3f82dd5c, 32'hc032626f} /* (8, 22, 17) {real, imag} */,
  {32'hbfd5e880, 32'hc0244b7b} /* (8, 22, 16) {real, imag} */,
  {32'h3e0f8fa6, 32'hbfde75e3} /* (8, 22, 15) {real, imag} */,
  {32'hbf7faed8, 32'hbf29a535} /* (8, 22, 14) {real, imag} */,
  {32'hbe75eed1, 32'h3e16a5f6} /* (8, 22, 13) {real, imag} */,
  {32'h4035c8e2, 32'h3db4806d} /* (8, 22, 12) {real, imag} */,
  {32'h400fb16e, 32'hbd60911a} /* (8, 22, 11) {real, imag} */,
  {32'hc02f8c10, 32'hc074f6af} /* (8, 22, 10) {real, imag} */,
  {32'h3fb0aac4, 32'h3fd1ecf9} /* (8, 22, 9) {real, imag} */,
  {32'h40064767, 32'h3e4dea37} /* (8, 22, 8) {real, imag} */,
  {32'hbff32d59, 32'h3f93188e} /* (8, 22, 7) {real, imag} */,
  {32'hc007f512, 32'hbf6f47fb} /* (8, 22, 6) {real, imag} */,
  {32'hbf955c89, 32'hc08ee877} /* (8, 22, 5) {real, imag} */,
  {32'h4027b998, 32'h40146060} /* (8, 22, 4) {real, imag} */,
  {32'hc01dd2ec, 32'hbf81ed4a} /* (8, 22, 3) {real, imag} */,
  {32'hbfdaa122, 32'hc08898f0} /* (8, 22, 2) {real, imag} */,
  {32'h409af695, 32'h3f9e5eec} /* (8, 22, 1) {real, imag} */,
  {32'hc00b6118, 32'h40501a1b} /* (8, 22, 0) {real, imag} */,
  {32'hbfd6e4cb, 32'hbfbc76c3} /* (8, 21, 31) {real, imag} */,
  {32'h3fcd0a29, 32'h3f866868} /* (8, 21, 30) {real, imag} */,
  {32'h401f9023, 32'h3e1b9154} /* (8, 21, 29) {real, imag} */,
  {32'hc07c68f4, 32'h40917a49} /* (8, 21, 28) {real, imag} */,
  {32'hbfb6c5e9, 32'hbf99a7bb} /* (8, 21, 27) {real, imag} */,
  {32'hbeb0587a, 32'h3f0071c6} /* (8, 21, 26) {real, imag} */,
  {32'h3fc32768, 32'hbfe59f91} /* (8, 21, 25) {real, imag} */,
  {32'hbe2bee7b, 32'hbf60bcda} /* (8, 21, 24) {real, imag} */,
  {32'h3dd42154, 32'h3f772725} /* (8, 21, 23) {real, imag} */,
  {32'hbf841672, 32'hc007947a} /* (8, 21, 22) {real, imag} */,
  {32'h3fde813e, 32'h3e1c825b} /* (8, 21, 21) {real, imag} */,
  {32'hc05c4bcc, 32'h3fcc9d13} /* (8, 21, 20) {real, imag} */,
  {32'h3f3c6f9f, 32'h3ea7ae1b} /* (8, 21, 19) {real, imag} */,
  {32'h3e766cd6, 32'h3c052ff8} /* (8, 21, 18) {real, imag} */,
  {32'h3f5b5e5f, 32'h3f5d0ea7} /* (8, 21, 17) {real, imag} */,
  {32'h3fca3ce5, 32'hbe40fc02} /* (8, 21, 16) {real, imag} */,
  {32'hbeab4d8d, 32'h3eb52eec} /* (8, 21, 15) {real, imag} */,
  {32'h3e9dc48c, 32'h3e503df9} /* (8, 21, 14) {real, imag} */,
  {32'hbf8758de, 32'hbff9920a} /* (8, 21, 13) {real, imag} */,
  {32'hbf9eed0e, 32'h3df7da54} /* (8, 21, 12) {real, imag} */,
  {32'h4015f1fd, 32'h4094cdb4} /* (8, 21, 11) {real, imag} */,
  {32'h3f8c5bed, 32'hbdacfb0e} /* (8, 21, 10) {real, imag} */,
  {32'h4015742b, 32'hbeb09856} /* (8, 21, 9) {real, imag} */,
  {32'hbfb490d2, 32'hbfb9d34e} /* (8, 21, 8) {real, imag} */,
  {32'hc00b7f64, 32'hbf2b26f5} /* (8, 21, 7) {real, imag} */,
  {32'hbe860f04, 32'h403728ef} /* (8, 21, 6) {real, imag} */,
  {32'h3f4c258f, 32'hbd2984e0} /* (8, 21, 5) {real, imag} */,
  {32'h3d8ba7d5, 32'hc0115e6f} /* (8, 21, 4) {real, imag} */,
  {32'hbf932217, 32'hbe902fea} /* (8, 21, 3) {real, imag} */,
  {32'h3e106350, 32'h3fafc8a9} /* (8, 21, 2) {real, imag} */,
  {32'h3fc1c473, 32'hc0050130} /* (8, 21, 1) {real, imag} */,
  {32'hbefd7ec7, 32'hbe0ac460} /* (8, 21, 0) {real, imag} */,
  {32'h3ff92039, 32'hbfb7902f} /* (8, 20, 31) {real, imag} */,
  {32'h3f8d1b81, 32'hc000edd7} /* (8, 20, 30) {real, imag} */,
  {32'hbebb454e, 32'h3fce4a4f} /* (8, 20, 29) {real, imag} */,
  {32'hbfd5aee4, 32'hbfbcd579} /* (8, 20, 28) {real, imag} */,
  {32'hbfc0aab0, 32'h3f7d943f} /* (8, 20, 27) {real, imag} */,
  {32'h3fa2c609, 32'hbf2e1460} /* (8, 20, 26) {real, imag} */,
  {32'hbeebc58a, 32'h405f9c22} /* (8, 20, 25) {real, imag} */,
  {32'h3f77a21f, 32'hbf5b80e4} /* (8, 20, 24) {real, imag} */,
  {32'h3f8702c4, 32'hbf977b6e} /* (8, 20, 23) {real, imag} */,
  {32'h40827bd9, 32'h4003ae30} /* (8, 20, 22) {real, imag} */,
  {32'hbed32ae7, 32'h3fc6f9a0} /* (8, 20, 21) {real, imag} */,
  {32'hbf3234c1, 32'h3f8772e6} /* (8, 20, 20) {real, imag} */,
  {32'h3fd17f4c, 32'hbfa063a1} /* (8, 20, 19) {real, imag} */,
  {32'h4056f8da, 32'hbf1ad316} /* (8, 20, 18) {real, imag} */,
  {32'hbfbb4735, 32'h3fe15654} /* (8, 20, 17) {real, imag} */,
  {32'hc004c911, 32'h3f86495a} /* (8, 20, 16) {real, imag} */,
  {32'h3dcb4322, 32'h4021d0a0} /* (8, 20, 15) {real, imag} */,
  {32'h3f222865, 32'hc02e2794} /* (8, 20, 14) {real, imag} */,
  {32'h3f0e1eb9, 32'hbfda5d67} /* (8, 20, 13) {real, imag} */,
  {32'h3f89b713, 32'hbe5ddbe9} /* (8, 20, 12) {real, imag} */,
  {32'hbffd7ebe, 32'hc01810e2} /* (8, 20, 11) {real, imag} */,
  {32'hbf58bffe, 32'hbf374fbb} /* (8, 20, 10) {real, imag} */,
  {32'hbd50bb57, 32'hc003373d} /* (8, 20, 9) {real, imag} */,
  {32'h3f93fc41, 32'hc067f84d} /* (8, 20, 8) {real, imag} */,
  {32'h3f739fdd, 32'hbf9f7a04} /* (8, 20, 7) {real, imag} */,
  {32'hbf99724c, 32'h403071b7} /* (8, 20, 6) {real, imag} */,
  {32'hbfbd3e19, 32'hbffa5eaa} /* (8, 20, 5) {real, imag} */,
  {32'hbfac1d89, 32'hc02c4c16} /* (8, 20, 4) {real, imag} */,
  {32'hbfb52bce, 32'h401b8ac4} /* (8, 20, 3) {real, imag} */,
  {32'hbfad98d1, 32'h3f2866dc} /* (8, 20, 2) {real, imag} */,
  {32'h3d33cf7c, 32'hbe419997} /* (8, 20, 1) {real, imag} */,
  {32'hbf95c6ad, 32'hc02d3695} /* (8, 20, 0) {real, imag} */,
  {32'hbfba2814, 32'h40435130} /* (8, 19, 31) {real, imag} */,
  {32'h3fa609fe, 32'h3c64e742} /* (8, 19, 30) {real, imag} */,
  {32'h3f4cb597, 32'hbfb9b6fd} /* (8, 19, 29) {real, imag} */,
  {32'h40050c77, 32'h3f70cb85} /* (8, 19, 28) {real, imag} */,
  {32'hbeb0e229, 32'h3e9b98c2} /* (8, 19, 27) {real, imag} */,
  {32'hbff1788c, 32'h3ebe577c} /* (8, 19, 26) {real, imag} */,
  {32'h3ff0d3c9, 32'h3fd6337c} /* (8, 19, 25) {real, imag} */,
  {32'h40250c4b, 32'hbf0757e6} /* (8, 19, 24) {real, imag} */,
  {32'h3ed3e0db, 32'hbf84d3da} /* (8, 19, 23) {real, imag} */,
  {32'h3e87697f, 32'h3f820af6} /* (8, 19, 22) {real, imag} */,
  {32'h4089be61, 32'h3ebdccfb} /* (8, 19, 21) {real, imag} */,
  {32'h404d6c90, 32'h406ad6d0} /* (8, 19, 20) {real, imag} */,
  {32'h3f82b0b5, 32'hc03d6369} /* (8, 19, 19) {real, imag} */,
  {32'hbf9a700d, 32'h3f778e12} /* (8, 19, 18) {real, imag} */,
  {32'hbd32a24b, 32'h3fc2716a} /* (8, 19, 17) {real, imag} */,
  {32'h3f37fa64, 32'h3f58ec4c} /* (8, 19, 16) {real, imag} */,
  {32'h3cca1103, 32'h3f408a04} /* (8, 19, 15) {real, imag} */,
  {32'hbfab34a0, 32'hbfe29321} /* (8, 19, 14) {real, imag} */,
  {32'h4080f25c, 32'h3fc59d19} /* (8, 19, 13) {real, imag} */,
  {32'hc0433a64, 32'hbeae040d} /* (8, 19, 12) {real, imag} */,
  {32'hc001f16e, 32'hbe455383} /* (8, 19, 11) {real, imag} */,
  {32'hbff6e22a, 32'h3f3696b6} /* (8, 19, 10) {real, imag} */,
  {32'hbf41fccd, 32'h3f430f7e} /* (8, 19, 9) {real, imag} */,
  {32'hbf6ed8cd, 32'hc02ada54} /* (8, 19, 8) {real, imag} */,
  {32'hbe2b1aed, 32'h3fc4a587} /* (8, 19, 7) {real, imag} */,
  {32'h3f897517, 32'hc03a39bb} /* (8, 19, 6) {real, imag} */,
  {32'h403a221c, 32'hbed2c3a1} /* (8, 19, 5) {real, imag} */,
  {32'h3eb65c48, 32'h3fde7a5f} /* (8, 19, 4) {real, imag} */,
  {32'h3ec8715b, 32'hbf6e1f72} /* (8, 19, 3) {real, imag} */,
  {32'h3fd08426, 32'hbffb5ae6} /* (8, 19, 2) {real, imag} */,
  {32'hbfa96b44, 32'hc01277f6} /* (8, 19, 1) {real, imag} */,
  {32'h3ff45703, 32'hbf2e1fe3} /* (8, 19, 0) {real, imag} */,
  {32'hbf89e306, 32'h3f187d8e} /* (8, 18, 31) {real, imag} */,
  {32'h3f5ab9e2, 32'h3fbf31e9} /* (8, 18, 30) {real, imag} */,
  {32'hbf227761, 32'h406692f3} /* (8, 18, 29) {real, imag} */,
  {32'h3e66eb59, 32'h3f901c7b} /* (8, 18, 28) {real, imag} */,
  {32'hbf20000d, 32'hbf452e64} /* (8, 18, 27) {real, imag} */,
  {32'hbfbc7eed, 32'hbe47e577} /* (8, 18, 26) {real, imag} */,
  {32'h3f9eae69, 32'h402ad165} /* (8, 18, 25) {real, imag} */,
  {32'h3fe262fa, 32'hbca09f9c} /* (8, 18, 24) {real, imag} */,
  {32'h3fd72362, 32'hc03deebd} /* (8, 18, 23) {real, imag} */,
  {32'hbfe828e3, 32'h3fa9efa3} /* (8, 18, 22) {real, imag} */,
  {32'h3f952608, 32'hc022c02a} /* (8, 18, 21) {real, imag} */,
  {32'h40211068, 32'hc0623e3f} /* (8, 18, 20) {real, imag} */,
  {32'hbe650d08, 32'hbf94f8b2} /* (8, 18, 19) {real, imag} */,
  {32'h3f0b2336, 32'hbd7afafe} /* (8, 18, 18) {real, imag} */,
  {32'h3e480091, 32'h3e2f722e} /* (8, 18, 17) {real, imag} */,
  {32'h3fe51e1c, 32'hbf868985} /* (8, 18, 16) {real, imag} */,
  {32'hbfc83d62, 32'h3f5364c2} /* (8, 18, 15) {real, imag} */,
  {32'hbefe3a91, 32'hc00e0952} /* (8, 18, 14) {real, imag} */,
  {32'hbf22f030, 32'h3f6033b6} /* (8, 18, 13) {real, imag} */,
  {32'h3fbb869f, 32'h3fb3c908} /* (8, 18, 12) {real, imag} */,
  {32'hbfa0d742, 32'hc050c68b} /* (8, 18, 11) {real, imag} */,
  {32'hbd10f733, 32'hbd7c138c} /* (8, 18, 10) {real, imag} */,
  {32'h408d8f22, 32'h3f079c3a} /* (8, 18, 9) {real, imag} */,
  {32'h40345720, 32'h3edaabe2} /* (8, 18, 8) {real, imag} */,
  {32'h3f47bdf4, 32'h3fd0de85} /* (8, 18, 7) {real, imag} */,
  {32'hc05124dd, 32'hbdc4d747} /* (8, 18, 6) {real, imag} */,
  {32'hbf780b09, 32'hbf5115f6} /* (8, 18, 5) {real, imag} */,
  {32'h401b619b, 32'h3f25bdbb} /* (8, 18, 4) {real, imag} */,
  {32'hbf88a7e1, 32'hbed91430} /* (8, 18, 3) {real, imag} */,
  {32'h3f08f130, 32'hbe6b9745} /* (8, 18, 2) {real, imag} */,
  {32'hbf5463b9, 32'hc018ed72} /* (8, 18, 1) {real, imag} */,
  {32'hc0103ba8, 32'hbf0a4c4a} /* (8, 18, 0) {real, imag} */,
  {32'hbf6f6293, 32'hbf312106} /* (8, 17, 31) {real, imag} */,
  {32'hbeadfdf7, 32'hbee20324} /* (8, 17, 30) {real, imag} */,
  {32'h3ed68f38, 32'hbf0635e6} /* (8, 17, 29) {real, imag} */,
  {32'h3def66cb, 32'h3e2e1468} /* (8, 17, 28) {real, imag} */,
  {32'h3ec88569, 32'h402c9471} /* (8, 17, 27) {real, imag} */,
  {32'hbfacadb5, 32'h404d72dd} /* (8, 17, 26) {real, imag} */,
  {32'hbeae338f, 32'hbf8332cd} /* (8, 17, 25) {real, imag} */,
  {32'h3e9c70f9, 32'h40445380} /* (8, 17, 24) {real, imag} */,
  {32'hbf1a2376, 32'h405b1945} /* (8, 17, 23) {real, imag} */,
  {32'h3f534955, 32'h4007747d} /* (8, 17, 22) {real, imag} */,
  {32'hbe38f35c, 32'h3f9574b5} /* (8, 17, 21) {real, imag} */,
  {32'hc02ce79d, 32'hbf2580c6} /* (8, 17, 20) {real, imag} */,
  {32'h3eb9f539, 32'hbff75057} /* (8, 17, 19) {real, imag} */,
  {32'h3f5c431d, 32'h3f600ad3} /* (8, 17, 18) {real, imag} */,
  {32'h3c8beecf, 32'hbeda28b1} /* (8, 17, 17) {real, imag} */,
  {32'hbf0175fb, 32'hbf326f2b} /* (8, 17, 16) {real, imag} */,
  {32'hbcf0d3c7, 32'hc0173e85} /* (8, 17, 15) {real, imag} */,
  {32'h3d471995, 32'h3d8ac1e0} /* (8, 17, 14) {real, imag} */,
  {32'h3faca6e5, 32'hbf30e0be} /* (8, 17, 13) {real, imag} */,
  {32'h3f647ed1, 32'hbf86fb99} /* (8, 17, 12) {real, imag} */,
  {32'hbfe7d3ac, 32'h3f917420} /* (8, 17, 11) {real, imag} */,
  {32'h3f8a7921, 32'h4023fd86} /* (8, 17, 10) {real, imag} */,
  {32'h3d8f889c, 32'hbd4991ca} /* (8, 17, 9) {real, imag} */,
  {32'hbf78c41a, 32'hc01c9a65} /* (8, 17, 8) {real, imag} */,
  {32'h3feb77e2, 32'hbedfdc00} /* (8, 17, 7) {real, imag} */,
  {32'h3f28b4a5, 32'h3f9585e3} /* (8, 17, 6) {real, imag} */,
  {32'h3ffee69b, 32'hbf5e1a92} /* (8, 17, 5) {real, imag} */,
  {32'hbf063c42, 32'h400c34ca} /* (8, 17, 4) {real, imag} */,
  {32'hc01a4a70, 32'hbf8346cc} /* (8, 17, 3) {real, imag} */,
  {32'hbf529a57, 32'hbe3f18e5} /* (8, 17, 2) {real, imag} */,
  {32'h4023c02f, 32'h3e70a683} /* (8, 17, 1) {real, imag} */,
  {32'hbe5e263f, 32'h3f16b252} /* (8, 17, 0) {real, imag} */,
  {32'hc02c2d4d, 32'hbefcfc6c} /* (8, 16, 31) {real, imag} */,
  {32'hbf90574e, 32'hbf432cb1} /* (8, 16, 30) {real, imag} */,
  {32'hbfd57071, 32'h3f6a4c3a} /* (8, 16, 29) {real, imag} */,
  {32'hbfc80ee1, 32'h3dd2eb79} /* (8, 16, 28) {real, imag} */,
  {32'hbfa8712e, 32'hbfce6892} /* (8, 16, 27) {real, imag} */,
  {32'h3feab74a, 32'hbe1741be} /* (8, 16, 26) {real, imag} */,
  {32'h3f907e5b, 32'h4001ef69} /* (8, 16, 25) {real, imag} */,
  {32'hbf481f85, 32'hbfc3862b} /* (8, 16, 24) {real, imag} */,
  {32'hbeed07e9, 32'h3f521e43} /* (8, 16, 23) {real, imag} */,
  {32'hbf1eb2c9, 32'h3e687bd3} /* (8, 16, 22) {real, imag} */,
  {32'hbf49d3e4, 32'h3fe4bfa1} /* (8, 16, 21) {real, imag} */,
  {32'h3ef5c081, 32'hbfee26d6} /* (8, 16, 20) {real, imag} */,
  {32'hbe11f38b, 32'h3f92f9ef} /* (8, 16, 19) {real, imag} */,
  {32'hc0570d8f, 32'h3f1731d6} /* (8, 16, 18) {real, imag} */,
  {32'h3f8ccddb, 32'h3e81a58a} /* (8, 16, 17) {real, imag} */,
  {32'h3fef6f04, 32'h3f1e8ccb} /* (8, 16, 16) {real, imag} */,
  {32'hbd7e0484, 32'hbf0fb677} /* (8, 16, 15) {real, imag} */,
  {32'hbe97d747, 32'hbee90fd4} /* (8, 16, 14) {real, imag} */,
  {32'h3f6d9bb8, 32'h3f3a79cc} /* (8, 16, 13) {real, imag} */,
  {32'h3e8581ee, 32'h3f8b4698} /* (8, 16, 12) {real, imag} */,
  {32'hbf325ef7, 32'hbe5dcca1} /* (8, 16, 11) {real, imag} */,
  {32'hc00b9683, 32'h3ea78e3b} /* (8, 16, 10) {real, imag} */,
  {32'hbde897ef, 32'hbf478540} /* (8, 16, 9) {real, imag} */,
  {32'h4024ecaf, 32'h3f73de37} /* (8, 16, 8) {real, imag} */,
  {32'h3f427337, 32'h3f0a2343} /* (8, 16, 7) {real, imag} */,
  {32'hbfd80e8f, 32'h40037466} /* (8, 16, 6) {real, imag} */,
  {32'h3ff44b76, 32'h3f2bf986} /* (8, 16, 5) {real, imag} */,
  {32'h3fb39b8a, 32'h3fe0a979} /* (8, 16, 4) {real, imag} */,
  {32'h3ffe6504, 32'h3fdaf5af} /* (8, 16, 3) {real, imag} */,
  {32'h3f590cbe, 32'hbf2da9f4} /* (8, 16, 2) {real, imag} */,
  {32'hbf135e8e, 32'h3e879e5d} /* (8, 16, 1) {real, imag} */,
  {32'hbef8eea7, 32'hc0419af0} /* (8, 16, 0) {real, imag} */,
  {32'h3d2f5f64, 32'hc007f9fe} /* (8, 15, 31) {real, imag} */,
  {32'h3f026bc5, 32'h400dae17} /* (8, 15, 30) {real, imag} */,
  {32'h3f81c89f, 32'hbd96fcbe} /* (8, 15, 29) {real, imag} */,
  {32'h3f472c16, 32'h3f8701f6} /* (8, 15, 28) {real, imag} */,
  {32'hbfaa386f, 32'hbf6ddac7} /* (8, 15, 27) {real, imag} */,
  {32'hbd889e3c, 32'h3f83c8d8} /* (8, 15, 26) {real, imag} */,
  {32'hbfb9be52, 32'hbffb5cf6} /* (8, 15, 25) {real, imag} */,
  {32'h3f0f4fbb, 32'hbf82ef82} /* (8, 15, 24) {real, imag} */,
  {32'h3e4927cc, 32'hbfee40f5} /* (8, 15, 23) {real, imag} */,
  {32'hc00ac5b9, 32'hbfbd086b} /* (8, 15, 22) {real, imag} */,
  {32'hbeb2cb8b, 32'hbf35b875} /* (8, 15, 21) {real, imag} */,
  {32'h3edcf558, 32'h3e30d9e3} /* (8, 15, 20) {real, imag} */,
  {32'hbf3b4e9d, 32'h3e33f57e} /* (8, 15, 19) {real, imag} */,
  {32'hbe9cfcac, 32'h3f186fbe} /* (8, 15, 18) {real, imag} */,
  {32'hbf8f85e9, 32'h3e901f1e} /* (8, 15, 17) {real, imag} */,
  {32'hbf60caad, 32'h3ea84d54} /* (8, 15, 16) {real, imag} */,
  {32'hbeaeb6f9, 32'h3f9b24be} /* (8, 15, 15) {real, imag} */,
  {32'hbe238a01, 32'hbf76c4a4} /* (8, 15, 14) {real, imag} */,
  {32'h3f0b315b, 32'h3f41bc62} /* (8, 15, 13) {real, imag} */,
  {32'hc025592f, 32'hc03b1793} /* (8, 15, 12) {real, imag} */,
  {32'h3e9ff539, 32'h3e9701cf} /* (8, 15, 11) {real, imag} */,
  {32'hbe976e30, 32'hbf38e918} /* (8, 15, 10) {real, imag} */,
  {32'hbf0926fd, 32'hbf2fe7a2} /* (8, 15, 9) {real, imag} */,
  {32'hbfa17cdd, 32'h3eb2660d} /* (8, 15, 8) {real, imag} */,
  {32'hbe9237ce, 32'hbe98325a} /* (8, 15, 7) {real, imag} */,
  {32'h3f88a362, 32'h3f83623b} /* (8, 15, 6) {real, imag} */,
  {32'hbfab280b, 32'h3ef96d96} /* (8, 15, 5) {real, imag} */,
  {32'hbf757321, 32'h3fe4c3ad} /* (8, 15, 4) {real, imag} */,
  {32'hbededf1d, 32'hbfec210f} /* (8, 15, 3) {real, imag} */,
  {32'h3e5b047e, 32'h3ff24546} /* (8, 15, 2) {real, imag} */,
  {32'hbe50f42d, 32'h3f10f437} /* (8, 15, 1) {real, imag} */,
  {32'h3f377a23, 32'hc01368ce} /* (8, 15, 0) {real, imag} */,
  {32'h3da699ab, 32'h3fb26a04} /* (8, 14, 31) {real, imag} */,
  {32'hbfbd2913, 32'h3f91895e} /* (8, 14, 30) {real, imag} */,
  {32'hbed1e355, 32'hc019ffbc} /* (8, 14, 29) {real, imag} */,
  {32'hbf63122f, 32'hc0672904} /* (8, 14, 28) {real, imag} */,
  {32'h4016931a, 32'hbf0704ad} /* (8, 14, 27) {real, imag} */,
  {32'hc0140df4, 32'h3fa32959} /* (8, 14, 26) {real, imag} */,
  {32'h3fa3442c, 32'h4020a9bf} /* (8, 14, 25) {real, imag} */,
  {32'h3f36e1bd, 32'h3f999b05} /* (8, 14, 24) {real, imag} */,
  {32'h4000d282, 32'h3f53c2bf} /* (8, 14, 23) {real, imag} */,
  {32'hc00d5af1, 32'hbfa439fb} /* (8, 14, 22) {real, imag} */,
  {32'h3f8c9ebc, 32'h3fe32244} /* (8, 14, 21) {real, imag} */,
  {32'hbfdef551, 32'h401984e9} /* (8, 14, 20) {real, imag} */,
  {32'hbdf6ad57, 32'hbf21d080} /* (8, 14, 19) {real, imag} */,
  {32'h3fbf7987, 32'hc0583443} /* (8, 14, 18) {real, imag} */,
  {32'hbfee118a, 32'h4010dc14} /* (8, 14, 17) {real, imag} */,
  {32'hbf896824, 32'hc01c6b14} /* (8, 14, 16) {real, imag} */,
  {32'hbf93a371, 32'hbfb73181} /* (8, 14, 15) {real, imag} */,
  {32'h3f935f9a, 32'h400a4831} /* (8, 14, 14) {real, imag} */,
  {32'h3f34121c, 32'hbebde759} /* (8, 14, 13) {real, imag} */,
  {32'h3ea73a72, 32'h3f5e9090} /* (8, 14, 12) {real, imag} */,
  {32'h3de19c10, 32'h40286923} /* (8, 14, 11) {real, imag} */,
  {32'h3f8919e9, 32'h3f88f9dc} /* (8, 14, 10) {real, imag} */,
  {32'hbf55a814, 32'hc01d97c8} /* (8, 14, 9) {real, imag} */,
  {32'hbfe0f7b6, 32'hc03103f4} /* (8, 14, 8) {real, imag} */,
  {32'h3f93c49d, 32'hbfb6d59b} /* (8, 14, 7) {real, imag} */,
  {32'hbea82c46, 32'hc026e974} /* (8, 14, 6) {real, imag} */,
  {32'hbdeca958, 32'h3f270547} /* (8, 14, 5) {real, imag} */,
  {32'h3fed9598, 32'h3f60e696} /* (8, 14, 4) {real, imag} */,
  {32'hbe6fb784, 32'h3f12b5e2} /* (8, 14, 3) {real, imag} */,
  {32'hbf01ca49, 32'hbde4bba7} /* (8, 14, 2) {real, imag} */,
  {32'h3ff19c16, 32'h3fc3bf13} /* (8, 14, 1) {real, imag} */,
  {32'h3fa0b741, 32'h3f551362} /* (8, 14, 0) {real, imag} */,
  {32'hbfcf5194, 32'h400ee17d} /* (8, 13, 31) {real, imag} */,
  {32'hbf2b1a5c, 32'hc0148d6c} /* (8, 13, 30) {real, imag} */,
  {32'h3fda295c, 32'h3fc9978b} /* (8, 13, 29) {real, imag} */,
  {32'h3fbd4122, 32'h3f900a0f} /* (8, 13, 28) {real, imag} */,
  {32'h3f957b21, 32'h3deb74c8} /* (8, 13, 27) {real, imag} */,
  {32'h3c965504, 32'h3fa771f4} /* (8, 13, 26) {real, imag} */,
  {32'hbf611c71, 32'h4013fe53} /* (8, 13, 25) {real, imag} */,
  {32'hc00e6082, 32'h3ec9f320} /* (8, 13, 24) {real, imag} */,
  {32'hc02214af, 32'h4053571b} /* (8, 13, 23) {real, imag} */,
  {32'hbf1d9da0, 32'hbff8fb68} /* (8, 13, 22) {real, imag} */,
  {32'h3f83e7cc, 32'hc0455803} /* (8, 13, 21) {real, imag} */,
  {32'h3fa59d32, 32'hbfee73a6} /* (8, 13, 20) {real, imag} */,
  {32'hbf892560, 32'h4024b617} /* (8, 13, 19) {real, imag} */,
  {32'h403a55ce, 32'hbee98418} /* (8, 13, 18) {real, imag} */,
  {32'h3feb3afb, 32'h3eb0a0bf} /* (8, 13, 17) {real, imag} */,
  {32'hc006c524, 32'h3f99e4fd} /* (8, 13, 16) {real, imag} */,
  {32'h3ee943b8, 32'hbfd9abad} /* (8, 13, 15) {real, imag} */,
  {32'h3da240d4, 32'hbfe358a1} /* (8, 13, 14) {real, imag} */,
  {32'h3e1b9b53, 32'hbe85417f} /* (8, 13, 13) {real, imag} */,
  {32'h400ca397, 32'hbdd42c51} /* (8, 13, 12) {real, imag} */,
  {32'hc086dca5, 32'hc0486a71} /* (8, 13, 11) {real, imag} */,
  {32'h3fb24392, 32'hbee0f0f5} /* (8, 13, 10) {real, imag} */,
  {32'h4038bf6f, 32'h3f230238} /* (8, 13, 9) {real, imag} */,
  {32'h40466d06, 32'hbf693eb9} /* (8, 13, 8) {real, imag} */,
  {32'h3eec2a32, 32'hbf7f0f4e} /* (8, 13, 7) {real, imag} */,
  {32'h3f8574d5, 32'h3ffb8d32} /* (8, 13, 6) {real, imag} */,
  {32'h3f2b4e12, 32'h4021e3ff} /* (8, 13, 5) {real, imag} */,
  {32'hbe91bfb9, 32'hc0380493} /* (8, 13, 4) {real, imag} */,
  {32'hbfb44685, 32'h3f4864f6} /* (8, 13, 3) {real, imag} */,
  {32'h3dd688f5, 32'hbfb71920} /* (8, 13, 2) {real, imag} */,
  {32'hbf598cc5, 32'h3ff77817} /* (8, 13, 1) {real, imag} */,
  {32'h3db2e204, 32'hc01a6733} /* (8, 13, 0) {real, imag} */,
  {32'hbf32d11e, 32'h4009c357} /* (8, 12, 31) {real, imag} */,
  {32'hbaa96760, 32'hc02948ee} /* (8, 12, 30) {real, imag} */,
  {32'hc02a5087, 32'h3fb7fc9f} /* (8, 12, 29) {real, imag} */,
  {32'hbe2f4b26, 32'hc071953a} /* (8, 12, 28) {real, imag} */,
  {32'h3ed305a9, 32'hbff9858d} /* (8, 12, 27) {real, imag} */,
  {32'hbffc0c83, 32'h3fb89fb5} /* (8, 12, 26) {real, imag} */,
  {32'hbcc77cc1, 32'hbf5652d2} /* (8, 12, 25) {real, imag} */,
  {32'h40264257, 32'hbf617911} /* (8, 12, 24) {real, imag} */,
  {32'hbfae74c2, 32'hbf11b9bd} /* (8, 12, 23) {real, imag} */,
  {32'h3fb75646, 32'hc015f6c3} /* (8, 12, 22) {real, imag} */,
  {32'hbff84502, 32'hc03bcfa5} /* (8, 12, 21) {real, imag} */,
  {32'hbf10a5fd, 32'hbfbd4745} /* (8, 12, 20) {real, imag} */,
  {32'h4033c770, 32'hbf1ebb7c} /* (8, 12, 19) {real, imag} */,
  {32'hc040078a, 32'hbfdb666e} /* (8, 12, 18) {real, imag} */,
  {32'h3fca8a87, 32'h3f16cbd8} /* (8, 12, 17) {real, imag} */,
  {32'h3fb0a15f, 32'h3fe711ae} /* (8, 12, 16) {real, imag} */,
  {32'h3dc82db8, 32'hc0a2e797} /* (8, 12, 15) {real, imag} */,
  {32'hbfd4c1f0, 32'hbed90c38} /* (8, 12, 14) {real, imag} */,
  {32'hbf933751, 32'hc00c1ce2} /* (8, 12, 13) {real, imag} */,
  {32'h3f258ca5, 32'h3e09da80} /* (8, 12, 12) {real, imag} */,
  {32'hbea596c7, 32'h3fd2e50b} /* (8, 12, 11) {real, imag} */,
  {32'hc0560cc0, 32'h3e1c9cc4} /* (8, 12, 10) {real, imag} */,
  {32'h3f2cb7b4, 32'hbf7a85ea} /* (8, 12, 9) {real, imag} */,
  {32'h3eec266d, 32'h40a44370} /* (8, 12, 8) {real, imag} */,
  {32'h4043421f, 32'h40651ca0} /* (8, 12, 7) {real, imag} */,
  {32'h3eec1e8d, 32'hbfa1b2f6} /* (8, 12, 6) {real, imag} */,
  {32'h3fd9e973, 32'hc01a2e21} /* (8, 12, 5) {real, imag} */,
  {32'hbf8a61ca, 32'h3fd2c996} /* (8, 12, 4) {real, imag} */,
  {32'h3d1b83ec, 32'hbfe1db5f} /* (8, 12, 3) {real, imag} */,
  {32'hbf2f7179, 32'hbe8cb1bb} /* (8, 12, 2) {real, imag} */,
  {32'hbf8279a2, 32'hbeaf209f} /* (8, 12, 1) {real, imag} */,
  {32'hbe8838ef, 32'h3f9c0eb9} /* (8, 12, 0) {real, imag} */,
  {32'h4080be94, 32'h3fea3cdb} /* (8, 11, 31) {real, imag} */,
  {32'h3f62f4be, 32'h3f3da8cd} /* (8, 11, 30) {real, imag} */,
  {32'h3c9724ff, 32'h3f784581} /* (8, 11, 29) {real, imag} */,
  {32'h3f4fb4c9, 32'hc04daed6} /* (8, 11, 28) {real, imag} */,
  {32'hbf4f0823, 32'hc042a404} /* (8, 11, 27) {real, imag} */,
  {32'h40037cce, 32'h3f624ae9} /* (8, 11, 26) {real, imag} */,
  {32'hbfcf4e0f, 32'hbfb12de0} /* (8, 11, 25) {real, imag} */,
  {32'h3e3dc0c0, 32'h4000d850} /* (8, 11, 24) {real, imag} */,
  {32'hbec8b6fc, 32'hbfb18ca4} /* (8, 11, 23) {real, imag} */,
  {32'h3fe7b713, 32'h3f88c911} /* (8, 11, 22) {real, imag} */,
  {32'hbea0a4c1, 32'h3fc08e29} /* (8, 11, 21) {real, imag} */,
  {32'h3ee16d17, 32'h4016954b} /* (8, 11, 20) {real, imag} */,
  {32'h3f8000ee, 32'hbf5c03b0} /* (8, 11, 19) {real, imag} */,
  {32'hbf327cd9, 32'h3f6783a1} /* (8, 11, 18) {real, imag} */,
  {32'hbfdc94a0, 32'h3e8e9272} /* (8, 11, 17) {real, imag} */,
  {32'h3ee55716, 32'h3f1f29c2} /* (8, 11, 16) {real, imag} */,
  {32'h3e1f8326, 32'h3fd2f1d3} /* (8, 11, 15) {real, imag} */,
  {32'h3f4ab007, 32'hc05dfcd7} /* (8, 11, 14) {real, imag} */,
  {32'hc042e537, 32'hbfdb83ad} /* (8, 11, 13) {real, imag} */,
  {32'hc003b553, 32'hbdeabc32} /* (8, 11, 12) {real, imag} */,
  {32'hbf47cc31, 32'h403cfb26} /* (8, 11, 11) {real, imag} */,
  {32'hc075588e, 32'h402c501a} /* (8, 11, 10) {real, imag} */,
  {32'h3fe8b6ae, 32'hbfbf5b15} /* (8, 11, 9) {real, imag} */,
  {32'hc00def69, 32'hc0076489} /* (8, 11, 8) {real, imag} */,
  {32'hc035fe4b, 32'h3fc103f5} /* (8, 11, 7) {real, imag} */,
  {32'h40087ea4, 32'hbf1e08d0} /* (8, 11, 6) {real, imag} */,
  {32'hbff1328a, 32'h3f31ad7c} /* (8, 11, 5) {real, imag} */,
  {32'h3ff379f0, 32'hbfd9a15f} /* (8, 11, 4) {real, imag} */,
  {32'h3fa3b437, 32'hc017a7df} /* (8, 11, 3) {real, imag} */,
  {32'hc00b5e67, 32'hc058a06a} /* (8, 11, 2) {real, imag} */,
  {32'h3f5cb411, 32'h3f83c0ce} /* (8, 11, 1) {real, imag} */,
  {32'h3fd70bc2, 32'h4042add0} /* (8, 11, 0) {real, imag} */,
  {32'hc03c600d, 32'hc060dbfe} /* (8, 10, 31) {real, imag} */,
  {32'h3e8d880e, 32'h40009b07} /* (8, 10, 30) {real, imag} */,
  {32'h3eb63b1c, 32'h3e976334} /* (8, 10, 29) {real, imag} */,
  {32'hbf9a1a75, 32'h3fa06d93} /* (8, 10, 28) {real, imag} */,
  {32'h3e6fa912, 32'hbfbe09a6} /* (8, 10, 27) {real, imag} */,
  {32'hbe7e8173, 32'h3d845900} /* (8, 10, 26) {real, imag} */,
  {32'hbd43f480, 32'hbe6ddeac} /* (8, 10, 25) {real, imag} */,
  {32'h3f81e806, 32'hbecb87f8} /* (8, 10, 24) {real, imag} */,
  {32'hc00eb0d6, 32'hbfa1e476} /* (8, 10, 23) {real, imag} */,
  {32'h3eb1e8a1, 32'hbefa7d30} /* (8, 10, 22) {real, imag} */,
  {32'h3feb0f79, 32'hbeb83c2c} /* (8, 10, 21) {real, imag} */,
  {32'hbf11c69f, 32'h3edc50a1} /* (8, 10, 20) {real, imag} */,
  {32'h40112eec, 32'h40080bdf} /* (8, 10, 19) {real, imag} */,
  {32'h3e18f5e8, 32'hbf621759} /* (8, 10, 18) {real, imag} */,
  {32'h3f5c84ac, 32'hbf8c31b5} /* (8, 10, 17) {real, imag} */,
  {32'hbe88c5f6, 32'hbeb8f584} /* (8, 10, 16) {real, imag} */,
  {32'h3fdb4698, 32'hbf83f81b} /* (8, 10, 15) {real, imag} */,
  {32'hbfee1522, 32'h3eb07a62} /* (8, 10, 14) {real, imag} */,
  {32'h3e18f290, 32'h4030f6c3} /* (8, 10, 13) {real, imag} */,
  {32'hbfcb4f09, 32'h3e2b2019} /* (8, 10, 12) {real, imag} */,
  {32'h3f9d53f7, 32'hbe5eecc6} /* (8, 10, 11) {real, imag} */,
  {32'h40471e73, 32'hbfbe68c4} /* (8, 10, 10) {real, imag} */,
  {32'h3fb82a01, 32'h3e6d2a88} /* (8, 10, 9) {real, imag} */,
  {32'hbff504e1, 32'h3f4c9af9} /* (8, 10, 8) {real, imag} */,
  {32'hbd6ec555, 32'hc001ad57} /* (8, 10, 7) {real, imag} */,
  {32'hbfd478cf, 32'hc00a4e20} /* (8, 10, 6) {real, imag} */,
  {32'h3f3c6ea9, 32'h3e665376} /* (8, 10, 5) {real, imag} */,
  {32'hbebd856d, 32'hbe516c04} /* (8, 10, 4) {real, imag} */,
  {32'hc02ddce5, 32'hbf0452bc} /* (8, 10, 3) {real, imag} */,
  {32'h40569bd2, 32'hbc8b304b} /* (8, 10, 2) {real, imag} */,
  {32'hbf7ea675, 32'h3fe17ac8} /* (8, 10, 1) {real, imag} */,
  {32'hbfff24c2, 32'h3da9eb87} /* (8, 10, 0) {real, imag} */,
  {32'hc0241804, 32'hc00c1be6} /* (8, 9, 31) {real, imag} */,
  {32'hbee6c34a, 32'hc05dfc54} /* (8, 9, 30) {real, imag} */,
  {32'h3f3c7f96, 32'hbfb0f10c} /* (8, 9, 29) {real, imag} */,
  {32'hc03a9209, 32'hbfc5c806} /* (8, 9, 28) {real, imag} */,
  {32'h3f73e45c, 32'h3fbfad9a} /* (8, 9, 27) {real, imag} */,
  {32'h3f54bdea, 32'h40274056} /* (8, 9, 26) {real, imag} */,
  {32'h3f38c7fd, 32'hbe80da89} /* (8, 9, 25) {real, imag} */,
  {32'hbec50a7f, 32'h3fd55e15} /* (8, 9, 24) {real, imag} */,
  {32'h3faf1104, 32'hc02ffeb1} /* (8, 9, 23) {real, imag} */,
  {32'h3ecbeb5f, 32'h3f00c43a} /* (8, 9, 22) {real, imag} */,
  {32'hbfd96a34, 32'hbf7906a8} /* (8, 9, 21) {real, imag} */,
  {32'h3f805f73, 32'h3f221fa6} /* (8, 9, 20) {real, imag} */,
  {32'h402d009f, 32'h4089d166} /* (8, 9, 19) {real, imag} */,
  {32'hc01325e6, 32'hbe1101b1} /* (8, 9, 18) {real, imag} */,
  {32'h40203f65, 32'h3ed30c46} /* (8, 9, 17) {real, imag} */,
  {32'hbee85efe, 32'hbf96275f} /* (8, 9, 16) {real, imag} */,
  {32'h4001d217, 32'h40120f4c} /* (8, 9, 15) {real, imag} */,
  {32'h3cc57f88, 32'hbf1c45b5} /* (8, 9, 14) {real, imag} */,
  {32'h406968f3, 32'hbe80bc31} /* (8, 9, 13) {real, imag} */,
  {32'h405b83d4, 32'h4004e773} /* (8, 9, 12) {real, imag} */,
  {32'hbef074b9, 32'hbfa96358} /* (8, 9, 11) {real, imag} */,
  {32'h3f38e9f0, 32'h4007db34} /* (8, 9, 10) {real, imag} */,
  {32'hc03647c2, 32'h40035c71} /* (8, 9, 9) {real, imag} */,
  {32'h3f8d6d1c, 32'hbf902b58} /* (8, 9, 8) {real, imag} */,
  {32'hbe74859b, 32'h3e7b85e4} /* (8, 9, 7) {real, imag} */,
  {32'hbfaf2bae, 32'h3f0ec0dd} /* (8, 9, 6) {real, imag} */,
  {32'hbf4d4aa1, 32'hbf581fe6} /* (8, 9, 5) {real, imag} */,
  {32'hbfec9c74, 32'h402eb491} /* (8, 9, 4) {real, imag} */,
  {32'h4037cdea, 32'hc0770a34} /* (8, 9, 3) {real, imag} */,
  {32'hbea9044d, 32'h3ecf1229} /* (8, 9, 2) {real, imag} */,
  {32'hbfcc3d0d, 32'hbe43d6fd} /* (8, 9, 1) {real, imag} */,
  {32'hc0211aa3, 32'hbfba1744} /* (8, 9, 0) {real, imag} */,
  {32'h404b198c, 32'hbf809cb8} /* (8, 8, 31) {real, imag} */,
  {32'h3f9cdc34, 32'h3ff71051} /* (8, 8, 30) {real, imag} */,
  {32'h4004d7cd, 32'hc05c72f6} /* (8, 8, 29) {real, imag} */,
  {32'h407bfe82, 32'hc0698e16} /* (8, 8, 28) {real, imag} */,
  {32'hbf7b0e35, 32'hbf3e0ef2} /* (8, 8, 27) {real, imag} */,
  {32'hbf88056b, 32'hc021cc99} /* (8, 8, 26) {real, imag} */,
  {32'h3c33ea20, 32'hc0878c8a} /* (8, 8, 25) {real, imag} */,
  {32'hbff905b6, 32'hbfc3e516} /* (8, 8, 24) {real, imag} */,
  {32'hbf69a182, 32'hc04af914} /* (8, 8, 23) {real, imag} */,
  {32'hbeb8e6b4, 32'h4083b0d7} /* (8, 8, 22) {real, imag} */,
  {32'h40152001, 32'h401e7f87} /* (8, 8, 21) {real, imag} */,
  {32'hbf91281c, 32'h3f36759f} /* (8, 8, 20) {real, imag} */,
  {32'hbf0f65b7, 32'hbf93cf7d} /* (8, 8, 19) {real, imag} */,
  {32'h3f6898c1, 32'h3e7ef864} /* (8, 8, 18) {real, imag} */,
  {32'hbf74f8b0, 32'h3df19db2} /* (8, 8, 17) {real, imag} */,
  {32'h3fc1f54f, 32'hc0591702} /* (8, 8, 16) {real, imag} */,
  {32'h4007035b, 32'hbe56f76f} /* (8, 8, 15) {real, imag} */,
  {32'hc054f896, 32'h409bdf91} /* (8, 8, 14) {real, imag} */,
  {32'hbfb09404, 32'hbef93d4f} /* (8, 8, 13) {real, imag} */,
  {32'h3edc8de6, 32'h3e98d82a} /* (8, 8, 12) {real, imag} */,
  {32'hc0851310, 32'hbe5401e1} /* (8, 8, 11) {real, imag} */,
  {32'h404c6632, 32'h40488414} /* (8, 8, 10) {real, imag} */,
  {32'h4096c2de, 32'hc0413db1} /* (8, 8, 9) {real, imag} */,
  {32'hbf95d52e, 32'hc03cb7f7} /* (8, 8, 8) {real, imag} */,
  {32'hc019521d, 32'h3f1dbd44} /* (8, 8, 7) {real, imag} */,
  {32'h3ff5f6dc, 32'hbfd1af33} /* (8, 8, 6) {real, imag} */,
  {32'h3fb7b7e7, 32'hbfbf33a7} /* (8, 8, 5) {real, imag} */,
  {32'h40470fbc, 32'hc0c8ecb4} /* (8, 8, 4) {real, imag} */,
  {32'hbe938e34, 32'hbfd86c34} /* (8, 8, 3) {real, imag} */,
  {32'hc104f28e, 32'h3e99b8d7} /* (8, 8, 2) {real, imag} */,
  {32'h3f85c819, 32'h3fb5249b} /* (8, 8, 1) {real, imag} */,
  {32'h40188965, 32'h3f138815} /* (8, 8, 0) {real, imag} */,
  {32'hc088c08e, 32'hbfe29bb3} /* (8, 7, 31) {real, imag} */,
  {32'hbe7c8d28, 32'hbf535da0} /* (8, 7, 30) {real, imag} */,
  {32'hc0353e6f, 32'hbf1ec191} /* (8, 7, 29) {real, imag} */,
  {32'h3f7a5c7d, 32'h3f06a091} /* (8, 7, 28) {real, imag} */,
  {32'hbfbd0f5e, 32'hbe3798d6} /* (8, 7, 27) {real, imag} */,
  {32'h3fa70676, 32'hc008755e} /* (8, 7, 26) {real, imag} */,
  {32'h3d846d97, 32'h403ee135} /* (8, 7, 25) {real, imag} */,
  {32'hbf8cfd78, 32'hbf6059fb} /* (8, 7, 24) {real, imag} */,
  {32'hbefe283b, 32'hbea5941b} /* (8, 7, 23) {real, imag} */,
  {32'h403438ba, 32'hbf4103ac} /* (8, 7, 22) {real, imag} */,
  {32'hc02e0cc5, 32'h400e3eab} /* (8, 7, 21) {real, imag} */,
  {32'h3f230410, 32'hbd8a31d7} /* (8, 7, 20) {real, imag} */,
  {32'h3e767820, 32'h3c1075ba} /* (8, 7, 19) {real, imag} */,
  {32'h3e3bb36c, 32'hc011e208} /* (8, 7, 18) {real, imag} */,
  {32'h3f5c9f8a, 32'h3fe8ea08} /* (8, 7, 17) {real, imag} */,
  {32'h3ef3e08c, 32'h3ee22356} /* (8, 7, 16) {real, imag} */,
  {32'hbe7c1b7a, 32'hbf0a7546} /* (8, 7, 15) {real, imag} */,
  {32'h4026762f, 32'h3fd0a03e} /* (8, 7, 14) {real, imag} */,
  {32'hc028cf20, 32'hbfc2ca47} /* (8, 7, 13) {real, imag} */,
  {32'hbef44718, 32'h3f0d3e21} /* (8, 7, 12) {real, imag} */,
  {32'h406a044b, 32'hbf0ab662} /* (8, 7, 11) {real, imag} */,
  {32'h3e24b456, 32'h3ede9741} /* (8, 7, 10) {real, imag} */,
  {32'h3f94e675, 32'hbfece42f} /* (8, 7, 9) {real, imag} */,
  {32'h3ee9c432, 32'h4098dc93} /* (8, 7, 8) {real, imag} */,
  {32'hbfe24565, 32'h40002fdb} /* (8, 7, 7) {real, imag} */,
  {32'hc012f825, 32'h3f1a6dd4} /* (8, 7, 6) {real, imag} */,
  {32'h40305f2a, 32'h401bd4bc} /* (8, 7, 5) {real, imag} */,
  {32'hbf7e4d55, 32'h40175b97} /* (8, 7, 4) {real, imag} */,
  {32'hc06b862a, 32'h40494699} /* (8, 7, 3) {real, imag} */,
  {32'h3c9da54a, 32'hbe5f8a8e} /* (8, 7, 2) {real, imag} */,
  {32'h3fd9924a, 32'hc0c3f90b} /* (8, 7, 1) {real, imag} */,
  {32'h3fe73424, 32'h4056de71} /* (8, 7, 0) {real, imag} */,
  {32'h409baee7, 32'hbfb92203} /* (8, 6, 31) {real, imag} */,
  {32'h4046c2f7, 32'h401fb7c4} /* (8, 6, 30) {real, imag} */,
  {32'h406bef34, 32'hc0560aee} /* (8, 6, 29) {real, imag} */,
  {32'hc00fcf0a, 32'h3feb0660} /* (8, 6, 28) {real, imag} */,
  {32'hc00a90d8, 32'h400602fb} /* (8, 6, 27) {real, imag} */,
  {32'hbf9dc94b, 32'hc0418e2f} /* (8, 6, 26) {real, imag} */,
  {32'h407da905, 32'h3fb59158} /* (8, 6, 25) {real, imag} */,
  {32'h3ef4b6bf, 32'hbfa79f68} /* (8, 6, 24) {real, imag} */,
  {32'h3f7e48e3, 32'h3f8fa671} /* (8, 6, 23) {real, imag} */,
  {32'h3f85f1fd, 32'h3f8f79a5} /* (8, 6, 22) {real, imag} */,
  {32'hbf3a63c9, 32'hbe3e7e0d} /* (8, 6, 21) {real, imag} */,
  {32'h3ecc39ae, 32'hc01f4638} /* (8, 6, 20) {real, imag} */,
  {32'hbf8b275e, 32'hbf848dc0} /* (8, 6, 19) {real, imag} */,
  {32'h3ea1071b, 32'hc01320f9} /* (8, 6, 18) {real, imag} */,
  {32'h40838c00, 32'h3fcd5331} /* (8, 6, 17) {real, imag} */,
  {32'hbf8bf209, 32'hbf600c2c} /* (8, 6, 16) {real, imag} */,
  {32'h3f1ceaa0, 32'hbe59d933} /* (8, 6, 15) {real, imag} */,
  {32'h3e8a8adf, 32'h3e207cc2} /* (8, 6, 14) {real, imag} */,
  {32'hbf39bef4, 32'hbfe26b52} /* (8, 6, 13) {real, imag} */,
  {32'h400c38e3, 32'hbfc23ddb} /* (8, 6, 12) {real, imag} */,
  {32'h3eaf4fcc, 32'h3ff74801} /* (8, 6, 11) {real, imag} */,
  {32'hbfda4d8a, 32'h3f2091ad} /* (8, 6, 10) {real, imag} */,
  {32'h3eb924fc, 32'hc090728a} /* (8, 6, 9) {real, imag} */,
  {32'hc01e96ba, 32'hc080184e} /* (8, 6, 8) {real, imag} */,
  {32'hc028b9c0, 32'h3fec431f} /* (8, 6, 7) {real, imag} */,
  {32'hc0031099, 32'hbf636265} /* (8, 6, 6) {real, imag} */,
  {32'h3fd066b7, 32'hbfbec40c} /* (8, 6, 5) {real, imag} */,
  {32'h3e030747, 32'hbf06cc79} /* (8, 6, 4) {real, imag} */,
  {32'hbfe48670, 32'h4051c608} /* (8, 6, 3) {real, imag} */,
  {32'h3f5a0750, 32'hbf28abfc} /* (8, 6, 2) {real, imag} */,
  {32'h4028e993, 32'h3f19d209} /* (8, 6, 1) {real, imag} */,
  {32'hbedd3871, 32'hc0342f26} /* (8, 6, 0) {real, imag} */,
  {32'h4089e028, 32'hc0d60d12} /* (8, 5, 31) {real, imag} */,
  {32'hc05de3e6, 32'h401d8cb4} /* (8, 5, 30) {real, imag} */,
  {32'h3f611447, 32'hbf083ae3} /* (8, 5, 29) {real, imag} */,
  {32'h4060b3c4, 32'h3e5f37c8} /* (8, 5, 28) {real, imag} */,
  {32'h3fb62130, 32'h400ffbf7} /* (8, 5, 27) {real, imag} */,
  {32'h3fc40b46, 32'hbe1500c6} /* (8, 5, 26) {real, imag} */,
  {32'h3ffcb912, 32'hbfd13dd8} /* (8, 5, 25) {real, imag} */,
  {32'h3fc575cb, 32'hbf85edd3} /* (8, 5, 24) {real, imag} */,
  {32'h3f8e29e2, 32'hbda6cb58} /* (8, 5, 23) {real, imag} */,
  {32'hbe9b35c2, 32'h4055a960} /* (8, 5, 22) {real, imag} */,
  {32'hbfb0e1b9, 32'hbe9ae9c1} /* (8, 5, 21) {real, imag} */,
  {32'hbf6c2a76, 32'h3f5b8c7c} /* (8, 5, 20) {real, imag} */,
  {32'hbf780e73, 32'h3fb3a2ec} /* (8, 5, 19) {real, imag} */,
  {32'h3f6ad938, 32'h3f7afd89} /* (8, 5, 18) {real, imag} */,
  {32'hbf21cec5, 32'hbe019198} /* (8, 5, 17) {real, imag} */,
  {32'h3f0d7b46, 32'h3f670f26} /* (8, 5, 16) {real, imag} */,
  {32'h402605b5, 32'h3f87fd7b} /* (8, 5, 15) {real, imag} */,
  {32'hbf637af7, 32'hc03d72bb} /* (8, 5, 14) {real, imag} */,
  {32'hbfd570e3, 32'hc0363173} /* (8, 5, 13) {real, imag} */,
  {32'h3f8b74d5, 32'h3ecc6a14} /* (8, 5, 12) {real, imag} */,
  {32'h4064c769, 32'hc003069f} /* (8, 5, 11) {real, imag} */,
  {32'h3f199ad3, 32'hbf8689f5} /* (8, 5, 10) {real, imag} */,
  {32'hbfd8b6d2, 32'h3e0716dc} /* (8, 5, 9) {real, imag} */,
  {32'hbf99c8a3, 32'h3ed6a4c7} /* (8, 5, 8) {real, imag} */,
  {32'h3ea9ec2d, 32'h3fc13ea6} /* (8, 5, 7) {real, imag} */,
  {32'hbfe5e3a3, 32'h3c773557} /* (8, 5, 6) {real, imag} */,
  {32'h40688344, 32'h403170d8} /* (8, 5, 5) {real, imag} */,
  {32'h40180b63, 32'h4096e41a} /* (8, 5, 4) {real, imag} */,
  {32'h4003d02c, 32'hc001146e} /* (8, 5, 3) {real, imag} */,
  {32'hc0251a4d, 32'hc01855a3} /* (8, 5, 2) {real, imag} */,
  {32'h40390c61, 32'h3fbdb0b6} /* (8, 5, 1) {real, imag} */,
  {32'h40c93c1a, 32'hc03a652f} /* (8, 5, 0) {real, imag} */,
  {32'hc0599ce1, 32'hc0542d74} /* (8, 4, 31) {real, imag} */,
  {32'h40e66195, 32'hbf059971} /* (8, 4, 30) {real, imag} */,
  {32'h401048ff, 32'hbfe150fd} /* (8, 4, 29) {real, imag} */,
  {32'hbf35cf2f, 32'h3f8a6164} /* (8, 4, 28) {real, imag} */,
  {32'h3f40ff95, 32'hbdcf327b} /* (8, 4, 27) {real, imag} */,
  {32'hbfd18b62, 32'hc04100e9} /* (8, 4, 26) {real, imag} */,
  {32'h405248c1, 32'hbfaeaab9} /* (8, 4, 25) {real, imag} */,
  {32'h3ff4c602, 32'hbe58d007} /* (8, 4, 24) {real, imag} */,
  {32'hbfdf6616, 32'hbf6fcaa0} /* (8, 4, 23) {real, imag} */,
  {32'h3ecd79bc, 32'hbec7357f} /* (8, 4, 22) {real, imag} */,
  {32'h401d7724, 32'h3f4c83c5} /* (8, 4, 21) {real, imag} */,
  {32'hbf6ed86f, 32'h3dd7df8f} /* (8, 4, 20) {real, imag} */,
  {32'h3fba181c, 32'hbe398389} /* (8, 4, 19) {real, imag} */,
  {32'h40391619, 32'h3fbfa436} /* (8, 4, 18) {real, imag} */,
  {32'hbf55d955, 32'h3fde7175} /* (8, 4, 17) {real, imag} */,
  {32'h400174bc, 32'hbf405fd3} /* (8, 4, 16) {real, imag} */,
  {32'hbe126820, 32'hbf86c7a1} /* (8, 4, 15) {real, imag} */,
  {32'hbfc1ce73, 32'h3fb4da9a} /* (8, 4, 14) {real, imag} */,
  {32'hc056d4e4, 32'h40303edd} /* (8, 4, 13) {real, imag} */,
  {32'h3e646fca, 32'h40100856} /* (8, 4, 12) {real, imag} */,
  {32'hbf84e837, 32'hc01ca4f9} /* (8, 4, 11) {real, imag} */,
  {32'h3e99094b, 32'hc047c216} /* (8, 4, 10) {real, imag} */,
  {32'hc031b069, 32'h3fe7d719} /* (8, 4, 9) {real, imag} */,
  {32'h405460ce, 32'hc0a9d0f5} /* (8, 4, 8) {real, imag} */,
  {32'hc0be84d6, 32'h3f4ea635} /* (8, 4, 7) {real, imag} */,
  {32'h40055f4c, 32'hc06b31fe} /* (8, 4, 6) {real, imag} */,
  {32'h3fc9b4ff, 32'h3df3a32a} /* (8, 4, 5) {real, imag} */,
  {32'hc00dec04, 32'hc0d61f2f} /* (8, 4, 4) {real, imag} */,
  {32'h3f886eda, 32'h4000c538} /* (8, 4, 3) {real, imag} */,
  {32'h40ea6c66, 32'hc014fc6d} /* (8, 4, 2) {real, imag} */,
  {32'hc0f7e71a, 32'h405d9d64} /* (8, 4, 1) {real, imag} */,
  {32'hbf5022cf, 32'hbf2af00b} /* (8, 4, 0) {real, imag} */,
  {32'hc01df710, 32'hc0bc59ec} /* (8, 3, 31) {real, imag} */,
  {32'h40068ba2, 32'h40110168} /* (8, 3, 30) {real, imag} */,
  {32'h4095af02, 32'hbe5d8c1c} /* (8, 3, 29) {real, imag} */,
  {32'hc0887583, 32'h3fd9c269} /* (8, 3, 28) {real, imag} */,
  {32'hbf8bbac1, 32'hbf63164f} /* (8, 3, 27) {real, imag} */,
  {32'hbfba1e2b, 32'h402f3d3b} /* (8, 3, 26) {real, imag} */,
  {32'hbf9af070, 32'h3fe3bc93} /* (8, 3, 25) {real, imag} */,
  {32'hbfa6af4d, 32'hc088221b} /* (8, 3, 24) {real, imag} */,
  {32'hbe1374f0, 32'h3eadd8af} /* (8, 3, 23) {real, imag} */,
  {32'h4072adae, 32'h3f8b2986} /* (8, 3, 22) {real, imag} */,
  {32'h3fef972a, 32'h3fdf9f27} /* (8, 3, 21) {real, imag} */,
  {32'h402a8bb7, 32'hbfb9e4d5} /* (8, 3, 20) {real, imag} */,
  {32'hc042e15e, 32'hc0058722} /* (8, 3, 19) {real, imag} */,
  {32'h3dbf5c17, 32'h402f4425} /* (8, 3, 18) {real, imag} */,
  {32'hc024318f, 32'hbf1bb01f} /* (8, 3, 17) {real, imag} */,
  {32'h3f1747c6, 32'h401254a4} /* (8, 3, 16) {real, imag} */,
  {32'hbf00ce95, 32'hbffaa248} /* (8, 3, 15) {real, imag} */,
  {32'hbfb8bb56, 32'hbee15383} /* (8, 3, 14) {real, imag} */,
  {32'hbff7bfd9, 32'hbfa54964} /* (8, 3, 13) {real, imag} */,
  {32'h3fdc1dff, 32'hbfcaa280} /* (8, 3, 12) {real, imag} */,
  {32'h40020bad, 32'hbfac8376} /* (8, 3, 11) {real, imag} */,
  {32'h3ff59577, 32'hc01d2d40} /* (8, 3, 10) {real, imag} */,
  {32'hc08634e1, 32'h4079383e} /* (8, 3, 9) {real, imag} */,
  {32'h3fe109ae, 32'h4058b63d} /* (8, 3, 8) {real, imag} */,
  {32'hbebf2ac9, 32'hc06364d2} /* (8, 3, 7) {real, imag} */,
  {32'hc00da0b2, 32'h3fcfc726} /* (8, 3, 6) {real, imag} */,
  {32'h3fa69ad1, 32'h3f5b36ff} /* (8, 3, 5) {real, imag} */,
  {32'h40049929, 32'hbfcbbfed} /* (8, 3, 4) {real, imag} */,
  {32'h3fb264fd, 32'hbf0dd07a} /* (8, 3, 3) {real, imag} */,
  {32'h40b25e52, 32'h3f605d75} /* (8, 3, 2) {real, imag} */,
  {32'hc0b46bec, 32'h3f7af1c3} /* (8, 3, 1) {real, imag} */,
  {32'hc0198b69, 32'hc01042fc} /* (8, 3, 0) {real, imag} */,
  {32'h418a52a7, 32'hc13f6e8b} /* (8, 2, 31) {real, imag} */,
  {32'hc1221985, 32'h41418729} /* (8, 2, 30) {real, imag} */,
  {32'hbfc37788, 32'hc04da494} /* (8, 2, 29) {real, imag} */,
  {32'hbf9b82ce, 32'hbfa5a21c} /* (8, 2, 28) {real, imag} */,
  {32'hbf22d783, 32'hbee1a093} /* (8, 2, 27) {real, imag} */,
  {32'hbf8dbe7e, 32'h3ffead18} /* (8, 2, 26) {real, imag} */,
  {32'h3faf3379, 32'hbf8c70e9} /* (8, 2, 25) {real, imag} */,
  {32'h3c56737c, 32'h4099a259} /* (8, 2, 24) {real, imag} */,
  {32'h3f143e2d, 32'h3f8e8829} /* (8, 2, 23) {real, imag} */,
  {32'h3f9a1990, 32'hbe2bdbf7} /* (8, 2, 22) {real, imag} */,
  {32'h3df24f8b, 32'h3f127d44} /* (8, 2, 21) {real, imag} */,
  {32'h3f6fcc0b, 32'hbfbdce65} /* (8, 2, 20) {real, imag} */,
  {32'hbfb43e18, 32'hbf1bbd2e} /* (8, 2, 19) {real, imag} */,
  {32'hbee81c9d, 32'h3ea420e6} /* (8, 2, 18) {real, imag} */,
  {32'hc01d141e, 32'h3f35fcd9} /* (8, 2, 17) {real, imag} */,
  {32'hbf90ac27, 32'h3ddc047a} /* (8, 2, 16) {real, imag} */,
  {32'hbaab9847, 32'h401d3488} /* (8, 2, 15) {real, imag} */,
  {32'hc01e1211, 32'h3f8f2e45} /* (8, 2, 14) {real, imag} */,
  {32'hbe771607, 32'hbfe483ef} /* (8, 2, 13) {real, imag} */,
  {32'hbfa7470d, 32'hbe7aef39} /* (8, 2, 12) {real, imag} */,
  {32'hc07d8d66, 32'hc0608f29} /* (8, 2, 11) {real, imag} */,
  {32'hbf6c0ee3, 32'hbf49f4d7} /* (8, 2, 10) {real, imag} */,
  {32'hc01b0b8e, 32'h3eaf3b58} /* (8, 2, 9) {real, imag} */,
  {32'hc0a93501, 32'h3fa62ed5} /* (8, 2, 8) {real, imag} */,
  {32'h3f6c0b40, 32'hbec4c56e} /* (8, 2, 7) {real, imag} */,
  {32'h402fbc48, 32'h3ef82051} /* (8, 2, 6) {real, imag} */,
  {32'hc0b39358, 32'hbff2ffb4} /* (8, 2, 5) {real, imag} */,
  {32'h40b5338d, 32'hc0aec42f} /* (8, 2, 4) {real, imag} */,
  {32'h3f0c0ff0, 32'hbff0ba2f} /* (8, 2, 3) {real, imag} */,
  {32'hc02e38c4, 32'h40a92edc} /* (8, 2, 2) {real, imag} */,
  {32'h41377b40, 32'hc13ddd4c} /* (8, 2, 1) {real, imag} */,
  {32'h413aa1d1, 32'hc0edd0d4} /* (8, 2, 0) {real, imag} */,
  {32'hc147f7b4, 32'h418d40ad} /* (8, 1, 31) {real, imag} */,
  {32'hbf850bac, 32'hc0eaa787} /* (8, 1, 30) {real, imag} */,
  {32'h3e833c93, 32'h3ff07022} /* (8, 1, 29) {real, imag} */,
  {32'hc0020e1d, 32'hbfe73d4c} /* (8, 1, 28) {real, imag} */,
  {32'h4067a85b, 32'hc08d3bcd} /* (8, 1, 27) {real, imag} */,
  {32'hc003e4b5, 32'h4007aa44} /* (8, 1, 26) {real, imag} */,
  {32'hc0acfdba, 32'h3ec1145b} /* (8, 1, 25) {real, imag} */,
  {32'hbf834267, 32'hc09c8e4e} /* (8, 1, 24) {real, imag} */,
  {32'hbddf95a5, 32'h4011f28f} /* (8, 1, 23) {real, imag} */,
  {32'hc016eb8d, 32'h3f21b606} /* (8, 1, 22) {real, imag} */,
  {32'hbf9f6ecc, 32'hc0ae318e} /* (8, 1, 21) {real, imag} */,
  {32'hc022e245, 32'hc01d890c} /* (8, 1, 20) {real, imag} */,
  {32'hc041e14e, 32'h3e97b355} /* (8, 1, 19) {real, imag} */,
  {32'h3ff8cb82, 32'hbf6fe752} /* (8, 1, 18) {real, imag} */,
  {32'h3eeb19c7, 32'h3edeb623} /* (8, 1, 17) {real, imag} */,
  {32'h3e999674, 32'h3ddee17a} /* (8, 1, 16) {real, imag} */,
  {32'h3e1ceff0, 32'h3f54ef32} /* (8, 1, 15) {real, imag} */,
  {32'h3f6625c5, 32'h3f701cff} /* (8, 1, 14) {real, imag} */,
  {32'hbfacb9cb, 32'h3e984056} /* (8, 1, 13) {real, imag} */,
  {32'hc015236b, 32'hc0919868} /* (8, 1, 12) {real, imag} */,
  {32'h3f1c52cb, 32'h3f933ad1} /* (8, 1, 11) {real, imag} */,
  {32'hbce7a44c, 32'h4022094d} /* (8, 1, 10) {real, imag} */,
  {32'h3d52b90d, 32'hc02c88d2} /* (8, 1, 9) {real, imag} */,
  {32'h40a13655, 32'h3efe2e55} /* (8, 1, 8) {real, imag} */,
  {32'hc0c442bb, 32'hbf6b9e72} /* (8, 1, 7) {real, imag} */,
  {32'h3fe642a9, 32'h3fc18be2} /* (8, 1, 6) {real, imag} */,
  {32'h40ebcf1f, 32'hbf368d25} /* (8, 1, 5) {real, imag} */,
  {32'h3f9a7777, 32'hc0bc6560} /* (8, 1, 4) {real, imag} */,
  {32'h3fd1614c, 32'h3fe58171} /* (8, 1, 3) {real, imag} */,
  {32'h418f193a, 32'hc01920a2} /* (8, 1, 2) {real, imag} */,
  {32'hc1d113d0, 32'h40be6938} /* (8, 1, 1) {real, imag} */,
  {32'hc11b6bdf, 32'h414197be} /* (8, 1, 0) {real, imag} */,
  {32'hc0d6af11, 32'h416fcae3} /* (8, 0, 31) {real, imag} */,
  {32'hbfa65c3b, 32'hc04fd79b} /* (8, 0, 30) {real, imag} */,
  {32'h40251ca1, 32'h3ff25aa9} /* (8, 0, 29) {real, imag} */,
  {32'hc0832be1, 32'hbf28d8af} /* (8, 0, 28) {real, imag} */,
  {32'hbe7c4009, 32'hc0887065} /* (8, 0, 27) {real, imag} */,
  {32'hbfc65bff, 32'hc02e2307} /* (8, 0, 26) {real, imag} */,
  {32'h40514d9d, 32'h4025df23} /* (8, 0, 25) {real, imag} */,
  {32'hc086ec75, 32'hbf329e91} /* (8, 0, 24) {real, imag} */,
  {32'h3fa571d1, 32'h3f91f7f5} /* (8, 0, 23) {real, imag} */,
  {32'hbeb77af3, 32'hbf189f6c} /* (8, 0, 22) {real, imag} */,
  {32'hc031ebdd, 32'hbf3becd8} /* (8, 0, 21) {real, imag} */,
  {32'hbfb4a37b, 32'hbdeb692b} /* (8, 0, 20) {real, imag} */,
  {32'h3e1abb31, 32'hbff820b6} /* (8, 0, 19) {real, imag} */,
  {32'hbf207fda, 32'h3f1d2b1d} /* (8, 0, 18) {real, imag} */,
  {32'hbf84a399, 32'h3e91a3a3} /* (8, 0, 17) {real, imag} */,
  {32'hbf823d68, 32'h3e9eb703} /* (8, 0, 16) {real, imag} */,
  {32'hc01750a2, 32'h4025af6f} /* (8, 0, 15) {real, imag} */,
  {32'h4065b005, 32'h4067e2b1} /* (8, 0, 14) {real, imag} */,
  {32'hbf9b72e1, 32'hbfe4c5ee} /* (8, 0, 13) {real, imag} */,
  {32'hbf86e8e7, 32'h3f970e3b} /* (8, 0, 12) {real, imag} */,
  {32'h3fe6fb1d, 32'hbf5a5215} /* (8, 0, 11) {real, imag} */,
  {32'hc081e7ed, 32'hc0737537} /* (8, 0, 10) {real, imag} */,
  {32'h3fb4db4a, 32'h3fc200f0} /* (8, 0, 9) {real, imag} */,
  {32'h4023b349, 32'hc014b47f} /* (8, 0, 8) {real, imag} */,
  {32'hc09c5354, 32'h40494d7f} /* (8, 0, 7) {real, imag} */,
  {32'h4062294a, 32'h40494b4b} /* (8, 0, 6) {real, imag} */,
  {32'h4085d9f2, 32'hc01066ce} /* (8, 0, 5) {real, imag} */,
  {32'hbec4f62b, 32'h3f992d77} /* (8, 0, 4) {real, imag} */,
  {32'h3f8078cd, 32'hc096e363} /* (8, 0, 3) {real, imag} */,
  {32'h40961550, 32'h4083fece} /* (8, 0, 2) {real, imag} */,
  {32'hc14d4dab, 32'h405f092b} /* (8, 0, 1) {real, imag} */,
  {32'hc0a7ed62, 32'h40ee2d8e} /* (8, 0, 0) {real, imag} */,
  {32'h4068e8f7, 32'hc0cb8ad7} /* (7, 31, 31) {real, imag} */,
  {32'h409be686, 32'h404c82c3} /* (7, 31, 30) {real, imag} */,
  {32'hc10aee11, 32'hbfa2da0b} /* (7, 31, 29) {real, imag} */,
  {32'h3f1acaa7, 32'hc0a3e10e} /* (7, 31, 28) {real, imag} */,
  {32'h400d777a, 32'h4070cacc} /* (7, 31, 27) {real, imag} */,
  {32'hbf0d4940, 32'h4085246d} /* (7, 31, 26) {real, imag} */,
  {32'hbecff1c8, 32'h3e991447} /* (7, 31, 25) {real, imag} */,
  {32'h40369024, 32'hbf8e8671} /* (7, 31, 24) {real, imag} */,
  {32'hc0a4dc9a, 32'hbe8ed65a} /* (7, 31, 23) {real, imag} */,
  {32'h401dff51, 32'hbec4ed4d} /* (7, 31, 22) {real, imag} */,
  {32'h3f61b173, 32'h3f376f89} /* (7, 31, 21) {real, imag} */,
  {32'h3ecb01ee, 32'h3ff0cb9c} /* (7, 31, 20) {real, imag} */,
  {32'h3fc2d836, 32'hbfa1c604} /* (7, 31, 19) {real, imag} */,
  {32'h3fa10d92, 32'hbef20f97} /* (7, 31, 18) {real, imag} */,
  {32'h3f382851, 32'hbf56d160} /* (7, 31, 17) {real, imag} */,
  {32'h3f262fb5, 32'hbe364841} /* (7, 31, 16) {real, imag} */,
  {32'h3f27a5ea, 32'h3e22938b} /* (7, 31, 15) {real, imag} */,
  {32'h3ff1fde2, 32'h3fb045b2} /* (7, 31, 14) {real, imag} */,
  {32'h3f8d5a4c, 32'h3f886406} /* (7, 31, 13) {real, imag} */,
  {32'hbf8d3655, 32'h3ee6f24d} /* (7, 31, 12) {real, imag} */,
  {32'hbfc110d1, 32'h3ffc17f1} /* (7, 31, 11) {real, imag} */,
  {32'hc01999c7, 32'hbf2e109f} /* (7, 31, 10) {real, imag} */,
  {32'h3e84f333, 32'h3fb37ced} /* (7, 31, 9) {real, imag} */,
  {32'hbf18776f, 32'h3f871c2f} /* (7, 31, 8) {real, imag} */,
  {32'hc0258f50, 32'hbea5b3f2} /* (7, 31, 7) {real, imag} */,
  {32'h3fb68ae1, 32'h402372a8} /* (7, 31, 6) {real, imag} */,
  {32'hc05213bc, 32'h3f496679} /* (7, 31, 5) {real, imag} */,
  {32'hc0a68f88, 32'hc0970734} /* (7, 31, 4) {real, imag} */,
  {32'hbbec520d, 32'hc0171c6d} /* (7, 31, 3) {real, imag} */,
  {32'h3f8cfb77, 32'h40bf5f84} /* (7, 31, 2) {real, imag} */,
  {32'hbfe2bdb8, 32'h4027109d} /* (7, 31, 1) {real, imag} */,
  {32'hc06de830, 32'hc0592fd6} /* (7, 31, 0) {real, imag} */,
  {32'hbfe79119, 32'h3f92dbe8} /* (7, 30, 31) {real, imag} */,
  {32'hbf813f21, 32'hbeba3ebf} /* (7, 30, 30) {real, imag} */,
  {32'h3f86a6ec, 32'hc0879d66} /* (7, 30, 29) {real, imag} */,
  {32'hbf8fbde9, 32'hc016e88b} /* (7, 30, 28) {real, imag} */,
  {32'h3fe0f596, 32'h3f2c02c5} /* (7, 30, 27) {real, imag} */,
  {32'h40700ad4, 32'h3ea14461} /* (7, 30, 26) {real, imag} */,
  {32'hc08f712b, 32'hc034d699} /* (7, 30, 25) {real, imag} */,
  {32'h401ad3e7, 32'hbfbc43bf} /* (7, 30, 24) {real, imag} */,
  {32'hbfd79df7, 32'hc037d647} /* (7, 30, 23) {real, imag} */,
  {32'hc0219a48, 32'h40589fe4} /* (7, 30, 22) {real, imag} */,
  {32'hbf73e0de, 32'h3ff8a3b5} /* (7, 30, 21) {real, imag} */,
  {32'hbf633759, 32'h4076ccbb} /* (7, 30, 20) {real, imag} */,
  {32'hbf33e7dd, 32'h3f8a925b} /* (7, 30, 19) {real, imag} */,
  {32'hbee92878, 32'h3e5ba02e} /* (7, 30, 18) {real, imag} */,
  {32'h3fc03d62, 32'hbfbdf331} /* (7, 30, 17) {real, imag} */,
  {32'h3f8129b8, 32'h3f1ee425} /* (7, 30, 16) {real, imag} */,
  {32'h3f94a303, 32'h3fd30bae} /* (7, 30, 15) {real, imag} */,
  {32'h405541c9, 32'h3edccee1} /* (7, 30, 14) {real, imag} */,
  {32'hbea63fe0, 32'hbd6c7ca7} /* (7, 30, 13) {real, imag} */,
  {32'hbede4394, 32'hbec6b798} /* (7, 30, 12) {real, imag} */,
  {32'h3dc28706, 32'h3f15f0b1} /* (7, 30, 11) {real, imag} */,
  {32'h403ca5ae, 32'hc01f28a5} /* (7, 30, 10) {real, imag} */,
  {32'h3f9e8aba, 32'h3ec566c7} /* (7, 30, 9) {real, imag} */,
  {32'h3f922a96, 32'hbf40fd02} /* (7, 30, 8) {real, imag} */,
  {32'hc0006a83, 32'h3fbe6090} /* (7, 30, 7) {real, imag} */,
  {32'hc0c1711c, 32'h3de3b5aa} /* (7, 30, 6) {real, imag} */,
  {32'h3ee0dc9a, 32'hbf15179d} /* (7, 30, 5) {real, imag} */,
  {32'hc051e869, 32'hc0976d45} /* (7, 30, 4) {real, imag} */,
  {32'h405bfcb1, 32'hc0215fcf} /* (7, 30, 3) {real, imag} */,
  {32'h3f0b72f8, 32'h40b2023a} /* (7, 30, 2) {real, imag} */,
  {32'h408aa45f, 32'h4098329c} /* (7, 30, 1) {real, imag} */,
  {32'hc04bdd0b, 32'h41062499} /* (7, 30, 0) {real, imag} */,
  {32'h3f0fd115, 32'h3fdf7a81} /* (7, 29, 31) {real, imag} */,
  {32'hc0a0f453, 32'hbee710bf} /* (7, 29, 30) {real, imag} */,
  {32'hc02a712f, 32'hbf6b5194} /* (7, 29, 29) {real, imag} */,
  {32'hc007f4f2, 32'hbf94fcc1} /* (7, 29, 28) {real, imag} */,
  {32'h40a3f6f6, 32'hbf43d54f} /* (7, 29, 27) {real, imag} */,
  {32'h3ee35f1a, 32'h4094bdc4} /* (7, 29, 26) {real, imag} */,
  {32'hc04dd678, 32'h3f32882b} /* (7, 29, 25) {real, imag} */,
  {32'h3f1ab382, 32'h3c3427f9} /* (7, 29, 24) {real, imag} */,
  {32'h3fc49393, 32'h3f49c880} /* (7, 29, 23) {real, imag} */,
  {32'hbfed66db, 32'hc06b0d21} /* (7, 29, 22) {real, imag} */,
  {32'h3e115a20, 32'hbf17388b} /* (7, 29, 21) {real, imag} */,
  {32'hbf0febdd, 32'h3be703ab} /* (7, 29, 20) {real, imag} */,
  {32'hbe061ac6, 32'h3fc94652} /* (7, 29, 19) {real, imag} */,
  {32'hbf607120, 32'hbfb19713} /* (7, 29, 18) {real, imag} */,
  {32'h3f186b3a, 32'h3dd57f25} /* (7, 29, 17) {real, imag} */,
  {32'h3fae9413, 32'h3f1b55bf} /* (7, 29, 16) {real, imag} */,
  {32'hbf9f0acb, 32'h3f98f736} /* (7, 29, 15) {real, imag} */,
  {32'hbd833d21, 32'hc0372b1d} /* (7, 29, 14) {real, imag} */,
  {32'hbeb18947, 32'h3fae9cf4} /* (7, 29, 13) {real, imag} */,
  {32'hbeba95ab, 32'h40251d64} /* (7, 29, 12) {real, imag} */,
  {32'hbfa70fd9, 32'h4019cbf9} /* (7, 29, 11) {real, imag} */,
  {32'hbe8b299f, 32'h3fb13bb7} /* (7, 29, 10) {real, imag} */,
  {32'hbff0c34a, 32'hc0216c6e} /* (7, 29, 9) {real, imag} */,
  {32'h3faa5918, 32'h3f84dc9a} /* (7, 29, 8) {real, imag} */,
  {32'h400080b8, 32'h405ec89a} /* (7, 29, 7) {real, imag} */,
  {32'hc028d608, 32'hbe6d5bf1} /* (7, 29, 6) {real, imag} */,
  {32'hbf7959e5, 32'h40bf3dfb} /* (7, 29, 5) {real, imag} */,
  {32'hc017ebe2, 32'hbfa3bcbe} /* (7, 29, 4) {real, imag} */,
  {32'h3f7ea417, 32'h3b94497a} /* (7, 29, 3) {real, imag} */,
  {32'h3f67d955, 32'hbfb6ea18} /* (7, 29, 2) {real, imag} */,
  {32'hbfbcb86f, 32'h3f92d748} /* (7, 29, 1) {real, imag} */,
  {32'hc0b21258, 32'h401a3c4c} /* (7, 29, 0) {real, imag} */,
  {32'hbf800a15, 32'h40347513} /* (7, 28, 31) {real, imag} */,
  {32'hbf8d3102, 32'h3fd7acfb} /* (7, 28, 30) {real, imag} */,
  {32'h3f3947e7, 32'hc0660463} /* (7, 28, 29) {real, imag} */,
  {32'h4097ffdf, 32'hbe25ad08} /* (7, 28, 28) {real, imag} */,
  {32'hc054cccf, 32'hbe8f006e} /* (7, 28, 27) {real, imag} */,
  {32'hbd1c1a5d, 32'h4062e029} /* (7, 28, 26) {real, imag} */,
  {32'h3f3606ab, 32'h4010762f} /* (7, 28, 25) {real, imag} */,
  {32'hc02c053c, 32'h404ec698} /* (7, 28, 24) {real, imag} */,
  {32'h401c334e, 32'hbe951e92} /* (7, 28, 23) {real, imag} */,
  {32'h4078b98c, 32'hbf1b4cf3} /* (7, 28, 22) {real, imag} */,
  {32'hc02bae47, 32'h3f5ac2b1} /* (7, 28, 21) {real, imag} */,
  {32'hbfea598b, 32'h3f554d1e} /* (7, 28, 20) {real, imag} */,
  {32'h3fadfc82, 32'hbfbec6c0} /* (7, 28, 19) {real, imag} */,
  {32'hbf6e8591, 32'hbf8477dd} /* (7, 28, 18) {real, imag} */,
  {32'h3f228e00, 32'h3f749824} /* (7, 28, 17) {real, imag} */,
  {32'hbf8c2c54, 32'h3ff2406c} /* (7, 28, 16) {real, imag} */,
  {32'hbeb2a973, 32'h3de4afa5} /* (7, 28, 15) {real, imag} */,
  {32'hbf1f3712, 32'h3f0709ff} /* (7, 28, 14) {real, imag} */,
  {32'h3e79e616, 32'h40266743} /* (7, 28, 13) {real, imag} */,
  {32'hbe9f457f, 32'h3f4418b5} /* (7, 28, 12) {real, imag} */,
  {32'h402e0489, 32'hc025f0c6} /* (7, 28, 11) {real, imag} */,
  {32'h3f669aae, 32'h4005facc} /* (7, 28, 10) {real, imag} */,
  {32'h3fcc925e, 32'hc0116460} /* (7, 28, 9) {real, imag} */,
  {32'hbfb40e98, 32'hbf40f46b} /* (7, 28, 8) {real, imag} */,
  {32'hbeab315d, 32'hbec52236} /* (7, 28, 7) {real, imag} */,
  {32'hbfa38abb, 32'hc0ad94f4} /* (7, 28, 6) {real, imag} */,
  {32'hbfcac4a3, 32'h40004c77} /* (7, 28, 5) {real, imag} */,
  {32'h4008dd6b, 32'hbe696de1} /* (7, 28, 4) {real, imag} */,
  {32'h3f4886bc, 32'h3fc2225a} /* (7, 28, 3) {real, imag} */,
  {32'h3c42d5f9, 32'hc004103e} /* (7, 28, 2) {real, imag} */,
  {32'hbf8afdc5, 32'hbfa31a5b} /* (7, 28, 1) {real, imag} */,
  {32'h3f5ff2dc, 32'hc0994c7c} /* (7, 28, 0) {real, imag} */,
  {32'hc03fbc73, 32'h4056ff46} /* (7, 27, 31) {real, imag} */,
  {32'h3f713ea1, 32'h3ff0373c} /* (7, 27, 30) {real, imag} */,
  {32'h3faceb19, 32'hc027a32c} /* (7, 27, 29) {real, imag} */,
  {32'hbe8ea19f, 32'hc0b92a0d} /* (7, 27, 28) {real, imag} */,
  {32'h3eac8b80, 32'h40113fe1} /* (7, 27, 27) {real, imag} */,
  {32'h3e79655b, 32'hbf2564c2} /* (7, 27, 26) {real, imag} */,
  {32'h3ef0185d, 32'h3feac28a} /* (7, 27, 25) {real, imag} */,
  {32'hbfd8510b, 32'h3ea1a95c} /* (7, 27, 24) {real, imag} */,
  {32'h3fc29a73, 32'h40ae67fa} /* (7, 27, 23) {real, imag} */,
  {32'h3c6a9c97, 32'hbf0fa9e5} /* (7, 27, 22) {real, imag} */,
  {32'hbfe46ccb, 32'hbfa8b3fd} /* (7, 27, 21) {real, imag} */,
  {32'hbfc147c5, 32'h3f9febb3} /* (7, 27, 20) {real, imag} */,
  {32'h3f1f9a8c, 32'hbf4936ad} /* (7, 27, 19) {real, imag} */,
  {32'h403f747b, 32'hbed3fa3c} /* (7, 27, 18) {real, imag} */,
  {32'hbe556e1c, 32'hbdfca2b6} /* (7, 27, 17) {real, imag} */,
  {32'hbf27abc3, 32'hbf286e1e} /* (7, 27, 16) {real, imag} */,
  {32'h3f185986, 32'hbe524a8e} /* (7, 27, 15) {real, imag} */,
  {32'h3d59f182, 32'hbe31fd63} /* (7, 27, 14) {real, imag} */,
  {32'hbfcbb8da, 32'hbf7f6ae8} /* (7, 27, 13) {real, imag} */,
  {32'hbfced8dd, 32'h4008dbf8} /* (7, 27, 12) {real, imag} */,
  {32'h3fe5848d, 32'hbf7fa0f7} /* (7, 27, 11) {real, imag} */,
  {32'hc038eecb, 32'h40162d06} /* (7, 27, 10) {real, imag} */,
  {32'h40394646, 32'hbf6d576d} /* (7, 27, 9) {real, imag} */,
  {32'hbe31e65e, 32'h403fef90} /* (7, 27, 8) {real, imag} */,
  {32'h3f238a05, 32'h3fe369b1} /* (7, 27, 7) {real, imag} */,
  {32'h40855bfa, 32'hc0ab1488} /* (7, 27, 6) {real, imag} */,
  {32'hc0199c66, 32'h3ed1dfe8} /* (7, 27, 5) {real, imag} */,
  {32'hc029aee3, 32'h40ab7e79} /* (7, 27, 4) {real, imag} */,
  {32'hbec1525b, 32'h402517d8} /* (7, 27, 3) {real, imag} */,
  {32'hc07db18d, 32'hc0185c1a} /* (7, 27, 2) {real, imag} */,
  {32'hc0720a53, 32'hc0485b11} /* (7, 27, 1) {real, imag} */,
  {32'h407281a3, 32'h40756d0d} /* (7, 27, 0) {real, imag} */,
  {32'hc03b792f, 32'h405c08c3} /* (7, 26, 31) {real, imag} */,
  {32'hbe8e1bbc, 32'hbf60c3ee} /* (7, 26, 30) {real, imag} */,
  {32'h3f80a608, 32'h3fbba8cd} /* (7, 26, 29) {real, imag} */,
  {32'hc04919a3, 32'hbebb88a5} /* (7, 26, 28) {real, imag} */,
  {32'hc002e719, 32'hc02cfe3e} /* (7, 26, 27) {real, imag} */,
  {32'hc016d649, 32'hc0013895} /* (7, 26, 26) {real, imag} */,
  {32'h40205d4a, 32'hbfad8b31} /* (7, 26, 25) {real, imag} */,
  {32'hbf9e549c, 32'h3c050659} /* (7, 26, 24) {real, imag} */,
  {32'h3e4941a2, 32'h3fbd7ecf} /* (7, 26, 23) {real, imag} */,
  {32'hc03c049b, 32'hc04e663f} /* (7, 26, 22) {real, imag} */,
  {32'hbe9c5afb, 32'hc05a0f47} /* (7, 26, 21) {real, imag} */,
  {32'h40701070, 32'hbfb220d4} /* (7, 26, 20) {real, imag} */,
  {32'hbff40732, 32'hbd9a4371} /* (7, 26, 19) {real, imag} */,
  {32'hbfd10fc3, 32'h4018bfda} /* (7, 26, 18) {real, imag} */,
  {32'h3e900ffe, 32'h3f3f5571} /* (7, 26, 17) {real, imag} */,
  {32'hbf926d46, 32'hbfb97530} /* (7, 26, 16) {real, imag} */,
  {32'hbf036fdb, 32'h3f135e27} /* (7, 26, 15) {real, imag} */,
  {32'h4010e53d, 32'h3f9073d9} /* (7, 26, 14) {real, imag} */,
  {32'h40898a11, 32'hbfba6daf} /* (7, 26, 13) {real, imag} */,
  {32'hbf488a66, 32'hc0376fd6} /* (7, 26, 12) {real, imag} */,
  {32'hbf44a57f, 32'h40055130} /* (7, 26, 11) {real, imag} */,
  {32'hbd0d4d99, 32'h3f9460b5} /* (7, 26, 10) {real, imag} */,
  {32'hc04525c2, 32'hbd9e1569} /* (7, 26, 9) {real, imag} */,
  {32'h3e728368, 32'h3fc47650} /* (7, 26, 8) {real, imag} */,
  {32'hc07046e4, 32'h3f4fc5d4} /* (7, 26, 7) {real, imag} */,
  {32'h3f8c5624, 32'h3fd1fee0} /* (7, 26, 6) {real, imag} */,
  {32'h401cdd73, 32'hbd2e1018} /* (7, 26, 5) {real, imag} */,
  {32'hbf88f9e8, 32'hc0870178} /* (7, 26, 4) {real, imag} */,
  {32'hc016845a, 32'h3fa59e29} /* (7, 26, 3) {real, imag} */,
  {32'h3de6eea5, 32'h3e7d0efb} /* (7, 26, 2) {real, imag} */,
  {32'hbf35bb0e, 32'h3f19fd84} /* (7, 26, 1) {real, imag} */,
  {32'hbceb9042, 32'h3ee33e1a} /* (7, 26, 0) {real, imag} */,
  {32'h4066b529, 32'h3fca23e8} /* (7, 25, 31) {real, imag} */,
  {32'hbfb15e50, 32'h3f8d2d8a} /* (7, 25, 30) {real, imag} */,
  {32'h3fc44635, 32'h3fa664e7} /* (7, 25, 29) {real, imag} */,
  {32'hc06a25e8, 32'hc04e9404} /* (7, 25, 28) {real, imag} */,
  {32'h3d34f8aa, 32'h400ee6c1} /* (7, 25, 27) {real, imag} */,
  {32'h3fee95e3, 32'hbfa2f374} /* (7, 25, 26) {real, imag} */,
  {32'hbff8c758, 32'hbe5fc453} /* (7, 25, 25) {real, imag} */,
  {32'hbfc8bb9f, 32'h3fef260c} /* (7, 25, 24) {real, imag} */,
  {32'h3f72c04d, 32'hc005451b} /* (7, 25, 23) {real, imag} */,
  {32'hc010031c, 32'hbf259c04} /* (7, 25, 22) {real, imag} */,
  {32'h3d6a1faa, 32'h3e2e1fc0} /* (7, 25, 21) {real, imag} */,
  {32'hbfc893b9, 32'hbfa784a3} /* (7, 25, 20) {real, imag} */,
  {32'hc063d9ab, 32'hbfb9a933} /* (7, 25, 19) {real, imag} */,
  {32'h3eef9cba, 32'hc03262bb} /* (7, 25, 18) {real, imag} */,
  {32'hbf2c2040, 32'h4012e86c} /* (7, 25, 17) {real, imag} */,
  {32'h401057f3, 32'h3f657e48} /* (7, 25, 16) {real, imag} */,
  {32'h40283944, 32'h3f002186} /* (7, 25, 15) {real, imag} */,
  {32'h3f1fddbb, 32'h3d14a311} /* (7, 25, 14) {real, imag} */,
  {32'h3f95c039, 32'hc02b94c7} /* (7, 25, 13) {real, imag} */,
  {32'h40339067, 32'h4034c106} /* (7, 25, 12) {real, imag} */,
  {32'hc00bc072, 32'hbf875cc3} /* (7, 25, 11) {real, imag} */,
  {32'h402fe286, 32'h403907de} /* (7, 25, 10) {real, imag} */,
  {32'h3f373123, 32'h3f76bd35} /* (7, 25, 9) {real, imag} */,
  {32'hbf483117, 32'hbfc0fcfa} /* (7, 25, 8) {real, imag} */,
  {32'hbf1b2a95, 32'h400524f1} /* (7, 25, 7) {real, imag} */,
  {32'h403ebdac, 32'h404c3564} /* (7, 25, 6) {real, imag} */,
  {32'hc0481e53, 32'hbe107608} /* (7, 25, 5) {real, imag} */,
  {32'h4042cb8a, 32'h409023b1} /* (7, 25, 4) {real, imag} */,
  {32'hbeffbd60, 32'h3f8e316f} /* (7, 25, 3) {real, imag} */,
  {32'hbfd850c5, 32'h3fe7a685} /* (7, 25, 2) {real, imag} */,
  {32'hc034d32b, 32'h3dfc8988} /* (7, 25, 1) {real, imag} */,
  {32'h4000264f, 32'hbf599dbf} /* (7, 25, 0) {real, imag} */,
  {32'hc037661b, 32'hbfd27834} /* (7, 24, 31) {real, imag} */,
  {32'h3d23f5aa, 32'h400ba12e} /* (7, 24, 30) {real, imag} */,
  {32'h3f3e9cc2, 32'h403b5d72} /* (7, 24, 29) {real, imag} */,
  {32'h400ce7f1, 32'hbe5d07bf} /* (7, 24, 28) {real, imag} */,
  {32'h4064e831, 32'h402c0855} /* (7, 24, 27) {real, imag} */,
  {32'h4014f1c4, 32'hbfaab159} /* (7, 24, 26) {real, imag} */,
  {32'h4101ce9f, 32'hbeae6215} /* (7, 24, 25) {real, imag} */,
  {32'hbefd97f8, 32'hbf874c03} /* (7, 24, 24) {real, imag} */,
  {32'h3ebab182, 32'hbd1debbb} /* (7, 24, 23) {real, imag} */,
  {32'hc0098752, 32'h3fc6d864} /* (7, 24, 22) {real, imag} */,
  {32'h3d904e1b, 32'h3efc1d03} /* (7, 24, 21) {real, imag} */,
  {32'h3f2ad0c8, 32'h402927cb} /* (7, 24, 20) {real, imag} */,
  {32'h3f43aa5e, 32'h3ecc9e77} /* (7, 24, 19) {real, imag} */,
  {32'hbd99ec20, 32'hc0668c58} /* (7, 24, 18) {real, imag} */,
  {32'hbf2b55b9, 32'h3e5fa53c} /* (7, 24, 17) {real, imag} */,
  {32'h3e5b46d3, 32'h3e95b079} /* (7, 24, 16) {real, imag} */,
  {32'h3f8a4fd2, 32'h401349e4} /* (7, 24, 15) {real, imag} */,
  {32'h3d8cb9f9, 32'h3d2d2ccd} /* (7, 24, 14) {real, imag} */,
  {32'h3fe03012, 32'hbfc2d7de} /* (7, 24, 13) {real, imag} */,
  {32'hbf874c59, 32'h40893d08} /* (7, 24, 12) {real, imag} */,
  {32'h3eb2194c, 32'hbfdacd19} /* (7, 24, 11) {real, imag} */,
  {32'hc074ad83, 32'hc087adbf} /* (7, 24, 10) {real, imag} */,
  {32'hc05d8ea6, 32'hbf86c429} /* (7, 24, 9) {real, imag} */,
  {32'hbfcd447b, 32'hbf964edf} /* (7, 24, 8) {real, imag} */,
  {32'h4088d6b5, 32'hc013b311} /* (7, 24, 7) {real, imag} */,
  {32'hbf8aaa69, 32'h3ffe393d} /* (7, 24, 6) {real, imag} */,
  {32'hc008191a, 32'h3edab1e6} /* (7, 24, 5) {real, imag} */,
  {32'hbffec264, 32'h400e16f1} /* (7, 24, 4) {real, imag} */,
  {32'h4039f3c6, 32'hbf910dc0} /* (7, 24, 3) {real, imag} */,
  {32'hc01d2db7, 32'h3eab2c8b} /* (7, 24, 2) {real, imag} */,
  {32'hbf8ee309, 32'h3fdf9817} /* (7, 24, 1) {real, imag} */,
  {32'h3e912429, 32'hc0801be2} /* (7, 24, 0) {real, imag} */,
  {32'hc0137502, 32'h4038c94a} /* (7, 23, 31) {real, imag} */,
  {32'h405087c9, 32'hbfdd0dd7} /* (7, 23, 30) {real, imag} */,
  {32'h3d6e8eb2, 32'hc08a21fe} /* (7, 23, 29) {real, imag} */,
  {32'h4040df5b, 32'h40005af6} /* (7, 23, 28) {real, imag} */,
  {32'hc02a38ee, 32'h3fb18aa0} /* (7, 23, 27) {real, imag} */,
  {32'hbfc737e8, 32'hc05da5f9} /* (7, 23, 26) {real, imag} */,
  {32'h3de2bb33, 32'hbfa4cd42} /* (7, 23, 25) {real, imag} */,
  {32'h3fa1c425, 32'hbf953a26} /* (7, 23, 24) {real, imag} */,
  {32'hc0891b86, 32'h4012b38e} /* (7, 23, 23) {real, imag} */,
  {32'h40915297, 32'hbfb5f3a4} /* (7, 23, 22) {real, imag} */,
  {32'hbe8ac951, 32'h3f94fa15} /* (7, 23, 21) {real, imag} */,
  {32'hbfcb1f91, 32'hbf2404b4} /* (7, 23, 20) {real, imag} */,
  {32'h4049b386, 32'hbf6555aa} /* (7, 23, 19) {real, imag} */,
  {32'h3ecb6a11, 32'h40380633} /* (7, 23, 18) {real, imag} */,
  {32'h3f870cc0, 32'h4017a7a2} /* (7, 23, 17) {real, imag} */,
  {32'h3f60a407, 32'hbe406be1} /* (7, 23, 16) {real, imag} */,
  {32'h3e0b1c4a, 32'hbea24a9d} /* (7, 23, 15) {real, imag} */,
  {32'hbf89432d, 32'hbf82aa9f} /* (7, 23, 14) {real, imag} */,
  {32'hc09258fc, 32'h3db4b317} /* (7, 23, 13) {real, imag} */,
  {32'hbefcafe0, 32'h3ea4da65} /* (7, 23, 12) {real, imag} */,
  {32'h3f2a71ff, 32'h3fa2a80d} /* (7, 23, 11) {real, imag} */,
  {32'hbf3f3152, 32'h3f999b27} /* (7, 23, 10) {real, imag} */,
  {32'h3f011a70, 32'h3ea82b33} /* (7, 23, 9) {real, imag} */,
  {32'h401144d9, 32'h3e01e74e} /* (7, 23, 8) {real, imag} */,
  {32'hbe939064, 32'hc0787d39} /* (7, 23, 7) {real, imag} */,
  {32'hbeb620a8, 32'h3f759de7} /* (7, 23, 6) {real, imag} */,
  {32'h3faa5e2b, 32'h3f0c2a22} /* (7, 23, 5) {real, imag} */,
  {32'hbf544b44, 32'hbdbcc4d1} /* (7, 23, 4) {real, imag} */,
  {32'hbecb3d53, 32'hbdcf21d9} /* (7, 23, 3) {real, imag} */,
  {32'h3fba631f, 32'h3f1b2d85} /* (7, 23, 2) {real, imag} */,
  {32'h402287bb, 32'h404295c9} /* (7, 23, 1) {real, imag} */,
  {32'hbf1da61d, 32'hbf37c8c9} /* (7, 23, 0) {real, imag} */,
  {32'h3fdb5fb2, 32'hc02480b0} /* (7, 22, 31) {real, imag} */,
  {32'h3fd37b96, 32'hc071d9d8} /* (7, 22, 30) {real, imag} */,
  {32'hc04029f9, 32'h4030f40a} /* (7, 22, 29) {real, imag} */,
  {32'h402bf9e0, 32'h40055c6d} /* (7, 22, 28) {real, imag} */,
  {32'hc00b7bc3, 32'h3f57fc91} /* (7, 22, 27) {real, imag} */,
  {32'hc02ca6ba, 32'hc00b549e} /* (7, 22, 26) {real, imag} */,
  {32'hbdc5c2b8, 32'hbe91df38} /* (7, 22, 25) {real, imag} */,
  {32'h3e362b96, 32'hc009c2b4} /* (7, 22, 24) {real, imag} */,
  {32'hbf4e0c87, 32'h40535a25} /* (7, 22, 23) {real, imag} */,
  {32'hbf9e1d1d, 32'h3f573d1b} /* (7, 22, 22) {real, imag} */,
  {32'h3f82231e, 32'hc02675fe} /* (7, 22, 21) {real, imag} */,
  {32'h3fb118f6, 32'h403cf0f3} /* (7, 22, 20) {real, imag} */,
  {32'hbfff7609, 32'hc0450184} /* (7, 22, 19) {real, imag} */,
  {32'h3edafee1, 32'h3fb00ecf} /* (7, 22, 18) {real, imag} */,
  {32'hbf824fef, 32'h3f106367} /* (7, 22, 17) {real, imag} */,
  {32'h3f9a75a0, 32'h402c1d35} /* (7, 22, 16) {real, imag} */,
  {32'h3f155a2c, 32'h3f831a1a} /* (7, 22, 15) {real, imag} */,
  {32'hc006521a, 32'h3efad008} /* (7, 22, 14) {real, imag} */,
  {32'hbf593cf1, 32'h401a08f9} /* (7, 22, 13) {real, imag} */,
  {32'h3fde7928, 32'h3ca010c6} /* (7, 22, 12) {real, imag} */,
  {32'hbf00dece, 32'hbe819277} /* (7, 22, 11) {real, imag} */,
  {32'hc0807991, 32'h3fc441f8} /* (7, 22, 10) {real, imag} */,
  {32'h4060c6d7, 32'hc08542cf} /* (7, 22, 9) {real, imag} */,
  {32'h3e030052, 32'hbf6cd4f3} /* (7, 22, 8) {real, imag} */,
  {32'h3cb2c4fe, 32'hc05e8a9f} /* (7, 22, 7) {real, imag} */,
  {32'h4007e108, 32'hbfcb18ba} /* (7, 22, 6) {real, imag} */,
  {32'hbe0a7780, 32'hbf7455dc} /* (7, 22, 5) {real, imag} */,
  {32'h3f9f7f62, 32'h4057c049} /* (7, 22, 4) {real, imag} */,
  {32'hbf113990, 32'h3fa03c48} /* (7, 22, 3) {real, imag} */,
  {32'h3e11cd5f, 32'h40aca365} /* (7, 22, 2) {real, imag} */,
  {32'h3dc81d00, 32'h3f35d16f} /* (7, 22, 1) {real, imag} */,
  {32'h3e90b0cc, 32'hbfa4d4e3} /* (7, 22, 0) {real, imag} */,
  {32'h403bf995, 32'hc0281c4f} /* (7, 21, 31) {real, imag} */,
  {32'hbfaa6f32, 32'hbd404f0d} /* (7, 21, 30) {real, imag} */,
  {32'hbf3a7f20, 32'hbff302e4} /* (7, 21, 29) {real, imag} */,
  {32'h3f544c06, 32'h400f0dc8} /* (7, 21, 28) {real, imag} */,
  {32'hc076fc7d, 32'hbdcfe68e} /* (7, 21, 27) {real, imag} */,
  {32'h3fa46ec4, 32'hbebd6389} /* (7, 21, 26) {real, imag} */,
  {32'hbf437ee5, 32'h40011797} /* (7, 21, 25) {real, imag} */,
  {32'hc0149d5f, 32'h3f9dfb61} /* (7, 21, 24) {real, imag} */,
  {32'h3fb09922, 32'hc07dff7a} /* (7, 21, 23) {real, imag} */,
  {32'h3ea7a224, 32'h40145936} /* (7, 21, 22) {real, imag} */,
  {32'h4061c0fd, 32'h3f15e517} /* (7, 21, 21) {real, imag} */,
  {32'hbfa23a02, 32'hc01f0ac7} /* (7, 21, 20) {real, imag} */,
  {32'h4003ce88, 32'hbf97f2d0} /* (7, 21, 19) {real, imag} */,
  {32'h3fccb2be, 32'h3f0d5a92} /* (7, 21, 18) {real, imag} */,
  {32'hc00af3fb, 32'hbef9b51d} /* (7, 21, 17) {real, imag} */,
  {32'hbf61a597, 32'hbfde0e2f} /* (7, 21, 16) {real, imag} */,
  {32'hbec2fdc3, 32'h40581fc3} /* (7, 21, 15) {real, imag} */,
  {32'hc0225058, 32'hc0450dc8} /* (7, 21, 14) {real, imag} */,
  {32'hbfaea4ab, 32'hbf3e32d2} /* (7, 21, 13) {real, imag} */,
  {32'hc01c233e, 32'h400012ac} /* (7, 21, 12) {real, imag} */,
  {32'hc00d2dfd, 32'hbf808387} /* (7, 21, 11) {real, imag} */,
  {32'h3f058c0d, 32'hbfd52d6c} /* (7, 21, 10) {real, imag} */,
  {32'h40639b7c, 32'h3ec594da} /* (7, 21, 9) {real, imag} */,
  {32'hbff34f11, 32'hbf5c461d} /* (7, 21, 8) {real, imag} */,
  {32'h40358be4, 32'h3ea2bc6d} /* (7, 21, 7) {real, imag} */,
  {32'h4009b8de, 32'hbfb596d2} /* (7, 21, 6) {real, imag} */,
  {32'hbe5933c7, 32'hbfc135a4} /* (7, 21, 5) {real, imag} */,
  {32'h400273bf, 32'h3ec692c8} /* (7, 21, 4) {real, imag} */,
  {32'hc0218a65, 32'hbe2eb095} /* (7, 21, 3) {real, imag} */,
  {32'h3f9f0110, 32'hbee4b66a} /* (7, 21, 2) {real, imag} */,
  {32'hbf59bd6f, 32'hbf1d2d3e} /* (7, 21, 1) {real, imag} */,
  {32'hbe36d0c6, 32'hbef2d20c} /* (7, 21, 0) {real, imag} */,
  {32'h3d918fd0, 32'hbe9ab044} /* (7, 20, 31) {real, imag} */,
  {32'hbebcfc20, 32'h3f38bb78} /* (7, 20, 30) {real, imag} */,
  {32'h3fbb9325, 32'h3f8d93bd} /* (7, 20, 29) {real, imag} */,
  {32'h3e11cbfa, 32'hc01aacff} /* (7, 20, 28) {real, imag} */,
  {32'h3fc0ad6b, 32'h3e2f8e16} /* (7, 20, 27) {real, imag} */,
  {32'hbfc02ce2, 32'h3f9e4b8d} /* (7, 20, 26) {real, imag} */,
  {32'hbed2e008, 32'hbf722a60} /* (7, 20, 25) {real, imag} */,
  {32'h3f513613, 32'h408b0214} /* (7, 20, 24) {real, imag} */,
  {32'h3e856b01, 32'hbe8e0ddb} /* (7, 20, 23) {real, imag} */,
  {32'h3fa7722d, 32'h40768dae} /* (7, 20, 22) {real, imag} */,
  {32'h3fb0f92a, 32'h3d6d9197} /* (7, 20, 21) {real, imag} */,
  {32'hc080d573, 32'h40021192} /* (7, 20, 20) {real, imag} */,
  {32'h3f0e0ad4, 32'hbe5fb4e4} /* (7, 20, 19) {real, imag} */,
  {32'hbeb0c5af, 32'h40472c74} /* (7, 20, 18) {real, imag} */,
  {32'hbfc0d69a, 32'hbfdf0c0f} /* (7, 20, 17) {real, imag} */,
  {32'h3fafa264, 32'h3e42cc09} /* (7, 20, 16) {real, imag} */,
  {32'hbe7ef06e, 32'hbf888aba} /* (7, 20, 15) {real, imag} */,
  {32'hbf047930, 32'h3f7a7ef3} /* (7, 20, 14) {real, imag} */,
  {32'hbfd707d0, 32'hbfb3238f} /* (7, 20, 13) {real, imag} */,
  {32'hbfd5d06b, 32'hc0a5364b} /* (7, 20, 12) {real, imag} */,
  {32'hc0045569, 32'h3fbdaed7} /* (7, 20, 11) {real, imag} */,
  {32'hbeb7b1a4, 32'h3fb7fc28} /* (7, 20, 10) {real, imag} */,
  {32'hc049f94c, 32'h40264cf7} /* (7, 20, 9) {real, imag} */,
  {32'hc029b92c, 32'hbf28da70} /* (7, 20, 8) {real, imag} */,
  {32'h3fafc5ef, 32'h404f6365} /* (7, 20, 7) {real, imag} */,
  {32'hc0432499, 32'hbe6e4534} /* (7, 20, 6) {real, imag} */,
  {32'h3ebcd6c9, 32'hbf2e195c} /* (7, 20, 5) {real, imag} */,
  {32'h3e60f4be, 32'hc02b78ad} /* (7, 20, 4) {real, imag} */,
  {32'hbf9ca249, 32'hbe55988b} /* (7, 20, 3) {real, imag} */,
  {32'h402821b8, 32'h3f40d907} /* (7, 20, 2) {real, imag} */,
  {32'hbf3af07c, 32'hbfe26905} /* (7, 20, 1) {real, imag} */,
  {32'h3f97e552, 32'h3f9d3c56} /* (7, 20, 0) {real, imag} */,
  {32'h3f262e97, 32'hbff0d895} /* (7, 19, 31) {real, imag} */,
  {32'h4084294f, 32'hbf840c9c} /* (7, 19, 30) {real, imag} */,
  {32'hbf89aabf, 32'h3fd6ba76} /* (7, 19, 29) {real, imag} */,
  {32'hbf23a618, 32'h3feb17d8} /* (7, 19, 28) {real, imag} */,
  {32'hbf0ddcfe, 32'hbf1f3417} /* (7, 19, 27) {real, imag} */,
  {32'hbf47a981, 32'hbf3924bb} /* (7, 19, 26) {real, imag} */,
  {32'hc027e3f3, 32'h40b1d856} /* (7, 19, 25) {real, imag} */,
  {32'hbe017fd9, 32'hbead39ea} /* (7, 19, 24) {real, imag} */,
  {32'h3fc5c3db, 32'h3fa13dcd} /* (7, 19, 23) {real, imag} */,
  {32'h402deb20, 32'h3fee7d63} /* (7, 19, 22) {real, imag} */,
  {32'hbf857d93, 32'hbf11d507} /* (7, 19, 21) {real, imag} */,
  {32'hbed4ee49, 32'hbfd6137e} /* (7, 19, 20) {real, imag} */,
  {32'hbeeba876, 32'h3e631e52} /* (7, 19, 19) {real, imag} */,
  {32'hbfd36005, 32'h3e01f51b} /* (7, 19, 18) {real, imag} */,
  {32'hbfbe03d8, 32'h3fc0088e} /* (7, 19, 17) {real, imag} */,
  {32'h3f4baf5c, 32'hc00e00e1} /* (7, 19, 16) {real, imag} */,
  {32'hbe077a2e, 32'hc00b8c51} /* (7, 19, 15) {real, imag} */,
  {32'h3e332537, 32'h3e59d887} /* (7, 19, 14) {real, imag} */,
  {32'hbed08cc3, 32'h400323ee} /* (7, 19, 13) {real, imag} */,
  {32'h40cb9fbc, 32'h3e2103d7} /* (7, 19, 12) {real, imag} */,
  {32'h3ff8721b, 32'h4009e436} /* (7, 19, 11) {real, imag} */,
  {32'h3f1f4344, 32'h3f297030} /* (7, 19, 10) {real, imag} */,
  {32'h3e8e7e07, 32'hbef00bc2} /* (7, 19, 9) {real, imag} */,
  {32'hbf79b1de, 32'hbf20ed1e} /* (7, 19, 8) {real, imag} */,
  {32'h3f024e7a, 32'h3f069717} /* (7, 19, 7) {real, imag} */,
  {32'h3f1673e2, 32'h40164f26} /* (7, 19, 6) {real, imag} */,
  {32'hbf987d1b, 32'hbf0af0f9} /* (7, 19, 5) {real, imag} */,
  {32'hbe57abb1, 32'h3f15eec7} /* (7, 19, 4) {real, imag} */,
  {32'hbf91308d, 32'h3fdeddd4} /* (7, 19, 3) {real, imag} */,
  {32'h3f6fb035, 32'hc043ed04} /* (7, 19, 2) {real, imag} */,
  {32'h3fa25e28, 32'hbe548924} /* (7, 19, 1) {real, imag} */,
  {32'h3eb5398c, 32'hbede21fe} /* (7, 19, 0) {real, imag} */,
  {32'hbf9afbf9, 32'h3faa0d60} /* (7, 18, 31) {real, imag} */,
  {32'hc01af198, 32'hbedca988} /* (7, 18, 30) {real, imag} */,
  {32'h3f4d6d30, 32'h3fbb7bef} /* (7, 18, 29) {real, imag} */,
  {32'h3fa95a1e, 32'h3f9c3a2d} /* (7, 18, 28) {real, imag} */,
  {32'hc04ea44b, 32'h406b25d1} /* (7, 18, 27) {real, imag} */,
  {32'hc0173f50, 32'hbe347af2} /* (7, 18, 26) {real, imag} */,
  {32'h3f01ae9a, 32'hbc209c8f} /* (7, 18, 25) {real, imag} */,
  {32'hbea58867, 32'h401f9997} /* (7, 18, 24) {real, imag} */,
  {32'hbf75fbf6, 32'h3f8b220b} /* (7, 18, 23) {real, imag} */,
  {32'hbd13bf43, 32'hc085d41a} /* (7, 18, 22) {real, imag} */,
  {32'h3f622db0, 32'h3f5c267d} /* (7, 18, 21) {real, imag} */,
  {32'h3e9906f7, 32'hbf06037e} /* (7, 18, 20) {real, imag} */,
  {32'h3fbbf043, 32'hbfa3010a} /* (7, 18, 19) {real, imag} */,
  {32'h3e2d2737, 32'h3e899ac5} /* (7, 18, 18) {real, imag} */,
  {32'hbe97cc0b, 32'h3fa05456} /* (7, 18, 17) {real, imag} */,
  {32'hbf8a56e9, 32'h3f723e58} /* (7, 18, 16) {real, imag} */,
  {32'hc003a7f0, 32'hbee89d27} /* (7, 18, 15) {real, imag} */,
  {32'h40796360, 32'h3f021318} /* (7, 18, 14) {real, imag} */,
  {32'h3ffe6a6d, 32'hbedc09d4} /* (7, 18, 13) {real, imag} */,
  {32'h3fdf6a80, 32'h3f90d508} /* (7, 18, 12) {real, imag} */,
  {32'h3fd96b3f, 32'hbef7b129} /* (7, 18, 11) {real, imag} */,
  {32'h3fa9b172, 32'h3f9af729} /* (7, 18, 10) {real, imag} */,
  {32'h401e250c, 32'hbf0f00a3} /* (7, 18, 9) {real, imag} */,
  {32'h3fdfb0d2, 32'h4009300b} /* (7, 18, 8) {real, imag} */,
  {32'h3e5f59b1, 32'h40564956} /* (7, 18, 7) {real, imag} */,
  {32'hbf877631, 32'hbfd23621} /* (7, 18, 6) {real, imag} */,
  {32'hbe329080, 32'h3e6f3313} /* (7, 18, 5) {real, imag} */,
  {32'hbffb3af8, 32'hbfa869c8} /* (7, 18, 4) {real, imag} */,
  {32'hc0223d72, 32'hbea20400} /* (7, 18, 3) {real, imag} */,
  {32'h3eed62fd, 32'h3faa0f87} /* (7, 18, 2) {real, imag} */,
  {32'hbf662bb9, 32'h3ef0c974} /* (7, 18, 1) {real, imag} */,
  {32'h3fe5e6c2, 32'h3f3787a5} /* (7, 18, 0) {real, imag} */,
  {32'h3ef15289, 32'hbf486477} /* (7, 17, 31) {real, imag} */,
  {32'h3e360d5f, 32'hbe2da011} /* (7, 17, 30) {real, imag} */,
  {32'hbf3aa749, 32'h3ebaeb17} /* (7, 17, 29) {real, imag} */,
  {32'h3ea37ec4, 32'h3f3c7c3e} /* (7, 17, 28) {real, imag} */,
  {32'h3e94c45a, 32'h3e02a6b6} /* (7, 17, 27) {real, imag} */,
  {32'h3ffaa34f, 32'h3fd5a930} /* (7, 17, 26) {real, imag} */,
  {32'h3ea3e728, 32'hbfbb78c5} /* (7, 17, 25) {real, imag} */,
  {32'h3f81070c, 32'hc00e346b} /* (7, 17, 24) {real, imag} */,
  {32'hbef9e0a7, 32'hbf06be46} /* (7, 17, 23) {real, imag} */,
  {32'hbf59370e, 32'hbf988d09} /* (7, 17, 22) {real, imag} */,
  {32'hc05b5b37, 32'hbc916eba} /* (7, 17, 21) {real, imag} */,
  {32'h3f364cd1, 32'h3f0bb3ee} /* (7, 17, 20) {real, imag} */,
  {32'hbfb8ff5a, 32'h3ff356bb} /* (7, 17, 19) {real, imag} */,
  {32'h3fb42991, 32'h3d7a5fba} /* (7, 17, 18) {real, imag} */,
  {32'hbf166896, 32'h3f6629a9} /* (7, 17, 17) {real, imag} */,
  {32'h3fb9237f, 32'hbed8a814} /* (7, 17, 16) {real, imag} */,
  {32'h3fba0dcf, 32'h4001a687} /* (7, 17, 15) {real, imag} */,
  {32'h3f911546, 32'h40347030} /* (7, 17, 14) {real, imag} */,
  {32'h405706dc, 32'hbff1c3bc} /* (7, 17, 13) {real, imag} */,
  {32'hbf5c21bf, 32'hbf05d98e} /* (7, 17, 12) {real, imag} */,
  {32'h3e811573, 32'hbfa8a98a} /* (7, 17, 11) {real, imag} */,
  {32'h3e2d7dc7, 32'h3f13ad2f} /* (7, 17, 10) {real, imag} */,
  {32'hbf34f635, 32'h400ac1a1} /* (7, 17, 9) {real, imag} */,
  {32'hbed7cbd3, 32'h3f74d578} /* (7, 17, 8) {real, imag} */,
  {32'hbeae7891, 32'hbf10c45f} /* (7, 17, 7) {real, imag} */,
  {32'hc01a8d6a, 32'h3ffe4c24} /* (7, 17, 6) {real, imag} */,
  {32'hbf694bbb, 32'h3e01bb0e} /* (7, 17, 5) {real, imag} */,
  {32'hbf56352f, 32'hbe9ea328} /* (7, 17, 4) {real, imag} */,
  {32'h3f3f6200, 32'hbf0755a2} /* (7, 17, 3) {real, imag} */,
  {32'h3f2284a5, 32'hc01c1511} /* (7, 17, 2) {real, imag} */,
  {32'hb9c1e304, 32'h3f7a7696} /* (7, 17, 1) {real, imag} */,
  {32'hc03876ba, 32'h3f497afe} /* (7, 17, 0) {real, imag} */,
  {32'h3f97c8bd, 32'h3f6fb3b0} /* (7, 16, 31) {real, imag} */,
  {32'hbfaf0435, 32'hbf9f4fc2} /* (7, 16, 30) {real, imag} */,
  {32'h3fbe6281, 32'hbf7fbcb4} /* (7, 16, 29) {real, imag} */,
  {32'h401ec460, 32'h3cc53534} /* (7, 16, 28) {real, imag} */,
  {32'hbf2035cd, 32'hbd1b7da2} /* (7, 16, 27) {real, imag} */,
  {32'hbfecb8ed, 32'hbf8d8dfd} /* (7, 16, 26) {real, imag} */,
  {32'h3f23bcfd, 32'hbf522bf7} /* (7, 16, 25) {real, imag} */,
  {32'h3f9f1295, 32'h3e5f0f1e} /* (7, 16, 24) {real, imag} */,
  {32'hbe9b7a05, 32'hbf193395} /* (7, 16, 23) {real, imag} */,
  {32'h3f231a3a, 32'h3ec9683c} /* (7, 16, 22) {real, imag} */,
  {32'h3f6feefb, 32'h3f910997} /* (7, 16, 21) {real, imag} */,
  {32'hbfc624e3, 32'hbf85be44} /* (7, 16, 20) {real, imag} */,
  {32'h3f9a0680, 32'hc00e57ed} /* (7, 16, 19) {real, imag} */,
  {32'hbf8f029d, 32'hbfa76cac} /* (7, 16, 18) {real, imag} */,
  {32'hbfd953f7, 32'h3ea42a8c} /* (7, 16, 17) {real, imag} */,
  {32'hbe9f30cd, 32'hbf4e425a} /* (7, 16, 16) {real, imag} */,
  {32'h3f05ec40, 32'hbe3497fe} /* (7, 16, 15) {real, imag} */,
  {32'hbf006ce2, 32'hbf5eb722} /* (7, 16, 14) {real, imag} */,
  {32'h3d9273be, 32'hbfc7d5d3} /* (7, 16, 13) {real, imag} */,
  {32'h3e8a2cb0, 32'h3e6b4a78} /* (7, 16, 12) {real, imag} */,
  {32'hbf2764eb, 32'h400c599c} /* (7, 16, 11) {real, imag} */,
  {32'hbf848481, 32'hc01523b5} /* (7, 16, 10) {real, imag} */,
  {32'h3e25f9b4, 32'h40128930} /* (7, 16, 9) {real, imag} */,
  {32'h3e456aa9, 32'h3fc232c7} /* (7, 16, 8) {real, imag} */,
  {32'hc0122a6c, 32'h3be52054} /* (7, 16, 7) {real, imag} */,
  {32'h3ede3b84, 32'h3f1018ed} /* (7, 16, 6) {real, imag} */,
  {32'h3f23ccd1, 32'h3f53eb2c} /* (7, 16, 5) {real, imag} */,
  {32'hbe2afca9, 32'h3f3c9573} /* (7, 16, 4) {real, imag} */,
  {32'h3e81a4d1, 32'hbf043e83} /* (7, 16, 3) {real, imag} */,
  {32'hbfd0a00f, 32'hbd80fa73} /* (7, 16, 2) {real, imag} */,
  {32'hbff80ce5, 32'hbf8a7217} /* (7, 16, 1) {real, imag} */,
  {32'h3eb7f7ac, 32'h3cf99927} /* (7, 16, 0) {real, imag} */,
  {32'h3f7b2db4, 32'hbf5d1e9d} /* (7, 15, 31) {real, imag} */,
  {32'hbfb2f9da, 32'hbf27b1a8} /* (7, 15, 30) {real, imag} */,
  {32'hbe862136, 32'h3f034495} /* (7, 15, 29) {real, imag} */,
  {32'hbe414179, 32'h3ff4910a} /* (7, 15, 28) {real, imag} */,
  {32'h3b640088, 32'h3fca3336} /* (7, 15, 27) {real, imag} */,
  {32'hbd3d5b74, 32'hbfc36fea} /* (7, 15, 26) {real, imag} */,
  {32'h405eacc1, 32'h3f20879c} /* (7, 15, 25) {real, imag} */,
  {32'hbf99b70b, 32'h3fb508f1} /* (7, 15, 24) {real, imag} */,
  {32'h3f8d8c16, 32'hbfa18e99} /* (7, 15, 23) {real, imag} */,
  {32'h3e86bc5f, 32'h4016d28b} /* (7, 15, 22) {real, imag} */,
  {32'h40153ee6, 32'hbf9964f3} /* (7, 15, 21) {real, imag} */,
  {32'hbf26a59a, 32'h3f19f8ad} /* (7, 15, 20) {real, imag} */,
  {32'h3f2e1f8d, 32'h3d783c9a} /* (7, 15, 19) {real, imag} */,
  {32'h3fc39922, 32'h3f1ec5f8} /* (7, 15, 18) {real, imag} */,
  {32'h3f91f03c, 32'hbeba9a7c} /* (7, 15, 17) {real, imag} */,
  {32'hbda9cc77, 32'h3ea4554b} /* (7, 15, 16) {real, imag} */,
  {32'h3eec6bae, 32'hbf028615} /* (7, 15, 15) {real, imag} */,
  {32'hbfe277dd, 32'hbbede588} /* (7, 15, 14) {real, imag} */,
  {32'h3e8c63df, 32'h3f98278b} /* (7, 15, 13) {real, imag} */,
  {32'hbf8439b6, 32'hbf13e63a} /* (7, 15, 12) {real, imag} */,
  {32'hbe9ddd8b, 32'h3fb22cff} /* (7, 15, 11) {real, imag} */,
  {32'hc01c61a6, 32'hbf42e323} /* (7, 15, 10) {real, imag} */,
  {32'h3fab7c65, 32'h3fff3ccf} /* (7, 15, 9) {real, imag} */,
  {32'hbd61144c, 32'hc009138e} /* (7, 15, 8) {real, imag} */,
  {32'h4007dd80, 32'h400b0c3d} /* (7, 15, 7) {real, imag} */,
  {32'hbdbce961, 32'h3f3368e2} /* (7, 15, 6) {real, imag} */,
  {32'h3e876d37, 32'h3ff9ec34} /* (7, 15, 5) {real, imag} */,
  {32'h3efb557a, 32'hc0081e1e} /* (7, 15, 4) {real, imag} */,
  {32'h3f435af4, 32'hbeb7508b} /* (7, 15, 3) {real, imag} */,
  {32'h3f0ff1a4, 32'hbf978770} /* (7, 15, 2) {real, imag} */,
  {32'h3e831aa6, 32'hc029a2db} /* (7, 15, 1) {real, imag} */,
  {32'hc0268683, 32'hbf329d11} /* (7, 15, 0) {real, imag} */,
  {32'hbe8ed0ef, 32'hbe15a1a1} /* (7, 14, 31) {real, imag} */,
  {32'h3ed1c043, 32'h3f67891c} /* (7, 14, 30) {real, imag} */,
  {32'h3fcce273, 32'h3f888e98} /* (7, 14, 29) {real, imag} */,
  {32'hbf23ce66, 32'hbfe68395} /* (7, 14, 28) {real, imag} */,
  {32'h3ffe556b, 32'hc07b378a} /* (7, 14, 27) {real, imag} */,
  {32'hc03d7015, 32'h3fa98cbe} /* (7, 14, 26) {real, imag} */,
  {32'h3fd501c7, 32'hbfdcf48f} /* (7, 14, 25) {real, imag} */,
  {32'hbed67745, 32'h3fcda9a3} /* (7, 14, 24) {real, imag} */,
  {32'hbed2744f, 32'h3f0fb9e0} /* (7, 14, 23) {real, imag} */,
  {32'hbea47d0a, 32'hbfcc4da8} /* (7, 14, 22) {real, imag} */,
  {32'hbf864bf2, 32'h3fed7c89} /* (7, 14, 21) {real, imag} */,
  {32'h3eee4c49, 32'hbfb0bd40} /* (7, 14, 20) {real, imag} */,
  {32'h3f31a221, 32'hbeffa280} /* (7, 14, 19) {real, imag} */,
  {32'h3ff43218, 32'h3f46f779} /* (7, 14, 18) {real, imag} */,
  {32'h4003bcb6, 32'hbd02ae1d} /* (7, 14, 17) {real, imag} */,
  {32'h3f2650a9, 32'h3e9c9530} /* (7, 14, 16) {real, imag} */,
  {32'hbe5d5e3f, 32'hbfaf99b5} /* (7, 14, 15) {real, imag} */,
  {32'hbf118ee8, 32'h3f620893} /* (7, 14, 14) {real, imag} */,
  {32'hbfaafe91, 32'h3f9ade1a} /* (7, 14, 13) {real, imag} */,
  {32'h400f3d49, 32'h3f699d75} /* (7, 14, 12) {real, imag} */,
  {32'h3f2d7ac7, 32'hbf441b1b} /* (7, 14, 11) {real, imag} */,
  {32'h3fba3072, 32'hbfc5c3c0} /* (7, 14, 10) {real, imag} */,
  {32'hbf257f75, 32'hbfa4c3cb} /* (7, 14, 9) {real, imag} */,
  {32'hbf9cc512, 32'hbecf681d} /* (7, 14, 8) {real, imag} */,
  {32'h4033d0e1, 32'hbf28f05e} /* (7, 14, 7) {real, imag} */,
  {32'h4059f775, 32'hbfb8a1a4} /* (7, 14, 6) {real, imag} */,
  {32'h3e4ec77c, 32'h3ea98952} /* (7, 14, 5) {real, imag} */,
  {32'hbe8d9d81, 32'h3f6768d9} /* (7, 14, 4) {real, imag} */,
  {32'h3f6db535, 32'h3e3849b4} /* (7, 14, 3) {real, imag} */,
  {32'hbf224c3f, 32'h3fe80e65} /* (7, 14, 2) {real, imag} */,
  {32'hc01a0610, 32'h3f63e6c0} /* (7, 14, 1) {real, imag} */,
  {32'hbf667ac2, 32'h3d992f4b} /* (7, 14, 0) {real, imag} */,
  {32'hbe3a8b13, 32'h3ed217f5} /* (7, 13, 31) {real, imag} */,
  {32'h3f888216, 32'h3f3f463c} /* (7, 13, 30) {real, imag} */,
  {32'hc029f1be, 32'hc0166653} /* (7, 13, 29) {real, imag} */,
  {32'hbfea11f1, 32'hbf8b20d2} /* (7, 13, 28) {real, imag} */,
  {32'h4018056d, 32'h3ee5da2c} /* (7, 13, 27) {real, imag} */,
  {32'hbfbbb70e, 32'hbf83fdbc} /* (7, 13, 26) {real, imag} */,
  {32'hbf0c2a30, 32'h3e61a092} /* (7, 13, 25) {real, imag} */,
  {32'h402af66a, 32'hbdc856f9} /* (7, 13, 24) {real, imag} */,
  {32'h3d183abb, 32'h3f831c5f} /* (7, 13, 23) {real, imag} */,
  {32'h3f27bb7e, 32'h3fd127f5} /* (7, 13, 22) {real, imag} */,
  {32'h3e9ac23b, 32'hc025ae06} /* (7, 13, 21) {real, imag} */,
  {32'hbf98f727, 32'h4054ac24} /* (7, 13, 20) {real, imag} */,
  {32'hbe5302fb, 32'hbff0f51c} /* (7, 13, 19) {real, imag} */,
  {32'hbe9f4233, 32'h40584bee} /* (7, 13, 18) {real, imag} */,
  {32'hbf5ba566, 32'h3df619a6} /* (7, 13, 17) {real, imag} */,
  {32'h402fc34c, 32'h3f176334} /* (7, 13, 16) {real, imag} */,
  {32'h3de9fa41, 32'h406c9397} /* (7, 13, 15) {real, imag} */,
  {32'hbfea4233, 32'hc048145b} /* (7, 13, 14) {real, imag} */,
  {32'h3fc91cc4, 32'hbffbd3ac} /* (7, 13, 13) {real, imag} */,
  {32'h3f4e893f, 32'h3f7a9da4} /* (7, 13, 12) {real, imag} */,
  {32'h40171035, 32'h3f10280a} /* (7, 13, 11) {real, imag} */,
  {32'h3f9e8f4d, 32'h3fa57906} /* (7, 13, 10) {real, imag} */,
  {32'h3f06957c, 32'h402c416f} /* (7, 13, 9) {real, imag} */,
  {32'hbf4f9ff1, 32'hbdd300d6} /* (7, 13, 8) {real, imag} */,
  {32'hc009039b, 32'h3fc1b0ba} /* (7, 13, 7) {real, imag} */,
  {32'hbf81af2e, 32'hc09b8d57} /* (7, 13, 6) {real, imag} */,
  {32'h3f96fbb2, 32'hbd7d0153} /* (7, 13, 5) {real, imag} */,
  {32'hbef111bc, 32'h3fa630fa} /* (7, 13, 4) {real, imag} */,
  {32'h3d1733f4, 32'hbea2bcbe} /* (7, 13, 3) {real, imag} */,
  {32'h3f8e9bed, 32'h3f091130} /* (7, 13, 2) {real, imag} */,
  {32'h403430c5, 32'hbf19b11e} /* (7, 13, 1) {real, imag} */,
  {32'hbfd2c82e, 32'hc013469e} /* (7, 13, 0) {real, imag} */,
  {32'h3e3779bd, 32'hbfdf4905} /* (7, 12, 31) {real, imag} */,
  {32'hbf0d2110, 32'hbf89cae3} /* (7, 12, 30) {real, imag} */,
  {32'hbf1aa9d7, 32'h40195999} /* (7, 12, 29) {real, imag} */,
  {32'hbd925de7, 32'hc05a310b} /* (7, 12, 28) {real, imag} */,
  {32'hbf9fe78d, 32'h3f9f9927} /* (7, 12, 27) {real, imag} */,
  {32'hbe3362e9, 32'hc096585f} /* (7, 12, 26) {real, imag} */,
  {32'hbf865ab2, 32'hbfc95300} /* (7, 12, 25) {real, imag} */,
  {32'hbff75c93, 32'h3fd3f5b7} /* (7, 12, 24) {real, imag} */,
  {32'h400f87c2, 32'h3d4a2d87} /* (7, 12, 23) {real, imag} */,
  {32'h3f88ee07, 32'h3f352065} /* (7, 12, 22) {real, imag} */,
  {32'h4036aa15, 32'h40a4b64c} /* (7, 12, 21) {real, imag} */,
  {32'h3eb5d95b, 32'hbf5789ce} /* (7, 12, 20) {real, imag} */,
  {32'h405feaac, 32'hbfe82c2f} /* (7, 12, 19) {real, imag} */,
  {32'h3f77bcda, 32'hc00bb020} /* (7, 12, 18) {real, imag} */,
  {32'hbfd942d3, 32'hc0250f22} /* (7, 12, 17) {real, imag} */,
  {32'hbf303f5b, 32'hbf662205} /* (7, 12, 16) {real, imag} */,
  {32'h3efbb759, 32'hbfcb7b51} /* (7, 12, 15) {real, imag} */,
  {32'hbff9f654, 32'hbfbb2b5f} /* (7, 12, 14) {real, imag} */,
  {32'h3f74a211, 32'hbf934a72} /* (7, 12, 13) {real, imag} */,
  {32'hbf40b06d, 32'h3feb6d64} /* (7, 12, 12) {real, imag} */,
  {32'hbda7b70e, 32'h3f778469} /* (7, 12, 11) {real, imag} */,
  {32'hbfe489be, 32'h3f8b01a2} /* (7, 12, 10) {real, imag} */,
  {32'h40703106, 32'h4014e6b3} /* (7, 12, 9) {real, imag} */,
  {32'h3eb7b0a3, 32'hc088fcb4} /* (7, 12, 8) {real, imag} */,
  {32'hc00d64db, 32'hbf8df64f} /* (7, 12, 7) {real, imag} */,
  {32'h3e45d243, 32'hbf0ccd11} /* (7, 12, 6) {real, imag} */,
  {32'h403e47e8, 32'h3fea3efe} /* (7, 12, 5) {real, imag} */,
  {32'hbf33493c, 32'hbee0e89f} /* (7, 12, 4) {real, imag} */,
  {32'h3e81c4bd, 32'h3e86d6b1} /* (7, 12, 3) {real, imag} */,
  {32'hbf5dcef1, 32'hbf1dbf4c} /* (7, 12, 2) {real, imag} */,
  {32'hbf104d9a, 32'h3fc46b2b} /* (7, 12, 1) {real, imag} */,
  {32'hbe62ab3b, 32'hbf517cde} /* (7, 12, 0) {real, imag} */,
  {32'hbfd780e9, 32'h3e6199e8} /* (7, 11, 31) {real, imag} */,
  {32'hbffc01d9, 32'hc022df3e} /* (7, 11, 30) {real, imag} */,
  {32'hc0263923, 32'h3fd3ba86} /* (7, 11, 29) {real, imag} */,
  {32'hbe642d64, 32'h3f1aaecf} /* (7, 11, 28) {real, imag} */,
  {32'h405fa76b, 32'h406b4251} /* (7, 11, 27) {real, imag} */,
  {32'hbe056a2a, 32'hbf993dd2} /* (7, 11, 26) {real, imag} */,
  {32'h3febd5a2, 32'hc00c500f} /* (7, 11, 25) {real, imag} */,
  {32'hbedfb4bb, 32'hc02db096} /* (7, 11, 24) {real, imag} */,
  {32'hbf90687e, 32'hc092aea5} /* (7, 11, 23) {real, imag} */,
  {32'h3f96caef, 32'hbef26764} /* (7, 11, 22) {real, imag} */,
  {32'h3f305e3b, 32'hbe71342c} /* (7, 11, 21) {real, imag} */,
  {32'h3f090b59, 32'h401a8b3c} /* (7, 11, 20) {real, imag} */,
  {32'hbfa964f7, 32'h4006b899} /* (7, 11, 19) {real, imag} */,
  {32'hbf7810be, 32'hbfc574c9} /* (7, 11, 18) {real, imag} */,
  {32'hbdaf0f96, 32'hbe75faa1} /* (7, 11, 17) {real, imag} */,
  {32'h3fe9da91, 32'hbfa9ce0d} /* (7, 11, 16) {real, imag} */,
  {32'hbf3ff85e, 32'h401b032e} /* (7, 11, 15) {real, imag} */,
  {32'h4047c21d, 32'hbe1bacd1} /* (7, 11, 14) {real, imag} */,
  {32'h3fda1f6f, 32'hc092c1df} /* (7, 11, 13) {real, imag} */,
  {32'h3e72b425, 32'hbfbea9ff} /* (7, 11, 12) {real, imag} */,
  {32'hbfeddba4, 32'hbf40d054} /* (7, 11, 11) {real, imag} */,
  {32'hc04e9b08, 32'hbf71ddfe} /* (7, 11, 10) {real, imag} */,
  {32'hc03560cc, 32'h3f95eda9} /* (7, 11, 9) {real, imag} */,
  {32'h3f51b686, 32'hbca25ebd} /* (7, 11, 8) {real, imag} */,
  {32'h40804333, 32'h3f0aab69} /* (7, 11, 7) {real, imag} */,
  {32'hc0153e0d, 32'h400e1857} /* (7, 11, 6) {real, imag} */,
  {32'hbede4b0e, 32'hbf854960} /* (7, 11, 5) {real, imag} */,
  {32'hbf96f087, 32'hbf1d441d} /* (7, 11, 4) {real, imag} */,
  {32'hbf8904f9, 32'h3fd10444} /* (7, 11, 3) {real, imag} */,
  {32'h404771ad, 32'hbfc87e5f} /* (7, 11, 2) {real, imag} */,
  {32'hc06e8f33, 32'hc01bb747} /* (7, 11, 1) {real, imag} */,
  {32'hbf639671, 32'hbf961d0c} /* (7, 11, 0) {real, imag} */,
  {32'h3e643d74, 32'hbfb32e90} /* (7, 10, 31) {real, imag} */,
  {32'hbfc3c00c, 32'hc0438ccd} /* (7, 10, 30) {real, imag} */,
  {32'hbfb1955a, 32'h4032c38a} /* (7, 10, 29) {real, imag} */,
  {32'hc049b161, 32'hbf3e1e78} /* (7, 10, 28) {real, imag} */,
  {32'h3f2d56ff, 32'h3ffee69e} /* (7, 10, 27) {real, imag} */,
  {32'h3f4f84ef, 32'h40650fad} /* (7, 10, 26) {real, imag} */,
  {32'h3ff991d7, 32'hc035c019} /* (7, 10, 25) {real, imag} */,
  {32'h3fbfd717, 32'h400fc79e} /* (7, 10, 24) {real, imag} */,
  {32'hbf4870b5, 32'hc04b4cdb} /* (7, 10, 23) {real, imag} */,
  {32'h4051141d, 32'hbfbab7e9} /* (7, 10, 22) {real, imag} */,
  {32'hc03d7d5d, 32'h3ffbb7aa} /* (7, 10, 21) {real, imag} */,
  {32'hc0372de5, 32'h3f379900} /* (7, 10, 20) {real, imag} */,
  {32'hc0881e30, 32'h3f720a2c} /* (7, 10, 19) {real, imag} */,
  {32'h3f01de98, 32'hbebe48e9} /* (7, 10, 18) {real, imag} */,
  {32'hbd76a4aa, 32'hc0230003} /* (7, 10, 17) {real, imag} */,
  {32'hbe38ae3b, 32'hbe885104} /* (7, 10, 16) {real, imag} */,
  {32'hbf9399d3, 32'h3f0e3783} /* (7, 10, 15) {real, imag} */,
  {32'hbec99b03, 32'hbfae5fc3} /* (7, 10, 14) {real, imag} */,
  {32'hbea2357e, 32'h3fe469c2} /* (7, 10, 13) {real, imag} */,
  {32'h403fc72d, 32'hbfad088f} /* (7, 10, 12) {real, imag} */,
  {32'hbf0dd4fe, 32'h3e6e0e23} /* (7, 10, 11) {real, imag} */,
  {32'h3ef8e661, 32'hc01fcd66} /* (7, 10, 10) {real, imag} */,
  {32'hbe059e56, 32'hbf84e753} /* (7, 10, 9) {real, imag} */,
  {32'hbf3b0651, 32'h3fac6cde} /* (7, 10, 8) {real, imag} */,
  {32'h3faaeb37, 32'h3c8417fd} /* (7, 10, 7) {real, imag} */,
  {32'hbf9b6b54, 32'h3feb90cb} /* (7, 10, 6) {real, imag} */,
  {32'hbfb7276d, 32'h3fb7faf5} /* (7, 10, 5) {real, imag} */,
  {32'hbffdf99e, 32'hbeed29a6} /* (7, 10, 4) {real, imag} */,
  {32'hbeafeff3, 32'hc048c269} /* (7, 10, 3) {real, imag} */,
  {32'h40161005, 32'h40298ee6} /* (7, 10, 2) {real, imag} */,
  {32'h3f0895d2, 32'hbf9073a0} /* (7, 10, 1) {real, imag} */,
  {32'h3fbcf87a, 32'h3e90c6aa} /* (7, 10, 0) {real, imag} */,
  {32'h3f62a0be, 32'hbfd201fb} /* (7, 9, 31) {real, imag} */,
  {32'h3fb9d499, 32'h3eef80d6} /* (7, 9, 30) {real, imag} */,
  {32'hbf42742c, 32'h3f9cf707} /* (7, 9, 29) {real, imag} */,
  {32'h400e4a37, 32'hbe87f8ae} /* (7, 9, 28) {real, imag} */,
  {32'hbf6d5ef7, 32'hbffe01bd} /* (7, 9, 27) {real, imag} */,
  {32'hbfcd55b6, 32'h3eb63c82} /* (7, 9, 26) {real, imag} */,
  {32'h4073acb9, 32'h3f40eaeb} /* (7, 9, 25) {real, imag} */,
  {32'hbbb6b89a, 32'hbfee16b4} /* (7, 9, 24) {real, imag} */,
  {32'h3f96a4e1, 32'hbf0218e5} /* (7, 9, 23) {real, imag} */,
  {32'h404a3bc5, 32'h401a2dee} /* (7, 9, 22) {real, imag} */,
  {32'hc050ea16, 32'h3f943498} /* (7, 9, 21) {real, imag} */,
  {32'hbf95889e, 32'h3ecd7cef} /* (7, 9, 20) {real, imag} */,
  {32'h3fe9b021, 32'hbfe6bb79} /* (7, 9, 19) {real, imag} */,
  {32'h3f6b6e98, 32'hc0008ace} /* (7, 9, 18) {real, imag} */,
  {32'hbf79342f, 32'h3ffa0c8f} /* (7, 9, 17) {real, imag} */,
  {32'h3ee8a782, 32'hbf9d10de} /* (7, 9, 16) {real, imag} */,
  {32'h3eea8939, 32'hbf8aefb8} /* (7, 9, 15) {real, imag} */,
  {32'h3f0b2845, 32'h3fa55e71} /* (7, 9, 14) {real, imag} */,
  {32'h40125509, 32'hbf0745dc} /* (7, 9, 13) {real, imag} */,
  {32'h3f9d821b, 32'h3ee2f59f} /* (7, 9, 12) {real, imag} */,
  {32'hc0112c65, 32'hbf84dfe0} /* (7, 9, 11) {real, imag} */,
  {32'h40389a42, 32'h4067df92} /* (7, 9, 10) {real, imag} */,
  {32'hbf000d26, 32'hc0797eb3} /* (7, 9, 9) {real, imag} */,
  {32'h3ff2d3d5, 32'h3fa065b0} /* (7, 9, 8) {real, imag} */,
  {32'hc00fbd00, 32'h40a88b3f} /* (7, 9, 7) {real, imag} */,
  {32'hbfab900a, 32'hc0666382} /* (7, 9, 6) {real, imag} */,
  {32'hbe131520, 32'hbea153bc} /* (7, 9, 5) {real, imag} */,
  {32'hbf8275d8, 32'h3f978c97} /* (7, 9, 4) {real, imag} */,
  {32'h3d70c82f, 32'h3f1af408} /* (7, 9, 3) {real, imag} */,
  {32'h40b38d30, 32'h3eb84ee4} /* (7, 9, 2) {real, imag} */,
  {32'h3fb97970, 32'h3fad2e6c} /* (7, 9, 1) {real, imag} */,
  {32'hbf826782, 32'h40363344} /* (7, 9, 0) {real, imag} */,
  {32'hbe843ca6, 32'h3f9430c8} /* (7, 8, 31) {real, imag} */,
  {32'hbfaea303, 32'h3f54c91b} /* (7, 8, 30) {real, imag} */,
  {32'h4073d52c, 32'hbe950630} /* (7, 8, 29) {real, imag} */,
  {32'hbf0e7b15, 32'h40549edb} /* (7, 8, 28) {real, imag} */,
  {32'h3fd4c5f4, 32'h40363099} /* (7, 8, 27) {real, imag} */,
  {32'h3f0ec09e, 32'hc07d27c5} /* (7, 8, 26) {real, imag} */,
  {32'hc00fa17b, 32'hbee9d406} /* (7, 8, 25) {real, imag} */,
  {32'hbfbb301d, 32'h3f4091b3} /* (7, 8, 24) {real, imag} */,
  {32'hc0826949, 32'hbf6a2e1e} /* (7, 8, 23) {real, imag} */,
  {32'hbfd30276, 32'hc0265717} /* (7, 8, 22) {real, imag} */,
  {32'hbf70c0dd, 32'h3e6dd0b4} /* (7, 8, 21) {real, imag} */,
  {32'h3efe382a, 32'hbf4cfe3d} /* (7, 8, 20) {real, imag} */,
  {32'h3fe7905f, 32'h3f066abb} /* (7, 8, 19) {real, imag} */,
  {32'hbee35ee8, 32'hbf6daf19} /* (7, 8, 18) {real, imag} */,
  {32'hc02332ab, 32'h3ed9cb7c} /* (7, 8, 17) {real, imag} */,
  {32'hbdde132e, 32'hbfb14b83} /* (7, 8, 16) {real, imag} */,
  {32'hbf1808e9, 32'hc0272339} /* (7, 8, 15) {real, imag} */,
  {32'hbf0cb0ac, 32'h3faaf334} /* (7, 8, 14) {real, imag} */,
  {32'hbe8fa90e, 32'hbf83435b} /* (7, 8, 13) {real, imag} */,
  {32'hc06a6491, 32'h3e3a5ccf} /* (7, 8, 12) {real, imag} */,
  {32'h40aed304, 32'h3f0589a7} /* (7, 8, 11) {real, imag} */,
  {32'h3fc524e9, 32'hc00db481} /* (7, 8, 10) {real, imag} */,
  {32'h405d6e0d, 32'h40412bee} /* (7, 8, 9) {real, imag} */,
  {32'h3f1bfa81, 32'hbe716631} /* (7, 8, 8) {real, imag} */,
  {32'h407b37da, 32'h3f1dfd67} /* (7, 8, 7) {real, imag} */,
  {32'h3fb4ac91, 32'h3f3021ca} /* (7, 8, 6) {real, imag} */,
  {32'hbfd8eb8a, 32'h3f8baa9e} /* (7, 8, 5) {real, imag} */,
  {32'h4021c0b3, 32'h3fc21381} /* (7, 8, 4) {real, imag} */,
  {32'hbc8d55f1, 32'h3e373fd8} /* (7, 8, 3) {real, imag} */,
  {32'hbf5a0c36, 32'hc0107047} /* (7, 8, 2) {real, imag} */,
  {32'hc00f4bed, 32'hc0338d18} /* (7, 8, 1) {real, imag} */,
  {32'h3f46e8bb, 32'h407cfcb6} /* (7, 8, 0) {real, imag} */,
  {32'h3f3b8faf, 32'hbf2438ef} /* (7, 7, 31) {real, imag} */,
  {32'h3fe4795c, 32'h4048b65d} /* (7, 7, 30) {real, imag} */,
  {32'h402d93f1, 32'h40431e13} /* (7, 7, 29) {real, imag} */,
  {32'h3f2478a7, 32'h3f43b812} /* (7, 7, 28) {real, imag} */,
  {32'hbf86a372, 32'h3f1d2347} /* (7, 7, 27) {real, imag} */,
  {32'hc01489d0, 32'hbd51e11c} /* (7, 7, 26) {real, imag} */,
  {32'h3e625e9b, 32'hc027a426} /* (7, 7, 25) {real, imag} */,
  {32'hbee59afd, 32'hbed50136} /* (7, 7, 24) {real, imag} */,
  {32'h3ee65d6b, 32'h3fb83b8d} /* (7, 7, 23) {real, imag} */,
  {32'h4013f104, 32'hbfea99f2} /* (7, 7, 22) {real, imag} */,
  {32'h3ffb70a2, 32'h403fbff3} /* (7, 7, 21) {real, imag} */,
  {32'h4029d02a, 32'hbf7e8993} /* (7, 7, 20) {real, imag} */,
  {32'hbf4a67cc, 32'hbefc7ebb} /* (7, 7, 19) {real, imag} */,
  {32'hbea046fb, 32'h4011ac94} /* (7, 7, 18) {real, imag} */,
  {32'h3f8c6f5a, 32'hbf272456} /* (7, 7, 17) {real, imag} */,
  {32'h3f3c6ba4, 32'h3c524cc6} /* (7, 7, 16) {real, imag} */,
  {32'h3f9d25cd, 32'h3fad5feb} /* (7, 7, 15) {real, imag} */,
  {32'hbdbe2227, 32'hbf70ecb3} /* (7, 7, 14) {real, imag} */,
  {32'h3fe81977, 32'hbf7a188c} /* (7, 7, 13) {real, imag} */,
  {32'hbfa3057b, 32'h3ee219a4} /* (7, 7, 12) {real, imag} */,
  {32'hbd86ed63, 32'h3f663317} /* (7, 7, 11) {real, imag} */,
  {32'hbe5e53c8, 32'hbe84f3a0} /* (7, 7, 10) {real, imag} */,
  {32'hbfea40ab, 32'hc038d59a} /* (7, 7, 9) {real, imag} */,
  {32'h3f339e92, 32'hbfca0900} /* (7, 7, 8) {real, imag} */,
  {32'h4002f005, 32'h3db33e6c} /* (7, 7, 7) {real, imag} */,
  {32'h3e1e7efa, 32'h400ace6b} /* (7, 7, 6) {real, imag} */,
  {32'h3ed9be5d, 32'h404ddeec} /* (7, 7, 5) {real, imag} */,
  {32'hbf8338f1, 32'hbf7a1b2a} /* (7, 7, 4) {real, imag} */,
  {32'hc045c3d9, 32'h3f19e8b0} /* (7, 7, 3) {real, imag} */,
  {32'h3fa5c054, 32'h3fb9ba53} /* (7, 7, 2) {real, imag} */,
  {32'h40161171, 32'hbf8c6339} /* (7, 7, 1) {real, imag} */,
  {32'hc00aba2c, 32'hbf95e35c} /* (7, 7, 0) {real, imag} */,
  {32'hbfee4a2b, 32'hbff72a9a} /* (7, 6, 31) {real, imag} */,
  {32'h408897d5, 32'h3f079b69} /* (7, 6, 30) {real, imag} */,
  {32'h3f128cc0, 32'h404cefe0} /* (7, 6, 29) {real, imag} */,
  {32'h3ed43ec5, 32'h3fcc866d} /* (7, 6, 28) {real, imag} */,
  {32'hc011e565, 32'h402e2e34} /* (7, 6, 27) {real, imag} */,
  {32'hbfd35fe4, 32'h3cebeab9} /* (7, 6, 26) {real, imag} */,
  {32'h4039cbac, 32'hbf39b60f} /* (7, 6, 25) {real, imag} */,
  {32'hbfad50d5, 32'h3f679588} /* (7, 6, 24) {real, imag} */,
  {32'h400ae0bd, 32'h3c996bfa} /* (7, 6, 23) {real, imag} */,
  {32'hc0599002, 32'h3fb4da83} /* (7, 6, 22) {real, imag} */,
  {32'h4020a027, 32'h403aea57} /* (7, 6, 21) {real, imag} */,
  {32'h3e526a36, 32'hbfb9fbc2} /* (7, 6, 20) {real, imag} */,
  {32'hbf8a010d, 32'hc0082647} /* (7, 6, 19) {real, imag} */,
  {32'hbe96ecb4, 32'hbef3f5b9} /* (7, 6, 18) {real, imag} */,
  {32'hbe5f9f43, 32'h3fc18d28} /* (7, 6, 17) {real, imag} */,
  {32'h3e9bfd4a, 32'hbf0b6536} /* (7, 6, 16) {real, imag} */,
  {32'h3ee3b1dc, 32'h3eee8b53} /* (7, 6, 15) {real, imag} */,
  {32'h3f59e21a, 32'hbed42ee7} /* (7, 6, 14) {real, imag} */,
  {32'h3e826534, 32'h40521c35} /* (7, 6, 13) {real, imag} */,
  {32'h3c4bb7a4, 32'hbf90ca8e} /* (7, 6, 12) {real, imag} */,
  {32'hbc3bb38b, 32'h403c6002} /* (7, 6, 11) {real, imag} */,
  {32'h3f46d172, 32'hbf0f966d} /* (7, 6, 10) {real, imag} */,
  {32'h3fa3cbcf, 32'hc01deea7} /* (7, 6, 9) {real, imag} */,
  {32'hc017f1e5, 32'h4006826b} /* (7, 6, 8) {real, imag} */,
  {32'hbf1e9f13, 32'hc009e43e} /* (7, 6, 7) {real, imag} */,
  {32'hbec408c3, 32'hbec9fa3b} /* (7, 6, 6) {real, imag} */,
  {32'hbfe2724e, 32'hbfa8b143} /* (7, 6, 5) {real, imag} */,
  {32'h3fd3a594, 32'h3ebbef6b} /* (7, 6, 4) {real, imag} */,
  {32'hbe87c8cb, 32'hbee06e91} /* (7, 6, 3) {real, imag} */,
  {32'hbfaad2ba, 32'hc048da45} /* (7, 6, 2) {real, imag} */,
  {32'h4084c039, 32'h3ff2eb66} /* (7, 6, 1) {real, imag} */,
  {32'hbe9d8e07, 32'hbf51abcf} /* (7, 6, 0) {real, imag} */,
  {32'h3fc45461, 32'h3fad402b} /* (7, 5, 31) {real, imag} */,
  {32'hbe5254aa, 32'h40e05c31} /* (7, 5, 30) {real, imag} */,
  {32'h3fa5982e, 32'h3ee52088} /* (7, 5, 29) {real, imag} */,
  {32'h3f6f6dcb, 32'hbfe73126} /* (7, 5, 28) {real, imag} */,
  {32'h409a441f, 32'hc036ef07} /* (7, 5, 27) {real, imag} */,
  {32'hc062a917, 32'h3f25012f} /* (7, 5, 26) {real, imag} */,
  {32'h4019b29f, 32'h4099d42b} /* (7, 5, 25) {real, imag} */,
  {32'hbe52d29a, 32'hbfa995b2} /* (7, 5, 24) {real, imag} */,
  {32'h404f4cc7, 32'h40475a97} /* (7, 5, 23) {real, imag} */,
  {32'h3f2b8109, 32'h3eb64880} /* (7, 5, 22) {real, imag} */,
  {32'hbffeec3a, 32'hbf7045b9} /* (7, 5, 21) {real, imag} */,
  {32'hbff78a89, 32'hbf298e58} /* (7, 5, 20) {real, imag} */,
  {32'hc08aca65, 32'h3f242182} /* (7, 5, 19) {real, imag} */,
  {32'h4073a847, 32'h3fb5c189} /* (7, 5, 18) {real, imag} */,
  {32'h3e56715e, 32'h3f75a46c} /* (7, 5, 17) {real, imag} */,
  {32'h3fae5f0b, 32'h3e2f4c76} /* (7, 5, 16) {real, imag} */,
  {32'h3fbb3296, 32'hbf5c0b5b} /* (7, 5, 15) {real, imag} */,
  {32'h3f924607, 32'h3ec87350} /* (7, 5, 14) {real, imag} */,
  {32'h3f8fd92f, 32'hbf8e8160} /* (7, 5, 13) {real, imag} */,
  {32'h3f07ac39, 32'hbfc6ad2c} /* (7, 5, 12) {real, imag} */,
  {32'hbd59ceb8, 32'hc025d394} /* (7, 5, 11) {real, imag} */,
  {32'hbf09a76b, 32'h40a89c3b} /* (7, 5, 10) {real, imag} */,
  {32'h3de9794a, 32'h405276c1} /* (7, 5, 9) {real, imag} */,
  {32'h3f3ff1af, 32'h3fd83755} /* (7, 5, 8) {real, imag} */,
  {32'h40227cc1, 32'hc040f060} /* (7, 5, 7) {real, imag} */,
  {32'hc019f548, 32'h3f1ed62b} /* (7, 5, 6) {real, imag} */,
  {32'hbf6426a4, 32'h3f9b8c82} /* (7, 5, 5) {real, imag} */,
  {32'h3fb4996e, 32'h3ff4ce17} /* (7, 5, 4) {real, imag} */,
  {32'hbf84621c, 32'hc03ea424} /* (7, 5, 3) {real, imag} */,
  {32'hc044a891, 32'h404357c8} /* (7, 5, 2) {real, imag} */,
  {32'hbffb6a83, 32'hbf610af9} /* (7, 5, 1) {real, imag} */,
  {32'h3f9f48c0, 32'hc0cc51fe} /* (7, 5, 0) {real, imag} */,
  {32'h3fdd7fbc, 32'hbff9aba1} /* (7, 4, 31) {real, imag} */,
  {32'h405dc3af, 32'hc091c81a} /* (7, 4, 30) {real, imag} */,
  {32'hbf6db6e9, 32'hc0249f7e} /* (7, 4, 29) {real, imag} */,
  {32'hc0162930, 32'h405439b7} /* (7, 4, 28) {real, imag} */,
  {32'h4071cd51, 32'hc041aad2} /* (7, 4, 27) {real, imag} */,
  {32'hbfcac594, 32'h400457c7} /* (7, 4, 26) {real, imag} */,
  {32'h3f6645d6, 32'h3ff24a22} /* (7, 4, 25) {real, imag} */,
  {32'h40343ddd, 32'h4005b946} /* (7, 4, 24) {real, imag} */,
  {32'hbd7704c9, 32'h3c8c7efa} /* (7, 4, 23) {real, imag} */,
  {32'hbf6d823d, 32'h40694904} /* (7, 4, 22) {real, imag} */,
  {32'hc06bd578, 32'hc002a3e3} /* (7, 4, 21) {real, imag} */,
  {32'h3ef2b476, 32'h3e5baa05} /* (7, 4, 20) {real, imag} */,
  {32'hbfa59aa2, 32'hbe2ac4c3} /* (7, 4, 19) {real, imag} */,
  {32'hbf6efca5, 32'h405997db} /* (7, 4, 18) {real, imag} */,
  {32'hbe80cda6, 32'hbf8cabe5} /* (7, 4, 17) {real, imag} */,
  {32'h3ec07c23, 32'h3ed6a5a2} /* (7, 4, 16) {real, imag} */,
  {32'h3eac0742, 32'hbdf922db} /* (7, 4, 15) {real, imag} */,
  {32'h3ef51379, 32'h40121b86} /* (7, 4, 14) {real, imag} */,
  {32'hc0803d18, 32'hbf7b7788} /* (7, 4, 13) {real, imag} */,
  {32'h3fb39e82, 32'hbfec99e6} /* (7, 4, 12) {real, imag} */,
  {32'h3f95f93d, 32'h40292bf4} /* (7, 4, 11) {real, imag} */,
  {32'h3eaa5e78, 32'hbf99d914} /* (7, 4, 10) {real, imag} */,
  {32'hbfdc52f5, 32'hc007ce17} /* (7, 4, 9) {real, imag} */,
  {32'h402b051e, 32'h4025c588} /* (7, 4, 8) {real, imag} */,
  {32'hc0443ea8, 32'hbfad079a} /* (7, 4, 7) {real, imag} */,
  {32'h3f326465, 32'h400cac98} /* (7, 4, 6) {real, imag} */,
  {32'h3f9b398a, 32'h3fa7aa30} /* (7, 4, 5) {real, imag} */,
  {32'h40a9cd28, 32'hbb8eb776} /* (7, 4, 4) {real, imag} */,
  {32'hc03ca09e, 32'h404abd27} /* (7, 4, 3) {real, imag} */,
  {32'h3fd81941, 32'hc0e6085e} /* (7, 4, 2) {real, imag} */,
  {32'hbedc56f7, 32'h401d25d2} /* (7, 4, 1) {real, imag} */,
  {32'hbf1a5b02, 32'h401fa95b} /* (7, 4, 0) {real, imag} */,
  {32'hc0c361d7, 32'hc097e66b} /* (7, 3, 31) {real, imag} */,
  {32'h3e56f5aa, 32'h403f10aa} /* (7, 3, 30) {real, imag} */,
  {32'hbe020d8f, 32'h40c90093} /* (7, 3, 29) {real, imag} */,
  {32'hbef4b4e7, 32'hc024fce1} /* (7, 3, 28) {real, imag} */,
  {32'h3de8c478, 32'hbfec5eb9} /* (7, 3, 27) {real, imag} */,
  {32'h3fa99b2b, 32'hc01b90fd} /* (7, 3, 26) {real, imag} */,
  {32'h3fb89379, 32'hbf4ed297} /* (7, 3, 25) {real, imag} */,
  {32'h3fdd2b4b, 32'hbe99839d} /* (7, 3, 24) {real, imag} */,
  {32'h3fa3b94b, 32'h40646ebd} /* (7, 3, 23) {real, imag} */,
  {32'hbf2bc28c, 32'h3fcfcb4e} /* (7, 3, 22) {real, imag} */,
  {32'hbe82ad2b, 32'hbf82c020} /* (7, 3, 21) {real, imag} */,
  {32'h404a8983, 32'hc09cb89d} /* (7, 3, 20) {real, imag} */,
  {32'hbf273200, 32'h404ed7f6} /* (7, 3, 19) {real, imag} */,
  {32'h3f6d3472, 32'hbf20433a} /* (7, 3, 18) {real, imag} */,
  {32'hbf1a62a5, 32'hbf50d116} /* (7, 3, 17) {real, imag} */,
  {32'hbf285bad, 32'hbee73729} /* (7, 3, 16) {real, imag} */,
  {32'h3f829fdf, 32'hbeaffe45} /* (7, 3, 15) {real, imag} */,
  {32'hc0897ba4, 32'hbfb37b14} /* (7, 3, 14) {real, imag} */,
  {32'hbe249acf, 32'h3e93e64a} /* (7, 3, 13) {real, imag} */,
  {32'h3f7e4ee4, 32'hc027b10c} /* (7, 3, 12) {real, imag} */,
  {32'h4018e8e9, 32'hbe904283} /* (7, 3, 11) {real, imag} */,
  {32'h3efb8eca, 32'hbfccc4de} /* (7, 3, 10) {real, imag} */,
  {32'h3ea813ed, 32'hc05b232f} /* (7, 3, 9) {real, imag} */,
  {32'h3ea498c6, 32'h3f879e63} /* (7, 3, 8) {real, imag} */,
  {32'hc0837067, 32'h3f11118c} /* (7, 3, 7) {real, imag} */,
  {32'hc026ac0d, 32'h4020d137} /* (7, 3, 6) {real, imag} */,
  {32'hc0145cc2, 32'hc0813cc0} /* (7, 3, 5) {real, imag} */,
  {32'h406b4b67, 32'hbe005b62} /* (7, 3, 4) {real, imag} */,
  {32'h40b7ea11, 32'h3e1bad15} /* (7, 3, 3) {real, imag} */,
  {32'h3fc6b4df, 32'hbfd239b9} /* (7, 3, 2) {real, imag} */,
  {32'h407002c3, 32'h3f5859f4} /* (7, 3, 1) {real, imag} */,
  {32'h40821060, 32'h3eeff27e} /* (7, 3, 0) {real, imag} */,
  {32'hc037f6c1, 32'h403d50d4} /* (7, 2, 31) {real, imag} */,
  {32'hbfeedbdc, 32'hc0bf490c} /* (7, 2, 30) {real, imag} */,
  {32'hc0d9afc8, 32'hc0addadc} /* (7, 2, 29) {real, imag} */,
  {32'h4075b2ad, 32'hc0a43eca} /* (7, 2, 28) {real, imag} */,
  {32'hc02f02fd, 32'h3ff2279f} /* (7, 2, 27) {real, imag} */,
  {32'hbfa52dea, 32'h3f445802} /* (7, 2, 26) {real, imag} */,
  {32'h3ea8ef7a, 32'h4041e13e} /* (7, 2, 25) {real, imag} */,
  {32'h3fadeef4, 32'hc08c29e1} /* (7, 2, 24) {real, imag} */,
  {32'h3fcd4468, 32'h3f169679} /* (7, 2, 23) {real, imag} */,
  {32'hbfcf3ef3, 32'h3f63649c} /* (7, 2, 22) {real, imag} */,
  {32'hc03b03ee, 32'hbef6e33f} /* (7, 2, 21) {real, imag} */,
  {32'h3fe4f444, 32'h3f3328db} /* (7, 2, 20) {real, imag} */,
  {32'hbeb9d596, 32'h3f7ad8ee} /* (7, 2, 19) {real, imag} */,
  {32'h3ea490c1, 32'hbfca6d9e} /* (7, 2, 18) {real, imag} */,
  {32'h3f3b34b3, 32'h40413ea5} /* (7, 2, 17) {real, imag} */,
  {32'h3ea74fbb, 32'hbf848bc9} /* (7, 2, 16) {real, imag} */,
  {32'hbd8fa4b4, 32'h3e5176d8} /* (7, 2, 15) {real, imag} */,
  {32'h3fbc6c46, 32'h3e93095b} /* (7, 2, 14) {real, imag} */,
  {32'hbeb4fcfe, 32'h3ef2b1a0} /* (7, 2, 13) {real, imag} */,
  {32'h3fd49c5f, 32'h3f18b534} /* (7, 2, 12) {real, imag} */,
  {32'hc091ad36, 32'hbff4a0aa} /* (7, 2, 11) {real, imag} */,
  {32'hc05169ec, 32'hbd5e8957} /* (7, 2, 10) {real, imag} */,
  {32'h40708586, 32'h3e861fc6} /* (7, 2, 9) {real, imag} */,
  {32'h3fa0cec5, 32'h3d617b9b} /* (7, 2, 8) {real, imag} */,
  {32'h3f86c24e, 32'hbdd29f9b} /* (7, 2, 7) {real, imag} */,
  {32'hbfd1690d, 32'h3fa3b5fd} /* (7, 2, 6) {real, imag} */,
  {32'h4065cc30, 32'hbfc3022d} /* (7, 2, 5) {real, imag} */,
  {32'h3fbc3799, 32'hbf84f7a0} /* (7, 2, 4) {real, imag} */,
  {32'h40778266, 32'hbe9af201} /* (7, 2, 3) {real, imag} */,
  {32'hc07895b2, 32'hc02c0f95} /* (7, 2, 2) {real, imag} */,
  {32'hbf6b7468, 32'h3fe6bd0a} /* (7, 2, 1) {real, imag} */,
  {32'hbf82554f, 32'h403e8a55} /* (7, 2, 0) {real, imag} */,
  {32'h3de7cae4, 32'hc0f47d5d} /* (7, 1, 31) {real, imag} */,
  {32'hc0c51e8f, 32'h40931558} /* (7, 1, 30) {real, imag} */,
  {32'h3ebcef90, 32'h4001a5cc} /* (7, 1, 29) {real, imag} */,
  {32'h40772e6c, 32'hbfa06ff3} /* (7, 1, 28) {real, imag} */,
  {32'h402b6528, 32'h40c76abe} /* (7, 1, 27) {real, imag} */,
  {32'h3f886cd6, 32'h3f4faf88} /* (7, 1, 26) {real, imag} */,
  {32'h3fe24452, 32'h409dbc5b} /* (7, 1, 25) {real, imag} */,
  {32'h3f461ace, 32'hbfe8a5a4} /* (7, 1, 24) {real, imag} */,
  {32'h3fc57399, 32'hc091676b} /* (7, 1, 23) {real, imag} */,
  {32'hc08dfb6f, 32'h3fb1550d} /* (7, 1, 22) {real, imag} */,
  {32'hbff1cbbb, 32'hbfbc7764} /* (7, 1, 21) {real, imag} */,
  {32'hbfc55d66, 32'h3fe21a43} /* (7, 1, 20) {real, imag} */,
  {32'h3f9db8d9, 32'hc00c15a5} /* (7, 1, 19) {real, imag} */,
  {32'hc00bad2c, 32'h3f809ccf} /* (7, 1, 18) {real, imag} */,
  {32'hbf02c5c8, 32'h3f9767f4} /* (7, 1, 17) {real, imag} */,
  {32'h3f197904, 32'hbee462f4} /* (7, 1, 16) {real, imag} */,
  {32'hbf279ac2, 32'h3f4069d9} /* (7, 1, 15) {real, imag} */,
  {32'h3e16bb1f, 32'hbfd336e0} /* (7, 1, 14) {real, imag} */,
  {32'h3fbc0a26, 32'h3f0f296c} /* (7, 1, 13) {real, imag} */,
  {32'h3d48f037, 32'h3fa65995} /* (7, 1, 12) {real, imag} */,
  {32'hbf836365, 32'hc0369d50} /* (7, 1, 11) {real, imag} */,
  {32'hc0556c23, 32'hbf9fa9ee} /* (7, 1, 10) {real, imag} */,
  {32'h3f008fc9, 32'hbda75a67} /* (7, 1, 9) {real, imag} */,
  {32'hbfa65773, 32'hbe97de3b} /* (7, 1, 8) {real, imag} */,
  {32'h3d16874d, 32'h3fdd2beb} /* (7, 1, 7) {real, imag} */,
  {32'h40629c76, 32'hc0d22625} /* (7, 1, 6) {real, imag} */,
  {32'hbf4d7b3e, 32'hbfa97efa} /* (7, 1, 5) {real, imag} */,
  {32'h3d3be098, 32'h3dcfd68d} /* (7, 1, 4) {real, imag} */,
  {32'hbdd3430e, 32'hc09a65ea} /* (7, 1, 3) {real, imag} */,
  {32'hc0490f6d, 32'h40a2cb24} /* (7, 1, 2) {real, imag} */,
  {32'h409763a3, 32'hc07a1664} /* (7, 1, 1) {real, imag} */,
  {32'h3f6fab2c, 32'h406c72c2} /* (7, 1, 0) {real, imag} */,
  {32'hbc38e6f5, 32'h40596853} /* (7, 0, 31) {real, imag} */,
  {32'hbf386261, 32'h3f9f3684} /* (7, 0, 30) {real, imag} */,
  {32'hbfbe7592, 32'h3fc9b686} /* (7, 0, 29) {real, imag} */,
  {32'hbfe22fa1, 32'h40b5d2c9} /* (7, 0, 28) {real, imag} */,
  {32'hbf689f13, 32'h40694b1d} /* (7, 0, 27) {real, imag} */,
  {32'h408d96a7, 32'hbfcba01b} /* (7, 0, 26) {real, imag} */,
  {32'h3f1aaa81, 32'hbbef4a07} /* (7, 0, 25) {real, imag} */,
  {32'h3fc5f2c2, 32'h402e0a14} /* (7, 0, 24) {real, imag} */,
  {32'hbfa9afed, 32'hbf07a34a} /* (7, 0, 23) {real, imag} */,
  {32'hc06963cd, 32'hbc837845} /* (7, 0, 22) {real, imag} */,
  {32'h3f95c853, 32'hbfa24fd5} /* (7, 0, 21) {real, imag} */,
  {32'h3fc8cd3d, 32'h3f867565} /* (7, 0, 20) {real, imag} */,
  {32'h3fddd953, 32'h3df4e206} /* (7, 0, 19) {real, imag} */,
  {32'hbeca1760, 32'hbe79220f} /* (7, 0, 18) {real, imag} */,
  {32'hbfea1094, 32'h404d2377} /* (7, 0, 17) {real, imag} */,
  {32'hbf89737c, 32'hbf9c7286} /* (7, 0, 16) {real, imag} */,
  {32'hbf6faf1f, 32'hbfc2275f} /* (7, 0, 15) {real, imag} */,
  {32'h3f7306fc, 32'hbf16bda2} /* (7, 0, 14) {real, imag} */,
  {32'hbfce0a37, 32'h403c9796} /* (7, 0, 13) {real, imag} */,
  {32'h3e917c57, 32'hc0879cbb} /* (7, 0, 12) {real, imag} */,
  {32'hc02726a4, 32'hbfc4fcdd} /* (7, 0, 11) {real, imag} */,
  {32'hbe2481f8, 32'hbfb968d7} /* (7, 0, 10) {real, imag} */,
  {32'hbea07ab2, 32'h401a5b47} /* (7, 0, 9) {real, imag} */,
  {32'h4000e5e6, 32'hbf895439} /* (7, 0, 8) {real, imag} */,
  {32'hbf532a8e, 32'hc023aabd} /* (7, 0, 7) {real, imag} */,
  {32'h40584196, 32'hbf2a0ad3} /* (7, 0, 6) {real, imag} */,
  {32'hc067b81c, 32'hbe9d8e39} /* (7, 0, 5) {real, imag} */,
  {32'h4098350f, 32'h4081118b} /* (7, 0, 4) {real, imag} */,
  {32'h404db148, 32'h3fceeaa4} /* (7, 0, 3) {real, imag} */,
  {32'hbfc9992d, 32'hc0af316a} /* (7, 0, 2) {real, imag} */,
  {32'h40215e4a, 32'h3fd92793} /* (7, 0, 1) {real, imag} */,
  {32'hbe9f7d7b, 32'hc0c1131b} /* (7, 0, 0) {real, imag} */,
  {32'hc0890c3e, 32'hc00c9d5f} /* (6, 31, 31) {real, imag} */,
  {32'hbf913e86, 32'hc036d137} /* (6, 31, 30) {real, imag} */,
  {32'h41382502, 32'h3fd3efca} /* (6, 31, 29) {real, imag} */,
  {32'hbf9058a9, 32'h40bbe310} /* (6, 31, 28) {real, imag} */,
  {32'hbeb8a664, 32'h3f6f2b14} /* (6, 31, 27) {real, imag} */,
  {32'hbf261d28, 32'hc041b257} /* (6, 31, 26) {real, imag} */,
  {32'h404074f6, 32'h3fb1156b} /* (6, 31, 25) {real, imag} */,
  {32'hc02cbc29, 32'hc00163d0} /* (6, 31, 24) {real, imag} */,
  {32'h40222462, 32'hbdc9cc69} /* (6, 31, 23) {real, imag} */,
  {32'hc02424cf, 32'h3f75d9de} /* (6, 31, 22) {real, imag} */,
  {32'hbf85adaa, 32'h3fb20aa0} /* (6, 31, 21) {real, imag} */,
  {32'hbf01a688, 32'hc024e197} /* (6, 31, 20) {real, imag} */,
  {32'h402ea663, 32'h4044d3a3} /* (6, 31, 19) {real, imag} */,
  {32'h3e5f49ad, 32'h3e416d2a} /* (6, 31, 18) {real, imag} */,
  {32'hbebb3906, 32'hc0147820} /* (6, 31, 17) {real, imag} */,
  {32'hbdf554ac, 32'h3e92891c} /* (6, 31, 16) {real, imag} */,
  {32'h3f06d585, 32'hbe0debbe} /* (6, 31, 15) {real, imag} */,
  {32'h3f8ca5b0, 32'hbfabfd79} /* (6, 31, 14) {real, imag} */,
  {32'hbf6273a7, 32'h3f5f23dd} /* (6, 31, 13) {real, imag} */,
  {32'h405e2c8c, 32'h400d2ddd} /* (6, 31, 12) {real, imag} */,
  {32'hc031eeac, 32'h3de4d6c1} /* (6, 31, 11) {real, imag} */,
  {32'hbfda0198, 32'h3f08c799} /* (6, 31, 10) {real, imag} */,
  {32'h405c55c0, 32'h3ffc686a} /* (6, 31, 9) {real, imag} */,
  {32'h3f61a052, 32'hbf97bf82} /* (6, 31, 8) {real, imag} */,
  {32'hc0035216, 32'h4042491f} /* (6, 31, 7) {real, imag} */,
  {32'hc02cc300, 32'hc0666ca5} /* (6, 31, 6) {real, imag} */,
  {32'h3fb9ab28, 32'h4008ef1a} /* (6, 31, 5) {real, imag} */,
  {32'hc0acfb26, 32'h40f6dc31} /* (6, 31, 4) {real, imag} */,
  {32'h3f29b795, 32'hc1053939} /* (6, 31, 3) {real, imag} */,
  {32'h40f09af1, 32'h40bbb4a9} /* (6, 31, 2) {real, imag} */,
  {32'hbee9b043, 32'hbfe851d9} /* (6, 31, 1) {real, imag} */,
  {32'hc112c05e, 32'hbef71cae} /* (6, 31, 0) {real, imag} */,
  {32'h410ac75d, 32'h3fd4ec1e} /* (6, 30, 31) {real, imag} */,
  {32'h40b15230, 32'h3f8b6a49} /* (6, 30, 30) {real, imag} */,
  {32'h40a89385, 32'hbfa2fea4} /* (6, 30, 29) {real, imag} */,
  {32'hc02c1aaa, 32'h4066b20a} /* (6, 30, 28) {real, imag} */,
  {32'h3ee4e156, 32'hbf799317} /* (6, 30, 27) {real, imag} */,
  {32'hbff8d806, 32'hbf4e5b6f} /* (6, 30, 26) {real, imag} */,
  {32'hbe9604e8, 32'h3edb0737} /* (6, 30, 25) {real, imag} */,
  {32'h3dfd3081, 32'h4018b9de} /* (6, 30, 24) {real, imag} */,
  {32'hc052e9b1, 32'hbfaf5b92} /* (6, 30, 23) {real, imag} */,
  {32'hc01a7233, 32'h3c690f17} /* (6, 30, 22) {real, imag} */,
  {32'h3c7a18c9, 32'h3fa4a40e} /* (6, 30, 21) {real, imag} */,
  {32'hc0878c23, 32'h402d828f} /* (6, 30, 20) {real, imag} */,
  {32'h3ec40815, 32'hc017bce9} /* (6, 30, 19) {real, imag} */,
  {32'hbf62826c, 32'hbebb04c4} /* (6, 30, 18) {real, imag} */,
  {32'hbf84de0b, 32'hbed6a8a5} /* (6, 30, 17) {real, imag} */,
  {32'hbf0d0276, 32'hbed022df} /* (6, 30, 16) {real, imag} */,
  {32'hbfd83313, 32'h3f8000fa} /* (6, 30, 15) {real, imag} */,
  {32'hbca002e4, 32'hbe5e7e03} /* (6, 30, 14) {real, imag} */,
  {32'hbe2f8d37, 32'h3f437bba} /* (6, 30, 13) {real, imag} */,
  {32'h3ea4bb1a, 32'hc017cd78} /* (6, 30, 12) {real, imag} */,
  {32'h3f0ce1e2, 32'h3dd00cf7} /* (6, 30, 11) {real, imag} */,
  {32'hc0891cb5, 32'hbfe84ce9} /* (6, 30, 10) {real, imag} */,
  {32'h3f6acf5c, 32'h3c28fcd2} /* (6, 30, 9) {real, imag} */,
  {32'h3fd048f8, 32'h40298a85} /* (6, 30, 8) {real, imag} */,
  {32'h3eb1aeed, 32'hbeb6fe7b} /* (6, 30, 7) {real, imag} */,
  {32'h3f48b696, 32'hc0808286} /* (6, 30, 6) {real, imag} */,
  {32'hc0a33c7a, 32'h40934697} /* (6, 30, 5) {real, imag} */,
  {32'h3ffeab76, 32'hc0c06cc7} /* (6, 30, 4) {real, imag} */,
  {32'hc01db557, 32'h40da2d9c} /* (6, 30, 3) {real, imag} */,
  {32'h40d651aa, 32'hc107dc6a} /* (6, 30, 2) {real, imag} */,
  {32'hc0ba9cbf, 32'h4029c230} /* (6, 30, 1) {real, imag} */,
  {32'hc0738015, 32'hbfb7635f} /* (6, 30, 0) {real, imag} */,
  {32'hbf9454f0, 32'hc0e51da8} /* (6, 29, 31) {real, imag} */,
  {32'h401e6c9b, 32'h40aebf2b} /* (6, 29, 30) {real, imag} */,
  {32'h40b9a660, 32'h3f98d99d} /* (6, 29, 29) {real, imag} */,
  {32'hc0434c4d, 32'h3f9afad8} /* (6, 29, 28) {real, imag} */,
  {32'hbf001827, 32'hbff5124b} /* (6, 29, 27) {real, imag} */,
  {32'h3ed96380, 32'h40084fcc} /* (6, 29, 26) {real, imag} */,
  {32'hc03840cd, 32'h3c486142} /* (6, 29, 25) {real, imag} */,
  {32'hbf351a67, 32'h4014e206} /* (6, 29, 24) {real, imag} */,
  {32'hc055f41c, 32'hc0405bf8} /* (6, 29, 23) {real, imag} */,
  {32'hbf6208d2, 32'hbf9a1052} /* (6, 29, 22) {real, imag} */,
  {32'h4058d8a9, 32'hc07c653c} /* (6, 29, 21) {real, imag} */,
  {32'h3ea2291c, 32'h402461bd} /* (6, 29, 20) {real, imag} */,
  {32'h4055d242, 32'h3fb6c20f} /* (6, 29, 19) {real, imag} */,
  {32'h401bc0c1, 32'h3f2745d1} /* (6, 29, 18) {real, imag} */,
  {32'h3f9673f1, 32'hbf581255} /* (6, 29, 17) {real, imag} */,
  {32'h3f6657b6, 32'hbf344b98} /* (6, 29, 16) {real, imag} */,
  {32'h3f3bbe94, 32'h3f5b9b76} /* (6, 29, 15) {real, imag} */,
  {32'hbffbf68b, 32'h402901b6} /* (6, 29, 14) {real, imag} */,
  {32'hbfb456be, 32'h3f78a949} /* (6, 29, 13) {real, imag} */,
  {32'h403ce0e8, 32'h3f67c354} /* (6, 29, 12) {real, imag} */,
  {32'h3fabc9e5, 32'hc0828371} /* (6, 29, 11) {real, imag} */,
  {32'hbfd2946c, 32'h3e812f16} /* (6, 29, 10) {real, imag} */,
  {32'h3f36b948, 32'hbfc0772a} /* (6, 29, 9) {real, imag} */,
  {32'h40a79437, 32'h3ee8172e} /* (6, 29, 8) {real, imag} */,
  {32'h3fb0290b, 32'hbfa1b565} /* (6, 29, 7) {real, imag} */,
  {32'h3f709778, 32'h3fd681c6} /* (6, 29, 6) {real, imag} */,
  {32'hc01b69dc, 32'hc0a82bd9} /* (6, 29, 5) {real, imag} */,
  {32'hc03d4aca, 32'hbec1944f} /* (6, 29, 4) {real, imag} */,
  {32'h4001e697, 32'h40afb0e1} /* (6, 29, 3) {real, imag} */,
  {32'hc022b852, 32'h40dfdcd3} /* (6, 29, 2) {real, imag} */,
  {32'h401b7bc4, 32'h3eca723c} /* (6, 29, 1) {real, imag} */,
  {32'h40e2155e, 32'hc12fc090} /* (6, 29, 0) {real, imag} */,
  {32'hc06e67b9, 32'hc0868ee7} /* (6, 28, 31) {real, imag} */,
  {32'hc0ba8a74, 32'h3f012ec4} /* (6, 28, 30) {real, imag} */,
  {32'h40d347eb, 32'hc08541d7} /* (6, 28, 29) {real, imag} */,
  {32'h3f626f31, 32'hc034ec67} /* (6, 28, 28) {real, imag} */,
  {32'h4077529e, 32'h40265fbf} /* (6, 28, 27) {real, imag} */,
  {32'hc09fcf94, 32'h3f33f96e} /* (6, 28, 26) {real, imag} */,
  {32'h401ed6ed, 32'h4014be2c} /* (6, 28, 25) {real, imag} */,
  {32'h40549c5e, 32'hbf40ce57} /* (6, 28, 24) {real, imag} */,
  {32'hbf044f67, 32'hbf83aff5} /* (6, 28, 23) {real, imag} */,
  {32'h3e40b5f3, 32'h3f4596f1} /* (6, 28, 22) {real, imag} */,
  {32'hbeaa11a7, 32'h3fded89e} /* (6, 28, 21) {real, imag} */,
  {32'h3ffdc406, 32'hbf86ba46} /* (6, 28, 20) {real, imag} */,
  {32'hc05b30cf, 32'h3face9bf} /* (6, 28, 19) {real, imag} */,
  {32'h3f066a41, 32'hbeb30d74} /* (6, 28, 18) {real, imag} */,
  {32'hbfd23211, 32'hc021431c} /* (6, 28, 17) {real, imag} */,
  {32'hbf36a517, 32'hbf82e1f2} /* (6, 28, 16) {real, imag} */,
  {32'h3fd02a02, 32'hbea72367} /* (6, 28, 15) {real, imag} */,
  {32'h3fd0a438, 32'hbea60d62} /* (6, 28, 14) {real, imag} */,
  {32'hbfdc5b77, 32'hc0914cb2} /* (6, 28, 13) {real, imag} */,
  {32'h402ef3a7, 32'hc0596042} /* (6, 28, 12) {real, imag} */,
  {32'hc02638d0, 32'h40117072} /* (6, 28, 11) {real, imag} */,
  {32'h3f09c873, 32'h3ffae799} /* (6, 28, 10) {real, imag} */,
  {32'h3f535b1a, 32'h3fe70b42} /* (6, 28, 9) {real, imag} */,
  {32'h4020486b, 32'h3ed47f04} /* (6, 28, 8) {real, imag} */,
  {32'h40b3868f, 32'hbf85b8f8} /* (6, 28, 7) {real, imag} */,
  {32'hbfb30897, 32'hc0b5c00a} /* (6, 28, 6) {real, imag} */,
  {32'h3bda0664, 32'hc0530912} /* (6, 28, 5) {real, imag} */,
  {32'h4053777a, 32'h3ffbf9e4} /* (6, 28, 4) {real, imag} */,
  {32'h408f1c6c, 32'h3fe20139} /* (6, 28, 3) {real, imag} */,
  {32'h40a1d87e, 32'h407236a8} /* (6, 28, 2) {real, imag} */,
  {32'hc07e77d3, 32'h3fd00d29} /* (6, 28, 1) {real, imag} */,
  {32'h3f37aa4c, 32'h3f173cee} /* (6, 28, 0) {real, imag} */,
  {32'hbf6ef52d, 32'h40015d19} /* (6, 27, 31) {real, imag} */,
  {32'h409d49e0, 32'hc022b966} /* (6, 27, 30) {real, imag} */,
  {32'hbeb7180a, 32'h3ffc4edb} /* (6, 27, 29) {real, imag} */,
  {32'hc08443cd, 32'hbf4cd1c0} /* (6, 27, 28) {real, imag} */,
  {32'hbfa23f54, 32'h3e0533d9} /* (6, 27, 27) {real, imag} */,
  {32'h3e8f34e1, 32'h3ec368d2} /* (6, 27, 26) {real, imag} */,
  {32'hc0400107, 32'h3f7dd6bc} /* (6, 27, 25) {real, imag} */,
  {32'h40401b54, 32'hc0316028} /* (6, 27, 24) {real, imag} */,
  {32'h3d7939d4, 32'h3e5e9dd1} /* (6, 27, 23) {real, imag} */,
  {32'h40389e5d, 32'h3fb2d19e} /* (6, 27, 22) {real, imag} */,
  {32'hbdc91340, 32'hbec19f91} /* (6, 27, 21) {real, imag} */,
  {32'h3fb997d7, 32'hbf844677} /* (6, 27, 20) {real, imag} */,
  {32'h3fb9b661, 32'hc07d0247} /* (6, 27, 19) {real, imag} */,
  {32'h3f1dc045, 32'h3f93c006} /* (6, 27, 18) {real, imag} */,
  {32'hbe1db2ab, 32'h3e72821c} /* (6, 27, 17) {real, imag} */,
  {32'hbf810d47, 32'hbfc71d3d} /* (6, 27, 16) {real, imag} */,
  {32'hbf2523d3, 32'h3f9742c8} /* (6, 27, 15) {real, imag} */,
  {32'h3e5d6c82, 32'h3f9cbac6} /* (6, 27, 14) {real, imag} */,
  {32'hbfbb0383, 32'hbf907eeb} /* (6, 27, 13) {real, imag} */,
  {32'h40955986, 32'h3fd4b328} /* (6, 27, 12) {real, imag} */,
  {32'h3fcc51cc, 32'h3f57b106} /* (6, 27, 11) {real, imag} */,
  {32'hc04b7dc0, 32'h3f736c29} /* (6, 27, 10) {real, imag} */,
  {32'h3f0045d0, 32'hc015d09b} /* (6, 27, 9) {real, imag} */,
  {32'hbea036cc, 32'hc023123b} /* (6, 27, 8) {real, imag} */,
  {32'h3fdf2eaa, 32'h3e48e60c} /* (6, 27, 7) {real, imag} */,
  {32'h3eb8c134, 32'h3e9735b3} /* (6, 27, 6) {real, imag} */,
  {32'h3e79dd38, 32'hc0a0714f} /* (6, 27, 5) {real, imag} */,
  {32'hc00edfc0, 32'hbf6a1740} /* (6, 27, 4) {real, imag} */,
  {32'hbfb3ae66, 32'h3f843f04} /* (6, 27, 3) {real, imag} */,
  {32'h3f6e1b5a, 32'h3e5ab591} /* (6, 27, 2) {real, imag} */,
  {32'hc041f344, 32'hc014fcb7} /* (6, 27, 1) {real, imag} */,
  {32'h3de67127, 32'hc079fc0a} /* (6, 27, 0) {real, imag} */,
  {32'h407fd40c, 32'hc0638119} /* (6, 26, 31) {real, imag} */,
  {32'hbf0cd021, 32'h3f657d6a} /* (6, 26, 30) {real, imag} */,
  {32'hbf74c9ad, 32'h407d73ba} /* (6, 26, 29) {real, imag} */,
  {32'hbeae2ceb, 32'hc07267fd} /* (6, 26, 28) {real, imag} */,
  {32'hbf512d37, 32'hbe9a2e06} /* (6, 26, 27) {real, imag} */,
  {32'h3f2ea376, 32'h3fa68235} /* (6, 26, 26) {real, imag} */,
  {32'h400c246d, 32'hbf83a9ef} /* (6, 26, 25) {real, imag} */,
  {32'h3e9c08aa, 32'h4080c27a} /* (6, 26, 24) {real, imag} */,
  {32'h401a09d1, 32'h40184347} /* (6, 26, 23) {real, imag} */,
  {32'hc025a35b, 32'h3e779edb} /* (6, 26, 22) {real, imag} */,
  {32'hbe98ff5f, 32'hbf3f18db} /* (6, 26, 21) {real, imag} */,
  {32'h3f51c390, 32'hbf8dfd1e} /* (6, 26, 20) {real, imag} */,
  {32'hbfe51150, 32'h408681b4} /* (6, 26, 19) {real, imag} */,
  {32'h3f38befd, 32'hbece0efa} /* (6, 26, 18) {real, imag} */,
  {32'hbec67627, 32'h3f89ad34} /* (6, 26, 17) {real, imag} */,
  {32'h3fb1222c, 32'hbcccc8db} /* (6, 26, 16) {real, imag} */,
  {32'hbf334d4c, 32'hbd1d3416} /* (6, 26, 15) {real, imag} */,
  {32'h3e2db08c, 32'hbfb1ade7} /* (6, 26, 14) {real, imag} */,
  {32'hc01b84ee, 32'hbfa0909b} /* (6, 26, 13) {real, imag} */,
  {32'h3f15ae96, 32'hbf5e6dc9} /* (6, 26, 12) {real, imag} */,
  {32'h3fe46e25, 32'h3f2d2557} /* (6, 26, 11) {real, imag} */,
  {32'hbff9459b, 32'hbf3452e9} /* (6, 26, 10) {real, imag} */,
  {32'h3da34456, 32'h3e282ce2} /* (6, 26, 9) {real, imag} */,
  {32'hbfbe5913, 32'hbf4227f8} /* (6, 26, 8) {real, imag} */,
  {32'hbfe90737, 32'hc0a0847b} /* (6, 26, 7) {real, imag} */,
  {32'h4082fd32, 32'h402d521c} /* (6, 26, 6) {real, imag} */,
  {32'h401e87aa, 32'h3e95b78d} /* (6, 26, 5) {real, imag} */,
  {32'h3fa0d772, 32'h407bbac4} /* (6, 26, 4) {real, imag} */,
  {32'h40bf994b, 32'hbd90861b} /* (6, 26, 3) {real, imag} */,
  {32'hc053b6dd, 32'h3e8e9dc6} /* (6, 26, 2) {real, imag} */,
  {32'h4012668f, 32'hbf9f6f37} /* (6, 26, 1) {real, imag} */,
  {32'h3f7bb9c8, 32'h40b5e67e} /* (6, 26, 0) {real, imag} */,
  {32'h4045a726, 32'hc0602031} /* (6, 25, 31) {real, imag} */,
  {32'hbebe0d19, 32'h3f7480b4} /* (6, 25, 30) {real, imag} */,
  {32'h3e0871a2, 32'h40bccca5} /* (6, 25, 29) {real, imag} */,
  {32'h3f52f834, 32'h3eb1e40b} /* (6, 25, 28) {real, imag} */,
  {32'h3f4486d6, 32'h3eeebb07} /* (6, 25, 27) {real, imag} */,
  {32'hbf8b2221, 32'hc041ba8d} /* (6, 25, 26) {real, imag} */,
  {32'hbea862c4, 32'hc01958cb} /* (6, 25, 25) {real, imag} */,
  {32'h3f798c15, 32'h403b54ca} /* (6, 25, 24) {real, imag} */,
  {32'hbf168e53, 32'h3f09e990} /* (6, 25, 23) {real, imag} */,
  {32'hbffd035f, 32'h3ee137d8} /* (6, 25, 22) {real, imag} */,
  {32'h3ff73552, 32'h3f7ad227} /* (6, 25, 21) {real, imag} */,
  {32'h3f5666d1, 32'hbd1b18f0} /* (6, 25, 20) {real, imag} */,
  {32'hbf3dd29c, 32'hbe388f19} /* (6, 25, 19) {real, imag} */,
  {32'hbdb19a6f, 32'hc0330e6d} /* (6, 25, 18) {real, imag} */,
  {32'hbea016c8, 32'hc0478830} /* (6, 25, 17) {real, imag} */,
  {32'hbfb0151c, 32'h3fb39029} /* (6, 25, 16) {real, imag} */,
  {32'h3f5a7ac4, 32'h3fc038d6} /* (6, 25, 15) {real, imag} */,
  {32'hc00d2086, 32'h3fd42523} /* (6, 25, 14) {real, imag} */,
  {32'hbee93d12, 32'hc00980f9} /* (6, 25, 13) {real, imag} */,
  {32'hbfe46db5, 32'h3d929421} /* (6, 25, 12) {real, imag} */,
  {32'h401ccabe, 32'hc046ed68} /* (6, 25, 11) {real, imag} */,
  {32'hbeaa2038, 32'h3fea8e85} /* (6, 25, 10) {real, imag} */,
  {32'h3efda3c1, 32'hbe0ea315} /* (6, 25, 9) {real, imag} */,
  {32'hc07deed9, 32'hbf4e598a} /* (6, 25, 8) {real, imag} */,
  {32'h3f85363c, 32'h3f8b8b2a} /* (6, 25, 7) {real, imag} */,
  {32'hbfa2af1e, 32'hbff0162f} /* (6, 25, 6) {real, imag} */,
  {32'h3e973b18, 32'h40345d9e} /* (6, 25, 5) {real, imag} */,
  {32'hc033060b, 32'hc02a7e9c} /* (6, 25, 4) {real, imag} */,
  {32'h3d275fd6, 32'hbfd15348} /* (6, 25, 3) {real, imag} */,
  {32'hbfc6efe9, 32'hbf1144a0} /* (6, 25, 2) {real, imag} */,
  {32'h4027f683, 32'hc07608ee} /* (6, 25, 1) {real, imag} */,
  {32'hbfd8c48a, 32'hc03cca96} /* (6, 25, 0) {real, imag} */,
  {32'hc0096f50, 32'h3fc23a5a} /* (6, 24, 31) {real, imag} */,
  {32'h402373d0, 32'hc0d1d23a} /* (6, 24, 30) {real, imag} */,
  {32'hbdd25c3e, 32'hc034d3d1} /* (6, 24, 29) {real, imag} */,
  {32'h401d8a31, 32'hbf6df5a4} /* (6, 24, 28) {real, imag} */,
  {32'hbfc31a28, 32'h3ed2055a} /* (6, 24, 27) {real, imag} */,
  {32'h3f1f4db1, 32'hbe955dc6} /* (6, 24, 26) {real, imag} */,
  {32'h408fa381, 32'h3f89addc} /* (6, 24, 25) {real, imag} */,
  {32'h3f81c9c4, 32'h3fab381c} /* (6, 24, 24) {real, imag} */,
  {32'h403fbe8c, 32'hbfcccaeb} /* (6, 24, 23) {real, imag} */,
  {32'hbf574be2, 32'hc053d54a} /* (6, 24, 22) {real, imag} */,
  {32'hbfb83cc4, 32'hc01a48e8} /* (6, 24, 21) {real, imag} */,
  {32'hbf62ea5c, 32'hbfa8f3a8} /* (6, 24, 20) {real, imag} */,
  {32'hc01bf957, 32'h3ff54035} /* (6, 24, 19) {real, imag} */,
  {32'h4022367a, 32'hbfccff81} /* (6, 24, 18) {real, imag} */,
  {32'hbf958a85, 32'hbfe752da} /* (6, 24, 17) {real, imag} */,
  {32'hbf8a5fc4, 32'h3fe1f0bd} /* (6, 24, 16) {real, imag} */,
  {32'h3e99dfcd, 32'h3f66cbaa} /* (6, 24, 15) {real, imag} */,
  {32'h3f261578, 32'hc0392448} /* (6, 24, 14) {real, imag} */,
  {32'hbf00c181, 32'h3f975ffe} /* (6, 24, 13) {real, imag} */,
  {32'h400e415c, 32'hbf86c9c9} /* (6, 24, 12) {real, imag} */,
  {32'hbffee716, 32'hc04139a2} /* (6, 24, 11) {real, imag} */,
  {32'h3fe70ff9, 32'h3fe9ae72} /* (6, 24, 10) {real, imag} */,
  {32'h3f23844b, 32'hbf993ecc} /* (6, 24, 9) {real, imag} */,
  {32'hc078ac17, 32'hbdb88990} /* (6, 24, 8) {real, imag} */,
  {32'h3ed166e2, 32'h3de0e576} /* (6, 24, 7) {real, imag} */,
  {32'hc026e30e, 32'hc06d2f8c} /* (6, 24, 6) {real, imag} */,
  {32'hbf1906b4, 32'h3e69efba} /* (6, 24, 5) {real, imag} */,
  {32'h3f848552, 32'h4004789d} /* (6, 24, 4) {real, imag} */,
  {32'hbe864b22, 32'hc04cd06a} /* (6, 24, 3) {real, imag} */,
  {32'hc095a5b9, 32'h40b53167} /* (6, 24, 2) {real, imag} */,
  {32'hbf8869c0, 32'hbf071898} /* (6, 24, 1) {real, imag} */,
  {32'h407f328e, 32'h3faf2abb} /* (6, 24, 0) {real, imag} */,
  {32'h3f239512, 32'hbf1431b0} /* (6, 23, 31) {real, imag} */,
  {32'h3ff5dcb1, 32'hbf93d682} /* (6, 23, 30) {real, imag} */,
  {32'h400684b4, 32'hbf0ed66a} /* (6, 23, 29) {real, imag} */,
  {32'h3f886811, 32'hbf9a6cf2} /* (6, 23, 28) {real, imag} */,
  {32'h3f2c97a3, 32'hbf44e224} /* (6, 23, 27) {real, imag} */,
  {32'h3e328e84, 32'h403e0b6e} /* (6, 23, 26) {real, imag} */,
  {32'h4027aea4, 32'hbe293302} /* (6, 23, 25) {real, imag} */,
  {32'hbf0962c6, 32'hbfbc6d64} /* (6, 23, 24) {real, imag} */,
  {32'h40803e4d, 32'h3f499bfb} /* (6, 23, 23) {real, imag} */,
  {32'hbf7055cd, 32'h4049c947} /* (6, 23, 22) {real, imag} */,
  {32'h3f80c8b6, 32'h4028c41a} /* (6, 23, 21) {real, imag} */,
  {32'hbfd1e4a7, 32'hbf21a59a} /* (6, 23, 20) {real, imag} */,
  {32'hbe8cf9b4, 32'hbf8fda35} /* (6, 23, 19) {real, imag} */,
  {32'h3fd7ce5b, 32'h3fbbecc9} /* (6, 23, 18) {real, imag} */,
  {32'hbfc50b5b, 32'hbf23a92a} /* (6, 23, 17) {real, imag} */,
  {32'hc02e4054, 32'hc02143eb} /* (6, 23, 16) {real, imag} */,
  {32'hbf8d9d1e, 32'hbf2702f6} /* (6, 23, 15) {real, imag} */,
  {32'hbf9f7053, 32'hc0608809} /* (6, 23, 14) {real, imag} */,
  {32'hbf38dd39, 32'h3f552b4c} /* (6, 23, 13) {real, imag} */,
  {32'h3feb4767, 32'hbfd7dfd5} /* (6, 23, 12) {real, imag} */,
  {32'h3f529885, 32'h404050e4} /* (6, 23, 11) {real, imag} */,
  {32'h3fbab614, 32'hc0480109} /* (6, 23, 10) {real, imag} */,
  {32'hbf12af5a, 32'hbfdea230} /* (6, 23, 9) {real, imag} */,
  {32'hc0000a3f, 32'h3edbf650} /* (6, 23, 8) {real, imag} */,
  {32'h3e756695, 32'h4003afb6} /* (6, 23, 7) {real, imag} */,
  {32'h3fce6dd5, 32'hbf26e700} /* (6, 23, 6) {real, imag} */,
  {32'h3fc753bf, 32'h404d25db} /* (6, 23, 5) {real, imag} */,
  {32'hc0136ac7, 32'h3f8f1f33} /* (6, 23, 4) {real, imag} */,
  {32'hbd937977, 32'h401adf6c} /* (6, 23, 3) {real, imag} */,
  {32'hbe1915bc, 32'hc067b636} /* (6, 23, 2) {real, imag} */,
  {32'h3ee28613, 32'h3f087f8c} /* (6, 23, 1) {real, imag} */,
  {32'h3ff85cd1, 32'hbfd4b9ea} /* (6, 23, 0) {real, imag} */,
  {32'h3badb1f8, 32'hbe8c3066} /* (6, 22, 31) {real, imag} */,
  {32'hbf4d1a99, 32'h3f7538be} /* (6, 22, 30) {real, imag} */,
  {32'h40367e17, 32'h4008ba84} /* (6, 22, 29) {real, imag} */,
  {32'hbf6943a7, 32'hc04a5ae7} /* (6, 22, 28) {real, imag} */,
  {32'h3f4694b8, 32'hbdd5e9ca} /* (6, 22, 27) {real, imag} */,
  {32'h40716def, 32'hbf4953f4} /* (6, 22, 26) {real, imag} */,
  {32'hbcf63948, 32'hbf754171} /* (6, 22, 25) {real, imag} */,
  {32'h400b0f64, 32'h40739fb8} /* (6, 22, 24) {real, imag} */,
  {32'hbeda8626, 32'hbfb9d406} /* (6, 22, 23) {real, imag} */,
  {32'hbfd56ea7, 32'hbf956477} /* (6, 22, 22) {real, imag} */,
  {32'hbf88875d, 32'h3f4292f7} /* (6, 22, 21) {real, imag} */,
  {32'h3f750440, 32'hbea9bfd9} /* (6, 22, 20) {real, imag} */,
  {32'hbf9a949f, 32'hbe4876b5} /* (6, 22, 19) {real, imag} */,
  {32'h3f2341e0, 32'h3fe6a8ba} /* (6, 22, 18) {real, imag} */,
  {32'hbe1ea961, 32'h3ea09db2} /* (6, 22, 17) {real, imag} */,
  {32'h4020a0ac, 32'h3f2f3994} /* (6, 22, 16) {real, imag} */,
  {32'hbd9654fe, 32'hc07163ec} /* (6, 22, 15) {real, imag} */,
  {32'h3f3863dc, 32'hbf336661} /* (6, 22, 14) {real, imag} */,
  {32'hbfad5b9d, 32'hbedc2110} /* (6, 22, 13) {real, imag} */,
  {32'h3fcd4c26, 32'hbe6a4486} /* (6, 22, 12) {real, imag} */,
  {32'hbf54d6b7, 32'hbe12720f} /* (6, 22, 11) {real, imag} */,
  {32'h3f0355dd, 32'h40540987} /* (6, 22, 10) {real, imag} */,
  {32'h3fbdd49b, 32'h3eefce2e} /* (6, 22, 9) {real, imag} */,
  {32'h40a1f8cd, 32'hbff049d1} /* (6, 22, 8) {real, imag} */,
  {32'hbfdde9d8, 32'h4000d3ac} /* (6, 22, 7) {real, imag} */,
  {32'hbeddbd5c, 32'hc0886e28} /* (6, 22, 6) {real, imag} */,
  {32'hbf93bbce, 32'h405b1249} /* (6, 22, 5) {real, imag} */,
  {32'hbe830664, 32'h3f3c6f5f} /* (6, 22, 4) {real, imag} */,
  {32'h4060e267, 32'h3df5a5e9} /* (6, 22, 3) {real, imag} */,
  {32'hc001c3de, 32'h3f7d26af} /* (6, 22, 2) {real, imag} */,
  {32'hbf0d93fd, 32'h3f98ab3e} /* (6, 22, 1) {real, imag} */,
  {32'hc01f3402, 32'hbfad6705} /* (6, 22, 0) {real, imag} */,
  {32'h3fac1e4d, 32'h3fc3bcaf} /* (6, 21, 31) {real, imag} */,
  {32'hbf430dea, 32'hbf01dec6} /* (6, 21, 30) {real, imag} */,
  {32'hc0542366, 32'h3f28de7a} /* (6, 21, 29) {real, imag} */,
  {32'h3f46f33d, 32'hc0469c0e} /* (6, 21, 28) {real, imag} */,
  {32'hbec700ce, 32'hbecf952d} /* (6, 21, 27) {real, imag} */,
  {32'hc0124191, 32'h3faf9aaa} /* (6, 21, 26) {real, imag} */,
  {32'h3e114a99, 32'h3fbe15a4} /* (6, 21, 25) {real, imag} */,
  {32'h3f94a603, 32'hc0157fcb} /* (6, 21, 24) {real, imag} */,
  {32'h3fa5731c, 32'hc095ddce} /* (6, 21, 23) {real, imag} */,
  {32'hbf648dc7, 32'h3f62ed24} /* (6, 21, 22) {real, imag} */,
  {32'hbfc9cd18, 32'h3ff3fa22} /* (6, 21, 21) {real, imag} */,
  {32'hbef7b444, 32'hc005ad85} /* (6, 21, 20) {real, imag} */,
  {32'hbfe83507, 32'hc04e0f68} /* (6, 21, 19) {real, imag} */,
  {32'h3f49e1b2, 32'h3dbfcedd} /* (6, 21, 18) {real, imag} */,
  {32'hbf6a35d3, 32'h40372cbe} /* (6, 21, 17) {real, imag} */,
  {32'hbf145e60, 32'hbfa853ee} /* (6, 21, 16) {real, imag} */,
  {32'h3f98d877, 32'h3f4348c0} /* (6, 21, 15) {real, imag} */,
  {32'hbf837a57, 32'h3fea750e} /* (6, 21, 14) {real, imag} */,
  {32'h3e9bdb81, 32'hc03db982} /* (6, 21, 13) {real, imag} */,
  {32'hc031df7a, 32'hc0129383} /* (6, 21, 12) {real, imag} */,
  {32'hbfb03abc, 32'h3fb8c295} /* (6, 21, 11) {real, imag} */,
  {32'h3ec40b2f, 32'hbf5a5371} /* (6, 21, 10) {real, imag} */,
  {32'h3f260b2b, 32'h3fdc5d6d} /* (6, 21, 9) {real, imag} */,
  {32'h3fd5816e, 32'h3eed123c} /* (6, 21, 8) {real, imag} */,
  {32'hbfea71ca, 32'hc01f788f} /* (6, 21, 7) {real, imag} */,
  {32'hbfa97466, 32'h3ea0b213} /* (6, 21, 6) {real, imag} */,
  {32'hc02a5ef7, 32'h3e259fa9} /* (6, 21, 5) {real, imag} */,
  {32'hbf9b2463, 32'hc0117b88} /* (6, 21, 4) {real, imag} */,
  {32'h3febaf6b, 32'hbf45c435} /* (6, 21, 3) {real, imag} */,
  {32'h405766be, 32'hbf76d3c1} /* (6, 21, 2) {real, imag} */,
  {32'hc0504d15, 32'h3f699093} /* (6, 21, 1) {real, imag} */,
  {32'h3fbc6fcb, 32'hbe9b7369} /* (6, 21, 0) {real, imag} */,
  {32'hbff2083c, 32'h3f882801} /* (6, 20, 31) {real, imag} */,
  {32'h4037584a, 32'h400c50b3} /* (6, 20, 30) {real, imag} */,
  {32'hbe265477, 32'hc000b218} /* (6, 20, 29) {real, imag} */,
  {32'hbead4053, 32'hbf7c74ac} /* (6, 20, 28) {real, imag} */,
  {32'hbe261fbd, 32'h3fc81b52} /* (6, 20, 27) {real, imag} */,
  {32'h3f1fddd5, 32'hbe9b97d1} /* (6, 20, 26) {real, imag} */,
  {32'h3d41d6ca, 32'h3f1fa7fc} /* (6, 20, 25) {real, imag} */,
  {32'h3ffaffac, 32'hc07b025b} /* (6, 20, 24) {real, imag} */,
  {32'hbfe52051, 32'h3fc61a3c} /* (6, 20, 23) {real, imag} */,
  {32'h3fe7de0c, 32'hc0285933} /* (6, 20, 22) {real, imag} */,
  {32'hbfb53590, 32'hbfb03673} /* (6, 20, 21) {real, imag} */,
  {32'h4022e10d, 32'h3eeb1bcb} /* (6, 20, 20) {real, imag} */,
  {32'h3f51acfb, 32'hbf8a2f8c} /* (6, 20, 19) {real, imag} */,
  {32'hbecaf370, 32'h40477a9b} /* (6, 20, 18) {real, imag} */,
  {32'hbd506d93, 32'h3e961172} /* (6, 20, 17) {real, imag} */,
  {32'hbf45f626, 32'h4017fc8b} /* (6, 20, 16) {real, imag} */,
  {32'h3f9da5e2, 32'h40201a49} /* (6, 20, 15) {real, imag} */,
  {32'hbddb1dda, 32'h3f952fc6} /* (6, 20, 14) {real, imag} */,
  {32'h4020e3fb, 32'hbf1444f3} /* (6, 20, 13) {real, imag} */,
  {32'hbff79a8c, 32'hbfb28dda} /* (6, 20, 12) {real, imag} */,
  {32'h40154f6e, 32'h3fff1eeb} /* (6, 20, 11) {real, imag} */,
  {32'h3fb3be00, 32'hbf9b6703} /* (6, 20, 10) {real, imag} */,
  {32'h3fb38ddb, 32'hbfc51eba} /* (6, 20, 9) {real, imag} */,
  {32'hc01877bf, 32'h3f3c385d} /* (6, 20, 8) {real, imag} */,
  {32'h3d825cce, 32'hbf8f5a4a} /* (6, 20, 7) {real, imag} */,
  {32'hc008aa14, 32'h3f91df3a} /* (6, 20, 6) {real, imag} */,
  {32'hbf82dd7b, 32'hc002f799} /* (6, 20, 5) {real, imag} */,
  {32'hbfdf0616, 32'h4001c05f} /* (6, 20, 4) {real, imag} */,
  {32'hbfddfd54, 32'h3fc2ffdd} /* (6, 20, 3) {real, imag} */,
  {32'h3f9ce3b0, 32'h3e981c9e} /* (6, 20, 2) {real, imag} */,
  {32'h3eeb8d7b, 32'hbf7df4f2} /* (6, 20, 1) {real, imag} */,
  {32'h3f1eb140, 32'h3fdce5da} /* (6, 20, 0) {real, imag} */,
  {32'hbf7c1efb, 32'h403c92b5} /* (6, 19, 31) {real, imag} */,
  {32'h3ed1cfe3, 32'hbfe88c4f} /* (6, 19, 30) {real, imag} */,
  {32'hbf8cbee6, 32'h3f3f4fcd} /* (6, 19, 29) {real, imag} */,
  {32'hbf9438be, 32'hbfb000d8} /* (6, 19, 28) {real, imag} */,
  {32'hbe8e7f84, 32'hbe1091c4} /* (6, 19, 27) {real, imag} */,
  {32'hbfbb4055, 32'h3f42ea02} /* (6, 19, 26) {real, imag} */,
  {32'hc05b2eab, 32'hbf03ac26} /* (6, 19, 25) {real, imag} */,
  {32'h4004a7c4, 32'hbf428274} /* (6, 19, 24) {real, imag} */,
  {32'hbfd5eb4f, 32'h3e8def72} /* (6, 19, 23) {real, imag} */,
  {32'hbefe5eb5, 32'h3fa3afcb} /* (6, 19, 22) {real, imag} */,
  {32'h3e89e04f, 32'hbfebc93a} /* (6, 19, 21) {real, imag} */,
  {32'h3ea3cff3, 32'hc0039d5c} /* (6, 19, 20) {real, imag} */,
  {32'h3fbe0ebf, 32'hc0150fe5} /* (6, 19, 19) {real, imag} */,
  {32'hbe1c8b0d, 32'h3fdb2093} /* (6, 19, 18) {real, imag} */,
  {32'h3f8cdc49, 32'h3f0499d8} /* (6, 19, 17) {real, imag} */,
  {32'h3e52b36e, 32'h3e5718ef} /* (6, 19, 16) {real, imag} */,
  {32'hc007c12f, 32'hbf8b1e37} /* (6, 19, 15) {real, imag} */,
  {32'hbf94ee72, 32'hc023de1e} /* (6, 19, 14) {real, imag} */,
  {32'hbfad80f7, 32'hbf118369} /* (6, 19, 13) {real, imag} */,
  {32'hc0458014, 32'hbd191575} /* (6, 19, 12) {real, imag} */,
  {32'hbf315308, 32'h3fdc900b} /* (6, 19, 11) {real, imag} */,
  {32'h402233c9, 32'hbfa6798a} /* (6, 19, 10) {real, imag} */,
  {32'h40594f19, 32'hbf8b6966} /* (6, 19, 9) {real, imag} */,
  {32'h3f378d9b, 32'h3f694958} /* (6, 19, 8) {real, imag} */,
  {32'hbf68c4d4, 32'hbeeb61bc} /* (6, 19, 7) {real, imag} */,
  {32'hbfc31db9, 32'h3f368514} /* (6, 19, 6) {real, imag} */,
  {32'h3fbe167c, 32'hbf6d150b} /* (6, 19, 5) {real, imag} */,
  {32'hbe89f65c, 32'hbfbff52f} /* (6, 19, 4) {real, imag} */,
  {32'hbfb9439c, 32'h3df3b881} /* (6, 19, 3) {real, imag} */,
  {32'h3f994a12, 32'h3facb539} /* (6, 19, 2) {real, imag} */,
  {32'hbf3da694, 32'h3c9e55a3} /* (6, 19, 1) {real, imag} */,
  {32'hbec3cee4, 32'hbfb5a5bb} /* (6, 19, 0) {real, imag} */,
  {32'hc016bc65, 32'hbf24580e} /* (6, 18, 31) {real, imag} */,
  {32'hbef06cb3, 32'h3ea1860f} /* (6, 18, 30) {real, imag} */,
  {32'h3fd6cb8b, 32'h402c5662} /* (6, 18, 29) {real, imag} */,
  {32'hbfe038f8, 32'h3fcae717} /* (6, 18, 28) {real, imag} */,
  {32'hbd4e43fd, 32'h3edb85ca} /* (6, 18, 27) {real, imag} */,
  {32'hbfea2f11, 32'hbfd49f8d} /* (6, 18, 26) {real, imag} */,
  {32'h3e823620, 32'h3f5e191a} /* (6, 18, 25) {real, imag} */,
  {32'h3e667988, 32'h3f221834} /* (6, 18, 24) {real, imag} */,
  {32'hc0418428, 32'hbe785146} /* (6, 18, 23) {real, imag} */,
  {32'h3f4184eb, 32'hbf589325} /* (6, 18, 22) {real, imag} */,
  {32'hbf751d56, 32'h3f874a55} /* (6, 18, 21) {real, imag} */,
  {32'hbf3072df, 32'hbff79f13} /* (6, 18, 20) {real, imag} */,
  {32'h3f3d53f5, 32'hbfd908a5} /* (6, 18, 19) {real, imag} */,
  {32'hc0380554, 32'hbdc6889f} /* (6, 18, 18) {real, imag} */,
  {32'hbf8038a0, 32'hbe927024} /* (6, 18, 17) {real, imag} */,
  {32'hbf168a00, 32'h3e8c3c4a} /* (6, 18, 16) {real, imag} */,
  {32'hc012f959, 32'h3e1ca029} /* (6, 18, 15) {real, imag} */,
  {32'h3f92d421, 32'h3ff79839} /* (6, 18, 14) {real, imag} */,
  {32'h3ec39bca, 32'hbf3a903e} /* (6, 18, 13) {real, imag} */,
  {32'hbe8bfcd2, 32'hbf1892a1} /* (6, 18, 12) {real, imag} */,
  {32'h3f5dd10c, 32'h3e4fb6ef} /* (6, 18, 11) {real, imag} */,
  {32'hc002c641, 32'h4030c47c} /* (6, 18, 10) {real, imag} */,
  {32'hbeccdaf9, 32'h3fd5014c} /* (6, 18, 9) {real, imag} */,
  {32'h3c859e7c, 32'h3fcb151f} /* (6, 18, 8) {real, imag} */,
  {32'h402e623d, 32'h3f6587ef} /* (6, 18, 7) {real, imag} */,
  {32'h400fed4f, 32'h3fe8e88d} /* (6, 18, 6) {real, imag} */,
  {32'hbdd0a57f, 32'h3f6b59b7} /* (6, 18, 5) {real, imag} */,
  {32'hc04bc63a, 32'h3edd9599} /* (6, 18, 4) {real, imag} */,
  {32'h3f5c2e80, 32'hc044a5aa} /* (6, 18, 3) {real, imag} */,
  {32'hbf042e7c, 32'h3eb00279} /* (6, 18, 2) {real, imag} */,
  {32'h3e9fd9d4, 32'h3fcc7d70} /* (6, 18, 1) {real, imag} */,
  {32'h3de8868e, 32'hbf411ca4} /* (6, 18, 0) {real, imag} */,
  {32'h3f2d8816, 32'h3e8a03c2} /* (6, 17, 31) {real, imag} */,
  {32'h4042ac02, 32'h40016be9} /* (6, 17, 30) {real, imag} */,
  {32'hbef575d9, 32'h3e44200e} /* (6, 17, 29) {real, imag} */,
  {32'hbfb273c1, 32'h3fa061b2} /* (6, 17, 28) {real, imag} */,
  {32'hbf8829d2, 32'hbfa5aee1} /* (6, 17, 27) {real, imag} */,
  {32'hc015095b, 32'hbf925327} /* (6, 17, 26) {real, imag} */,
  {32'h3e998e6b, 32'h3f417655} /* (6, 17, 25) {real, imag} */,
  {32'h3d5f333c, 32'h3f7e0439} /* (6, 17, 24) {real, imag} */,
  {32'h3fc6191b, 32'h3f3ee991} /* (6, 17, 23) {real, imag} */,
  {32'hbf6ba6b5, 32'hbad3ba65} /* (6, 17, 22) {real, imag} */,
  {32'hbf2edd01, 32'h3fd6cb25} /* (6, 17, 21) {real, imag} */,
  {32'h3f9baa6a, 32'hbf608416} /* (6, 17, 20) {real, imag} */,
  {32'hbf88480a, 32'hbfe22591} /* (6, 17, 19) {real, imag} */,
  {32'h3e98cc4c, 32'h400fb219} /* (6, 17, 18) {real, imag} */,
  {32'hbe89eddc, 32'hbfaf980b} /* (6, 17, 17) {real, imag} */,
  {32'hc054a131, 32'h3efdb083} /* (6, 17, 16) {real, imag} */,
  {32'h4004be78, 32'hbf29917d} /* (6, 17, 15) {real, imag} */,
  {32'h3fc56e47, 32'hbf13f363} /* (6, 17, 14) {real, imag} */,
  {32'hbfbbddab, 32'hbfae14a1} /* (6, 17, 13) {real, imag} */,
  {32'hbe8942a7, 32'h3f5ebf31} /* (6, 17, 12) {real, imag} */,
  {32'h3b7ae2f8, 32'h3e251ab8} /* (6, 17, 11) {real, imag} */,
  {32'hc02a7f44, 32'hc009b310} /* (6, 17, 10) {real, imag} */,
  {32'h3dbebc79, 32'hbf2d760d} /* (6, 17, 9) {real, imag} */,
  {32'hbf380e44, 32'hbfe63b13} /* (6, 17, 8) {real, imag} */,
  {32'hbfb71c6f, 32'h3fc984f0} /* (6, 17, 7) {real, imag} */,
  {32'hbea643d8, 32'h3f62c195} /* (6, 17, 6) {real, imag} */,
  {32'hbfb069b5, 32'hbf4e7655} /* (6, 17, 5) {real, imag} */,
  {32'h3fe1e99a, 32'hbe1c870c} /* (6, 17, 4) {real, imag} */,
  {32'h3f994a48, 32'h3ffe731f} /* (6, 17, 3) {real, imag} */,
  {32'hc0873980, 32'h3f1f1471} /* (6, 17, 2) {real, imag} */,
  {32'hbf119c35, 32'h3e265ed7} /* (6, 17, 1) {real, imag} */,
  {32'hbfecfbd8, 32'hbe519dbd} /* (6, 17, 0) {real, imag} */,
  {32'h3f04af00, 32'hbf234812} /* (6, 16, 31) {real, imag} */,
  {32'h3f52bab8, 32'h3ee2161a} /* (6, 16, 30) {real, imag} */,
  {32'h3f7f6698, 32'h3ed273fc} /* (6, 16, 29) {real, imag} */,
  {32'hbf419a01, 32'hbde68fde} /* (6, 16, 28) {real, imag} */,
  {32'hbf4567b9, 32'hbf7bb584} /* (6, 16, 27) {real, imag} */,
  {32'hbeffb8fe, 32'h3f9a68cb} /* (6, 16, 26) {real, imag} */,
  {32'h3e8ce073, 32'hbf21d4f5} /* (6, 16, 25) {real, imag} */,
  {32'h3f68e110, 32'hbf77f78a} /* (6, 16, 24) {real, imag} */,
  {32'h3e8794ef, 32'h3d5d73cc} /* (6, 16, 23) {real, imag} */,
  {32'h3e9a932f, 32'h3d11b5bd} /* (6, 16, 22) {real, imag} */,
  {32'h3eee18f4, 32'h3fa1bb8f} /* (6, 16, 21) {real, imag} */,
  {32'h3fd8bb47, 32'h3e24ed12} /* (6, 16, 20) {real, imag} */,
  {32'h3f8226ca, 32'h3eac4c09} /* (6, 16, 19) {real, imag} */,
  {32'h3fc366ef, 32'hbfe4bef3} /* (6, 16, 18) {real, imag} */,
  {32'h4008dee3, 32'h3f87d890} /* (6, 16, 17) {real, imag} */,
  {32'h3e6d240d, 32'hbf93f0e0} /* (6, 16, 16) {real, imag} */,
  {32'hbecbcf9d, 32'hbf1ce9d1} /* (6, 16, 15) {real, imag} */,
  {32'h3fa611b0, 32'hc0313ba3} /* (6, 16, 14) {real, imag} */,
  {32'h3fb39c2a, 32'hbf513fd9} /* (6, 16, 13) {real, imag} */,
  {32'hbf8f14e2, 32'h3fafb8dd} /* (6, 16, 12) {real, imag} */,
  {32'h3e894f2a, 32'h3eeb3811} /* (6, 16, 11) {real, imag} */,
  {32'hbde653c5, 32'hbffa72ea} /* (6, 16, 10) {real, imag} */,
  {32'hbf694e32, 32'h3f8be399} /* (6, 16, 9) {real, imag} */,
  {32'hbe1ef30b, 32'hbe16fff3} /* (6, 16, 8) {real, imag} */,
  {32'h3e1e94ae, 32'hbea21f18} /* (6, 16, 7) {real, imag} */,
  {32'hbec1dbcb, 32'hbf78dbbb} /* (6, 16, 6) {real, imag} */,
  {32'hbf680666, 32'h3fbb4748} /* (6, 16, 5) {real, imag} */,
  {32'hbffb8f4f, 32'h3dc571fa} /* (6, 16, 4) {real, imag} */,
  {32'h3f1efb02, 32'hbf0e6195} /* (6, 16, 3) {real, imag} */,
  {32'h3dd3e79e, 32'h3f763cb5} /* (6, 16, 2) {real, imag} */,
  {32'h3b086186, 32'hbf831dc3} /* (6, 16, 1) {real, imag} */,
  {32'h3ed7c19c, 32'h3ebed2fa} /* (6, 16, 0) {real, imag} */,
  {32'h3f7d0699, 32'hbfc13c5e} /* (6, 15, 31) {real, imag} */,
  {32'h3f61a2ad, 32'h3f8dbb7f} /* (6, 15, 30) {real, imag} */,
  {32'h3e6f0adc, 32'hc00d5533} /* (6, 15, 29) {real, imag} */,
  {32'h3e3837b7, 32'h3f9e54db} /* (6, 15, 28) {real, imag} */,
  {32'hbfc2348e, 32'hbfdaac1e} /* (6, 15, 27) {real, imag} */,
  {32'h3fbfb7a8, 32'h3fc9581e} /* (6, 15, 26) {real, imag} */,
  {32'h3fa0197c, 32'hc015222a} /* (6, 15, 25) {real, imag} */,
  {32'hc04217eb, 32'hc00eb1b3} /* (6, 15, 24) {real, imag} */,
  {32'h3e94d305, 32'hbf45c660} /* (6, 15, 23) {real, imag} */,
  {32'hbef5bbac, 32'hbf6d7ac8} /* (6, 15, 22) {real, imag} */,
  {32'hc0341d61, 32'hbebdc9d7} /* (6, 15, 21) {real, imag} */,
  {32'hbe7f5604, 32'h3d8302ac} /* (6, 15, 20) {real, imag} */,
  {32'hbe94eac7, 32'h4010c9d9} /* (6, 15, 19) {real, imag} */,
  {32'hc00fa6b2, 32'hbf37226b} /* (6, 15, 18) {real, imag} */,
  {32'hbf3acb9a, 32'h3e65a00f} /* (6, 15, 17) {real, imag} */,
  {32'h3f932be9, 32'h3f409762} /* (6, 15, 16) {real, imag} */,
  {32'h3d0b1cbf, 32'hbfb77db6} /* (6, 15, 15) {real, imag} */,
  {32'hbf2da467, 32'hbf7620fd} /* (6, 15, 14) {real, imag} */,
  {32'h3f3d1716, 32'h3f9e4fbe} /* (6, 15, 13) {real, imag} */,
  {32'h3ea2aa1a, 32'h3d94c268} /* (6, 15, 12) {real, imag} */,
  {32'hc00440b5, 32'h3dda8ea2} /* (6, 15, 11) {real, imag} */,
  {32'h3fcdba1b, 32'h402c493d} /* (6, 15, 10) {real, imag} */,
  {32'hc02d3103, 32'h3fffccb4} /* (6, 15, 9) {real, imag} */,
  {32'hbfbac3f3, 32'hbfb89c13} /* (6, 15, 8) {real, imag} */,
  {32'h3f45cc8a, 32'hc000760d} /* (6, 15, 7) {real, imag} */,
  {32'hbdc57d2f, 32'h3f38738e} /* (6, 15, 6) {real, imag} */,
  {32'h3cc4560f, 32'hbfc64234} /* (6, 15, 5) {real, imag} */,
  {32'hbfe33081, 32'h3fddd7f2} /* (6, 15, 4) {real, imag} */,
  {32'h40319c8e, 32'h3dd2aa9a} /* (6, 15, 3) {real, imag} */,
  {32'hbd504e96, 32'h3ead53e2} /* (6, 15, 2) {real, imag} */,
  {32'hbf5982d9, 32'hbf570e0c} /* (6, 15, 1) {real, imag} */,
  {32'h401fd2ae, 32'h3f6d758d} /* (6, 15, 0) {real, imag} */,
  {32'hc028ee9c, 32'hbf6561e9} /* (6, 14, 31) {real, imag} */,
  {32'hbe55e0ee, 32'h400051b0} /* (6, 14, 30) {real, imag} */,
  {32'hbf29fe59, 32'h3e89bcc9} /* (6, 14, 29) {real, imag} */,
  {32'hbd1ab65e, 32'h3f803288} /* (6, 14, 28) {real, imag} */,
  {32'hbec1a9af, 32'h3f5bf4b6} /* (6, 14, 27) {real, imag} */,
  {32'hbd1fe17a, 32'h404c42a4} /* (6, 14, 26) {real, imag} */,
  {32'hbf2fba6f, 32'hbe0f1b6d} /* (6, 14, 25) {real, imag} */,
  {32'hc03b5feb, 32'hbfcc43e4} /* (6, 14, 24) {real, imag} */,
  {32'h3f952fa4, 32'hbfdf0b84} /* (6, 14, 23) {real, imag} */,
  {32'hbf9439b6, 32'hbf183f97} /* (6, 14, 22) {real, imag} */,
  {32'h3f1b2bc9, 32'h4029c36b} /* (6, 14, 21) {real, imag} */,
  {32'hbfe977f1, 32'hbfb125c6} /* (6, 14, 20) {real, imag} */,
  {32'hc00eea61, 32'hbfaa7d5e} /* (6, 14, 19) {real, imag} */,
  {32'hbfb52932, 32'hc020bf4e} /* (6, 14, 18) {real, imag} */,
  {32'h3f0b1f49, 32'h3f965de3} /* (6, 14, 17) {real, imag} */,
  {32'hbf3e5208, 32'h3fb33f8a} /* (6, 14, 16) {real, imag} */,
  {32'hbeb2e298, 32'hbf87adff} /* (6, 14, 15) {real, imag} */,
  {32'h40071fb9, 32'h3f7ee161} /* (6, 14, 14) {real, imag} */,
  {32'hbf4b0c1f, 32'h3f5eaaa8} /* (6, 14, 13) {real, imag} */,
  {32'hbf7709fa, 32'h3f81690c} /* (6, 14, 12) {real, imag} */,
  {32'hbf68e93a, 32'h3f6da19f} /* (6, 14, 11) {real, imag} */,
  {32'h3f981212, 32'h3fcbf117} /* (6, 14, 10) {real, imag} */,
  {32'h3fbc7d27, 32'h3f2abefe} /* (6, 14, 9) {real, imag} */,
  {32'hbeba69d1, 32'h402da327} /* (6, 14, 8) {real, imag} */,
  {32'h3f448e4d, 32'hbf0b3899} /* (6, 14, 7) {real, imag} */,
  {32'hc033066e, 32'h3f55ecec} /* (6, 14, 6) {real, imag} */,
  {32'h3fa69792, 32'h404a0da1} /* (6, 14, 5) {real, imag} */,
  {32'hbf349af8, 32'h3df6a3ac} /* (6, 14, 4) {real, imag} */,
  {32'h3f400449, 32'hbeb77228} /* (6, 14, 3) {real, imag} */,
  {32'h3fc2b17d, 32'h3f4ea1a1} /* (6, 14, 2) {real, imag} */,
  {32'hbef688cf, 32'hbef2ee15} /* (6, 14, 1) {real, imag} */,
  {32'hc00b42a1, 32'h3ff6ec47} /* (6, 14, 0) {real, imag} */,
  {32'h401ca526, 32'hc0376a08} /* (6, 13, 31) {real, imag} */,
  {32'hbe76248d, 32'h3f7b9ad3} /* (6, 13, 30) {real, imag} */,
  {32'h3ff77fbe, 32'hbd812b2b} /* (6, 13, 29) {real, imag} */,
  {32'h3e2a8c3b, 32'hbf660c32} /* (6, 13, 28) {real, imag} */,
  {32'h3f9c4bc2, 32'hbfcb2067} /* (6, 13, 27) {real, imag} */,
  {32'hc0276e1c, 32'hbfb14633} /* (6, 13, 26) {real, imag} */,
  {32'hbcade284, 32'hbf55eb01} /* (6, 13, 25) {real, imag} */,
  {32'h3f3a2df7, 32'hbe0db93a} /* (6, 13, 24) {real, imag} */,
  {32'h3efe2e66, 32'hbfeecee2} /* (6, 13, 23) {real, imag} */,
  {32'hbde94372, 32'h3efe1bfb} /* (6, 13, 22) {real, imag} */,
  {32'h3fc9481e, 32'h400c3ed6} /* (6, 13, 21) {real, imag} */,
  {32'h3f381e14, 32'hbfec833a} /* (6, 13, 20) {real, imag} */,
  {32'hc04a8a81, 32'hbf679101} /* (6, 13, 19) {real, imag} */,
  {32'h3fb7e5a6, 32'h3f0bcfed} /* (6, 13, 18) {real, imag} */,
  {32'h3f1c93c8, 32'h3df462de} /* (6, 13, 17) {real, imag} */,
  {32'hbebd3ea8, 32'hbfe2f582} /* (6, 13, 16) {real, imag} */,
  {32'h3f3916c9, 32'hc01029ac} /* (6, 13, 15) {real, imag} */,
  {32'h3fda6630, 32'h40c13e60} /* (6, 13, 14) {real, imag} */,
  {32'h3f83b336, 32'hbfd65d88} /* (6, 13, 13) {real, imag} */,
  {32'hc011d3c7, 32'hc01761e4} /* (6, 13, 12) {real, imag} */,
  {32'hbf715124, 32'h3e29a128} /* (6, 13, 11) {real, imag} */,
  {32'hbe3365d9, 32'h3ffde375} /* (6, 13, 10) {real, imag} */,
  {32'h3f125029, 32'hbe612b79} /* (6, 13, 9) {real, imag} */,
  {32'h3f290e11, 32'h3fce0f40} /* (6, 13, 8) {real, imag} */,
  {32'hc0320e5d, 32'hc006b8d9} /* (6, 13, 7) {real, imag} */,
  {32'hbf683461, 32'h400f1574} /* (6, 13, 6) {real, imag} */,
  {32'hc0381fc7, 32'hbfd8b0af} /* (6, 13, 5) {real, imag} */,
  {32'h40179cde, 32'h3ec6d125} /* (6, 13, 4) {real, imag} */,
  {32'hc002fd50, 32'hbea51556} /* (6, 13, 3) {real, imag} */,
  {32'hbff8bdfd, 32'hbe058189} /* (6, 13, 2) {real, imag} */,
  {32'h3e9be9d1, 32'hc016e70f} /* (6, 13, 1) {real, imag} */,
  {32'hbe2aea41, 32'hbf5e9988} /* (6, 13, 0) {real, imag} */,
  {32'hbfc0440b, 32'h3eabe591} /* (6, 12, 31) {real, imag} */,
  {32'hc060e4bc, 32'hbfd6b9b0} /* (6, 12, 30) {real, imag} */,
  {32'hbf6d6874, 32'hbe60f095} /* (6, 12, 29) {real, imag} */,
  {32'h3df04810, 32'h3fcd5b49} /* (6, 12, 28) {real, imag} */,
  {32'h3fa9ca0f, 32'h3f76d525} /* (6, 12, 27) {real, imag} */,
  {32'h3f72289c, 32'hc01fb4d1} /* (6, 12, 26) {real, imag} */,
  {32'h3fc7e1ac, 32'h4057a324} /* (6, 12, 25) {real, imag} */,
  {32'h3fc3012f, 32'hbf9aac2c} /* (6, 12, 24) {real, imag} */,
  {32'h3fcbc3ec, 32'hbe58ce91} /* (6, 12, 23) {real, imag} */,
  {32'h403a7efc, 32'h3fa8f06d} /* (6, 12, 22) {real, imag} */,
  {32'hbf7df7b5, 32'hbec2286f} /* (6, 12, 21) {real, imag} */,
  {32'h3f922ec0, 32'h3e8480ce} /* (6, 12, 20) {real, imag} */,
  {32'h4038b87a, 32'h400397ff} /* (6, 12, 19) {real, imag} */,
  {32'h3fa2108f, 32'h4009ca51} /* (6, 12, 18) {real, imag} */,
  {32'hbedba813, 32'h4001d1fa} /* (6, 12, 17) {real, imag} */,
  {32'hbf53b9e7, 32'h3df1a81f} /* (6, 12, 16) {real, imag} */,
  {32'h3daf6fd4, 32'h3f39d966} /* (6, 12, 15) {real, imag} */,
  {32'hbea2cd98, 32'h3d9752d2} /* (6, 12, 14) {real, imag} */,
  {32'h401195aa, 32'hbfa1f89e} /* (6, 12, 13) {real, imag} */,
  {32'hbf6318af, 32'h3f913d9f} /* (6, 12, 12) {real, imag} */,
  {32'h3fdbeaef, 32'h3fc560e4} /* (6, 12, 11) {real, imag} */,
  {32'h3f092773, 32'hc081fccf} /* (6, 12, 10) {real, imag} */,
  {32'h3ebc2b87, 32'hbe7bfba7} /* (6, 12, 9) {real, imag} */,
  {32'hbf2e173e, 32'h3d2ae7eb} /* (6, 12, 8) {real, imag} */,
  {32'hbf073c36, 32'h40039a42} /* (6, 12, 7) {real, imag} */,
  {32'hbfbce0c3, 32'hbf006f9b} /* (6, 12, 6) {real, imag} */,
  {32'h403c5d32, 32'h3e8f7e59} /* (6, 12, 5) {real, imag} */,
  {32'hc0058252, 32'hbf3c84f8} /* (6, 12, 4) {real, imag} */,
  {32'hbddc0b06, 32'h3db7873a} /* (6, 12, 3) {real, imag} */,
  {32'h3f4c1ddd, 32'h3ec5d8af} /* (6, 12, 2) {real, imag} */,
  {32'hc00c9537, 32'hbf298ab3} /* (6, 12, 1) {real, imag} */,
  {32'hbfceacd1, 32'hbf25738f} /* (6, 12, 0) {real, imag} */,
  {32'h3eee10cd, 32'hc0627459} /* (6, 11, 31) {real, imag} */,
  {32'h3f192d92, 32'hc0263abf} /* (6, 11, 30) {real, imag} */,
  {32'h3ead7971, 32'h3d8bf1b2} /* (6, 11, 29) {real, imag} */,
  {32'hbf42ba99, 32'h3faac074} /* (6, 11, 28) {real, imag} */,
  {32'hc08830e8, 32'hbf9cb904} /* (6, 11, 27) {real, imag} */,
  {32'h3fd8b5e3, 32'hc08ff45e} /* (6, 11, 26) {real, imag} */,
  {32'hc0118f2e, 32'h4029e430} /* (6, 11, 25) {real, imag} */,
  {32'h3ff643f7, 32'h400149fe} /* (6, 11, 24) {real, imag} */,
  {32'h3f8d18a0, 32'h3faf40de} /* (6, 11, 23) {real, imag} */,
  {32'h3f7eadef, 32'hc026a3f6} /* (6, 11, 22) {real, imag} */,
  {32'hc0462074, 32'hbfb099f6} /* (6, 11, 21) {real, imag} */,
  {32'hbfd371f0, 32'h3feb0f70} /* (6, 11, 20) {real, imag} */,
  {32'h3fa32567, 32'hbf77df1b} /* (6, 11, 19) {real, imag} */,
  {32'h3f691425, 32'h40212d42} /* (6, 11, 18) {real, imag} */,
  {32'hbf8cea31, 32'hc023b7d8} /* (6, 11, 17) {real, imag} */,
  {32'hbe73cdbf, 32'h4009f769} /* (6, 11, 16) {real, imag} */,
  {32'h402e4454, 32'hbe26c7c2} /* (6, 11, 15) {real, imag} */,
  {32'hbde40550, 32'h3fc52922} /* (6, 11, 14) {real, imag} */,
  {32'hbeaa298a, 32'h400c538c} /* (6, 11, 13) {real, imag} */,
  {32'h3fc2aecf, 32'h3fd21616} /* (6, 11, 12) {real, imag} */,
  {32'hbeb01961, 32'h3f93bdc1} /* (6, 11, 11) {real, imag} */,
  {32'hbf4ae3ad, 32'hbfb35790} /* (6, 11, 10) {real, imag} */,
  {32'h3ddf5117, 32'hbf69f1b6} /* (6, 11, 9) {real, imag} */,
  {32'hbf777948, 32'h3f2aa832} /* (6, 11, 8) {real, imag} */,
  {32'hc040561c, 32'hc0076d76} /* (6, 11, 7) {real, imag} */,
  {32'h3f558e34, 32'h3fbbc2e2} /* (6, 11, 6) {real, imag} */,
  {32'h3ebe83b6, 32'h3fe378dd} /* (6, 11, 5) {real, imag} */,
  {32'hbfe3986a, 32'h3f498b18} /* (6, 11, 4) {real, imag} */,
  {32'h3f9d2159, 32'hc0254345} /* (6, 11, 3) {real, imag} */,
  {32'h40505a04, 32'h3fc20c6f} /* (6, 11, 2) {real, imag} */,
  {32'hbf038ff5, 32'h3f2a517b} /* (6, 11, 1) {real, imag} */,
  {32'h3fe4870c, 32'h4008d44d} /* (6, 11, 0) {real, imag} */,
  {32'hbf8785c5, 32'h4011c163} /* (6, 10, 31) {real, imag} */,
  {32'h3f23cb6d, 32'h3f3fed04} /* (6, 10, 30) {real, imag} */,
  {32'hc03d4a07, 32'h3f5b3529} /* (6, 10, 29) {real, imag} */,
  {32'hbf9400ea, 32'hc01af297} /* (6, 10, 28) {real, imag} */,
  {32'hbf90ba6f, 32'h402edf8f} /* (6, 10, 27) {real, imag} */,
  {32'hbfd7ade7, 32'hbf791533} /* (6, 10, 26) {real, imag} */,
  {32'hc0367c75, 32'h3f969aed} /* (6, 10, 25) {real, imag} */,
  {32'h3c757c37, 32'hc005b9ef} /* (6, 10, 24) {real, imag} */,
  {32'h3fa6e25a, 32'h3fe1ebed} /* (6, 10, 23) {real, imag} */,
  {32'h3fe1ddfc, 32'h405075b9} /* (6, 10, 22) {real, imag} */,
  {32'hbf817183, 32'hbff27ea5} /* (6, 10, 21) {real, imag} */,
  {32'hbf5e6c0d, 32'hc00eb868} /* (6, 10, 20) {real, imag} */,
  {32'hbf2bdd08, 32'hc005e02f} /* (6, 10, 19) {real, imag} */,
  {32'h3f40c29a, 32'hbcd04858} /* (6, 10, 18) {real, imag} */,
  {32'h3f5d68e8, 32'h406cd765} /* (6, 10, 17) {real, imag} */,
  {32'h3f44890e, 32'h3dbaa56c} /* (6, 10, 16) {real, imag} */,
  {32'hbeb42c24, 32'hbf465244} /* (6, 10, 15) {real, imag} */,
  {32'hc03ff4a9, 32'h400476b6} /* (6, 10, 14) {real, imag} */,
  {32'h40432b93, 32'h3fbc4587} /* (6, 10, 13) {real, imag} */,
  {32'hbfd900c7, 32'hc0181ce5} /* (6, 10, 12) {real, imag} */,
  {32'hc0774731, 32'h402ce653} /* (6, 10, 11) {real, imag} */,
  {32'h3f1d23ec, 32'hbe277789} /* (6, 10, 10) {real, imag} */,
  {32'hbf82f6c9, 32'hc023aaca} /* (6, 10, 9) {real, imag} */,
  {32'h3f85db20, 32'h4001ed28} /* (6, 10, 8) {real, imag} */,
  {32'hbfe0a6a8, 32'h3f9a4e30} /* (6, 10, 7) {real, imag} */,
  {32'h4013b9a3, 32'h403fcedf} /* (6, 10, 6) {real, imag} */,
  {32'h3f7bcbec, 32'hc044e55c} /* (6, 10, 5) {real, imag} */,
  {32'h40811e0a, 32'h3f68e049} /* (6, 10, 4) {real, imag} */,
  {32'hbd03211b, 32'h3f996a0a} /* (6, 10, 3) {real, imag} */,
  {32'hbea63c9a, 32'hbdfa37a3} /* (6, 10, 2) {real, imag} */,
  {32'h3ef6d77d, 32'h40017ade} /* (6, 10, 1) {real, imag} */,
  {32'h3f6e59db, 32'hc004ea7d} /* (6, 10, 0) {real, imag} */,
  {32'hbf9dd291, 32'h3ffc7194} /* (6, 9, 31) {real, imag} */,
  {32'hbd522cc1, 32'hc0876fdc} /* (6, 9, 30) {real, imag} */,
  {32'hc0923c50, 32'h4007525c} /* (6, 9, 29) {real, imag} */,
  {32'hbf41ef51, 32'h3da394f7} /* (6, 9, 28) {real, imag} */,
  {32'h4050453b, 32'h3fc32053} /* (6, 9, 27) {real, imag} */,
  {32'h3f41c6dd, 32'h3f0010b3} /* (6, 9, 26) {real, imag} */,
  {32'h3f5086da, 32'h40886732} /* (6, 9, 25) {real, imag} */,
  {32'h404e8bf4, 32'h3e4c9b3b} /* (6, 9, 24) {real, imag} */,
  {32'h3f9745db, 32'hbee3b0ea} /* (6, 9, 23) {real, imag} */,
  {32'hc05120f2, 32'hbf528d3b} /* (6, 9, 22) {real, imag} */,
  {32'h3f27e291, 32'hbfb72aab} /* (6, 9, 21) {real, imag} */,
  {32'hbfe18918, 32'h400dfee2} /* (6, 9, 20) {real, imag} */,
  {32'hbf310ad0, 32'hc00259e5} /* (6, 9, 19) {real, imag} */,
  {32'h3eea3c57, 32'hbf70ced5} /* (6, 9, 18) {real, imag} */,
  {32'h3f880573, 32'h3fa25030} /* (6, 9, 17) {real, imag} */,
  {32'h3f21a260, 32'h3ec5552d} /* (6, 9, 16) {real, imag} */,
  {32'h40116019, 32'h3eb4dd5c} /* (6, 9, 15) {real, imag} */,
  {32'h3d2837fd, 32'hc0653f65} /* (6, 9, 14) {real, imag} */,
  {32'h3fd8c8d7, 32'h3fad7993} /* (6, 9, 13) {real, imag} */,
  {32'h3fee31c3, 32'hbe585e73} /* (6, 9, 12) {real, imag} */,
  {32'h3e0d6009, 32'h3ff3ecf1} /* (6, 9, 11) {real, imag} */,
  {32'hbe867f2b, 32'hbe363727} /* (6, 9, 10) {real, imag} */,
  {32'h408bbaec, 32'hbfb75de9} /* (6, 9, 9) {real, imag} */,
  {32'h3f8db2d6, 32'h3e70adc2} /* (6, 9, 8) {real, imag} */,
  {32'h40778d07, 32'hc04d752e} /* (6, 9, 7) {real, imag} */,
  {32'h3f1e1dcc, 32'h3fd2a41a} /* (6, 9, 6) {real, imag} */,
  {32'h3f177b88, 32'h3fba4309} /* (6, 9, 5) {real, imag} */,
  {32'hbfdba76f, 32'hbfac408b} /* (6, 9, 4) {real, imag} */,
  {32'h40754288, 32'h4000d935} /* (6, 9, 3) {real, imag} */,
  {32'h40641196, 32'h3e4053c9} /* (6, 9, 2) {real, imag} */,
  {32'hbf20550a, 32'h3e3efe72} /* (6, 9, 1) {real, imag} */,
  {32'hbe992be7, 32'h40e18d71} /* (6, 9, 0) {real, imag} */,
  {32'h3ea1b563, 32'h4026e9af} /* (6, 8, 31) {real, imag} */,
  {32'h400b176a, 32'hbfb3371c} /* (6, 8, 30) {real, imag} */,
  {32'hbfcd5d8f, 32'h40507b88} /* (6, 8, 29) {real, imag} */,
  {32'hc0388e5e, 32'hc04764a2} /* (6, 8, 28) {real, imag} */,
  {32'hc066521e, 32'hc008485e} /* (6, 8, 27) {real, imag} */,
  {32'hbfe63b45, 32'h408d0b30} /* (6, 8, 26) {real, imag} */,
  {32'hbf2a19bd, 32'hbffd715d} /* (6, 8, 25) {real, imag} */,
  {32'h3f1aca0c, 32'h40256bef} /* (6, 8, 24) {real, imag} */,
  {32'h405e4209, 32'hc08cf861} /* (6, 8, 23) {real, imag} */,
  {32'hbfba8024, 32'h3ff5484a} /* (6, 8, 22) {real, imag} */,
  {32'hbfa750ad, 32'hbf2746f3} /* (6, 8, 21) {real, imag} */,
  {32'hbde3d9b7, 32'hbf798e3c} /* (6, 8, 20) {real, imag} */,
  {32'hc00af6a5, 32'hc00df1db} /* (6, 8, 19) {real, imag} */,
  {32'hbf985a73, 32'hbeacc059} /* (6, 8, 18) {real, imag} */,
  {32'h3f630c4b, 32'h3f5c30c6} /* (6, 8, 17) {real, imag} */,
  {32'h3eca2b8b, 32'hbf4338cd} /* (6, 8, 16) {real, imag} */,
  {32'h3ded34e9, 32'hbf6f47ad} /* (6, 8, 15) {real, imag} */,
  {32'hc004c6f0, 32'h3e7809d0} /* (6, 8, 14) {real, imag} */,
  {32'hbec3c69c, 32'h40925b33} /* (6, 8, 13) {real, imag} */,
  {32'h3f7d154a, 32'hc067c5d5} /* (6, 8, 12) {real, imag} */,
  {32'hbf47e9dc, 32'hbfa32ca7} /* (6, 8, 11) {real, imag} */,
  {32'hc003d8d9, 32'hbf19c529} /* (6, 8, 10) {real, imag} */,
  {32'h3f31eade, 32'h3fffbab3} /* (6, 8, 9) {real, imag} */,
  {32'h4004a31f, 32'hc01e0f5a} /* (6, 8, 8) {real, imag} */,
  {32'h401e9261, 32'hbdd0774a} /* (6, 8, 7) {real, imag} */,
  {32'hbf4c1b81, 32'h400d3d7e} /* (6, 8, 6) {real, imag} */,
  {32'hc025376b, 32'hbe1fef39} /* (6, 8, 5) {real, imag} */,
  {32'hc089f3b5, 32'hbf9be7d7} /* (6, 8, 4) {real, imag} */,
  {32'hbf978c2b, 32'hc0269671} /* (6, 8, 3) {real, imag} */,
  {32'h3e5620ff, 32'h3fbc79a3} /* (6, 8, 2) {real, imag} */,
  {32'hbfaf2cd4, 32'h407a0d19} /* (6, 8, 1) {real, imag} */,
  {32'h3ec5eb66, 32'hbf4bc3cc} /* (6, 8, 0) {real, imag} */,
  {32'h3fc324c6, 32'h40b210e1} /* (6, 7, 31) {real, imag} */,
  {32'h4074d4ba, 32'hc0a6e606} /* (6, 7, 30) {real, imag} */,
  {32'h3ff36b32, 32'h40088079} /* (6, 7, 29) {real, imag} */,
  {32'h40630b8f, 32'hbf1fe4e8} /* (6, 7, 28) {real, imag} */,
  {32'hc02406f5, 32'hc0338707} /* (6, 7, 27) {real, imag} */,
  {32'h3edbccf1, 32'h4056a618} /* (6, 7, 26) {real, imag} */,
  {32'h40a1982b, 32'hbf359295} /* (6, 7, 25) {real, imag} */,
  {32'hc008d310, 32'h3df059c9} /* (6, 7, 24) {real, imag} */,
  {32'hbff55c28, 32'hbe8a5d77} /* (6, 7, 23) {real, imag} */,
  {32'h4000b0e4, 32'h3e8ffa3e} /* (6, 7, 22) {real, imag} */,
  {32'h40886654, 32'hbf3e7491} /* (6, 7, 21) {real, imag} */,
  {32'hbfd46c0c, 32'hbf98f295} /* (6, 7, 20) {real, imag} */,
  {32'h3f67505f, 32'h3f6af4aa} /* (6, 7, 19) {real, imag} */,
  {32'hbd915c9d, 32'h3e35d4de} /* (6, 7, 18) {real, imag} */,
  {32'hc07b2d16, 32'h3f64ab32} /* (6, 7, 17) {real, imag} */,
  {32'h3f8bc452, 32'h3fd897c7} /* (6, 7, 16) {real, imag} */,
  {32'hc01fac40, 32'hc00fc751} /* (6, 7, 15) {real, imag} */,
  {32'hbfe55b7b, 32'hc0087eac} /* (6, 7, 14) {real, imag} */,
  {32'hc01539cd, 32'h3da27fd2} /* (6, 7, 13) {real, imag} */,
  {32'hc01c73d2, 32'hbfaa3ea6} /* (6, 7, 12) {real, imag} */,
  {32'hc032baf8, 32'hbe9a5d9f} /* (6, 7, 11) {real, imag} */,
  {32'h405b7d15, 32'hc00624bb} /* (6, 7, 10) {real, imag} */,
  {32'h401b37c6, 32'hbef01082} /* (6, 7, 9) {real, imag} */,
  {32'hbfeb9576, 32'hbfa7ac6c} /* (6, 7, 8) {real, imag} */,
  {32'hbe077fe5, 32'h3db4d627} /* (6, 7, 7) {real, imag} */,
  {32'h3e901b9b, 32'h3f6e4e26} /* (6, 7, 6) {real, imag} */,
  {32'hc015fa14, 32'h3eef3a1f} /* (6, 7, 5) {real, imag} */,
  {32'h40e1cb89, 32'hbfa81189} /* (6, 7, 4) {real, imag} */,
  {32'h40cda99a, 32'h3fd4dcc3} /* (6, 7, 3) {real, imag} */,
  {32'hc06abe98, 32'h400a08c2} /* (6, 7, 2) {real, imag} */,
  {32'h3f1d0cae, 32'hbfddd69a} /* (6, 7, 1) {real, imag} */,
  {32'hc0135aa7, 32'hc0ba7ca0} /* (6, 7, 0) {real, imag} */,
  {32'hbf6c405a, 32'hbf6497c5} /* (6, 6, 31) {real, imag} */,
  {32'hc0b8876e, 32'hc01ff751} /* (6, 6, 30) {real, imag} */,
  {32'h3fec65f6, 32'hbf3ef286} /* (6, 6, 29) {real, imag} */,
  {32'h401a30bb, 32'h406574e7} /* (6, 6, 28) {real, imag} */,
  {32'h401c4a3d, 32'hc03ba499} /* (6, 6, 27) {real, imag} */,
  {32'h3f1744d3, 32'hbf6add00} /* (6, 6, 26) {real, imag} */,
  {32'h4006d6a2, 32'hbfd2e224} /* (6, 6, 25) {real, imag} */,
  {32'h3f920603, 32'h3e884d98} /* (6, 6, 24) {real, imag} */,
  {32'hc0764b54, 32'h3f2f4879} /* (6, 6, 23) {real, imag} */,
  {32'h3e6664ea, 32'h3ea287c6} /* (6, 6, 22) {real, imag} */,
  {32'h3fd0943b, 32'h3fb1554a} /* (6, 6, 21) {real, imag} */,
  {32'hc01c9ce9, 32'hc0739c27} /* (6, 6, 20) {real, imag} */,
  {32'hbe7793a8, 32'hc0002282} /* (6, 6, 19) {real, imag} */,
  {32'hbf1b1d84, 32'h40605020} /* (6, 6, 18) {real, imag} */,
  {32'h3fcbe06d, 32'hbf36d20a} /* (6, 6, 17) {real, imag} */,
  {32'hbe93a315, 32'h4025a53d} /* (6, 6, 16) {real, imag} */,
  {32'hbfa7e70e, 32'h3fa0b9ce} /* (6, 6, 15) {real, imag} */,
  {32'hbf5238cf, 32'h3f5c9230} /* (6, 6, 14) {real, imag} */,
  {32'h3fc8a97a, 32'hbeaf817f} /* (6, 6, 13) {real, imag} */,
  {32'h3e3fe59e, 32'hbf4049a4} /* (6, 6, 12) {real, imag} */,
  {32'hbfde75c1, 32'h3e7ac317} /* (6, 6, 11) {real, imag} */,
  {32'hc0977cdf, 32'h408c6e64} /* (6, 6, 10) {real, imag} */,
  {32'h402dfd9c, 32'hc004a85a} /* (6, 6, 9) {real, imag} */,
  {32'hc0377333, 32'hbfa7f883} /* (6, 6, 8) {real, imag} */,
  {32'h40114447, 32'hc0df1fa6} /* (6, 6, 7) {real, imag} */,
  {32'hbf6b6f7a, 32'h3fc556d9} /* (6, 6, 6) {real, imag} */,
  {32'hbf9e28c8, 32'h409f3e10} /* (6, 6, 5) {real, imag} */,
  {32'hc00136ed, 32'hc01ce551} /* (6, 6, 4) {real, imag} */,
  {32'h3f652bc5, 32'hc037b723} /* (6, 6, 3) {real, imag} */,
  {32'h3f40747d, 32'h3fe58c61} /* (6, 6, 2) {real, imag} */,
  {32'h3faa677d, 32'h40009b89} /* (6, 6, 1) {real, imag} */,
  {32'hbf1908b5, 32'hc0595e66} /* (6, 6, 0) {real, imag} */,
  {32'h3f3b570a, 32'h3fa61197} /* (6, 5, 31) {real, imag} */,
  {32'h408baa81, 32'h3df9e99a} /* (6, 5, 30) {real, imag} */,
  {32'hc0b0fc94, 32'h40204bbc} /* (6, 5, 29) {real, imag} */,
  {32'h3e554d58, 32'h40f401f8} /* (6, 5, 28) {real, imag} */,
  {32'h3f9ed637, 32'hc00f332f} /* (6, 5, 27) {real, imag} */,
  {32'hbfe5678a, 32'h3e84dbb4} /* (6, 5, 26) {real, imag} */,
  {32'hbfe8ec74, 32'hbfc71690} /* (6, 5, 25) {real, imag} */,
  {32'hc05553a0, 32'hbf99a487} /* (6, 5, 24) {real, imag} */,
  {32'hbfa2d56b, 32'hc019b1dc} /* (6, 5, 23) {real, imag} */,
  {32'h3ba9ee3b, 32'hbfcecced} /* (6, 5, 22) {real, imag} */,
  {32'hc03564fc, 32'hc053665b} /* (6, 5, 21) {real, imag} */,
  {32'h3fc2c72e, 32'hc0155204} /* (6, 5, 20) {real, imag} */,
  {32'h3d87cd45, 32'hbf4600d6} /* (6, 5, 19) {real, imag} */,
  {32'h3fa837c3, 32'hbe9be891} /* (6, 5, 18) {real, imag} */,
  {32'hbed6e592, 32'hc01f99f7} /* (6, 5, 17) {real, imag} */,
  {32'hc0515bef, 32'hbfaa0599} /* (6, 5, 16) {real, imag} */,
  {32'hbc39cecd, 32'h4005cc26} /* (6, 5, 15) {real, imag} */,
  {32'h3e609241, 32'h3f6e2563} /* (6, 5, 14) {real, imag} */,
  {32'h40298669, 32'h3f84df96} /* (6, 5, 13) {real, imag} */,
  {32'hc06c0f0b, 32'hbe8a40fe} /* (6, 5, 12) {real, imag} */,
  {32'h3ffa659c, 32'h3ee53f81} /* (6, 5, 11) {real, imag} */,
  {32'hc057289c, 32'h3ff8f978} /* (6, 5, 10) {real, imag} */,
  {32'hbec5d478, 32'hc08d1901} /* (6, 5, 9) {real, imag} */,
  {32'hbf89d831, 32'hbec66967} /* (6, 5, 8) {real, imag} */,
  {32'h3fed661f, 32'h40922340} /* (6, 5, 7) {real, imag} */,
  {32'h3f7cdaa0, 32'hbe0fa616} /* (6, 5, 6) {real, imag} */,
  {32'h3f5c9302, 32'hbf524488} /* (6, 5, 5) {real, imag} */,
  {32'h4006fad8, 32'h3fc51e82} /* (6, 5, 4) {real, imag} */,
  {32'hbf06a079, 32'h3d372c5d} /* (6, 5, 3) {real, imag} */,
  {32'hbfbf8687, 32'hc08ac48e} /* (6, 5, 2) {real, imag} */,
  {32'h4067b859, 32'hc06af89b} /* (6, 5, 1) {real, imag} */,
  {32'hc0a5ff76, 32'h400cf3cd} /* (6, 5, 0) {real, imag} */,
  {32'h3e2b9e70, 32'h40694071} /* (6, 4, 31) {real, imag} */,
  {32'h3dad635a, 32'hbf0cf19e} /* (6, 4, 30) {real, imag} */,
  {32'h3f31c94d, 32'hc0d09fc5} /* (6, 4, 29) {real, imag} */,
  {32'hc0993046, 32'h408de49c} /* (6, 4, 28) {real, imag} */,
  {32'h4007c61c, 32'hc0108763} /* (6, 4, 27) {real, imag} */,
  {32'hbcee8db6, 32'hc0904e26} /* (6, 4, 26) {real, imag} */,
  {32'hc057ab43, 32'h3fa53ff3} /* (6, 4, 25) {real, imag} */,
  {32'h3fad1275, 32'hbfab780a} /* (6, 4, 24) {real, imag} */,
  {32'hbff4d61d, 32'h407d1a78} /* (6, 4, 23) {real, imag} */,
  {32'h401ea21c, 32'h4000137f} /* (6, 4, 22) {real, imag} */,
  {32'hc02b9eae, 32'h3f96eb80} /* (6, 4, 21) {real, imag} */,
  {32'h401e087c, 32'h3f516b46} /* (6, 4, 20) {real, imag} */,
  {32'h3fb50ce1, 32'h4031ca38} /* (6, 4, 19) {real, imag} */,
  {32'h3e50d875, 32'hbe495b8d} /* (6, 4, 18) {real, imag} */,
  {32'hc003b0e1, 32'hbd593a13} /* (6, 4, 17) {real, imag} */,
  {32'h3ee8d7ce, 32'hbfb067e6} /* (6, 4, 16) {real, imag} */,
  {32'h3ec6baa1, 32'h3f298374} /* (6, 4, 15) {real, imag} */,
  {32'hbd641b5b, 32'h3e087ced} /* (6, 4, 14) {real, imag} */,
  {32'hbeecfcd8, 32'hbeeb253e} /* (6, 4, 13) {real, imag} */,
  {32'hbf97d385, 32'h3e5315fc} /* (6, 4, 12) {real, imag} */,
  {32'h3fdf4300, 32'h3f132931} /* (6, 4, 11) {real, imag} */,
  {32'h4017486a, 32'hbf5bb70d} /* (6, 4, 10) {real, imag} */,
  {32'hc0950b40, 32'h400c2721} /* (6, 4, 9) {real, imag} */,
  {32'hc0245e40, 32'h3ec46166} /* (6, 4, 8) {real, imag} */,
  {32'hc03e9322, 32'hbda085d5} /* (6, 4, 7) {real, imag} */,
  {32'h3f88ae55, 32'hbfe1c387} /* (6, 4, 6) {real, imag} */,
  {32'h3f65fc91, 32'h40012ccc} /* (6, 4, 5) {real, imag} */,
  {32'h3fdc2c2b, 32'hc028e9bc} /* (6, 4, 4) {real, imag} */,
  {32'hc04fc698, 32'hc0d783f5} /* (6, 4, 3) {real, imag} */,
  {32'hbfd45848, 32'h40060e3e} /* (6, 4, 2) {real, imag} */,
  {32'h408c4afe, 32'h3fd16813} /* (6, 4, 1) {real, imag} */,
  {32'h40796794, 32'hbfd6a601} /* (6, 4, 0) {real, imag} */,
  {32'h4003a051, 32'h40db2f83} /* (6, 3, 31) {real, imag} */,
  {32'h4039cad5, 32'hc036926a} /* (6, 3, 30) {real, imag} */,
  {32'h3f62ba39, 32'h3f8e6837} /* (6, 3, 29) {real, imag} */,
  {32'h3f74e174, 32'h3fb99042} /* (6, 3, 28) {real, imag} */,
  {32'hbe90aad0, 32'hbfaeb037} /* (6, 3, 27) {real, imag} */,
  {32'h3fa31404, 32'h40420fb4} /* (6, 3, 26) {real, imag} */,
  {32'h3e975dd1, 32'hc0629c63} /* (6, 3, 25) {real, imag} */,
  {32'h3eb0fa07, 32'hbe07b6b6} /* (6, 3, 24) {real, imag} */,
  {32'h3fb52286, 32'hc0256647} /* (6, 3, 23) {real, imag} */,
  {32'h3edaa3b0, 32'hc083f50e} /* (6, 3, 22) {real, imag} */,
  {32'h400a163a, 32'h409ee6fa} /* (6, 3, 21) {real, imag} */,
  {32'hbfddb37b, 32'h3f16d481} /* (6, 3, 20) {real, imag} */,
  {32'h3fd21d92, 32'h3ee0d861} /* (6, 3, 19) {real, imag} */,
  {32'hbdfc664c, 32'hbfc8e794} /* (6, 3, 18) {real, imag} */,
  {32'h3ef2480e, 32'h3f8a7ea8} /* (6, 3, 17) {real, imag} */,
  {32'h4000a010, 32'h3fb2bfb8} /* (6, 3, 16) {real, imag} */,
  {32'hbd1e3d90, 32'h3f5faab7} /* (6, 3, 15) {real, imag} */,
  {32'h3f460090, 32'hc040bb10} /* (6, 3, 14) {real, imag} */,
  {32'h3de224b2, 32'hbf45a578} /* (6, 3, 13) {real, imag} */,
  {32'hc0029e8b, 32'hbee2df02} /* (6, 3, 12) {real, imag} */,
  {32'hbd84e2fa, 32'hbff69bc3} /* (6, 3, 11) {real, imag} */,
  {32'hbd9430d8, 32'hbf17bf8b} /* (6, 3, 10) {real, imag} */,
  {32'hbf4e15d5, 32'hbf320b60} /* (6, 3, 9) {real, imag} */,
  {32'hbfb15f48, 32'hbeb4a96e} /* (6, 3, 8) {real, imag} */,
  {32'hbfac9b5f, 32'hbf5467b3} /* (6, 3, 7) {real, imag} */,
  {32'hbfcaa794, 32'h3f076948} /* (6, 3, 6) {real, imag} */,
  {32'h3f4b099e, 32'hc0cde56b} /* (6, 3, 5) {real, imag} */,
  {32'h400ea393, 32'hbf3af0db} /* (6, 3, 4) {real, imag} */,
  {32'hc0ac7eaf, 32'h40363480} /* (6, 3, 3) {real, imag} */,
  {32'h40818f2c, 32'h3e64e367} /* (6, 3, 2) {real, imag} */,
  {32'h409e1ac8, 32'hc09c9657} /* (6, 3, 1) {real, imag} */,
  {32'hbfe5c67b, 32'h406f525c} /* (6, 3, 0) {real, imag} */,
  {32'h4177f004, 32'h3f45dfa0} /* (6, 2, 31) {real, imag} */,
  {32'h40111794, 32'hbf6a094c} /* (6, 2, 30) {real, imag} */,
  {32'hc08aa37f, 32'hbf8961d1} /* (6, 2, 29) {real, imag} */,
  {32'hc0732384, 32'hc0bbbcdd} /* (6, 2, 28) {real, imag} */,
  {32'hc00519da, 32'h4051c7be} /* (6, 2, 27) {real, imag} */,
  {32'hc0540ec3, 32'h3f08e127} /* (6, 2, 26) {real, imag} */,
  {32'h408d016f, 32'hbf2f1e01} /* (6, 2, 25) {real, imag} */,
  {32'hc086f4a6, 32'h4072a58f} /* (6, 2, 24) {real, imag} */,
  {32'hbe91cc60, 32'h4063b0f8} /* (6, 2, 23) {real, imag} */,
  {32'h3d3d5e44, 32'hc02df3d3} /* (6, 2, 22) {real, imag} */,
  {32'hbf45b2b5, 32'hc04cd1b1} /* (6, 2, 21) {real, imag} */,
  {32'h3e956e2b, 32'h400327d7} /* (6, 2, 20) {real, imag} */,
  {32'h3f64a396, 32'hbf1596ac} /* (6, 2, 19) {real, imag} */,
  {32'hbe659c17, 32'h3ed4bd46} /* (6, 2, 18) {real, imag} */,
  {32'h3f17f216, 32'hbdf3b102} /* (6, 2, 17) {real, imag} */,
  {32'h3f0bec93, 32'h3f2fe88e} /* (6, 2, 16) {real, imag} */,
  {32'h3d608073, 32'h3f3c1301} /* (6, 2, 15) {real, imag} */,
  {32'h3e1f833e, 32'hbfc1092a} /* (6, 2, 14) {real, imag} */,
  {32'hbebaee0e, 32'h3f3ee320} /* (6, 2, 13) {real, imag} */,
  {32'hbf9ddb82, 32'h400b93bc} /* (6, 2, 12) {real, imag} */,
  {32'hbd780b4c, 32'h3f00bad3} /* (6, 2, 11) {real, imag} */,
  {32'hbf3c4a28, 32'hbf5a84b0} /* (6, 2, 10) {real, imag} */,
  {32'hc00260d3, 32'hbcea575b} /* (6, 2, 9) {real, imag} */,
  {32'h40337ebb, 32'h3fc2ca4a} /* (6, 2, 8) {real, imag} */,
  {32'hc01384c3, 32'h402ac462} /* (6, 2, 7) {real, imag} */,
  {32'h40174786, 32'h4021126d} /* (6, 2, 6) {real, imag} */,
  {32'hc07814a4, 32'h4029bbc2} /* (6, 2, 5) {real, imag} */,
  {32'h3f45075f, 32'h4045920f} /* (6, 2, 4) {real, imag} */,
  {32'h408ed09f, 32'hc097124e} /* (6, 2, 3) {real, imag} */,
  {32'hc021b009, 32'hc08f9777} /* (6, 2, 2) {real, imag} */,
  {32'hc094fde1, 32'h400574d0} /* (6, 2, 1) {real, imag} */,
  {32'hc04bb2ad, 32'hc0d9123d} /* (6, 2, 0) {real, imag} */,
  {32'hc00d659d, 32'hbffdb69d} /* (6, 1, 31) {real, imag} */,
  {32'hbfa02e9b, 32'hc02730e6} /* (6, 1, 30) {real, imag} */,
  {32'hbfc7890e, 32'hc09daa5a} /* (6, 1, 29) {real, imag} */,
  {32'h409a9625, 32'h408eb14c} /* (6, 1, 28) {real, imag} */,
  {32'h3f17178b, 32'hbeaf24de} /* (6, 1, 27) {real, imag} */,
  {32'h402c43b9, 32'hbfec328e} /* (6, 1, 26) {real, imag} */,
  {32'hbf8a8852, 32'hbe42121d} /* (6, 1, 25) {real, imag} */,
  {32'hbda22654, 32'hc077f0bf} /* (6, 1, 24) {real, imag} */,
  {32'hc031aec7, 32'hc022b2d0} /* (6, 1, 23) {real, imag} */,
  {32'h405cc29b, 32'h3f831b1f} /* (6, 1, 22) {real, imag} */,
  {32'hc0244862, 32'h3eb538b9} /* (6, 1, 21) {real, imag} */,
  {32'h4003492a, 32'h4060efa2} /* (6, 1, 20) {real, imag} */,
  {32'hbf274220, 32'h3f4c7075} /* (6, 1, 19) {real, imag} */,
  {32'h40553579, 32'h3f45d2db} /* (6, 1, 18) {real, imag} */,
  {32'h3f50d2f5, 32'h3ed5c50a} /* (6, 1, 17) {real, imag} */,
  {32'hbf970166, 32'h3b70d60b} /* (6, 1, 16) {real, imag} */,
  {32'h3f630e27, 32'h3f20c22e} /* (6, 1, 15) {real, imag} */,
  {32'h3dc3d062, 32'hc06662a7} /* (6, 1, 14) {real, imag} */,
  {32'hbf94b634, 32'h4092b145} /* (6, 1, 13) {real, imag} */,
  {32'hbfe927c5, 32'hbfbe7e27} /* (6, 1, 12) {real, imag} */,
  {32'hbfcf6ced, 32'h3f841dee} /* (6, 1, 11) {real, imag} */,
  {32'hbeca6573, 32'hbf457d48} /* (6, 1, 10) {real, imag} */,
  {32'h3d8ea803, 32'h3e844276} /* (6, 1, 9) {real, imag} */,
  {32'hbfe38f38, 32'h3dea8ccb} /* (6, 1, 8) {real, imag} */,
  {32'hc00cdb3f, 32'hbf047097} /* (6, 1, 7) {real, imag} */,
  {32'hbfdc08f6, 32'hbf86795b} /* (6, 1, 6) {real, imag} */,
  {32'h3fd042bf, 32'h3f547200} /* (6, 1, 5) {real, imag} */,
  {32'h405ef213, 32'h3eee749f} /* (6, 1, 4) {real, imag} */,
  {32'hbfddd0c4, 32'h3fc5c2f0} /* (6, 1, 3) {real, imag} */,
  {32'hc0a165ba, 32'h3fd8d645} /* (6, 1, 2) {real, imag} */,
  {32'h40254c21, 32'h4010b9cb} /* (6, 1, 1) {real, imag} */,
  {32'h40da89fd, 32'hc0ada06d} /* (6, 1, 0) {real, imag} */,
  {32'h3f381d16, 32'h40c43062} /* (6, 0, 31) {real, imag} */,
  {32'hc0dc3da7, 32'hbf64887e} /* (6, 0, 30) {real, imag} */,
  {32'h3e1fd7e6, 32'h3d5d435f} /* (6, 0, 29) {real, imag} */,
  {32'hbf97bb6a, 32'hc084127d} /* (6, 0, 28) {real, imag} */,
  {32'h4092bdb7, 32'h410bbc7b} /* (6, 0, 27) {real, imag} */,
  {32'h3e4b256f, 32'h3fe8122e} /* (6, 0, 26) {real, imag} */,
  {32'h3fae9a81, 32'hbfc39489} /* (6, 0, 25) {real, imag} */,
  {32'hbf7c3987, 32'hc09b274a} /* (6, 0, 24) {real, imag} */,
  {32'hbfe42acf, 32'h3f66f86b} /* (6, 0, 23) {real, imag} */,
  {32'h3fedc330, 32'h3fde1e51} /* (6, 0, 22) {real, imag} */,
  {32'hbf45ebd9, 32'hbf04edc0} /* (6, 0, 21) {real, imag} */,
  {32'h3f7d94d2, 32'h3eae23dd} /* (6, 0, 20) {real, imag} */,
  {32'h3f3c2d37, 32'h3fb4a9e9} /* (6, 0, 19) {real, imag} */,
  {32'hbfdd25f5, 32'h3e6d4e17} /* (6, 0, 18) {real, imag} */,
  {32'hbff50780, 32'h3e8f0233} /* (6, 0, 17) {real, imag} */,
  {32'hbef56a0b, 32'h400732f1} /* (6, 0, 16) {real, imag} */,
  {32'hbf111999, 32'hbf271b7e} /* (6, 0, 15) {real, imag} */,
  {32'h3fbb126b, 32'h402da3b5} /* (6, 0, 14) {real, imag} */,
  {32'hc05269f2, 32'hbff7c591} /* (6, 0, 13) {real, imag} */,
  {32'h3ee38372, 32'hbfe61ccd} /* (6, 0, 12) {real, imag} */,
  {32'h3f2e2b6b, 32'hc052b595} /* (6, 0, 11) {real, imag} */,
  {32'hbf990497, 32'hc028456c} /* (6, 0, 10) {real, imag} */,
  {32'hbf7a539e, 32'hbfadfb1a} /* (6, 0, 9) {real, imag} */,
  {32'hbf968e29, 32'hbf50adcd} /* (6, 0, 8) {real, imag} */,
  {32'h40a61a8b, 32'hc019199d} /* (6, 0, 7) {real, imag} */,
  {32'hbf0c8e4a, 32'h3fd787ce} /* (6, 0, 6) {real, imag} */,
  {32'hbfc27fa9, 32'hc06aae23} /* (6, 0, 5) {real, imag} */,
  {32'hc02b48eb, 32'hc095414c} /* (6, 0, 4) {real, imag} */,
  {32'h3e7dbb0b, 32'h4007a621} /* (6, 0, 3) {real, imag} */,
  {32'h40bc2028, 32'h40db7cb5} /* (6, 0, 2) {real, imag} */,
  {32'h40737003, 32'h3fa344c0} /* (6, 0, 1) {real, imag} */,
  {32'h40fce6ce, 32'h40e29fd0} /* (6, 0, 0) {real, imag} */,
  {32'h3f566ac7, 32'hc20fff4d} /* (5, 31, 31) {real, imag} */,
  {32'h412302a0, 32'h41a09a80} /* (5, 31, 30) {real, imag} */,
  {32'hbd4191cf, 32'h412f0c18} /* (5, 31, 29) {real, imag} */,
  {32'hbfb114fa, 32'hc079456f} /* (5, 31, 28) {real, imag} */,
  {32'hbfc70060, 32'h4018e11d} /* (5, 31, 27) {real, imag} */,
  {32'h405d669e, 32'h3dc0627e} /* (5, 31, 26) {real, imag} */,
  {32'h405a8f36, 32'hc082c89c} /* (5, 31, 25) {real, imag} */,
  {32'h3f96c8fb, 32'h40ef1ee6} /* (5, 31, 24) {real, imag} */,
  {32'hbf51b2b5, 32'h3ff66049} /* (5, 31, 23) {real, imag} */,
  {32'h3e617b9a, 32'h3ea7a5d4} /* (5, 31, 22) {real, imag} */,
  {32'hbecfac62, 32'h403b0c96} /* (5, 31, 21) {real, imag} */,
  {32'h3f327c75, 32'hbf28ada2} /* (5, 31, 20) {real, imag} */,
  {32'h3fd97a92, 32'hbfd8e425} /* (5, 31, 19) {real, imag} */,
  {32'h3fd33820, 32'hc0286d7f} /* (5, 31, 18) {real, imag} */,
  {32'hbf6d8895, 32'h3ff7cc2c} /* (5, 31, 17) {real, imag} */,
  {32'h3f7377e9, 32'hbecec20d} /* (5, 31, 16) {real, imag} */,
  {32'h3e38d079, 32'h3fad38c6} /* (5, 31, 15) {real, imag} */,
  {32'h3e44b447, 32'h3fdd867e} /* (5, 31, 14) {real, imag} */,
  {32'h3eef630c, 32'h3f0b56b3} /* (5, 31, 13) {real, imag} */,
  {32'hbf294eac, 32'hc00e3b14} /* (5, 31, 12) {real, imag} */,
  {32'hbfb3cb61, 32'h3e486256} /* (5, 31, 11) {real, imag} */,
  {32'h3f310329, 32'hbebb188b} /* (5, 31, 10) {real, imag} */,
  {32'hbf2c7b1b, 32'hbe36ccf8} /* (5, 31, 9) {real, imag} */,
  {32'hc0735bea, 32'h4000afaa} /* (5, 31, 8) {real, imag} */,
  {32'hbf168fc2, 32'hc0dc7c6e} /* (5, 31, 7) {real, imag} */,
  {32'hbfdd9fcb, 32'h3a02e6c4} /* (5, 31, 6) {real, imag} */,
  {32'hc11d150a, 32'h40adf41d} /* (5, 31, 5) {real, imag} */,
  {32'h409b6c95, 32'hbe5219cc} /* (5, 31, 4) {real, imag} */,
  {32'h402ad420, 32'hbff72679} /* (5, 31, 3) {real, imag} */,
  {32'hc0e75f58, 32'h40ea406e} /* (5, 31, 2) {real, imag} */,
  {32'h41da5ff9, 32'hc19094fc} /* (5, 31, 1) {real, imag} */,
  {32'h4119c833, 32'hc1f9609c} /* (5, 31, 0) {real, imag} */,
  {32'hc11282a5, 32'h41938103} /* (5, 30, 31) {real, imag} */,
  {32'h413d996e, 32'hc1975b94} /* (5, 30, 30) {real, imag} */,
  {32'h3f0e996d, 32'hbf4d643d} /* (5, 30, 29) {real, imag} */,
  {32'hc01541ec, 32'h40b22f88} /* (5, 30, 28) {real, imag} */,
  {32'hc0567007, 32'hc0e2ed8a} /* (5, 30, 27) {real, imag} */,
  {32'h40508184, 32'h403df438} /* (5, 30, 26) {real, imag} */,
  {32'hc027a38e, 32'h3fe5d850} /* (5, 30, 25) {real, imag} */,
  {32'h3f10ba7f, 32'h402f5192} /* (5, 30, 24) {real, imag} */,
  {32'hbfc42388, 32'h3f87605b} /* (5, 30, 23) {real, imag} */,
  {32'h3fa17119, 32'h3f7ca388} /* (5, 30, 22) {real, imag} */,
  {32'hbeabc85a, 32'h3da4229a} /* (5, 30, 21) {real, imag} */,
  {32'hbd7cce16, 32'h3f377f67} /* (5, 30, 20) {real, imag} */,
  {32'hbfbffae9, 32'hbe670592} /* (5, 30, 19) {real, imag} */,
  {32'h400ff890, 32'hc017f52d} /* (5, 30, 18) {real, imag} */,
  {32'h3f1eebc2, 32'h3e96032d} /* (5, 30, 17) {real, imag} */,
  {32'h3ee1cc05, 32'h3f6279c4} /* (5, 30, 16) {real, imag} */,
  {32'hbf3da239, 32'hbfdb4bd5} /* (5, 30, 15) {real, imag} */,
  {32'h3f5c026b, 32'h3fdb7718} /* (5, 30, 14) {real, imag} */,
  {32'h3e98d62b, 32'h3fe45646} /* (5, 30, 13) {real, imag} */,
  {32'h3f52c271, 32'hbe40a0eb} /* (5, 30, 12) {real, imag} */,
  {32'h3fbe1424, 32'h400aa8dc} /* (5, 30, 11) {real, imag} */,
  {32'h3f6e2f07, 32'h3e807e23} /* (5, 30, 10) {real, imag} */,
  {32'h408144c1, 32'h4026f217} /* (5, 30, 9) {real, imag} */,
  {32'h409ae812, 32'h3d72b0d9} /* (5, 30, 8) {real, imag} */,
  {32'hc0c699f9, 32'hbfd28b11} /* (5, 30, 7) {real, imag} */,
  {32'h40c4968c, 32'hbf73ad20} /* (5, 30, 6) {real, imag} */,
  {32'h402c482e, 32'hbf94c0cc} /* (5, 30, 5) {real, imag} */,
  {32'hc0f8113a, 32'h3faa624d} /* (5, 30, 4) {real, imag} */,
  {32'hc10b551f, 32'h40c6d987} /* (5, 30, 3) {real, imag} */,
  {32'h41162c06, 32'hc158debb} /* (5, 30, 2) {real, imag} */,
  {32'hc1a82d7f, 32'h41c7bc0f} /* (5, 30, 1) {real, imag} */,
  {32'h408f6436, 32'h41d11684} /* (5, 30, 0) {real, imag} */,
  {32'hc0568e65, 32'hc0c03f11} /* (5, 29, 31) {real, imag} */,
  {32'h40bceed7, 32'h4098f1f8} /* (5, 29, 30) {real, imag} */,
  {32'h3ee62d79, 32'h3ebee5d6} /* (5, 29, 29) {real, imag} */,
  {32'hc0593fcc, 32'hbf376669} /* (5, 29, 28) {real, imag} */,
  {32'hbeb857db, 32'hc06bee5c} /* (5, 29, 27) {real, imag} */,
  {32'h409c0eea, 32'h40a6b752} /* (5, 29, 26) {real, imag} */,
  {32'hc01f906b, 32'hc0ba0525} /* (5, 29, 25) {real, imag} */,
  {32'hbfed8ecc, 32'h40253476} /* (5, 29, 24) {real, imag} */,
  {32'hbe95d50a, 32'h40840704} /* (5, 29, 23) {real, imag} */,
  {32'hbfa37384, 32'h3f537098} /* (5, 29, 22) {real, imag} */,
  {32'h3ec3eef8, 32'hbf5a83fb} /* (5, 29, 21) {real, imag} */,
  {32'h3fab9341, 32'hc072a760} /* (5, 29, 20) {real, imag} */,
  {32'hbdc33c44, 32'h3fc9ed6c} /* (5, 29, 19) {real, imag} */,
  {32'hbff6e634, 32'h3f6cb042} /* (5, 29, 18) {real, imag} */,
  {32'hbfb13587, 32'h3f9ffe99} /* (5, 29, 17) {real, imag} */,
  {32'hbf1179e7, 32'hbf486f0e} /* (5, 29, 16) {real, imag} */,
  {32'h3fcedf2a, 32'hbeccac7f} /* (5, 29, 15) {real, imag} */,
  {32'h4002a637, 32'h3fa0c9f3} /* (5, 29, 14) {real, imag} */,
  {32'h3fb75ce3, 32'hbffd8a3e} /* (5, 29, 13) {real, imag} */,
  {32'hbffcdf3b, 32'h3f1257e2} /* (5, 29, 12) {real, imag} */,
  {32'h3de76713, 32'hbf3fcdbe} /* (5, 29, 11) {real, imag} */,
  {32'hc069cb85, 32'hbfec087f} /* (5, 29, 10) {real, imag} */,
  {32'h4064cb4c, 32'hbf0ed7ff} /* (5, 29, 9) {real, imag} */,
  {32'h4052654c, 32'h40b6088c} /* (5, 29, 8) {real, imag} */,
  {32'h3fc8e2c0, 32'h401fca64} /* (5, 29, 7) {real, imag} */,
  {32'hc06b7706, 32'hbfc648d3} /* (5, 29, 6) {real, imag} */,
  {32'hc057d16d, 32'h4099f7ff} /* (5, 29, 5) {real, imag} */,
  {32'h408c3375, 32'hc099fe23} /* (5, 29, 4) {real, imag} */,
  {32'h40408634, 32'h3fc1ad07} /* (5, 29, 3) {real, imag} */,
  {32'h4125b26e, 32'hc0a16882} /* (5, 29, 2) {real, imag} */,
  {32'hc166aef6, 32'h40414338} /* (5, 29, 1) {real, imag} */,
  {32'h40c7d274, 32'hc0e61689} /* (5, 29, 0) {real, imag} */,
  {32'hbdd0dbce, 32'hc148be4f} /* (5, 28, 31) {real, imag} */,
  {32'hc0b2ce47, 32'h410f0c40} /* (5, 28, 30) {real, imag} */,
  {32'hbfefce2f, 32'h40691709} /* (5, 28, 29) {real, imag} */,
  {32'hbe6709e5, 32'hbfc4be96} /* (5, 28, 28) {real, imag} */,
  {32'h400c33ef, 32'h400a9010} /* (5, 28, 27) {real, imag} */,
  {32'h3f217938, 32'hc0b5d367} /* (5, 28, 26) {real, imag} */,
  {32'h3f588417, 32'h3d366576} /* (5, 28, 25) {real, imag} */,
  {32'h3f09d70c, 32'hbf894a95} /* (5, 28, 24) {real, imag} */,
  {32'h4020881a, 32'hbfb9f7c4} /* (5, 28, 23) {real, imag} */,
  {32'hc0277fba, 32'h3d9492cd} /* (5, 28, 22) {real, imag} */,
  {32'hbfd88994, 32'hbf9e343f} /* (5, 28, 21) {real, imag} */,
  {32'h3d58b60f, 32'hbf949e16} /* (5, 28, 20) {real, imag} */,
  {32'h3f4fb661, 32'hbd790902} /* (5, 28, 19) {real, imag} */,
  {32'hbedf2730, 32'h40387066} /* (5, 28, 18) {real, imag} */,
  {32'hbf586f08, 32'h3ff66f32} /* (5, 28, 17) {real, imag} */,
  {32'h3f2e4e5d, 32'hbfec6afd} /* (5, 28, 16) {real, imag} */,
  {32'h4008ceb7, 32'h3d1ecb70} /* (5, 28, 15) {real, imag} */,
  {32'hbf6df517, 32'hbf1c8534} /* (5, 28, 14) {real, imag} */,
  {32'hbf1b8849, 32'h4004eb2a} /* (5, 28, 13) {real, imag} */,
  {32'hbfb824da, 32'h3f5900cf} /* (5, 28, 12) {real, imag} */,
  {32'h3d5de636, 32'hbe9f9b6d} /* (5, 28, 11) {real, imag} */,
  {32'h40459902, 32'hbfd1c407} /* (5, 28, 10) {real, imag} */,
  {32'hbf60b185, 32'h40376772} /* (5, 28, 9) {real, imag} */,
  {32'hc0469bcb, 32'h40386780} /* (5, 28, 8) {real, imag} */,
  {32'h3f3acb9e, 32'hc030dfde} /* (5, 28, 7) {real, imag} */,
  {32'hc01add25, 32'h402bb02e} /* (5, 28, 6) {real, imag} */,
  {32'hbf00df38, 32'h3fdcec75} /* (5, 28, 5) {real, imag} */,
  {32'hc0200b31, 32'hc0c356a9} /* (5, 28, 4) {real, imag} */,
  {32'h3f8742c5, 32'h4097b284} /* (5, 28, 3) {real, imag} */,
  {32'h408fa855, 32'h409a1b25} /* (5, 28, 2) {real, imag} */,
  {32'hc107038a, 32'hc09d7308} /* (5, 28, 1) {real, imag} */,
  {32'h4033948a, 32'h40bef1c9} /* (5, 28, 0) {real, imag} */,
  {32'hc11ac09a, 32'h40fc55fb} /* (5, 27, 31) {real, imag} */,
  {32'hbf90a631, 32'hc023b676} /* (5, 27, 30) {real, imag} */,
  {32'h3fb4ad8d, 32'h3f4e50af} /* (5, 27, 29) {real, imag} */,
  {32'h3ea3e1e5, 32'h3f306ac2} /* (5, 27, 28) {real, imag} */,
  {32'h400f7287, 32'hc064ae49} /* (5, 27, 27) {real, imag} */,
  {32'hbf075d88, 32'hc08f49a9} /* (5, 27, 26) {real, imag} */,
  {32'h3fdaf5f4, 32'h40001acf} /* (5, 27, 25) {real, imag} */,
  {32'hbf11f288, 32'h406e393d} /* (5, 27, 24) {real, imag} */,
  {32'h3f8d666e, 32'hbfc54d96} /* (5, 27, 23) {real, imag} */,
  {32'h40028719, 32'hc04b8737} /* (5, 27, 22) {real, imag} */,
  {32'h3f01d9ad, 32'hbaa9764a} /* (5, 27, 21) {real, imag} */,
  {32'h40265e21, 32'h4063ac2b} /* (5, 27, 20) {real, imag} */,
  {32'h3e5dffe2, 32'hbfe6923d} /* (5, 27, 19) {real, imag} */,
  {32'hc002687f, 32'h3e81e47a} /* (5, 27, 18) {real, imag} */,
  {32'hbf9815e2, 32'h3d3c0c47} /* (5, 27, 17) {real, imag} */,
  {32'h3fc2b545, 32'h3f8274f3} /* (5, 27, 16) {real, imag} */,
  {32'h3f627bb8, 32'hbf154524} /* (5, 27, 15) {real, imag} */,
  {32'h3fc87c99, 32'hbff4d531} /* (5, 27, 14) {real, imag} */,
  {32'h3f4ae9e3, 32'h3ecbe975} /* (5, 27, 13) {real, imag} */,
  {32'h3fe3e395, 32'h3f530f71} /* (5, 27, 12) {real, imag} */,
  {32'h3ecd6be8, 32'hbf0888ac} /* (5, 27, 11) {real, imag} */,
  {32'h3f38dd2c, 32'hbea246a1} /* (5, 27, 10) {real, imag} */,
  {32'hc0221747, 32'hbf967fd6} /* (5, 27, 9) {real, imag} */,
  {32'hbf6bb8d8, 32'h3e0c72fc} /* (5, 27, 8) {real, imag} */,
  {32'hbef1bdb8, 32'h403f7d86} /* (5, 27, 7) {real, imag} */,
  {32'h3fbd669f, 32'h40017847} /* (5, 27, 6) {real, imag} */,
  {32'h40a64ae3, 32'h3f645568} /* (5, 27, 5) {real, imag} */,
  {32'hbec4796c, 32'hc006750a} /* (5, 27, 4) {real, imag} */,
  {32'hc09e9e35, 32'hc08b27d3} /* (5, 27, 3) {real, imag} */,
  {32'h40e04304, 32'hc0caa814} /* (5, 27, 2) {real, imag} */,
  {32'h402e0763, 32'h40e47694} /* (5, 27, 1) {real, imag} */,
  {32'hc09603b5, 32'h402a6ebb} /* (5, 27, 0) {real, imag} */,
  {32'hc0a71829, 32'h3fe58fd8} /* (5, 26, 31) {real, imag} */,
  {32'h3f2015d5, 32'hbcb9a8cd} /* (5, 26, 30) {real, imag} */,
  {32'h3fcb9bf1, 32'hbfd1e184} /* (5, 26, 29) {real, imag} */,
  {32'hbfad30ee, 32'h3fd4e0b6} /* (5, 26, 28) {real, imag} */,
  {32'h3f46fcec, 32'h4082aee8} /* (5, 26, 27) {real, imag} */,
  {32'h3faba6b1, 32'h40618351} /* (5, 26, 26) {real, imag} */,
  {32'hbf983560, 32'h40245e4e} /* (5, 26, 25) {real, imag} */,
  {32'h405607b1, 32'hc0ac1ec9} /* (5, 26, 24) {real, imag} */,
  {32'hc0882f43, 32'hbe1a63f7} /* (5, 26, 23) {real, imag} */,
  {32'hbe93be9a, 32'hbf5afcac} /* (5, 26, 22) {real, imag} */,
  {32'h401f3757, 32'hbfbe0315} /* (5, 26, 21) {real, imag} */,
  {32'hc01845d5, 32'h3f899229} /* (5, 26, 20) {real, imag} */,
  {32'h3d4d75b2, 32'h3f68b209} /* (5, 26, 19) {real, imag} */,
  {32'hbf6d01c5, 32'h404d98aa} /* (5, 26, 18) {real, imag} */,
  {32'h3fd9cd71, 32'hbfdfab86} /* (5, 26, 17) {real, imag} */,
  {32'h3f19bf7c, 32'h3f20c466} /* (5, 26, 16) {real, imag} */,
  {32'hbfb75c59, 32'h3fd77077} /* (5, 26, 15) {real, imag} */,
  {32'hbed9f72d, 32'h3f52516b} /* (5, 26, 14) {real, imag} */,
  {32'h3f8cf68e, 32'h3f89c0ae} /* (5, 26, 13) {real, imag} */,
  {32'h3f8e30b4, 32'h3e9ca189} /* (5, 26, 12) {real, imag} */,
  {32'hbf91532d, 32'hbdecd91e} /* (5, 26, 11) {real, imag} */,
  {32'h40846292, 32'hbf8e5ae1} /* (5, 26, 10) {real, imag} */,
  {32'hbff40f35, 32'hbda50418} /* (5, 26, 9) {real, imag} */,
  {32'hbf81ccc7, 32'h3f82fd5b} /* (5, 26, 8) {real, imag} */,
  {32'h3fd94627, 32'h4081368e} /* (5, 26, 7) {real, imag} */,
  {32'h40437847, 32'hc025f2d6} /* (5, 26, 6) {real, imag} */,
  {32'h40ddab85, 32'hbf52dc1c} /* (5, 26, 5) {real, imag} */,
  {32'h4026d152, 32'h3e8d984f} /* (5, 26, 4) {real, imag} */,
  {32'hc096f727, 32'h3edb3d77} /* (5, 26, 3) {real, imag} */,
  {32'hc02e3f92, 32'hbf2342c0} /* (5, 26, 2) {real, imag} */,
  {32'hc0bb4b55, 32'h4081f36d} /* (5, 26, 1) {real, imag} */,
  {32'h3f9b8565, 32'h40b65cb7} /* (5, 26, 0) {real, imag} */,
  {32'hbfc4b3da, 32'hc086646e} /* (5, 25, 31) {real, imag} */,
  {32'h40a3b2ba, 32'h404ef264} /* (5, 25, 30) {real, imag} */,
  {32'h3fed553e, 32'hc029dcf3} /* (5, 25, 29) {real, imag} */,
  {32'h3fd34ece, 32'h40006f9f} /* (5, 25, 28) {real, imag} */,
  {32'h3f2f0650, 32'hc0083c63} /* (5, 25, 27) {real, imag} */,
  {32'hbfae8b6e, 32'h3ed81cad} /* (5, 25, 26) {real, imag} */,
  {32'hc0169c4f, 32'h3e07855a} /* (5, 25, 25) {real, imag} */,
  {32'h3fa3b06d, 32'h3f9bd9e7} /* (5, 25, 24) {real, imag} */,
  {32'h3bd5b41d, 32'h3e8c52b9} /* (5, 25, 23) {real, imag} */,
  {32'hbf3bc1c1, 32'h3d075f86} /* (5, 25, 22) {real, imag} */,
  {32'hbf2ab465, 32'h401de006} /* (5, 25, 21) {real, imag} */,
  {32'h3fd7be94, 32'h3fb70916} /* (5, 25, 20) {real, imag} */,
  {32'h3fafde29, 32'hbe4b4162} /* (5, 25, 19) {real, imag} */,
  {32'h3fe1e8fe, 32'hbfa42c9b} /* (5, 25, 18) {real, imag} */,
  {32'h3fb60222, 32'hbff66af9} /* (5, 25, 17) {real, imag} */,
  {32'hc05751a2, 32'hbdfdc26e} /* (5, 25, 16) {real, imag} */,
  {32'h3d4c65fa, 32'hc01656d2} /* (5, 25, 15) {real, imag} */,
  {32'h3e6a62ff, 32'h3c698fbc} /* (5, 25, 14) {real, imag} */,
  {32'hbfa8aa49, 32'hc041f33f} /* (5, 25, 13) {real, imag} */,
  {32'h400b12c9, 32'hc00a363e} /* (5, 25, 12) {real, imag} */,
  {32'h40119f08, 32'h40548cba} /* (5, 25, 11) {real, imag} */,
  {32'hbee8f595, 32'hbfaf993a} /* (5, 25, 10) {real, imag} */,
  {32'h3f5c08a1, 32'h3fb952a5} /* (5, 25, 9) {real, imag} */,
  {32'h404d0c11, 32'h3f73713d} /* (5, 25, 8) {real, imag} */,
  {32'hc0214c0c, 32'h3f5e018f} /* (5, 25, 7) {real, imag} */,
  {32'hc0053779, 32'h3e882c43} /* (5, 25, 6) {real, imag} */,
  {32'hbbb0cb30, 32'h4006984c} /* (5, 25, 5) {real, imag} */,
  {32'hbf3e9330, 32'hc021d07b} /* (5, 25, 4) {real, imag} */,
  {32'h4018f901, 32'h4017b318} /* (5, 25, 3) {real, imag} */,
  {32'h40ad7551, 32'h3f05d6b1} /* (5, 25, 2) {real, imag} */,
  {32'h3eeed053, 32'h403c1047} /* (5, 25, 1) {real, imag} */,
  {32'hc0020a27, 32'hc080b46c} /* (5, 25, 0) {real, imag} */,
  {32'hbe788339, 32'h3e67282a} /* (5, 24, 31) {real, imag} */,
  {32'h3fe11007, 32'hc0067ed2} /* (5, 24, 30) {real, imag} */,
  {32'hc02440a0, 32'hc058e83f} /* (5, 24, 29) {real, imag} */,
  {32'hc0154ed6, 32'h3f7d92c0} /* (5, 24, 28) {real, imag} */,
  {32'hbf9a6e9e, 32'h3f31b8a3} /* (5, 24, 27) {real, imag} */,
  {32'h404b2687, 32'h4052268c} /* (5, 24, 26) {real, imag} */,
  {32'hc0380f4a, 32'hbd25b993} /* (5, 24, 25) {real, imag} */,
  {32'hbfce4d9f, 32'hbf787213} /* (5, 24, 24) {real, imag} */,
  {32'hbfd5a14b, 32'h3fe75ba6} /* (5, 24, 23) {real, imag} */,
  {32'hc08487ff, 32'h406251f1} /* (5, 24, 22) {real, imag} */,
  {32'h40a48e5a, 32'hbfa562e8} /* (5, 24, 21) {real, imag} */,
  {32'h4011a9e5, 32'h40054996} /* (5, 24, 20) {real, imag} */,
  {32'h3f306094, 32'h3f37a66b} /* (5, 24, 19) {real, imag} */,
  {32'hbe235597, 32'h3f0132f4} /* (5, 24, 18) {real, imag} */,
  {32'h40039008, 32'h3f328b9a} /* (5, 24, 17) {real, imag} */,
  {32'hbfd6e331, 32'hbe510f03} /* (5, 24, 16) {real, imag} */,
  {32'hbf9441cb, 32'hbed41270} /* (5, 24, 15) {real, imag} */,
  {32'hbf0c2630, 32'h3f3c2ac0} /* (5, 24, 14) {real, imag} */,
  {32'h3fa1e5d6, 32'hbf9f3a02} /* (5, 24, 13) {real, imag} */,
  {32'hc01ff298, 32'h3fa3cac9} /* (5, 24, 12) {real, imag} */,
  {32'hbda298e0, 32'h3f2ff646} /* (5, 24, 11) {real, imag} */,
  {32'hbeca444a, 32'hbfbb2755} /* (5, 24, 10) {real, imag} */,
  {32'h40125a82, 32'hbf455dc4} /* (5, 24, 9) {real, imag} */,
  {32'h409b4674, 32'hc02d7a92} /* (5, 24, 8) {real, imag} */,
  {32'hbe7d66ea, 32'h3fb5af90} /* (5, 24, 7) {real, imag} */,
  {32'hbf1d3044, 32'hbff8701f} /* (5, 24, 6) {real, imag} */,
  {32'h408564d6, 32'h3f84a23e} /* (5, 24, 5) {real, imag} */,
  {32'hc04e51e0, 32'hc02ad5c7} /* (5, 24, 4) {real, imag} */,
  {32'h40abb0cd, 32'hbf78abd3} /* (5, 24, 3) {real, imag} */,
  {32'hbf4f1e09, 32'hc0474cc4} /* (5, 24, 2) {real, imag} */,
  {32'h3fb3496f, 32'h40e3aac5} /* (5, 24, 1) {real, imag} */,
  {32'h3ef4ce51, 32'h407c5a6d} /* (5, 24, 0) {real, imag} */,
  {32'h3ec7d51a, 32'h3cdd3235} /* (5, 23, 31) {real, imag} */,
  {32'hbf532417, 32'hc01bdff9} /* (5, 23, 30) {real, imag} */,
  {32'hbf23b245, 32'h4083808a} /* (5, 23, 29) {real, imag} */,
  {32'hc04b0959, 32'hbee3ad60} /* (5, 23, 28) {real, imag} */,
  {32'h40882a84, 32'hc030df36} /* (5, 23, 27) {real, imag} */,
  {32'h3f44b2fa, 32'h3ffdaa94} /* (5, 23, 26) {real, imag} */,
  {32'hbfd85180, 32'h3f77d8d2} /* (5, 23, 25) {real, imag} */,
  {32'hbfb44cd8, 32'h3f471c6b} /* (5, 23, 24) {real, imag} */,
  {32'hbfaa981b, 32'hc016483c} /* (5, 23, 23) {real, imag} */,
  {32'hbe406c9c, 32'h3f6f3394} /* (5, 23, 22) {real, imag} */,
  {32'hbec6535d, 32'hc08a14b7} /* (5, 23, 21) {real, imag} */,
  {32'hbfcc486b, 32'hbeeae6ae} /* (5, 23, 20) {real, imag} */,
  {32'h401193df, 32'hbf92e5af} /* (5, 23, 19) {real, imag} */,
  {32'h3fe0369c, 32'h3f3911ef} /* (5, 23, 18) {real, imag} */,
  {32'hbf062c23, 32'h3ff8cc56} /* (5, 23, 17) {real, imag} */,
  {32'hc09056ce, 32'hbf6b4aa8} /* (5, 23, 16) {real, imag} */,
  {32'h40905394, 32'hbf85a276} /* (5, 23, 15) {real, imag} */,
  {32'hbf44332c, 32'h3f266de2} /* (5, 23, 14) {real, imag} */,
  {32'h3f705267, 32'hbfa00a1e} /* (5, 23, 13) {real, imag} */,
  {32'h3f9cb88f, 32'hbf088a0c} /* (5, 23, 12) {real, imag} */,
  {32'hc0453144, 32'h3ffeb768} /* (5, 23, 11) {real, imag} */,
  {32'h3f502d83, 32'hbe8563ee} /* (5, 23, 10) {real, imag} */,
  {32'h4028d329, 32'hbfc651ea} /* (5, 23, 9) {real, imag} */,
  {32'h3f942f7e, 32'h400020de} /* (5, 23, 8) {real, imag} */,
  {32'h4017a41c, 32'hc00bda81} /* (5, 23, 7) {real, imag} */,
  {32'hc05027b7, 32'h408230ce} /* (5, 23, 6) {real, imag} */,
  {32'hbf202c70, 32'h4053a9a6} /* (5, 23, 5) {real, imag} */,
  {32'hc0032d92, 32'h4078ea99} /* (5, 23, 4) {real, imag} */,
  {32'h401c687a, 32'hbe41c2a0} /* (5, 23, 3) {real, imag} */,
  {32'h3fc644ec, 32'hc0553d71} /* (5, 23, 2) {real, imag} */,
  {32'hbfe24110, 32'hc002e75b} /* (5, 23, 1) {real, imag} */,
  {32'hbf16f9e4, 32'hbf181959} /* (5, 23, 0) {real, imag} */,
  {32'h4070e1c2, 32'hc041a511} /* (5, 22, 31) {real, imag} */,
  {32'hc045f8eb, 32'h404bb80e} /* (5, 22, 30) {real, imag} */,
  {32'hc04f1fe4, 32'hc07ebaca} /* (5, 22, 29) {real, imag} */,
  {32'hbf45891e, 32'hc00b2fa3} /* (5, 22, 28) {real, imag} */,
  {32'h3f6e1fc0, 32'h3f3c50cf} /* (5, 22, 27) {real, imag} */,
  {32'hc05314f3, 32'h3f2a4d29} /* (5, 22, 26) {real, imag} */,
  {32'h40826f7e, 32'hbfee9773} /* (5, 22, 25) {real, imag} */,
  {32'hbf179172, 32'h4013f253} /* (5, 22, 24) {real, imag} */,
  {32'h3f0fac16, 32'hbdcb4e38} /* (5, 22, 23) {real, imag} */,
  {32'hbe7cd5b5, 32'hbeeaf798} /* (5, 22, 22) {real, imag} */,
  {32'h40018e37, 32'h3fa66817} /* (5, 22, 21) {real, imag} */,
  {32'hc06d6841, 32'h3f3c72b5} /* (5, 22, 20) {real, imag} */,
  {32'h3ff82404, 32'h3f1c13a9} /* (5, 22, 19) {real, imag} */,
  {32'h3f306f3a, 32'hbea2eab7} /* (5, 22, 18) {real, imag} */,
  {32'h3c54781e, 32'hbfb38557} /* (5, 22, 17) {real, imag} */,
  {32'hbe0ac5f7, 32'hbee5adf6} /* (5, 22, 16) {real, imag} */,
  {32'h3f943218, 32'h403f2a7e} /* (5, 22, 15) {real, imag} */,
  {32'hbea7dff0, 32'h3edfcad1} /* (5, 22, 14) {real, imag} */,
  {32'h3e21e46c, 32'hbf9feadb} /* (5, 22, 13) {real, imag} */,
  {32'h3f7530c5, 32'hbf7f6d4b} /* (5, 22, 12) {real, imag} */,
  {32'hbe349673, 32'hc03b1da1} /* (5, 22, 11) {real, imag} */,
  {32'h40346a3f, 32'h4006702d} /* (5, 22, 10) {real, imag} */,
  {32'hbf759a5e, 32'hc0093e0c} /* (5, 22, 9) {real, imag} */,
  {32'hc002424f, 32'hbf636df5} /* (5, 22, 8) {real, imag} */,
  {32'h3fbf170e, 32'h4022114a} /* (5, 22, 7) {real, imag} */,
  {32'hbfb0461a, 32'h3e36d040} /* (5, 22, 6) {real, imag} */,
  {32'h40291ab7, 32'h3f300d66} /* (5, 22, 5) {real, imag} */,
  {32'h3fd9b4ae, 32'h3fb12229} /* (5, 22, 4) {real, imag} */,
  {32'hbfdf3c7b, 32'h3f299875} /* (5, 22, 3) {real, imag} */,
  {32'hbe2e4f19, 32'h3fbfe55a} /* (5, 22, 2) {real, imag} */,
  {32'hc046147a, 32'hbfd58e0a} /* (5, 22, 1) {real, imag} */,
  {32'hbff015df, 32'hc0268bc1} /* (5, 22, 0) {real, imag} */,
  {32'h3fab1855, 32'h3dea4e0c} /* (5, 21, 31) {real, imag} */,
  {32'hbf8e85de, 32'h3fda826f} /* (5, 21, 30) {real, imag} */,
  {32'h3f8bc9ee, 32'h3fa7b1ca} /* (5, 21, 29) {real, imag} */,
  {32'h409ea013, 32'h3f00c09f} /* (5, 21, 28) {real, imag} */,
  {32'hc009222b, 32'h3f284b67} /* (5, 21, 27) {real, imag} */,
  {32'h3f64ccad, 32'hbcf147bb} /* (5, 21, 26) {real, imag} */,
  {32'h3f1f8b64, 32'h3dcb4795} /* (5, 21, 25) {real, imag} */,
  {32'hbf80ac3a, 32'hbed259d9} /* (5, 21, 24) {real, imag} */,
  {32'h3ebf331c, 32'h40301d27} /* (5, 21, 23) {real, imag} */,
  {32'hc0535fce, 32'h4055ea4f} /* (5, 21, 22) {real, imag} */,
  {32'h3ef763fd, 32'h4023d47a} /* (5, 21, 21) {real, imag} */,
  {32'hc0180ddc, 32'hbe628dcc} /* (5, 21, 20) {real, imag} */,
  {32'hbf9c5260, 32'h402e9ae5} /* (5, 21, 19) {real, imag} */,
  {32'hbf893eeb, 32'hc00b5439} /* (5, 21, 18) {real, imag} */,
  {32'hbf38874f, 32'hc0132243} /* (5, 21, 17) {real, imag} */,
  {32'hbe0aaa25, 32'h401cb5e9} /* (5, 21, 16) {real, imag} */,
  {32'hbf90a454, 32'h3d12eea5} /* (5, 21, 15) {real, imag} */,
  {32'h404361ca, 32'hbfa56707} /* (5, 21, 14) {real, imag} */,
  {32'h40374aab, 32'h3fe0200a} /* (5, 21, 13) {real, imag} */,
  {32'h3ef47941, 32'hbe1503a8} /* (5, 21, 12) {real, imag} */,
  {32'h3f808ba7, 32'hbfeee766} /* (5, 21, 11) {real, imag} */,
  {32'hbf32661f, 32'hbeeebbfe} /* (5, 21, 10) {real, imag} */,
  {32'h3f835bf0, 32'hbfe13111} /* (5, 21, 9) {real, imag} */,
  {32'hbd925911, 32'hc007e676} /* (5, 21, 8) {real, imag} */,
  {32'h3d16777c, 32'h4091ea22} /* (5, 21, 7) {real, imag} */,
  {32'hbe125a4e, 32'hbf4e80b6} /* (5, 21, 6) {real, imag} */,
  {32'hbf8e103d, 32'hc084e02b} /* (5, 21, 5) {real, imag} */,
  {32'hbfa41bf3, 32'h40249dd5} /* (5, 21, 4) {real, imag} */,
  {32'h3f60776d, 32'h3eb71427} /* (5, 21, 3) {real, imag} */,
  {32'hbf04d3d9, 32'h3f9805c1} /* (5, 21, 2) {real, imag} */,
  {32'hbd4f2ca0, 32'h404d1ce8} /* (5, 21, 1) {real, imag} */,
  {32'h3f8239f4, 32'h4065110e} /* (5, 21, 0) {real, imag} */,
  {32'h3fec3568, 32'hbfede6dc} /* (5, 20, 31) {real, imag} */,
  {32'h3f017388, 32'hbfb20dcf} /* (5, 20, 30) {real, imag} */,
  {32'hbf771c42, 32'h3f047229} /* (5, 20, 29) {real, imag} */,
  {32'h4011dacd, 32'hbfc7fb4b} /* (5, 20, 28) {real, imag} */,
  {32'hc031db2d, 32'hc016cefd} /* (5, 20, 27) {real, imag} */,
  {32'hc043896a, 32'h3b1057d2} /* (5, 20, 26) {real, imag} */,
  {32'h3c96aae1, 32'h3e7cc52b} /* (5, 20, 25) {real, imag} */,
  {32'h3f8ba5a8, 32'h3f24c5f9} /* (5, 20, 24) {real, imag} */,
  {32'hbf64a03b, 32'hc02d76cb} /* (5, 20, 23) {real, imag} */,
  {32'h3f5b9abb, 32'hc0441966} /* (5, 20, 22) {real, imag} */,
  {32'hbecbf366, 32'hbf8c0ae2} /* (5, 20, 21) {real, imag} */,
  {32'h3f99093f, 32'h4046d039} /* (5, 20, 20) {real, imag} */,
  {32'hbf9a1caa, 32'hbe8e85bd} /* (5, 20, 19) {real, imag} */,
  {32'hbeb3db66, 32'h3f188428} /* (5, 20, 18) {real, imag} */,
  {32'h3f072c7e, 32'hbf3208a8} /* (5, 20, 17) {real, imag} */,
  {32'h3f1e630f, 32'h3f78794e} /* (5, 20, 16) {real, imag} */,
  {32'hbfbc7b50, 32'hbfa8037f} /* (5, 20, 15) {real, imag} */,
  {32'hc0102707, 32'h3f6ee016} /* (5, 20, 14) {real, imag} */,
  {32'hc017ba11, 32'hbf0c9d01} /* (5, 20, 13) {real, imag} */,
  {32'h3e8308d4, 32'h3cda7e9c} /* (5, 20, 12) {real, imag} */,
  {32'h3fde74b9, 32'hbff76a7d} /* (5, 20, 11) {real, imag} */,
  {32'hbfa5fc4a, 32'hbfb93d80} /* (5, 20, 10) {real, imag} */,
  {32'h40566376, 32'hbfb33bdb} /* (5, 20, 9) {real, imag} */,
  {32'hbed49f0a, 32'h3f0a6c4b} /* (5, 20, 8) {real, imag} */,
  {32'h3ee6b39a, 32'hc0647faf} /* (5, 20, 7) {real, imag} */,
  {32'h4018846c, 32'h3f4a4877} /* (5, 20, 6) {real, imag} */,
  {32'hbf766380, 32'hbff1e2fe} /* (5, 20, 5) {real, imag} */,
  {32'hc073cf27, 32'h4030c764} /* (5, 20, 4) {real, imag} */,
  {32'h3fed27ef, 32'h3f8c739c} /* (5, 20, 3) {real, imag} */,
  {32'hbe61dbdd, 32'h3e8b2bee} /* (5, 20, 2) {real, imag} */,
  {32'h3f6cb9fd, 32'hbff0a08c} /* (5, 20, 1) {real, imag} */,
  {32'h3fffa6b6, 32'hbf83da9b} /* (5, 20, 0) {real, imag} */,
  {32'hbec99177, 32'hbe987a26} /* (5, 19, 31) {real, imag} */,
  {32'h3f5355ca, 32'h3fb5206e} /* (5, 19, 30) {real, imag} */,
  {32'hbfc477c0, 32'hbf8da572} /* (5, 19, 29) {real, imag} */,
  {32'hbfe34d10, 32'hbed0cf67} /* (5, 19, 28) {real, imag} */,
  {32'h3fd84010, 32'hbfa13fca} /* (5, 19, 27) {real, imag} */,
  {32'hbfd699b0, 32'h3f8ff6ec} /* (5, 19, 26) {real, imag} */,
  {32'h40457e48, 32'hc024bd87} /* (5, 19, 25) {real, imag} */,
  {32'h3ef36f94, 32'hbd4cb3f6} /* (5, 19, 24) {real, imag} */,
  {32'h3fa88a6d, 32'hc0434a5f} /* (5, 19, 23) {real, imag} */,
  {32'h3f565a8a, 32'h3f4a1cd5} /* (5, 19, 22) {real, imag} */,
  {32'h40336db6, 32'hc0010629} /* (5, 19, 21) {real, imag} */,
  {32'hbeeb3d57, 32'hbe8a1290} /* (5, 19, 20) {real, imag} */,
  {32'h3f00d326, 32'h3fa659fa} /* (5, 19, 19) {real, imag} */,
  {32'hbfb04eb0, 32'h3edfe41b} /* (5, 19, 18) {real, imag} */,
  {32'hbf0fb343, 32'h4006bcbf} /* (5, 19, 17) {real, imag} */,
  {32'h3ff6ca54, 32'hbf84d977} /* (5, 19, 16) {real, imag} */,
  {32'hbfc6592c, 32'hbf691dc9} /* (5, 19, 15) {real, imag} */,
  {32'h3eebf40d, 32'h3fc430e3} /* (5, 19, 14) {real, imag} */,
  {32'h3f0df1be, 32'h40279810} /* (5, 19, 13) {real, imag} */,
  {32'hbec45608, 32'h3ff36cea} /* (5, 19, 12) {real, imag} */,
  {32'hc006e756, 32'h3e9a4d89} /* (5, 19, 11) {real, imag} */,
  {32'h402d6d13, 32'hbfaffebe} /* (5, 19, 10) {real, imag} */,
  {32'hbfff00f3, 32'h40004707} /* (5, 19, 9) {real, imag} */,
  {32'hc0199763, 32'hbf612b74} /* (5, 19, 8) {real, imag} */,
  {32'hbf4d9e14, 32'h3fa1cf32} /* (5, 19, 7) {real, imag} */,
  {32'h3ee30f62, 32'hbe317e98} /* (5, 19, 6) {real, imag} */,
  {32'hc08cfcd4, 32'hbf51fe2d} /* (5, 19, 5) {real, imag} */,
  {32'h403c642f, 32'h3ebac3d7} /* (5, 19, 4) {real, imag} */,
  {32'hbff8d255, 32'h3e403044} /* (5, 19, 3) {real, imag} */,
  {32'h3f0de3d6, 32'hbf339c2d} /* (5, 19, 2) {real, imag} */,
  {32'h3fc53417, 32'hbf2eddc6} /* (5, 19, 1) {real, imag} */,
  {32'hc00233ee, 32'hbe154b6e} /* (5, 19, 0) {real, imag} */,
  {32'hbec1d39b, 32'hbf677abd} /* (5, 18, 31) {real, imag} */,
  {32'h3c630062, 32'h406216cb} /* (5, 18, 30) {real, imag} */,
  {32'h3fa1b1ca, 32'hc04ed7bb} /* (5, 18, 29) {real, imag} */,
  {32'hbeff8478, 32'hbf1f2e1b} /* (5, 18, 28) {real, imag} */,
  {32'h3fdf4870, 32'hbc11d1b2} /* (5, 18, 27) {real, imag} */,
  {32'h3ef94f67, 32'h3eeac5e3} /* (5, 18, 26) {real, imag} */,
  {32'h3f895c5d, 32'hbedb605d} /* (5, 18, 25) {real, imag} */,
  {32'hbf1df981, 32'h3d2b3a26} /* (5, 18, 24) {real, imag} */,
  {32'hc02a7f1f, 32'h3f4637e7} /* (5, 18, 23) {real, imag} */,
  {32'h4085aabf, 32'hc01ebd1f} /* (5, 18, 22) {real, imag} */,
  {32'h3fd95279, 32'h3f583309} /* (5, 18, 21) {real, imag} */,
  {32'h3f6433ed, 32'hc0680cc3} /* (5, 18, 20) {real, imag} */,
  {32'h3fb11e7b, 32'h3f2f909e} /* (5, 18, 19) {real, imag} */,
  {32'hbf034b87, 32'h3ee92175} /* (5, 18, 18) {real, imag} */,
  {32'h3fa3687b, 32'hc0096edf} /* (5, 18, 17) {real, imag} */,
  {32'hbf13dc09, 32'hbe5093b3} /* (5, 18, 16) {real, imag} */,
  {32'h3f26bb51, 32'h3f55f0e5} /* (5, 18, 15) {real, imag} */,
  {32'hbfa15d40, 32'hbf05c707} /* (5, 18, 14) {real, imag} */,
  {32'h3f9392ec, 32'hbfb8035a} /* (5, 18, 13) {real, imag} */,
  {32'h3f35441c, 32'hc03e1220} /* (5, 18, 12) {real, imag} */,
  {32'h3fa5b91f, 32'hbca42698} /* (5, 18, 11) {real, imag} */,
  {32'h3f718fe8, 32'h406fe94e} /* (5, 18, 10) {real, imag} */,
  {32'h3f40d98f, 32'h3f2bcfd2} /* (5, 18, 9) {real, imag} */,
  {32'hbfc8f6ff, 32'h4007fae2} /* (5, 18, 8) {real, imag} */,
  {32'hc02d2c78, 32'hbf8b4d74} /* (5, 18, 7) {real, imag} */,
  {32'h401778ad, 32'hc029776e} /* (5, 18, 6) {real, imag} */,
  {32'hbefd831f, 32'hbe4bf915} /* (5, 18, 5) {real, imag} */,
  {32'hbf4cbbcf, 32'hc05017fb} /* (5, 18, 4) {real, imag} */,
  {32'h3f1ffd36, 32'hbf3793bf} /* (5, 18, 3) {real, imag} */,
  {32'hbf68fffc, 32'hbfd0de96} /* (5, 18, 2) {real, imag} */,
  {32'hbd2446c6, 32'h404b67f8} /* (5, 18, 1) {real, imag} */,
  {32'h3e9abafa, 32'h3f8bce1e} /* (5, 18, 0) {real, imag} */,
  {32'hbd8a66e3, 32'hc0031d5c} /* (5, 17, 31) {real, imag} */,
  {32'hbf0f7d1d, 32'hbfbdce1a} /* (5, 17, 30) {real, imag} */,
  {32'h3ee99e9c, 32'h3db37548} /* (5, 17, 29) {real, imag} */,
  {32'hbfae0b34, 32'h3f69fc8b} /* (5, 17, 28) {real, imag} */,
  {32'h406e160c, 32'h3e381dbe} /* (5, 17, 27) {real, imag} */,
  {32'hbfa46434, 32'h4010f8cc} /* (5, 17, 26) {real, imag} */,
  {32'hbfeb535f, 32'hbeeb29a9} /* (5, 17, 25) {real, imag} */,
  {32'h40098117, 32'hbf23d31e} /* (5, 17, 24) {real, imag} */,
  {32'hbf43dc07, 32'h3f80c5fd} /* (5, 17, 23) {real, imag} */,
  {32'h3f84d324, 32'hbf464d45} /* (5, 17, 22) {real, imag} */,
  {32'h3ea5ba1a, 32'hc0270535} /* (5, 17, 21) {real, imag} */,
  {32'hbdee3616, 32'h3f8a9baf} /* (5, 17, 20) {real, imag} */,
  {32'h3f68ec5f, 32'hbd60ed97} /* (5, 17, 19) {real, imag} */,
  {32'hbf3233b3, 32'h3c8fe803} /* (5, 17, 18) {real, imag} */,
  {32'hbeed27b9, 32'hbf076289} /* (5, 17, 17) {real, imag} */,
  {32'h3fc65ea4, 32'hbf8f236f} /* (5, 17, 16) {real, imag} */,
  {32'h3e407555, 32'h3da0f4e5} /* (5, 17, 15) {real, imag} */,
  {32'hc004ebae, 32'h401bf860} /* (5, 17, 14) {real, imag} */,
  {32'hbee89856, 32'h3fd10549} /* (5, 17, 13) {real, imag} */,
  {32'hbfa84386, 32'h3f133e6f} /* (5, 17, 12) {real, imag} */,
  {32'h3f0ecb66, 32'h3dad275e} /* (5, 17, 11) {real, imag} */,
  {32'hbfb0865f, 32'h3f79abde} /* (5, 17, 10) {real, imag} */,
  {32'hbf91aa07, 32'hbf5efc56} /* (5, 17, 9) {real, imag} */,
  {32'h3c840ad9, 32'h3d8f1982} /* (5, 17, 8) {real, imag} */,
  {32'hbfc41e23, 32'hbf1bb780} /* (5, 17, 7) {real, imag} */,
  {32'hbe94ae1f, 32'h3fbd9c14} /* (5, 17, 6) {real, imag} */,
  {32'h3dc4fe2e, 32'h3e782fc5} /* (5, 17, 5) {real, imag} */,
  {32'h3ea76196, 32'hbf3454c9} /* (5, 17, 4) {real, imag} */,
  {32'hbf131738, 32'h3ecee514} /* (5, 17, 3) {real, imag} */,
  {32'hbe0dfde1, 32'h3f3f53df} /* (5, 17, 2) {real, imag} */,
  {32'hc003050b, 32'h3e46e20e} /* (5, 17, 1) {real, imag} */,
  {32'h3cfd026f, 32'hbed856f7} /* (5, 17, 0) {real, imag} */,
  {32'h3d800434, 32'h3f18b804} /* (5, 16, 31) {real, imag} */,
  {32'h3881167f, 32'h3df0ab10} /* (5, 16, 30) {real, imag} */,
  {32'h3e3d0c71, 32'hbfa41233} /* (5, 16, 29) {real, imag} */,
  {32'hbf421cd5, 32'h3fa42fbd} /* (5, 16, 28) {real, imag} */,
  {32'h3d6d4a89, 32'h3f856c50} /* (5, 16, 27) {real, imag} */,
  {32'h3e523392, 32'hbdded9aa} /* (5, 16, 26) {real, imag} */,
  {32'h3f0816e6, 32'hbe52b0a0} /* (5, 16, 25) {real, imag} */,
  {32'hbe256b50, 32'h403644ac} /* (5, 16, 24) {real, imag} */,
  {32'hbd7b1d81, 32'h3dbc97da} /* (5, 16, 23) {real, imag} */,
  {32'h3fa2d87b, 32'hbf9a2c78} /* (5, 16, 22) {real, imag} */,
  {32'hbf70482f, 32'hbf7b03df} /* (5, 16, 21) {real, imag} */,
  {32'hc076b2ee, 32'h3f8a6c35} /* (5, 16, 20) {real, imag} */,
  {32'hc02e8748, 32'hbe172af4} /* (5, 16, 19) {real, imag} */,
  {32'h3ef7bf25, 32'h3ee23ad0} /* (5, 16, 18) {real, imag} */,
  {32'h3f11a220, 32'h3cbea816} /* (5, 16, 17) {real, imag} */,
  {32'hbf55ca0a, 32'hbfda67d5} /* (5, 16, 16) {real, imag} */,
  {32'hbd0dc93a, 32'hbf7f4540} /* (5, 16, 15) {real, imag} */,
  {32'hbf378ce3, 32'h3fa0da6e} /* (5, 16, 14) {real, imag} */,
  {32'h3f74bb90, 32'h3ebb313b} /* (5, 16, 13) {real, imag} */,
  {32'h3f3354fa, 32'h3e1cb779} /* (5, 16, 12) {real, imag} */,
  {32'h3fc5b3f1, 32'hbf88631c} /* (5, 16, 11) {real, imag} */,
  {32'hbf0b72f7, 32'hbfb5b82f} /* (5, 16, 10) {real, imag} */,
  {32'h3fcdafa5, 32'h3ff4bcbc} /* (5, 16, 9) {real, imag} */,
  {32'h3f16d58e, 32'hbf2ecbed} /* (5, 16, 8) {real, imag} */,
  {32'h3f462552, 32'h3f3540c3} /* (5, 16, 7) {real, imag} */,
  {32'hbf5220cb, 32'h3e3fec29} /* (5, 16, 6) {real, imag} */,
  {32'hbd803875, 32'h3e424207} /* (5, 16, 5) {real, imag} */,
  {32'h3e9ac01c, 32'hbeb448d7} /* (5, 16, 4) {real, imag} */,
  {32'hbe3f42da, 32'h3fb3e0e6} /* (5, 16, 3) {real, imag} */,
  {32'hbf6f8795, 32'hbf4f1682} /* (5, 16, 2) {real, imag} */,
  {32'hbf747d8b, 32'h3f4fe89b} /* (5, 16, 1) {real, imag} */,
  {32'h3f21364b, 32'h3b816a99} /* (5, 16, 0) {real, imag} */,
  {32'hbf1f4a4f, 32'hbefa6754} /* (5, 15, 31) {real, imag} */,
  {32'hbea57944, 32'h405748c3} /* (5, 15, 30) {real, imag} */,
  {32'h3c571ccc, 32'hbe714429} /* (5, 15, 29) {real, imag} */,
  {32'hbee080a4, 32'hbf266e4a} /* (5, 15, 28) {real, imag} */,
  {32'hc00ef763, 32'h3f2d0dcc} /* (5, 15, 27) {real, imag} */,
  {32'hbe72c29d, 32'h3f6386b5} /* (5, 15, 26) {real, imag} */,
  {32'hbfe0749c, 32'hbeea7c07} /* (5, 15, 25) {real, imag} */,
  {32'hc026de24, 32'hbe81d4b1} /* (5, 15, 24) {real, imag} */,
  {32'h3f7c5297, 32'h3e077448} /* (5, 15, 23) {real, imag} */,
  {32'h3fbd5660, 32'h3fe17856} /* (5, 15, 22) {real, imag} */,
  {32'h3ea4cc4a, 32'hbee74c0d} /* (5, 15, 21) {real, imag} */,
  {32'h3f29167c, 32'hbdc82eac} /* (5, 15, 20) {real, imag} */,
  {32'hc003eea9, 32'hbf7df29e} /* (5, 15, 19) {real, imag} */,
  {32'hbfdc3959, 32'hbe0a7f8f} /* (5, 15, 18) {real, imag} */,
  {32'h3fcddc9f, 32'hbfa6af97} /* (5, 15, 17) {real, imag} */,
  {32'hbf9e2443, 32'h4016650c} /* (5, 15, 16) {real, imag} */,
  {32'h3f505a21, 32'h3f63f3a4} /* (5, 15, 15) {real, imag} */,
  {32'h3e5c7b59, 32'h3fd90a45} /* (5, 15, 14) {real, imag} */,
  {32'h3f80c508, 32'h3fc231b9} /* (5, 15, 13) {real, imag} */,
  {32'hbf0bf606, 32'h403b39e3} /* (5, 15, 12) {real, imag} */,
  {32'h3edfe4c8, 32'h3f76ddc1} /* (5, 15, 11) {real, imag} */,
  {32'h40340cf0, 32'hbff90c07} /* (5, 15, 10) {real, imag} */,
  {32'hbe9651e6, 32'h3e9468b6} /* (5, 15, 9) {real, imag} */,
  {32'hc030d357, 32'h3d27467d} /* (5, 15, 8) {real, imag} */,
  {32'h3eedfe4a, 32'hbbb84b36} /* (5, 15, 7) {real, imag} */,
  {32'h3df30846, 32'hbf36a2cf} /* (5, 15, 6) {real, imag} */,
  {32'h3eb7008d, 32'h3f26e790} /* (5, 15, 5) {real, imag} */,
  {32'h3f3c26e5, 32'h3e748840} /* (5, 15, 4) {real, imag} */,
  {32'hbf28fd6b, 32'h3d43fc18} /* (5, 15, 3) {real, imag} */,
  {32'hbf822b48, 32'hbf12f6ac} /* (5, 15, 2) {real, imag} */,
  {32'h3fafb58e, 32'h3f11e280} /* (5, 15, 1) {real, imag} */,
  {32'h402cafd7, 32'h4063f311} /* (5, 15, 0) {real, imag} */,
  {32'hbf942db1, 32'h3eb29ac0} /* (5, 14, 31) {real, imag} */,
  {32'hbeb0cd0b, 32'h3ef222e8} /* (5, 14, 30) {real, imag} */,
  {32'hbfc1e97b, 32'h3f937552} /* (5, 14, 29) {real, imag} */,
  {32'hbf7c4ff5, 32'h3ed16666} /* (5, 14, 28) {real, imag} */,
  {32'hc04774cf, 32'hbefb3592} /* (5, 14, 27) {real, imag} */,
  {32'hc01df9ee, 32'h3f7054c6} /* (5, 14, 26) {real, imag} */,
  {32'hc03533a0, 32'hc02e4ff3} /* (5, 14, 25) {real, imag} */,
  {32'hbfac8f5b, 32'hbfd3bf51} /* (5, 14, 24) {real, imag} */,
  {32'h3f3f994b, 32'h3ff5d793} /* (5, 14, 23) {real, imag} */,
  {32'hbfefd602, 32'h3f6c0f28} /* (5, 14, 22) {real, imag} */,
  {32'h4014ce64, 32'hbf392ac0} /* (5, 14, 21) {real, imag} */,
  {32'h3d43a662, 32'hc00a4167} /* (5, 14, 20) {real, imag} */,
  {32'h3e8d1fcd, 32'hbe95c01e} /* (5, 14, 19) {real, imag} */,
  {32'h3ed9ea0d, 32'hbfdb0cc8} /* (5, 14, 18) {real, imag} */,
  {32'h3fcfeb1a, 32'hc02f3dcf} /* (5, 14, 17) {real, imag} */,
  {32'h3f40e3a9, 32'h3fd1ac27} /* (5, 14, 16) {real, imag} */,
  {32'hbf9bc091, 32'hbf269a77} /* (5, 14, 15) {real, imag} */,
  {32'h3ee50b9b, 32'hbfdd43a5} /* (5, 14, 14) {real, imag} */,
  {32'h3f9d8633, 32'h3fbe0e67} /* (5, 14, 13) {real, imag} */,
  {32'h40098b50, 32'hbfc17466} /* (5, 14, 12) {real, imag} */,
  {32'hc02d05d1, 32'hc02595b7} /* (5, 14, 11) {real, imag} */,
  {32'h3f9c9100, 32'h3fcd32cd} /* (5, 14, 10) {real, imag} */,
  {32'hbeba3c6c, 32'h403c90cc} /* (5, 14, 9) {real, imag} */,
  {32'h3fe8be4d, 32'h3f837988} /* (5, 14, 8) {real, imag} */,
  {32'hbebd436d, 32'h3fa7c023} /* (5, 14, 7) {real, imag} */,
  {32'h3ea59b4e, 32'h3fa64bd1} /* (5, 14, 6) {real, imag} */,
  {32'h3e08dec3, 32'h4019c64c} /* (5, 14, 5) {real, imag} */,
  {32'hc0162f48, 32'hbf97068e} /* (5, 14, 4) {real, imag} */,
  {32'h3f46f243, 32'hbeabd956} /* (5, 14, 3) {real, imag} */,
  {32'h40512989, 32'h3f93e7de} /* (5, 14, 2) {real, imag} */,
  {32'hc032010f, 32'h3f0fbe3a} /* (5, 14, 1) {real, imag} */,
  {32'h3f7647c4, 32'h3fbf52f9} /* (5, 14, 0) {real, imag} */,
  {32'h3e8a999b, 32'hbfda5709} /* (5, 13, 31) {real, imag} */,
  {32'hbe3ae9fc, 32'h3fba0139} /* (5, 13, 30) {real, imag} */,
  {32'h4028577e, 32'h3f772884} /* (5, 13, 29) {real, imag} */,
  {32'h3e3ada87, 32'hbf9f2377} /* (5, 13, 28) {real, imag} */,
  {32'hc0238465, 32'hbfc4aead} /* (5, 13, 27) {real, imag} */,
  {32'h4006cd13, 32'h3efcb7da} /* (5, 13, 26) {real, imag} */,
  {32'h3fd82137, 32'hc00f5e48} /* (5, 13, 25) {real, imag} */,
  {32'h3f179cb0, 32'hbea9b76a} /* (5, 13, 24) {real, imag} */,
  {32'hbfc96116, 32'hc05836e5} /* (5, 13, 23) {real, imag} */,
  {32'h3ff1c1b4, 32'h408ec3a7} /* (5, 13, 22) {real, imag} */,
  {32'hc01aa770, 32'h400f59bc} /* (5, 13, 21) {real, imag} */,
  {32'h3fe3f62c, 32'hbf013d3e} /* (5, 13, 20) {real, imag} */,
  {32'hbd62c332, 32'hbea56690} /* (5, 13, 19) {real, imag} */,
  {32'hbfb3ad3d, 32'h3fd32c24} /* (5, 13, 18) {real, imag} */,
  {32'h3f975547, 32'h3e9d70ce} /* (5, 13, 17) {real, imag} */,
  {32'h3da4954b, 32'hbee3a2ca} /* (5, 13, 16) {real, imag} */,
  {32'h3f09fecd, 32'h3f92e69c} /* (5, 13, 15) {real, imag} */,
  {32'hbf01c955, 32'hc09b55ad} /* (5, 13, 14) {real, imag} */,
  {32'hbfe4263f, 32'hbf8fb466} /* (5, 13, 13) {real, imag} */,
  {32'hbedc322c, 32'h3fcd0a86} /* (5, 13, 12) {real, imag} */,
  {32'h3f8a97dc, 32'h3f36b6db} /* (5, 13, 11) {real, imag} */,
  {32'h3d6d70a5, 32'hbf91bf6d} /* (5, 13, 10) {real, imag} */,
  {32'h3f98e492, 32'h3f005669} /* (5, 13, 9) {real, imag} */,
  {32'h3fb4c84a, 32'hc030b606} /* (5, 13, 8) {real, imag} */,
  {32'h3fad94e0, 32'h3e5707d1} /* (5, 13, 7) {real, imag} */,
  {32'hbfbf2f28, 32'h3fdaf5d3} /* (5, 13, 6) {real, imag} */,
  {32'h3fd4213e, 32'hbe1bc280} /* (5, 13, 5) {real, imag} */,
  {32'h3ecc0e99, 32'h3f020344} /* (5, 13, 4) {real, imag} */,
  {32'h4011aa42, 32'h3f640024} /* (5, 13, 3) {real, imag} */,
  {32'h3e74479b, 32'hbfa0795d} /* (5, 13, 2) {real, imag} */,
  {32'hbfad07e9, 32'h3f9c1afd} /* (5, 13, 1) {real, imag} */,
  {32'hc0087b36, 32'h40136a0c} /* (5, 13, 0) {real, imag} */,
  {32'hbfb9a7f7, 32'hbf3c284e} /* (5, 12, 31) {real, imag} */,
  {32'hbff82369, 32'hc0057cfb} /* (5, 12, 30) {real, imag} */,
  {32'hbf5b0193, 32'hbfe863aa} /* (5, 12, 29) {real, imag} */,
  {32'hbf8c6c8a, 32'hbfb1fafc} /* (5, 12, 28) {real, imag} */,
  {32'h400900bb, 32'h3faa7226} /* (5, 12, 27) {real, imag} */,
  {32'hbfa13b05, 32'h3fee11f9} /* (5, 12, 26) {real, imag} */,
  {32'h3ebff6b9, 32'h3fc718af} /* (5, 12, 25) {real, imag} */,
  {32'h4034fad4, 32'h3fd05d66} /* (5, 12, 24) {real, imag} */,
  {32'h3fd0fb73, 32'hc0018b83} /* (5, 12, 23) {real, imag} */,
  {32'hbfdf3f0c, 32'hbefd44dd} /* (5, 12, 22) {real, imag} */,
  {32'h3e95204c, 32'hc01f2b56} /* (5, 12, 21) {real, imag} */,
  {32'h3f862225, 32'h3d6527c5} /* (5, 12, 20) {real, imag} */,
  {32'h3f3ff40f, 32'h3f51d6c7} /* (5, 12, 19) {real, imag} */,
  {32'hbe6a2e64, 32'hbf8ae92c} /* (5, 12, 18) {real, imag} */,
  {32'h3f3ca4de, 32'h402e0353} /* (5, 12, 17) {real, imag} */,
  {32'h3ec41525, 32'hbecccb72} /* (5, 12, 16) {real, imag} */,
  {32'h3f0557b2, 32'h3df189f7} /* (5, 12, 15) {real, imag} */,
  {32'h3fd5ad9e, 32'h401835d3} /* (5, 12, 14) {real, imag} */,
  {32'h3c6b81df, 32'hbfe0cb13} /* (5, 12, 13) {real, imag} */,
  {32'hbfb74f4b, 32'hbe52b13f} /* (5, 12, 12) {real, imag} */,
  {32'hc0520705, 32'h3fd98205} /* (5, 12, 11) {real, imag} */,
  {32'h3ec00ed7, 32'hbf07758a} /* (5, 12, 10) {real, imag} */,
  {32'h3f9a10b0, 32'h3f5d4e92} /* (5, 12, 9) {real, imag} */,
  {32'h3f0029f4, 32'h3f9f5f8c} /* (5, 12, 8) {real, imag} */,
  {32'h4039ac44, 32'h4002e359} /* (5, 12, 7) {real, imag} */,
  {32'hc00533b6, 32'hbe8a66b0} /* (5, 12, 6) {real, imag} */,
  {32'hbd8a3259, 32'hc02f83f1} /* (5, 12, 5) {real, imag} */,
  {32'hbf496fd9, 32'hbf4e93a7} /* (5, 12, 4) {real, imag} */,
  {32'hbe415c79, 32'h3f117062} /* (5, 12, 3) {real, imag} */,
  {32'hbf6b018f, 32'h3fc44c6b} /* (5, 12, 2) {real, imag} */,
  {32'h3fbe8eca, 32'hbecda98e} /* (5, 12, 1) {real, imag} */,
  {32'h4020fad2, 32'hbf983e67} /* (5, 12, 0) {real, imag} */,
  {32'h4017d5e3, 32'h3ec488b1} /* (5, 11, 31) {real, imag} */,
  {32'h3fc94a29, 32'h4023bd4d} /* (5, 11, 30) {real, imag} */,
  {32'hbec97f4e, 32'hbfb41a08} /* (5, 11, 29) {real, imag} */,
  {32'hbfde736b, 32'h3fdf34d9} /* (5, 11, 28) {real, imag} */,
  {32'h40479bd2, 32'h3d9af95c} /* (5, 11, 27) {real, imag} */,
  {32'hbf48f719, 32'hbfe0e37d} /* (5, 11, 26) {real, imag} */,
  {32'hbfdc3560, 32'hbefdf25a} /* (5, 11, 25) {real, imag} */,
  {32'hc013f3ff, 32'hbe567170} /* (5, 11, 24) {real, imag} */,
  {32'h3f818db5, 32'hbe6f3c5b} /* (5, 11, 23) {real, imag} */,
  {32'h3f7714d4, 32'hbe7ada90} /* (5, 11, 22) {real, imag} */,
  {32'h3edbaf5f, 32'hc005f873} /* (5, 11, 21) {real, imag} */,
  {32'h3fca881c, 32'h3f802ca8} /* (5, 11, 20) {real, imag} */,
  {32'h3fe51997, 32'hbc94d058} /* (5, 11, 19) {real, imag} */,
  {32'hbf97b6d0, 32'hc01db7cf} /* (5, 11, 18) {real, imag} */,
  {32'h3f5bb3e5, 32'h3f47ec73} /* (5, 11, 17) {real, imag} */,
  {32'h3f61d80d, 32'hbead965d} /* (5, 11, 16) {real, imag} */,
  {32'hbf6d71a8, 32'hc038ae65} /* (5, 11, 15) {real, imag} */,
  {32'h3f8c76a5, 32'h3e0a75b0} /* (5, 11, 14) {real, imag} */,
  {32'h3fcfe771, 32'h3f4b7a9e} /* (5, 11, 13) {real, imag} */,
  {32'h3f3f1553, 32'hbe76daea} /* (5, 11, 12) {real, imag} */,
  {32'h3f3d226f, 32'h40916bad} /* (5, 11, 11) {real, imag} */,
  {32'hc04cba86, 32'hbf5c0d4c} /* (5, 11, 10) {real, imag} */,
  {32'hbc6a7e41, 32'hc09f9c6b} /* (5, 11, 9) {real, imag} */,
  {32'h3e2bff6f, 32'h3f507e74} /* (5, 11, 8) {real, imag} */,
  {32'hbfa1e2bc, 32'hbf1d4dae} /* (5, 11, 7) {real, imag} */,
  {32'h402ff600, 32'hc013e432} /* (5, 11, 6) {real, imag} */,
  {32'h3fa11385, 32'h3e039194} /* (5, 11, 5) {real, imag} */,
  {32'hbe9c77fb, 32'h3ff002b3} /* (5, 11, 4) {real, imag} */,
  {32'h3cd5c127, 32'hbd2d495d} /* (5, 11, 3) {real, imag} */,
  {32'hbf9329b7, 32'hbf831c0c} /* (5, 11, 2) {real, imag} */,
  {32'hbfee2c20, 32'hbfe016db} /* (5, 11, 1) {real, imag} */,
  {32'hc02204ea, 32'h401cdce3} /* (5, 11, 0) {real, imag} */,
  {32'hc051ab04, 32'h3f0131c8} /* (5, 10, 31) {real, imag} */,
  {32'hbe249ea4, 32'hbfa481a2} /* (5, 10, 30) {real, imag} */,
  {32'h3f628772, 32'hc0454d46} /* (5, 10, 29) {real, imag} */,
  {32'h40245036, 32'h400fa842} /* (5, 10, 28) {real, imag} */,
  {32'hbede51ce, 32'h3f17ddb3} /* (5, 10, 27) {real, imag} */,
  {32'hbe2f80b5, 32'hbe4e9b7d} /* (5, 10, 26) {real, imag} */,
  {32'h3fe7fced, 32'h3e95b110} /* (5, 10, 25) {real, imag} */,
  {32'hbe8bc86e, 32'hc001cae0} /* (5, 10, 24) {real, imag} */,
  {32'hbf06d8ce, 32'h40198881} /* (5, 10, 23) {real, imag} */,
  {32'hbf5257ea, 32'hbf334998} /* (5, 10, 22) {real, imag} */,
  {32'h3f2d385e, 32'h3e83c52b} /* (5, 10, 21) {real, imag} */,
  {32'hc00c7958, 32'hbe403587} /* (5, 10, 20) {real, imag} */,
  {32'h3fcf4747, 32'h40146463} /* (5, 10, 19) {real, imag} */,
  {32'h3f751cb9, 32'h3ef832ee} /* (5, 10, 18) {real, imag} */,
  {32'hbeeeeb59, 32'hbe1f1827} /* (5, 10, 17) {real, imag} */,
  {32'h3f803f66, 32'hc04a80ff} /* (5, 10, 16) {real, imag} */,
  {32'hbe84dacf, 32'h4047cca7} /* (5, 10, 15) {real, imag} */,
  {32'h3ea89044, 32'hbcd4cada} /* (5, 10, 14) {real, imag} */,
  {32'hc039bb14, 32'h3e0d027e} /* (5, 10, 13) {real, imag} */,
  {32'hbf212563, 32'h3f4ddfad} /* (5, 10, 12) {real, imag} */,
  {32'h400e2585, 32'hbfa85ae8} /* (5, 10, 11) {real, imag} */,
  {32'hbfd8e992, 32'hc03d3ec2} /* (5, 10, 10) {real, imag} */,
  {32'hc0385d8a, 32'hc020fef0} /* (5, 10, 9) {real, imag} */,
  {32'h40670953, 32'h3f8294ac} /* (5, 10, 8) {real, imag} */,
  {32'hbf444414, 32'h3e862679} /* (5, 10, 7) {real, imag} */,
  {32'hbff4988d, 32'hc01c594d} /* (5, 10, 6) {real, imag} */,
  {32'h3ecea807, 32'h40300066} /* (5, 10, 5) {real, imag} */,
  {32'h3f8643f3, 32'hbee4817b} /* (5, 10, 4) {real, imag} */,
  {32'hbfa62d74, 32'hbeb64c4c} /* (5, 10, 3) {real, imag} */,
  {32'h3fd59a25, 32'h3e115172} /* (5, 10, 2) {real, imag} */,
  {32'h40539100, 32'hbfcba251} /* (5, 10, 1) {real, imag} */,
  {32'h40a09d74, 32'h40630413} /* (5, 10, 0) {real, imag} */,
  {32'h40abc1b7, 32'h401ce76e} /* (5, 9, 31) {real, imag} */,
  {32'hc05c621c, 32'h3f61d454} /* (5, 9, 30) {real, imag} */,
  {32'hbee01ea8, 32'h3fa148ed} /* (5, 9, 29) {real, imag} */,
  {32'hbec2bb50, 32'hbff906ae} /* (5, 9, 28) {real, imag} */,
  {32'hc0336e72, 32'h400f84ad} /* (5, 9, 27) {real, imag} */,
  {32'hc06f1d8e, 32'hc006f92e} /* (5, 9, 26) {real, imag} */,
  {32'hbf09a3fe, 32'hbf0acad6} /* (5, 9, 25) {real, imag} */,
  {32'hbf1a746c, 32'h3e930b38} /* (5, 9, 24) {real, imag} */,
  {32'hbfa04efc, 32'h3e985573} /* (5, 9, 23) {real, imag} */,
  {32'h4058406a, 32'h400b3912} /* (5, 9, 22) {real, imag} */,
  {32'h4050c463, 32'h400f0951} /* (5, 9, 21) {real, imag} */,
  {32'hc01a8be7, 32'h3fabb8e5} /* (5, 9, 20) {real, imag} */,
  {32'h3f111837, 32'h3fe97a9c} /* (5, 9, 19) {real, imag} */,
  {32'hbf2f1d76, 32'hc00f1755} /* (5, 9, 18) {real, imag} */,
  {32'hc013e270, 32'h3fa35734} /* (5, 9, 17) {real, imag} */,
  {32'h3fe898a1, 32'h3f94b62a} /* (5, 9, 16) {real, imag} */,
  {32'hc01f9b3c, 32'hc03942f4} /* (5, 9, 15) {real, imag} */,
  {32'h3fe0f21e, 32'hbf6e37f5} /* (5, 9, 14) {real, imag} */,
  {32'hbf6ea113, 32'hbf92a2ad} /* (5, 9, 13) {real, imag} */,
  {32'h3fa6bc4e, 32'h3eb6ea12} /* (5, 9, 12) {real, imag} */,
  {32'h3f6f426e, 32'hbf291b72} /* (5, 9, 11) {real, imag} */,
  {32'hbfbb6337, 32'hbef38df4} /* (5, 9, 10) {real, imag} */,
  {32'h3da16d77, 32'hbe81f1fa} /* (5, 9, 9) {real, imag} */,
  {32'hbf37efeb, 32'hbef6272c} /* (5, 9, 8) {real, imag} */,
  {32'h40490474, 32'h3fff9c75} /* (5, 9, 7) {real, imag} */,
  {32'hbf5c842a, 32'h40449b4d} /* (5, 9, 6) {real, imag} */,
  {32'h3fc24979, 32'h3e46bd8c} /* (5, 9, 5) {real, imag} */,
  {32'h404026a1, 32'hbf340ccf} /* (5, 9, 4) {real, imag} */,
  {32'h3fc606b8, 32'hc045b338} /* (5, 9, 3) {real, imag} */,
  {32'h3f83ff41, 32'hc0462b80} /* (5, 9, 2) {real, imag} */,
  {32'hbfc6cb47, 32'h403c9fe1} /* (5, 9, 1) {real, imag} */,
  {32'hc03370e3, 32'h3eed0818} /* (5, 9, 0) {real, imag} */,
  {32'hbfee2973, 32'h40a0dfab} /* (5, 8, 31) {real, imag} */,
  {32'h3fce8ef6, 32'h3eb33a66} /* (5, 8, 30) {real, imag} */,
  {32'h3f89a3af, 32'hbfdec7b5} /* (5, 8, 29) {real, imag} */,
  {32'hbfcb0572, 32'h3fa8ad70} /* (5, 8, 28) {real, imag} */,
  {32'h3fbc4363, 32'h3f68de19} /* (5, 8, 27) {real, imag} */,
  {32'hbf91f928, 32'hc02b1978} /* (5, 8, 26) {real, imag} */,
  {32'h408a7d9d, 32'hbf1e5827} /* (5, 8, 25) {real, imag} */,
  {32'h408c3f64, 32'hc05a3a91} /* (5, 8, 24) {real, imag} */,
  {32'hbe6f3d14, 32'hc00061da} /* (5, 8, 23) {real, imag} */,
  {32'hc057e571, 32'h4021db4f} /* (5, 8, 22) {real, imag} */,
  {32'h3f77e49b, 32'hc04d86b0} /* (5, 8, 21) {real, imag} */,
  {32'h3fd292fb, 32'h3fdd6393} /* (5, 8, 20) {real, imag} */,
  {32'hbf67f26d, 32'h3fc0c93e} /* (5, 8, 19) {real, imag} */,
  {32'hbfb0ee06, 32'h3f93f940} /* (5, 8, 18) {real, imag} */,
  {32'hbf4c0a7e, 32'h3fe0441e} /* (5, 8, 17) {real, imag} */,
  {32'h3f870503, 32'h3fc88c85} /* (5, 8, 16) {real, imag} */,
  {32'h3dc903a1, 32'hbde9a344} /* (5, 8, 15) {real, imag} */,
  {32'h4021a876, 32'hbe34b07b} /* (5, 8, 14) {real, imag} */,
  {32'hbebee095, 32'hbf826334} /* (5, 8, 13) {real, imag} */,
  {32'hbfb9a342, 32'h3e8673a1} /* (5, 8, 12) {real, imag} */,
  {32'h3f885d6d, 32'hc01fa70e} /* (5, 8, 11) {real, imag} */,
  {32'hbfc56cbb, 32'h3fa446b6} /* (5, 8, 10) {real, imag} */,
  {32'h3fe93622, 32'h3f63d655} /* (5, 8, 9) {real, imag} */,
  {32'h3e0fcca6, 32'h3f9b61e9} /* (5, 8, 8) {real, imag} */,
  {32'h3fa54d06, 32'hbf811eb5} /* (5, 8, 7) {real, imag} */,
  {32'hc0277f0f, 32'h3fcbc753} /* (5, 8, 6) {real, imag} */,
  {32'hbfa80aad, 32'h3ea94e13} /* (5, 8, 5) {real, imag} */,
  {32'hc05c5d2c, 32'h3fa2d2e7} /* (5, 8, 4) {real, imag} */,
  {32'h3d54cad2, 32'hbfc152b0} /* (5, 8, 3) {real, imag} */,
  {32'hc017bb41, 32'hbf7d76b0} /* (5, 8, 2) {real, imag} */,
  {32'hc01cef36, 32'h3eba0d0e} /* (5, 8, 1) {real, imag} */,
  {32'hc0516c3f, 32'h3eb3b691} /* (5, 8, 0) {real, imag} */,
  {32'hbd4bd0c0, 32'hc05ec0af} /* (5, 7, 31) {real, imag} */,
  {32'hbf8fc1ff, 32'hbf8627ea} /* (5, 7, 30) {real, imag} */,
  {32'hbfdbcada, 32'hc04daef7} /* (5, 7, 29) {real, imag} */,
  {32'hbf42f68e, 32'h3f87126e} /* (5, 7, 28) {real, imag} */,
  {32'h407b4371, 32'h3e0cc8a0} /* (5, 7, 27) {real, imag} */,
  {32'h3fbbc27a, 32'h3de26aa3} /* (5, 7, 26) {real, imag} */,
  {32'h40b898cf, 32'h4035fbcf} /* (5, 7, 25) {real, imag} */,
  {32'h4090bf8b, 32'hc08804c1} /* (5, 7, 24) {real, imag} */,
  {32'hbf698581, 32'h40828555} /* (5, 7, 23) {real, imag} */,
  {32'hbf9ade38, 32'h3ff5d54a} /* (5, 7, 22) {real, imag} */,
  {32'hc001cdb3, 32'hc021d753} /* (5, 7, 21) {real, imag} */,
  {32'h3f2ed021, 32'h401ae579} /* (5, 7, 20) {real, imag} */,
  {32'hc022efd2, 32'hbfad5e61} /* (5, 7, 19) {real, imag} */,
  {32'hbfe687e5, 32'h3fac1dbd} /* (5, 7, 18) {real, imag} */,
  {32'h3f96d2d2, 32'h3fe88aac} /* (5, 7, 17) {real, imag} */,
  {32'hbfdf2bee, 32'hbf128fbc} /* (5, 7, 16) {real, imag} */,
  {32'h3d62b7de, 32'hbf8718ba} /* (5, 7, 15) {real, imag} */,
  {32'hbdf25361, 32'hbf608bb5} /* (5, 7, 14) {real, imag} */,
  {32'h4024690b, 32'h3f77fc15} /* (5, 7, 13) {real, imag} */,
  {32'h3f08916d, 32'hbdb71cc2} /* (5, 7, 12) {real, imag} */,
  {32'h3f0aca99, 32'h407f2085} /* (5, 7, 11) {real, imag} */,
  {32'h3f632e9e, 32'hbf26b4b5} /* (5, 7, 10) {real, imag} */,
  {32'h4046c4df, 32'hbf9cb95d} /* (5, 7, 9) {real, imag} */,
  {32'hc03e6fef, 32'h401102e8} /* (5, 7, 8) {real, imag} */,
  {32'hc0878dfb, 32'hbeb40064} /* (5, 7, 7) {real, imag} */,
  {32'h402c0ae2, 32'h40a96982} /* (5, 7, 6) {real, imag} */,
  {32'hbfc528cc, 32'hc00afc01} /* (5, 7, 5) {real, imag} */,
  {32'hbef6e11f, 32'h4093ade1} /* (5, 7, 4) {real, imag} */,
  {32'h402bee61, 32'hbf7c0ab8} /* (5, 7, 3) {real, imag} */,
  {32'hc04a77ee, 32'h3fcbc35b} /* (5, 7, 2) {real, imag} */,
  {32'h40e38bbf, 32'hc05d41b7} /* (5, 7, 1) {real, imag} */,
  {32'hc01f65cc, 32'h3ed500df} /* (5, 7, 0) {real, imag} */,
  {32'h3f1ae0b8, 32'h40b3aa13} /* (5, 6, 31) {real, imag} */,
  {32'h3fb37722, 32'hc04f20e0} /* (5, 6, 30) {real, imag} */,
  {32'h3e6f5746, 32'hbf51ff86} /* (5, 6, 29) {real, imag} */,
  {32'hbfc8e110, 32'h40649cfb} /* (5, 6, 28) {real, imag} */,
  {32'h3f418cc0, 32'hbeecbbf2} /* (5, 6, 27) {real, imag} */,
  {32'hbf764cb1, 32'hbf05d391} /* (5, 6, 26) {real, imag} */,
  {32'hc01f10c4, 32'hbd6f3431} /* (5, 6, 25) {real, imag} */,
  {32'h3f8921ea, 32'hbf4f8e42} /* (5, 6, 24) {real, imag} */,
  {32'h3fd8386f, 32'hbf2a26f6} /* (5, 6, 23) {real, imag} */,
  {32'h3f116813, 32'hbf8d8c2b} /* (5, 6, 22) {real, imag} */,
  {32'h3fc543ac, 32'hbf1fd771} /* (5, 6, 21) {real, imag} */,
  {32'h3fabd762, 32'h3fd1a2d4} /* (5, 6, 20) {real, imag} */,
  {32'hbf84bad3, 32'hbed76af8} /* (5, 6, 19) {real, imag} */,
  {32'hc0446eb9, 32'hbdfe8523} /* (5, 6, 18) {real, imag} */,
  {32'hbf6e1eb2, 32'hc03a6208} /* (5, 6, 17) {real, imag} */,
  {32'h3ea5105e, 32'h40410c77} /* (5, 6, 16) {real, imag} */,
  {32'hbf98fccc, 32'hbe426bc2} /* (5, 6, 15) {real, imag} */,
  {32'h3f1b3d98, 32'hbec87fb9} /* (5, 6, 14) {real, imag} */,
  {32'hbf925132, 32'hc00a0770} /* (5, 6, 13) {real, imag} */,
  {32'h3f1d57c3, 32'h3f63911a} /* (5, 6, 12) {real, imag} */,
  {32'hbda0fdb6, 32'hc0612fbc} /* (5, 6, 11) {real, imag} */,
  {32'h40909daa, 32'hbfe10b9c} /* (5, 6, 10) {real, imag} */,
  {32'h3f6d8a42, 32'h3e880aa6} /* (5, 6, 9) {real, imag} */,
  {32'h403fe0e8, 32'h401c6eb1} /* (5, 6, 8) {real, imag} */,
  {32'hbfe249bf, 32'hbe6ffc0f} /* (5, 6, 7) {real, imag} */,
  {32'h40510580, 32'hc03a86c0} /* (5, 6, 6) {real, imag} */,
  {32'hc03b5608, 32'h3e4eec0a} /* (5, 6, 5) {real, imag} */,
  {32'hbfc5c414, 32'h3f9e479f} /* (5, 6, 4) {real, imag} */,
  {32'hbeb7cc61, 32'hc0412712} /* (5, 6, 3) {real, imag} */,
  {32'h403a9f94, 32'h3fc82ef9} /* (5, 6, 2) {real, imag} */,
  {32'hc0b84561, 32'hbed7c82b} /* (5, 6, 1) {real, imag} */,
  {32'h3f20dc05, 32'hbfc0e2b4} /* (5, 6, 0) {real, imag} */,
  {32'hc0272efd, 32'h401246b0} /* (5, 5, 31) {real, imag} */,
  {32'h40281f28, 32'hbe885dee} /* (5, 5, 30) {real, imag} */,
  {32'h4050b7a0, 32'h40217033} /* (5, 5, 29) {real, imag} */,
  {32'hc04d8572, 32'h3f024562} /* (5, 5, 28) {real, imag} */,
  {32'hbf0739ee, 32'hbfb27c4c} /* (5, 5, 27) {real, imag} */,
  {32'h3ee1a944, 32'h40262d57} /* (5, 5, 26) {real, imag} */,
  {32'h402c385e, 32'hbe910810} /* (5, 5, 25) {real, imag} */,
  {32'h4078f31b, 32'hc0595302} /* (5, 5, 24) {real, imag} */,
  {32'h3fcadd4b, 32'h401fa993} /* (5, 5, 23) {real, imag} */,
  {32'h400e096f, 32'h3fc3376d} /* (5, 5, 22) {real, imag} */,
  {32'hbecef7eb, 32'hbffa7f68} /* (5, 5, 21) {real, imag} */,
  {32'h3ec27b29, 32'hbf28fde9} /* (5, 5, 20) {real, imag} */,
  {32'h3c8257ef, 32'h3fa27efc} /* (5, 5, 19) {real, imag} */,
  {32'hbfa71920, 32'hbce9454c} /* (5, 5, 18) {real, imag} */,
  {32'hbecab523, 32'h3f043559} /* (5, 5, 17) {real, imag} */,
  {32'hbefc070f, 32'hbebdf3eb} /* (5, 5, 16) {real, imag} */,
  {32'h3f4b842b, 32'hbf16d0f2} /* (5, 5, 15) {real, imag} */,
  {32'hbfc1a4a4, 32'h40200d61} /* (5, 5, 14) {real, imag} */,
  {32'hbfafe74d, 32'h3ff7d59f} /* (5, 5, 13) {real, imag} */,
  {32'hbfc683a0, 32'hbec2022a} /* (5, 5, 12) {real, imag} */,
  {32'h40033778, 32'h3f1d0c8a} /* (5, 5, 11) {real, imag} */,
  {32'hbe4f32f7, 32'h3e832ddd} /* (5, 5, 10) {real, imag} */,
  {32'hbfa9e7a7, 32'hbea1c918} /* (5, 5, 9) {real, imag} */,
  {32'hbee496a6, 32'h3de6a6af} /* (5, 5, 8) {real, imag} */,
  {32'h40652a28, 32'h3fffcab4} /* (5, 5, 7) {real, imag} */,
  {32'h40664fe6, 32'hbe561a66} /* (5, 5, 6) {real, imag} */,
  {32'h3fea0327, 32'hc01b0258} /* (5, 5, 5) {real, imag} */,
  {32'hbd5fa857, 32'hc0974581} /* (5, 5, 4) {real, imag} */,
  {32'hbf503096, 32'h3f88b712} /* (5, 5, 3) {real, imag} */,
  {32'hc0909846, 32'h3ef19a38} /* (5, 5, 2) {real, imag} */,
  {32'hc0f4dcc6, 32'h40c1b4ae} /* (5, 5, 1) {real, imag} */,
  {32'hc1122386, 32'h407b6cf7} /* (5, 5, 0) {real, imag} */,
  {32'h402fd995, 32'hbee1e5cb} /* (5, 4, 31) {real, imag} */,
  {32'hc12ccdc3, 32'hc10117d8} /* (5, 4, 30) {real, imag} */,
  {32'hbf6512a6, 32'hbf549fd3} /* (5, 4, 29) {real, imag} */,
  {32'h40a1dd7a, 32'hc0956ca2} /* (5, 4, 28) {real, imag} */,
  {32'h40823a65, 32'hbfdce113} /* (5, 4, 27) {real, imag} */,
  {32'h3f21a316, 32'hc0d3b4f0} /* (5, 4, 26) {real, imag} */,
  {32'h401f2b4d, 32'h40a3e6ef} /* (5, 4, 25) {real, imag} */,
  {32'hbfef9a82, 32'h40024658} /* (5, 4, 24) {real, imag} */,
  {32'hbfbf75bb, 32'h3f94de1d} /* (5, 4, 23) {real, imag} */,
  {32'h3e837953, 32'hbf9e4f82} /* (5, 4, 22) {real, imag} */,
  {32'hbf1d5bd1, 32'h40025c36} /* (5, 4, 21) {real, imag} */,
  {32'hbed2ea8a, 32'h3f85115f} /* (5, 4, 20) {real, imag} */,
  {32'h3ddbf666, 32'h3ffdff5c} /* (5, 4, 19) {real, imag} */,
  {32'hbebd6b4f, 32'h3ecdab2f} /* (5, 4, 18) {real, imag} */,
  {32'hbecceedd, 32'h3fdc2dbd} /* (5, 4, 17) {real, imag} */,
  {32'h3e2445be, 32'hbf409260} /* (5, 4, 16) {real, imag} */,
  {32'hbec9cb55, 32'hbf669be9} /* (5, 4, 15) {real, imag} */,
  {32'hc02c2cdc, 32'h3fa0875f} /* (5, 4, 14) {real, imag} */,
  {32'h4035cc54, 32'hbf323201} /* (5, 4, 13) {real, imag} */,
  {32'h3f077251, 32'h3fbbb9bd} /* (5, 4, 12) {real, imag} */,
  {32'h3fc6a016, 32'h3fbf70c6} /* (5, 4, 11) {real, imag} */,
  {32'hbf184884, 32'hbf7bdc25} /* (5, 4, 10) {real, imag} */,
  {32'hbfed25d4, 32'hc0276d15} /* (5, 4, 9) {real, imag} */,
  {32'hbfb6185f, 32'h3e06a849} /* (5, 4, 8) {real, imag} */,
  {32'h3f58d8c9, 32'hbf79e9b4} /* (5, 4, 7) {real, imag} */,
  {32'hc09d94e5, 32'h3eb312c1} /* (5, 4, 6) {real, imag} */,
  {32'hbf728cb8, 32'h3f53e868} /* (5, 4, 5) {real, imag} */,
  {32'hc005bdb6, 32'h3fca8684} /* (5, 4, 4) {real, imag} */,
  {32'h3c847f3f, 32'h3fdda250} /* (5, 4, 3) {real, imag} */,
  {32'hc1104b52, 32'h4011871f} /* (5, 4, 2) {real, imag} */,
  {32'h40d167ae, 32'hc011a9c7} /* (5, 4, 1) {real, imag} */,
  {32'h41312030, 32'hc035a22a} /* (5, 4, 0) {real, imag} */,
  {32'hc113464c, 32'h3f850d83} /* (5, 3, 31) {real, imag} */,
  {32'hc064c0c9, 32'hc060ef6b} /* (5, 3, 30) {real, imag} */,
  {32'h3f72a659, 32'h4097a7c7} /* (5, 3, 29) {real, imag} */,
  {32'h3fde757e, 32'hbf3c18d0} /* (5, 3, 28) {real, imag} */,
  {32'hbf131618, 32'h408f01f5} /* (5, 3, 27) {real, imag} */,
  {32'hc02cc475, 32'hc034d93e} /* (5, 3, 26) {real, imag} */,
  {32'h3cb6057a, 32'h406b8ee1} /* (5, 3, 25) {real, imag} */,
  {32'hbfce2121, 32'h400a8a83} /* (5, 3, 24) {real, imag} */,
  {32'h40163d8f, 32'h4019e6b1} /* (5, 3, 23) {real, imag} */,
  {32'h3fa56779, 32'hbff95acc} /* (5, 3, 22) {real, imag} */,
  {32'h3f95a72e, 32'hbe940fa9} /* (5, 3, 21) {real, imag} */,
  {32'hbe3718b0, 32'hbff9d36a} /* (5, 3, 20) {real, imag} */,
  {32'h3fadbfd4, 32'hbfbe038d} /* (5, 3, 19) {real, imag} */,
  {32'hc01c5a30, 32'h3b737b2c} /* (5, 3, 18) {real, imag} */,
  {32'hbe0006cd, 32'h3fbaec90} /* (5, 3, 17) {real, imag} */,
  {32'hbf905fad, 32'h3fd3d5e1} /* (5, 3, 16) {real, imag} */,
  {32'hbfcad96b, 32'h3f37486f} /* (5, 3, 15) {real, imag} */,
  {32'h402ec3d2, 32'h3e33bd40} /* (5, 3, 14) {real, imag} */,
  {32'h3f8b2bcd, 32'h3f012f23} /* (5, 3, 13) {real, imag} */,
  {32'h3fd09b47, 32'hc0737cc2} /* (5, 3, 12) {real, imag} */,
  {32'h3f6862d5, 32'hbf81f1d3} /* (5, 3, 11) {real, imag} */,
  {32'h4004257d, 32'hbf16f761} /* (5, 3, 10) {real, imag} */,
  {32'h3e8afb8d, 32'hbe9b9b31} /* (5, 3, 9) {real, imag} */,
  {32'h401c83ce, 32'hbf5cbf02} /* (5, 3, 8) {real, imag} */,
  {32'hbf0c92a6, 32'h3dcea0f7} /* (5, 3, 7) {real, imag} */,
  {32'h3e3670a5, 32'h406f508c} /* (5, 3, 6) {real, imag} */,
  {32'h40c70d87, 32'hc01f3264} /* (5, 3, 5) {real, imag} */,
  {32'h3e04b724, 32'h40a2c8c7} /* (5, 3, 4) {real, imag} */,
  {32'h40b09664, 32'hbece51df} /* (5, 3, 3) {real, imag} */,
  {32'hc0c3df69, 32'h4065fbcb} /* (5, 3, 2) {real, imag} */,
  {32'h41a1700a, 32'hbf8d8ff1} /* (5, 3, 1) {real, imag} */,
  {32'hc0be0f01, 32'h404e89a2} /* (5, 3, 0) {real, imag} */,
  {32'hc136e0ad, 32'h41fb6439} /* (5, 2, 31) {real, imag} */,
  {32'h4097097e, 32'hc1cf2c64} /* (5, 2, 30) {real, imag} */,
  {32'hc038effb, 32'h40a97526} /* (5, 2, 29) {real, imag} */,
  {32'h40f84785, 32'h40c819f0} /* (5, 2, 28) {real, imag} */,
  {32'h4073739d, 32'hc105d7a4} /* (5, 2, 27) {real, imag} */,
  {32'h3f33072a, 32'hc06a7b7a} /* (5, 2, 26) {real, imag} */,
  {32'hc0079ac3, 32'h40025595} /* (5, 2, 25) {real, imag} */,
  {32'h3e39bfc9, 32'h40821c3b} /* (5, 2, 24) {real, imag} */,
  {32'h3f908d58, 32'hc017a708} /* (5, 2, 23) {real, imag} */,
  {32'hbfd269ff, 32'hbfe6cbec} /* (5, 2, 22) {real, imag} */,
  {32'h3f9764fa, 32'h3e0c1de5} /* (5, 2, 21) {real, imag} */,
  {32'hbf99e90d, 32'hc046f0dc} /* (5, 2, 20) {real, imag} */,
  {32'h3e3bade1, 32'h3fa6613f} /* (5, 2, 19) {real, imag} */,
  {32'hbfb3f172, 32'hbe99989e} /* (5, 2, 18) {real, imag} */,
  {32'h40470f29, 32'hbf30cd4a} /* (5, 2, 17) {real, imag} */,
  {32'hbfa54b41, 32'h3fd7d883} /* (5, 2, 16) {real, imag} */,
  {32'h3e0cbd60, 32'h3c72ed7d} /* (5, 2, 15) {real, imag} */,
  {32'h3f213394, 32'hbee044e4} /* (5, 2, 14) {real, imag} */,
  {32'hbe2310a7, 32'hbd322e36} /* (5, 2, 13) {real, imag} */,
  {32'hbf22afa0, 32'h3eded270} /* (5, 2, 12) {real, imag} */,
  {32'h3fbb3e14, 32'hbfca6bc1} /* (5, 2, 11) {real, imag} */,
  {32'h3eaabd67, 32'hbfd53c84} /* (5, 2, 10) {real, imag} */,
  {32'hc007738b, 32'hbfab94ef} /* (5, 2, 9) {real, imag} */,
  {32'h401c05ae, 32'hc02c3680} /* (5, 2, 8) {real, imag} */,
  {32'h3e06d04c, 32'h4081bd4c} /* (5, 2, 7) {real, imag} */,
  {32'hc017585c, 32'h403f7f11} /* (5, 2, 6) {real, imag} */,
  {32'h4100a4de, 32'hbf6c5326} /* (5, 2, 5) {real, imag} */,
  {32'hc10634bc, 32'h3fed488a} /* (5, 2, 4) {real, imag} */,
  {32'hbfedf73f, 32'h4105c269} /* (5, 2, 3) {real, imag} */,
  {32'h404f8a8b, 32'hc1a00a3f} /* (5, 2, 2) {real, imag} */,
  {32'hc093818b, 32'h413a6913} /* (5, 2, 1) {real, imag} */,
  {32'hc008cb01, 32'h3fd00d3f} /* (5, 2, 0) {real, imag} */,
  {32'h41122117, 32'hc1b0298d} /* (5, 1, 31) {real, imag} */,
  {32'hc057f2af, 32'h402372a3} /* (5, 1, 30) {real, imag} */,
  {32'h3ffed1bc, 32'h407cfbf3} /* (5, 1, 29) {real, imag} */,
  {32'h40c3c742, 32'h3f60b2ec} /* (5, 1, 28) {real, imag} */,
  {32'hc0c948a1, 32'h409b7a59} /* (5, 1, 27) {real, imag} */,
  {32'hbfcb4d0b, 32'hbf4bff48} /* (5, 1, 26) {real, imag} */,
  {32'hbfd91ea6, 32'hbef8bb81} /* (5, 1, 25) {real, imag} */,
  {32'hbfd81ed3, 32'h4036b250} /* (5, 1, 24) {real, imag} */,
  {32'h3f5f104f, 32'hbfc50179} /* (5, 1, 23) {real, imag} */,
  {32'h4005cc47, 32'h3fb53b23} /* (5, 1, 22) {real, imag} */,
  {32'h3fb7df63, 32'h3ff775b8} /* (5, 1, 21) {real, imag} */,
  {32'hbfc5472d, 32'hbf14f934} /* (5, 1, 20) {real, imag} */,
  {32'hbeec0151, 32'hbe577fa0} /* (5, 1, 19) {real, imag} */,
  {32'h409e1ee8, 32'hbf9b1a93} /* (5, 1, 18) {real, imag} */,
  {32'hc004e58c, 32'h3f2f0935} /* (5, 1, 17) {real, imag} */,
  {32'hbf801fb0, 32'hbdc45d4a} /* (5, 1, 16) {real, imag} */,
  {32'hbdb1ecd5, 32'hbf2fe896} /* (5, 1, 15) {real, imag} */,
  {32'hbf3373a9, 32'hbf8a30ac} /* (5, 1, 14) {real, imag} */,
  {32'hbeb92a98, 32'h3cc8b997} /* (5, 1, 13) {real, imag} */,
  {32'h3e0aee17, 32'h4027db4c} /* (5, 1, 12) {real, imag} */,
  {32'hc04d1370, 32'hbf5dfee8} /* (5, 1, 11) {real, imag} */,
  {32'h400626f2, 32'h3efdd859} /* (5, 1, 10) {real, imag} */,
  {32'hc04e1db6, 32'hbf6ad560} /* (5, 1, 9) {real, imag} */,
  {32'hc014941d, 32'hbfd30dd7} /* (5, 1, 8) {real, imag} */,
  {32'h3f4948e3, 32'h403d81ec} /* (5, 1, 7) {real, imag} */,
  {32'h40025ce8, 32'hbf495afd} /* (5, 1, 6) {real, imag} */,
  {32'hc0607d42, 32'h3c802d18} /* (5, 1, 5) {real, imag} */,
  {32'h4018f32d, 32'hc08c1844} /* (5, 1, 4) {real, imag} */,
  {32'hbfb3d9f7, 32'hc04ff685} /* (5, 1, 3) {real, imag} */,
  {32'hc1c3a727, 32'h41362d5a} /* (5, 1, 2) {real, imag} */,
  {32'h41f0874a, 32'hc13b802b} /* (5, 1, 1) {real, imag} */,
  {32'h41459674, 32'hc19a32ba} /* (5, 1, 0) {real, imag} */,
  {32'h3ebdfd1d, 32'hc1dc1fd6} /* (5, 0, 31) {real, imag} */,
  {32'h408e1be2, 32'h40ebf752} /* (5, 0, 30) {real, imag} */,
  {32'hc09d2a03, 32'hbfe69f80} /* (5, 0, 29) {real, imag} */,
  {32'h3f7e5061, 32'h40b994c0} /* (5, 0, 28) {real, imag} */,
  {32'h3ee28906, 32'h41039572} /* (5, 0, 27) {real, imag} */,
  {32'hc001eb1b, 32'hbf98fbe5} /* (5, 0, 26) {real, imag} */,
  {32'hbfc4af65, 32'hc0100ce9} /* (5, 0, 25) {real, imag} */,
  {32'h3f697f93, 32'hc0b1186f} /* (5, 0, 24) {real, imag} */,
  {32'hc0862a32, 32'hbeb7f0c6} /* (5, 0, 23) {real, imag} */,
  {32'hc046c0e9, 32'hbf664861} /* (5, 0, 22) {real, imag} */,
  {32'hbe4f03d4, 32'h40286376} /* (5, 0, 21) {real, imag} */,
  {32'hbe8342f9, 32'hc078eb62} /* (5, 0, 20) {real, imag} */,
  {32'h3ea1555c, 32'h3fb35a7a} /* (5, 0, 19) {real, imag} */,
  {32'h402e143d, 32'h3ec36a3e} /* (5, 0, 18) {real, imag} */,
  {32'hbddbc3a8, 32'h3fa05ea2} /* (5, 0, 17) {real, imag} */,
  {32'h40203f1d, 32'hbf2dbd3d} /* (5, 0, 16) {real, imag} */,
  {32'hbe1f8122, 32'h3ecd5c71} /* (5, 0, 15) {real, imag} */,
  {32'hbf4d7535, 32'h3fcdcc67} /* (5, 0, 14) {real, imag} */,
  {32'h4018a80e, 32'hc00d4a76} /* (5, 0, 13) {real, imag} */,
  {32'h3fb3ff8e, 32'hc033920e} /* (5, 0, 12) {real, imag} */,
  {32'hbf7722d3, 32'hbf264e94} /* (5, 0, 11) {real, imag} */,
  {32'hc063744f, 32'h3e8423e7} /* (5, 0, 10) {real, imag} */,
  {32'hbffd0919, 32'hbfac93ef} /* (5, 0, 9) {real, imag} */,
  {32'hc06d38ef, 32'h400658f4} /* (5, 0, 8) {real, imag} */,
  {32'hbfddc9c2, 32'h3fd3b395} /* (5, 0, 7) {real, imag} */,
  {32'h400b9005, 32'h3f77f103} /* (5, 0, 6) {real, imag} */,
  {32'h3fd4f815, 32'h3f82b3d8} /* (5, 0, 5) {real, imag} */,
  {32'h3f5f5806, 32'h3ec6de7a} /* (5, 0, 4) {real, imag} */,
  {32'h4014e698, 32'h40c71ffa} /* (5, 0, 3) {real, imag} */,
  {32'hc155d1fa, 32'h408f3c4a} /* (5, 0, 2) {real, imag} */,
  {32'h41bf434e, 32'hc06a13f0} /* (5, 0, 1) {real, imag} */,
  {32'h402bf908, 32'hc1a493ea} /* (5, 0, 0) {real, imag} */,
  {32'h40e7006a, 32'h42e4c5b8} /* (4, 31, 31) {real, imag} */,
  {32'hc1c317df, 32'hc25ee6e3} /* (4, 31, 30) {real, imag} */,
  {32'h4071ea86, 32'hc0fa3c9f} /* (4, 31, 29) {real, imag} */,
  {32'h40be14b6, 32'h4101d080} /* (4, 31, 28) {real, imag} */,
  {32'h3ecf40a8, 32'hc1172f38} /* (4, 31, 27) {real, imag} */,
  {32'h3fb848df, 32'hc09bbce7} /* (4, 31, 26) {real, imag} */,
  {32'h40927df3, 32'h403ce5d6} /* (4, 31, 25) {real, imag} */,
  {32'hc0b37989, 32'hc088a5be} /* (4, 31, 24) {real, imag} */,
  {32'h400ef6bf, 32'h40868bec} /* (4, 31, 23) {real, imag} */,
  {32'hbf42b01e, 32'h3eaacc9d} /* (4, 31, 22) {real, imag} */,
  {32'hc03dc3b7, 32'hbf7687af} /* (4, 31, 21) {real, imag} */,
  {32'hbdd0917f, 32'h404048e9} /* (4, 31, 20) {real, imag} */,
  {32'h3e972fce, 32'h3e4cc2f4} /* (4, 31, 19) {real, imag} */,
  {32'hc0484c0c, 32'h3f4a479a} /* (4, 31, 18) {real, imag} */,
  {32'hbeff0de6, 32'hbf3f81bf} /* (4, 31, 17) {real, imag} */,
  {32'hbfceb193, 32'hbeee13dd} /* (4, 31, 16) {real, imag} */,
  {32'hbfba89d8, 32'h3d7e8d30} /* (4, 31, 15) {real, imag} */,
  {32'h3c4986f2, 32'hc081babf} /* (4, 31, 14) {real, imag} */,
  {32'h3f94715b, 32'hbfe70035} /* (4, 31, 13) {real, imag} */,
  {32'hbf2544dc, 32'h3fe95c1e} /* (4, 31, 12) {real, imag} */,
  {32'h40d54d63, 32'h3f7b1802} /* (4, 31, 11) {real, imag} */,
  {32'hc0823008, 32'h408b7f47} /* (4, 31, 10) {real, imag} */,
  {32'h3fa937a6, 32'hbfef9820} /* (4, 31, 9) {real, imag} */,
  {32'h40814e4e, 32'hc02646a6} /* (4, 31, 8) {real, imag} */,
  {32'hbfeb043e, 32'hbfe931bb} /* (4, 31, 7) {real, imag} */,
  {32'hbe31e5bb, 32'hc0781325} /* (4, 31, 6) {real, imag} */,
  {32'h414e30bd, 32'hc1608355} /* (4, 31, 5) {real, imag} */,
  {32'hc078edbc, 32'h40b0b6e9} /* (4, 31, 4) {real, imag} */,
  {32'h40782d77, 32'h401fddc9} /* (4, 31, 3) {real, imag} */,
  {32'h3f86e60b, 32'hc1ead033} /* (4, 31, 2) {real, imag} */,
  {32'hc1f846e9, 32'h4297ad61} /* (4, 31, 1) {real, imag} */,
  {32'hc1c80f1d, 32'h426f6af6} /* (4, 31, 0) {real, imag} */,
  {32'h41540e86, 32'hc229ffb7} /* (4, 30, 31) {real, imag} */,
  {32'hc128dc08, 32'h41ad4b29} /* (4, 30, 30) {real, imag} */,
  {32'hbfec2131, 32'h40476acc} /* (4, 30, 29) {real, imag} */,
  {32'h41397d6a, 32'hc16014e9} /* (4, 30, 28) {real, imag} */,
  {32'hbe9a6503, 32'h415e1578} /* (4, 30, 27) {real, imag} */,
  {32'h40a4b623, 32'hbfb86729} /* (4, 30, 26) {real, imag} */,
  {32'hc04c536e, 32'hc0412846} /* (4, 30, 25) {real, imag} */,
  {32'hbe46dd04, 32'h40694703} /* (4, 30, 24) {real, imag} */,
  {32'h3ff7d26a, 32'h3f821546} /* (4, 30, 23) {real, imag} */,
  {32'h3f54dd40, 32'h3fb26a98} /* (4, 30, 22) {real, imag} */,
  {32'h400fb283, 32'h409889f8} /* (4, 30, 21) {real, imag} */,
  {32'hbfab0afe, 32'h3d164d32} /* (4, 30, 20) {real, imag} */,
  {32'h3f78674e, 32'hbefef6ef} /* (4, 30, 19) {real, imag} */,
  {32'h3e077e67, 32'h4013ca58} /* (4, 30, 18) {real, imag} */,
  {32'h3fc5a361, 32'hbfa0233c} /* (4, 30, 17) {real, imag} */,
  {32'hbfffdf68, 32'hbfe9bf47} /* (4, 30, 16) {real, imag} */,
  {32'h3ea5eba1, 32'h3ec08774} /* (4, 30, 15) {real, imag} */,
  {32'hc0392a72, 32'hbfe9e4d1} /* (4, 30, 14) {real, imag} */,
  {32'h3fe25252, 32'h3ccc0ea2} /* (4, 30, 13) {real, imag} */,
  {32'h3f9c8fb1, 32'h3fa5037d} /* (4, 30, 12) {real, imag} */,
  {32'hc04ab0f1, 32'h40006b50} /* (4, 30, 11) {real, imag} */,
  {32'h405b96e1, 32'h400b9834} /* (4, 30, 10) {real, imag} */,
  {32'h4011f205, 32'hc069d4b3} /* (4, 30, 9) {real, imag} */,
  {32'hc087c7f0, 32'h4093bbe7} /* (4, 30, 8) {real, imag} */,
  {32'hbf54daa7, 32'hc040ca0e} /* (4, 30, 7) {real, imag} */,
  {32'h3e0b00fd, 32'h3e84a4e7} /* (4, 30, 6) {real, imag} */,
  {32'hbfc36d5f, 32'hc00c0275} /* (4, 30, 5) {real, imag} */,
  {32'h414b7da9, 32'hc1037185} /* (4, 30, 4) {real, imag} */,
  {32'h406d31cc, 32'hc0b9549b} /* (4, 30, 3) {real, imag} */,
  {32'hc1be7cca, 32'h4237fb5b} /* (4, 30, 2) {real, imag} */,
  {32'h41847eef, 32'hc299b604} /* (4, 30, 1) {real, imag} */,
  {32'h40bddd35, 32'hc22f47c3} /* (4, 30, 0) {real, imag} */,
  {32'h4126716e, 32'h41ee3c59} /* (4, 29, 31) {real, imag} */,
  {32'hc12a4cb1, 32'hc13675b7} /* (4, 29, 30) {real, imag} */,
  {32'h4070aadc, 32'h412a09aa} /* (4, 29, 29) {real, imag} */,
  {32'hc0dc7505, 32'hc08ecc45} /* (4, 29, 28) {real, imag} */,
  {32'hc04292dd, 32'h408f6722} /* (4, 29, 27) {real, imag} */,
  {32'hc05ecff1, 32'hc04bc3a7} /* (4, 29, 26) {real, imag} */,
  {32'hc0dc7eec, 32'h3ff1c779} /* (4, 29, 25) {real, imag} */,
  {32'h3eeacea7, 32'h40666f30} /* (4, 29, 24) {real, imag} */,
  {32'h3e7dbd14, 32'hc0474690} /* (4, 29, 23) {real, imag} */,
  {32'hbfe8ce6e, 32'hc0401d89} /* (4, 29, 22) {real, imag} */,
  {32'h4017a4c9, 32'h3e43c503} /* (4, 29, 21) {real, imag} */,
  {32'h3e298183, 32'hbf705d2e} /* (4, 29, 20) {real, imag} */,
  {32'hbe59bacd, 32'h3f974f89} /* (4, 29, 19) {real, imag} */,
  {32'h3e252ff7, 32'h3f64ae63} /* (4, 29, 18) {real, imag} */,
  {32'h3e46ea41, 32'hbf875574} /* (4, 29, 17) {real, imag} */,
  {32'hbf683918, 32'hbe9a769e} /* (4, 29, 16) {real, imag} */,
  {32'h40372d01, 32'hbe775184} /* (4, 29, 15) {real, imag} */,
  {32'h3ef2723d, 32'hbf7fe4c0} /* (4, 29, 14) {real, imag} */,
  {32'h400624bc, 32'h3f88f456} /* (4, 29, 13) {real, imag} */,
  {32'hbf522cae, 32'h3dae6340} /* (4, 29, 12) {real, imag} */,
  {32'h3fc76b7b, 32'hbe575774} /* (4, 29, 11) {real, imag} */,
  {32'h3e92aeaf, 32'h3eb7e8ee} /* (4, 29, 10) {real, imag} */,
  {32'hc050ea24, 32'hbedc8c1e} /* (4, 29, 9) {real, imag} */,
  {32'hc0bfdd3c, 32'hc05eba9f} /* (4, 29, 8) {real, imag} */,
  {32'hc08f357f, 32'h4007a2b1} /* (4, 29, 7) {real, imag} */,
  {32'hc082049d, 32'hc048f17b} /* (4, 29, 6) {real, imag} */,
  {32'h404c7d1a, 32'hc0046f1e} /* (4, 29, 5) {real, imag} */,
  {32'hbda3f672, 32'h4037d2a5} /* (4, 29, 4) {real, imag} */,
  {32'h40f4506e, 32'h3e069131} /* (4, 29, 3) {real, imag} */,
  {32'hc186eb88, 32'hbebe6c21} /* (4, 29, 2) {real, imag} */,
  {32'h41d2b196, 32'hc12aff60} /* (4, 29, 1) {real, imag} */,
  {32'h41336d8d, 32'h3fd50841} /* (4, 29, 0) {real, imag} */,
  {32'h40a15b95, 32'h41b065c4} /* (4, 28, 31) {real, imag} */,
  {32'hc16e7d42, 32'hc179cf63} /* (4, 28, 30) {real, imag} */,
  {32'hc0410f25, 32'hc028b712} /* (4, 28, 29) {real, imag} */,
  {32'hbce8de18, 32'h3f81e48f} /* (4, 28, 28) {real, imag} */,
  {32'hc1020aac, 32'hbf89661c} /* (4, 28, 27) {real, imag} */,
  {32'hbfb7eced, 32'h3f09694d} /* (4, 28, 26) {real, imag} */,
  {32'h3fc16cc6, 32'h3f977432} /* (4, 28, 25) {real, imag} */,
  {32'hbeca6dc6, 32'hbf9f8fc5} /* (4, 28, 24) {real, imag} */,
  {32'hbe0baf7a, 32'h3cd3abdb} /* (4, 28, 23) {real, imag} */,
  {32'h40bc5284, 32'hbf6fab6e} /* (4, 28, 22) {real, imag} */,
  {32'h3fe48a25, 32'h3f42d7c4} /* (4, 28, 21) {real, imag} */,
  {32'h3fc9e7ee, 32'h3ea7d92e} /* (4, 28, 20) {real, imag} */,
  {32'hc03d947f, 32'hbfe8381f} /* (4, 28, 19) {real, imag} */,
  {32'hbf96e9aa, 32'hbe6292da} /* (4, 28, 18) {real, imag} */,
  {32'h3fbd7c0d, 32'h3e24e5dd} /* (4, 28, 17) {real, imag} */,
  {32'h3ed289c6, 32'hbf07dae8} /* (4, 28, 16) {real, imag} */,
  {32'h3e2aa35c, 32'h4018b69e} /* (4, 28, 15) {real, imag} */,
  {32'h408c5787, 32'h402c4799} /* (4, 28, 14) {real, imag} */,
  {32'hbfc0032f, 32'hbf3abadf} /* (4, 28, 13) {real, imag} */,
  {32'h3cb7e85c, 32'hbde5e575} /* (4, 28, 12) {real, imag} */,
  {32'hbfb527e4, 32'hc05f8d07} /* (4, 28, 11) {real, imag} */,
  {32'hbf898d35, 32'hbe88198c} /* (4, 28, 10) {real, imag} */,
  {32'hbf1c108f, 32'hbf4f27e3} /* (4, 28, 9) {real, imag} */,
  {32'h40596cd9, 32'h3e8e15df} /* (4, 28, 8) {real, imag} */,
  {32'hbf2132df, 32'hc01500bc} /* (4, 28, 7) {real, imag} */,
  {32'h3fc8d40f, 32'h3fa9dc95} /* (4, 28, 6) {real, imag} */,
  {32'h3e60b2d4, 32'hc0e4b1be} /* (4, 28, 5) {real, imag} */,
  {32'h40419bd6, 32'h41312b4f} /* (4, 28, 4) {real, imag} */,
  {32'h404aa862, 32'h40e699af} /* (4, 28, 3) {real, imag} */,
  {32'hc06b3588, 32'hc0e44e7e} /* (4, 28, 2) {real, imag} */,
  {32'h408e88b4, 32'h413490eb} /* (4, 28, 1) {real, imag} */,
  {32'h40a1d8c4, 32'h417c9e3a} /* (4, 28, 0) {real, imag} */,
  {32'hc0ea40ea, 32'hc19535ba} /* (4, 27, 31) {real, imag} */,
  {32'h40cd7f53, 32'h40f3b139} /* (4, 27, 30) {real, imag} */,
  {32'hbf62f4c1, 32'h40973345} /* (4, 27, 29) {real, imag} */,
  {32'hc00a00a7, 32'hc08a66ea} /* (4, 27, 28) {real, imag} */,
  {32'h40765dfa, 32'hbfa7e5ad} /* (4, 27, 27) {real, imag} */,
  {32'h3ffe57af, 32'h40869a9c} /* (4, 27, 26) {real, imag} */,
  {32'hc071abe9, 32'hbf16fa45} /* (4, 27, 25) {real, imag} */,
  {32'h3f776bf0, 32'hbec6960d} /* (4, 27, 24) {real, imag} */,
  {32'hbfa30339, 32'hbf3e5da0} /* (4, 27, 23) {real, imag} */,
  {32'h3d86f96f, 32'h3fb6e87d} /* (4, 27, 22) {real, imag} */,
  {32'hbf80a6a5, 32'hbfc6c642} /* (4, 27, 21) {real, imag} */,
  {32'hbfb35aeb, 32'hc0032483} /* (4, 27, 20) {real, imag} */,
  {32'hc00d7367, 32'hbfc30b93} /* (4, 27, 19) {real, imag} */,
  {32'h3e1a312a, 32'hbf2289cd} /* (4, 27, 18) {real, imag} */,
  {32'h3ed1cb8e, 32'hbdf3d72e} /* (4, 27, 17) {real, imag} */,
  {32'h3de246a6, 32'hbf5ff73d} /* (4, 27, 16) {real, imag} */,
  {32'hc003fafc, 32'h3e527bda} /* (4, 27, 15) {real, imag} */,
  {32'hbf79296e, 32'h3f5d4b3e} /* (4, 27, 14) {real, imag} */,
  {32'h3ff7d555, 32'h3f71547f} /* (4, 27, 13) {real, imag} */,
  {32'hbea1c70c, 32'h3f1075dc} /* (4, 27, 12) {real, imag} */,
  {32'hbfdad2b2, 32'h40642c35} /* (4, 27, 11) {real, imag} */,
  {32'hbd8d0dce, 32'h3e6c5352} /* (4, 27, 10) {real, imag} */,
  {32'hbf9a1513, 32'h3feebc8c} /* (4, 27, 9) {real, imag} */,
  {32'h401641df, 32'hbff2230d} /* (4, 27, 8) {real, imag} */,
  {32'hc086ab95, 32'hc0057588} /* (4, 27, 7) {real, imag} */,
  {32'h3f9cfacd, 32'hc08d0954} /* (4, 27, 6) {real, imag} */,
  {32'hc0090f67, 32'h405cf097} /* (4, 27, 5) {real, imag} */,
  {32'hbfd0d1df, 32'h3fd49da7} /* (4, 27, 4) {real, imag} */,
  {32'h3e0df25f, 32'hc040e73f} /* (4, 27, 3) {real, imag} */,
  {32'hc013a504, 32'h40f7df37} /* (4, 27, 2) {real, imag} */,
  {32'h4190779a, 32'hc17d56a4} /* (4, 27, 1) {real, imag} */,
  {32'hc0086bf0, 32'hc1494cfd} /* (4, 27, 0) {real, imag} */,
  {32'h404bd348, 32'hc0ca37ce} /* (4, 26, 31) {real, imag} */,
  {32'h4003a936, 32'h3f0573b5} /* (4, 26, 30) {real, imag} */,
  {32'hbf3c757f, 32'hc00b8af5} /* (4, 26, 29) {real, imag} */,
  {32'h4067b802, 32'h3f3f83c2} /* (4, 26, 28) {real, imag} */,
  {32'h4008468b, 32'hc02fddb2} /* (4, 26, 27) {real, imag} */,
  {32'h3f8ab697, 32'hc0ac9ac2} /* (4, 26, 26) {real, imag} */,
  {32'hbd6a3f72, 32'hbf83627d} /* (4, 26, 25) {real, imag} */,
  {32'h3fb4d835, 32'h3fa88c20} /* (4, 26, 24) {real, imag} */,
  {32'h40886f94, 32'h3c419dbb} /* (4, 26, 23) {real, imag} */,
  {32'hbed0f436, 32'hbf8c1334} /* (4, 26, 22) {real, imag} */,
  {32'h4014f598, 32'hbd655cf5} /* (4, 26, 21) {real, imag} */,
  {32'hbc91c8fe, 32'h3d590fbf} /* (4, 26, 20) {real, imag} */,
  {32'hbf9b09f6, 32'h40307474} /* (4, 26, 19) {real, imag} */,
  {32'h3ffdaa5e, 32'hbfe7c17f} /* (4, 26, 18) {real, imag} */,
  {32'h3f8667fd, 32'hbee1b908} /* (4, 26, 17) {real, imag} */,
  {32'h3e03923d, 32'hbf2037fe} /* (4, 26, 16) {real, imag} */,
  {32'hbfaaf57a, 32'hbfcba35d} /* (4, 26, 15) {real, imag} */,
  {32'h3f34962f, 32'h4002696c} /* (4, 26, 14) {real, imag} */,
  {32'hbfa14995, 32'hbf3d3efb} /* (4, 26, 13) {real, imag} */,
  {32'h3da30289, 32'hbfb2fd23} /* (4, 26, 12) {real, imag} */,
  {32'h3e6cd0c5, 32'hc075163b} /* (4, 26, 11) {real, imag} */,
  {32'hc0110ce3, 32'hbfa5667a} /* (4, 26, 10) {real, imag} */,
  {32'hbfb2c32b, 32'hbf520d4a} /* (4, 26, 9) {real, imag} */,
  {32'h3f0211f4, 32'h409c2a86} /* (4, 26, 8) {real, imag} */,
  {32'h3fdba8df, 32'hbf9f811d} /* (4, 26, 7) {real, imag} */,
  {32'hc01f36e7, 32'hc0cd044a} /* (4, 26, 6) {real, imag} */,
  {32'h40b14066, 32'hbf36719a} /* (4, 26, 5) {real, imag} */,
  {32'h3fce4fd9, 32'hc0a1a0c0} /* (4, 26, 4) {real, imag} */,
  {32'hc049b4a2, 32'h3fb0f998} /* (4, 26, 3) {real, imag} */,
  {32'hc0d9d2fe, 32'h3faef098} /* (4, 26, 2) {real, imag} */,
  {32'h40a5fd73, 32'hbf349049} /* (4, 26, 1) {real, imag} */,
  {32'hc07b48ec, 32'h406f52a1} /* (4, 26, 0) {real, imag} */,
  {32'hbfc898a5, 32'hbeb47eea} /* (4, 25, 31) {real, imag} */,
  {32'hc0c04ffe, 32'h40f9d384} /* (4, 25, 30) {real, imag} */,
  {32'hbfa4ad75, 32'hc04ad35f} /* (4, 25, 29) {real, imag} */,
  {32'h4093fb78, 32'hc01a5ccd} /* (4, 25, 28) {real, imag} */,
  {32'hbed8f2e5, 32'h408304b8} /* (4, 25, 27) {real, imag} */,
  {32'hbfc54346, 32'h3ef1bc8f} /* (4, 25, 26) {real, imag} */,
  {32'hbf5c6220, 32'h402cd9e2} /* (4, 25, 25) {real, imag} */,
  {32'hbea5d736, 32'hbfa83128} /* (4, 25, 24) {real, imag} */,
  {32'hc0113eae, 32'hc00496dc} /* (4, 25, 23) {real, imag} */,
  {32'h3f7fe3ed, 32'h3f6e7884} /* (4, 25, 22) {real, imag} */,
  {32'h4042ee7e, 32'hbf89b3fc} /* (4, 25, 21) {real, imag} */,
  {32'hbfad2662, 32'hbf5561c5} /* (4, 25, 20) {real, imag} */,
  {32'h401700f1, 32'h3e3d275e} /* (4, 25, 19) {real, imag} */,
  {32'h3ffbd4cc, 32'hbf9ae7e2} /* (4, 25, 18) {real, imag} */,
  {32'hbf65ee18, 32'hbea89a25} /* (4, 25, 17) {real, imag} */,
  {32'hbfbae3ba, 32'h3f921620} /* (4, 25, 16) {real, imag} */,
  {32'h3f65dd1f, 32'h3fe18916} /* (4, 25, 15) {real, imag} */,
  {32'hbf9fdfcf, 32'h3fea44b2} /* (4, 25, 14) {real, imag} */,
  {32'h3f3ec830, 32'h4002aa3f} /* (4, 25, 13) {real, imag} */,
  {32'hc05927d5, 32'hbf7b78ed} /* (4, 25, 12) {real, imag} */,
  {32'hbfd1b067, 32'h3f15c220} /* (4, 25, 11) {real, imag} */,
  {32'h3d7dce85, 32'hbf820ad8} /* (4, 25, 10) {real, imag} */,
  {32'hbf83a962, 32'h3ff1c73d} /* (4, 25, 9) {real, imag} */,
  {32'h40b99d2b, 32'h3ef1ebdd} /* (4, 25, 8) {real, imag} */,
  {32'hbe6c13f1, 32'h3f85f4a6} /* (4, 25, 7) {real, imag} */,
  {32'h4044163c, 32'hbfee0c64} /* (4, 25, 6) {real, imag} */,
  {32'hc007cc51, 32'h3f0b0101} /* (4, 25, 5) {real, imag} */,
  {32'hc0190a04, 32'hc093e1ff} /* (4, 25, 4) {real, imag} */,
  {32'hbf62fb5e, 32'h3f417e5a} /* (4, 25, 3) {real, imag} */,
  {32'h407bc3b4, 32'h3f875e90} /* (4, 25, 2) {real, imag} */,
  {32'hc0211cb3, 32'hbfaf36b2} /* (4, 25, 1) {real, imag} */,
  {32'h3f7cb4d9, 32'h3f47fbc3} /* (4, 25, 0) {real, imag} */,
  {32'hc00d24a4, 32'hc101b241} /* (4, 24, 31) {real, imag} */,
  {32'h40759d92, 32'h40060cd3} /* (4, 24, 30) {real, imag} */,
  {32'hc0915586, 32'h3f168c9c} /* (4, 24, 29) {real, imag} */,
  {32'hbf343a0c, 32'hc0081829} /* (4, 24, 28) {real, imag} */,
  {32'h3fc5b72a, 32'hc071f2cf} /* (4, 24, 27) {real, imag} */,
  {32'h3f8e1766, 32'h3fe3016d} /* (4, 24, 26) {real, imag} */,
  {32'h3f9bd4c6, 32'hc03654c3} /* (4, 24, 25) {real, imag} */,
  {32'h3f8547c9, 32'h40693079} /* (4, 24, 24) {real, imag} */,
  {32'h3fd64dd1, 32'hbfbd6146} /* (4, 24, 23) {real, imag} */,
  {32'h3fb29765, 32'hbf84ad9b} /* (4, 24, 22) {real, imag} */,
  {32'h3e3c9fa6, 32'hbe530964} /* (4, 24, 21) {real, imag} */,
  {32'hbe4050e7, 32'hc044ac53} /* (4, 24, 20) {real, imag} */,
  {32'hbf11cd46, 32'h3f3e4a05} /* (4, 24, 19) {real, imag} */,
  {32'hbfaa325b, 32'h3f67f300} /* (4, 24, 18) {real, imag} */,
  {32'h3ef7686a, 32'h3f6e726a} /* (4, 24, 17) {real, imag} */,
  {32'h3f21b1c1, 32'hbe6cb8fa} /* (4, 24, 16) {real, imag} */,
  {32'h3e9fa726, 32'h3f55fb8d} /* (4, 24, 15) {real, imag} */,
  {32'hbf950cb7, 32'hbf5445c4} /* (4, 24, 14) {real, imag} */,
  {32'hbf96b5df, 32'hbda91710} /* (4, 24, 13) {real, imag} */,
  {32'hbf895bd7, 32'hc0bf00b4} /* (4, 24, 12) {real, imag} */,
  {32'hbf381b0a, 32'h3fae6ac5} /* (4, 24, 11) {real, imag} */,
  {32'h3f9e9d57, 32'h408b57d8} /* (4, 24, 10) {real, imag} */,
  {32'h400f1b12, 32'hbf828a35} /* (4, 24, 9) {real, imag} */,
  {32'hc086a581, 32'h4001bf7e} /* (4, 24, 8) {real, imag} */,
  {32'h3ee6ec84, 32'hbf9d4f38} /* (4, 24, 7) {real, imag} */,
  {32'hc043b5d4, 32'h407685ee} /* (4, 24, 6) {real, imag} */,
  {32'h3f9d2b4a, 32'h3e8ca92a} /* (4, 24, 5) {real, imag} */,
  {32'hbe4fb669, 32'hbf1d7811} /* (4, 24, 4) {real, imag} */,
  {32'h3f8464f7, 32'h40250a53} /* (4, 24, 3) {real, imag} */,
  {32'hc06295a1, 32'h40e2f547} /* (4, 24, 2) {real, imag} */,
  {32'hc033ada7, 32'hc1181725} /* (4, 24, 1) {real, imag} */,
  {32'hc06ad888, 32'hc10a298c} /* (4, 24, 0) {real, imag} */,
  {32'h3fc08a5b, 32'h3ed8ee8e} /* (4, 23, 31) {real, imag} */,
  {32'hbfdbd98d, 32'hc096984e} /* (4, 23, 30) {real, imag} */,
  {32'hbe9245e5, 32'hbe3ce781} /* (4, 23, 29) {real, imag} */,
  {32'h403f20da, 32'h3fb4ae58} /* (4, 23, 28) {real, imag} */,
  {32'hc02b0222, 32'h407571a4} /* (4, 23, 27) {real, imag} */,
  {32'hbf56308f, 32'hbf59e19c} /* (4, 23, 26) {real, imag} */,
  {32'hbfe355d0, 32'h3f824fe0} /* (4, 23, 25) {real, imag} */,
  {32'h4018d338, 32'h3dedf27e} /* (4, 23, 24) {real, imag} */,
  {32'h3d9430b5, 32'h400bcfb2} /* (4, 23, 23) {real, imag} */,
  {32'hbfe8a169, 32'hc007d171} /* (4, 23, 22) {real, imag} */,
  {32'hc0075137, 32'h3fac046c} /* (4, 23, 21) {real, imag} */,
  {32'h3f725ddc, 32'h3f7acc24} /* (4, 23, 20) {real, imag} */,
  {32'h401be979, 32'hbcb8ef85} /* (4, 23, 19) {real, imag} */,
  {32'hbdc00a17, 32'h3f973ca5} /* (4, 23, 18) {real, imag} */,
  {32'hbf4532a5, 32'h3eed04ee} /* (4, 23, 17) {real, imag} */,
  {32'h3e915dde, 32'hbf8e01cd} /* (4, 23, 16) {real, imag} */,
  {32'hbf2b41e4, 32'hbfa67a0e} /* (4, 23, 15) {real, imag} */,
  {32'hbe6ef564, 32'hbfd7ff4c} /* (4, 23, 14) {real, imag} */,
  {32'hbf56aca9, 32'h3de6a04d} /* (4, 23, 13) {real, imag} */,
  {32'h3f3b92c7, 32'h40220a1a} /* (4, 23, 12) {real, imag} */,
  {32'h3fed58ce, 32'hc0447b56} /* (4, 23, 11) {real, imag} */,
  {32'h4090b68a, 32'hbf8359d2} /* (4, 23, 10) {real, imag} */,
  {32'hbf74748f, 32'h3e477d9d} /* (4, 23, 9) {real, imag} */,
  {32'h3f005ee1, 32'h3f4ca706} /* (4, 23, 8) {real, imag} */,
  {32'hbfe17dfe, 32'h4049886b} /* (4, 23, 7) {real, imag} */,
  {32'h40218bdc, 32'h40508525} /* (4, 23, 6) {real, imag} */,
  {32'h3ff2e5b3, 32'hc06b8948} /* (4, 23, 5) {real, imag} */,
  {32'h406fcb32, 32'h3fda2b9e} /* (4, 23, 4) {real, imag} */,
  {32'hbf9496ca, 32'hc0534b9f} /* (4, 23, 3) {real, imag} */,
  {32'hc0bce4e9, 32'h3f8af65f} /* (4, 23, 2) {real, imag} */,
  {32'h3fbbb751, 32'h4007a556} /* (4, 23, 1) {real, imag} */,
  {32'h3fe3ee44, 32'h3ffe17a8} /* (4, 23, 0) {real, imag} */,
  {32'h3f259192, 32'h407db59b} /* (4, 22, 31) {real, imag} */,
  {32'hc016a007, 32'hc0274b08} /* (4, 22, 30) {real, imag} */,
  {32'hbdff1f40, 32'hbfa06c05} /* (4, 22, 29) {real, imag} */,
  {32'hbfef864e, 32'h3fc31565} /* (4, 22, 28) {real, imag} */,
  {32'hbff9839d, 32'hbf916e3a} /* (4, 22, 27) {real, imag} */,
  {32'h3d09571e, 32'hc0255b6e} /* (4, 22, 26) {real, imag} */,
  {32'h405249a1, 32'h4020cc01} /* (4, 22, 25) {real, imag} */,
  {32'hbdc5bafa, 32'hbb55281d} /* (4, 22, 24) {real, imag} */,
  {32'h3f80cba6, 32'h40156a34} /* (4, 22, 23) {real, imag} */,
  {32'h3f986544, 32'hbe7c278b} /* (4, 22, 22) {real, imag} */,
  {32'hbfd038b9, 32'h400faeac} /* (4, 22, 21) {real, imag} */,
  {32'h401cf79e, 32'hbf285c0f} /* (4, 22, 20) {real, imag} */,
  {32'h4094ce2b, 32'h3fbe7ced} /* (4, 22, 19) {real, imag} */,
  {32'hbf8fd182, 32'hbf951148} /* (4, 22, 18) {real, imag} */,
  {32'hbf53aca8, 32'h3fa70d84} /* (4, 22, 17) {real, imag} */,
  {32'hbfb34f4c, 32'hbfe62484} /* (4, 22, 16) {real, imag} */,
  {32'hbdc11fc4, 32'hbf3bfa82} /* (4, 22, 15) {real, imag} */,
  {32'hbf81e910, 32'h3eb8b617} /* (4, 22, 14) {real, imag} */,
  {32'h3f4f3e3a, 32'h3f4fc331} /* (4, 22, 13) {real, imag} */,
  {32'h3e43960d, 32'h400e7aaf} /* (4, 22, 12) {real, imag} */,
  {32'hbf7be1d6, 32'hbf10d108} /* (4, 22, 11) {real, imag} */,
  {32'hbf7a2359, 32'hbd5f644c} /* (4, 22, 10) {real, imag} */,
  {32'h3fe45b1b, 32'h40060b1c} /* (4, 22, 9) {real, imag} */,
  {32'hbf615943, 32'h3f1e4c1e} /* (4, 22, 8) {real, imag} */,
  {32'h3f87ae71, 32'h3fa1859e} /* (4, 22, 7) {real, imag} */,
  {32'hbf293d1a, 32'h3f000ad2} /* (4, 22, 6) {real, imag} */,
  {32'hbea40b57, 32'h3ec7b3d3} /* (4, 22, 5) {real, imag} */,
  {32'hc0151e2f, 32'h3fac7fd1} /* (4, 22, 4) {real, imag} */,
  {32'hc034a9ae, 32'h40302868} /* (4, 22, 3) {real, imag} */,
  {32'hc0091ea6, 32'hc093b8e5} /* (4, 22, 2) {real, imag} */,
  {32'hbf99d3ba, 32'h3ffec947} /* (4, 22, 1) {real, imag} */,
  {32'h40543155, 32'hc084879a} /* (4, 22, 0) {real, imag} */,
  {32'hc0051d94, 32'hbf35ab0a} /* (4, 21, 31) {real, imag} */,
  {32'h40c0dc4f, 32'h3f9f0f44} /* (4, 21, 30) {real, imag} */,
  {32'hc04f1c07, 32'h4036eb5b} /* (4, 21, 29) {real, imag} */,
  {32'h3eb89dd4, 32'hbfae0401} /* (4, 21, 28) {real, imag} */,
  {32'h3fa39311, 32'h3fde37c0} /* (4, 21, 27) {real, imag} */,
  {32'h3fd26cdd, 32'hbee3638e} /* (4, 21, 26) {real, imag} */,
  {32'hbfaae917, 32'h3feacbf7} /* (4, 21, 25) {real, imag} */,
  {32'hbfc44395, 32'hbfda59d4} /* (4, 21, 24) {real, imag} */,
  {32'hbf6393ad, 32'h3e6df008} /* (4, 21, 23) {real, imag} */,
  {32'hc02e8fb9, 32'hbfe48fbe} /* (4, 21, 22) {real, imag} */,
  {32'h3f410f8f, 32'hbfccda4c} /* (4, 21, 21) {real, imag} */,
  {32'h3f889bbf, 32'h3f68d333} /* (4, 21, 20) {real, imag} */,
  {32'hbdc93c18, 32'h4004bc1d} /* (4, 21, 19) {real, imag} */,
  {32'hbf1eaf87, 32'hbe5fe6a5} /* (4, 21, 18) {real, imag} */,
  {32'h3f46a2fc, 32'hbebaa2ea} /* (4, 21, 17) {real, imag} */,
  {32'h4002c145, 32'hbf8097bc} /* (4, 21, 16) {real, imag} */,
  {32'hbf753314, 32'hbf3db492} /* (4, 21, 15) {real, imag} */,
  {32'h3fa259a1, 32'hbdb93eac} /* (4, 21, 14) {real, imag} */,
  {32'hbfadf3d0, 32'h3edcdb93} /* (4, 21, 13) {real, imag} */,
  {32'h3f361cfc, 32'hbd976a36} /* (4, 21, 12) {real, imag} */,
  {32'h3f460a39, 32'h3f961da7} /* (4, 21, 11) {real, imag} */,
  {32'hbfc42222, 32'hc008b443} /* (4, 21, 10) {real, imag} */,
  {32'h3fd9ee66, 32'h3f8666b2} /* (4, 21, 9) {real, imag} */,
  {32'h3f954a1a, 32'hbf63330c} /* (4, 21, 8) {real, imag} */,
  {32'hbf6abe51, 32'hc014c4ec} /* (4, 21, 7) {real, imag} */,
  {32'h400d1ccf, 32'h3f8bb339} /* (4, 21, 6) {real, imag} */,
  {32'hbf66046e, 32'h4053d3b8} /* (4, 21, 5) {real, imag} */,
  {32'h3eaa5dea, 32'hbedd1316} /* (4, 21, 4) {real, imag} */,
  {32'h3f9d6471, 32'hbff2dbb8} /* (4, 21, 3) {real, imag} */,
  {32'h409380a9, 32'h3fb45ca5} /* (4, 21, 2) {real, imag} */,
  {32'h3e8e9075, 32'hc02e9585} /* (4, 21, 1) {real, imag} */,
  {32'hc07c47e9, 32'hbff5a1a6} /* (4, 21, 0) {real, imag} */,
  {32'h3fdcc14b, 32'h3f74f1d0} /* (4, 20, 31) {real, imag} */,
  {32'h3d949bd2, 32'h3bee8f8e} /* (4, 20, 30) {real, imag} */,
  {32'hc0042199, 32'h3f5184f1} /* (4, 20, 29) {real, imag} */,
  {32'hbea3befb, 32'h3fa656d9} /* (4, 20, 28) {real, imag} */,
  {32'h3ef08dde, 32'hc019db4d} /* (4, 20, 27) {real, imag} */,
  {32'h3eab286a, 32'h3f2544bb} /* (4, 20, 26) {real, imag} */,
  {32'h3f739bd8, 32'h3f188815} /* (4, 20, 25) {real, imag} */,
  {32'h400f024b, 32'hbff883ce} /* (4, 20, 24) {real, imag} */,
  {32'hbe28b58f, 32'h400019a5} /* (4, 20, 23) {real, imag} */,
  {32'h3edee188, 32'hbf05d50b} /* (4, 20, 22) {real, imag} */,
  {32'h3f67886f, 32'hbf1a4157} /* (4, 20, 21) {real, imag} */,
  {32'hbe6fa3bd, 32'h3fca008a} /* (4, 20, 20) {real, imag} */,
  {32'hc013395a, 32'h3d89b6b4} /* (4, 20, 19) {real, imag} */,
  {32'hbecf1ed3, 32'hbfae31a9} /* (4, 20, 18) {real, imag} */,
  {32'hbf67c15b, 32'hbfc19cb2} /* (4, 20, 17) {real, imag} */,
  {32'h3e37ef9b, 32'h3f34faff} /* (4, 20, 16) {real, imag} */,
  {32'hbf821d3a, 32'h40069c22} /* (4, 20, 15) {real, imag} */,
  {32'hbf82f9b1, 32'hbfe4f536} /* (4, 20, 14) {real, imag} */,
  {32'h3efeeb6c, 32'hbf9adfa3} /* (4, 20, 13) {real, imag} */,
  {32'hbf3aabaa, 32'hbfda90ef} /* (4, 20, 12) {real, imag} */,
  {32'hbf8dd9c4, 32'h40870963} /* (4, 20, 11) {real, imag} */,
  {32'h3e3f72ee, 32'hc062eba9} /* (4, 20, 10) {real, imag} */,
  {32'h3e8816dc, 32'hbfdefc0e} /* (4, 20, 9) {real, imag} */,
  {32'hc04e99ef, 32'h3eed9636} /* (4, 20, 8) {real, imag} */,
  {32'h3f9e3dd2, 32'hbfee0a6d} /* (4, 20, 7) {real, imag} */,
  {32'h3f7f1770, 32'h3f345bd5} /* (4, 20, 6) {real, imag} */,
  {32'hbfbbe502, 32'h40897102} /* (4, 20, 5) {real, imag} */,
  {32'hbf755ca4, 32'h3f000153} /* (4, 20, 4) {real, imag} */,
  {32'hbe27ba99, 32'h3ff2296a} /* (4, 20, 3) {real, imag} */,
  {32'h40bc88b1, 32'h3e268ad9} /* (4, 20, 2) {real, imag} */,
  {32'hbfa8047c, 32'hbef544d3} /* (4, 20, 1) {real, imag} */,
  {32'h3fb6509d, 32'hbf696db0} /* (4, 20, 0) {real, imag} */,
  {32'hbef4a09f, 32'h3fca3657} /* (4, 19, 31) {real, imag} */,
  {32'hc00da3dc, 32'h3f36a67a} /* (4, 19, 30) {real, imag} */,
  {32'h3fc24f4e, 32'hbfa47113} /* (4, 19, 29) {real, imag} */,
  {32'hc00c3bdd, 32'h40302fe4} /* (4, 19, 28) {real, imag} */,
  {32'hbe67c916, 32'hc029b02b} /* (4, 19, 27) {real, imag} */,
  {32'h3fffb60f, 32'h3e7dc6a3} /* (4, 19, 26) {real, imag} */,
  {32'h3ee2c745, 32'hbfc1ff86} /* (4, 19, 25) {real, imag} */,
  {32'h40294e46, 32'h3fb07ec8} /* (4, 19, 24) {real, imag} */,
  {32'hbfad25c9, 32'h3e5592be} /* (4, 19, 23) {real, imag} */,
  {32'h40131133, 32'hc02efde6} /* (4, 19, 22) {real, imag} */,
  {32'hbf88ba7f, 32'hbf088d20} /* (4, 19, 21) {real, imag} */,
  {32'hbf5dde6c, 32'hbf941aa6} /* (4, 19, 20) {real, imag} */,
  {32'h3f3f18fb, 32'h3e6f160f} /* (4, 19, 19) {real, imag} */,
  {32'hbf102b24, 32'h3f152220} /* (4, 19, 18) {real, imag} */,
  {32'h3cac67e2, 32'hbfc7db63} /* (4, 19, 17) {real, imag} */,
  {32'h3fb101cf, 32'h3fa4a6c9} /* (4, 19, 16) {real, imag} */,
  {32'h3f4429b5, 32'hc0079742} /* (4, 19, 15) {real, imag} */,
  {32'hbd266330, 32'hc035c5fe} /* (4, 19, 14) {real, imag} */,
  {32'hbfe6bcb7, 32'hbff972b2} /* (4, 19, 13) {real, imag} */,
  {32'h3f27f2e7, 32'h3facb6c2} /* (4, 19, 12) {real, imag} */,
  {32'hc04d0ace, 32'h3fa85cf0} /* (4, 19, 11) {real, imag} */,
  {32'hc062d755, 32'hbe1e31f1} /* (4, 19, 10) {real, imag} */,
  {32'hbfa7f3cf, 32'h3ea60e71} /* (4, 19, 9) {real, imag} */,
  {32'h3f73c722, 32'hbef1a336} /* (4, 19, 8) {real, imag} */,
  {32'hbdab9ef6, 32'hc00014be} /* (4, 19, 7) {real, imag} */,
  {32'h3e1c28c6, 32'h3eefc298} /* (4, 19, 6) {real, imag} */,
  {32'h3f8141f3, 32'hbf1408c6} /* (4, 19, 5) {real, imag} */,
  {32'hbea29449, 32'h3dda5533} /* (4, 19, 4) {real, imag} */,
  {32'h400f4878, 32'hbdf6281b} /* (4, 19, 3) {real, imag} */,
  {32'hbfaccff6, 32'hc000a4f2} /* (4, 19, 2) {real, imag} */,
  {32'h3f688ae3, 32'hbe3dc453} /* (4, 19, 1) {real, imag} */,
  {32'h40045fad, 32'h3e991342} /* (4, 19, 0) {real, imag} */,
  {32'h3fca307f, 32'hbfbdda2e} /* (4, 18, 31) {real, imag} */,
  {32'h3fa3cd07, 32'h4016d243} /* (4, 18, 30) {real, imag} */,
  {32'h3e68014d, 32'h3f598c1b} /* (4, 18, 29) {real, imag} */,
  {32'h3fb010b0, 32'hbfb3d69d} /* (4, 18, 28) {real, imag} */,
  {32'h3fca4511, 32'h3e05e599} /* (4, 18, 27) {real, imag} */,
  {32'h4004e3e8, 32'h3f86bcbb} /* (4, 18, 26) {real, imag} */,
  {32'h3fa76325, 32'hbef3c4a4} /* (4, 18, 25) {real, imag} */,
  {32'hc00bd9ee, 32'h3fb58b4f} /* (4, 18, 24) {real, imag} */,
  {32'h3e49b43e, 32'h3fa1dd08} /* (4, 18, 23) {real, imag} */,
  {32'hc0860799, 32'h400489ba} /* (4, 18, 22) {real, imag} */,
  {32'h3fad8327, 32'h3efa426b} /* (4, 18, 21) {real, imag} */,
  {32'hbedcaa5c, 32'hbb0eee0e} /* (4, 18, 20) {real, imag} */,
  {32'hbf4c7723, 32'h3a48f653} /* (4, 18, 19) {real, imag} */,
  {32'h3eb626c5, 32'hbe86404b} /* (4, 18, 18) {real, imag} */,
  {32'hbfe3c94a, 32'h3fbf7c80} /* (4, 18, 17) {real, imag} */,
  {32'hbef04334, 32'hbf2a949e} /* (4, 18, 16) {real, imag} */,
  {32'hbefd2816, 32'hbf967e08} /* (4, 18, 15) {real, imag} */,
  {32'hbf592ffd, 32'hbfc0e1fe} /* (4, 18, 14) {real, imag} */,
  {32'h3fae4ff7, 32'h3f3577d2} /* (4, 18, 13) {real, imag} */,
  {32'h3fa61d56, 32'hbf7ec496} /* (4, 18, 12) {real, imag} */,
  {32'hbf6df43c, 32'hbf4a3cee} /* (4, 18, 11) {real, imag} */,
  {32'h3f592577, 32'hbfe4b1a7} /* (4, 18, 10) {real, imag} */,
  {32'h3f605405, 32'hbf1c6036} /* (4, 18, 9) {real, imag} */,
  {32'hbfd0d80c, 32'hbfb14802} /* (4, 18, 8) {real, imag} */,
  {32'hc0086ae4, 32'h3ca2f146} /* (4, 18, 7) {real, imag} */,
  {32'h4049f721, 32'h4029a84b} /* (4, 18, 6) {real, imag} */,
  {32'hbf0ff506, 32'hbe44634e} /* (4, 18, 5) {real, imag} */,
  {32'h3fb08d51, 32'h3ed99a26} /* (4, 18, 4) {real, imag} */,
  {32'h3eb087c5, 32'hbf4a781b} /* (4, 18, 3) {real, imag} */,
  {32'h3f56b248, 32'hbf09a328} /* (4, 18, 2) {real, imag} */,
  {32'hc03c3619, 32'hbe7b98e0} /* (4, 18, 1) {real, imag} */,
  {32'hc005dcf7, 32'hbfb4b309} /* (4, 18, 0) {real, imag} */,
  {32'h3fc3e42c, 32'h3fc2cb7c} /* (4, 17, 31) {real, imag} */,
  {32'h3e59ecb7, 32'hbe6440db} /* (4, 17, 30) {real, imag} */,
  {32'hbf3ecba7, 32'hc00aa8f8} /* (4, 17, 29) {real, imag} */,
  {32'h3ed3c0ac, 32'hbf3dac7a} /* (4, 17, 28) {real, imag} */,
  {32'hbf0a152e, 32'hbfad6811} /* (4, 17, 27) {real, imag} */,
  {32'hbf82e25e, 32'hbf10b3a4} /* (4, 17, 26) {real, imag} */,
  {32'hbf196f37, 32'hbffc4fae} /* (4, 17, 25) {real, imag} */,
  {32'hbf7745af, 32'h3ff7a638} /* (4, 17, 24) {real, imag} */,
  {32'hbf3f8b0a, 32'h3f3f2702} /* (4, 17, 23) {real, imag} */,
  {32'hbf0e2b04, 32'hbd0994f6} /* (4, 17, 22) {real, imag} */,
  {32'h404229c2, 32'h3fa0d16e} /* (4, 17, 21) {real, imag} */,
  {32'hbfc733b5, 32'h40115872} /* (4, 17, 20) {real, imag} */,
  {32'h3f91208b, 32'hbf22029b} /* (4, 17, 19) {real, imag} */,
  {32'h4001c6a2, 32'hbe763e3b} /* (4, 17, 18) {real, imag} */,
  {32'h3f8b5662, 32'h3f0a91bf} /* (4, 17, 17) {real, imag} */,
  {32'hbf122511, 32'h3e048ea5} /* (4, 17, 16) {real, imag} */,
  {32'h3e2a55a6, 32'h3fff8c82} /* (4, 17, 15) {real, imag} */,
  {32'h3f5526f6, 32'hbf821958} /* (4, 17, 14) {real, imag} */,
  {32'hbf9b01ae, 32'hc036f703} /* (4, 17, 13) {real, imag} */,
  {32'h403a495f, 32'hbecd2344} /* (4, 17, 12) {real, imag} */,
  {32'hbf8012fb, 32'h3c47e3f0} /* (4, 17, 11) {real, imag} */,
  {32'hbe418edc, 32'h3e99a965} /* (4, 17, 10) {real, imag} */,
  {32'h3e5f8b0b, 32'h3f688ebb} /* (4, 17, 9) {real, imag} */,
  {32'hbf3065bf, 32'h40016621} /* (4, 17, 8) {real, imag} */,
  {32'hbec7a204, 32'hbf89ccdb} /* (4, 17, 7) {real, imag} */,
  {32'h3f327ca8, 32'hc024a8df} /* (4, 17, 6) {real, imag} */,
  {32'h3fc3441b, 32'h3e2c2713} /* (4, 17, 5) {real, imag} */,
  {32'h3f63d961, 32'hbf19b2ff} /* (4, 17, 4) {real, imag} */,
  {32'h3d848438, 32'h4039de8b} /* (4, 17, 3) {real, imag} */,
  {32'h3ee56730, 32'h3effec71} /* (4, 17, 2) {real, imag} */,
  {32'h3e5a6c8d, 32'h3f060890} /* (4, 17, 1) {real, imag} */,
  {32'hbf08f434, 32'hbfba38b5} /* (4, 17, 0) {real, imag} */,
  {32'h3f8bdc65, 32'h3e5370ba} /* (4, 16, 31) {real, imag} */,
  {32'h3f28950c, 32'hbf570baa} /* (4, 16, 30) {real, imag} */,
  {32'h3f2903c2, 32'h3f9093d9} /* (4, 16, 29) {real, imag} */,
  {32'hbe801ac5, 32'hbfcb0508} /* (4, 16, 28) {real, imag} */,
  {32'hc01ec4fc, 32'hbe0bfe47} /* (4, 16, 27) {real, imag} */,
  {32'h3e9da2f0, 32'h3f97e984} /* (4, 16, 26) {real, imag} */,
  {32'hbf1b103a, 32'h3f7b277d} /* (4, 16, 25) {real, imag} */,
  {32'hbed18232, 32'h3fe10177} /* (4, 16, 24) {real, imag} */,
  {32'hbfdab5c0, 32'h3f46d0d0} /* (4, 16, 23) {real, imag} */,
  {32'hbf396cf8, 32'h3f0e0552} /* (4, 16, 22) {real, imag} */,
  {32'h3f8ce44b, 32'h3ed93c86} /* (4, 16, 21) {real, imag} */,
  {32'h3ef5c42d, 32'hbf0f674e} /* (4, 16, 20) {real, imag} */,
  {32'hbf4c0294, 32'h3fd08ae6} /* (4, 16, 19) {real, imag} */,
  {32'hbf725fc5, 32'h3f20023e} /* (4, 16, 18) {real, imag} */,
  {32'hbec9877e, 32'h3f0025e6} /* (4, 16, 17) {real, imag} */,
  {32'h3fe78f22, 32'hbe1ab163} /* (4, 16, 16) {real, imag} */,
  {32'hbf7ede65, 32'h3ee7d674} /* (4, 16, 15) {real, imag} */,
  {32'hbeed59e9, 32'h3f80281e} /* (4, 16, 14) {real, imag} */,
  {32'h4081afce, 32'h3d3b0c5a} /* (4, 16, 13) {real, imag} */,
  {32'hbf88156e, 32'hbf0def1b} /* (4, 16, 12) {real, imag} */,
  {32'hbea221ad, 32'h3fb4d365} /* (4, 16, 11) {real, imag} */,
  {32'hbfa080e5, 32'h3d167db6} /* (4, 16, 10) {real, imag} */,
  {32'hbf398267, 32'h3ee7af6c} /* (4, 16, 9) {real, imag} */,
  {32'hbecb4894, 32'hbf22b414} /* (4, 16, 8) {real, imag} */,
  {32'h3f7db075, 32'hbefd1ba0} /* (4, 16, 7) {real, imag} */,
  {32'h3f56260f, 32'hbfd88531} /* (4, 16, 6) {real, imag} */,
  {32'hbf9d87b4, 32'h3f84030d} /* (4, 16, 5) {real, imag} */,
  {32'h3ec8e32e, 32'hbff0ef53} /* (4, 16, 4) {real, imag} */,
  {32'hbfbf0126, 32'hbddf52d8} /* (4, 16, 3) {real, imag} */,
  {32'h3e42b288, 32'h3f7ec8a6} /* (4, 16, 2) {real, imag} */,
  {32'h3f80c595, 32'h3dcc2d01} /* (4, 16, 1) {real, imag} */,
  {32'h3eed3bdf, 32'h400b8bd5} /* (4, 16, 0) {real, imag} */,
  {32'hbf87b66a, 32'h3efe4a66} /* (4, 15, 31) {real, imag} */,
  {32'hbbe311d7, 32'h3fdaf243} /* (4, 15, 30) {real, imag} */,
  {32'hbffec727, 32'hbf46a8ca} /* (4, 15, 29) {real, imag} */,
  {32'hbfd98c37, 32'hbfb5c1c8} /* (4, 15, 28) {real, imag} */,
  {32'hbdbafa89, 32'hbe7414e9} /* (4, 15, 27) {real, imag} */,
  {32'hbed24904, 32'h3fe19913} /* (4, 15, 26) {real, imag} */,
  {32'h40135186, 32'h3ee14e64} /* (4, 15, 25) {real, imag} */,
  {32'h40055808, 32'hc05cbc06} /* (4, 15, 24) {real, imag} */,
  {32'h402cf4dd, 32'hbfb6b210} /* (4, 15, 23) {real, imag} */,
  {32'h401e2b6b, 32'hbf894a5b} /* (4, 15, 22) {real, imag} */,
  {32'hc04aa4cd, 32'h3ebac52c} /* (4, 15, 21) {real, imag} */,
  {32'h3f87d565, 32'hbeb2f728} /* (4, 15, 20) {real, imag} */,
  {32'hbf73d121, 32'h3f3d37b4} /* (4, 15, 19) {real, imag} */,
  {32'hbe6842a6, 32'h3f457f54} /* (4, 15, 18) {real, imag} */,
  {32'h3f409de2, 32'hbf167e35} /* (4, 15, 17) {real, imag} */,
  {32'h3e0acbf8, 32'h3f65d9f9} /* (4, 15, 16) {real, imag} */,
  {32'hbea641d3, 32'h3e640677} /* (4, 15, 15) {real, imag} */,
  {32'h3f961a3c, 32'h3db313d7} /* (4, 15, 14) {real, imag} */,
  {32'hbd5395de, 32'hbe1762d0} /* (4, 15, 13) {real, imag} */,
  {32'hbf903a61, 32'h3fb553b8} /* (4, 15, 12) {real, imag} */,
  {32'hc0368fb0, 32'h3f6474a6} /* (4, 15, 11) {real, imag} */,
  {32'h3ee306df, 32'h3f27ed57} /* (4, 15, 10) {real, imag} */,
  {32'h3f151b3b, 32'hbfc36ca2} /* (4, 15, 9) {real, imag} */,
  {32'h3ea2a18d, 32'hbefc9787} /* (4, 15, 8) {real, imag} */,
  {32'h3c9643d8, 32'hbfe3e0e6} /* (4, 15, 7) {real, imag} */,
  {32'h3fb8d515, 32'h3e82569d} /* (4, 15, 6) {real, imag} */,
  {32'h401137b3, 32'hbf613839} /* (4, 15, 5) {real, imag} */,
  {32'h3eb495c8, 32'h3feaef46} /* (4, 15, 4) {real, imag} */,
  {32'hbfbe30fe, 32'h3f9ebfcb} /* (4, 15, 3) {real, imag} */,
  {32'h3fa858cf, 32'h3f1f03ce} /* (4, 15, 2) {real, imag} */,
  {32'hc0280c4c, 32'h3f7324ec} /* (4, 15, 1) {real, imag} */,
  {32'hbf3a5c64, 32'hbe20f418} /* (4, 15, 0) {real, imag} */,
  {32'h406aaa4d, 32'hbcc1166d} /* (4, 14, 31) {real, imag} */,
  {32'h3ea12fab, 32'h3edc24e4} /* (4, 14, 30) {real, imag} */,
  {32'h3df86fb8, 32'hbefed998} /* (4, 14, 29) {real, imag} */,
  {32'h3f3f8812, 32'hbfb52800} /* (4, 14, 28) {real, imag} */,
  {32'hbf429b73, 32'h3f99c2f2} /* (4, 14, 27) {real, imag} */,
  {32'h3f936fc2, 32'h3f4bcd87} /* (4, 14, 26) {real, imag} */,
  {32'h3fd8eca4, 32'h3fcd1dbc} /* (4, 14, 25) {real, imag} */,
  {32'h4006a048, 32'hbfc98b95} /* (4, 14, 24) {real, imag} */,
  {32'hbe109740, 32'h3f85c466} /* (4, 14, 23) {real, imag} */,
  {32'hbdbb1c14, 32'hc0111c92} /* (4, 14, 22) {real, imag} */,
  {32'h3e568f5f, 32'hbfa77a38} /* (4, 14, 21) {real, imag} */,
  {32'hc01cc6df, 32'hbee0d517} /* (4, 14, 20) {real, imag} */,
  {32'h3f1d784c, 32'hc04af479} /* (4, 14, 19) {real, imag} */,
  {32'hbed61d58, 32'h401dd523} /* (4, 14, 18) {real, imag} */,
  {32'h3f6c66c8, 32'h3f4480bf} /* (4, 14, 17) {real, imag} */,
  {32'hbe5e5c07, 32'h3f9c8951} /* (4, 14, 16) {real, imag} */,
  {32'hbe022f65, 32'hbf97ca49} /* (4, 14, 15) {real, imag} */,
  {32'hbf866575, 32'h3fad2587} /* (4, 14, 14) {real, imag} */,
  {32'hbe66f262, 32'h3e86946a} /* (4, 14, 13) {real, imag} */,
  {32'hbd977b99, 32'h3f9d261e} /* (4, 14, 12) {real, imag} */,
  {32'h3f8bd469, 32'hbfbb5965} /* (4, 14, 11) {real, imag} */,
  {32'h3eb7f41c, 32'hbcefc3b4} /* (4, 14, 10) {real, imag} */,
  {32'hbedd9ac7, 32'hbfd1f8a1} /* (4, 14, 9) {real, imag} */,
  {32'h3f3ad753, 32'h3ff10793} /* (4, 14, 8) {real, imag} */,
  {32'hbfa0eee2, 32'hbfbebaf4} /* (4, 14, 7) {real, imag} */,
  {32'h3f346962, 32'h3fb2f3de} /* (4, 14, 6) {real, imag} */,
  {32'hbf6b610f, 32'hbe07c57b} /* (4, 14, 5) {real, imag} */,
  {32'h4004934f, 32'hbec8a8a7} /* (4, 14, 4) {real, imag} */,
  {32'hbf39dee9, 32'h3ec0741f} /* (4, 14, 3) {real, imag} */,
  {32'hbfcc131c, 32'hc03b753b} /* (4, 14, 2) {real, imag} */,
  {32'h40120b7d, 32'h3f98c784} /* (4, 14, 1) {real, imag} */,
  {32'h3f1919b1, 32'h3f808e9d} /* (4, 14, 0) {real, imag} */,
  {32'hbf65a805, 32'h3ff3f9d9} /* (4, 13, 31) {real, imag} */,
  {32'hbf1d4bd3, 32'hc016b9e6} /* (4, 13, 30) {real, imag} */,
  {32'hbf1ecc27, 32'h3fc87f04} /* (4, 13, 29) {real, imag} */,
  {32'h3f78986a, 32'h4015b7f5} /* (4, 13, 28) {real, imag} */,
  {32'h40141f80, 32'hbda45921} /* (4, 13, 27) {real, imag} */,
  {32'h401fb089, 32'h3f1e214c} /* (4, 13, 26) {real, imag} */,
  {32'hbfb1c963, 32'h40068f93} /* (4, 13, 25) {real, imag} */,
  {32'hbfc082c6, 32'h3f1ab088} /* (4, 13, 24) {real, imag} */,
  {32'h3fde985b, 32'hbf9cd431} /* (4, 13, 23) {real, imag} */,
  {32'hbee0fcef, 32'h3edf8e08} /* (4, 13, 22) {real, imag} */,
  {32'h3ee85fa3, 32'hbf3ec0ee} /* (4, 13, 21) {real, imag} */,
  {32'h3fb17dbc, 32'h4018ef63} /* (4, 13, 20) {real, imag} */,
  {32'h4042099e, 32'h3e289413} /* (4, 13, 19) {real, imag} */,
  {32'hbfe522f8, 32'hbf5e7995} /* (4, 13, 18) {real, imag} */,
  {32'h3f9c8e31, 32'hbf288f64} /* (4, 13, 17) {real, imag} */,
  {32'hbf27cf22, 32'h3df7ec96} /* (4, 13, 16) {real, imag} */,
  {32'hbe772da3, 32'hbe353280} /* (4, 13, 15) {real, imag} */,
  {32'hbf9b55bb, 32'h3f9daa51} /* (4, 13, 14) {real, imag} */,
  {32'hc030a9ad, 32'hbf8f6d84} /* (4, 13, 13) {real, imag} */,
  {32'hbf064ecb, 32'hbee8d718} /* (4, 13, 12) {real, imag} */,
  {32'hbe9f51ec, 32'h3fe79158} /* (4, 13, 11) {real, imag} */,
  {32'h40218688, 32'hbfbdd1bb} /* (4, 13, 10) {real, imag} */,
  {32'h3f7a5be0, 32'h3fa86078} /* (4, 13, 9) {real, imag} */,
  {32'h3f0f6814, 32'hc084fc28} /* (4, 13, 8) {real, imag} */,
  {32'h3d8b5bc7, 32'h3fc0aa81} /* (4, 13, 7) {real, imag} */,
  {32'h3f028175, 32'h4013c14d} /* (4, 13, 6) {real, imag} */,
  {32'h3cadb9ef, 32'hc0055e28} /* (4, 13, 5) {real, imag} */,
  {32'hbf62b581, 32'h3faed179} /* (4, 13, 4) {real, imag} */,
  {32'hbf1ff6c6, 32'h3f80295a} /* (4, 13, 3) {real, imag} */,
  {32'h3fb96083, 32'h3fc575ea} /* (4, 13, 2) {real, imag} */,
  {32'hbf0e1e0f, 32'h4050aff7} /* (4, 13, 1) {real, imag} */,
  {32'hc0425d6b, 32'hbfe00a38} /* (4, 13, 0) {real, imag} */,
  {32'hbffc1300, 32'hc02dc558} /* (4, 12, 31) {real, imag} */,
  {32'h3ef65f3d, 32'h3f86f31e} /* (4, 12, 30) {real, imag} */,
  {32'h3f42e556, 32'h3f82ff4a} /* (4, 12, 29) {real, imag} */,
  {32'h3f7c320e, 32'h3edc4408} /* (4, 12, 28) {real, imag} */,
  {32'h3fa5ec41, 32'hc04a4e62} /* (4, 12, 27) {real, imag} */,
  {32'h40779d32, 32'hc010010f} /* (4, 12, 26) {real, imag} */,
  {32'h3e7b1165, 32'h3fd58dc4} /* (4, 12, 25) {real, imag} */,
  {32'hbf78c178, 32'h3e8ca19c} /* (4, 12, 24) {real, imag} */,
  {32'hbfbcc756, 32'h3fdde237} /* (4, 12, 23) {real, imag} */,
  {32'h3f586bce, 32'h4078b071} /* (4, 12, 22) {real, imag} */,
  {32'h3bbadd0d, 32'h401a1c67} /* (4, 12, 21) {real, imag} */,
  {32'hbf552a95, 32'hc0302acb} /* (4, 12, 20) {real, imag} */,
  {32'hbe78b5c1, 32'h3f934bfd} /* (4, 12, 19) {real, imag} */,
  {32'h40626763, 32'hbfef22a7} /* (4, 12, 18) {real, imag} */,
  {32'h3eef6f5d, 32'h3e6644e1} /* (4, 12, 17) {real, imag} */,
  {32'hbe964693, 32'h3eb3a858} /* (4, 12, 16) {real, imag} */,
  {32'h3f55c58d, 32'h3f309354} /* (4, 12, 15) {real, imag} */,
  {32'h3e9b48bb, 32'h3f98a939} /* (4, 12, 14) {real, imag} */,
  {32'hc058fdfb, 32'h3eee7a83} /* (4, 12, 13) {real, imag} */,
  {32'h3fbd91ce, 32'hbf6e707b} /* (4, 12, 12) {real, imag} */,
  {32'hbf99036f, 32'hc01aa869} /* (4, 12, 11) {real, imag} */,
  {32'hbfbcf0f3, 32'hbf2330dd} /* (4, 12, 10) {real, imag} */,
  {32'hc088eacb, 32'h3d97ce63} /* (4, 12, 9) {real, imag} */,
  {32'hc00fffcc, 32'hc025d88e} /* (4, 12, 8) {real, imag} */,
  {32'hbffe9a14, 32'h402ce580} /* (4, 12, 7) {real, imag} */,
  {32'hbc3e84f3, 32'h4002bc8d} /* (4, 12, 6) {real, imag} */,
  {32'hbf852eeb, 32'h3d06574a} /* (4, 12, 5) {real, imag} */,
  {32'h3fdf9347, 32'h3f946c9a} /* (4, 12, 4) {real, imag} */,
  {32'hbf90858b, 32'hbf8ea72a} /* (4, 12, 3) {real, imag} */,
  {32'h3fb774e4, 32'hc01b53b4} /* (4, 12, 2) {real, imag} */,
  {32'hbee8cee5, 32'hbf0ae55e} /* (4, 12, 1) {real, imag} */,
  {32'hbfafaf59, 32'hbf5bf710} /* (4, 12, 0) {real, imag} */,
  {32'h40240363, 32'hbf850734} /* (4, 11, 31) {real, imag} */,
  {32'hc0861605, 32'hbfbec722} /* (4, 11, 30) {real, imag} */,
  {32'hbfa6b8fc, 32'h3fcadd48} /* (4, 11, 29) {real, imag} */,
  {32'h3fdc3e72, 32'hbe560e89} /* (4, 11, 28) {real, imag} */,
  {32'h3e497105, 32'hbf7572ce} /* (4, 11, 27) {real, imag} */,
  {32'h40077799, 32'hbf744a58} /* (4, 11, 26) {real, imag} */,
  {32'hbea05ad5, 32'hbff3b3f2} /* (4, 11, 25) {real, imag} */,
  {32'h3edb81f1, 32'h4027934f} /* (4, 11, 24) {real, imag} */,
  {32'hc00263a9, 32'h3f942af2} /* (4, 11, 23) {real, imag} */,
  {32'h40466326, 32'hbf41948e} /* (4, 11, 22) {real, imag} */,
  {32'hbfe79f49, 32'hbf2e9dae} /* (4, 11, 21) {real, imag} */,
  {32'hc037db67, 32'h408292dd} /* (4, 11, 20) {real, imag} */,
  {32'hc04fcb4b, 32'hbff1e093} /* (4, 11, 19) {real, imag} */,
  {32'h3f74bc0c, 32'h3fc3120b} /* (4, 11, 18) {real, imag} */,
  {32'hbfc589fc, 32'hbf3ecad1} /* (4, 11, 17) {real, imag} */,
  {32'h3f8cec99, 32'hbf99b96d} /* (4, 11, 16) {real, imag} */,
  {32'h3f2627b6, 32'h401232d7} /* (4, 11, 15) {real, imag} */,
  {32'hc00a2132, 32'hbfb66002} /* (4, 11, 14) {real, imag} */,
  {32'hc021da80, 32'h3f246f60} /* (4, 11, 13) {real, imag} */,
  {32'h3cba5a73, 32'h3d0167f2} /* (4, 11, 12) {real, imag} */,
  {32'h3fbac362, 32'hbec6f49a} /* (4, 11, 11) {real, imag} */,
  {32'hbf3438c4, 32'h40605f69} /* (4, 11, 10) {real, imag} */,
  {32'hbfa176fe, 32'h3fb0bf3e} /* (4, 11, 9) {real, imag} */,
  {32'hbfc0710c, 32'h3f72b120} /* (4, 11, 8) {real, imag} */,
  {32'hbf6db495, 32'hbf33a646} /* (4, 11, 7) {real, imag} */,
  {32'hbf35661e, 32'hc006d69f} /* (4, 11, 6) {real, imag} */,
  {32'hc08dadab, 32'hbfc8faf0} /* (4, 11, 5) {real, imag} */,
  {32'hbde7de12, 32'h3f3621ee} /* (4, 11, 4) {real, imag} */,
  {32'h407219de, 32'h3ed2fdb1} /* (4, 11, 3) {real, imag} */,
  {32'h3f2a8bae, 32'hc090e89b} /* (4, 11, 2) {real, imag} */,
  {32'h40c4f597, 32'hbee0def7} /* (4, 11, 1) {real, imag} */,
  {32'h3fe3816e, 32'hbf50b365} /* (4, 11, 0) {real, imag} */,
  {32'hc0005cad, 32'hc00627b2} /* (4, 10, 31) {real, imag} */,
  {32'h3fda92f9, 32'h408d9ae1} /* (4, 10, 30) {real, imag} */,
  {32'h4017d97b, 32'hbf366b18} /* (4, 10, 29) {real, imag} */,
  {32'hbf0c2bb8, 32'h3e4bb2cf} /* (4, 10, 28) {real, imag} */,
  {32'hbf91f6f5, 32'h3f578439} /* (4, 10, 27) {real, imag} */,
  {32'hc052101f, 32'h402ee1d2} /* (4, 10, 26) {real, imag} */,
  {32'hbfef55d0, 32'h4011a2fc} /* (4, 10, 25) {real, imag} */,
  {32'h3f3b9b4c, 32'hbdd93fbe} /* (4, 10, 24) {real, imag} */,
  {32'h3fc1f4fb, 32'hc0b84927} /* (4, 10, 23) {real, imag} */,
  {32'hbed04182, 32'hbe512868} /* (4, 10, 22) {real, imag} */,
  {32'h40269995, 32'hbfc1863e} /* (4, 10, 21) {real, imag} */,
  {32'h3f872626, 32'h40009178} /* (4, 10, 20) {real, imag} */,
  {32'h3eb80f8e, 32'h3f5ce9e6} /* (4, 10, 19) {real, imag} */,
  {32'hbe73be23, 32'h3f96c78f} /* (4, 10, 18) {real, imag} */,
  {32'h3f1eb52e, 32'h3d2296a3} /* (4, 10, 17) {real, imag} */,
  {32'hbf3c4ba9, 32'hbf90d99b} /* (4, 10, 16) {real, imag} */,
  {32'hc03c24fd, 32'h3e6f738d} /* (4, 10, 15) {real, imag} */,
  {32'hbf6e0ee6, 32'hbff4cbc4} /* (4, 10, 14) {real, imag} */,
  {32'hbe47f782, 32'h3fa482a1} /* (4, 10, 13) {real, imag} */,
  {32'hc0130e31, 32'h3fc8d618} /* (4, 10, 12) {real, imag} */,
  {32'hbfbcb373, 32'h3f073de9} /* (4, 10, 11) {real, imag} */,
  {32'hbf963542, 32'hbd4d6542} /* (4, 10, 10) {real, imag} */,
  {32'h40909e3e, 32'hc01a416b} /* (4, 10, 9) {real, imag} */,
  {32'h4049b0f1, 32'hc04f4612} /* (4, 10, 8) {real, imag} */,
  {32'hc008f060, 32'hbed97695} /* (4, 10, 7) {real, imag} */,
  {32'hbfdcf3c7, 32'h400e56f2} /* (4, 10, 6) {real, imag} */,
  {32'h3fce53e6, 32'h3fcaffed} /* (4, 10, 5) {real, imag} */,
  {32'h3fd4ca0a, 32'hc0243aae} /* (4, 10, 4) {real, imag} */,
  {32'h40327463, 32'hbfe43631} /* (4, 10, 3) {real, imag} */,
  {32'h409cbc3d, 32'h3ea44f25} /* (4, 10, 2) {real, imag} */,
  {32'h3ea86129, 32'h3e38cfc1} /* (4, 10, 1) {real, imag} */,
  {32'hc054d540, 32'hbe371ff7} /* (4, 10, 0) {real, imag} */,
  {32'h3f94f384, 32'hc01fe32c} /* (4, 9, 31) {real, imag} */,
  {32'h40166f44, 32'h4023ce49} /* (4, 9, 30) {real, imag} */,
  {32'h3ed68390, 32'hbfc4b25e} /* (4, 9, 29) {real, imag} */,
  {32'hc0cac31e, 32'h40447286} /* (4, 9, 28) {real, imag} */,
  {32'h3ffe6500, 32'hbfd562d7} /* (4, 9, 27) {real, imag} */,
  {32'hbf2fcd1f, 32'hbe9750b0} /* (4, 9, 26) {real, imag} */,
  {32'h3ff1a975, 32'hbfcf9a28} /* (4, 9, 25) {real, imag} */,
  {32'h401775cd, 32'hbf3b3853} /* (4, 9, 24) {real, imag} */,
  {32'h3ff3c38a, 32'h3dbb7700} /* (4, 9, 23) {real, imag} */,
  {32'hbf1c5928, 32'h3fbe1b9e} /* (4, 9, 22) {real, imag} */,
  {32'h40616539, 32'h3ee6d828} /* (4, 9, 21) {real, imag} */,
  {32'hbd971eb5, 32'h3ed9bfc1} /* (4, 9, 20) {real, imag} */,
  {32'hbf2a1f84, 32'hbf223627} /* (4, 9, 19) {real, imag} */,
  {32'hbeb4a93e, 32'hbf530304} /* (4, 9, 18) {real, imag} */,
  {32'h3f184cf4, 32'hbfb4b63d} /* (4, 9, 17) {real, imag} */,
  {32'h3f8eed85, 32'hbf26cba1} /* (4, 9, 16) {real, imag} */,
  {32'h3fa69a84, 32'h3e7fda12} /* (4, 9, 15) {real, imag} */,
  {32'hbf7fff97, 32'hbf862180} /* (4, 9, 14) {real, imag} */,
  {32'h3fc2f901, 32'h3f8748f0} /* (4, 9, 13) {real, imag} */,
  {32'h3f6b93c6, 32'h402148d5} /* (4, 9, 12) {real, imag} */,
  {32'h3f09735b, 32'h3f80f578} /* (4, 9, 11) {real, imag} */,
  {32'h401d0f85, 32'h3f7ec0bc} /* (4, 9, 10) {real, imag} */,
  {32'hbf8ecb38, 32'h3fc6d569} /* (4, 9, 9) {real, imag} */,
  {32'hc07c17be, 32'h403aab6b} /* (4, 9, 8) {real, imag} */,
  {32'hbe887da2, 32'h40528a84} /* (4, 9, 7) {real, imag} */,
  {32'h40b7a914, 32'hc08475b6} /* (4, 9, 6) {real, imag} */,
  {32'hbf3f8367, 32'h3f5da665} /* (4, 9, 5) {real, imag} */,
  {32'hbfa59298, 32'h400a7a3b} /* (4, 9, 4) {real, imag} */,
  {32'hc087a579, 32'h3ff3817a} /* (4, 9, 3) {real, imag} */,
  {32'h400f13c1, 32'hbfa468f9} /* (4, 9, 2) {real, imag} */,
  {32'hc0c542a9, 32'hbf942ea8} /* (4, 9, 1) {real, imag} */,
  {32'hbfdf855f, 32'hc0029399} /* (4, 9, 0) {real, imag} */,
  {32'h40f9bfbb, 32'hc0e9cc1c} /* (4, 8, 31) {real, imag} */,
  {32'hc04fdc1b, 32'h4093aa16} /* (4, 8, 30) {real, imag} */,
  {32'hc084bf9e, 32'h40c966e2} /* (4, 8, 29) {real, imag} */,
  {32'h4083a5cf, 32'hc01cd06c} /* (4, 8, 28) {real, imag} */,
  {32'h40490168, 32'h4094a619} /* (4, 8, 27) {real, imag} */,
  {32'h3ea194b5, 32'h4013ad3a} /* (4, 8, 26) {real, imag} */,
  {32'h40375430, 32'hc03d33ad} /* (4, 8, 25) {real, imag} */,
  {32'h4002310a, 32'h3e753c80} /* (4, 8, 24) {real, imag} */,
  {32'h402a56b7, 32'h400bf837} /* (4, 8, 23) {real, imag} */,
  {32'h3f9c2a37, 32'hbfad1e9d} /* (4, 8, 22) {real, imag} */,
  {32'hc03d1744, 32'h4050333e} /* (4, 8, 21) {real, imag} */,
  {32'hbe1c7c19, 32'h3ff19bb2} /* (4, 8, 20) {real, imag} */,
  {32'hbfe04118, 32'h3f60cebe} /* (4, 8, 19) {real, imag} */,
  {32'hbf845fe0, 32'hbd4f1088} /* (4, 8, 18) {real, imag} */,
  {32'hbd695a67, 32'h3e10608d} /* (4, 8, 17) {real, imag} */,
  {32'hbe84735b, 32'hbff4517c} /* (4, 8, 16) {real, imag} */,
  {32'h40088128, 32'hbe79a066} /* (4, 8, 15) {real, imag} */,
  {32'h4036db56, 32'hbf7a0b2c} /* (4, 8, 14) {real, imag} */,
  {32'hc00d94f4, 32'h3f538ab9} /* (4, 8, 13) {real, imag} */,
  {32'hc001f06b, 32'hc0747d13} /* (4, 8, 12) {real, imag} */,
  {32'hbf918368, 32'h3f8c270f} /* (4, 8, 11) {real, imag} */,
  {32'hbfde9834, 32'h3efc46e9} /* (4, 8, 10) {real, imag} */,
  {32'h3fd5fefe, 32'hbefaaeb8} /* (4, 8, 9) {real, imag} */,
  {32'hbf118345, 32'hbdb97a45} /* (4, 8, 8) {real, imag} */,
  {32'h407bfadd, 32'h40560785} /* (4, 8, 7) {real, imag} */,
  {32'hc0668c5a, 32'hbfab1618} /* (4, 8, 6) {real, imag} */,
  {32'hc00db859, 32'hc0ce739c} /* (4, 8, 5) {real, imag} */,
  {32'h40901f6d, 32'h3fbfcfd5} /* (4, 8, 4) {real, imag} */,
  {32'hbf5d449a, 32'h3f7b6921} /* (4, 8, 3) {real, imag} */,
  {32'hc07eff2f, 32'h40b830a9} /* (4, 8, 2) {real, imag} */,
  {32'h4132a3a2, 32'hc06ef32a} /* (4, 8, 1) {real, imag} */,
  {32'h40024a59, 32'hbf877adf} /* (4, 8, 0) {real, imag} */,
  {32'h3f90a002, 32'h40a49773} /* (4, 7, 31) {real, imag} */,
  {32'h401228c5, 32'hc080f5ec} /* (4, 7, 30) {real, imag} */,
  {32'hc0179b29, 32'h403000ad} /* (4, 7, 29) {real, imag} */,
  {32'h400203f5, 32'h403bd5d9} /* (4, 7, 28) {real, imag} */,
  {32'hbf2c604b, 32'hc0c52dcc} /* (4, 7, 27) {real, imag} */,
  {32'hc02ec76e, 32'hbfa9fb9b} /* (4, 7, 26) {real, imag} */,
  {32'hc011806b, 32'hc0268217} /* (4, 7, 25) {real, imag} */,
  {32'hbed279eb, 32'hbf7ecc48} /* (4, 7, 24) {real, imag} */,
  {32'h406ea534, 32'h40165a6d} /* (4, 7, 23) {real, imag} */,
  {32'hbefbcde7, 32'hbea8b1b9} /* (4, 7, 22) {real, imag} */,
  {32'hbed3432b, 32'hbebbb186} /* (4, 7, 21) {real, imag} */,
  {32'h40068999, 32'h4007e3f5} /* (4, 7, 20) {real, imag} */,
  {32'hbede77dd, 32'hc06392e0} /* (4, 7, 19) {real, imag} */,
  {32'hbfaa8fc9, 32'h3d3e15a9} /* (4, 7, 18) {real, imag} */,
  {32'h3fbdd93d, 32'hbf626fad} /* (4, 7, 17) {real, imag} */,
  {32'h3ff9ade5, 32'hbf8e4a98} /* (4, 7, 16) {real, imag} */,
  {32'hbf9531ad, 32'hbf939686} /* (4, 7, 15) {real, imag} */,
  {32'h400d307c, 32'h3fce0ddd} /* (4, 7, 14) {real, imag} */,
  {32'h3fca2df4, 32'hbd45506f} /* (4, 7, 13) {real, imag} */,
  {32'hbf4bccf6, 32'hbf8eea51} /* (4, 7, 12) {real, imag} */,
  {32'h400bfb3c, 32'hc010a173} /* (4, 7, 11) {real, imag} */,
  {32'hc06ce5d0, 32'h40369534} /* (4, 7, 10) {real, imag} */,
  {32'h3fa7ce63, 32'hbf034421} /* (4, 7, 9) {real, imag} */,
  {32'hbdbe2c17, 32'h3fec7ae2} /* (4, 7, 8) {real, imag} */,
  {32'h40a2e4f3, 32'hc00a6e7e} /* (4, 7, 7) {real, imag} */,
  {32'hc0a87f67, 32'h401df0d8} /* (4, 7, 6) {real, imag} */,
  {32'hbfbf5d6f, 32'h409e6d43} /* (4, 7, 5) {real, imag} */,
  {32'hbf0e68e3, 32'hc0204f41} /* (4, 7, 4) {real, imag} */,
  {32'hc0313c59, 32'hbfe8d68c} /* (4, 7, 3) {real, imag} */,
  {32'h40b1c70e, 32'h3e9990e9} /* (4, 7, 2) {real, imag} */,
  {32'hc10b524d, 32'hbf61f465} /* (4, 7, 1) {real, imag} */,
  {32'hc037cb8f, 32'h405ad442} /* (4, 7, 0) {real, imag} */,
  {32'hc0872809, 32'h3daf95a4} /* (4, 6, 31) {real, imag} */,
  {32'hc0c505f6, 32'h4065ac28} /* (4, 6, 30) {real, imag} */,
  {32'hbf113567, 32'hc00b1602} /* (4, 6, 29) {real, imag} */,
  {32'hc016d383, 32'h4043559b} /* (4, 6, 28) {real, imag} */,
  {32'hc03b7bd0, 32'hbf28cafd} /* (4, 6, 27) {real, imag} */,
  {32'hbffadc81, 32'h3fc5a99d} /* (4, 6, 26) {real, imag} */,
  {32'hbe940f9d, 32'h40302897} /* (4, 6, 25) {real, imag} */,
  {32'h406dfb40, 32'hbf987903} /* (4, 6, 24) {real, imag} */,
  {32'h4039ed8b, 32'hbf1d8bab} /* (4, 6, 23) {real, imag} */,
  {32'hbfb15884, 32'hc08e39b6} /* (4, 6, 22) {real, imag} */,
  {32'h401a7ff6, 32'hbfd43620} /* (4, 6, 21) {real, imag} */,
  {32'h3e171f0d, 32'hc0972812} /* (4, 6, 20) {real, imag} */,
  {32'h3f84dab4, 32'hbfcf3d8b} /* (4, 6, 19) {real, imag} */,
  {32'h3f2a8b39, 32'h3e67a37a} /* (4, 6, 18) {real, imag} */,
  {32'h3f9da833, 32'h3eca6984} /* (4, 6, 17) {real, imag} */,
  {32'h3f0038f6, 32'h3cc65452} /* (4, 6, 16) {real, imag} */,
  {32'h3c8c41c0, 32'h3f7b5302} /* (4, 6, 15) {real, imag} */,
  {32'hbfa47b83, 32'h3f77401b} /* (4, 6, 14) {real, imag} */,
  {32'hbf20c614, 32'hbfdadb42} /* (4, 6, 13) {real, imag} */,
  {32'hbfc2014f, 32'h3ffff70a} /* (4, 6, 12) {real, imag} */,
  {32'hc0194e3e, 32'hbf5dcfd7} /* (4, 6, 11) {real, imag} */,
  {32'hbf1d800e, 32'h4005c35c} /* (4, 6, 10) {real, imag} */,
  {32'h402138d3, 32'hbfbe7e35} /* (4, 6, 9) {real, imag} */,
  {32'h3f9ab373, 32'h3ff48743} /* (4, 6, 8) {real, imag} */,
  {32'hbd7878f6, 32'hbfd2741a} /* (4, 6, 7) {real, imag} */,
  {32'hbe4a8a10, 32'hc07b7110} /* (4, 6, 6) {real, imag} */,
  {32'h3fe89a5d, 32'h3fba08ac} /* (4, 6, 5) {real, imag} */,
  {32'h3fe13c31, 32'hbf01e0f1} /* (4, 6, 4) {real, imag} */,
  {32'h3ebd04bb, 32'h3fd1c5e1} /* (4, 6, 3) {real, imag} */,
  {32'hc0584f04, 32'hc09755f6} /* (4, 6, 2) {real, imag} */,
  {32'hbf870635, 32'hc03be1cd} /* (4, 6, 1) {real, imag} */,
  {32'hc00e91e8, 32'hc09b6666} /* (4, 6, 0) {real, imag} */,
  {32'h4016f3b3, 32'hc10013c3} /* (4, 5, 31) {real, imag} */,
  {32'hbef3f08f, 32'h402a723c} /* (4, 5, 30) {real, imag} */,
  {32'h401b2a21, 32'hbf2e7c37} /* (4, 5, 29) {real, imag} */,
  {32'h40be5549, 32'hc01f5275} /* (4, 5, 28) {real, imag} */,
  {32'hc002ad9a, 32'h4098a706} /* (4, 5, 27) {real, imag} */,
  {32'hbf01d6e2, 32'hbe0bbbdf} /* (4, 5, 26) {real, imag} */,
  {32'hc073f349, 32'hc08d0571} /* (4, 5, 25) {real, imag} */,
  {32'hbf767709, 32'hbfed0b80} /* (4, 5, 24) {real, imag} */,
  {32'h3fd4f557, 32'hbf81a135} /* (4, 5, 23) {real, imag} */,
  {32'hbf18d197, 32'hbf2528de} /* (4, 5, 22) {real, imag} */,
  {32'hbf91d970, 32'h4011ef71} /* (4, 5, 21) {real, imag} */,
  {32'h3dc9a26b, 32'hc01e3010} /* (4, 5, 20) {real, imag} */,
  {32'h4087d218, 32'hbf573a3a} /* (4, 5, 19) {real, imag} */,
  {32'h3f6a543c, 32'h3fa86e68} /* (4, 5, 18) {real, imag} */,
  {32'hbf2c3805, 32'h3c955d1e} /* (4, 5, 17) {real, imag} */,
  {32'h3f687a3d, 32'hbecc82c3} /* (4, 5, 16) {real, imag} */,
  {32'h3edd8c4d, 32'hbe65d09a} /* (4, 5, 15) {real, imag} */,
  {32'h3f0bcf74, 32'hbeaf5479} /* (4, 5, 14) {real, imag} */,
  {32'h3ff2028b, 32'hbe8f6aab} /* (4, 5, 13) {real, imag} */,
  {32'h3e98f05f, 32'h3e6faaf9} /* (4, 5, 12) {real, imag} */,
  {32'hbfc93fe1, 32'h3f059275} /* (4, 5, 11) {real, imag} */,
  {32'h3ee65f48, 32'hc08a34b3} /* (4, 5, 10) {real, imag} */,
  {32'hc031be0e, 32'hbe931244} /* (4, 5, 9) {real, imag} */,
  {32'h3f241ad8, 32'hc03a7b93} /* (4, 5, 8) {real, imag} */,
  {32'h3fb1c5f8, 32'hbe9a601d} /* (4, 5, 7) {real, imag} */,
  {32'hbfc3a1d2, 32'h40f18960} /* (4, 5, 6) {real, imag} */,
  {32'h3cd622be, 32'h3f396928} /* (4, 5, 5) {real, imag} */,
  {32'hc039dd74, 32'h3fae8f0b} /* (4, 5, 4) {real, imag} */,
  {32'hc0746d4c, 32'h3f59642e} /* (4, 5, 3) {real, imag} */,
  {32'hc094879a, 32'h408c62be} /* (4, 5, 2) {real, imag} */,
  {32'h41425323, 32'hc0b0aa2b} /* (4, 5, 1) {real, imag} */,
  {32'h40dde50e, 32'hc0c1c34a} /* (4, 5, 0) {real, imag} */,
  {32'hc174f041, 32'h412dee90} /* (4, 4, 31) {real, imag} */,
  {32'h414abae3, 32'h40369d72} /* (4, 4, 30) {real, imag} */,
  {32'hc04cbbe0, 32'hc0a030b9} /* (4, 4, 29) {real, imag} */,
  {32'hc1474531, 32'h40e2b654} /* (4, 4, 28) {real, imag} */,
  {32'hbe838c20, 32'hc0a0ff43} /* (4, 4, 27) {real, imag} */,
  {32'h4022a9ca, 32'h40301058} /* (4, 4, 26) {real, imag} */,
  {32'hc07aa49a, 32'hbe1775a2} /* (4, 4, 25) {real, imag} */,
  {32'hbf686f11, 32'hbf8aa181} /* (4, 4, 24) {real, imag} */,
  {32'h4063e850, 32'hbfdb589a} /* (4, 4, 23) {real, imag} */,
  {32'hbf93486b, 32'h3f8f6941} /* (4, 4, 22) {real, imag} */,
  {32'h3fce843c, 32'hc003daa3} /* (4, 4, 21) {real, imag} */,
  {32'h3acd0892, 32'h3f59c098} /* (4, 4, 20) {real, imag} */,
  {32'hbfc89136, 32'h403a7128} /* (4, 4, 19) {real, imag} */,
  {32'hbefddd7d, 32'h3f38e123} /* (4, 4, 18) {real, imag} */,
  {32'hbf94d277, 32'hbeadb9c8} /* (4, 4, 17) {real, imag} */,
  {32'h3ee2f0bd, 32'hbefb5d21} /* (4, 4, 16) {real, imag} */,
  {32'h3f15d200, 32'hbd099f7a} /* (4, 4, 15) {real, imag} */,
  {32'h3f4d997b, 32'hbf7aa0a6} /* (4, 4, 14) {real, imag} */,
  {32'h406ce146, 32'h3f73d46b} /* (4, 4, 13) {real, imag} */,
  {32'hbf0fa309, 32'hbefc582a} /* (4, 4, 12) {real, imag} */,
  {32'h3ff49769, 32'h3f285f7b} /* (4, 4, 11) {real, imag} */,
  {32'h3f47164e, 32'hbfceeec5} /* (4, 4, 10) {real, imag} */,
  {32'h404ad63d, 32'h403cc251} /* (4, 4, 9) {real, imag} */,
  {32'h40122a80, 32'hbdf0d213} /* (4, 4, 8) {real, imag} */,
  {32'hc044de01, 32'h3f873b32} /* (4, 4, 7) {real, imag} */,
  {32'h40493917, 32'hc069414b} /* (4, 4, 6) {real, imag} */,
  {32'h3df37b9b, 32'hbf3abe2d} /* (4, 4, 5) {real, imag} */,
  {32'hc08b4c23, 32'hbf9bcfa0} /* (4, 4, 4) {real, imag} */,
  {32'hc0213521, 32'h409431cd} /* (4, 4, 3) {real, imag} */,
  {32'h41708f1e, 32'hc082c799} /* (4, 4, 2) {real, imag} */,
  {32'hc17f0f95, 32'h41c55b5a} /* (4, 4, 1) {real, imag} */,
  {32'hc0db90c1, 32'h4062319f} /* (4, 4, 0) {real, imag} */,
  {32'h3fdc962d, 32'hc195b01c} /* (4, 3, 31) {real, imag} */,
  {32'h415dd7c4, 32'h41242df6} /* (4, 3, 30) {real, imag} */,
  {32'h3fec68c3, 32'h40a2d561} /* (4, 3, 29) {real, imag} */,
  {32'hc036eac3, 32'hc054920d} /* (4, 3, 28) {real, imag} */,
  {32'h402fe671, 32'h408da99c} /* (4, 3, 27) {real, imag} */,
  {32'h3d5a7b3c, 32'hbfbb473b} /* (4, 3, 26) {real, imag} */,
  {32'h3ffa16f1, 32'hc005e67a} /* (4, 3, 25) {real, imag} */,
  {32'h3f4781fc, 32'h3fca1226} /* (4, 3, 24) {real, imag} */,
  {32'hc08cd733, 32'h3e8523d7} /* (4, 3, 23) {real, imag} */,
  {32'hbf87a913, 32'h400b4825} /* (4, 3, 22) {real, imag} */,
  {32'h3fbd8b15, 32'hc064362b} /* (4, 3, 21) {real, imag} */,
  {32'hc06e3c89, 32'h4006bace} /* (4, 3, 20) {real, imag} */,
  {32'h40022d2b, 32'h3f6e8a9c} /* (4, 3, 19) {real, imag} */,
  {32'h3fb702e4, 32'h3fc5adf0} /* (4, 3, 18) {real, imag} */,
  {32'hbfd16e68, 32'hc03001d0} /* (4, 3, 17) {real, imag} */,
  {32'hbe8c67a4, 32'h40009711} /* (4, 3, 16) {real, imag} */,
  {32'hbed0a859, 32'h3ea95d13} /* (4, 3, 15) {real, imag} */,
  {32'hbf138d5c, 32'h3fc152f7} /* (4, 3, 14) {real, imag} */,
  {32'hc02418d1, 32'h3f262597} /* (4, 3, 13) {real, imag} */,
  {32'h3dc3bf9c, 32'hc020503d} /* (4, 3, 12) {real, imag} */,
  {32'h3e015fbf, 32'h3fda031e} /* (4, 3, 11) {real, imag} */,
  {32'hbf6e16c2, 32'hc04c1b17} /* (4, 3, 10) {real, imag} */,
  {32'h3fe227be, 32'hc0051c41} /* (4, 3, 9) {real, imag} */,
  {32'h3e835fa0, 32'hbe929c85} /* (4, 3, 8) {real, imag} */,
  {32'hc0b1e5a5, 32'h40a86f08} /* (4, 3, 7) {real, imag} */,
  {32'h3f929d97, 32'h40b067e5} /* (4, 3, 6) {real, imag} */,
  {32'h3fe0ef12, 32'h407193af} /* (4, 3, 5) {real, imag} */,
  {32'h4028bb93, 32'hbf06a61d} /* (4, 3, 4) {real, imag} */,
  {32'hc0e2339b, 32'h3e63cc90} /* (4, 3, 3) {real, imag} */,
  {32'h410ff4b0, 32'hbf99ecb4} /* (4, 3, 2) {real, imag} */,
  {32'hc17761d3, 32'hbfb4b744} /* (4, 3, 1) {real, imag} */,
  {32'h3fe52126, 32'hbf8d7d16} /* (4, 3, 0) {real, imag} */,
  {32'h4202aeb2, 32'hc295499b} /* (4, 2, 31) {real, imag} */,
  {32'hc13c128f, 32'h42468722} /* (4, 2, 30) {real, imag} */,
  {32'h40618cda, 32'hc1168dc2} /* (4, 2, 29) {real, imag} */,
  {32'hc08cb6ee, 32'hc1529b05} /* (4, 2, 28) {real, imag} */,
  {32'h404ea0ce, 32'h41065381} /* (4, 2, 27) {real, imag} */,
  {32'hc02c7ab4, 32'hc034fd57} /* (4, 2, 26) {real, imag} */,
  {32'h3f43795b, 32'hc00b0930} /* (4, 2, 25) {real, imag} */,
  {32'h3fdc27e3, 32'h40fc2d8d} /* (4, 2, 24) {real, imag} */,
  {32'h400a6410, 32'h3f82cc7e} /* (4, 2, 23) {real, imag} */,
  {32'hc08d7904, 32'h3f3de555} /* (4, 2, 22) {real, imag} */,
  {32'h40658017, 32'h403530f2} /* (4, 2, 21) {real, imag} */,
  {32'hbfc33504, 32'hbf8c2fa4} /* (4, 2, 20) {real, imag} */,
  {32'h3e47920c, 32'h3ea5855f} /* (4, 2, 19) {real, imag} */,
  {32'h3f2910be, 32'hbe89bcd4} /* (4, 2, 18) {real, imag} */,
  {32'hbea6b8e9, 32'hb9dc551e} /* (4, 2, 17) {real, imag} */,
  {32'hbfc8505e, 32'h3f8b2399} /* (4, 2, 16) {real, imag} */,
  {32'hbf7fa5d2, 32'hbf826fab} /* (4, 2, 15) {real, imag} */,
  {32'hbff52692, 32'h40379659} /* (4, 2, 14) {real, imag} */,
  {32'h3ed39cea, 32'hbf75867f} /* (4, 2, 13) {real, imag} */,
  {32'h3e6f6f84, 32'hc00a52ec} /* (4, 2, 12) {real, imag} */,
  {32'hc0310ebe, 32'h3e58f34c} /* (4, 2, 11) {real, imag} */,
  {32'h3d0dd17a, 32'hc00a8a19} /* (4, 2, 10) {real, imag} */,
  {32'hc03f6dea, 32'h3f6339b5} /* (4, 2, 9) {real, imag} */,
  {32'hc056644a, 32'h40c53aa0} /* (4, 2, 8) {real, imag} */,
  {32'h4056e43c, 32'hbf1b3850} /* (4, 2, 7) {real, imag} */,
  {32'hc0321fd8, 32'hbf8f70a1} /* (4, 2, 6) {real, imag} */,
  {32'hc0f3c0ef, 32'h410248da} /* (4, 2, 5) {real, imag} */,
  {32'hbff383fd, 32'hc117c94b} /* (4, 2, 4) {real, imag} */,
  {32'h404847a9, 32'hc0ced8c3} /* (4, 2, 3) {real, imag} */,
  {32'hbed63da6, 32'h42090cdb} /* (4, 2, 2) {real, imag} */,
  {32'h40f21c1a, 32'hc22f8b17} /* (4, 2, 1) {real, imag} */,
  {32'h41b0c404, 32'hc21e4bbc} /* (4, 2, 0) {real, imag} */,
  {32'hc0391f02, 32'h42848756} /* (4, 1, 31) {real, imag} */,
  {32'h413ecfd2, 32'hc1e14199} /* (4, 1, 30) {real, imag} */,
  {32'hbf616836, 32'h40f36c88} /* (4, 1, 29) {real, imag} */,
  {32'hc033a82e, 32'h414c6779} /* (4, 1, 28) {real, imag} */,
  {32'h40f7fd93, 32'hc19d40e3} /* (4, 1, 27) {real, imag} */,
  {32'hc08b297c, 32'h404fa4d0} /* (4, 1, 26) {real, imag} */,
  {32'h4098dac9, 32'h3f511f23} /* (4, 1, 25) {real, imag} */,
  {32'hc04b0976, 32'hc0d8bdd4} /* (4, 1, 24) {real, imag} */,
  {32'h3e9aa20a, 32'h3ef528e8} /* (4, 1, 23) {real, imag} */,
  {32'h3f0a3475, 32'h3fd88f48} /* (4, 1, 22) {real, imag} */,
  {32'hc10e6297, 32'hc0b68869} /* (4, 1, 21) {real, imag} */,
  {32'h40939630, 32'h3faca6e8} /* (4, 1, 20) {real, imag} */,
  {32'hbfcf6a6a, 32'h3f2647fc} /* (4, 1, 19) {real, imag} */,
  {32'hc064db7c, 32'h3e8ab14c} /* (4, 1, 18) {real, imag} */,
  {32'hbf3b3760, 32'hbeb46be6} /* (4, 1, 17) {real, imag} */,
  {32'h3ff1b942, 32'h3f59a416} /* (4, 1, 16) {real, imag} */,
  {32'hbfe7244e, 32'hbfcfdb2c} /* (4, 1, 15) {real, imag} */,
  {32'h3e6d7d40, 32'h3fbc7029} /* (4, 1, 14) {real, imag} */,
  {32'hbf4f52d2, 32'hbf112b16} /* (4, 1, 13) {real, imag} */,
  {32'hbd4c28e7, 32'hc022a943} /* (4, 1, 12) {real, imag} */,
  {32'h402b2cad, 32'hbf4b5145} /* (4, 1, 11) {real, imag} */,
  {32'hbfde5996, 32'hc00a8812} /* (4, 1, 10) {real, imag} */,
  {32'h40147b07, 32'h403d9252} /* (4, 1, 9) {real, imag} */,
  {32'h40d90411, 32'hbea579ca} /* (4, 1, 8) {real, imag} */,
  {32'hbf6cce40, 32'hbe876091} /* (4, 1, 7) {real, imag} */,
  {32'h409c706f, 32'h4044e51c} /* (4, 1, 6) {real, imag} */,
  {32'h413448a3, 32'hc0e0e8ab} /* (4, 1, 5) {real, imag} */,
  {32'hc0012445, 32'hbf3de2c2} /* (4, 1, 4) {real, imag} */,
  {32'hc009aebc, 32'hc12060b2} /* (4, 1, 3) {real, imag} */,
  {32'h4273320d, 32'hc17c37e8} /* (4, 1, 2) {real, imag} */,
  {32'hc2a2aa6d, 32'h42805593} /* (4, 1, 1) {real, imag} */,
  {32'hc242fdcf, 32'h42655ace} /* (4, 1, 0) {real, imag} */,
  {32'h419928ba, 32'h42766e9a} /* (4, 0, 31) {real, imag} */,
  {32'hc18101bc, 32'hc04ddff0} /* (4, 0, 30) {real, imag} */,
  {32'h3f91e829, 32'h40b50e8f} /* (4, 0, 29) {real, imag} */,
  {32'hc0475a4e, 32'hc0a7bf94} /* (4, 0, 28) {real, imag} */,
  {32'h40ecbeb1, 32'hc1014cc7} /* (4, 0, 27) {real, imag} */,
  {32'h405a41ca, 32'h3d32855c} /* (4, 0, 26) {real, imag} */,
  {32'h40a9dbd3, 32'h404be6d4} /* (4, 0, 25) {real, imag} */,
  {32'hbfe685ad, 32'hc03bcf93} /* (4, 0, 24) {real, imag} */,
  {32'hc09478e6, 32'hc0be9dcc} /* (4, 0, 23) {real, imag} */,
  {32'h4042ef8d, 32'hbf6b0428} /* (4, 0, 22) {real, imag} */,
  {32'h3f0467b7, 32'hc0978442} /* (4, 0, 21) {real, imag} */,
  {32'h3f550d7c, 32'hbe4384fe} /* (4, 0, 20) {real, imag} */,
  {32'hbe99f321, 32'h3e4554b0} /* (4, 0, 19) {real, imag} */,
  {32'hc084a11f, 32'hbf923215} /* (4, 0, 18) {real, imag} */,
  {32'hbfcd545c, 32'h3f2c61e7} /* (4, 0, 17) {real, imag} */,
  {32'h3f99023b, 32'hbef26135} /* (4, 0, 16) {real, imag} */,
  {32'h3f5f462e, 32'hbef13711} /* (4, 0, 15) {real, imag} */,
  {32'h3fd3de62, 32'hbee5505b} /* (4, 0, 14) {real, imag} */,
  {32'hbea3a473, 32'hc03d9d20} /* (4, 0, 13) {real, imag} */,
  {32'hbe2ade7a, 32'hbee71309} /* (4, 0, 12) {real, imag} */,
  {32'h40190d63, 32'hbfb221e0} /* (4, 0, 11) {real, imag} */,
  {32'hba70eff8, 32'hc072353f} /* (4, 0, 10) {real, imag} */,
  {32'h40a0f3b0, 32'h40311608} /* (4, 0, 9) {real, imag} */,
  {32'h4087034b, 32'hbf1312f6} /* (4, 0, 8) {real, imag} */,
  {32'hc0a99bc5, 32'hbfd59e07} /* (4, 0, 7) {real, imag} */,
  {32'hbfcfaba1, 32'hc04bc282} /* (4, 0, 6) {real, imag} */,
  {32'h3efd30e6, 32'hc0d831b1} /* (4, 0, 5) {real, imag} */,
  {32'h4047d27e, 32'h40905c56} /* (4, 0, 4) {real, imag} */,
  {32'h40967372, 32'hc11ba78e} /* (4, 0, 3) {real, imag} */,
  {32'h418b47f7, 32'h3fdbe539} /* (4, 0, 2) {real, imag} */,
  {32'hc25be04b, 32'h4202f6bb} /* (4, 0, 1) {real, imag} */,
  {32'hc1c0d8dc, 32'h42292b7d} /* (4, 0, 0) {real, imag} */,
  {32'h41ffaae4, 32'h4339b71d} /* (3, 31, 31) {real, imag} */,
  {32'hc21431e3, 32'hc2934ac6} /* (3, 31, 30) {real, imag} */,
  {32'h41946661, 32'hc1927a72} /* (3, 31, 29) {real, imag} */,
  {32'hc090f8dd, 32'h416d854f} /* (3, 31, 28) {real, imag} */,
  {32'hc10fb5df, 32'hc18ea5a3} /* (3, 31, 27) {real, imag} */,
  {32'h40484aee, 32'hc0844f2f} /* (3, 31, 26) {real, imag} */,
  {32'h3ff0c035, 32'h405f6f85} /* (3, 31, 25) {real, imag} */,
  {32'hc0a729fe, 32'h3db36117} /* (3, 31, 24) {real, imag} */,
  {32'h4020d2df, 32'hbf17818a} /* (3, 31, 23) {real, imag} */,
  {32'h3ee34bf7, 32'h3d6088e0} /* (3, 31, 22) {real, imag} */,
  {32'hbf872020, 32'hbfbabbee} /* (3, 31, 21) {real, imag} */,
  {32'h3f9648a7, 32'hbf96d530} /* (3, 31, 20) {real, imag} */,
  {32'h3f254958, 32'hbf0f8a12} /* (3, 31, 19) {real, imag} */,
  {32'hc08126ce, 32'hbf74d79c} /* (3, 31, 18) {real, imag} */,
  {32'h3ff6b0f8, 32'hbe2a66f6} /* (3, 31, 17) {real, imag} */,
  {32'h3f07853d, 32'hbfd6b7cb} /* (3, 31, 16) {real, imag} */,
  {32'h3f1630a9, 32'h3f0da003} /* (3, 31, 15) {real, imag} */,
  {32'h406f70d3, 32'hc0025a78} /* (3, 31, 14) {real, imag} */,
  {32'hbf0c5dcf, 32'h3fbd4055} /* (3, 31, 13) {real, imag} */,
  {32'hbef65b42, 32'h3f3cebfd} /* (3, 31, 12) {real, imag} */,
  {32'h409b5841, 32'hc0dc4b6c} /* (3, 31, 11) {real, imag} */,
  {32'h401e0688, 32'hbf957027} /* (3, 31, 10) {real, imag} */,
  {32'h3e370693, 32'h4088d0c7} /* (3, 31, 9) {real, imag} */,
  {32'h40316663, 32'hc07ed12c} /* (3, 31, 8) {real, imag} */,
  {32'hbf92f272, 32'h40f12eed} /* (3, 31, 7) {real, imag} */,
  {32'hbe3b91d1, 32'hc0576db5} /* (3, 31, 6) {real, imag} */,
  {32'h412ee02a, 32'hc155195a} /* (3, 31, 5) {real, imag} */,
  {32'h405ceea8, 32'h413ac18d} /* (3, 31, 4) {real, imag} */,
  {32'hc110ec6c, 32'hc091a928} /* (3, 31, 3) {real, imag} */,
  {32'h4112c960, 32'hc21f2440} /* (3, 31, 2) {real, imag} */,
  {32'hc287da1a, 32'h42a18326} /* (3, 31, 1) {real, imag} */,
  {32'hc187b308, 32'h42f1e859} /* (3, 31, 0) {real, imag} */,
  {32'h41c9b592, 32'hc28a68f0} /* (3, 30, 31) {real, imag} */,
  {32'hc1ecc9da, 32'h4246c764} /* (3, 30, 30) {real, imag} */,
  {32'h407676ce, 32'h408a4197} /* (3, 30, 29) {real, imag} */,
  {32'h400ef944, 32'hc1cc64b1} /* (3, 30, 28) {real, imag} */,
  {32'hc0f5717c, 32'h4116a8c5} /* (3, 30, 27) {real, imag} */,
  {32'hbfbe2f5c, 32'h40578355} /* (3, 30, 26) {real, imag} */,
  {32'hc0b61a4a, 32'hc0806ffc} /* (3, 30, 25) {real, imag} */,
  {32'hc0c72788, 32'h40a376ad} /* (3, 30, 24) {real, imag} */,
  {32'h4058f7ed, 32'h40918067} /* (3, 30, 23) {real, imag} */,
  {32'hbf50ca93, 32'hc03b9e7d} /* (3, 30, 22) {real, imag} */,
  {32'h4015fd27, 32'h407da490} /* (3, 30, 21) {real, imag} */,
  {32'h3ecf1a0f, 32'hbfa54d67} /* (3, 30, 20) {real, imag} */,
  {32'hbf5c8aa6, 32'hbf1a5cb9} /* (3, 30, 19) {real, imag} */,
  {32'h3f843619, 32'hc007737c} /* (3, 30, 18) {real, imag} */,
  {32'h3dc549cb, 32'hbe923cf3} /* (3, 30, 17) {real, imag} */,
  {32'h3d967779, 32'hbaa137b0} /* (3, 30, 16) {real, imag} */,
  {32'hbf3f620b, 32'h4002edbe} /* (3, 30, 15) {real, imag} */,
  {32'hc03b4e11, 32'h3f558f5c} /* (3, 30, 14) {real, imag} */,
  {32'hbf9b560e, 32'h3f045551} /* (3, 30, 13) {real, imag} */,
  {32'hbf48e669, 32'hbf3e4c58} /* (3, 30, 12) {real, imag} */,
  {32'hbfa0103a, 32'hbf0af5da} /* (3, 30, 11) {real, imag} */,
  {32'hbf1db8d3, 32'hbf146883} /* (3, 30, 10) {real, imag} */,
  {32'hbfc83ae4, 32'h3f9dff91} /* (3, 30, 9) {real, imag} */,
  {32'hc058ce96, 32'h40da5840} /* (3, 30, 8) {real, imag} */,
  {32'hbf91f0e0, 32'h4088e116} /* (3, 30, 7) {real, imag} */,
  {32'h40030d2b, 32'h40c94930} /* (3, 30, 6) {real, imag} */,
  {32'hc08e76cd, 32'h40f8e770} /* (3, 30, 5) {real, imag} */,
  {32'h41236e3b, 32'hbf8aa78f} /* (3, 30, 4) {real, imag} */,
  {32'h40d874a9, 32'h3f54f58e} /* (3, 30, 3) {real, imag} */,
  {32'hc2245837, 32'h422f4217} /* (3, 30, 2) {real, imag} */,
  {32'h4194c473, 32'hc2e58a99} /* (3, 30, 1) {real, imag} */,
  {32'hc09bbc3f, 32'hc298f038} /* (3, 30, 0) {real, imag} */,
  {32'h3f2d62c8, 32'h41b9b95b} /* (3, 29, 31) {real, imag} */,
  {32'hc1ebd41e, 32'h3f29d3a3} /* (3, 29, 30) {real, imag} */,
  {32'h4040e80e, 32'h40c09d7a} /* (3, 29, 29) {real, imag} */,
  {32'h40f5b294, 32'hbf84e2cc} /* (3, 29, 28) {real, imag} */,
  {32'hc0c7a80a, 32'h3f8df81d} /* (3, 29, 27) {real, imag} */,
  {32'hbdb91586, 32'hc035e84b} /* (3, 29, 26) {real, imag} */,
  {32'h40a92bba, 32'hbcb01ffc} /* (3, 29, 25) {real, imag} */,
  {32'hc022cca5, 32'hc0908aab} /* (3, 29, 24) {real, imag} */,
  {32'h3f8ae3f0, 32'h4017846f} /* (3, 29, 23) {real, imag} */,
  {32'h3fde6473, 32'hc056cb2f} /* (3, 29, 22) {real, imag} */,
  {32'hbe431877, 32'hbfe62129} /* (3, 29, 21) {real, imag} */,
  {32'h4005a478, 32'hc0694227} /* (3, 29, 20) {real, imag} */,
  {32'hbfd59ab9, 32'hbf6c7aac} /* (3, 29, 19) {real, imag} */,
  {32'hbff9de2e, 32'h3f932d03} /* (3, 29, 18) {real, imag} */,
  {32'h3f52faae, 32'h3f3b20ca} /* (3, 29, 17) {real, imag} */,
  {32'h3f88ed77, 32'hbf7b076b} /* (3, 29, 16) {real, imag} */,
  {32'hbffa7a1c, 32'h3f5ce193} /* (3, 29, 15) {real, imag} */,
  {32'h3f190b0c, 32'h3e465fa9} /* (3, 29, 14) {real, imag} */,
  {32'h3fb1cfbb, 32'hbd24e6c0} /* (3, 29, 13) {real, imag} */,
  {32'hbf9758b0, 32'h3f61e54c} /* (3, 29, 12) {real, imag} */,
  {32'h4035dbf5, 32'hbfe29b29} /* (3, 29, 11) {real, imag} */,
  {32'hc0aabc6e, 32'h3fa031c5} /* (3, 29, 10) {real, imag} */,
  {32'h4028500d, 32'h407ba9a5} /* (3, 29, 9) {real, imag} */,
  {32'hc003d391, 32'hc0702555} /* (3, 29, 8) {real, imag} */,
  {32'h40bce19d, 32'hbed36b08} /* (3, 29, 7) {real, imag} */,
  {32'h3fc79d13, 32'h3f4a3453} /* (3, 29, 6) {real, imag} */,
  {32'hc1006436, 32'hc10f77e1} /* (3, 29, 5) {real, imag} */,
  {32'h3f89ea0f, 32'h409f186d} /* (3, 29, 4) {real, imag} */,
  {32'h3f4f8cb4, 32'h3f69a11a} /* (3, 29, 3) {real, imag} */,
  {32'hc1a5cc30, 32'h40fba628} /* (3, 29, 2) {real, imag} */,
  {32'h415b38a8, 32'hc1d60566} /* (3, 29, 1) {real, imag} */,
  {32'hc05d9b3d, 32'hc0b2ffd9} /* (3, 29, 0) {real, imag} */,
  {32'h414f1384, 32'h41f5161b} /* (3, 28, 31) {real, imag} */,
  {32'hc0fd30dc, 32'hc197ed6d} /* (3, 28, 30) {real, imag} */,
  {32'hc0007116, 32'hc0b68917} /* (3, 28, 29) {real, imag} */,
  {32'h407c800b, 32'h3e1ab0b3} /* (3, 28, 28) {real, imag} */,
  {32'h4080a58e, 32'h40053475} /* (3, 28, 27) {real, imag} */,
  {32'h402f992b, 32'h408da8fa} /* (3, 28, 26) {real, imag} */,
  {32'hbeaab2ff, 32'h40dbef37} /* (3, 28, 25) {real, imag} */,
  {32'hbfe27f1f, 32'h400f6193} /* (3, 28, 24) {real, imag} */,
  {32'hbfaa4fc4, 32'hbfb510a6} /* (3, 28, 23) {real, imag} */,
  {32'hbf2d1e44, 32'hc087b9b3} /* (3, 28, 22) {real, imag} */,
  {32'hc01f68dd, 32'h3f745f9f} /* (3, 28, 21) {real, imag} */,
  {32'hbf103123, 32'hbe511a02} /* (3, 28, 20) {real, imag} */,
  {32'hbf1a3be3, 32'h402275e9} /* (3, 28, 19) {real, imag} */,
  {32'h3fe9f432, 32'hbede3477} /* (3, 28, 18) {real, imag} */,
  {32'h3fb7c8b5, 32'h3ee34892} /* (3, 28, 17) {real, imag} */,
  {32'h3c0576be, 32'hbf76f8bc} /* (3, 28, 16) {real, imag} */,
  {32'hbf15e826, 32'hbf027613} /* (3, 28, 15) {real, imag} */,
  {32'hbf74cb8f, 32'hc03ff773} /* (3, 28, 14) {real, imag} */,
  {32'h3f8f9288, 32'h3f60340f} /* (3, 28, 13) {real, imag} */,
  {32'hbf0ec1c5, 32'h3f996950} /* (3, 28, 12) {real, imag} */,
  {32'hc004e689, 32'hc014e404} /* (3, 28, 11) {real, imag} */,
  {32'hc0157474, 32'h4043f5ce} /* (3, 28, 10) {real, imag} */,
  {32'h402815ff, 32'h402f1676} /* (3, 28, 9) {real, imag} */,
  {32'hbeb0e402, 32'hc0169c1d} /* (3, 28, 8) {real, imag} */,
  {32'h404ddeff, 32'h3ffd5c1d} /* (3, 28, 7) {real, imag} */,
  {32'h40a2ae10, 32'h3ee800ba} /* (3, 28, 6) {real, imag} */,
  {32'hc033fb9b, 32'h3f7602bf} /* (3, 28, 5) {real, imag} */,
  {32'h400593b5, 32'h400b72cf} /* (3, 28, 4) {real, imag} */,
  {32'h3e7d10e7, 32'hbce4c7f9} /* (3, 28, 3) {real, imag} */,
  {32'hc158e69e, 32'hc195de58} /* (3, 28, 2) {real, imag} */,
  {32'h41450b21, 32'h40dd6827} /* (3, 28, 1) {real, imag} */,
  {32'h412b451a, 32'h40aaf819} /* (3, 28, 0) {real, imag} */,
  {32'hc118768c, 32'hc107a8d0} /* (3, 27, 31) {real, imag} */,
  {32'h402ee25d, 32'h40a42b00} /* (3, 27, 30) {real, imag} */,
  {32'hbed3f32b, 32'hc016d08d} /* (3, 27, 29) {real, imag} */,
  {32'hc04e22fb, 32'hc080e270} /* (3, 27, 28) {real, imag} */,
  {32'h410c5983, 32'h407e87c5} /* (3, 27, 27) {real, imag} */,
  {32'hbffcbf33, 32'h3f854e73} /* (3, 27, 26) {real, imag} */,
  {32'h400f4e6f, 32'h40843d78} /* (3, 27, 25) {real, imag} */,
  {32'hbf1600ea, 32'hbed4f729} /* (3, 27, 24) {real, imag} */,
  {32'h3eadb976, 32'hc0054f4c} /* (3, 27, 23) {real, imag} */,
  {32'hbf295958, 32'hc01c97ca} /* (3, 27, 22) {real, imag} */,
  {32'hbfbea8f2, 32'h3f27930c} /* (3, 27, 21) {real, imag} */,
  {32'hbf819448, 32'hbf8a5e8b} /* (3, 27, 20) {real, imag} */,
  {32'h402050d3, 32'h3eeb67fe} /* (3, 27, 19) {real, imag} */,
  {32'h3f694081, 32'hbe9836f1} /* (3, 27, 18) {real, imag} */,
  {32'h3eaadfd5, 32'h3fe665ec} /* (3, 27, 17) {real, imag} */,
  {32'hbf294277, 32'hbea059ab} /* (3, 27, 16) {real, imag} */,
  {32'h3f740595, 32'h3f7e7b2a} /* (3, 27, 15) {real, imag} */,
  {32'hbf8e5633, 32'hbfc5ef5e} /* (3, 27, 14) {real, imag} */,
  {32'h3f80ea06, 32'hbf964e86} /* (3, 27, 13) {real, imag} */,
  {32'hbf7f3e07, 32'hbf052055} /* (3, 27, 12) {real, imag} */,
  {32'hbed9d6fd, 32'h3fc56f45} /* (3, 27, 11) {real, imag} */,
  {32'hc0009519, 32'h3ef07d34} /* (3, 27, 10) {real, imag} */,
  {32'h3f95e49e, 32'hbf4bca09} /* (3, 27, 9) {real, imag} */,
  {32'h4018534e, 32'h405473d5} /* (3, 27, 8) {real, imag} */,
  {32'h4065f808, 32'hbf62a152} /* (3, 27, 7) {real, imag} */,
  {32'h3faa53cc, 32'hbfa0d492} /* (3, 27, 6) {real, imag} */,
  {32'hc09f7f55, 32'h40c9d929} /* (3, 27, 5) {real, imag} */,
  {32'h4042e185, 32'hc087bcf0} /* (3, 27, 4) {real, imag} */,
  {32'hbf4bedf7, 32'h3fa76212} /* (3, 27, 3) {real, imag} */,
  {32'hc104dcb9, 32'h40d7ca2a} /* (3, 27, 2) {real, imag} */,
  {32'hbfa53227, 32'hc15f877d} /* (3, 27, 1) {real, imag} */,
  {32'h409b5e1d, 32'hc18c1f9a} /* (3, 27, 0) {real, imag} */,
  {32'hbe510fc5, 32'hc0805452} /* (3, 26, 31) {real, imag} */,
  {32'hc011bdef, 32'hc0108219} /* (3, 26, 30) {real, imag} */,
  {32'h3fbc5b66, 32'h3e95a4fa} /* (3, 26, 29) {real, imag} */,
  {32'h40641de8, 32'h3fcae0a0} /* (3, 26, 28) {real, imag} */,
  {32'h3ff69762, 32'h3f55db08} /* (3, 26, 27) {real, imag} */,
  {32'h40058633, 32'h40b41a1f} /* (3, 26, 26) {real, imag} */,
  {32'hc067987d, 32'h407a6bf3} /* (3, 26, 25) {real, imag} */,
  {32'h407e06ba, 32'h3fad576e} /* (3, 26, 24) {real, imag} */,
  {32'hc08f3d36, 32'hc05a82a9} /* (3, 26, 23) {real, imag} */,
  {32'h3eebc1fb, 32'hbe0095f1} /* (3, 26, 22) {real, imag} */,
  {32'hbfff8106, 32'h40819498} /* (3, 26, 21) {real, imag} */,
  {32'h3eb05a8b, 32'h3e4aa71a} /* (3, 26, 20) {real, imag} */,
  {32'hbfe44311, 32'hbe989ca2} /* (3, 26, 19) {real, imag} */,
  {32'hbfb9712d, 32'hbfba2898} /* (3, 26, 18) {real, imag} */,
  {32'h3db04820, 32'hbf6b353f} /* (3, 26, 17) {real, imag} */,
  {32'hbeb56cbf, 32'hbf22c8a3} /* (3, 26, 16) {real, imag} */,
  {32'h3fe410c2, 32'hbf5f6214} /* (3, 26, 15) {real, imag} */,
  {32'h3fb5906f, 32'hbeea608c} /* (3, 26, 14) {real, imag} */,
  {32'hc014850c, 32'hc04d6778} /* (3, 26, 13) {real, imag} */,
  {32'hbf6d70de, 32'hbfa8dd03} /* (3, 26, 12) {real, imag} */,
  {32'h3ee92302, 32'h3f1fff3f} /* (3, 26, 11) {real, imag} */,
  {32'hbe124e47, 32'h406a1d05} /* (3, 26, 10) {real, imag} */,
  {32'hbf5d426d, 32'hbed07e43} /* (3, 26, 9) {real, imag} */,
  {32'hbfb2a01c, 32'hbf374b37} /* (3, 26, 8) {real, imag} */,
  {32'h401c1439, 32'h4099b8ed} /* (3, 26, 7) {real, imag} */,
  {32'hbfb8f00c, 32'h3eabd345} /* (3, 26, 6) {real, imag} */,
  {32'h400f3c84, 32'h3f91377d} /* (3, 26, 5) {real, imag} */,
  {32'h400783f1, 32'h406afb2d} /* (3, 26, 4) {real, imag} */,
  {32'h407f5110, 32'hbfa67f5c} /* (3, 26, 3) {real, imag} */,
  {32'h3fa4570c, 32'hbf691bea} /* (3, 26, 2) {real, imag} */,
  {32'h3fbd0033, 32'hbf8526ed} /* (3, 26, 1) {real, imag} */,
  {32'h40296a32, 32'hc08b4469} /* (3, 26, 0) {real, imag} */,
  {32'h40979fb9, 32'h40da823d} /* (3, 25, 31) {real, imag} */,
  {32'hc0c581cd, 32'h402708de} /* (3, 25, 30) {real, imag} */,
  {32'h3f94e39a, 32'hc00e2e11} /* (3, 25, 29) {real, imag} */,
  {32'h4003a2d5, 32'h404a54eb} /* (3, 25, 28) {real, imag} */,
  {32'hc04c39d2, 32'h3fcd3a61} /* (3, 25, 27) {real, imag} */,
  {32'hc0390e10, 32'h3ff8addf} /* (3, 25, 26) {real, imag} */,
  {32'hbfa46db7, 32'hbf1b823b} /* (3, 25, 25) {real, imag} */,
  {32'h3f616f30, 32'hc0bad4d6} /* (3, 25, 24) {real, imag} */,
  {32'h3fd55819, 32'h3fefc7f3} /* (3, 25, 23) {real, imag} */,
  {32'hc01f4648, 32'h40102a09} /* (3, 25, 22) {real, imag} */,
  {32'h3fd30c5b, 32'hbf5b5700} /* (3, 25, 21) {real, imag} */,
  {32'hbf891ff0, 32'h3fba7cf5} /* (3, 25, 20) {real, imag} */,
  {32'h3f25a7ea, 32'hbff95b86} /* (3, 25, 19) {real, imag} */,
  {32'hbeecfead, 32'hbee8a575} /* (3, 25, 18) {real, imag} */,
  {32'h3f6c6876, 32'hbfb1085b} /* (3, 25, 17) {real, imag} */,
  {32'hbffc8f02, 32'h3f66c8e7} /* (3, 25, 16) {real, imag} */,
  {32'hbea4098e, 32'hc033a229} /* (3, 25, 15) {real, imag} */,
  {32'hbf9b1fd8, 32'h3fa3b318} /* (3, 25, 14) {real, imag} */,
  {32'h3f9f1402, 32'h3f107ce9} /* (3, 25, 13) {real, imag} */,
  {32'h3e0fea22, 32'hc05d6e45} /* (3, 25, 12) {real, imag} */,
  {32'h3facb872, 32'h4014ec57} /* (3, 25, 11) {real, imag} */,
  {32'hbffc3631, 32'hbf77eb87} /* (3, 25, 10) {real, imag} */,
  {32'hbf8b0bec, 32'h3f8efeea} /* (3, 25, 9) {real, imag} */,
  {32'hbeeaf237, 32'hbfb04e84} /* (3, 25, 8) {real, imag} */,
  {32'h3f01d1d1, 32'hc0adf394} /* (3, 25, 7) {real, imag} */,
  {32'h3f5f808a, 32'hbfbda42b} /* (3, 25, 6) {real, imag} */,
  {32'hc003fea2, 32'h3fddff3f} /* (3, 25, 5) {real, imag} */,
  {32'h40a21fcc, 32'hc07aab26} /* (3, 25, 4) {real, imag} */,
  {32'h408793fd, 32'hc03eeb1a} /* (3, 25, 3) {real, imag} */,
  {32'h3e031459, 32'h3fc25400} /* (3, 25, 2) {real, imag} */,
  {32'h3f8b9872, 32'h4087f436} /* (3, 25, 1) {real, imag} */,
  {32'h3ff0c19f, 32'h40f16b33} /* (3, 25, 0) {real, imag} */,
  {32'hc0a9e787, 32'hc0a03b31} /* (3, 24, 31) {real, imag} */,
  {32'h404b968b, 32'hc00846c9} /* (3, 24, 30) {real, imag} */,
  {32'h4023808f, 32'h406aaa5a} /* (3, 24, 29) {real, imag} */,
  {32'hbf7b7c0d, 32'h3fa2c5ea} /* (3, 24, 28) {real, imag} */,
  {32'h3ed1ad44, 32'h40acbf54} /* (3, 24, 27) {real, imag} */,
  {32'h405a6f54, 32'hbfa9b800} /* (3, 24, 26) {real, imag} */,
  {32'h4065981d, 32'hbfdfa151} /* (3, 24, 25) {real, imag} */,
  {32'h3feaccaf, 32'hbff7a712} /* (3, 24, 24) {real, imag} */,
  {32'hc04647a1, 32'h3fd53ee6} /* (3, 24, 23) {real, imag} */,
  {32'hbf1b6b9c, 32'hc099d531} /* (3, 24, 22) {real, imag} */,
  {32'h40a1dbf7, 32'h3f8fab7f} /* (3, 24, 21) {real, imag} */,
  {32'hbdd03108, 32'h3ff91c23} /* (3, 24, 20) {real, imag} */,
  {32'hc0192f1c, 32'h3f0b64f5} /* (3, 24, 19) {real, imag} */,
  {32'h3f674755, 32'h3f9aa3e4} /* (3, 24, 18) {real, imag} */,
  {32'hc05556e2, 32'hbeb0ca37} /* (3, 24, 17) {real, imag} */,
  {32'hbed5d46e, 32'h3e92e09a} /* (3, 24, 16) {real, imag} */,
  {32'h3fd43ab4, 32'hbeef01a9} /* (3, 24, 15) {real, imag} */,
  {32'h3ed197cf, 32'h3f5231a9} /* (3, 24, 14) {real, imag} */,
  {32'h3f7fbff1, 32'h3fc8e866} /* (3, 24, 13) {real, imag} */,
  {32'hbfa2d17d, 32'hbf4492a0} /* (3, 24, 12) {real, imag} */,
  {32'hbf2e7e65, 32'hc0151356} /* (3, 24, 11) {real, imag} */,
  {32'h3fda9f9e, 32'h3f189195} /* (3, 24, 10) {real, imag} */,
  {32'h3f7af86b, 32'hc0a6cd17} /* (3, 24, 9) {real, imag} */,
  {32'hc027f2c8, 32'hbf06dda0} /* (3, 24, 8) {real, imag} */,
  {32'h3f267825, 32'hc0276162} /* (3, 24, 7) {real, imag} */,
  {32'hbecd92d3, 32'hbf9cf727} /* (3, 24, 6) {real, imag} */,
  {32'hc0047e8f, 32'hc057981a} /* (3, 24, 5) {real, imag} */,
  {32'h4050ef37, 32'hbfe6d226} /* (3, 24, 4) {real, imag} */,
  {32'hc0d78b74, 32'h3f5a018d} /* (3, 24, 3) {real, imag} */,
  {32'h3f2408b6, 32'h41052180} /* (3, 24, 2) {real, imag} */,
  {32'h3f239ee9, 32'hc120d26f} /* (3, 24, 1) {real, imag} */,
  {32'hbd176c8a, 32'hc07c3f61} /* (3, 24, 0) {real, imag} */,
  {32'hc02db620, 32'h403d5a47} /* (3, 23, 31) {real, imag} */,
  {32'hbd462a9f, 32'hc0193ff0} /* (3, 23, 30) {real, imag} */,
  {32'hbe9a7d33, 32'h3ca68d07} /* (3, 23, 29) {real, imag} */,
  {32'hbfe2dd39, 32'hbf2bdc69} /* (3, 23, 28) {real, imag} */,
  {32'h40025dde, 32'h3ed854b6} /* (3, 23, 27) {real, imag} */,
  {32'hc0205876, 32'h3eef2ffd} /* (3, 23, 26) {real, imag} */,
  {32'hbf8ab9dd, 32'h403d4cc5} /* (3, 23, 25) {real, imag} */,
  {32'hc023b575, 32'hbfce6c6d} /* (3, 23, 24) {real, imag} */,
  {32'h3eb7562a, 32'h3d246c66} /* (3, 23, 23) {real, imag} */,
  {32'h3ff00d24, 32'hbfb95e19} /* (3, 23, 22) {real, imag} */,
  {32'hbf1b4cae, 32'h4008ef81} /* (3, 23, 21) {real, imag} */,
  {32'h3c73b8ad, 32'h4021f5a8} /* (3, 23, 20) {real, imag} */,
  {32'hbff6497d, 32'h3f8c1629} /* (3, 23, 19) {real, imag} */,
  {32'h3f6751d8, 32'h3fd1a2cf} /* (3, 23, 18) {real, imag} */,
  {32'h40261193, 32'h3f163843} /* (3, 23, 17) {real, imag} */,
  {32'h3e8e6524, 32'h3fadc811} /* (3, 23, 16) {real, imag} */,
  {32'h3f75cd59, 32'h4043e2b8} /* (3, 23, 15) {real, imag} */,
  {32'hbf05f899, 32'hbf81fe11} /* (3, 23, 14) {real, imag} */,
  {32'h408071ec, 32'hbff1b9c8} /* (3, 23, 13) {real, imag} */,
  {32'hbda82ec8, 32'h40500d4d} /* (3, 23, 12) {real, imag} */,
  {32'hc0000967, 32'hbf9d3222} /* (3, 23, 11) {real, imag} */,
  {32'hbfa4a644, 32'hbe7df0a9} /* (3, 23, 10) {real, imag} */,
  {32'h402313f7, 32'hbf05fc8a} /* (3, 23, 9) {real, imag} */,
  {32'hbff66746, 32'h3dc05568} /* (3, 23, 8) {real, imag} */,
  {32'h3dc88c71, 32'hbe878877} /* (3, 23, 7) {real, imag} */,
  {32'h3f26fda4, 32'hbfedf074} /* (3, 23, 6) {real, imag} */,
  {32'hc08b7cb2, 32'hbff506f6} /* (3, 23, 5) {real, imag} */,
  {32'h400bd30b, 32'hbfb355f8} /* (3, 23, 4) {real, imag} */,
  {32'h3fd4f7ff, 32'h3f18b9e0} /* (3, 23, 3) {real, imag} */,
  {32'hbfe81209, 32'hbf9983e8} /* (3, 23, 2) {real, imag} */,
  {32'h40d30aea, 32'hc03317cf} /* (3, 23, 1) {real, imag} */,
  {32'h3fbd1da9, 32'h3fffc696} /* (3, 23, 0) {real, imag} */,
  {32'hbfcf2c1c, 32'hbe8f0960} /* (3, 22, 31) {real, imag} */,
  {32'h4056c07d, 32'hbe3d80d4} /* (3, 22, 30) {real, imag} */,
  {32'h40b6edaa, 32'hc068460f} /* (3, 22, 29) {real, imag} */,
  {32'hbf0cec6c, 32'hc0901a8e} /* (3, 22, 28) {real, imag} */,
  {32'hc018eecf, 32'hc0103dbd} /* (3, 22, 27) {real, imag} */,
  {32'hc00afb57, 32'h3e93fa92} /* (3, 22, 26) {real, imag} */,
  {32'hc050fbc9, 32'hbf6627d3} /* (3, 22, 25) {real, imag} */,
  {32'h3ed2e8d2, 32'h3fcfad12} /* (3, 22, 24) {real, imag} */,
  {32'h3ff701fe, 32'hc05076fd} /* (3, 22, 23) {real, imag} */,
  {32'h3fd00c92, 32'hbe43d882} /* (3, 22, 22) {real, imag} */,
  {32'hbf0ed199, 32'h40006cb9} /* (3, 22, 21) {real, imag} */,
  {32'hbedaf5d2, 32'h3fd68117} /* (3, 22, 20) {real, imag} */,
  {32'h40371cb5, 32'hc0878ab1} /* (3, 22, 19) {real, imag} */,
  {32'h3fb0e7f7, 32'h3fcafbbc} /* (3, 22, 18) {real, imag} */,
  {32'hbf5809b8, 32'hbf476f28} /* (3, 22, 17) {real, imag} */,
  {32'hbfb1e1b7, 32'h3e969af5} /* (3, 22, 16) {real, imag} */,
  {32'hbf398aff, 32'hbe1a7346} /* (3, 22, 15) {real, imag} */,
  {32'hc0448abf, 32'h3fdeee58} /* (3, 22, 14) {real, imag} */,
  {32'hbf9151e2, 32'hbc58370a} /* (3, 22, 13) {real, imag} */,
  {32'hbe1199da, 32'h3fc98058} /* (3, 22, 12) {real, imag} */,
  {32'h40616794, 32'hbf9fa4d2} /* (3, 22, 11) {real, imag} */,
  {32'hbf11ae5e, 32'h3fb0424e} /* (3, 22, 10) {real, imag} */,
  {32'hbfa0efef, 32'hbf01b3e3} /* (3, 22, 9) {real, imag} */,
  {32'h401fd116, 32'hbf3b227e} /* (3, 22, 8) {real, imag} */,
  {32'hc09e3d94, 32'h3e9e0f11} /* (3, 22, 7) {real, imag} */,
  {32'hbe7c455b, 32'hbf035924} /* (3, 22, 6) {real, imag} */,
  {32'hc05bf3f1, 32'h3f6aafcb} /* (3, 22, 5) {real, imag} */,
  {32'h3fdf16f1, 32'h40c857b5} /* (3, 22, 4) {real, imag} */,
  {32'hbd01198b, 32'h402c7112} /* (3, 22, 3) {real, imag} */,
  {32'hc0ba47c1, 32'hc093c12e} /* (3, 22, 2) {real, imag} */,
  {32'h4068891e, 32'h3fd882d4} /* (3, 22, 1) {real, imag} */,
  {32'h4019aa3c, 32'h400fb0c7} /* (3, 22, 0) {real, imag} */,
  {32'hc05ece4f, 32'hbfe6b75e} /* (3, 21, 31) {real, imag} */,
  {32'h403619c6, 32'h3fa46289} /* (3, 21, 30) {real, imag} */,
  {32'h406166c6, 32'h3ea38925} /* (3, 21, 29) {real, imag} */,
  {32'h403000f7, 32'h3e8ab97c} /* (3, 21, 28) {real, imag} */,
  {32'hbfc5391b, 32'hbfbdb286} /* (3, 21, 27) {real, imag} */,
  {32'h401fcbd3, 32'h40429d41} /* (3, 21, 26) {real, imag} */,
  {32'hbe390945, 32'hbf24491b} /* (3, 21, 25) {real, imag} */,
  {32'hbd089bcc, 32'hbedb3540} /* (3, 21, 24) {real, imag} */,
  {32'h3f23a9af, 32'h3facb08a} /* (3, 21, 23) {real, imag} */,
  {32'h40139faa, 32'h3ea676c2} /* (3, 21, 22) {real, imag} */,
  {32'hc002dc43, 32'h3e1838a6} /* (3, 21, 21) {real, imag} */,
  {32'hbec3e153, 32'hc02b8f5a} /* (3, 21, 20) {real, imag} */,
  {32'h3feba3b4, 32'hbf02890c} /* (3, 21, 19) {real, imag} */,
  {32'hc05626b4, 32'hc00667ef} /* (3, 21, 18) {real, imag} */,
  {32'hbf3f051a, 32'h3fc05928} /* (3, 21, 17) {real, imag} */,
  {32'h3dee8838, 32'h3d2ddb5f} /* (3, 21, 16) {real, imag} */,
  {32'h3f8c2c92, 32'hbfeb7d36} /* (3, 21, 15) {real, imag} */,
  {32'hc0217535, 32'h3f259d26} /* (3, 21, 14) {real, imag} */,
  {32'hbfb255dc, 32'h3ede9ee0} /* (3, 21, 13) {real, imag} */,
  {32'h3f706995, 32'h3f6c161d} /* (3, 21, 12) {real, imag} */,
  {32'hbf504858, 32'h40344af2} /* (3, 21, 11) {real, imag} */,
  {32'h3f86bdd3, 32'hbf641b1e} /* (3, 21, 10) {real, imag} */,
  {32'h3e675383, 32'hc00ba37c} /* (3, 21, 9) {real, imag} */,
  {32'h401fb101, 32'hc041ab36} /* (3, 21, 8) {real, imag} */,
  {32'hc02dd570, 32'hc0077429} /* (3, 21, 7) {real, imag} */,
  {32'hbfae1640, 32'hc0094f11} /* (3, 21, 6) {real, imag} */,
  {32'h4011d379, 32'hbfca5d9e} /* (3, 21, 5) {real, imag} */,
  {32'hc04967a3, 32'h403ebd41} /* (3, 21, 4) {real, imag} */,
  {32'h3e9b52a0, 32'h3f685c64} /* (3, 21, 3) {real, imag} */,
  {32'h400acfb2, 32'h4095caf1} /* (3, 21, 2) {real, imag} */,
  {32'hbf8f65e5, 32'hbfb766ee} /* (3, 21, 1) {real, imag} */,
  {32'hc05bfe06, 32'hc005d76c} /* (3, 21, 0) {real, imag} */,
  {32'h3f0c58b2, 32'h3f892c06} /* (3, 20, 31) {real, imag} */,
  {32'h3ec8e986, 32'hc004f041} /* (3, 20, 30) {real, imag} */,
  {32'hbc15d4b2, 32'h3f213b10} /* (3, 20, 29) {real, imag} */,
  {32'h3f04ee13, 32'h3f54018f} /* (3, 20, 28) {real, imag} */,
  {32'h3fcb5d26, 32'hbf205133} /* (3, 20, 27) {real, imag} */,
  {32'h3f9f1f45, 32'h3eed64bd} /* (3, 20, 26) {real, imag} */,
  {32'hc0b931d4, 32'hc02bfbf4} /* (3, 20, 25) {real, imag} */,
  {32'h4037589b, 32'h3e205053} /* (3, 20, 24) {real, imag} */,
  {32'h3d377092, 32'h3d26edaf} /* (3, 20, 23) {real, imag} */,
  {32'h4013ee33, 32'hbe03e858} /* (3, 20, 22) {real, imag} */,
  {32'hbfd70437, 32'hbe8ec548} /* (3, 20, 21) {real, imag} */,
  {32'h3fc27083, 32'hc01a3065} /* (3, 20, 20) {real, imag} */,
  {32'hbf87e13c, 32'hbff92bfa} /* (3, 20, 19) {real, imag} */,
  {32'h3ee22726, 32'hbfc8d36a} /* (3, 20, 18) {real, imag} */,
  {32'h3de4178f, 32'h4013ce90} /* (3, 20, 17) {real, imag} */,
  {32'h3d946752, 32'hbe89e6c8} /* (3, 20, 16) {real, imag} */,
  {32'h3e36d29a, 32'h3fa18dbc} /* (3, 20, 15) {real, imag} */,
  {32'h3f28f55b, 32'h3f458025} /* (3, 20, 14) {real, imag} */,
  {32'hc03ca1eb, 32'hc0164ade} /* (3, 20, 13) {real, imag} */,
  {32'h3ee9985c, 32'hbe593939} /* (3, 20, 12) {real, imag} */,
  {32'h3f966488, 32'hbfca9487} /* (3, 20, 11) {real, imag} */,
  {32'hbd8f1fe1, 32'hbf2c8057} /* (3, 20, 10) {real, imag} */,
  {32'h3f2f721d, 32'hc05b3252} /* (3, 20, 9) {real, imag} */,
  {32'h3d17670b, 32'h3f12a7d8} /* (3, 20, 8) {real, imag} */,
  {32'h4067f208, 32'hbfc4a26d} /* (3, 20, 7) {real, imag} */,
  {32'hbec063de, 32'hbf26b9cf} /* (3, 20, 6) {real, imag} */,
  {32'hbbdaf5d3, 32'hbeb109ab} /* (3, 20, 5) {real, imag} */,
  {32'h3f110b75, 32'hbeb5c29a} /* (3, 20, 4) {real, imag} */,
  {32'h40863b71, 32'hbfdf89a9} /* (3, 20, 3) {real, imag} */,
  {32'hc01433f8, 32'h3fc00f3e} /* (3, 20, 2) {real, imag} */,
  {32'hc01a98ae, 32'h4024b903} /* (3, 20, 1) {real, imag} */,
  {32'h3febec95, 32'hbfb93cb3} /* (3, 20, 0) {real, imag} */,
  {32'hbe63a0f1, 32'hbe429669} /* (3, 19, 31) {real, imag} */,
  {32'hc03ac04e, 32'hbf46256e} /* (3, 19, 30) {real, imag} */,
  {32'hbf724e0e, 32'h3ffff77d} /* (3, 19, 29) {real, imag} */,
  {32'hbf4d9128, 32'h3e3e4c90} /* (3, 19, 28) {real, imag} */,
  {32'hbf59be1e, 32'h3eb1c8d4} /* (3, 19, 27) {real, imag} */,
  {32'h3f32ba70, 32'h3f9cba1e} /* (3, 19, 26) {real, imag} */,
  {32'h3ea529e5, 32'hbf899e6f} /* (3, 19, 25) {real, imag} */,
  {32'hc0307939, 32'h4065370e} /* (3, 19, 24) {real, imag} */,
  {32'h3ff39d05, 32'hc0267260} /* (3, 19, 23) {real, imag} */,
  {32'hbf74b723, 32'h3f4c333b} /* (3, 19, 22) {real, imag} */,
  {32'hbd455834, 32'hbe20ac2c} /* (3, 19, 21) {real, imag} */,
  {32'hbfdc1b19, 32'h3e41f404} /* (3, 19, 20) {real, imag} */,
  {32'hbe8b9889, 32'h3fe2658d} /* (3, 19, 19) {real, imag} */,
  {32'hbf40f0a1, 32'h3efba9d5} /* (3, 19, 18) {real, imag} */,
  {32'hbf804f3b, 32'h3f1b8258} /* (3, 19, 17) {real, imag} */,
  {32'hbd9884a2, 32'h3fb8f4f5} /* (3, 19, 16) {real, imag} */,
  {32'hbe5d751e, 32'h3ef5d5bf} /* (3, 19, 15) {real, imag} */,
  {32'h3f61f0fa, 32'h3eb82a6f} /* (3, 19, 14) {real, imag} */,
  {32'hbeea7738, 32'h401bf43a} /* (3, 19, 13) {real, imag} */,
  {32'hbf9710bb, 32'hbee328be} /* (3, 19, 12) {real, imag} */,
  {32'hbf83214b, 32'h40123cc2} /* (3, 19, 11) {real, imag} */,
  {32'hbfdbf469, 32'hbf42aed8} /* (3, 19, 10) {real, imag} */,
  {32'h4077de13, 32'h401efdbb} /* (3, 19, 9) {real, imag} */,
  {32'hbdf55df3, 32'hbf9ee859} /* (3, 19, 8) {real, imag} */,
  {32'hbf7ce6c1, 32'hbf51049e} /* (3, 19, 7) {real, imag} */,
  {32'hbf5716c7, 32'h3fcb4fca} /* (3, 19, 6) {real, imag} */,
  {32'hbe8d18e7, 32'h3fb4f2e4} /* (3, 19, 5) {real, imag} */,
  {32'hbfc0001d, 32'hbf300a04} /* (3, 19, 4) {real, imag} */,
  {32'h3fc609b4, 32'hbf847545} /* (3, 19, 3) {real, imag} */,
  {32'h3e73835b, 32'hbf3499c3} /* (3, 19, 2) {real, imag} */,
  {32'h40588c99, 32'h3ff38cc2} /* (3, 19, 1) {real, imag} */,
  {32'hbf5c9b6f, 32'h3fb20ddb} /* (3, 19, 0) {real, imag} */,
  {32'hc00e0096, 32'h3f00e6a2} /* (3, 18, 31) {real, imag} */,
  {32'hbeb32c97, 32'h3fc5c6bb} /* (3, 18, 30) {real, imag} */,
  {32'hbed6ef37, 32'hbf3bcf4c} /* (3, 18, 29) {real, imag} */,
  {32'hbfa16c17, 32'hbe3eba11} /* (3, 18, 28) {real, imag} */,
  {32'h3fdb78cf, 32'hbda9545f} /* (3, 18, 27) {real, imag} */,
  {32'hbeb7135e, 32'hbf067c63} /* (3, 18, 26) {real, imag} */,
  {32'h3f881e06, 32'hbf122bfb} /* (3, 18, 25) {real, imag} */,
  {32'h402a0056, 32'h3f165bac} /* (3, 18, 24) {real, imag} */,
  {32'hc07526b9, 32'hbf7e1eb6} /* (3, 18, 23) {real, imag} */,
  {32'h3fc123bd, 32'hc0211f79} /* (3, 18, 22) {real, imag} */,
  {32'h3f2fd6e0, 32'hc0473a73} /* (3, 18, 21) {real, imag} */,
  {32'h3fae3eae, 32'h3f7ef999} /* (3, 18, 20) {real, imag} */,
  {32'h3fd3d4ef, 32'hbfafd71a} /* (3, 18, 19) {real, imag} */,
  {32'hbfa021c1, 32'h3fac7201} /* (3, 18, 18) {real, imag} */,
  {32'hbf51acef, 32'hbf5022c9} /* (3, 18, 17) {real, imag} */,
  {32'h3fce004a, 32'hbe8820b0} /* (3, 18, 16) {real, imag} */,
  {32'h3e97cb20, 32'hbf5023ff} /* (3, 18, 15) {real, imag} */,
  {32'hbf2e56e3, 32'hbfa2c76c} /* (3, 18, 14) {real, imag} */,
  {32'h3fb0006f, 32'hbfaced48} /* (3, 18, 13) {real, imag} */,
  {32'hbe7d80fa, 32'hbf1d1d64} /* (3, 18, 12) {real, imag} */,
  {32'hc0600f28, 32'hbee6ca44} /* (3, 18, 11) {real, imag} */,
  {32'h3f525efa, 32'hbfdc9aa5} /* (3, 18, 10) {real, imag} */,
  {32'h3f16703a, 32'hbf9e327c} /* (3, 18, 9) {real, imag} */,
  {32'hbf8007c4, 32'h40536366} /* (3, 18, 8) {real, imag} */,
  {32'h4017085d, 32'h3f6831ce} /* (3, 18, 7) {real, imag} */,
  {32'hbf9723d5, 32'h3e0fabe7} /* (3, 18, 6) {real, imag} */,
  {32'hbce7ddff, 32'h3dd08929} /* (3, 18, 5) {real, imag} */,
  {32'hbe411eb4, 32'hbfa0a940} /* (3, 18, 4) {real, imag} */,
  {32'hbfcf9644, 32'hbf167e11} /* (3, 18, 3) {real, imag} */,
  {32'hbe93bb90, 32'h4030c050} /* (3, 18, 2) {real, imag} */,
  {32'hc04ebba2, 32'hbffe631a} /* (3, 18, 1) {real, imag} */,
  {32'hc037dfcf, 32'h3f431e85} /* (3, 18, 0) {real, imag} */,
  {32'h3f2390a4, 32'h3f373077} /* (3, 17, 31) {real, imag} */,
  {32'hbf309309, 32'h3ef0af2b} /* (3, 17, 30) {real, imag} */,
  {32'hbf26fa04, 32'h3edf2b3d} /* (3, 17, 29) {real, imag} */,
  {32'hbe523f73, 32'hbfd5dda8} /* (3, 17, 28) {real, imag} */,
  {32'h3f64e83c, 32'h3f7f9281} /* (3, 17, 27) {real, imag} */,
  {32'hbed4ea9e, 32'hbf5440ac} /* (3, 17, 26) {real, imag} */,
  {32'h3f82c651, 32'hbf202b01} /* (3, 17, 25) {real, imag} */,
  {32'hbf674865, 32'hbfa55e4b} /* (3, 17, 24) {real, imag} */,
  {32'h3e812acb, 32'hbfa267fd} /* (3, 17, 23) {real, imag} */,
  {32'hbfb53341, 32'h3f9f9211} /* (3, 17, 22) {real, imag} */,
  {32'hbb37cefe, 32'hbe16330e} /* (3, 17, 21) {real, imag} */,
  {32'hbf3ce433, 32'hbf171a69} /* (3, 17, 20) {real, imag} */,
  {32'h3db821e8, 32'h3ec0e8d2} /* (3, 17, 19) {real, imag} */,
  {32'hbb8b218b, 32'hc0245f10} /* (3, 17, 18) {real, imag} */,
  {32'hbf0541a3, 32'h3e4fddc1} /* (3, 17, 17) {real, imag} */,
  {32'hbff056f1, 32'h3e5b9e7f} /* (3, 17, 16) {real, imag} */,
  {32'h3f42097b, 32'h3f5a7f06} /* (3, 17, 15) {real, imag} */,
  {32'hbfb0dd9d, 32'h3f9330a6} /* (3, 17, 14) {real, imag} */,
  {32'hbfdf5e4d, 32'h40164642} /* (3, 17, 13) {real, imag} */,
  {32'hbfab9f40, 32'h400c82d5} /* (3, 17, 12) {real, imag} */,
  {32'hbf8b92f3, 32'hc00242c2} /* (3, 17, 11) {real, imag} */,
  {32'h3fa9427d, 32'hbf8bd9aa} /* (3, 17, 10) {real, imag} */,
  {32'h3f98b4b5, 32'hbe9b3de1} /* (3, 17, 9) {real, imag} */,
  {32'h3fa218fd, 32'h3da36cdc} /* (3, 17, 8) {real, imag} */,
  {32'h3f9fe945, 32'hbdbe7ecf} /* (3, 17, 7) {real, imag} */,
  {32'h3f765d32, 32'hbdded79f} /* (3, 17, 6) {real, imag} */,
  {32'h3fb46db7, 32'hbd88787a} /* (3, 17, 5) {real, imag} */,
  {32'hbf1ee632, 32'hbe9b7c50} /* (3, 17, 4) {real, imag} */,
  {32'hc02b689f, 32'h3f89eef1} /* (3, 17, 3) {real, imag} */,
  {32'hbf3e848b, 32'h3eccc229} /* (3, 17, 2) {real, imag} */,
  {32'h404a11c4, 32'hbfd1936a} /* (3, 17, 1) {real, imag} */,
  {32'hbfded959, 32'h3f5c665c} /* (3, 17, 0) {real, imag} */,
  {32'hbe44ba32, 32'hbdd32852} /* (3, 16, 31) {real, imag} */,
  {32'h3e79f529, 32'hbca8bed9} /* (3, 16, 30) {real, imag} */,
  {32'h3f8d257f, 32'h3fd14f91} /* (3, 16, 29) {real, imag} */,
  {32'h3ec708bf, 32'hbdb2de16} /* (3, 16, 28) {real, imag} */,
  {32'h3f0f254c, 32'hbf23846e} /* (3, 16, 27) {real, imag} */,
  {32'h3e37ba2f, 32'hbf3c45c2} /* (3, 16, 26) {real, imag} */,
  {32'hbf94058c, 32'h3f97ba66} /* (3, 16, 25) {real, imag} */,
  {32'h3ff273fa, 32'hbfb763eb} /* (3, 16, 24) {real, imag} */,
  {32'h3e978e9d, 32'h3ee1c9b7} /* (3, 16, 23) {real, imag} */,
  {32'hbf56aa10, 32'h3fd2987f} /* (3, 16, 22) {real, imag} */,
  {32'hbf2e79b3, 32'hbf5c1159} /* (3, 16, 21) {real, imag} */,
  {32'hbee98c1d, 32'h3f93ebec} /* (3, 16, 20) {real, imag} */,
  {32'h3eb1b425, 32'h3f38d2d8} /* (3, 16, 19) {real, imag} */,
  {32'h3faf79b2, 32'h3f3c4d7d} /* (3, 16, 18) {real, imag} */,
  {32'hbe8b0286, 32'hbed385fa} /* (3, 16, 17) {real, imag} */,
  {32'h3e5e0899, 32'hbee978f8} /* (3, 16, 16) {real, imag} */,
  {32'h3fd4d416, 32'hbe6a4452} /* (3, 16, 15) {real, imag} */,
  {32'h3f849911, 32'hbfab3f16} /* (3, 16, 14) {real, imag} */,
  {32'hbf4f9155, 32'h3f535912} /* (3, 16, 13) {real, imag} */,
  {32'hbfa2127d, 32'h3ee32dde} /* (3, 16, 12) {real, imag} */,
  {32'hc0347a74, 32'h3ecdf961} /* (3, 16, 11) {real, imag} */,
  {32'hbd307ada, 32'hbe816f4d} /* (3, 16, 10) {real, imag} */,
  {32'h3e544c41, 32'hbe16fd9a} /* (3, 16, 9) {real, imag} */,
  {32'h3f631e0b, 32'hbf4bce93} /* (3, 16, 8) {real, imag} */,
  {32'hbf4bb3fd, 32'hbed5f114} /* (3, 16, 7) {real, imag} */,
  {32'h3e048498, 32'h3f483315} /* (3, 16, 6) {real, imag} */,
  {32'h3e79a41e, 32'h3f2ca988} /* (3, 16, 5) {real, imag} */,
  {32'hbf94dd90, 32'hbfb97693} /* (3, 16, 4) {real, imag} */,
  {32'hbfaae10f, 32'h3ef2c36b} /* (3, 16, 3) {real, imag} */,
  {32'h3f34fe48, 32'hbebb495d} /* (3, 16, 2) {real, imag} */,
  {32'hbe4a68b7, 32'hbf58ef6f} /* (3, 16, 1) {real, imag} */,
  {32'h3f4c1dc6, 32'hbfd43828} /* (3, 16, 0) {real, imag} */,
  {32'hbfa762a9, 32'h3f44c9df} /* (3, 15, 31) {real, imag} */,
  {32'h40275438, 32'h3f2c5b78} /* (3, 15, 30) {real, imag} */,
  {32'hbf7865ce, 32'h3f50679c} /* (3, 15, 29) {real, imag} */,
  {32'hbf488ad2, 32'h3ebd3558} /* (3, 15, 28) {real, imag} */,
  {32'h3decdbae, 32'h3d9d0677} /* (3, 15, 27) {real, imag} */,
  {32'hbfb5b1a1, 32'hbf8059d0} /* (3, 15, 26) {real, imag} */,
  {32'hbe3b8c07, 32'h3fbe9a41} /* (3, 15, 25) {real, imag} */,
  {32'hbfacdaf1, 32'h3f1fdcd8} /* (3, 15, 24) {real, imag} */,
  {32'h3ef70fc1, 32'hbf49e99c} /* (3, 15, 23) {real, imag} */,
  {32'hc07f57c6, 32'hc01840e3} /* (3, 15, 22) {real, imag} */,
  {32'h400569f4, 32'hbec98163} /* (3, 15, 21) {real, imag} */,
  {32'hbf1f3c3d, 32'hbfe33c5e} /* (3, 15, 20) {real, imag} */,
  {32'hbfa951ee, 32'h3e4fcd1f} /* (3, 15, 19) {real, imag} */,
  {32'hbed8e380, 32'h3fadb8fc} /* (3, 15, 18) {real, imag} */,
  {32'h3f8695b4, 32'h3f10414c} /* (3, 15, 17) {real, imag} */,
  {32'hbfa85a60, 32'h3ed881c4} /* (3, 15, 16) {real, imag} */,
  {32'h3ed5d220, 32'hbeb511e7} /* (3, 15, 15) {real, imag} */,
  {32'h3dfb7a8b, 32'h3fbb5699} /* (3, 15, 14) {real, imag} */,
  {32'h3f9d2975, 32'hbfa3ad7d} /* (3, 15, 13) {real, imag} */,
  {32'h3f49c3cc, 32'hbe09c72b} /* (3, 15, 12) {real, imag} */,
  {32'h3e036e4c, 32'h4042f3fb} /* (3, 15, 11) {real, imag} */,
  {32'hbf5639d0, 32'hbef3feb7} /* (3, 15, 10) {real, imag} */,
  {32'h3e9f04b7, 32'h3fb4a5ef} /* (3, 15, 9) {real, imag} */,
  {32'hbf905e43, 32'h3dfaf710} /* (3, 15, 8) {real, imag} */,
  {32'hbf3f90e2, 32'hbf3b91f3} /* (3, 15, 7) {real, imag} */,
  {32'h3f7522f6, 32'hbe0ebe80} /* (3, 15, 6) {real, imag} */,
  {32'hbff032f4, 32'h3fa4a978} /* (3, 15, 5) {real, imag} */,
  {32'hbf011f08, 32'hbfb17fde} /* (3, 15, 4) {real, imag} */,
  {32'h3cb5cdad, 32'h3f80074e} /* (3, 15, 3) {real, imag} */,
  {32'h4082c94f, 32'h3f6eb0c0} /* (3, 15, 2) {real, imag} */,
  {32'hbfc2ee23, 32'h3f8d7b80} /* (3, 15, 1) {real, imag} */,
  {32'hbd32f800, 32'h3f0b13ee} /* (3, 15, 0) {real, imag} */,
  {32'h401a4490, 32'h3f42ce48} /* (3, 14, 31) {real, imag} */,
  {32'hbff33bd2, 32'h3f850070} /* (3, 14, 30) {real, imag} */,
  {32'hbe8df4b0, 32'hbebb022d} /* (3, 14, 29) {real, imag} */,
  {32'h3f50a0ab, 32'hbf3db0b2} /* (3, 14, 28) {real, imag} */,
  {32'hbff85413, 32'h3f4368e3} /* (3, 14, 27) {real, imag} */,
  {32'h3f2b225b, 32'hbf6cd580} /* (3, 14, 26) {real, imag} */,
  {32'h3fc05634, 32'h3ee1a1a3} /* (3, 14, 25) {real, imag} */,
  {32'h3fee803e, 32'h3f4fefa6} /* (3, 14, 24) {real, imag} */,
  {32'hbfbd0880, 32'h3fd68714} /* (3, 14, 23) {real, imag} */,
  {32'h4008c0c8, 32'h3f3b67f7} /* (3, 14, 22) {real, imag} */,
  {32'hbc7913de, 32'h4023f77c} /* (3, 14, 21) {real, imag} */,
  {32'h3fde4a4e, 32'hbdbc5896} /* (3, 14, 20) {real, imag} */,
  {32'hc00438fa, 32'h40023de7} /* (3, 14, 19) {real, imag} */,
  {32'hbe8972f2, 32'hbebee70b} /* (3, 14, 18) {real, imag} */,
  {32'hc00966a3, 32'hbfe83a17} /* (3, 14, 17) {real, imag} */,
  {32'hbe9e9381, 32'hbf239fde} /* (3, 14, 16) {real, imag} */,
  {32'h3f26a8e0, 32'h3f0a8ec2} /* (3, 14, 15) {real, imag} */,
  {32'hbf620dfb, 32'hbe4c9218} /* (3, 14, 14) {real, imag} */,
  {32'hc0058451, 32'h3fa56953} /* (3, 14, 13) {real, imag} */,
  {32'h3e8061bc, 32'hbfcdd507} /* (3, 14, 12) {real, imag} */,
  {32'hbe754814, 32'hbfa3b26f} /* (3, 14, 11) {real, imag} */,
  {32'hbdbb3b8c, 32'h402717d6} /* (3, 14, 10) {real, imag} */,
  {32'h3fafd817, 32'hbef1a359} /* (3, 14, 9) {real, imag} */,
  {32'hbf51cc45, 32'h3e579328} /* (3, 14, 8) {real, imag} */,
  {32'hbf02c8a5, 32'h401e70f1} /* (3, 14, 7) {real, imag} */,
  {32'hbf1c6b34, 32'hc01bf9dc} /* (3, 14, 6) {real, imag} */,
  {32'hc02449b0, 32'hbfd512b8} /* (3, 14, 5) {real, imag} */,
  {32'h3f7ecba1, 32'hbff2303a} /* (3, 14, 4) {real, imag} */,
  {32'hbed08289, 32'hbf83168c} /* (3, 14, 3) {real, imag} */,
  {32'hc03a8403, 32'h3f289af3} /* (3, 14, 2) {real, imag} */,
  {32'h3f673561, 32'h3f1a3c4e} /* (3, 14, 1) {real, imag} */,
  {32'h3ee24657, 32'hbf1f3b1d} /* (3, 14, 0) {real, imag} */,
  {32'h3ee91e81, 32'hbea7b2e1} /* (3, 13, 31) {real, imag} */,
  {32'hc0494ed7, 32'h3edee00b} /* (3, 13, 30) {real, imag} */,
  {32'hbfb2c330, 32'h3d7d7eb3} /* (3, 13, 29) {real, imag} */,
  {32'h3f32866b, 32'hbf4e7484} /* (3, 13, 28) {real, imag} */,
  {32'h3e320476, 32'hbea922f5} /* (3, 13, 27) {real, imag} */,
  {32'h402deeca, 32'hbf51bd96} /* (3, 13, 26) {real, imag} */,
  {32'h3fc3b785, 32'h3f3f196e} /* (3, 13, 25) {real, imag} */,
  {32'h3fc8984f, 32'hbf115164} /* (3, 13, 24) {real, imag} */,
  {32'hbf30919a, 32'h3fae6bea} /* (3, 13, 23) {real, imag} */,
  {32'h3f5a7621, 32'hbe0039f8} /* (3, 13, 22) {real, imag} */,
  {32'h3fd72bd4, 32'h3f1351d3} /* (3, 13, 21) {real, imag} */,
  {32'hbfc48bf5, 32'hbf9b2433} /* (3, 13, 20) {real, imag} */,
  {32'hbfee7941, 32'h40237bc9} /* (3, 13, 19) {real, imag} */,
  {32'hbf1ac461, 32'hbe883e90} /* (3, 13, 18) {real, imag} */,
  {32'h3f605dae, 32'hbf959e22} /* (3, 13, 17) {real, imag} */,
  {32'h3f6ecf5a, 32'h3faf8b91} /* (3, 13, 16) {real, imag} */,
  {32'hbee1f1ff, 32'h3fe4848b} /* (3, 13, 15) {real, imag} */,
  {32'h3f620b19, 32'h3edb4a93} /* (3, 13, 14) {real, imag} */,
  {32'h3f480b55, 32'h3f5dd4cf} /* (3, 13, 13) {real, imag} */,
  {32'hc01866ed, 32'hbf287d6c} /* (3, 13, 12) {real, imag} */,
  {32'hc028fa43, 32'hc0403bad} /* (3, 13, 11) {real, imag} */,
  {32'h4000b2f3, 32'h3f875e64} /* (3, 13, 10) {real, imag} */,
  {32'h3ecba86f, 32'hbe20fcf6} /* (3, 13, 9) {real, imag} */,
  {32'hbf5b99bd, 32'hbf30192f} /* (3, 13, 8) {real, imag} */,
  {32'h3f554613, 32'h3f8d4464} /* (3, 13, 7) {real, imag} */,
  {32'hbf9896b1, 32'h401929f1} /* (3, 13, 6) {real, imag} */,
  {32'h3f8f3b1f, 32'hc0074401} /* (3, 13, 5) {real, imag} */,
  {32'h3f6935a5, 32'h40061f4c} /* (3, 13, 4) {real, imag} */,
  {32'hbe77af20, 32'hbda1dd58} /* (3, 13, 3) {real, imag} */,
  {32'h402fbbcf, 32'hbf9e735c} /* (3, 13, 2) {real, imag} */,
  {32'hbf1bb909, 32'hbf99834d} /* (3, 13, 1) {real, imag} */,
  {32'hbf5977df, 32'h3fbcf13b} /* (3, 13, 0) {real, imag} */,
  {32'hbc63d6f1, 32'h3f8ae325} /* (3, 12, 31) {real, imag} */,
  {32'h3ff9b196, 32'hbfa824c2} /* (3, 12, 30) {real, imag} */,
  {32'hbfe2ef4f, 32'hbf8351af} /* (3, 12, 29) {real, imag} */,
  {32'hbfa65484, 32'h3f6b65cc} /* (3, 12, 28) {real, imag} */,
  {32'hbfcddf7c, 32'hc0295be0} /* (3, 12, 27) {real, imag} */,
  {32'h3c8077d1, 32'h4039f8b7} /* (3, 12, 26) {real, imag} */,
  {32'h3e42de42, 32'hbf22ba8a} /* (3, 12, 25) {real, imag} */,
  {32'hc011dcbd, 32'hbfa999db} /* (3, 12, 24) {real, imag} */,
  {32'h3f29e8d7, 32'h3fb43cbe} /* (3, 12, 23) {real, imag} */,
  {32'hbf23c813, 32'h3f0e59ca} /* (3, 12, 22) {real, imag} */,
  {32'h3f5734dd, 32'h3fdf2ac9} /* (3, 12, 21) {real, imag} */,
  {32'h3fac99f8, 32'hbf4ecb9d} /* (3, 12, 20) {real, imag} */,
  {32'hbf06c8bb, 32'hc080263b} /* (3, 12, 19) {real, imag} */,
  {32'h3e7babab, 32'hbecfd3ec} /* (3, 12, 18) {real, imag} */,
  {32'h3fecb634, 32'h403d43e5} /* (3, 12, 17) {real, imag} */,
  {32'h3f751ed5, 32'hbfbf36ed} /* (3, 12, 16) {real, imag} */,
  {32'hbf827b91, 32'hbe3e616e} /* (3, 12, 15) {real, imag} */,
  {32'h3f80c4ad, 32'h3ae2bab3} /* (3, 12, 14) {real, imag} */,
  {32'h3e63cb5f, 32'h3fac2cbf} /* (3, 12, 13) {real, imag} */,
  {32'h3e7e2b02, 32'h409001c2} /* (3, 12, 12) {real, imag} */,
  {32'hbf244c9e, 32'h3fb00dcf} /* (3, 12, 11) {real, imag} */,
  {32'h3fb9e2ac, 32'hbf74d70d} /* (3, 12, 10) {real, imag} */,
  {32'h3e2e8886, 32'h3fd3bf81} /* (3, 12, 9) {real, imag} */,
  {32'hbfbc94ee, 32'hbfb1069e} /* (3, 12, 8) {real, imag} */,
  {32'h3f778bfe, 32'hc0178742} /* (3, 12, 7) {real, imag} */,
  {32'h3d944ea3, 32'h3d32f524} /* (3, 12, 6) {real, imag} */,
  {32'hc043de2d, 32'h3fe83c4d} /* (3, 12, 5) {real, imag} */,
  {32'h408a27cb, 32'h3e0d931a} /* (3, 12, 4) {real, imag} */,
  {32'h3dc080d8, 32'hbfef6603} /* (3, 12, 3) {real, imag} */,
  {32'h3f949b8d, 32'hbde5c5d7} /* (3, 12, 2) {real, imag} */,
  {32'h3ee9496f, 32'hc00bf4ed} /* (3, 12, 1) {real, imag} */,
  {32'h3e67fde9, 32'h3ec4bc0b} /* (3, 12, 0) {real, imag} */,
  {32'h4096aabb, 32'hbece73a9} /* (3, 11, 31) {real, imag} */,
  {32'hbffc5481, 32'h3fee7920} /* (3, 11, 30) {real, imag} */,
  {32'hbfeb2d86, 32'h404e5477} /* (3, 11, 29) {real, imag} */,
  {32'hbfc137d5, 32'hbf0a4870} /* (3, 11, 28) {real, imag} */,
  {32'hbf12a33a, 32'h3e66d25b} /* (3, 11, 27) {real, imag} */,
  {32'hc00bbac0, 32'hbf58fdda} /* (3, 11, 26) {real, imag} */,
  {32'hc08289e0, 32'h3f37cdb0} /* (3, 11, 25) {real, imag} */,
  {32'hbf17e641, 32'hc0480bab} /* (3, 11, 24) {real, imag} */,
  {32'hbe9edb48, 32'hbff62f2b} /* (3, 11, 23) {real, imag} */,
  {32'hbec7e146, 32'hc029aa4f} /* (3, 11, 22) {real, imag} */,
  {32'h408cbb0c, 32'h3f936635} /* (3, 11, 21) {real, imag} */,
  {32'h3f0f5f87, 32'h3f0eebf7} /* (3, 11, 20) {real, imag} */,
  {32'hbd91b779, 32'h3f940a93} /* (3, 11, 19) {real, imag} */,
  {32'h4033c2fe, 32'h40421c84} /* (3, 11, 18) {real, imag} */,
  {32'hbda4ca61, 32'hbe07e2a6} /* (3, 11, 17) {real, imag} */,
  {32'hbdd9e18c, 32'hbe0e9955} /* (3, 11, 16) {real, imag} */,
  {32'hbf7a69dc, 32'hbf420dba} /* (3, 11, 15) {real, imag} */,
  {32'h3eab5090, 32'hc00307e0} /* (3, 11, 14) {real, imag} */,
  {32'h3fe7faa7, 32'hc003b30d} /* (3, 11, 13) {real, imag} */,
  {32'hbf9a147e, 32'h3e006371} /* (3, 11, 12) {real, imag} */,
  {32'hc03e036c, 32'hbea95202} /* (3, 11, 11) {real, imag} */,
  {32'hc02b6683, 32'h4017f3aa} /* (3, 11, 10) {real, imag} */,
  {32'hbf5420a8, 32'hbf8a26e1} /* (3, 11, 9) {real, imag} */,
  {32'hbe447e93, 32'hbf9000ba} /* (3, 11, 8) {real, imag} */,
  {32'h40519300, 32'h3fb6ecf2} /* (3, 11, 7) {real, imag} */,
  {32'hbf64711c, 32'hc02ed046} /* (3, 11, 6) {real, imag} */,
  {32'hbe43a040, 32'h3f960ea0} /* (3, 11, 5) {real, imag} */,
  {32'h3f8231e7, 32'hc005576d} /* (3, 11, 4) {real, imag} */,
  {32'h3f907739, 32'hbf5a2d09} /* (3, 11, 3) {real, imag} */,
  {32'hc0829c46, 32'h3f5af039} /* (3, 11, 2) {real, imag} */,
  {32'h4077a877, 32'h3fc7e879} /* (3, 11, 1) {real, imag} */,
  {32'h3faec751, 32'hbf110f10} /* (3, 11, 0) {real, imag} */,
  {32'hbe0b72db, 32'h3f0df828} /* (3, 10, 31) {real, imag} */,
  {32'h4041e4bf, 32'h40381928} /* (3, 10, 30) {real, imag} */,
  {32'hbf9759b0, 32'h3f33d793} /* (3, 10, 29) {real, imag} */,
  {32'hbf39d105, 32'h3f5c28cd} /* (3, 10, 28) {real, imag} */,
  {32'h3f8a7ec3, 32'h3f852291} /* (3, 10, 27) {real, imag} */,
  {32'hbf3a619f, 32'hbe8bc337} /* (3, 10, 26) {real, imag} */,
  {32'h3eac2612, 32'hbd96c174} /* (3, 10, 25) {real, imag} */,
  {32'h40afa642, 32'h3ee22a6b} /* (3, 10, 24) {real, imag} */,
  {32'hbf945c1f, 32'hc0695d60} /* (3, 10, 23) {real, imag} */,
  {32'h4007c179, 32'hc026aedb} /* (3, 10, 22) {real, imag} */,
  {32'hc0556e64, 32'h40768a08} /* (3, 10, 21) {real, imag} */,
  {32'h3e8b8882, 32'h40818ec6} /* (3, 10, 20) {real, imag} */,
  {32'hbfc5b79a, 32'hbf9f00e1} /* (3, 10, 19) {real, imag} */,
  {32'h3ecce083, 32'h3ebd89ec} /* (3, 10, 18) {real, imag} */,
  {32'hbf8a868a, 32'hbf437d3f} /* (3, 10, 17) {real, imag} */,
  {32'h3f129543, 32'hbf64da3b} /* (3, 10, 16) {real, imag} */,
  {32'h3ff8d4bd, 32'h3f896060} /* (3, 10, 15) {real, imag} */,
  {32'hbf740269, 32'hbee35052} /* (3, 10, 14) {real, imag} */,
  {32'hbf2cb94a, 32'h404dd813} /* (3, 10, 13) {real, imag} */,
  {32'hc0108dca, 32'h3df0e7a6} /* (3, 10, 12) {real, imag} */,
  {32'hbd18f747, 32'hbf5270f4} /* (3, 10, 11) {real, imag} */,
  {32'hbfb4aed6, 32'hc01acd7b} /* (3, 10, 10) {real, imag} */,
  {32'h3f807290, 32'hbf2e9e8e} /* (3, 10, 9) {real, imag} */,
  {32'hc02481a5, 32'hbdeca734} /* (3, 10, 8) {real, imag} */,
  {32'h3f25c5c0, 32'hbfe5a3ae} /* (3, 10, 7) {real, imag} */,
  {32'h3fb749c1, 32'hc094dd39} /* (3, 10, 6) {real, imag} */,
  {32'h3f245149, 32'hc04ff351} /* (3, 10, 5) {real, imag} */,
  {32'h3d219c9a, 32'h3df66766} /* (3, 10, 4) {real, imag} */,
  {32'h40470e3c, 32'hbffb6932} /* (3, 10, 3) {real, imag} */,
  {32'h403af073, 32'h40137a86} /* (3, 10, 2) {real, imag} */,
  {32'hc0763e19, 32'h3f1fc4f5} /* (3, 10, 1) {real, imag} */,
  {32'hc01d8daa, 32'hc0dce454} /* (3, 10, 0) {real, imag} */,
  {32'hc00d905c, 32'hc087c143} /* (3, 9, 31) {real, imag} */,
  {32'h4040c6d4, 32'h3f4f3770} /* (3, 9, 30) {real, imag} */,
  {32'hc09e1285, 32'h3fc16734} /* (3, 9, 29) {real, imag} */,
  {32'h3fd97e89, 32'hc0b617ab} /* (3, 9, 28) {real, imag} */,
  {32'h404762b9, 32'hc03e6069} /* (3, 9, 27) {real, imag} */,
  {32'hbf91c9d5, 32'hc04ea6b2} /* (3, 9, 26) {real, imag} */,
  {32'hc00df3f1, 32'hbf0c6194} /* (3, 9, 25) {real, imag} */,
  {32'hbf1d90e8, 32'h3f3dbfb0} /* (3, 9, 24) {real, imag} */,
  {32'h3f87ea77, 32'hbfa5c48a} /* (3, 9, 23) {real, imag} */,
  {32'h3fbc68d5, 32'h3ff47aa6} /* (3, 9, 22) {real, imag} */,
  {32'hbfcc039c, 32'h4000eef6} /* (3, 9, 21) {real, imag} */,
  {32'h3f526379, 32'hc0221241} /* (3, 9, 20) {real, imag} */,
  {32'hbf9a3517, 32'hc08433a9} /* (3, 9, 19) {real, imag} */,
  {32'h3ff94224, 32'h3f46c065} /* (3, 9, 18) {real, imag} */,
  {32'hbf2f84fb, 32'hbd726d33} /* (3, 9, 17) {real, imag} */,
  {32'hbef68c41, 32'h3eeaa077} /* (3, 9, 16) {real, imag} */,
  {32'hbe928ee1, 32'h3eb68f9f} /* (3, 9, 15) {real, imag} */,
  {32'hbfda4ee0, 32'hbef2e015} /* (3, 9, 14) {real, imag} */,
  {32'hbfcbf6a4, 32'hbf8a4f78} /* (3, 9, 13) {real, imag} */,
  {32'h3f3a9bc0, 32'hbee4a463} /* (3, 9, 12) {real, imag} */,
  {32'h3fbd1c22, 32'h3efe1ad8} /* (3, 9, 11) {real, imag} */,
  {32'h3fe736ac, 32'h4029a599} /* (3, 9, 10) {real, imag} */,
  {32'h3ed8e5ad, 32'hbffdec9b} /* (3, 9, 9) {real, imag} */,
  {32'h3ee45f1b, 32'h3faa9888} /* (3, 9, 8) {real, imag} */,
  {32'h3fc1f29c, 32'hbf19495f} /* (3, 9, 7) {real, imag} */,
  {32'hbff98d5a, 32'hbfb336fd} /* (3, 9, 6) {real, imag} */,
  {32'hc0863403, 32'hbfb4941f} /* (3, 9, 5) {real, imag} */,
  {32'hbf379ba9, 32'h40032a00} /* (3, 9, 4) {real, imag} */,
  {32'h3f5575b1, 32'hbfdcc5c0} /* (3, 9, 3) {real, imag} */,
  {32'hc0043b2d, 32'hbf153de8} /* (3, 9, 2) {real, imag} */,
  {32'hbf39ddb7, 32'h40da730a} /* (3, 9, 1) {real, imag} */,
  {32'h3fce5bf5, 32'hbf9e872c} /* (3, 9, 0) {real, imag} */,
  {32'h407042a5, 32'hc0bcee6f} /* (3, 8, 31) {real, imag} */,
  {32'hbda6c9d5, 32'h40a9084a} /* (3, 8, 30) {real, imag} */,
  {32'hbfcf7554, 32'hbfc25c17} /* (3, 8, 29) {real, imag} */,
  {32'hbf5a648c, 32'h3f95de39} /* (3, 8, 28) {real, imag} */,
  {32'hbea48db3, 32'hbf1f061c} /* (3, 8, 27) {real, imag} */,
  {32'h4072f5cd, 32'hbf832d9a} /* (3, 8, 26) {real, imag} */,
  {32'h408f2518, 32'hc0020a47} /* (3, 8, 25) {real, imag} */,
  {32'h3fa92dbc, 32'hbf25fbaa} /* (3, 8, 24) {real, imag} */,
  {32'h3fb102fe, 32'h3cf84efa} /* (3, 8, 23) {real, imag} */,
  {32'hbe979af9, 32'h3fe478e7} /* (3, 8, 22) {real, imag} */,
  {32'hc01854f0, 32'hbfc5c7c6} /* (3, 8, 21) {real, imag} */,
  {32'hbec61305, 32'h3ecb3cf0} /* (3, 8, 20) {real, imag} */,
  {32'h3fefbdfa, 32'h3f3d6fc5} /* (3, 8, 19) {real, imag} */,
  {32'h3f4b61be, 32'hbf5892fb} /* (3, 8, 18) {real, imag} */,
  {32'h3e871995, 32'hbfdf8de8} /* (3, 8, 17) {real, imag} */,
  {32'hbf9199b0, 32'h3df53c33} /* (3, 8, 16) {real, imag} */,
  {32'h3e0a31e8, 32'hbf345b05} /* (3, 8, 15) {real, imag} */,
  {32'h3e496e5a, 32'hbf35f8dd} /* (3, 8, 14) {real, imag} */,
  {32'hbfe143a3, 32'h3e332f46} /* (3, 8, 13) {real, imag} */,
  {32'h3f916923, 32'hbfafee2d} /* (3, 8, 12) {real, imag} */,
  {32'hc09be87a, 32'hc06c9191} /* (3, 8, 11) {real, imag} */,
  {32'hbeaf0e6a, 32'h409ec0de} /* (3, 8, 10) {real, imag} */,
  {32'h3f7b1c18, 32'hc02a4d01} /* (3, 8, 9) {real, imag} */,
  {32'hc09623d0, 32'hbf775233} /* (3, 8, 8) {real, imag} */,
  {32'hc054d775, 32'hbee8c705} /* (3, 8, 7) {real, imag} */,
  {32'h3d7353f4, 32'h3fe13940} /* (3, 8, 6) {real, imag} */,
  {32'hbf2ebb89, 32'hc02e15c6} /* (3, 8, 5) {real, imag} */,
  {32'h3f9b0c69, 32'h408436d0} /* (3, 8, 4) {real, imag} */,
  {32'hc08efb8f, 32'hc03d6df5} /* (3, 8, 3) {real, imag} */,
  {32'hbf4a5e6e, 32'h405bd5ac} /* (3, 8, 2) {real, imag} */,
  {32'h408656ba, 32'hbeaaa2b5} /* (3, 8, 1) {real, imag} */,
  {32'h402d1bdd, 32'hc087f2e5} /* (3, 8, 0) {real, imag} */,
  {32'h3fd75b98, 32'hbfda3262} /* (3, 7, 31) {real, imag} */,
  {32'h3d8f0b8d, 32'hbde1614d} /* (3, 7, 30) {real, imag} */,
  {32'h3f840823, 32'h401138c7} /* (3, 7, 29) {real, imag} */,
  {32'h401bb393, 32'h404f664a} /* (3, 7, 28) {real, imag} */,
  {32'h3f17a4f5, 32'hbf93c984} /* (3, 7, 27) {real, imag} */,
  {32'h3f07a552, 32'h406d30f5} /* (3, 7, 26) {real, imag} */,
  {32'h3fd1cdc7, 32'hbf9a509d} /* (3, 7, 25) {real, imag} */,
  {32'hbfa6a23e, 32'h3f81f8de} /* (3, 7, 24) {real, imag} */,
  {32'h3e81c838, 32'hbfefcd7e} /* (3, 7, 23) {real, imag} */,
  {32'hbff4a5ff, 32'h3bc9904c} /* (3, 7, 22) {real, imag} */,
  {32'hc01714f8, 32'h3e723c75} /* (3, 7, 21) {real, imag} */,
  {32'hc026796d, 32'hbfcde374} /* (3, 7, 20) {real, imag} */,
  {32'h3f9f2459, 32'h4078ad53} /* (3, 7, 19) {real, imag} */,
  {32'h3f207332, 32'h403f1754} /* (3, 7, 18) {real, imag} */,
  {32'h3fe77170, 32'hbf7008dc} /* (3, 7, 17) {real, imag} */,
  {32'h3e6fb714, 32'h3f16de8e} /* (3, 7, 16) {real, imag} */,
  {32'h4001665c, 32'h3e00aacf} /* (3, 7, 15) {real, imag} */,
  {32'hc0080ea3, 32'h3efe3aca} /* (3, 7, 14) {real, imag} */,
  {32'h40079594, 32'hbf173295} /* (3, 7, 13) {real, imag} */,
  {32'h3f8d7aa6, 32'hbed1681e} /* (3, 7, 12) {real, imag} */,
  {32'hbf12d479, 32'h3f8f16c2} /* (3, 7, 11) {real, imag} */,
  {32'h40980f9c, 32'h3f89e9b3} /* (3, 7, 10) {real, imag} */,
  {32'hc02b0197, 32'hbcaec191} /* (3, 7, 9) {real, imag} */,
  {32'h3f1f4136, 32'hbf879f5b} /* (3, 7, 8) {real, imag} */,
  {32'hbfc72b43, 32'hbf867dbf} /* (3, 7, 7) {real, imag} */,
  {32'h3f45aaec, 32'h3f8842ac} /* (3, 7, 6) {real, imag} */,
  {32'h405e7499, 32'h402c37ef} /* (3, 7, 5) {real, imag} */,
  {32'hc07e78ad, 32'h405afbcf} /* (3, 7, 4) {real, imag} */,
  {32'h404dea96, 32'h3fbd2870} /* (3, 7, 3) {real, imag} */,
  {32'h4022ae4b, 32'hbfe65434} /* (3, 7, 2) {real, imag} */,
  {32'hbe8e2bbc, 32'h3fa5f9aa} /* (3, 7, 1) {real, imag} */,
  {32'h3f2151c2, 32'h40905de5} /* (3, 7, 0) {real, imag} */,
  {32'hc0544b3e, 32'hc03439f2} /* (3, 6, 31) {real, imag} */,
  {32'h3ff5cfb9, 32'hc04b9900} /* (3, 6, 30) {real, imag} */,
  {32'hbf499fb3, 32'hbee6bc7d} /* (3, 6, 29) {real, imag} */,
  {32'hbe49cc70, 32'hbf8d9687} /* (3, 6, 28) {real, imag} */,
  {32'h3f99d84c, 32'hc095512a} /* (3, 6, 27) {real, imag} */,
  {32'h40243e8d, 32'h40863a4d} /* (3, 6, 26) {real, imag} */,
  {32'hc0348af6, 32'hbfc0acd3} /* (3, 6, 25) {real, imag} */,
  {32'h3e29e194, 32'hbf1586cd} /* (3, 6, 24) {real, imag} */,
  {32'hbda36846, 32'h40d11e32} /* (3, 6, 23) {real, imag} */,
  {32'h3f0abd42, 32'hc05eeb20} /* (3, 6, 22) {real, imag} */,
  {32'h3f899e2c, 32'h3f8ebbc8} /* (3, 6, 21) {real, imag} */,
  {32'h4024d7d3, 32'hbf9a1cd0} /* (3, 6, 20) {real, imag} */,
  {32'h400cf67c, 32'h3f648ea2} /* (3, 6, 19) {real, imag} */,
  {32'hc02b2552, 32'h3f522f3f} /* (3, 6, 18) {real, imag} */,
  {32'h3f3a6790, 32'hbf90e7a5} /* (3, 6, 17) {real, imag} */,
  {32'hbfb1ced6, 32'hbf502797} /* (3, 6, 16) {real, imag} */,
  {32'hbf368527, 32'hbfcd4995} /* (3, 6, 15) {real, imag} */,
  {32'h3f1bf115, 32'hbe365f7d} /* (3, 6, 14) {real, imag} */,
  {32'hbf9b96e4, 32'h3ef45485} /* (3, 6, 13) {real, imag} */,
  {32'hc056c37d, 32'h3f8de583} /* (3, 6, 12) {real, imag} */,
  {32'hbf894c35, 32'h3f80bf34} /* (3, 6, 11) {real, imag} */,
  {32'hbf417089, 32'hbfb04aae} /* (3, 6, 10) {real, imag} */,
  {32'hbf63524f, 32'hbe45e47a} /* (3, 6, 9) {real, imag} */,
  {32'h3f9de225, 32'hc00cd59b} /* (3, 6, 8) {real, imag} */,
  {32'hc0f4274b, 32'h408b2ab0} /* (3, 6, 7) {real, imag} */,
  {32'hc024436a, 32'h3f7c6631} /* (3, 6, 6) {real, imag} */,
  {32'hc000b00f, 32'hbe4e020f} /* (3, 6, 5) {real, imag} */,
  {32'hbf99900a, 32'h3ef7e6b0} /* (3, 6, 4) {real, imag} */,
  {32'h40497701, 32'hbf894c1d} /* (3, 6, 3) {real, imag} */,
  {32'h3feb47b3, 32'hc0d209da} /* (3, 6, 2) {real, imag} */,
  {32'hbe3b6f49, 32'hc0b73fb9} /* (3, 6, 1) {real, imag} */,
  {32'h3fedd97d, 32'h406ec828} /* (3, 6, 0) {real, imag} */,
  {32'h40cf63af, 32'hc1b550d2} /* (3, 5, 31) {real, imag} */,
  {32'hc05ba367, 32'h41290779} /* (3, 5, 30) {real, imag} */,
  {32'hbf224813, 32'h40ac12f7} /* (3, 5, 29) {real, imag} */,
  {32'h3f2f2677, 32'hc00f3bb8} /* (3, 5, 28) {real, imag} */,
  {32'hbfc373a5, 32'h40dec2c2} /* (3, 5, 27) {real, imag} */,
  {32'hc04ee3ed, 32'hbfc699b2} /* (3, 5, 26) {real, imag} */,
  {32'hc0af9a51, 32'hbff4604d} /* (3, 5, 25) {real, imag} */,
  {32'h406540c7, 32'hc029490a} /* (3, 5, 24) {real, imag} */,
  {32'h3fc33f49, 32'hbf81d43a} /* (3, 5, 23) {real, imag} */,
  {32'hbfc9a999, 32'hbe614d9c} /* (3, 5, 22) {real, imag} */,
  {32'h3fcc7169, 32'h3fd27998} /* (3, 5, 21) {real, imag} */,
  {32'h3fd6e36a, 32'hbf3d41fd} /* (3, 5, 20) {real, imag} */,
  {32'h40413538, 32'hbe9df0c6} /* (3, 5, 19) {real, imag} */,
  {32'hbfbdf442, 32'h3f995e5f} /* (3, 5, 18) {real, imag} */,
  {32'hbd4551f2, 32'h3f855491} /* (3, 5, 17) {real, imag} */,
  {32'hbf4077c7, 32'h401105e6} /* (3, 5, 16) {real, imag} */,
  {32'hbf078f01, 32'h3eceb292} /* (3, 5, 15) {real, imag} */,
  {32'hc012ba9f, 32'hbe3a3257} /* (3, 5, 14) {real, imag} */,
  {32'h3e8bdf78, 32'hbe093580} /* (3, 5, 13) {real, imag} */,
  {32'h3fa898e7, 32'h401745fc} /* (3, 5, 12) {real, imag} */,
  {32'h3ebda071, 32'hc018e76f} /* (3, 5, 11) {real, imag} */,
  {32'hc012e072, 32'h401b205e} /* (3, 5, 10) {real, imag} */,
  {32'h4027f69c, 32'h3ff97103} /* (3, 5, 9) {real, imag} */,
  {32'hbf9fa26f, 32'h400d12f9} /* (3, 5, 8) {real, imag} */,
  {32'h408b521f, 32'h3eefd78e} /* (3, 5, 7) {real, imag} */,
  {32'h3fc0ca1f, 32'h402f167c} /* (3, 5, 6) {real, imag} */,
  {32'hc0d57fcd, 32'hc086c11d} /* (3, 5, 5) {real, imag} */,
  {32'hbf849c7c, 32'hbfa770f0} /* (3, 5, 4) {real, imag} */,
  {32'hc0818064, 32'hbf64a0f2} /* (3, 5, 3) {real, imag} */,
  {32'hbfb6d6cb, 32'h40ea0352} /* (3, 5, 2) {real, imag} */,
  {32'h41a2e425, 32'hc10092fa} /* (3, 5, 1) {real, imag} */,
  {32'h40e0630f, 32'hc13cbcad} /* (3, 5, 0) {real, imag} */,
  {32'hc18c773f, 32'h4125908f} /* (3, 4, 31) {real, imag} */,
  {32'h415e52e1, 32'hc1308ece} /* (3, 4, 30) {real, imag} */,
  {32'hc098c676, 32'h3fd71129} /* (3, 4, 29) {real, imag} */,
  {32'hbd57e5e4, 32'h40aa5fc9} /* (3, 4, 28) {real, imag} */,
  {32'h3e98ca41, 32'hc0e00290} /* (3, 4, 27) {real, imag} */,
  {32'hbfaeadc4, 32'hc088e21a} /* (3, 4, 26) {real, imag} */,
  {32'h402e92fa, 32'hbfd45ca4} /* (3, 4, 25) {real, imag} */,
  {32'h400b8e5d, 32'hbf11cf15} /* (3, 4, 24) {real, imag} */,
  {32'hbdf4fc27, 32'hbfc6245d} /* (3, 4, 23) {real, imag} */,
  {32'hbfc9cf76, 32'h400c2427} /* (3, 4, 22) {real, imag} */,
  {32'hbf717df2, 32'hc003cf8a} /* (3, 4, 21) {real, imag} */,
  {32'h3f87c16d, 32'h3fb85295} /* (3, 4, 20) {real, imag} */,
  {32'h3e5eeefc, 32'h3f3b27fa} /* (3, 4, 19) {real, imag} */,
  {32'h3f0e5ad8, 32'hbf4d64ed} /* (3, 4, 18) {real, imag} */,
  {32'h3f41a6c4, 32'h3f669b9f} /* (3, 4, 17) {real, imag} */,
  {32'h3e1d6b4e, 32'h3d9cf8ce} /* (3, 4, 16) {real, imag} */,
  {32'h3f1b672b, 32'hc01ba190} /* (3, 4, 15) {real, imag} */,
  {32'h40050d63, 32'hbfaa71fb} /* (3, 4, 14) {real, imag} */,
  {32'h3f1e239e, 32'hbee2b1df} /* (3, 4, 13) {real, imag} */,
  {32'hbd17ee89, 32'hbf8463df} /* (3, 4, 12) {real, imag} */,
  {32'h400c31b2, 32'h3fb0f8f9} /* (3, 4, 11) {real, imag} */,
  {32'hc047901e, 32'h3f639236} /* (3, 4, 10) {real, imag} */,
  {32'h4038f582, 32'hbf09a6ff} /* (3, 4, 9) {real, imag} */,
  {32'h403b200c, 32'hc05720fb} /* (3, 4, 8) {real, imag} */,
  {32'h405a0273, 32'hbd3c5b72} /* (3, 4, 7) {real, imag} */,
  {32'hbdf96e97, 32'h402e5f4d} /* (3, 4, 6) {real, imag} */,
  {32'h40cfad1b, 32'hbfc22649} /* (3, 4, 5) {real, imag} */,
  {32'hc11c79da, 32'h40b4e4e0} /* (3, 4, 4) {real, imag} */,
  {32'h40cbbe5d, 32'hc05685f9} /* (3, 4, 3) {real, imag} */,
  {32'h419e7eed, 32'hc108a5d4} /* (3, 4, 2) {real, imag} */,
  {32'hc16327ba, 32'h418e6c47} /* (3, 4, 1) {real, imag} */,
  {32'hc08fda18, 32'h41bf6cb2} /* (3, 4, 0) {real, imag} */,
  {32'hc08c98ce, 32'hc1b50186} /* (3, 3, 31) {real, imag} */,
  {32'h3f9367d1, 32'h412c782d} /* (3, 3, 30) {real, imag} */,
  {32'hbeaf6fb8, 32'hbed57494} /* (3, 3, 29) {real, imag} */,
  {32'hc0900e9d, 32'h3eaceec9} /* (3, 3, 28) {real, imag} */,
  {32'h405402ad, 32'hc00d712c} /* (3, 3, 27) {real, imag} */,
  {32'h40bd73a7, 32'h3cb8ac42} /* (3, 3, 26) {real, imag} */,
  {32'hc018a876, 32'hc0dbf8b8} /* (3, 3, 25) {real, imag} */,
  {32'h4124b160, 32'h3fe6d2ea} /* (3, 3, 24) {real, imag} */,
  {32'hc0874862, 32'h3f309b80} /* (3, 3, 23) {real, imag} */,
  {32'hbfc6dcc2, 32'hc01b7a6c} /* (3, 3, 22) {real, imag} */,
  {32'h3e83226d, 32'hbe5b57ca} /* (3, 3, 21) {real, imag} */,
  {32'h3f978cfa, 32'h3f26c8b3} /* (3, 3, 20) {real, imag} */,
  {32'hc0997ba9, 32'h3f4cafc6} /* (3, 3, 19) {real, imag} */,
  {32'h4017f213, 32'h3f846594} /* (3, 3, 18) {real, imag} */,
  {32'h40067646, 32'h3f8dbb0a} /* (3, 3, 17) {real, imag} */,
  {32'h3ff78287, 32'hbfb2d139} /* (3, 3, 16) {real, imag} */,
  {32'hbfd4efd5, 32'hbf40fcbe} /* (3, 3, 15) {real, imag} */,
  {32'h3ef6bd0a, 32'hbfb405c4} /* (3, 3, 14) {real, imag} */,
  {32'h3f66ab3b, 32'h3fccf8bc} /* (3, 3, 13) {real, imag} */,
  {32'h401b7461, 32'h40219d5d} /* (3, 3, 12) {real, imag} */,
  {32'h3e49adc0, 32'h3ffb1ec5} /* (3, 3, 11) {real, imag} */,
  {32'h400b7aaf, 32'h3fd4571a} /* (3, 3, 10) {real, imag} */,
  {32'hc086b745, 32'hbe8ef1ab} /* (3, 3, 9) {real, imag} */,
  {32'h3ef1d2cc, 32'h402680b9} /* (3, 3, 8) {real, imag} */,
  {32'hc07f4c49, 32'hc020f3c7} /* (3, 3, 7) {real, imag} */,
  {32'h4097c6df, 32'h401c03b8} /* (3, 3, 6) {real, imag} */,
  {32'hc02a8370, 32'h40c94701} /* (3, 3, 5) {real, imag} */,
  {32'hc08dd30f, 32'hc15fc88b} /* (3, 3, 4) {real, imag} */,
  {32'hbffe0a78, 32'h41013dbd} /* (3, 3, 3) {real, imag} */,
  {32'h4152d32d, 32'h414c7491} /* (3, 3, 2) {real, imag} */,
  {32'hc1672ddb, 32'h40348f70} /* (3, 3, 1) {real, imag} */,
  {32'hc05308e2, 32'hc168914e} /* (3, 3, 0) {real, imag} */,
  {32'h42350981, 32'hc2fa7b46} /* (3, 2, 31) {real, imag} */,
  {32'hc122bd67, 32'h4285d676} /* (3, 2, 30) {real, imag} */,
  {32'h3f2497ba, 32'hc0ffd906} /* (3, 2, 29) {real, imag} */,
  {32'hc13f49f0, 32'hc09d3dd2} /* (3, 2, 28) {real, imag} */,
  {32'h40b3d60d, 32'h411e1b0e} /* (3, 2, 27) {real, imag} */,
  {32'h3fe8e697, 32'h3ff13430} /* (3, 2, 26) {real, imag} */,
  {32'h3eb6a0e3, 32'h3e167ddd} /* (3, 2, 25) {real, imag} */,
  {32'h3ff86345, 32'h40ba86e4} /* (3, 2, 24) {real, imag} */,
  {32'hc00d2dab, 32'h3fff3ef1} /* (3, 2, 23) {real, imag} */,
  {32'hc0ae287e, 32'hbf3287fb} /* (3, 2, 22) {real, imag} */,
  {32'h402646cc, 32'hc023e261} /* (3, 2, 21) {real, imag} */,
  {32'hbf70da12, 32'h40154323} /* (3, 2, 20) {real, imag} */,
  {32'h40139edf, 32'h3f484c37} /* (3, 2, 19) {real, imag} */,
  {32'h3eeeddca, 32'hbf0555ec} /* (3, 2, 18) {real, imag} */,
  {32'hbfa64b0d, 32'hbe9da80f} /* (3, 2, 17) {real, imag} */,
  {32'h3d0b7e42, 32'h3fb3f94a} /* (3, 2, 16) {real, imag} */,
  {32'hbd9e4d98, 32'hbfc6489a} /* (3, 2, 15) {real, imag} */,
  {32'hbdfbab29, 32'hbf637d52} /* (3, 2, 14) {real, imag} */,
  {32'hbe1a92ea, 32'h3f26b3a5} /* (3, 2, 13) {real, imag} */,
  {32'h401b2741, 32'hbff88e6f} /* (3, 2, 12) {real, imag} */,
  {32'hbfdeb1e8, 32'h3f332e49} /* (3, 2, 11) {real, imag} */,
  {32'h401a2f6b, 32'hc01010a1} /* (3, 2, 10) {real, imag} */,
  {32'hc0261f69, 32'h3f82e819} /* (3, 2, 9) {real, imag} */,
  {32'hbe725135, 32'hbd92f1a9} /* (3, 2, 8) {real, imag} */,
  {32'h4061550d, 32'hbfe4fa8b} /* (3, 2, 7) {real, imag} */,
  {32'h3f2677fd, 32'hbfaa731c} /* (3, 2, 6) {real, imag} */,
  {32'hc0978e0e, 32'h41031486} /* (3, 2, 5) {real, imag} */,
  {32'h410ddbb4, 32'hc0ed8c99} /* (3, 2, 4) {real, imag} */,
  {32'hc09c3ece, 32'hc0a52078} /* (3, 2, 3) {real, imag} */,
  {32'hbf461e4e, 32'h4237bc33} /* (3, 2, 2) {real, imag} */,
  {32'h3e0edecd, 32'hc2797067} /* (3, 2, 1) {real, imag} */,
  {32'h41eb9fff, 32'hc22de765} /* (3, 2, 0) {real, imag} */,
  {32'hc156cbdc, 32'h4309411e} /* (3, 1, 31) {real, imag} */,
  {32'h41a54c6d, 32'hc1ea1b89} /* (3, 1, 30) {real, imag} */,
  {32'hc09296ea, 32'hc18fe05d} /* (3, 1, 29) {real, imag} */,
  {32'hc17a3ebd, 32'h417a5bdf} /* (3, 1, 28) {real, imag} */,
  {32'h40eaa911, 32'hc1a48fdb} /* (3, 1, 27) {real, imag} */,
  {32'hbfb12724, 32'hc05b4a53} /* (3, 1, 26) {real, imag} */,
  {32'h40eed908, 32'h3ff1df49} /* (3, 1, 25) {real, imag} */,
  {32'hc0489e6d, 32'hc0bc6647} /* (3, 1, 24) {real, imag} */,
  {32'h3fa8c932, 32'hbf75c066} /* (3, 1, 23) {real, imag} */,
  {32'h40029cc3, 32'h40245fd5} /* (3, 1, 22) {real, imag} */,
  {32'hbefa3260, 32'hc077ab16} /* (3, 1, 21) {real, imag} */,
  {32'hc00139ae, 32'h4004f27e} /* (3, 1, 20) {real, imag} */,
  {32'hc0054d15, 32'h3eddf50e} /* (3, 1, 19) {real, imag} */,
  {32'hc03cb5ad, 32'hbe6c8d9a} /* (3, 1, 18) {real, imag} */,
  {32'hbf3c2eb6, 32'hbfb3cac4} /* (3, 1, 17) {real, imag} */,
  {32'h3fc807aa, 32'h3f869e0c} /* (3, 1, 16) {real, imag} */,
  {32'hbe779aa0, 32'hbfa174b7} /* (3, 1, 15) {real, imag} */,
  {32'h3fac38ab, 32'h40214903} /* (3, 1, 14) {real, imag} */,
  {32'hc090fd2b, 32'hbfb65adf} /* (3, 1, 13) {real, imag} */,
  {32'h3fa44955, 32'h3fb4bb7b} /* (3, 1, 12) {real, imag} */,
  {32'h40a92429, 32'hbf813282} /* (3, 1, 11) {real, imag} */,
  {32'hbfcb5f66, 32'hc0aabdd2} /* (3, 1, 10) {real, imag} */,
  {32'h40a6e3db, 32'h3f186961} /* (3, 1, 9) {real, imag} */,
  {32'h40c1d97f, 32'hbf086677} /* (3, 1, 8) {real, imag} */,
  {32'hc05c90f7, 32'hc0c03355} /* (3, 1, 7) {real, imag} */,
  {32'hc0bfab25, 32'hc087bef7} /* (3, 1, 6) {real, imag} */,
  {32'h410bd82b, 32'hc15ef585} /* (3, 1, 5) {real, imag} */,
  {32'h3fb9c2f0, 32'h4112524c} /* (3, 1, 4) {real, imag} */,
  {32'h4193d282, 32'h410acee1} /* (3, 1, 3) {real, imag} */,
  {32'h428de949, 32'hc236a51c} /* (3, 1, 2) {real, imag} */,
  {32'hc305191c, 32'h4312a991} /* (3, 1, 1) {real, imag} */,
  {32'hc239a83e, 32'h42edf486} /* (3, 1, 0) {real, imag} */,
  {32'h4269be17, 32'h42acb596} /* (3, 0, 31) {real, imag} */,
  {32'hc1b61ee2, 32'hc1b35bfc} /* (3, 0, 30) {real, imag} */,
  {32'hc16924d5, 32'hc00e3985} /* (3, 0, 29) {real, imag} */,
  {32'hc17286fd, 32'hbf8b7f3e} /* (3, 0, 28) {real, imag} */,
  {32'h4092e3ce, 32'hc14aeba8} /* (3, 0, 27) {real, imag} */,
  {32'hc08cb2df, 32'hc027c2ac} /* (3, 0, 26) {real, imag} */,
  {32'h4085c387, 32'h402ef542} /* (3, 0, 25) {real, imag} */,
  {32'hc08369a4, 32'h401527fe} /* (3, 0, 24) {real, imag} */,
  {32'h3f60c307, 32'h404d9cd9} /* (3, 0, 23) {real, imag} */,
  {32'h3fadff49, 32'h40196d95} /* (3, 0, 22) {real, imag} */,
  {32'hbeb31e99, 32'hc01efc6a} /* (3, 0, 21) {real, imag} */,
  {32'h3ff2d6c4, 32'h40179a91} /* (3, 0, 20) {real, imag} */,
  {32'hbe83853f, 32'hbf41b6b2} /* (3, 0, 19) {real, imag} */,
  {32'h3e9bce9e, 32'hbff4208b} /* (3, 0, 18) {real, imag} */,
  {32'hbf10ad08, 32'hbfa08fc0} /* (3, 0, 17) {real, imag} */,
  {32'hbecafaff, 32'hbfad3113} /* (3, 0, 16) {real, imag} */,
  {32'hbfd09e88, 32'h3f0cadb8} /* (3, 0, 15) {real, imag} */,
  {32'h3fdf6a58, 32'h40585fcc} /* (3, 0, 14) {real, imag} */,
  {32'hbf27a437, 32'h404c0374} /* (3, 0, 13) {real, imag} */,
  {32'hc0831a9d, 32'h3e2dfe7c} /* (3, 0, 12) {real, imag} */,
  {32'h4014b00d, 32'h3f8f131d} /* (3, 0, 11) {real, imag} */,
  {32'h40960c17, 32'h4036364e} /* (3, 0, 10) {real, imag} */,
  {32'h3f6ef582, 32'hbfc5057f} /* (3, 0, 9) {real, imag} */,
  {32'h408531ba, 32'hbf826c82} /* (3, 0, 8) {real, imag} */,
  {32'hc0c2bbe2, 32'hc0db86dd} /* (3, 0, 7) {real, imag} */,
  {32'hc10fe016, 32'h401d2c13} /* (3, 0, 6) {real, imag} */,
  {32'h416a7091, 32'hc133b17c} /* (3, 0, 5) {real, imag} */,
  {32'h412f7f39, 32'hbff187ea} /* (3, 0, 4) {real, imag} */,
  {32'hc131d470, 32'hc1984692} /* (3, 0, 3) {real, imag} */,
  {32'h41a48bbe, 32'hc0572dd9} /* (3, 0, 2) {real, imag} */,
  {32'hc28e7e07, 32'h4289abac} /* (3, 0, 1) {real, imag} */,
  {32'hc1f2f479, 32'h42797e12} /* (3, 0, 0) {real, imag} */,
  {32'h43750664, 32'h444999dc} /* (2, 31, 31) {real, imag} */,
  {32'hc32b295f, 32'hc383799c} /* (2, 31, 30) {real, imag} */,
  {32'h408f793e, 32'hc1b34366} /* (2, 31, 29) {real, imag} */,
  {32'h4184de41, 32'h40132bcb} /* (2, 31, 28) {real, imag} */,
  {32'hc11c1686, 32'hc200ba84} /* (2, 31, 27) {real, imag} */,
  {32'h3f136497, 32'hc03b6f8e} /* (2, 31, 26) {real, imag} */,
  {32'h40d2f533, 32'h40ab4cf5} /* (2, 31, 25) {real, imag} */,
  {32'hc17bcab0, 32'hc12bbe0e} /* (2, 31, 24) {real, imag} */,
  {32'hbfc18ac4, 32'hbf2e0329} /* (2, 31, 23) {real, imag} */,
  {32'h3fa39e56, 32'hc08111d6} /* (2, 31, 22) {real, imag} */,
  {32'hc0812554, 32'hc0ad2f43} /* (2, 31, 21) {real, imag} */,
  {32'hbefb618f, 32'h3fd6b4cd} /* (2, 31, 20) {real, imag} */,
  {32'h3f18767d, 32'h3fab01c8} /* (2, 31, 19) {real, imag} */,
  {32'hc0a2af1c, 32'h3fe25a27} /* (2, 31, 18) {real, imag} */,
  {32'h4016b34f, 32'hbf9f0ffb} /* (2, 31, 17) {real, imag} */,
  {32'h3f04ee2a, 32'h3f65538a} /* (2, 31, 16) {real, imag} */,
  {32'hbd1fdad1, 32'hbea4843d} /* (2, 31, 15) {real, imag} */,
  {32'h40915d2f, 32'h3f826d14} /* (2, 31, 14) {real, imag} */,
  {32'h3dfb848c, 32'hc05320f9} /* (2, 31, 13) {real, imag} */,
  {32'hbf024f6d, 32'hbf1a84bd} /* (2, 31, 12) {real, imag} */,
  {32'h411efae8, 32'hc0b5b8a4} /* (2, 31, 11) {real, imag} */,
  {32'h3f098a48, 32'h3eb21c95} /* (2, 31, 10) {real, imag} */,
  {32'hbee60919, 32'hc067ab3a} /* (2, 31, 9) {real, imag} */,
  {32'h4127ee15, 32'hc0afc6a7} /* (2, 31, 8) {real, imag} */,
  {32'hc0a5e6b7, 32'h4093b168} /* (2, 31, 7) {real, imag} */,
  {32'h41409e32, 32'hc0be798d} /* (2, 31, 6) {real, imag} */,
  {32'h41823857, 32'hc2740455} /* (2, 31, 5) {real, imag} */,
  {32'h41c155f6, 32'h424df572} /* (2, 31, 4) {real, imag} */,
  {32'h41356100, 32'hc1a7a084} /* (2, 31, 3) {real, imag} */,
  {32'h41cb8a6c, 32'hc307b885} /* (2, 31, 2) {real, imag} */,
  {32'hc363a405, 32'h43ffa953} /* (2, 31, 1) {real, imag} */,
  {32'hc2afa8fc, 32'h441443e2} /* (2, 31, 0) {real, imag} */,
  {32'h42b31a1f, 32'hc373a611} /* (2, 30, 31) {real, imag} */,
  {32'hc2c3eebb, 32'h430de680} /* (2, 30, 30) {real, imag} */,
  {32'h40588da8, 32'h4048bf4e} /* (2, 30, 29) {real, imag} */,
  {32'h406a5d3b, 32'hc218f3d9} /* (2, 30, 28) {real, imag} */,
  {32'h41e1e526, 32'h41e8055c} /* (2, 30, 27) {real, imag} */,
  {32'h3cea1769, 32'hc086813e} /* (2, 30, 26) {real, imag} */,
  {32'h400b45ac, 32'hc069f3c3} /* (2, 30, 25) {real, imag} */,
  {32'h41054c07, 32'h4163ceec} /* (2, 30, 24) {real, imag} */,
  {32'hc0361ebd, 32'hbfdad88c} /* (2, 30, 23) {real, imag} */,
  {32'hc056f322, 32'hc0ac9f26} /* (2, 30, 22) {real, imag} */,
  {32'h40c2724c, 32'h403d34a1} /* (2, 30, 21) {real, imag} */,
  {32'h3e5a3e1b, 32'hbfc3c554} /* (2, 30, 20) {real, imag} */,
  {32'hbee2b415, 32'hbf8e3691} /* (2, 30, 19) {real, imag} */,
  {32'h40ae8274, 32'h3fd6e77e} /* (2, 30, 18) {real, imag} */,
  {32'hbf6e0795, 32'hbfdc31f2} /* (2, 30, 17) {real, imag} */,
  {32'h3fa4594b, 32'h40082653} /* (2, 30, 16) {real, imag} */,
  {32'h4088cfe2, 32'h3efa9d54} /* (2, 30, 15) {real, imag} */,
  {32'hc040907e, 32'h400c3f86} /* (2, 30, 14) {real, imag} */,
  {32'hbd67eb86, 32'h3f392de4} /* (2, 30, 13) {real, imag} */,
  {32'hbea260df, 32'hc075d5ec} /* (2, 30, 12) {real, imag} */,
  {32'hc1194fd8, 32'h3f5c6638} /* (2, 30, 11) {real, imag} */,
  {32'h40046152, 32'h3e7d2a0e} /* (2, 30, 10) {real, imag} */,
  {32'hbf5f8718, 32'h4009e7fb} /* (2, 30, 9) {real, imag} */,
  {32'hc1b859c7, 32'h412fa83a} /* (2, 30, 8) {real, imag} */,
  {32'h413d7688, 32'hc0001b9d} /* (2, 30, 7) {real, imag} */,
  {32'hc02f33ca, 32'h40a7683c} /* (2, 30, 6) {real, imag} */,
  {32'hc1cb41b3, 32'h41581812} /* (2, 30, 5) {real, imag} */,
  {32'h42170128, 32'hc1905b99} /* (2, 30, 4) {real, imag} */,
  {32'h410f371c, 32'hbfebe84c} /* (2, 30, 3) {real, imag} */,
  {32'hc2f4b5f1, 32'h4359f467} /* (2, 30, 2) {real, imag} */,
  {32'h42b01dd2, 32'hc3ddbab4} /* (2, 30, 1) {real, imag} */,
  {32'h40e32513, 32'hc37acf45} /* (2, 30, 0) {real, imag} */,
  {32'h420f5519, 32'h428b2aea} /* (2, 29, 31) {real, imag} */,
  {32'hc24dc073, 32'hc14ebf45} /* (2, 29, 30) {real, imag} */,
  {32'h415fa31a, 32'h4097a24d} /* (2, 29, 29) {real, imag} */,
  {32'h413d366f, 32'hc198c15d} /* (2, 29, 28) {real, imag} */,
  {32'h3f16ca90, 32'hc026b9c5} /* (2, 29, 27) {real, imag} */,
  {32'h401c68de, 32'hbe548867} /* (2, 29, 26) {real, imag} */,
  {32'h40b2bb25, 32'h402a185c} /* (2, 29, 25) {real, imag} */,
  {32'hbebe3edd, 32'h40880148} /* (2, 29, 24) {real, imag} */,
  {32'h3ed00f30, 32'h3e83ec3c} /* (2, 29, 23) {real, imag} */,
  {32'h3f0e56ae, 32'hbe71b180} /* (2, 29, 22) {real, imag} */,
  {32'h3fd3017f, 32'h40280b06} /* (2, 29, 21) {real, imag} */,
  {32'hbf51984e, 32'hc00f0d6e} /* (2, 29, 20) {real, imag} */,
  {32'hbf811ef4, 32'h3e9f15a9} /* (2, 29, 19) {real, imag} */,
  {32'hc01fe22e, 32'hbf9e4649} /* (2, 29, 18) {real, imag} */,
  {32'h3eee5477, 32'h3fccc76a} /* (2, 29, 17) {real, imag} */,
  {32'hbf7850ed, 32'hbd733db1} /* (2, 29, 16) {real, imag} */,
  {32'h3f0f198c, 32'h3ec7404d} /* (2, 29, 15) {real, imag} */,
  {32'hc010b8a6, 32'h3f84f826} /* (2, 29, 14) {real, imag} */,
  {32'hc08e5650, 32'hbf91cf40} /* (2, 29, 13) {real, imag} */,
  {32'hbfbbaf96, 32'hc03f77c3} /* (2, 29, 12) {real, imag} */,
  {32'hbe7d8f60, 32'hbd64b515} /* (2, 29, 11) {real, imag} */,
  {32'h40b0f982, 32'h3ff7436a} /* (2, 29, 10) {real, imag} */,
  {32'h3ff02b19, 32'h3e488e19} /* (2, 29, 9) {real, imag} */,
  {32'hc0d38e5a, 32'hc08d7dfe} /* (2, 29, 8) {real, imag} */,
  {32'hbd82f28d, 32'h3f968ceb} /* (2, 29, 7) {real, imag} */,
  {32'h4090069a, 32'h40891573} /* (2, 29, 6) {real, imag} */,
  {32'h408a97f6, 32'hc0dc955f} /* (2, 29, 5) {real, imag} */,
  {32'h4102690d, 32'h41558dd1} /* (2, 29, 4) {real, imag} */,
  {32'h3fd87d79, 32'h405f7f8b} /* (2, 29, 3) {real, imag} */,
  {32'hc24c371c, 32'h414b8448} /* (2, 29, 2) {real, imag} */,
  {32'h425b74d8, 32'hc2638df0} /* (2, 29, 1) {real, imag} */,
  {32'hc130fc6f, 32'hbfb71427} /* (2, 29, 0) {real, imag} */,
  {32'h4175143c, 32'h42a5023a} /* (2, 28, 31) {real, imag} */,
  {32'hc1dfbd95, 32'hc24e6be5} /* (2, 28, 30) {real, imag} */,
  {32'h404ed4f1, 32'h403bda0a} /* (2, 28, 29) {real, imag} */,
  {32'h3f828e05, 32'hc0566f0e} /* (2, 28, 28) {real, imag} */,
  {32'hc1498394, 32'hc0347a7c} /* (2, 28, 27) {real, imag} */,
  {32'h3f0c4fe9, 32'hbf966e0c} /* (2, 28, 26) {real, imag} */,
  {32'h401474ef, 32'h4051069c} /* (2, 28, 25) {real, imag} */,
  {32'hc0899c17, 32'hc0baa25c} /* (2, 28, 24) {real, imag} */,
  {32'h4011c8dc, 32'hbfaba89a} /* (2, 28, 23) {real, imag} */,
  {32'h40a54489, 32'hbffc9286} /* (2, 28, 22) {real, imag} */,
  {32'hbfbb2b8e, 32'h3f137266} /* (2, 28, 21) {real, imag} */,
  {32'h3ee5f52b, 32'h3fe99149} /* (2, 28, 20) {real, imag} */,
  {32'h3eb27d7d, 32'hbe1a6413} /* (2, 28, 19) {real, imag} */,
  {32'hc079075d, 32'hbfb7d87d} /* (2, 28, 18) {real, imag} */,
  {32'h402cc952, 32'hbf6760dc} /* (2, 28, 17) {real, imag} */,
  {32'hbe6985b0, 32'h3fbcbfad} /* (2, 28, 16) {real, imag} */,
  {32'hbf166b92, 32'h400cfca8} /* (2, 28, 15) {real, imag} */,
  {32'hbdb29236, 32'hc06b5298} /* (2, 28, 14) {real, imag} */,
  {32'hbf14a898, 32'h3f43133f} /* (2, 28, 13) {real, imag} */,
  {32'hc08f4a4b, 32'h40598d7b} /* (2, 28, 12) {real, imag} */,
  {32'h40838147, 32'hc0a21e4c} /* (2, 28, 11) {real, imag} */,
  {32'hbfc0efa1, 32'h3f114708} /* (2, 28, 10) {real, imag} */,
  {32'hc0969cb8, 32'h3ff274a8} /* (2, 28, 9) {real, imag} */,
  {32'hbfc32460, 32'hc000d33f} /* (2, 28, 8) {real, imag} */,
  {32'hbffd56c5, 32'hbe103e98} /* (2, 28, 7) {real, imag} */,
  {32'h40c46e43, 32'h3fa9b31c} /* (2, 28, 6) {real, imag} */,
  {32'h40850ebc, 32'hc14b986a} /* (2, 28, 5) {real, imag} */,
  {32'h40011c6a, 32'h41370ca3} /* (2, 28, 4) {real, imag} */,
  {32'hbf980553, 32'hbfd32861} /* (2, 28, 3) {real, imag} */,
  {32'hc1ffefef, 32'hc225b0ce} /* (2, 28, 2) {real, imag} */,
  {32'h42275d2f, 32'h4209eaa5} /* (2, 28, 1) {real, imag} */,
  {32'h3ee369fa, 32'h41ebd48a} /* (2, 28, 0) {real, imag} */,
  {32'hc20d9a00, 32'hc223aa24} /* (2, 27, 31) {real, imag} */,
  {32'h41377ad8, 32'h412bb034} /* (2, 27, 30) {real, imag} */,
  {32'hc09490dc, 32'hc0a33c4e} /* (2, 27, 29) {real, imag} */,
  {32'hc0546cb6, 32'h40041a87} /* (2, 27, 28) {real, imag} */,
  {32'hbf5fd5a8, 32'h4108ab9a} /* (2, 27, 27) {real, imag} */,
  {32'h40733d33, 32'h40061f0e} /* (2, 27, 26) {real, imag} */,
  {32'hbfdfe2be, 32'hc00fa790} /* (2, 27, 25) {real, imag} */,
  {32'h3ef73f07, 32'hc01c649f} /* (2, 27, 24) {real, imag} */,
  {32'h3faf5049, 32'h3f2c3552} /* (2, 27, 23) {real, imag} */,
  {32'hbf83f3f3, 32'hbf1ff5e1} /* (2, 27, 22) {real, imag} */,
  {32'h4081403c, 32'hbf89dce2} /* (2, 27, 21) {real, imag} */,
  {32'h3faa924b, 32'h3f9ba8a7} /* (2, 27, 20) {real, imag} */,
  {32'h3fe19cd7, 32'hc00646dc} /* (2, 27, 19) {real, imag} */,
  {32'h403e4f88, 32'hbf5918c9} /* (2, 27, 18) {real, imag} */,
  {32'h400d84ed, 32'h3e52e36d} /* (2, 27, 17) {real, imag} */,
  {32'hc0167def, 32'hbf800322} /* (2, 27, 16) {real, imag} */,
  {32'hbecabed2, 32'hbe3e83b4} /* (2, 27, 15) {real, imag} */,
  {32'hbfd9c08a, 32'hbfc23917} /* (2, 27, 14) {real, imag} */,
  {32'h3f98e479, 32'h4001d2a9} /* (2, 27, 13) {real, imag} */,
  {32'hbf4d7003, 32'h3f3ac034} /* (2, 27, 12) {real, imag} */,
  {32'hc0703673, 32'h3f9069a8} /* (2, 27, 11) {real, imag} */,
  {32'hbf22efd5, 32'h40bf93dd} /* (2, 27, 10) {real, imag} */,
  {32'h3f05603b, 32'hbdb55d5a} /* (2, 27, 9) {real, imag} */,
  {32'hc077c079, 32'h3fca8aad} /* (2, 27, 8) {real, imag} */,
  {32'hc046458f, 32'hc053e3f9} /* (2, 27, 7) {real, imag} */,
  {32'hc05e7122, 32'h403d15bd} /* (2, 27, 6) {real, imag} */,
  {32'h41018ed1, 32'h410c01f0} /* (2, 27, 5) {real, imag} */,
  {32'h41263bef, 32'hbfa41740} /* (2, 27, 4) {real, imag} */,
  {32'hc0828427, 32'hc03ae6bd} /* (2, 27, 3) {real, imag} */,
  {32'hc0d6a900, 32'h416ce489} /* (2, 27, 2) {real, imag} */,
  {32'hbfb52aa4, 32'hc2430ab8} /* (2, 27, 1) {real, imag} */,
  {32'hc10f778f, 32'hc20a52cb} /* (2, 27, 0) {real, imag} */,
  {32'hbfbbbb74, 32'hbf383793} /* (2, 26, 31) {real, imag} */,
  {32'h400ba8e4, 32'h40df54e4} /* (2, 26, 30) {real, imag} */,
  {32'h40a52d29, 32'hc00ab742} /* (2, 26, 29) {real, imag} */,
  {32'hc02423f4, 32'hc02631ea} /* (2, 26, 28) {real, imag} */,
  {32'hc00ea5dc, 32'h40c639e6} /* (2, 26, 27) {real, imag} */,
  {32'hbff1eee6, 32'h3d583b31} /* (2, 26, 26) {real, imag} */,
  {32'h3f89ed43, 32'h3f0d0a17} /* (2, 26, 25) {real, imag} */,
  {32'hbfac4e54, 32'h404f757f} /* (2, 26, 24) {real, imag} */,
  {32'hc038f59b, 32'hc01ac9e3} /* (2, 26, 23) {real, imag} */,
  {32'hbf9152c7, 32'hbec5c348} /* (2, 26, 22) {real, imag} */,
  {32'h3f891814, 32'h40145d13} /* (2, 26, 21) {real, imag} */,
  {32'h3f9d4690, 32'h3e14d980} /* (2, 26, 20) {real, imag} */,
  {32'h3f341a9e, 32'h3f8d1a94} /* (2, 26, 19) {real, imag} */,
  {32'hbf81ecea, 32'h3ef75bfa} /* (2, 26, 18) {real, imag} */,
  {32'hbf8b6022, 32'h3f22f123} /* (2, 26, 17) {real, imag} */,
  {32'h40104f9c, 32'hbf26f9d3} /* (2, 26, 16) {real, imag} */,
  {32'h3f7ecd65, 32'h3f383201} /* (2, 26, 15) {real, imag} */,
  {32'hbd3554cf, 32'h3fe6bcef} /* (2, 26, 14) {real, imag} */,
  {32'hbf269f85, 32'h3ff8603c} /* (2, 26, 13) {real, imag} */,
  {32'hbfde9023, 32'hbfe520e5} /* (2, 26, 12) {real, imag} */,
  {32'h3fb2f880, 32'h401c30e8} /* (2, 26, 11) {real, imag} */,
  {32'h3f4552a2, 32'h3f204697} /* (2, 26, 10) {real, imag} */,
  {32'hbf38d4c1, 32'h40868cf5} /* (2, 26, 9) {real, imag} */,
  {32'h40533e14, 32'h3f8a23d2} /* (2, 26, 8) {real, imag} */,
  {32'h3ee0afa2, 32'h3f74096a} /* (2, 26, 7) {real, imag} */,
  {32'h40dfd167, 32'h40285a08} /* (2, 26, 6) {real, imag} */,
  {32'h3e42bb59, 32'h3fedf71c} /* (2, 26, 5) {real, imag} */,
  {32'hc1082d4b, 32'hbf7ffdf3} /* (2, 26, 4) {real, imag} */,
  {32'hbfb39035, 32'h40934042} /* (2, 26, 3) {real, imag} */,
  {32'hbeeca322, 32'h407cd97b} /* (2, 26, 2) {real, imag} */,
  {32'hc0ab581b, 32'hc0cfaf15} /* (2, 26, 1) {real, imag} */,
  {32'h400ee842, 32'h401f88dd} /* (2, 26, 0) {real, imag} */,
  {32'h4116344d, 32'h409cb3fa} /* (2, 25, 31) {real, imag} */,
  {32'hbff72b1a, 32'h3e8c437b} /* (2, 25, 30) {real, imag} */,
  {32'hbf971acd, 32'h4045bb99} /* (2, 25, 29) {real, imag} */,
  {32'hbe8e4c8c, 32'hc000cd59} /* (2, 25, 28) {real, imag} */,
  {32'hc08c1e31, 32'hc05dc5dd} /* (2, 25, 27) {real, imag} */,
  {32'hc09f42e2, 32'h3fdf6b29} /* (2, 25, 26) {real, imag} */,
  {32'hbf44fa0e, 32'h3e35d3fe} /* (2, 25, 25) {real, imag} */,
  {32'hc021cd31, 32'h4035456d} /* (2, 25, 24) {real, imag} */,
  {32'hc02007eb, 32'hbf4b65de} /* (2, 25, 23) {real, imag} */,
  {32'h3e93d9f0, 32'hbfe76b22} /* (2, 25, 22) {real, imag} */,
  {32'h3e4d70cb, 32'h40094139} /* (2, 25, 21) {real, imag} */,
  {32'h3f1c0a62, 32'hbe7f6c42} /* (2, 25, 20) {real, imag} */,
  {32'hc02cd315, 32'h3e46d0db} /* (2, 25, 19) {real, imag} */,
  {32'h3f0ee549, 32'h3f91924d} /* (2, 25, 18) {real, imag} */,
  {32'hbf02a778, 32'h3fa4d687} /* (2, 25, 17) {real, imag} */,
  {32'h404db097, 32'hbfd9263f} /* (2, 25, 16) {real, imag} */,
  {32'hbf633a9a, 32'hc0132e0c} /* (2, 25, 15) {real, imag} */,
  {32'h3fa5eeb8, 32'hc0365c4e} /* (2, 25, 14) {real, imag} */,
  {32'h3fe53981, 32'h40b639a8} /* (2, 25, 13) {real, imag} */,
  {32'hbeebc2a7, 32'h3f6be4c8} /* (2, 25, 12) {real, imag} */,
  {32'hbe9c68da, 32'hbeaa2c27} /* (2, 25, 11) {real, imag} */,
  {32'h3fa5b05d, 32'h3fb79661} /* (2, 25, 10) {real, imag} */,
  {32'hc002b430, 32'hbf9fed16} /* (2, 25, 9) {real, imag} */,
  {32'hbfb65369, 32'hc0390a79} /* (2, 25, 8) {real, imag} */,
  {32'hbe940ca3, 32'h3fcd007a} /* (2, 25, 7) {real, imag} */,
  {32'h3fcb83ca, 32'h3f2d80c7} /* (2, 25, 6) {real, imag} */,
  {32'h3f60cf7f, 32'hbf8cecab} /* (2, 25, 5) {real, imag} */,
  {32'hbfc8589e, 32'hc0588919} /* (2, 25, 4) {real, imag} */,
  {32'hbf317449, 32'h3fe9fd1c} /* (2, 25, 3) {real, imag} */,
  {32'hbfb05b43, 32'hbfa0895a} /* (2, 25, 2) {real, imag} */,
  {32'h409d099d, 32'h406de482} /* (2, 25, 1) {real, imag} */,
  {32'h410132a3, 32'h407580f2} /* (2, 25, 0) {real, imag} */,
  {32'hc103c893, 32'hc14d30fa} /* (2, 24, 31) {real, imag} */,
  {32'h4086c307, 32'h40c036a3} /* (2, 24, 30) {real, imag} */,
  {32'h3f44582d, 32'hbf07b39f} /* (2, 24, 29) {real, imag} */,
  {32'hc00541e7, 32'hc0c45195} /* (2, 24, 28) {real, imag} */,
  {32'h40cf66e5, 32'h40a13f24} /* (2, 24, 27) {real, imag} */,
  {32'h3fadc060, 32'h404ac2b4} /* (2, 24, 26) {real, imag} */,
  {32'hc050fe38, 32'h3f7923c6} /* (2, 24, 25) {real, imag} */,
  {32'h400b8f47, 32'h401068ad} /* (2, 24, 24) {real, imag} */,
  {32'hbf0bf646, 32'hbdace64b} /* (2, 24, 23) {real, imag} */,
  {32'hc05fd871, 32'h3c836b41} /* (2, 24, 22) {real, imag} */,
  {32'h3ffea7ee, 32'h3fc87bd5} /* (2, 24, 21) {real, imag} */,
  {32'h3fe7d96a, 32'hbf9b98c4} /* (2, 24, 20) {real, imag} */,
  {32'h3f6df20d, 32'hbe4e80a3} /* (2, 24, 19) {real, imag} */,
  {32'h3e963049, 32'hbc35f2d2} /* (2, 24, 18) {real, imag} */,
  {32'hbec4b6de, 32'hbe1429a9} /* (2, 24, 17) {real, imag} */,
  {32'hbf35f79b, 32'hbe14305f} /* (2, 24, 16) {real, imag} */,
  {32'h3fe17cab, 32'h3f4f63af} /* (2, 24, 15) {real, imag} */,
  {32'h3f6958db, 32'h3dc5f7eb} /* (2, 24, 14) {real, imag} */,
  {32'h3f5aaa70, 32'h3cb30945} /* (2, 24, 13) {real, imag} */,
  {32'hbd5ad07f, 32'h402eb31a} /* (2, 24, 12) {real, imag} */,
  {32'hbf37e79f, 32'h40676381} /* (2, 24, 11) {real, imag} */,
  {32'h3be8df56, 32'h40d389f4} /* (2, 24, 10) {real, imag} */,
  {32'hbcc6f69c, 32'hc043fa8b} /* (2, 24, 9) {real, imag} */,
  {32'hbfd0148f, 32'h3fb0463e} /* (2, 24, 8) {real, imag} */,
  {32'hc08317a4, 32'hbfd22a32} /* (2, 24, 7) {real, imag} */,
  {32'h3dcd6d0a, 32'hc0822c24} /* (2, 24, 6) {real, imag} */,
  {32'h4028d0d0, 32'h40051b57} /* (2, 24, 5) {real, imag} */,
  {32'hc00cdcc6, 32'hbf7c7aef} /* (2, 24, 4) {real, imag} */,
  {32'hc0aec216, 32'h3fa60cd1} /* (2, 24, 3) {real, imag} */,
  {32'hc0446717, 32'h414d5f80} /* (2, 24, 2) {real, imag} */,
  {32'hc14b4257, 32'hc1d1e713} /* (2, 24, 1) {real, imag} */,
  {32'hc0141188, 32'hc1585f96} /* (2, 24, 0) {real, imag} */,
  {32'h40dae08a, 32'h40d349c8} /* (2, 23, 31) {real, imag} */,
  {32'hc0bdf112, 32'hbec35aff} /* (2, 23, 30) {real, imag} */,
  {32'hc0efe04f, 32'hbfff1d3a} /* (2, 23, 29) {real, imag} */,
  {32'h40b4c74b, 32'hbe9b86a6} /* (2, 23, 28) {real, imag} */,
  {32'h404371d9, 32'h401c770e} /* (2, 23, 27) {real, imag} */,
  {32'h3f1b2971, 32'h3fe8a3f1} /* (2, 23, 26) {real, imag} */,
  {32'h3fb0cd85, 32'h3d8a4d7d} /* (2, 23, 25) {real, imag} */,
  {32'hc0a95a81, 32'hbf35b6fe} /* (2, 23, 24) {real, imag} */,
  {32'h3fe4181b, 32'h3f7fcba9} /* (2, 23, 23) {real, imag} */,
  {32'hbf957808, 32'hc058f46d} /* (2, 23, 22) {real, imag} */,
  {32'hc0434cfd, 32'h3e5fee32} /* (2, 23, 21) {real, imag} */,
  {32'hbefb7c7f, 32'h3f7dcb42} /* (2, 23, 20) {real, imag} */,
  {32'h4027ea93, 32'hc024e155} /* (2, 23, 19) {real, imag} */,
  {32'hbf1b88f5, 32'h3fdb43b0} /* (2, 23, 18) {real, imag} */,
  {32'hbfae2354, 32'hbf8fb503} /* (2, 23, 17) {real, imag} */,
  {32'h3fdbb862, 32'hbf1a24b7} /* (2, 23, 16) {real, imag} */,
  {32'h3fc0eefd, 32'h3ed820ee} /* (2, 23, 15) {real, imag} */,
  {32'h3f6fac7e, 32'h401a3bdf} /* (2, 23, 14) {real, imag} */,
  {32'hbf639d48, 32'h407a5b1d} /* (2, 23, 13) {real, imag} */,
  {32'hc0586504, 32'h402dfbdd} /* (2, 23, 12) {real, imag} */,
  {32'h3fc2820a, 32'hc0333c39} /* (2, 23, 11) {real, imag} */,
  {32'hc00697b3, 32'hc07cea2f} /* (2, 23, 10) {real, imag} */,
  {32'h3ff1bb0f, 32'h3fb7a355} /* (2, 23, 9) {real, imag} */,
  {32'hbf96fcc7, 32'hbfa6bdf0} /* (2, 23, 8) {real, imag} */,
  {32'h3f5b71b7, 32'h3f441f96} /* (2, 23, 7) {real, imag} */,
  {32'h4072dca3, 32'hc004fa01} /* (2, 23, 6) {real, imag} */,
  {32'hbfd18ba2, 32'hbe82b654} /* (2, 23, 5) {real, imag} */,
  {32'h3fe8f894, 32'h4013d56a} /* (2, 23, 4) {real, imag} */,
  {32'h4042ff08, 32'h3e2cbe72} /* (2, 23, 3) {real, imag} */,
  {32'hc0e5553c, 32'hbf9546d4} /* (2, 23, 2) {real, imag} */,
  {32'h403cc6c1, 32'hc0d871fc} /* (2, 23, 1) {real, imag} */,
  {32'h3f80f19a, 32'h3b8ff004} /* (2, 23, 0) {real, imag} */,
  {32'h402067ee, 32'h40af85d4} /* (2, 22, 31) {real, imag} */,
  {32'hc0524f54, 32'hc0c8bcf9} /* (2, 22, 30) {real, imag} */,
  {32'h3f9bda61, 32'h3f89f92e} /* (2, 22, 29) {real, imag} */,
  {32'h402ce9c2, 32'h3ffac0c9} /* (2, 22, 28) {real, imag} */,
  {32'hbec3f03b, 32'h40234dca} /* (2, 22, 27) {real, imag} */,
  {32'hbea6e9ce, 32'h4087ab9c} /* (2, 22, 26) {real, imag} */,
  {32'hbf81f3c4, 32'h3f318ace} /* (2, 22, 25) {real, imag} */,
  {32'hc01bd342, 32'hbfc24fb5} /* (2, 22, 24) {real, imag} */,
  {32'hbd8b9551, 32'h4003df4f} /* (2, 22, 23) {real, imag} */,
  {32'h4011b23f, 32'hbff5dc9c} /* (2, 22, 22) {real, imag} */,
  {32'h3f7926ce, 32'hc0032794} /* (2, 22, 21) {real, imag} */,
  {32'hc01e31c8, 32'hbf7a67c0} /* (2, 22, 20) {real, imag} */,
  {32'hbfa26805, 32'h4016608f} /* (2, 22, 19) {real, imag} */,
  {32'hbff030f7, 32'h3ee4d820} /* (2, 22, 18) {real, imag} */,
  {32'h3f0261cc, 32'hbf3e72b9} /* (2, 22, 17) {real, imag} */,
  {32'h3fe302b1, 32'hc003d098} /* (2, 22, 16) {real, imag} */,
  {32'h3f6a7b94, 32'h3fd81380} /* (2, 22, 15) {real, imag} */,
  {32'h3fed0775, 32'h3f879a89} /* (2, 22, 14) {real, imag} */,
  {32'h401def0d, 32'h3f13c16c} /* (2, 22, 13) {real, imag} */,
  {32'hbf1e2bd6, 32'hbea57529} /* (2, 22, 12) {real, imag} */,
  {32'hc0624645, 32'h3fcf80a3} /* (2, 22, 11) {real, imag} */,
  {32'hbfaebed2, 32'h3fd1c02f} /* (2, 22, 10) {real, imag} */,
  {32'h3db9be4b, 32'hbd8e55e5} /* (2, 22, 9) {real, imag} */,
  {32'hbf9ed3a4, 32'hc03843ca} /* (2, 22, 8) {real, imag} */,
  {32'h3ffee535, 32'hc0080e2b} /* (2, 22, 7) {real, imag} */,
  {32'hbf1edca7, 32'hc017460f} /* (2, 22, 6) {real, imag} */,
  {32'hbf330c93, 32'hc05e96a0} /* (2, 22, 5) {real, imag} */,
  {32'hbfda24c3, 32'h3f0077d1} /* (2, 22, 4) {real, imag} */,
  {32'h404154b9, 32'h3fc513ca} /* (2, 22, 3) {real, imag} */,
  {32'hbf36eab4, 32'h401f84ca} /* (2, 22, 2) {real, imag} */,
  {32'h40edf53b, 32'hc010c10c} /* (2, 22, 1) {real, imag} */,
  {32'h401e1d87, 32'h3ed9ff22} /* (2, 22, 0) {real, imag} */,
  {32'hc11634fd, 32'hc0a70247} /* (2, 21, 31) {real, imag} */,
  {32'h40b6f6bf, 32'h3f54f47d} /* (2, 21, 30) {real, imag} */,
  {32'hbf2e1987, 32'h401023f8} /* (2, 21, 29) {real, imag} */,
  {32'hbfb8da4c, 32'h3fbc551d} /* (2, 21, 28) {real, imag} */,
  {32'h408e3ba2, 32'h400511be} /* (2, 21, 27) {real, imag} */,
  {32'h3fe2611d, 32'hc00a8cb7} /* (2, 21, 26) {real, imag} */,
  {32'hbef1ead0, 32'h400c3875} /* (2, 21, 25) {real, imag} */,
  {32'h406546bd, 32'h3e96d5c4} /* (2, 21, 24) {real, imag} */,
  {32'hbfc0ad53, 32'h3ffce433} /* (2, 21, 23) {real, imag} */,
  {32'h405ad45e, 32'h40c3f160} /* (2, 21, 22) {real, imag} */,
  {32'h3ff61c0f, 32'h3ff6a365} /* (2, 21, 21) {real, imag} */,
  {32'hc06e3e5c, 32'h3c23d8d9} /* (2, 21, 20) {real, imag} */,
  {32'h3f86bad5, 32'hbd590e49} /* (2, 21, 19) {real, imag} */,
  {32'hbf2afb14, 32'hbf77d69a} /* (2, 21, 18) {real, imag} */,
  {32'hbea223ca, 32'h3eca8b92} /* (2, 21, 17) {real, imag} */,
  {32'hc02c0bcf, 32'hbfb3676b} /* (2, 21, 16) {real, imag} */,
  {32'h401df63e, 32'hbef08ec5} /* (2, 21, 15) {real, imag} */,
  {32'h3e85e50a, 32'h3e683e83} /* (2, 21, 14) {real, imag} */,
  {32'hbf361a24, 32'h3e8c92ac} /* (2, 21, 13) {real, imag} */,
  {32'hbf9a3255, 32'hbfc54290} /* (2, 21, 12) {real, imag} */,
  {32'h3f653a69, 32'h405f38dd} /* (2, 21, 11) {real, imag} */,
  {32'h3fd1c944, 32'hbfad667b} /* (2, 21, 10) {real, imag} */,
  {32'h3f52bea4, 32'h3fa3ae8f} /* (2, 21, 9) {real, imag} */,
  {32'hbe152fa2, 32'h4071c05e} /* (2, 21, 8) {real, imag} */,
  {32'hbfbbf7e2, 32'h3f2a9c4d} /* (2, 21, 7) {real, imag} */,
  {32'h3f9909d3, 32'hc03abf95} /* (2, 21, 6) {real, imag} */,
  {32'h401b59f1, 32'h4042d322} /* (2, 21, 5) {real, imag} */,
  {32'h4051feca, 32'hbd1ed3b3} /* (2, 21, 4) {real, imag} */,
  {32'hbfc382f3, 32'h4080ca19} /* (2, 21, 3) {real, imag} */,
  {32'h40161f93, 32'h4000055f} /* (2, 21, 2) {real, imag} */,
  {32'hc0d83fd2, 32'hc0fd7c8f} /* (2, 21, 1) {real, imag} */,
  {32'hc087d318, 32'hc1142422} /* (2, 21, 0) {real, imag} */,
  {32'h3f830da1, 32'hbf64442d} /* (2, 20, 31) {real, imag} */,
  {32'hbfef002e, 32'h3e60a826} /* (2, 20, 30) {real, imag} */,
  {32'h4003f506, 32'h3fd5646f} /* (2, 20, 29) {real, imag} */,
  {32'hbfa1da36, 32'h3fc38145} /* (2, 20, 28) {real, imag} */,
  {32'h3d5ab544, 32'h3fb682e5} /* (2, 20, 27) {real, imag} */,
  {32'h3dc9fff4, 32'h4024c2fd} /* (2, 20, 26) {real, imag} */,
  {32'hbf97ea64, 32'hbf315d5e} /* (2, 20, 25) {real, imag} */,
  {32'h3f10e1b9, 32'h3f3cd8d9} /* (2, 20, 24) {real, imag} */,
  {32'hbf166e1a, 32'hc0b0ba38} /* (2, 20, 23) {real, imag} */,
  {32'h3f7b2998, 32'h402d0035} /* (2, 20, 22) {real, imag} */,
  {32'h3f8367aa, 32'h3fa6ada0} /* (2, 20, 21) {real, imag} */,
  {32'hc01ad6b7, 32'hbf96e081} /* (2, 20, 20) {real, imag} */,
  {32'hbfeb9f85, 32'h3fe3d686} /* (2, 20, 19) {real, imag} */,
  {32'hbf184a9e, 32'hc03ebb59} /* (2, 20, 18) {real, imag} */,
  {32'h3e3b7ffe, 32'h3e7717d1} /* (2, 20, 17) {real, imag} */,
  {32'hbea27dd6, 32'hbd5e071b} /* (2, 20, 16) {real, imag} */,
  {32'hc016a76f, 32'hbf903f42} /* (2, 20, 15) {real, imag} */,
  {32'hbed449eb, 32'hbfea7604} /* (2, 20, 14) {real, imag} */,
  {32'h3f803f17, 32'h3eb969b8} /* (2, 20, 13) {real, imag} */,
  {32'h3f48252b, 32'hc04e2a35} /* (2, 20, 12) {real, imag} */,
  {32'h3db5c9d1, 32'hbe4f6297} /* (2, 20, 11) {real, imag} */,
  {32'hbf45576f, 32'h3f480a09} /* (2, 20, 10) {real, imag} */,
  {32'hc0404ab5, 32'hbfec11f4} /* (2, 20, 9) {real, imag} */,
  {32'h40144552, 32'hbf9416e1} /* (2, 20, 8) {real, imag} */,
  {32'hbe22386b, 32'h3dfd29f3} /* (2, 20, 7) {real, imag} */,
  {32'hbfaa89f7, 32'h3faee495} /* (2, 20, 6) {real, imag} */,
  {32'h3f49aed2, 32'hbfd5a8cc} /* (2, 20, 5) {real, imag} */,
  {32'hbf0ce45a, 32'h3ece7084} /* (2, 20, 4) {real, imag} */,
  {32'hbdd920d6, 32'hbf1023bb} /* (2, 20, 3) {real, imag} */,
  {32'h400f9ab1, 32'h3e4e5192} /* (2, 20, 2) {real, imag} */,
  {32'h4041e90d, 32'hbf45d973} /* (2, 20, 1) {real, imag} */,
  {32'hc0188b30, 32'h403abde7} /* (2, 20, 0) {real, imag} */,
  {32'h4027c2bf, 32'h408de4f8} /* (2, 19, 31) {real, imag} */,
  {32'hbe4aa8c2, 32'hbf85c364} /* (2, 19, 30) {real, imag} */,
  {32'hbf18dde4, 32'hbefe5ffa} /* (2, 19, 29) {real, imag} */,
  {32'h3fad63c0, 32'h401a8e24} /* (2, 19, 28) {real, imag} */,
  {32'hbf347e71, 32'hc0105b3c} /* (2, 19, 27) {real, imag} */,
  {32'hbfa33dcf, 32'hc000a268} /* (2, 19, 26) {real, imag} */,
  {32'hbf98f65e, 32'h407fcefa} /* (2, 19, 25) {real, imag} */,
  {32'hc001d2f1, 32'hbed6ba79} /* (2, 19, 24) {real, imag} */,
  {32'h3fad5921, 32'hbf7f5e28} /* (2, 19, 23) {real, imag} */,
  {32'hbf2594ea, 32'hbd415764} /* (2, 19, 22) {real, imag} */,
  {32'hbf6a1753, 32'hbf2181c4} /* (2, 19, 21) {real, imag} */,
  {32'hbfde8cd1, 32'h3f82afc9} /* (2, 19, 20) {real, imag} */,
  {32'h3e7955c6, 32'h3f3691ce} /* (2, 19, 19) {real, imag} */,
  {32'hbf808ba9, 32'h404d7bd5} /* (2, 19, 18) {real, imag} */,
  {32'h3f6e3d1f, 32'h3e981ea9} /* (2, 19, 17) {real, imag} */,
  {32'h4009719f, 32'h3a8a8aa1} /* (2, 19, 16) {real, imag} */,
  {32'hbe207fe6, 32'hbf53daef} /* (2, 19, 15) {real, imag} */,
  {32'h400ca525, 32'hbfbd6807} /* (2, 19, 14) {real, imag} */,
  {32'h3e020355, 32'hbe8d346d} /* (2, 19, 13) {real, imag} */,
  {32'h400af863, 32'h3e0c32f9} /* (2, 19, 12) {real, imag} */,
  {32'h3c0fa1fb, 32'hbfabf2aa} /* (2, 19, 11) {real, imag} */,
  {32'h3f558019, 32'h40164741} /* (2, 19, 10) {real, imag} */,
  {32'h3fb63967, 32'h3f90f324} /* (2, 19, 9) {real, imag} */,
  {32'hbf7225a6, 32'hbf8acfb0} /* (2, 19, 8) {real, imag} */,
  {32'hc0017bf5, 32'h3d811f65} /* (2, 19, 7) {real, imag} */,
  {32'hc0663078, 32'h406e35a3} /* (2, 19, 6) {real, imag} */,
  {32'h3ed760a5, 32'h40181080} /* (2, 19, 5) {real, imag} */,
  {32'h3f9c36c9, 32'h404fb744} /* (2, 19, 4) {real, imag} */,
  {32'hbf8d9f0f, 32'h3e9a720f} /* (2, 19, 3) {real, imag} */,
  {32'h3c3a7e8b, 32'h3f0c9e01} /* (2, 19, 2) {real, imag} */,
  {32'h3f167f77, 32'h3f6fd0d9} /* (2, 19, 1) {real, imag} */,
  {32'h4024e6a6, 32'h3f62951e} /* (2, 19, 0) {real, imag} */,
  {32'hc039f520, 32'h3fbd2dc4} /* (2, 18, 31) {real, imag} */,
  {32'h3ef7e8ab, 32'hbf999573} /* (2, 18, 30) {real, imag} */,
  {32'h3f34918f, 32'h3e1f1117} /* (2, 18, 29) {real, imag} */,
  {32'h3ce1a10c, 32'hbfbe9973} /* (2, 18, 28) {real, imag} */,
  {32'h3fb93c7f, 32'hbfd757a5} /* (2, 18, 27) {real, imag} */,
  {32'h40144aac, 32'h3f7e1e67} /* (2, 18, 26) {real, imag} */,
  {32'h3f8c4433, 32'h3e91bfd9} /* (2, 18, 25) {real, imag} */,
  {32'h3f84a796, 32'h3f227935} /* (2, 18, 24) {real, imag} */,
  {32'h3e375f59, 32'h4020995b} /* (2, 18, 23) {real, imag} */,
  {32'hbf970306, 32'h40235455} /* (2, 18, 22) {real, imag} */,
  {32'h3f986ef5, 32'hbeabe36b} /* (2, 18, 21) {real, imag} */,
  {32'h3fe3501d, 32'hbfc89809} /* (2, 18, 20) {real, imag} */,
  {32'hc00baa15, 32'h3d9bafc8} /* (2, 18, 19) {real, imag} */,
  {32'h3f9f1164, 32'h3f95fc4f} /* (2, 18, 18) {real, imag} */,
  {32'hbe3b1b0d, 32'hbf809acd} /* (2, 18, 17) {real, imag} */,
  {32'hbfcc525d, 32'h3eabfa8d} /* (2, 18, 16) {real, imag} */,
  {32'h3f46311f, 32'h3f8a90e7} /* (2, 18, 15) {real, imag} */,
  {32'h3fc2d00f, 32'hbecef339} /* (2, 18, 14) {real, imag} */,
  {32'h3fbdb3f7, 32'hbffd256c} /* (2, 18, 13) {real, imag} */,
  {32'hbf97c1fe, 32'hbe374f27} /* (2, 18, 12) {real, imag} */,
  {32'hbd267e65, 32'h3f0e2d65} /* (2, 18, 11) {real, imag} */,
  {32'h3ed4d428, 32'h3f67edb7} /* (2, 18, 10) {real, imag} */,
  {32'h3e00b2ee, 32'hbf72030c} /* (2, 18, 9) {real, imag} */,
  {32'h3fce23ee, 32'h405d582c} /* (2, 18, 8) {real, imag} */,
  {32'hbf5f0621, 32'h3d9115b9} /* (2, 18, 7) {real, imag} */,
  {32'h3f874b47, 32'h3f8b94cf} /* (2, 18, 6) {real, imag} */,
  {32'hbe4f082e, 32'h3fdb740a} /* (2, 18, 5) {real, imag} */,
  {32'hc04ac1a3, 32'hc0ae0cff} /* (2, 18, 4) {real, imag} */,
  {32'h3ffcbf43, 32'hbf919b54} /* (2, 18, 3) {real, imag} */,
  {32'h3fc5d93d, 32'h404e9c1d} /* (2, 18, 2) {real, imag} */,
  {32'hc0819833, 32'hc0940d7e} /* (2, 18, 1) {real, imag} */,
  {32'hc051c253, 32'h3fd38a5d} /* (2, 18, 0) {real, imag} */,
  {32'h3fed4cc6, 32'h3f86f184} /* (2, 17, 31) {real, imag} */,
  {32'hc01d685a, 32'h3f1035ad} /* (2, 17, 30) {real, imag} */,
  {32'hbec63898, 32'hbdf43195} /* (2, 17, 29) {real, imag} */,
  {32'h3fb129a9, 32'hc0048c79} /* (2, 17, 28) {real, imag} */,
  {32'hbf2c1aa8, 32'h3f832976} /* (2, 17, 27) {real, imag} */,
  {32'h3fcee70e, 32'hbfdd1bcb} /* (2, 17, 26) {real, imag} */,
  {32'h3b52da9e, 32'h4036722c} /* (2, 17, 25) {real, imag} */,
  {32'hbf64a18c, 32'h3f6f5abd} /* (2, 17, 24) {real, imag} */,
  {32'h3fd13bc1, 32'h3e38cfb0} /* (2, 17, 23) {real, imag} */,
  {32'h3fc862b8, 32'hbfb6139f} /* (2, 17, 22) {real, imag} */,
  {32'h3eca1e25, 32'h3ffb9fad} /* (2, 17, 21) {real, imag} */,
  {32'hbf378cbe, 32'hc001e98b} /* (2, 17, 20) {real, imag} */,
  {32'h3e36842d, 32'h3d841183} /* (2, 17, 19) {real, imag} */,
  {32'hc0514631, 32'h3f54ac0d} /* (2, 17, 18) {real, imag} */,
  {32'hbf962a58, 32'hbd634a7c} /* (2, 17, 17) {real, imag} */,
  {32'h3e8b3d63, 32'hbfb1706e} /* (2, 17, 16) {real, imag} */,
  {32'hbf7ea8cd, 32'h4016321b} /* (2, 17, 15) {real, imag} */,
  {32'h3ede5885, 32'hc021e01a} /* (2, 17, 14) {real, imag} */,
  {32'hbeb83b4f, 32'h3e4f7675} /* (2, 17, 13) {real, imag} */,
  {32'hbead762c, 32'h3dd9efe1} /* (2, 17, 12) {real, imag} */,
  {32'hbf1913e5, 32'h3f5c19cd} /* (2, 17, 11) {real, imag} */,
  {32'h3fe2f660, 32'hbefbe3af} /* (2, 17, 10) {real, imag} */,
  {32'hbf308bb1, 32'hbee0ce75} /* (2, 17, 9) {real, imag} */,
  {32'h3f8426c4, 32'h3f1f4ffd} /* (2, 17, 8) {real, imag} */,
  {32'hbe52aa6a, 32'hbf8f971e} /* (2, 17, 7) {real, imag} */,
  {32'h3f8fe955, 32'h3f9b4580} /* (2, 17, 6) {real, imag} */,
  {32'h3f9b2e0d, 32'h3c8f4fce} /* (2, 17, 5) {real, imag} */,
  {32'hbe63ec37, 32'h40137263} /* (2, 17, 4) {real, imag} */,
  {32'h3d090f9b, 32'h3f5f4cc2} /* (2, 17, 3) {real, imag} */,
  {32'hc03989f2, 32'hbe4cdd42} /* (2, 17, 2) {real, imag} */,
  {32'h408264ae, 32'hbfa46882} /* (2, 17, 1) {real, imag} */,
  {32'h403cc802, 32'hbfc9221a} /* (2, 17, 0) {real, imag} */,
  {32'hbfc11956, 32'hbfb36792} /* (2, 16, 31) {real, imag} */,
  {32'hbe9b09e2, 32'h3c23c428} /* (2, 16, 30) {real, imag} */,
  {32'h3f535c47, 32'hbe216b3d} /* (2, 16, 29) {real, imag} */,
  {32'h3dbce757, 32'h3e844ff9} /* (2, 16, 28) {real, imag} */,
  {32'hbf5b97de, 32'h3f9021bf} /* (2, 16, 27) {real, imag} */,
  {32'hbfe45997, 32'h3efe6e89} /* (2, 16, 26) {real, imag} */,
  {32'hbf1dec47, 32'h3f59efa8} /* (2, 16, 25) {real, imag} */,
  {32'h3fdce25e, 32'hbf813f15} /* (2, 16, 24) {real, imag} */,
  {32'h3f50a68f, 32'hbeff9adf} /* (2, 16, 23) {real, imag} */,
  {32'hbd22b248, 32'h403f956f} /* (2, 16, 22) {real, imag} */,
  {32'h3fb2a05e, 32'h3f80d188} /* (2, 16, 21) {real, imag} */,
  {32'hbeefe73a, 32'h3e9dae99} /* (2, 16, 20) {real, imag} */,
  {32'hbf96c174, 32'hbe11cd9d} /* (2, 16, 19) {real, imag} */,
  {32'h3f903413, 32'h3f51521f} /* (2, 16, 18) {real, imag} */,
  {32'hbf153aa6, 32'h3f8245c7} /* (2, 16, 17) {real, imag} */,
  {32'hbeb8eca6, 32'h3f6609bd} /* (2, 16, 16) {real, imag} */,
  {32'hbfc3e2ff, 32'h4005a201} /* (2, 16, 15) {real, imag} */,
  {32'h3e19b8b7, 32'h3e5f7184} /* (2, 16, 14) {real, imag} */,
  {32'hbfa0d6a2, 32'hc036ebde} /* (2, 16, 13) {real, imag} */,
  {32'hbd400c2e, 32'hbfb1e9be} /* (2, 16, 12) {real, imag} */,
  {32'hbf93c723, 32'h3e9a27bf} /* (2, 16, 11) {real, imag} */,
  {32'h3fe4ca01, 32'h3f200283} /* (2, 16, 10) {real, imag} */,
  {32'h3f3e7f8d, 32'h3f8ae11f} /* (2, 16, 9) {real, imag} */,
  {32'hbed7b09e, 32'h3f75ec2b} /* (2, 16, 8) {real, imag} */,
  {32'hbe67cc25, 32'hbdd75498} /* (2, 16, 7) {real, imag} */,
  {32'h3f64b4d5, 32'hbf2a2c1d} /* (2, 16, 6) {real, imag} */,
  {32'h3f9b1824, 32'h3e8661d1} /* (2, 16, 5) {real, imag} */,
  {32'h3fd1cd1f, 32'h3ff36b99} /* (2, 16, 4) {real, imag} */,
  {32'hbf6ee17e, 32'h3f35a41e} /* (2, 16, 3) {real, imag} */,
  {32'hbf95846a, 32'hbf2e5dc4} /* (2, 16, 2) {real, imag} */,
  {32'h3d2a8ef2, 32'h3f0b27ee} /* (2, 16, 1) {real, imag} */,
  {32'hbfbd63ef, 32'hbf1c93f1} /* (2, 16, 0) {real, imag} */,
  {32'hbf87beba, 32'hbfc0b241} /* (2, 15, 31) {real, imag} */,
  {32'h3f499053, 32'hbfbaadcf} /* (2, 15, 30) {real, imag} */,
  {32'h3fa055cc, 32'h402e91d4} /* (2, 15, 29) {real, imag} */,
  {32'hbe973e0f, 32'h3f219783} /* (2, 15, 28) {real, imag} */,
  {32'h3f7893a9, 32'hbed54d85} /* (2, 15, 27) {real, imag} */,
  {32'hc0237e66, 32'h3eea66a0} /* (2, 15, 26) {real, imag} */,
  {32'h3e0da0c3, 32'h3ef5fb57} /* (2, 15, 25) {real, imag} */,
  {32'h3f87ed2e, 32'h3f26f9ca} /* (2, 15, 24) {real, imag} */,
  {32'h3fd241c1, 32'h3ff9c11c} /* (2, 15, 23) {real, imag} */,
  {32'h3fe98f3b, 32'h3fbefbe2} /* (2, 15, 22) {real, imag} */,
  {32'h3f8a79e4, 32'h3e42fda9} /* (2, 15, 21) {real, imag} */,
  {32'h3f4dbaf0, 32'hbe99a59d} /* (2, 15, 20) {real, imag} */,
  {32'hbf290bf8, 32'hbf98aea4} /* (2, 15, 19) {real, imag} */,
  {32'hbf1dc105, 32'h3ed29d0c} /* (2, 15, 18) {real, imag} */,
  {32'h3e61fc98, 32'h3ebf007a} /* (2, 15, 17) {real, imag} */,
  {32'hbeb61216, 32'hbf190227} /* (2, 15, 16) {real, imag} */,
  {32'h3f99762f, 32'hbf4db926} /* (2, 15, 15) {real, imag} */,
  {32'hbf302cb2, 32'h3f1c0c3e} /* (2, 15, 14) {real, imag} */,
  {32'h3ec18d89, 32'hbf3b481f} /* (2, 15, 13) {real, imag} */,
  {32'h400b4d36, 32'h3edb924e} /* (2, 15, 12) {real, imag} */,
  {32'h3fb281e5, 32'h3fb785a1} /* (2, 15, 11) {real, imag} */,
  {32'hbda8d4c4, 32'hbfcd6ddb} /* (2, 15, 10) {real, imag} */,
  {32'h3f738082, 32'hbec75fb0} /* (2, 15, 9) {real, imag} */,
  {32'hbf9d4eda, 32'h3ed8f8de} /* (2, 15, 8) {real, imag} */,
  {32'h4025073f, 32'hbfbfd775} /* (2, 15, 7) {real, imag} */,
  {32'hc089e295, 32'hbe6af85e} /* (2, 15, 6) {real, imag} */,
  {32'hbe8f61ef, 32'h3f4c832f} /* (2, 15, 5) {real, imag} */,
  {32'h400921f4, 32'hbee9a74a} /* (2, 15, 4) {real, imag} */,
  {32'hbeb9abda, 32'h3fb41cb9} /* (2, 15, 3) {real, imag} */,
  {32'h3ffdff6d, 32'hbfd64126} /* (2, 15, 2) {real, imag} */,
  {32'hc0275bc6, 32'hc00bd609} /* (2, 15, 1) {real, imag} */,
  {32'hbfd39531, 32'hbf2f58f4} /* (2, 15, 0) {real, imag} */,
  {32'h4095b446, 32'hc04728ae} /* (2, 14, 31) {real, imag} */,
  {32'hc0856d79, 32'h3fe3a18f} /* (2, 14, 30) {real, imag} */,
  {32'hbfa73ed6, 32'hc00448b9} /* (2, 14, 29) {real, imag} */,
  {32'h400f191e, 32'h3f16e86f} /* (2, 14, 28) {real, imag} */,
  {32'hc011dcb3, 32'h3e5c4feb} /* (2, 14, 27) {real, imag} */,
  {32'h40920ed7, 32'hbeff3c88} /* (2, 14, 26) {real, imag} */,
  {32'h3dc90418, 32'h3fbddf0e} /* (2, 14, 25) {real, imag} */,
  {32'h3e862827, 32'h3fa64f07} /* (2, 14, 24) {real, imag} */,
  {32'h3f60ef85, 32'hbf155e4f} /* (2, 14, 23) {real, imag} */,
  {32'hbf7a8ea2, 32'hbe9ff295} /* (2, 14, 22) {real, imag} */,
  {32'h3f01c0b1, 32'hbf806591} /* (2, 14, 21) {real, imag} */,
  {32'h400eed84, 32'hbf08801f} /* (2, 14, 20) {real, imag} */,
  {32'h3f993cb2, 32'h402a1f5c} /* (2, 14, 19) {real, imag} */,
  {32'hbf569975, 32'h3dbd897a} /* (2, 14, 18) {real, imag} */,
  {32'h3f51c217, 32'h3fd05436} /* (2, 14, 17) {real, imag} */,
  {32'h3f3c6ac0, 32'h3f84fc21} /* (2, 14, 16) {real, imag} */,
  {32'h3f9cc3d5, 32'hbfac8da3} /* (2, 14, 15) {real, imag} */,
  {32'h3f93e4fb, 32'hbf124506} /* (2, 14, 14) {real, imag} */,
  {32'h3f6ee5ad, 32'hbe206ed3} /* (2, 14, 13) {real, imag} */,
  {32'h3f3512f6, 32'h3df1ad91} /* (2, 14, 12) {real, imag} */,
  {32'h3fc3bf37, 32'hc024d126} /* (2, 14, 11) {real, imag} */,
  {32'h3c60277b, 32'hbebb346d} /* (2, 14, 10) {real, imag} */,
  {32'hbf4be799, 32'hbf4be052} /* (2, 14, 9) {real, imag} */,
  {32'hbf671e1c, 32'hbf3f2154} /* (2, 14, 8) {real, imag} */,
  {32'h4029df99, 32'hbefd6d1a} /* (2, 14, 7) {real, imag} */,
  {32'hbfb11a5c, 32'h3e0df049} /* (2, 14, 6) {real, imag} */,
  {32'hbf888358, 32'hbe8c922d} /* (2, 14, 5) {real, imag} */,
  {32'h40648148, 32'hc0796f1b} /* (2, 14, 4) {real, imag} */,
  {32'hbf8fe52f, 32'hbdce051e} /* (2, 14, 3) {real, imag} */,
  {32'hc06c1028, 32'h3e8b2706} /* (2, 14, 2) {real, imag} */,
  {32'h4071b038, 32'h3f406ef5} /* (2, 14, 1) {real, imag} */,
  {32'h40679b7a, 32'h3f12f625} /* (2, 14, 0) {real, imag} */,
  {32'h3d87f1c7, 32'hbf94acf3} /* (2, 13, 31) {real, imag} */,
  {32'h4016249b, 32'h3fda266c} /* (2, 13, 30) {real, imag} */,
  {32'hbf684ed6, 32'h3d915c11} /* (2, 13, 29) {real, imag} */,
  {32'h3ee560b9, 32'h3f45e288} /* (2, 13, 28) {real, imag} */,
  {32'hbf91f709, 32'hbf1f2254} /* (2, 13, 27) {real, imag} */,
  {32'hbf1ff56d, 32'h3e846584} /* (2, 13, 26) {real, imag} */,
  {32'h3ff1cfb7, 32'hbf846642} /* (2, 13, 25) {real, imag} */,
  {32'hbf192290, 32'h3f8897a3} /* (2, 13, 24) {real, imag} */,
  {32'hbfaf0d8c, 32'hbda2993d} /* (2, 13, 23) {real, imag} */,
  {32'hbea8a7bb, 32'hbfa629ad} /* (2, 13, 22) {real, imag} */,
  {32'hbd15af26, 32'h3e223007} /* (2, 13, 21) {real, imag} */,
  {32'h3f251e72, 32'h3f11f805} /* (2, 13, 20) {real, imag} */,
  {32'hbf00f903, 32'hbf23f217} /* (2, 13, 19) {real, imag} */,
  {32'hbd837598, 32'hbfb323c2} /* (2, 13, 18) {real, imag} */,
  {32'hbe994fc6, 32'h3f9f8d6b} /* (2, 13, 17) {real, imag} */,
  {32'h3f1c5c45, 32'h3ea8beff} /* (2, 13, 16) {real, imag} */,
  {32'h3edb208e, 32'hbeade901} /* (2, 13, 15) {real, imag} */,
  {32'hbea9eae6, 32'h404c2600} /* (2, 13, 14) {real, imag} */,
  {32'hbeb81d64, 32'h3fa151b2} /* (2, 13, 13) {real, imag} */,
  {32'h3e3a3e03, 32'hc03085b7} /* (2, 13, 12) {real, imag} */,
  {32'h3f5e4a31, 32'h3f753208} /* (2, 13, 11) {real, imag} */,
  {32'hbea494ea, 32'h3eded19e} /* (2, 13, 10) {real, imag} */,
  {32'h3ed75885, 32'hbe2f0b51} /* (2, 13, 9) {real, imag} */,
  {32'h3eaa56c2, 32'hbfc8ab17} /* (2, 13, 8) {real, imag} */,
  {32'hbdd70d4c, 32'h4073100a} /* (2, 13, 7) {real, imag} */,
  {32'h3f8de987, 32'hbf8c99a5} /* (2, 13, 6) {real, imag} */,
  {32'hc00a1492, 32'hbdd1c659} /* (2, 13, 5) {real, imag} */,
  {32'hbf948cb3, 32'hbfdcf08a} /* (2, 13, 4) {real, imag} */,
  {32'hbd64f06c, 32'hbf0a2adb} /* (2, 13, 3) {real, imag} */,
  {32'hbfb6d199, 32'hbf14cf3d} /* (2, 13, 2) {real, imag} */,
  {32'hbfc53271, 32'hbeb9a809} /* (2, 13, 1) {real, imag} */,
  {32'h3ea36205, 32'h3fcf19ae} /* (2, 13, 0) {real, imag} */,
  {32'hbf51c6c6, 32'h3fc55aaf} /* (2, 12, 31) {real, imag} */,
  {32'h3f600548, 32'h401a4eb5} /* (2, 12, 30) {real, imag} */,
  {32'h3fcd2e63, 32'hc081f2fe} /* (2, 12, 29) {real, imag} */,
  {32'hbe86f8e4, 32'hbf363068} /* (2, 12, 28) {real, imag} */,
  {32'hbf9a5334, 32'h3fe84c42} /* (2, 12, 27) {real, imag} */,
  {32'h3fee84ea, 32'hc04239ad} /* (2, 12, 26) {real, imag} */,
  {32'hc001c4bd, 32'hbf8a893b} /* (2, 12, 25) {real, imag} */,
  {32'h401f4d75, 32'h3e6b58fd} /* (2, 12, 24) {real, imag} */,
  {32'h3ecd4d3c, 32'h3cbbbd92} /* (2, 12, 23) {real, imag} */,
  {32'hbfa0ca4b, 32'h3fe53003} /* (2, 12, 22) {real, imag} */,
  {32'h3f1e3824, 32'hbf728698} /* (2, 12, 21) {real, imag} */,
  {32'hbf87a7ba, 32'hbe2ea960} /* (2, 12, 20) {real, imag} */,
  {32'hc0072257, 32'hbd3942a2} /* (2, 12, 19) {real, imag} */,
  {32'hbcb80cfa, 32'h3ff0b890} /* (2, 12, 18) {real, imag} */,
  {32'hbfafabda, 32'hbfce57c0} /* (2, 12, 17) {real, imag} */,
  {32'hbd3d68a9, 32'h3f63e5b6} /* (2, 12, 16) {real, imag} */,
  {32'hbf0189ff, 32'hbf60a596} /* (2, 12, 15) {real, imag} */,
  {32'hbf62b5d7, 32'hbff69330} /* (2, 12, 14) {real, imag} */,
  {32'h3ff531d8, 32'h3f9aedee} /* (2, 12, 13) {real, imag} */,
  {32'hbfed576a, 32'hbfb68ee0} /* (2, 12, 12) {real, imag} */,
  {32'h3f5f4ba3, 32'h3fa1c197} /* (2, 12, 11) {real, imag} */,
  {32'hbf805a4c, 32'h4042b7c7} /* (2, 12, 10) {real, imag} */,
  {32'h3f75a34d, 32'hbed05fd0} /* (2, 12, 9) {real, imag} */,
  {32'h404a452c, 32'hc0538745} /* (2, 12, 8) {real, imag} */,
  {32'hbe2c4b4f, 32'hbdc432d0} /* (2, 12, 7) {real, imag} */,
  {32'h3ff0e87e, 32'hbfbe53b7} /* (2, 12, 6) {real, imag} */,
  {32'hbf3b984a, 32'hc03ea07e} /* (2, 12, 5) {real, imag} */,
  {32'hbf257e10, 32'hbfe19a1e} /* (2, 12, 4) {real, imag} */,
  {32'hbfd2457b, 32'h406dc6dc} /* (2, 12, 3) {real, imag} */,
  {32'hbf10ce1c, 32'hbfad2953} /* (2, 12, 2) {real, imag} */,
  {32'h3f2d7aa5, 32'h3ffd3363} /* (2, 12, 1) {real, imag} */,
  {32'hbf7bfbb2, 32'h3e700dbf} /* (2, 12, 0) {real, imag} */,
  {32'h40aeaf72, 32'hc09553f5} /* (2, 11, 31) {real, imag} */,
  {32'hc097ba39, 32'h40bdb837} /* (2, 11, 30) {real, imag} */,
  {32'h3dc8369d, 32'h40174600} /* (2, 11, 29) {real, imag} */,
  {32'hbff18544, 32'h3fc52931} /* (2, 11, 28) {real, imag} */,
  {32'hbf10a447, 32'hbf3a1691} /* (2, 11, 27) {real, imag} */,
  {32'h4035ff47, 32'h4008ef82} /* (2, 11, 26) {real, imag} */,
  {32'h3fdb5843, 32'h3eb255f4} /* (2, 11, 25) {real, imag} */,
  {32'hbe6cc9f7, 32'hbf71f8de} /* (2, 11, 24) {real, imag} */,
  {32'h4023b5a1, 32'hc01dc97a} /* (2, 11, 23) {real, imag} */,
  {32'h3f97c63e, 32'hbf742f40} /* (2, 11, 22) {real, imag} */,
  {32'hbf1a43b3, 32'h402a7ae5} /* (2, 11, 21) {real, imag} */,
  {32'hc0016e2d, 32'h3f873c1f} /* (2, 11, 20) {real, imag} */,
  {32'hc0024b73, 32'hbfdc7722} /* (2, 11, 19) {real, imag} */,
  {32'h3fe48f97, 32'hc008f1cc} /* (2, 11, 18) {real, imag} */,
  {32'h3df9183f, 32'h3eaf0472} /* (2, 11, 17) {real, imag} */,
  {32'hbf279864, 32'hbf92f11b} /* (2, 11, 16) {real, imag} */,
  {32'h3f9f6b74, 32'h3f166674} /* (2, 11, 15) {real, imag} */,
  {32'h3e84ae6e, 32'h403fd7fb} /* (2, 11, 14) {real, imag} */,
  {32'h3f60d02c, 32'hbfa747bb} /* (2, 11, 13) {real, imag} */,
  {32'hbfebb5b5, 32'h40036bba} /* (2, 11, 12) {real, imag} */,
  {32'hbfde87e3, 32'hc088ccaa} /* (2, 11, 11) {real, imag} */,
  {32'h402ffe7e, 32'h3b180c4c} /* (2, 11, 10) {real, imag} */,
  {32'hc00cf8c0, 32'h4086a73a} /* (2, 11, 9) {real, imag} */,
  {32'h3ed51a4a, 32'h3faf05c1} /* (2, 11, 8) {real, imag} */,
  {32'h3e305409, 32'hbffd4f3e} /* (2, 11, 7) {real, imag} */,
  {32'h3fc02eab, 32'hbf46f7be} /* (2, 11, 6) {real, imag} */,
  {32'hbfcc48e4, 32'hbeb7c760} /* (2, 11, 5) {real, imag} */,
  {32'hbf28cb1d, 32'hbf99c103} /* (2, 11, 4) {real, imag} */,
  {32'hc059715e, 32'h40122ab5} /* (2, 11, 3) {real, imag} */,
  {32'hc1029f2a, 32'hc07d0d03} /* (2, 11, 2) {real, imag} */,
  {32'h41166d0e, 32'hbe7daeec} /* (2, 11, 1) {real, imag} */,
  {32'h4121d09a, 32'hc1115250} /* (2, 11, 0) {real, imag} */,
  {32'hc0e89c19, 32'h4014e960} /* (2, 10, 31) {real, imag} */,
  {32'h408cb370, 32'hbefde828} /* (2, 10, 30) {real, imag} */,
  {32'hbf83bf4a, 32'h40860765} /* (2, 10, 29) {real, imag} */,
  {32'h3f7eaa66, 32'h3fef38a1} /* (2, 10, 28) {real, imag} */,
  {32'h3f27d14f, 32'hc04970a9} /* (2, 10, 27) {real, imag} */,
  {32'h3fa67089, 32'h4012ed46} /* (2, 10, 26) {real, imag} */,
  {32'hbd483500, 32'hbf1892b8} /* (2, 10, 25) {real, imag} */,
  {32'h40226636, 32'hbf62f228} /* (2, 10, 24) {real, imag} */,
  {32'hc03c32e3, 32'h4006a7fd} /* (2, 10, 23) {real, imag} */,
  {32'hbdda7a25, 32'h403ec3da} /* (2, 10, 22) {real, imag} */,
  {32'hc01d897c, 32'hbfa9fcc3} /* (2, 10, 21) {real, imag} */,
  {32'hbfb4301e, 32'hbff7e4cf} /* (2, 10, 20) {real, imag} */,
  {32'h3fff0565, 32'hc004c592} /* (2, 10, 19) {real, imag} */,
  {32'h4000c9de, 32'hbf560d0f} /* (2, 10, 18) {real, imag} */,
  {32'hbffc6049, 32'h3fd17e7b} /* (2, 10, 17) {real, imag} */,
  {32'hbfd7c82d, 32'h3d7250b7} /* (2, 10, 16) {real, imag} */,
  {32'hc01b9be4, 32'hbfa3ff80} /* (2, 10, 15) {real, imag} */,
  {32'h3f34b0e5, 32'hbec45672} /* (2, 10, 14) {real, imag} */,
  {32'h40165474, 32'hbfe402ac} /* (2, 10, 13) {real, imag} */,
  {32'hc0656dbf, 32'h3f05e75c} /* (2, 10, 12) {real, imag} */,
  {32'h3e2c0539, 32'h40165883} /* (2, 10, 11) {real, imag} */,
  {32'h409eae66, 32'hbff19a02} /* (2, 10, 10) {real, imag} */,
  {32'h401789b3, 32'h4052604d} /* (2, 10, 9) {real, imag} */,
  {32'hc0199f4c, 32'h3fe61655} /* (2, 10, 8) {real, imag} */,
  {32'h3f19e2df, 32'h409b6fca} /* (2, 10, 7) {real, imag} */,
  {32'h3fd5329b, 32'hc017534f} /* (2, 10, 6) {real, imag} */,
  {32'h3be6d593, 32'h3f7fb755} /* (2, 10, 5) {real, imag} */,
  {32'hc05fddc0, 32'hbfe1eb4a} /* (2, 10, 4) {real, imag} */,
  {32'hbe5499ed, 32'hbfefe13c} /* (2, 10, 3) {real, imag} */,
  {32'h40ca3399, 32'hbf7cf704} /* (2, 10, 2) {real, imag} */,
  {32'hc055e24b, 32'h40c04817} /* (2, 10, 1) {real, imag} */,
  {32'hbfa41854, 32'h3ffee284} /* (2, 10, 0) {real, imag} */,
  {32'hc08d956f, 32'hc0fe74a5} /* (2, 9, 31) {real, imag} */,
  {32'h40daef62, 32'h40c21e1c} /* (2, 9, 30) {real, imag} */,
  {32'hc0256bd3, 32'h404505af} /* (2, 9, 29) {real, imag} */,
  {32'hbfb61e3f, 32'h3f5cc55e} /* (2, 9, 28) {real, imag} */,
  {32'h3f36d268, 32'hc0d82942} /* (2, 9, 27) {real, imag} */,
  {32'h4011be92, 32'h3f85e969} /* (2, 9, 26) {real, imag} */,
  {32'h3f862c69, 32'h3fc58c72} /* (2, 9, 25) {real, imag} */,
  {32'h400725ae, 32'hc021748e} /* (2, 9, 24) {real, imag} */,
  {32'hc01b239b, 32'h401b133e} /* (2, 9, 23) {real, imag} */,
  {32'hbef11a1d, 32'hbf3f43d8} /* (2, 9, 22) {real, imag} */,
  {32'h3e945fae, 32'hbfd5e613} /* (2, 9, 21) {real, imag} */,
  {32'h3f78b39c, 32'hc01b27c7} /* (2, 9, 20) {real, imag} */,
  {32'hbe8daafd, 32'h402c120f} /* (2, 9, 19) {real, imag} */,
  {32'h40497aa0, 32'hbfbb4ae7} /* (2, 9, 18) {real, imag} */,
  {32'h3f89dd3d, 32'hc0137581} /* (2, 9, 17) {real, imag} */,
  {32'hbf80ebe6, 32'h3f754af4} /* (2, 9, 16) {real, imag} */,
  {32'h3f2416ef, 32'h3f20d197} /* (2, 9, 15) {real, imag} */,
  {32'hc022b762, 32'h3f0320cb} /* (2, 9, 14) {real, imag} */,
  {32'h3fd913c2, 32'h3f81c364} /* (2, 9, 13) {real, imag} */,
  {32'hbf9d1d6d, 32'hbe1da932} /* (2, 9, 12) {real, imag} */,
  {32'hbfb954fa, 32'h3f68b539} /* (2, 9, 11) {real, imag} */,
  {32'hc06db83e, 32'hc03877aa} /* (2, 9, 10) {real, imag} */,
  {32'h40358163, 32'hbfa2e287} /* (2, 9, 9) {real, imag} */,
  {32'hbf18b5e1, 32'h3ece7eb5} /* (2, 9, 8) {real, imag} */,
  {32'hbfb42236, 32'hc004d0bd} /* (2, 9, 7) {real, imag} */,
  {32'h3f199939, 32'hbf0617c5} /* (2, 9, 6) {real, imag} */,
  {32'hc04c6bcd, 32'hbfc2a556} /* (2, 9, 5) {real, imag} */,
  {32'hc01d3f72, 32'hbfafa453} /* (2, 9, 4) {real, imag} */,
  {32'hbfa4ff1f, 32'hbf855fa1} /* (2, 9, 3) {real, imag} */,
  {32'h40460be4, 32'h407fc8d5} /* (2, 9, 2) {real, imag} */,
  {32'hc028eaae, 32'h40d2b6a8} /* (2, 9, 1) {real, imag} */,
  {32'h3fe6aa3a, 32'hbfa10770} /* (2, 9, 0) {real, imag} */,
  {32'h4154b7ac, 32'hc1a9e599} /* (2, 8, 31) {real, imag} */,
  {32'hc0de3753, 32'h41726839} /* (2, 8, 30) {real, imag} */,
  {32'h3ff43654, 32'hc079815b} /* (2, 8, 29) {real, imag} */,
  {32'h3d775cf6, 32'h3f67e0b4} /* (2, 8, 28) {real, imag} */,
  {32'hbf906945, 32'h401cccc6} /* (2, 8, 27) {real, imag} */,
  {32'hc08aa8c3, 32'h3f60e139} /* (2, 8, 26) {real, imag} */,
  {32'h409cf4d5, 32'h3f3138e0} /* (2, 8, 25) {real, imag} */,
  {32'hc05e7ebf, 32'h40bb1f41} /* (2, 8, 24) {real, imag} */,
  {32'h40397b0b, 32'h3f6b4a8f} /* (2, 8, 23) {real, imag} */,
  {32'hc002f45a, 32'hbf59c352} /* (2, 8, 22) {real, imag} */,
  {32'h3fc694bd, 32'h400b5e85} /* (2, 8, 21) {real, imag} */,
  {32'hbff72724, 32'h3fb2ee79} /* (2, 8, 20) {real, imag} */,
  {32'h3e9ea54d, 32'hbfbc711c} /* (2, 8, 19) {real, imag} */,
  {32'h3fd47777, 32'h3f506108} /* (2, 8, 18) {real, imag} */,
  {32'hbd30e27d, 32'h3f31edd0} /* (2, 8, 17) {real, imag} */,
  {32'hbfea807a, 32'h3fbd26e9} /* (2, 8, 16) {real, imag} */,
  {32'h3f874e11, 32'hbfc5b43c} /* (2, 8, 15) {real, imag} */,
  {32'h3f250ecc, 32'h3f59cca0} /* (2, 8, 14) {real, imag} */,
  {32'hbf662476, 32'h3d59a64b} /* (2, 8, 13) {real, imag} */,
  {32'hbfcd36b5, 32'h3eb02dd2} /* (2, 8, 12) {real, imag} */,
  {32'hc013c0dc, 32'h3f42146b} /* (2, 8, 11) {real, imag} */,
  {32'hbea13ce6, 32'h3f2268e3} /* (2, 8, 10) {real, imag} */,
  {32'h40218c45, 32'hbf9f36f7} /* (2, 8, 9) {real, imag} */,
  {32'h4056f660, 32'h3e8fb5fa} /* (2, 8, 8) {real, imag} */,
  {32'hc090ba36, 32'h400de5ba} /* (2, 8, 7) {real, imag} */,
  {32'h3bf8e284, 32'hbe6ad753} /* (2, 8, 6) {real, imag} */,
  {32'hbffa1cf2, 32'h40adffa5} /* (2, 8, 5) {real, imag} */,
  {32'h40473fe4, 32'hc0c0d3a0} /* (2, 8, 4) {real, imag} */,
  {32'hc089f15e, 32'h402564b9} /* (2, 8, 3) {real, imag} */,
  {32'hc0ad8628, 32'h40f40b15} /* (2, 8, 2) {real, imag} */,
  {32'h41289ab7, 32'hc0c029c6} /* (2, 8, 1) {real, imag} */,
  {32'h40deb631, 32'hc0a83d2b} /* (2, 8, 0) {real, imag} */,
  {32'hbf31d5e5, 32'h40d6cb0f} /* (2, 7, 31) {real, imag} */,
  {32'h408f15c2, 32'hc065677e} /* (2, 7, 30) {real, imag} */,
  {32'hbfcb3b67, 32'h3c1a4fd3} /* (2, 7, 29) {real, imag} */,
  {32'hbf8ba9ce, 32'hbeae69d9} /* (2, 7, 28) {real, imag} */,
  {32'h3fb26ac5, 32'hc027bce3} /* (2, 7, 27) {real, imag} */,
  {32'h3f02cfbb, 32'hbf682430} /* (2, 7, 26) {real, imag} */,
  {32'hc00d0b7e, 32'hbeb9f4ec} /* (2, 7, 25) {real, imag} */,
  {32'h4008b29b, 32'hbe8c398b} /* (2, 7, 24) {real, imag} */,
  {32'h408182b7, 32'h3f21fd47} /* (2, 7, 23) {real, imag} */,
  {32'hbeaa7cf2, 32'hbf8681e6} /* (2, 7, 22) {real, imag} */,
  {32'h3fb0f6f3, 32'h408eb314} /* (2, 7, 21) {real, imag} */,
  {32'hbfdfe10c, 32'hbefba5af} /* (2, 7, 20) {real, imag} */,
  {32'hbdf28afb, 32'h3fca0434} /* (2, 7, 19) {real, imag} */,
  {32'hc038e7a0, 32'hbf4912eb} /* (2, 7, 18) {real, imag} */,
  {32'h3da4052b, 32'hbf3d2c56} /* (2, 7, 17) {real, imag} */,
  {32'hbe857fd8, 32'h3f0095ee} /* (2, 7, 16) {real, imag} */,
  {32'h3fb87925, 32'h3f5959ad} /* (2, 7, 15) {real, imag} */,
  {32'hbd576c77, 32'h3fc76369} /* (2, 7, 14) {real, imag} */,
  {32'h3e45a926, 32'hbf4caef3} /* (2, 7, 13) {real, imag} */,
  {32'h3f9f5592, 32'h3f92480d} /* (2, 7, 12) {real, imag} */,
  {32'h402175b8, 32'h404ce749} /* (2, 7, 11) {real, imag} */,
  {32'h3f3c43fa, 32'h3f84fd2b} /* (2, 7, 10) {real, imag} */,
  {32'hbf5ae840, 32'hc027a841} /* (2, 7, 9) {real, imag} */,
  {32'h3f03472b, 32'hc0235838} /* (2, 7, 8) {real, imag} */,
  {32'hbec72a5c, 32'h40d30df8} /* (2, 7, 7) {real, imag} */,
  {32'hbfc98102, 32'hbef89af1} /* (2, 7, 6) {real, imag} */,
  {32'h4022c710, 32'hc04a8afc} /* (2, 7, 5) {real, imag} */,
  {32'hc00d6311, 32'hbe05ba3f} /* (2, 7, 4) {real, imag} */,
  {32'h4037e9fa, 32'hc1004d3a} /* (2, 7, 3) {real, imag} */,
  {32'h40274e72, 32'hbf530a15} /* (2, 7, 2) {real, imag} */,
  {32'hc1167e39, 32'h40a44690} /* (2, 7, 1) {real, imag} */,
  {32'hc0902899, 32'h40dbe2db} /* (2, 7, 0) {real, imag} */,
  {32'h404bb3b6, 32'h40277838} /* (2, 6, 31) {real, imag} */,
  {32'hc051de7a, 32'h40a1caec} /* (2, 6, 30) {real, imag} */,
  {32'h3f60b55b, 32'hc0179db9} /* (2, 6, 29) {real, imag} */,
  {32'hc017f02a, 32'h400ecb35} /* (2, 6, 28) {real, imag} */,
  {32'hc01e9d42, 32'hc0170f2b} /* (2, 6, 27) {real, imag} */,
  {32'hc00cb8f6, 32'h3f0ff9e0} /* (2, 6, 26) {real, imag} */,
  {32'hbef86617, 32'hbfb44006} /* (2, 6, 25) {real, imag} */,
  {32'hc03f8c37, 32'h3fd0db2f} /* (2, 6, 24) {real, imag} */,
  {32'hbf06f21d, 32'h3dff462b} /* (2, 6, 23) {real, imag} */,
  {32'h3e920a76, 32'h3f65d316} /* (2, 6, 22) {real, imag} */,
  {32'hc006ebfd, 32'h40142b5a} /* (2, 6, 21) {real, imag} */,
  {32'hbf15bcf3, 32'h3fbf2ee7} /* (2, 6, 20) {real, imag} */,
  {32'h3fb8331e, 32'hbe67160f} /* (2, 6, 19) {real, imag} */,
  {32'h3ead0d58, 32'hbe52d7f9} /* (2, 6, 18) {real, imag} */,
  {32'h3e6907f6, 32'hbf259052} /* (2, 6, 17) {real, imag} */,
  {32'hbf606ef8, 32'h3ecd8e21} /* (2, 6, 16) {real, imag} */,
  {32'h3f1625de, 32'h3e80581e} /* (2, 6, 15) {real, imag} */,
  {32'h3f267245, 32'hbfdefdf0} /* (2, 6, 14) {real, imag} */,
  {32'hc037e0fd, 32'h3f7c8ae1} /* (2, 6, 13) {real, imag} */,
  {32'h3f346531, 32'hbf9fd1fa} /* (2, 6, 12) {real, imag} */,
  {32'hbf3c6d95, 32'h3ff9dc8c} /* (2, 6, 11) {real, imag} */,
  {32'h3e9df42b, 32'hc08041fe} /* (2, 6, 10) {real, imag} */,
  {32'h4012321f, 32'h3fd9d84b} /* (2, 6, 9) {real, imag} */,
  {32'hbfe1e2a0, 32'h40707d6f} /* (2, 6, 8) {real, imag} */,
  {32'h3ffad705, 32'hbf785683} /* (2, 6, 7) {real, imag} */,
  {32'hc029fed6, 32'h40365bf5} /* (2, 6, 6) {real, imag} */,
  {32'h3fa1cc06, 32'h3ff49ab2} /* (2, 6, 5) {real, imag} */,
  {32'h3f539fc9, 32'h3fd635a2} /* (2, 6, 4) {real, imag} */,
  {32'hc080c0d5, 32'h402c802b} /* (2, 6, 3) {real, imag} */,
  {32'h409c197e, 32'h4101e3d7} /* (2, 6, 2) {real, imag} */,
  {32'h40238bd0, 32'hc0626806} /* (2, 6, 1) {real, imag} */,
  {32'hc06274b9, 32'hc0494e40} /* (2, 6, 0) {real, imag} */,
  {32'h4184c940, 32'hc22cd933} /* (2, 5, 31) {real, imag} */,
  {32'hc07ca3ca, 32'h4178ce92} /* (2, 5, 30) {real, imag} */,
  {32'hbf7a62fd, 32'h40a326cb} /* (2, 5, 29) {real, imag} */,
  {32'hc0d86bdf, 32'hc0a1507a} /* (2, 5, 28) {real, imag} */,
  {32'h408db01e, 32'h41309096} /* (2, 5, 27) {real, imag} */,
  {32'h4023dbed, 32'h3fa1c822} /* (2, 5, 26) {real, imag} */,
  {32'hbfaabacc, 32'hbdecf768} /* (2, 5, 25) {real, imag} */,
  {32'h40062f23, 32'h408db10c} /* (2, 5, 24) {real, imag} */,
  {32'hc0044ac7, 32'hbf1fd613} /* (2, 5, 23) {real, imag} */,
  {32'h3fbe7311, 32'h40575d63} /* (2, 5, 22) {real, imag} */,
  {32'h3f728b52, 32'h40cd0e8d} /* (2, 5, 21) {real, imag} */,
  {32'hbfb33d31, 32'h3dfcf8d0} /* (2, 5, 20) {real, imag} */,
  {32'hbfd83f11, 32'hbf04cc68} /* (2, 5, 19) {real, imag} */,
  {32'h4030b8aa, 32'h401527bd} /* (2, 5, 18) {real, imag} */,
  {32'h4004d570, 32'h3ed95fef} /* (2, 5, 17) {real, imag} */,
  {32'h3ece6f24, 32'h3e83ad69} /* (2, 5, 16) {real, imag} */,
  {32'hbfc1c7bd, 32'hbfbd16c8} /* (2, 5, 15) {real, imag} */,
  {32'hbfa2d2ee, 32'hc00c3b95} /* (2, 5, 14) {real, imag} */,
  {32'h3fa781d6, 32'hbf916e84} /* (2, 5, 13) {real, imag} */,
  {32'hbfc6e97a, 32'h40395d3a} /* (2, 5, 12) {real, imag} */,
  {32'hc09a86b1, 32'h3f6f4cd9} /* (2, 5, 11) {real, imag} */,
  {32'hbe846cea, 32'hc042ae19} /* (2, 5, 10) {real, imag} */,
  {32'h3f38bee6, 32'h4008e1d3} /* (2, 5, 9) {real, imag} */,
  {32'hc09eda4b, 32'h403a9c8b} /* (2, 5, 8) {real, imag} */,
  {32'h401d0abf, 32'h3e1539b8} /* (2, 5, 7) {real, imag} */,
  {32'hc04d3532, 32'hc087f054} /* (2, 5, 6) {real, imag} */,
  {32'hc178083c, 32'h41528df3} /* (2, 5, 5) {real, imag} */,
  {32'h40d0eb07, 32'hc09d4fcb} /* (2, 5, 4) {real, imag} */,
  {32'h407f3888, 32'hbfbd380d} /* (2, 5, 3) {real, imag} */,
  {32'hc1032788, 32'h4066c6c3} /* (2, 5, 2) {real, imag} */,
  {32'h41e55b7c, 32'hc1d6dbc5} /* (2, 5, 1) {real, imag} */,
  {32'h419be0a5, 32'hc1f47949} /* (2, 5, 0) {real, imag} */,
  {32'hc22100bd, 32'h4158cb75} /* (2, 4, 31) {real, imag} */,
  {32'h42056b8e, 32'hc1d47a65} /* (2, 4, 30) {real, imag} */,
  {32'h3f0dc41a, 32'hbfca41d4} /* (2, 4, 29) {real, imag} */,
  {32'hc08bf3ec, 32'h4186f7d9} /* (2, 4, 28) {real, imag} */,
  {32'hc0437c1f, 32'hc103c120} /* (2, 4, 27) {real, imag} */,
  {32'hc0b1319c, 32'h4063b132} /* (2, 4, 26) {real, imag} */,
  {32'hc02834fd, 32'h3e561384} /* (2, 4, 25) {real, imag} */,
  {32'hbe74efa5, 32'hc09558ab} /* (2, 4, 24) {real, imag} */,
  {32'hc0436d89, 32'h402f2b8f} /* (2, 4, 23) {real, imag} */,
  {32'h3fc5ff71, 32'h40763dec} /* (2, 4, 22) {real, imag} */,
  {32'hc057ea9f, 32'hc0e54ae2} /* (2, 4, 21) {real, imag} */,
  {32'h3fea8b98, 32'hbf08cd6d} /* (2, 4, 20) {real, imag} */,
  {32'h3ce79ce5, 32'hbdbfd9d3} /* (2, 4, 19) {real, imag} */,
  {32'h3f199c76, 32'hbf0d89cf} /* (2, 4, 18) {real, imag} */,
  {32'hc032094c, 32'h3eab797b} /* (2, 4, 17) {real, imag} */,
  {32'h3f61ed2b, 32'hbf6bc1da} /* (2, 4, 16) {real, imag} */,
  {32'h3f8217db, 32'hbfbee9ee} /* (2, 4, 15) {real, imag} */,
  {32'h3ff2fbc1, 32'h3e3c0b9e} /* (2, 4, 14) {real, imag} */,
  {32'h3e8edc62, 32'h3fce630c} /* (2, 4, 13) {real, imag} */,
  {32'h40780b6c, 32'hc002b7bc} /* (2, 4, 12) {real, imag} */,
  {32'hbdf5a8a0, 32'hbe33810d} /* (2, 4, 11) {real, imag} */,
  {32'hc026b2c3, 32'hbfde8d7e} /* (2, 4, 10) {real, imag} */,
  {32'h3f8da545, 32'h3ecb32f8} /* (2, 4, 9) {real, imag} */,
  {32'h40bdeeae, 32'h3e113cdc} /* (2, 4, 8) {real, imag} */,
  {32'hbea03c27, 32'h405d341d} /* (2, 4, 7) {real, imag} */,
  {32'h3e138acb, 32'hc02ea893} /* (2, 4, 6) {real, imag} */,
  {32'h40f80ab1, 32'h402964dd} /* (2, 4, 5) {real, imag} */,
  {32'hc13891ad, 32'h40c41e17} /* (2, 4, 4) {real, imag} */,
  {32'hc01e7dd8, 32'h40d147ee} /* (2, 4, 3) {real, imag} */,
  {32'h4223e130, 32'hc1e534a5} /* (2, 4, 2) {real, imag} */,
  {32'hc2029c05, 32'h428c1420} /* (2, 4, 1) {real, imag} */,
  {32'hc0e6cae1, 32'h4164deb8} /* (2, 4, 0) {real, imag} */,
  {32'hc1882d18, 32'hc286fa98} /* (2, 3, 31) {real, imag} */,
  {32'h4231fed4, 32'h42705097} /* (2, 3, 30) {real, imag} */,
  {32'hc0b1d76b, 32'hbed3156f} /* (2, 3, 29) {real, imag} */,
  {32'hc168e66a, 32'h4177c4a0} /* (2, 3, 28) {real, imag} */,
  {32'h40222ddc, 32'hc13a6e7c} /* (2, 3, 27) {real, imag} */,
  {32'hc096839a, 32'h3f5ae6e3} /* (2, 3, 26) {real, imag} */,
  {32'hbdf0c3e7, 32'h40a249d9} /* (2, 3, 25) {real, imag} */,
  {32'h40aba62d, 32'h3db8d9c4} /* (2, 3, 24) {real, imag} */,
  {32'hc0aadeca, 32'h400b87e7} /* (2, 3, 23) {real, imag} */,
  {32'hc0a91d20, 32'h401148db} /* (2, 3, 22) {real, imag} */,
  {32'hbfc7d9f5, 32'hc06de4f2} /* (2, 3, 21) {real, imag} */,
  {32'hbf3c9cc2, 32'hbf177697} /* (2, 3, 20) {real, imag} */,
  {32'hbeb58590, 32'hc003fffc} /* (2, 3, 19) {real, imag} */,
  {32'hbea1592c, 32'h3e2f88b1} /* (2, 3, 18) {real, imag} */,
  {32'hbd35b7e3, 32'hbf2cd7fc} /* (2, 3, 17) {real, imag} */,
  {32'hc00e7b81, 32'h3e2a1814} /* (2, 3, 16) {real, imag} */,
  {32'h3e95bfb2, 32'hbe0f53a6} /* (2, 3, 15) {real, imag} */,
  {32'h403c6233, 32'h3f0d8472} /* (2, 3, 14) {real, imag} */,
  {32'h3fa44cbe, 32'h3f24fe37} /* (2, 3, 13) {real, imag} */,
  {32'h3f3c8752, 32'h3f0ee040} /* (2, 3, 12) {real, imag} */,
  {32'hbfe1a2cc, 32'h4091394e} /* (2, 3, 11) {real, imag} */,
  {32'h4025c4f6, 32'hc08c9c69} /* (2, 3, 10) {real, imag} */,
  {32'hbfae8848, 32'hc01bd7e2} /* (2, 3, 9) {real, imag} */,
  {32'h40b0cbef, 32'hbf668333} /* (2, 3, 8) {real, imag} */,
  {32'hc0071bfc, 32'h401f9fa9} /* (2, 3, 7) {real, imag} */,
  {32'hc06a24fb, 32'hc0ab177a} /* (2, 3, 6) {real, imag} */,
  {32'hc0ee4e4f, 32'h4128e4bb} /* (2, 3, 5) {real, imag} */,
  {32'hc0022452, 32'hc04c88ea} /* (2, 3, 4) {real, imag} */,
  {32'hbfe61e01, 32'hc0f037cf} /* (2, 3, 3) {real, imag} */,
  {32'h4267b321, 32'h3f6fec37} /* (2, 3, 2) {real, imag} */,
  {32'hc236ad6f, 32'h41ec813b} /* (2, 3, 1) {real, imag} */,
  {32'hc0d00007, 32'hc0591057} /* (2, 3, 0) {real, imag} */,
  {32'h42e44b9b, 32'hc3e66b07} /* (2, 2, 31) {real, imag} */,
  {32'h41b0175f, 32'h43675454} /* (2, 2, 30) {real, imag} */,
  {32'h413993e9, 32'hc02f159a} /* (2, 2, 29) {real, imag} */,
  {32'hc2144f00, 32'hc19ebd67} /* (2, 2, 28) {real, imag} */,
  {32'h4115c006, 32'h421209b1} /* (2, 2, 27) {real, imag} */,
  {32'h400fa093, 32'h4106bdf4} /* (2, 2, 26) {real, imag} */,
  {32'hc123b7aa, 32'hc13e340a} /* (2, 2, 25) {real, imag} */,
  {32'h411c647d, 32'h40f24b1f} /* (2, 2, 24) {real, imag} */,
  {32'hc0629fca, 32'h401dc65f} /* (2, 2, 23) {real, imag} */,
  {32'hbfb2b7f5, 32'h3e2f4c53} /* (2, 2, 22) {real, imag} */,
  {32'h40d793ef, 32'h40cf1038} /* (2, 2, 21) {real, imag} */,
  {32'hc02f2d66, 32'hc044eadf} /* (2, 2, 20) {real, imag} */,
  {32'hbfa333ba, 32'h3e5b3062} /* (2, 2, 19) {real, imag} */,
  {32'h404b2c9a, 32'h403714ee} /* (2, 2, 18) {real, imag} */,
  {32'hc02a7867, 32'h3d21f263} /* (2, 2, 17) {real, imag} */,
  {32'h3f027bee, 32'hbf9f59a4} /* (2, 2, 16) {real, imag} */,
  {32'hbeb622ac, 32'hc029f31c} /* (2, 2, 15) {real, imag} */,
  {32'hc07e05c3, 32'h3f055f9c} /* (2, 2, 14) {real, imag} */,
  {32'h3e850304, 32'h3d7b589b} /* (2, 2, 13) {real, imag} */,
  {32'h3f2b1183, 32'h3f54a96f} /* (2, 2, 12) {real, imag} */,
  {32'hc0f430c6, 32'h3ff0ecf6} /* (2, 2, 11) {real, imag} */,
  {32'h4001e860, 32'hc080d7d0} /* (2, 2, 10) {real, imag} */,
  {32'hbf71539b, 32'hc02f79f4} /* (2, 2, 9) {real, imag} */,
  {32'hc0f6d6f1, 32'h40bf46f4} /* (2, 2, 8) {real, imag} */,
  {32'h3f1c0eb5, 32'hc082a530} /* (2, 2, 7) {real, imag} */,
  {32'hbfe854dd, 32'h408d9de9} /* (2, 2, 6) {real, imag} */,
  {32'hc20a4c56, 32'h41863c08} /* (2, 2, 5) {real, imag} */,
  {32'h420753db, 32'hc240b24b} /* (2, 2, 4) {real, imag} */,
  {32'h40a3258e, 32'hc08fdef4} /* (2, 2, 3) {real, imag} */,
  {32'h41508195, 32'h43389c33} /* (2, 2, 2) {real, imag} */,
  {32'hc06c0445, 32'hc38e9193} /* (2, 2, 1) {real, imag} */,
  {32'h42a9df32, 32'hc34c8af2} /* (2, 2, 0) {real, imag} */,
  {32'h41c4e950, 32'h44068a5c} /* (2, 1, 31) {real, imag} */,
  {32'h4182779c, 32'hc33b15b1} /* (2, 1, 30) {real, imag} */,
  {32'hc18b5e36, 32'h3ef0691d} /* (2, 1, 29) {real, imag} */,
  {32'hc1ef9c2f, 32'h41a61ab4} /* (2, 1, 28) {real, imag} */,
  {32'h4140e774, 32'hc24ccf86} /* (2, 1, 27) {real, imag} */,
  {32'h40cd96a8, 32'hc12d74c5} /* (2, 1, 26) {real, imag} */,
  {32'h40393b16, 32'h40fa62ca} /* (2, 1, 25) {real, imag} */,
  {32'hc0a7e4eb, 32'hc0f9ef3a} /* (2, 1, 24) {real, imag} */,
  {32'hc0d06433, 32'hc0a1773a} /* (2, 1, 23) {real, imag} */,
  {32'hc076eec8, 32'h403ea4ce} /* (2, 1, 22) {real, imag} */,
  {32'hc01b7283, 32'hc128e89c} /* (2, 1, 21) {real, imag} */,
  {32'hbf91004d, 32'h3e975261} /* (2, 1, 20) {real, imag} */,
  {32'hbf8d1f42, 32'h3fe3a8a2} /* (2, 1, 19) {real, imag} */,
  {32'hc07d6086, 32'hbcee3d61} /* (2, 1, 18) {real, imag} */,
  {32'hbc8e9d8b, 32'hbeb72f54} /* (2, 1, 17) {real, imag} */,
  {32'hbf83b9c4, 32'hbc452f02} /* (2, 1, 16) {real, imag} */,
  {32'hbec74663, 32'hbfb32487} /* (2, 1, 15) {real, imag} */,
  {32'h4089e5d6, 32'h402b9ee3} /* (2, 1, 14) {real, imag} */,
  {32'hbffeae5d, 32'h4092e7f4} /* (2, 1, 13) {real, imag} */,
  {32'h4023af26, 32'h3db2de06} /* (2, 1, 12) {real, imag} */,
  {32'h40d4e124, 32'hbf2db7d1} /* (2, 1, 11) {real, imag} */,
  {32'h40972715, 32'hc05577cd} /* (2, 1, 10) {real, imag} */,
  {32'h3e8c5ffe, 32'h3f251469} /* (2, 1, 9) {real, imag} */,
  {32'h4195e005, 32'hc0258639} /* (2, 1, 8) {real, imag} */,
  {32'hc10a7bb7, 32'h40660183} /* (2, 1, 7) {real, imag} */,
  {32'h40b49222, 32'hbf0ef6cc} /* (2, 1, 6) {real, imag} */,
  {32'h41deaa82, 32'hc1ed0171} /* (2, 1, 5) {real, imag} */,
  {32'hc1f3bc94, 32'h4171ecc8} /* (2, 1, 4) {real, imag} */,
  {32'hc15e74e7, 32'hc15d584f} /* (2, 1, 3) {real, imag} */,
  {32'h438094da, 32'hc3321858} /* (2, 1, 2) {real, imag} */,
  {32'hc4101db2, 32'h44259730} /* (2, 1, 1) {real, imag} */,
  {32'hc3392074, 32'h440d4f55} /* (2, 1, 0) {real, imag} */,
  {32'h43625fb0, 32'h43ddd790} /* (2, 0, 31) {real, imag} */,
  {32'hc2dd8506, 32'hc2c375da} /* (2, 0, 30) {real, imag} */,
  {32'h3f6de1f0, 32'hc18b0cfa} /* (2, 0, 29) {real, imag} */,
  {32'hc1fcdbb5, 32'h3fe29442} /* (2, 0, 28) {real, imag} */,
  {32'h40a57bae, 32'hc1e2251c} /* (2, 0, 27) {real, imag} */,
  {32'hbf925047, 32'hc0b5e02c} /* (2, 0, 26) {real, imag} */,
  {32'h4048b250, 32'h401dd484} /* (2, 0, 25) {real, imag} */,
  {32'hc10566f5, 32'hbf0b4d1d} /* (2, 0, 24) {real, imag} */,
  {32'h3e9bea89, 32'hc0538dc6} /* (2, 0, 23) {real, imag} */,
  {32'hbfadbb07, 32'hc04d6fa9} /* (2, 0, 22) {real, imag} */,
  {32'hbf4a8bc6, 32'hc05b4cde} /* (2, 0, 21) {real, imag} */,
  {32'h407182b2, 32'h40956e94} /* (2, 0, 20) {real, imag} */,
  {32'h3ff47b1d, 32'hbf723380} /* (2, 0, 19) {real, imag} */,
  {32'hbf6fa3d0, 32'hbe38170d} /* (2, 0, 18) {real, imag} */,
  {32'h3f98a979, 32'h3fddf0aa} /* (2, 0, 17) {real, imag} */,
  {32'hbf22ff31, 32'hbf595a4f} /* (2, 0, 16) {real, imag} */,
  {32'h3f2b66b0, 32'h3e88768f} /* (2, 0, 15) {real, imag} */,
  {32'hbf513d6f, 32'h3f1e8120} /* (2, 0, 14) {real, imag} */,
  {32'hc01b6059, 32'hc0158a47} /* (2, 0, 13) {real, imag} */,
  {32'h400e87a5, 32'hbfa5e5d4} /* (2, 0, 12) {real, imag} */,
  {32'h404f99ba, 32'h3e829f24} /* (2, 0, 11) {real, imag} */,
  {32'h40200834, 32'h400fe783} /* (2, 0, 10) {real, imag} */,
  {32'h3fd1e90f, 32'hc085a126} /* (2, 0, 9) {real, imag} */,
  {32'h414aaaf1, 32'h4010aea1} /* (2, 0, 8) {real, imag} */,
  {32'hc1802800, 32'hc03ca201} /* (2, 0, 7) {real, imag} */,
  {32'hc09510c4, 32'hc0338645} /* (2, 0, 6) {real, imag} */,
  {32'h40a975c8, 32'hc1d4565e} /* (2, 0, 5) {real, imag} */,
  {32'h4155c923, 32'hbfcb0799} /* (2, 0, 4) {real, imag} */,
  {32'h415f0961, 32'hc19a76a0} /* (2, 0, 3) {real, imag} */,
  {32'h42eeccbe, 32'hc229bd12} /* (2, 0, 2) {real, imag} */,
  {32'hc3c36af0, 32'h43a7593f} /* (2, 0, 1) {real, imag} */,
  {32'hc2d25a25, 32'h43eb6535} /* (2, 0, 0) {real, imag} */,
  {32'hc3aa13d4, 32'hc44b82a2} /* (1, 31, 31) {real, imag} */,
  {32'h431af7b3, 32'h43604a4c} /* (1, 31, 30) {real, imag} */,
  {32'h4199b3d9, 32'h411cdff7} /* (1, 31, 29) {real, imag} */,
  {32'h40710768, 32'hc0b73d3c} /* (1, 31, 28) {real, imag} */,
  {32'h40b8e41b, 32'h41bde69e} /* (1, 31, 27) {real, imag} */,
  {32'h4033a287, 32'h40563815} /* (1, 31, 26) {real, imag} */,
  {32'hc0f30270, 32'hc109ff6e} /* (1, 31, 25) {real, imag} */,
  {32'h411ba76c, 32'h40e0464c} /* (1, 31, 24) {real, imag} */,
  {32'hc079e560, 32'h3ffce1a2} /* (1, 31, 23) {real, imag} */,
  {32'h3f890c71, 32'h3cf948e1} /* (1, 31, 22) {real, imag} */,
  {32'h40c7ea4c, 32'h40658ced} /* (1, 31, 21) {real, imag} */,
  {32'h40644c9e, 32'hbfdf108e} /* (1, 31, 20) {real, imag} */,
  {32'h3f567d6d, 32'hbf0f7361} /* (1, 31, 19) {real, imag} */,
  {32'h400b8735, 32'h3ff3a28a} /* (1, 31, 18) {real, imag} */,
  {32'hbf694cc0, 32'hbf5228da} /* (1, 31, 17) {real, imag} */,
  {32'hbfb0b248, 32'hbe97b39a} /* (1, 31, 16) {real, imag} */,
  {32'hbe2dce92, 32'h3eb0c51c} /* (1, 31, 15) {real, imag} */,
  {32'hc09b8aef, 32'h402bf1ce} /* (1, 31, 14) {real, imag} */,
  {32'hbf8a6cf8, 32'h3febc496} /* (1, 31, 13) {real, imag} */,
  {32'h402fa83a, 32'hc009ea39} /* (1, 31, 12) {real, imag} */,
  {32'hc0569840, 32'h40b538bc} /* (1, 31, 11) {real, imag} */,
  {32'hc0ca7963, 32'h3dd5e25f} /* (1, 31, 10) {real, imag} */,
  {32'hbf5fd1f8, 32'h4052c65b} /* (1, 31, 9) {real, imag} */,
  {32'h3dd47b1f, 32'h40924b6c} /* (1, 31, 8) {real, imag} */,
  {32'h3f2b8969, 32'h4080824f} /* (1, 31, 7) {real, imag} */,
  {32'hc124507e, 32'hc00cf5e9} /* (1, 31, 6) {real, imag} */,
  {32'hc075fc07, 32'h41ea5854} /* (1, 31, 5) {real, imag} */,
  {32'hc19fbc62, 32'hc20de9c4} /* (1, 31, 4) {real, imag} */,
  {32'h409e9d0a, 32'h40f53094} /* (1, 31, 3) {real, imag} */,
  {32'hc11b89ec, 32'h42e5de86} /* (1, 31, 2) {real, imag} */,
  {32'h4344c965, 32'hc407fd22} /* (1, 31, 1) {real, imag} */,
  {32'hc1c9a61e, 32'hc4599db9} /* (1, 31, 0) {real, imag} */,
  {32'hc28ed767, 32'h433e6304} /* (1, 30, 31) {real, imag} */,
  {32'h4214d5ee, 32'hc2f14415} /* (1, 30, 30) {real, imag} */,
  {32'hc1b29041, 32'h40c0787d} /* (1, 30, 29) {real, imag} */,
  {32'h40997199, 32'h4191f598} /* (1, 30, 28) {real, imag} */,
  {32'hc138aa0b, 32'hc1a988e3} /* (1, 30, 27) {real, imag} */,
  {32'hc00efc93, 32'h403166a0} /* (1, 30, 26) {real, imag} */,
  {32'h409c2598, 32'h4059de92} /* (1, 30, 25) {real, imag} */,
  {32'hc0c4a3b8, 32'hc11381e9} /* (1, 30, 24) {real, imag} */,
  {32'hbf300945, 32'h3f1966f0} /* (1, 30, 23) {real, imag} */,
  {32'h3f72c956, 32'h3fec808d} /* (1, 30, 22) {real, imag} */,
  {32'hc08e23c1, 32'hc01c2de0} /* (1, 30, 21) {real, imag} */,
  {32'h3e2d14dd, 32'hbf6a9b87} /* (1, 30, 20) {real, imag} */,
  {32'hbe921cb7, 32'h4013b4f0} /* (1, 30, 19) {real, imag} */,
  {32'hbe4ceadd, 32'h3ed984e4} /* (1, 30, 18) {real, imag} */,
  {32'h3f22aa12, 32'h3f7b38cc} /* (1, 30, 17) {real, imag} */,
  {32'h3f46cfb2, 32'hbf59ea01} /* (1, 30, 16) {real, imag} */,
  {32'h3e4ca095, 32'hbf8a50e5} /* (1, 30, 15) {real, imag} */,
  {32'h4006ab3e, 32'h3f2c8dd2} /* (1, 30, 14) {real, imag} */,
  {32'h40125f90, 32'h3f9ba7e8} /* (1, 30, 13) {real, imag} */,
  {32'h3ed309c2, 32'hc00e74a5} /* (1, 30, 12) {real, imag} */,
  {32'h3f074bd4, 32'h3fa03e0e} /* (1, 30, 11) {real, imag} */,
  {32'hbe41a295, 32'h3f745af2} /* (1, 30, 10) {real, imag} */,
  {32'h3ed092ea, 32'h40962649} /* (1, 30, 9) {real, imag} */,
  {32'h40d7a494, 32'hc1013c1b} /* (1, 30, 8) {real, imag} */,
  {32'h3faa2123, 32'hbf9e8617} /* (1, 30, 7) {real, imag} */,
  {32'h4066d6b6, 32'hc0842024} /* (1, 30, 6) {real, imag} */,
  {32'h41248f9c, 32'hc18cce9a} /* (1, 30, 5) {real, imag} */,
  {32'hc19bc397, 32'h4021b15a} /* (1, 30, 4) {real, imag} */,
  {32'hc1b2542c, 32'h41032ab9} /* (1, 30, 3) {real, imag} */,
  {32'h42967d5a, 32'hc32231dd} /* (1, 30, 2) {real, imag} */,
  {32'hc1d1658e, 32'h43be0ad6} /* (1, 30, 1) {real, imag} */,
  {32'h41042068, 32'h43624196} /* (1, 30, 0) {real, imag} */,
  {32'hc1fd1b4e, 32'hc27592a6} /* (1, 29, 31) {real, imag} */,
  {32'h41991450, 32'hbeb04014} /* (1, 29, 30) {real, imag} */,
  {32'hc0afe47e, 32'h41499d63} /* (1, 29, 29) {real, imag} */,
  {32'hc0824e77, 32'h411d1293} /* (1, 29, 28) {real, imag} */,
  {32'hc0c8180d, 32'hbff635ec} /* (1, 29, 27) {real, imag} */,
  {32'hc04fd972, 32'h3f03e6bd} /* (1, 29, 26) {real, imag} */,
  {32'h40512162, 32'h4027c274} /* (1, 29, 25) {real, imag} */,
  {32'hc00adf51, 32'hbfb08c70} /* (1, 29, 24) {real, imag} */,
  {32'h40449654, 32'hc07082b6} /* (1, 29, 23) {real, imag} */,
  {32'hbf6d8af1, 32'h400f2aee} /* (1, 29, 22) {real, imag} */,
  {32'hbf359e7c, 32'h3fe4a69f} /* (1, 29, 21) {real, imag} */,
  {32'h3f7821e0, 32'hbe82d4c7} /* (1, 29, 20) {real, imag} */,
  {32'hbeae5878, 32'h3edbc459} /* (1, 29, 19) {real, imag} */,
  {32'h3ffac8d9, 32'hc0a8032a} /* (1, 29, 18) {real, imag} */,
  {32'hbe9736fd, 32'h3f72194d} /* (1, 29, 17) {real, imag} */,
  {32'hbf0b18cc, 32'h400b49d0} /* (1, 29, 16) {real, imag} */,
  {32'hbdd3a65f, 32'h3e82cdb3} /* (1, 29, 15) {real, imag} */,
  {32'h3f5252d7, 32'h4006bde9} /* (1, 29, 14) {real, imag} */,
  {32'hbf2340ad, 32'hc0076875} /* (1, 29, 13) {real, imag} */,
  {32'hc006d944, 32'hbde46237} /* (1, 29, 12) {real, imag} */,
  {32'hbf9c2d66, 32'hbe89aaad} /* (1, 29, 11) {real, imag} */,
  {32'h4039d039, 32'hc034e648} /* (1, 29, 10) {real, imag} */,
  {32'h3fd15431, 32'h3f6ba67a} /* (1, 29, 9) {real, imag} */,
  {32'h3f7be866, 32'hc0863b2b} /* (1, 29, 8) {real, imag} */,
  {32'hbfe349ad, 32'h3f9b4af4} /* (1, 29, 7) {real, imag} */,
  {32'hbf2a284e, 32'h40169c76} /* (1, 29, 6) {real, imag} */,
  {32'hbf7a25c9, 32'h412c52a2} /* (1, 29, 5) {real, imag} */,
  {32'hc0fbe03a, 32'hc1649e61} /* (1, 29, 4) {real, imag} */,
  {32'h40b5caa4, 32'h40271096} /* (1, 29, 3) {real, imag} */,
  {32'h4232533d, 32'hbea2e905} /* (1, 29, 2) {real, imag} */,
  {32'hc1dcd3c0, 32'h41e98d21} /* (1, 29, 1) {real, imag} */,
  {32'h4090b3f6, 32'h414b4f84} /* (1, 29, 0) {real, imag} */,
  {32'hc1a40cb3, 32'hc24b03c4} /* (1, 28, 31) {real, imag} */,
  {32'h416296ad, 32'h41e646ec} /* (1, 28, 30) {real, imag} */,
  {32'hc0f1dc53, 32'hbd2c52e7} /* (1, 28, 29) {real, imag} */,
  {32'hc14baf62, 32'h40bf47f6} /* (1, 28, 28) {real, imag} */,
  {32'h412cd2c8, 32'h405fd2a8} /* (1, 28, 27) {real, imag} */,
  {32'h408835b6, 32'hc04c9d00} /* (1, 28, 26) {real, imag} */,
  {32'h4028620d, 32'hc06a9dd5} /* (1, 28, 25) {real, imag} */,
  {32'h40334fcb, 32'hbe91bf1f} /* (1, 28, 24) {real, imag} */,
  {32'hbd2faf67, 32'hbf6259d6} /* (1, 28, 23) {real, imag} */,
  {32'hbf4cdf4c, 32'h3f0d5328} /* (1, 28, 22) {real, imag} */,
  {32'h409ee958, 32'hc0573855} /* (1, 28, 21) {real, imag} */,
  {32'hc04adafa, 32'h3fd3cb34} /* (1, 28, 20) {real, imag} */,
  {32'h3fc18595, 32'h3f676f87} /* (1, 28, 19) {real, imag} */,
  {32'h4009636c, 32'hc043b2ba} /* (1, 28, 18) {real, imag} */,
  {32'hbffd382e, 32'h3e076b7d} /* (1, 28, 17) {real, imag} */,
  {32'hbd311964, 32'hbe9a6b5c} /* (1, 28, 16) {real, imag} */,
  {32'h3f63682b, 32'h3deb48e5} /* (1, 28, 15) {real, imag} */,
  {32'h3f423fa8, 32'h3fa52da9} /* (1, 28, 14) {real, imag} */,
  {32'hbe74f736, 32'hbd95eefc} /* (1, 28, 13) {real, imag} */,
  {32'hbf83541f, 32'hbe79f3df} /* (1, 28, 12) {real, imag} */,
  {32'h4038f6a4, 32'hbfc26fbb} /* (1, 28, 11) {real, imag} */,
  {32'h4053fbf8, 32'h3f236671} /* (1, 28, 10) {real, imag} */,
  {32'hbfbde391, 32'hc04c37b0} /* (1, 28, 9) {real, imag} */,
  {32'hbed370e1, 32'h404699dc} /* (1, 28, 8) {real, imag} */,
  {32'hbf449144, 32'h4013b834} /* (1, 28, 7) {real, imag} */,
  {32'h3eaed6ac, 32'h4088a1b8} /* (1, 28, 6) {real, imag} */,
  {32'hc04a9d28, 32'h4033df8d} /* (1, 28, 5) {real, imag} */,
  {32'hbf941fb1, 32'hc110a117} /* (1, 28, 4) {real, imag} */,
  {32'hbf7ec318, 32'hc0ce076f} /* (1, 28, 3) {real, imag} */,
  {32'h41962fc0, 32'h4198500d} /* (1, 28, 2) {real, imag} */,
  {32'hc1ffdd89, 32'hc19af120} /* (1, 28, 1) {real, imag} */,
  {32'h41591b99, 32'hc1c60966} /* (1, 28, 0) {real, imag} */,
  {32'h41b323c8, 32'h41694fe3} /* (1, 27, 31) {real, imag} */,
  {32'hc149838f, 32'hc12e51e9} /* (1, 27, 30) {real, imag} */,
  {32'hc09b04c9, 32'h4096f027} /* (1, 27, 29) {real, imag} */,
  {32'h4078abcb, 32'h3f247139} /* (1, 27, 28) {real, imag} */,
  {32'hc02d4540, 32'hbfe3e8c9} /* (1, 27, 27) {real, imag} */,
  {32'hbfc9a6d9, 32'h3ad4afe7} /* (1, 27, 26) {real, imag} */,
  {32'h3f81447a, 32'h40c2487e} /* (1, 27, 25) {real, imag} */,
  {32'hc00cbfa6, 32'h3fd4ce88} /* (1, 27, 24) {real, imag} */,
  {32'hbfe1144a, 32'hc04f1cc2} /* (1, 27, 23) {real, imag} */,
  {32'hc0251677, 32'h3f08976c} /* (1, 27, 22) {real, imag} */,
  {32'hc0859cf4, 32'hbf95e244} /* (1, 27, 21) {real, imag} */,
  {32'hbfec6c1f, 32'hc043077e} /* (1, 27, 20) {real, imag} */,
  {32'h3edcbdcc, 32'hbfd8b700} /* (1, 27, 19) {real, imag} */,
  {32'hbfaf1175, 32'h3facdc48} /* (1, 27, 18) {real, imag} */,
  {32'h3d2fbc86, 32'hbe96f1f1} /* (1, 27, 17) {real, imag} */,
  {32'hbb1f4c75, 32'hbf0aa8da} /* (1, 27, 16) {real, imag} */,
  {32'hbfec6098, 32'h3b9fb68b} /* (1, 27, 15) {real, imag} */,
  {32'h3f18c3a2, 32'h3f8ffebb} /* (1, 27, 14) {real, imag} */,
  {32'h3edd3926, 32'h3f01fc3a} /* (1, 27, 13) {real, imag} */,
  {32'h3fe3c4f1, 32'h4058b754} /* (1, 27, 12) {real, imag} */,
  {32'hbee9e59a, 32'hbffd3401} /* (1, 27, 11) {real, imag} */,
  {32'h3f00bc85, 32'hbea48cfa} /* (1, 27, 10) {real, imag} */,
  {32'hbf4e4e91, 32'h3fb49a44} /* (1, 27, 9) {real, imag} */,
  {32'h40839c46, 32'hc08521e5} /* (1, 27, 8) {real, imag} */,
  {32'hc01607b3, 32'hbf8c333d} /* (1, 27, 7) {real, imag} */,
  {32'hbeb9ae1c, 32'h404ac8c2} /* (1, 27, 6) {real, imag} */,
  {32'hbfc9c2ad, 32'hc02d131a} /* (1, 27, 5) {real, imag} */,
  {32'h3fc77e5d, 32'h4083d14c} /* (1, 27, 4) {real, imag} */,
  {32'hc09bba7b, 32'h41231e52} /* (1, 27, 3) {real, imag} */,
  {32'h40096907, 32'hc0f4ab44} /* (1, 27, 2) {real, imag} */,
  {32'hc0d7eb7e, 32'h4209fd83} /* (1, 27, 1) {real, imag} */,
  {32'h4185105b, 32'h41935b84} /* (1, 27, 0) {real, imag} */,
  {32'hc087e8dd, 32'hbf7b487c} /* (1, 26, 31) {real, imag} */,
  {32'hc03e7dfe, 32'h4113bc74} /* (1, 26, 30) {real, imag} */,
  {32'hc0c8e7f2, 32'h40a5019b} /* (1, 26, 29) {real, imag} */,
  {32'h4040c5e2, 32'h407a7709} /* (1, 26, 28) {real, imag} */,
  {32'h40416002, 32'hc068641a} /* (1, 26, 27) {real, imag} */,
  {32'hc0c3b93f, 32'hc02948fd} /* (1, 26, 26) {real, imag} */,
  {32'h3f120f4c, 32'hc0791f53} /* (1, 26, 25) {real, imag} */,
  {32'h40164ffd, 32'hbff44446} /* (1, 26, 24) {real, imag} */,
  {32'h3fa8c8fa, 32'h40020797} /* (1, 26, 23) {real, imag} */,
  {32'h40880b00, 32'hbfc0de55} /* (1, 26, 22) {real, imag} */,
  {32'h3f34880e, 32'hbff2110c} /* (1, 26, 21) {real, imag} */,
  {32'hc026e127, 32'h3e9630f1} /* (1, 26, 20) {real, imag} */,
  {32'hbf9f8af4, 32'hbf721ec0} /* (1, 26, 19) {real, imag} */,
  {32'hbf730fde, 32'hbfd07ff5} /* (1, 26, 18) {real, imag} */,
  {32'hbe605592, 32'h3e7d11d8} /* (1, 26, 17) {real, imag} */,
  {32'h3fafc11b, 32'h4029d477} /* (1, 26, 16) {real, imag} */,
  {32'hbecc838c, 32'h3f7999ed} /* (1, 26, 15) {real, imag} */,
  {32'h3f75d0cc, 32'hbfd7f082} /* (1, 26, 14) {real, imag} */,
  {32'hc07e97b6, 32'h3f8c37c4} /* (1, 26, 13) {real, imag} */,
  {32'hbe9479e9, 32'h3f85b5e9} /* (1, 26, 12) {real, imag} */,
  {32'hbf542c75, 32'h3f1cda0f} /* (1, 26, 11) {real, imag} */,
  {32'hbf2ec3b3, 32'hbfba202c} /* (1, 26, 10) {real, imag} */,
  {32'hbfefbe55, 32'h3f8004d0} /* (1, 26, 9) {real, imag} */,
  {32'h3fa3ec49, 32'hbff8f65f} /* (1, 26, 8) {real, imag} */,
  {32'h4053a2da, 32'hc053606d} /* (1, 26, 7) {real, imag} */,
  {32'h3cb29b46, 32'hc05d5fd4} /* (1, 26, 6) {real, imag} */,
  {32'hbf5dfc92, 32'hc02dbc61} /* (1, 26, 5) {real, imag} */,
  {32'h3f611383, 32'h4041d314} /* (1, 26, 4) {real, imag} */,
  {32'h40a5628d, 32'hc0291bc8} /* (1, 26, 3) {real, imag} */,
  {32'h3f33a0fe, 32'hc0c54a3c} /* (1, 26, 2) {real, imag} */,
  {32'hc02e5067, 32'hc1095004} /* (1, 26, 1) {real, imag} */,
  {32'h40079cb4, 32'h401d0230} /* (1, 26, 0) {real, imag} */,
  {32'hc0865ac8, 32'h40b5f1bd} /* (1, 25, 31) {real, imag} */,
  {32'h409433c2, 32'h3fecd3dd} /* (1, 25, 30) {real, imag} */,
  {32'h3fa8c72e, 32'h4084a4db} /* (1, 25, 29) {real, imag} */,
  {32'hc0a3fc5c, 32'h40bfb318} /* (1, 25, 28) {real, imag} */,
  {32'h3ff03f72, 32'hc08d2d3a} /* (1, 25, 27) {real, imag} */,
  {32'h3fba4c78, 32'hc053653b} /* (1, 25, 26) {real, imag} */,
  {32'hbf02dbd2, 32'hbf8daa93} /* (1, 25, 25) {real, imag} */,
  {32'h3fb15b5a, 32'hbfa52b02} /* (1, 25, 24) {real, imag} */,
  {32'h3f811bec, 32'hbfc4bcc0} /* (1, 25, 23) {real, imag} */,
  {32'h3e8d7b52, 32'hc08b38b0} /* (1, 25, 22) {real, imag} */,
  {32'hbf8d8f81, 32'hc03f7d9e} /* (1, 25, 21) {real, imag} */,
  {32'h3fcb3157, 32'h40320b20} /* (1, 25, 20) {real, imag} */,
  {32'hbf67930d, 32'hbe843c66} /* (1, 25, 19) {real, imag} */,
  {32'h3f9100bf, 32'h40059e95} /* (1, 25, 18) {real, imag} */,
  {32'h3fe334b9, 32'h3fab317c} /* (1, 25, 17) {real, imag} */,
  {32'hbfa603f2, 32'h3ff2c167} /* (1, 25, 16) {real, imag} */,
  {32'hbfbf52db, 32'hbf55f455} /* (1, 25, 15) {real, imag} */,
  {32'h3ecf1fec, 32'hbfad74e2} /* (1, 25, 14) {real, imag} */,
  {32'hbfe64dcf, 32'hbf6f94d1} /* (1, 25, 13) {real, imag} */,
  {32'h3e49120b, 32'hbf655fed} /* (1, 25, 12) {real, imag} */,
  {32'hc012f2d6, 32'hbfe528ed} /* (1, 25, 11) {real, imag} */,
  {32'hc0355e50, 32'hbdd94058} /* (1, 25, 10) {real, imag} */,
  {32'h3fa75486, 32'h40a63d7e} /* (1, 25, 9) {real, imag} */,
  {32'h4025c705, 32'h3ff4c3bd} /* (1, 25, 8) {real, imag} */,
  {32'h4012c406, 32'hc065e631} /* (1, 25, 7) {real, imag} */,
  {32'h403c520d, 32'hbfd370ab} /* (1, 25, 6) {real, imag} */,
  {32'h3eb273fb, 32'hbf52edd4} /* (1, 25, 5) {real, imag} */,
  {32'hc0424b77, 32'h40747af2} /* (1, 25, 4) {real, imag} */,
  {32'hc0137a9c, 32'h405140fe} /* (1, 25, 3) {real, imag} */,
  {32'hc0080fce, 32'hc05bfd5a} /* (1, 25, 2) {real, imag} */,
  {32'hc0ab4394, 32'hc1203d89} /* (1, 25, 1) {real, imag} */,
  {32'h3e033c9c, 32'h3f3c350a} /* (1, 25, 0) {real, imag} */,
  {32'h409012a4, 32'h4124ce92} /* (1, 24, 31) {real, imag} */,
  {32'hbedd2a7a, 32'hc13f2f4f} /* (1, 24, 30) {real, imag} */,
  {32'h3e94e96b, 32'hbf62f008} /* (1, 24, 29) {real, imag} */,
  {32'h407f7b55, 32'h401de680} /* (1, 24, 28) {real, imag} */,
  {32'hbd98e0c1, 32'hc037683f} /* (1, 24, 27) {real, imag} */,
  {32'hc04c072f, 32'h3f0e3375} /* (1, 24, 26) {real, imag} */,
  {32'hc017e22d, 32'h40831359} /* (1, 24, 25) {real, imag} */,
  {32'hc01a5cfc, 32'hc0301769} /* (1, 24, 24) {real, imag} */,
  {32'hc0268734, 32'h3e2ea78f} /* (1, 24, 23) {real, imag} */,
  {32'h401383f9, 32'hbeeeb6f8} /* (1, 24, 22) {real, imag} */,
  {32'hbffb15b0, 32'h3fb6159a} /* (1, 24, 21) {real, imag} */,
  {32'hbfda68a7, 32'hbf9741be} /* (1, 24, 20) {real, imag} */,
  {32'h3ff700bc, 32'h3fcecc69} /* (1, 24, 19) {real, imag} */,
  {32'hbf803946, 32'hbef7b605} /* (1, 24, 18) {real, imag} */,
  {32'h3f81926d, 32'hbec3a324} /* (1, 24, 17) {real, imag} */,
  {32'hc011db6a, 32'h3f50b664} /* (1, 24, 16) {real, imag} */,
  {32'h4001ac78, 32'hbf59cd53} /* (1, 24, 15) {real, imag} */,
  {32'h3e608ecf, 32'hbfbd7cce} /* (1, 24, 14) {real, imag} */,
  {32'h3dce2417, 32'hbf2bb6f9} /* (1, 24, 13) {real, imag} */,
  {32'hbeaf9f0d, 32'h4008dc47} /* (1, 24, 12) {real, imag} */,
  {32'hbf24fe94, 32'h3f305a18} /* (1, 24, 11) {real, imag} */,
  {32'hbfc1453c, 32'h4043ea12} /* (1, 24, 10) {real, imag} */,
  {32'h402324b4, 32'h3faacd16} /* (1, 24, 9) {real, imag} */,
  {32'h3f2ec070, 32'hc08017f8} /* (1, 24, 8) {real, imag} */,
  {32'hc007ec91, 32'h3d08c4b5} /* (1, 24, 7) {real, imag} */,
  {32'hbc980722, 32'hbfecb148} /* (1, 24, 6) {real, imag} */,
  {32'h3eeebc28, 32'hc11b8949} /* (1, 24, 5) {real, imag} */,
  {32'hc06afd8d, 32'hbebee1e7} /* (1, 24, 4) {real, imag} */,
  {32'hbfd1c0e0, 32'h3efcf5f0} /* (1, 24, 3) {real, imag} */,
  {32'hbf558af0, 32'hc0c2d984} /* (1, 24, 2) {real, imag} */,
  {32'h40f77750, 32'h417d5cf5} /* (1, 24, 1) {real, imag} */,
  {32'h3fffbc67, 32'h4060332b} /* (1, 24, 0) {real, imag} */,
  {32'hc0a50389, 32'hbfe12bc7} /* (1, 23, 31) {real, imag} */,
  {32'h4084a20a, 32'h407a483d} /* (1, 23, 30) {real, imag} */,
  {32'hc0da4716, 32'hc0959960} /* (1, 23, 29) {real, imag} */,
  {32'h404224fc, 32'h401a7b20} /* (1, 23, 28) {real, imag} */,
  {32'h40937619, 32'h3fc52b0f} /* (1, 23, 27) {real, imag} */,
  {32'hbf51f932, 32'hbf8f0f40} /* (1, 23, 26) {real, imag} */,
  {32'hbf850ade, 32'h4016490c} /* (1, 23, 25) {real, imag} */,
  {32'h403bf4e9, 32'h405e7c3e} /* (1, 23, 24) {real, imag} */,
  {32'hc095a14c, 32'h40008bb4} /* (1, 23, 23) {real, imag} */,
  {32'h401ca27c, 32'h3da0535b} /* (1, 23, 22) {real, imag} */,
  {32'h3f626ab5, 32'h3f3919e5} /* (1, 23, 21) {real, imag} */,
  {32'h40080c20, 32'hbce14c5d} /* (1, 23, 20) {real, imag} */,
  {32'h3f9beece, 32'h3dafef2d} /* (1, 23, 19) {real, imag} */,
  {32'hbfb15442, 32'hbf45b389} /* (1, 23, 18) {real, imag} */,
  {32'hc0203cf3, 32'h3fc6898d} /* (1, 23, 17) {real, imag} */,
  {32'h3fa36f1b, 32'hbc12efba} /* (1, 23, 16) {real, imag} */,
  {32'hbfcbe414, 32'h401323e9} /* (1, 23, 15) {real, imag} */,
  {32'h3feade6b, 32'hbfc3e7c2} /* (1, 23, 14) {real, imag} */,
  {32'hc03468c5, 32'hbe31d07e} /* (1, 23, 13) {real, imag} */,
  {32'hc011f9e6, 32'h3f88c66e} /* (1, 23, 12) {real, imag} */,
  {32'h4015d319, 32'h3f5c0df1} /* (1, 23, 11) {real, imag} */,
  {32'h3f6b771b, 32'hbf9fef8c} /* (1, 23, 10) {real, imag} */,
  {32'h3ed15b5c, 32'h404549fd} /* (1, 23, 9) {real, imag} */,
  {32'hbf5538db, 32'h40837560} /* (1, 23, 8) {real, imag} */,
  {32'hbde78b33, 32'h3f9f11fe} /* (1, 23, 7) {real, imag} */,
  {32'h404f7ec0, 32'hc066db77} /* (1, 23, 6) {real, imag} */,
  {32'h3b9f5322, 32'h3e4e7deb} /* (1, 23, 5) {real, imag} */,
  {32'h4006569f, 32'hc032d870} /* (1, 23, 4) {real, imag} */,
  {32'hc0af2c39, 32'h3f042b04} /* (1, 23, 3) {real, imag} */,
  {32'h410c94f4, 32'hbfe34491} /* (1, 23, 2) {real, imag} */,
  {32'hc036eeb4, 32'h4042bffc} /* (1, 23, 1) {real, imag} */,
  {32'hc035798d, 32'h3f0ba218} /* (1, 23, 0) {real, imag} */,
  {32'hc02f4fed, 32'hc03a3ddf} /* (1, 22, 31) {real, imag} */,
  {32'h3ebab4e9, 32'hc0460128} /* (1, 22, 30) {real, imag} */,
  {32'h3f7d441a, 32'hbf66f25a} /* (1, 22, 29) {real, imag} */,
  {32'hbfc08022, 32'hc01761ff} /* (1, 22, 28) {real, imag} */,
  {32'h3fd5ea44, 32'hc052bc3c} /* (1, 22, 27) {real, imag} */,
  {32'hbda456c8, 32'h3f6e1c7c} /* (1, 22, 26) {real, imag} */,
  {32'h3f92b86a, 32'h3eb08718} /* (1, 22, 25) {real, imag} */,
  {32'h3f069ad1, 32'h40264a68} /* (1, 22, 24) {real, imag} */,
  {32'h3ee5c44c, 32'hc06614ab} /* (1, 22, 23) {real, imag} */,
  {32'h3f19270c, 32'h3fb484d6} /* (1, 22, 22) {real, imag} */,
  {32'hbef0eb05, 32'hbed4e984} /* (1, 22, 21) {real, imag} */,
  {32'h3f91022e, 32'hbe759bf4} /* (1, 22, 20) {real, imag} */,
  {32'h3fa52b4c, 32'h3ee5f5ee} /* (1, 22, 19) {real, imag} */,
  {32'h3fab335f, 32'h3e7d7e79} /* (1, 22, 18) {real, imag} */,
  {32'h3f35b320, 32'hbe8ec475} /* (1, 22, 17) {real, imag} */,
  {32'h3f3cf0ec, 32'h3ec17661} /* (1, 22, 16) {real, imag} */,
  {32'h3e779b25, 32'hbf3ff222} /* (1, 22, 15) {real, imag} */,
  {32'h3fa8bbe4, 32'h3fddc73c} /* (1, 22, 14) {real, imag} */,
  {32'h3f04105b, 32'h3fac391a} /* (1, 22, 13) {real, imag} */,
  {32'hbeefda1f, 32'hc010059e} /* (1, 22, 12) {real, imag} */,
  {32'hbff9eabb, 32'h3f3816d6} /* (1, 22, 11) {real, imag} */,
  {32'hbfbdf5fc, 32'hbf067274} /* (1, 22, 10) {real, imag} */,
  {32'h3f28ff38, 32'h3f05ef27} /* (1, 22, 9) {real, imag} */,
  {32'hc01802ec, 32'h3f8f1919} /* (1, 22, 8) {real, imag} */,
  {32'hbf90c833, 32'h4031e12a} /* (1, 22, 7) {real, imag} */,
  {32'h3e1555a5, 32'h3d39978e} /* (1, 22, 6) {real, imag} */,
  {32'hbe2de58e, 32'h3e1b7526} /* (1, 22, 5) {real, imag} */,
  {32'hbe3b261b, 32'hbf95466b} /* (1, 22, 4) {real, imag} */,
  {32'hbe452f11, 32'hbfba2053} /* (1, 22, 3) {real, imag} */,
  {32'h408bde3d, 32'h3fa8c1db} /* (1, 22, 2) {real, imag} */,
  {32'hc05d0fb1, 32'hbe3dfefe} /* (1, 22, 1) {real, imag} */,
  {32'hc04b00eb, 32'h4035e07c} /* (1, 22, 0) {real, imag} */,
  {32'h40bedc32, 32'h3fccc3ec} /* (1, 21, 31) {real, imag} */,
  {32'hc089599e, 32'hbf313a2a} /* (1, 21, 30) {real, imag} */,
  {32'h3f0aa5f2, 32'hbfbfb9d7} /* (1, 21, 29) {real, imag} */,
  {32'h4055d6d1, 32'hbecf1599} /* (1, 21, 28) {real, imag} */,
  {32'hbf836dd4, 32'hbf20dc90} /* (1, 21, 27) {real, imag} */,
  {32'hbea25769, 32'hc038d41f} /* (1, 21, 26) {real, imag} */,
  {32'h3f400336, 32'h3fe81d6b} /* (1, 21, 25) {real, imag} */,
  {32'hbebe1c1a, 32'h3e9d3c00} /* (1, 21, 24) {real, imag} */,
  {32'h4021fbdc, 32'hbf5055c7} /* (1, 21, 23) {real, imag} */,
  {32'hbffcd3fa, 32'h3ef088a4} /* (1, 21, 22) {real, imag} */,
  {32'h3f50bb0c, 32'hbd8b16ac} /* (1, 21, 21) {real, imag} */,
  {32'h4066e3c7, 32'h400935ff} /* (1, 21, 20) {real, imag} */,
  {32'hbf8eef61, 32'hbebf1a05} /* (1, 21, 19) {real, imag} */,
  {32'h3f73d978, 32'h3d10fd8f} /* (1, 21, 18) {real, imag} */,
  {32'hbdc7c23f, 32'hbe198f9f} /* (1, 21, 17) {real, imag} */,
  {32'h3f54e978, 32'hbfd7e4fb} /* (1, 21, 16) {real, imag} */,
  {32'h3f6dcaa7, 32'h3f711393} /* (1, 21, 15) {real, imag} */,
  {32'hc02e2546, 32'h3e4cec1e} /* (1, 21, 14) {real, imag} */,
  {32'h3e0d22ec, 32'h3ef86db1} /* (1, 21, 13) {real, imag} */,
  {32'hbe84a8b7, 32'hbfcecd1f} /* (1, 21, 12) {real, imag} */,
  {32'hbeaafb00, 32'h3cdc6ca8} /* (1, 21, 11) {real, imag} */,
  {32'hbf2a2131, 32'hbfc9852b} /* (1, 21, 10) {real, imag} */,
  {32'hbf86ec8d, 32'hbfa9ad8f} /* (1, 21, 9) {real, imag} */,
  {32'h3f860255, 32'hc0671f87} /* (1, 21, 8) {real, imag} */,
  {32'h3f63b330, 32'hbd1f410a} /* (1, 21, 7) {real, imag} */,
  {32'hbf04b0fa, 32'hc0a18fd0} /* (1, 21, 6) {real, imag} */,
  {32'hc04cdea8, 32'hc0488b06} /* (1, 21, 5) {real, imag} */,
  {32'hbdee9fc7, 32'h3e368694} /* (1, 21, 4) {real, imag} */,
  {32'hbfdc56ce, 32'h3f41a365} /* (1, 21, 3) {real, imag} */,
  {32'hc034fd9d, 32'hbfefbf6d} /* (1, 21, 2) {real, imag} */,
  {32'h40a493c2, 32'h40483920} /* (1, 21, 1) {real, imag} */,
  {32'h406a26be, 32'h40535263} /* (1, 21, 0) {real, imag} */,
  {32'h3fd6b639, 32'hbf37ee69} /* (1, 20, 31) {real, imag} */,
  {32'hbfeba609, 32'hbeb78c4f} /* (1, 20, 30) {real, imag} */,
  {32'h40190d68, 32'h3e8ad0d2} /* (1, 20, 29) {real, imag} */,
  {32'hbefdcfd1, 32'hc0101e32} /* (1, 20, 28) {real, imag} */,
  {32'h4004b40c, 32'h3dae78e1} /* (1, 20, 27) {real, imag} */,
  {32'h3ed34790, 32'hbf7da26e} /* (1, 20, 26) {real, imag} */,
  {32'hbf351fa4, 32'hbf81da52} /* (1, 20, 25) {real, imag} */,
  {32'hbf9342e4, 32'hbfedecb5} /* (1, 20, 24) {real, imag} */,
  {32'hbd69cbdf, 32'h3fb57a88} /* (1, 20, 23) {real, imag} */,
  {32'hbfb97606, 32'h402f62e0} /* (1, 20, 22) {real, imag} */,
  {32'h3d6a8969, 32'h3fb5874e} /* (1, 20, 21) {real, imag} */,
  {32'hbf2dd5ea, 32'hbfd902e8} /* (1, 20, 20) {real, imag} */,
  {32'h3f1bb97e, 32'h3f33e980} /* (1, 20, 19) {real, imag} */,
  {32'hbf797fe9, 32'h3f580c88} /* (1, 20, 18) {real, imag} */,
  {32'h3e9fef79, 32'hbeab0d4c} /* (1, 20, 17) {real, imag} */,
  {32'hbe1362a6, 32'hbff35833} /* (1, 20, 16) {real, imag} */,
  {32'h3f6619c7, 32'hbfc8841b} /* (1, 20, 15) {real, imag} */,
  {32'hc022a534, 32'hbf616e5c} /* (1, 20, 14) {real, imag} */,
  {32'hbf8f6302, 32'h3f84dca6} /* (1, 20, 13) {real, imag} */,
  {32'h3fedd6db, 32'hc0229ff0} /* (1, 20, 12) {real, imag} */,
  {32'h4023c2d9, 32'hc02266fe} /* (1, 20, 11) {real, imag} */,
  {32'h3ff2d38f, 32'h3f9156c1} /* (1, 20, 10) {real, imag} */,
  {32'h3e3b45da, 32'h3fa5b396} /* (1, 20, 9) {real, imag} */,
  {32'h3fa219bb, 32'h3fa9efa6} /* (1, 20, 8) {real, imag} */,
  {32'h3e0b26df, 32'h3dbdd786} /* (1, 20, 7) {real, imag} */,
  {32'h3d704fc2, 32'h4070b2fa} /* (1, 20, 6) {real, imag} */,
  {32'h3ec8c9c5, 32'hc040cb53} /* (1, 20, 5) {real, imag} */,
  {32'hbf6263f8, 32'hbfc1f4bd} /* (1, 20, 4) {real, imag} */,
  {32'hbf8b32d2, 32'h3eceaf9c} /* (1, 20, 3) {real, imag} */,
  {32'h3db1c527, 32'hbe849477} /* (1, 20, 2) {real, imag} */,
  {32'h407382be, 32'hbfb82010} /* (1, 20, 1) {real, imag} */,
  {32'hc09d0661, 32'h405715cd} /* (1, 20, 0) {real, imag} */,
  {32'h402f5fe5, 32'hc030c423} /* (1, 19, 31) {real, imag} */,
  {32'hbda9de6a, 32'hbf794a6e} /* (1, 19, 30) {real, imag} */,
  {32'h3fa7fcde, 32'h3fcc9b00} /* (1, 19, 29) {real, imag} */,
  {32'hc02ef729, 32'h3eb4365e} /* (1, 19, 28) {real, imag} */,
  {32'hbfe14f29, 32'hc0322daa} /* (1, 19, 27) {real, imag} */,
  {32'h3f1e9206, 32'h3f3bfbd2} /* (1, 19, 26) {real, imag} */,
  {32'h3e3c90cc, 32'h3f06602a} /* (1, 19, 25) {real, imag} */,
  {32'hbef6b690, 32'h3f5f7b52} /* (1, 19, 24) {real, imag} */,
  {32'h3fe6fe05, 32'h401548fe} /* (1, 19, 23) {real, imag} */,
  {32'hbfc7a384, 32'h3fe3f73f} /* (1, 19, 22) {real, imag} */,
  {32'h3f101259, 32'hbffb9515} /* (1, 19, 21) {real, imag} */,
  {32'h3fa0af57, 32'hbf88de2e} /* (1, 19, 20) {real, imag} */,
  {32'hc032bfcf, 32'hbf7cccbf} /* (1, 19, 19) {real, imag} */,
  {32'hbf9dab7c, 32'hbd63623e} /* (1, 19, 18) {real, imag} */,
  {32'h3faf6e2e, 32'h3f4c4b95} /* (1, 19, 17) {real, imag} */,
  {32'hbed0a384, 32'h3f4b93f5} /* (1, 19, 16) {real, imag} */,
  {32'hbeab23b5, 32'h3fbb2c7f} /* (1, 19, 15) {real, imag} */,
  {32'hbf7dc642, 32'h3fdfa624} /* (1, 19, 14) {real, imag} */,
  {32'hbf294d70, 32'h3d134101} /* (1, 19, 13) {real, imag} */,
  {32'hbf9b5291, 32'h3e9c4a0a} /* (1, 19, 12) {real, imag} */,
  {32'hbe61a32b, 32'hbe8311f3} /* (1, 19, 11) {real, imag} */,
  {32'h3fd93500, 32'h40158e9c} /* (1, 19, 10) {real, imag} */,
  {32'hbf86d0c5, 32'h3f93ddb4} /* (1, 19, 9) {real, imag} */,
  {32'h3f3ba730, 32'hbfe67f4d} /* (1, 19, 8) {real, imag} */,
  {32'h3ffb223b, 32'hc082d8db} /* (1, 19, 7) {real, imag} */,
  {32'h40665c13, 32'h3f9c669f} /* (1, 19, 6) {real, imag} */,
  {32'h3ecc777f, 32'h3f5e0468} /* (1, 19, 5) {real, imag} */,
  {32'hbe957ee5, 32'h3f0cbb5e} /* (1, 19, 4) {real, imag} */,
  {32'hbf46de87, 32'hbf609c20} /* (1, 19, 3) {real, imag} */,
  {32'hbf6bea67, 32'hbf93e232} /* (1, 19, 2) {real, imag} */,
  {32'hc00cf4b2, 32'h40360934} /* (1, 19, 1) {real, imag} */,
  {32'hbff01b4e, 32'h3ea75fae} /* (1, 19, 0) {real, imag} */,
  {32'h4072e479, 32'hbfb1aecb} /* (1, 18, 31) {real, imag} */,
  {32'hbf0b8032, 32'hbf81b975} /* (1, 18, 30) {real, imag} */,
  {32'h3fcb772f, 32'h3d4b9d6f} /* (1, 18, 29) {real, imag} */,
  {32'hc00270c8, 32'hbf2973c7} /* (1, 18, 28) {real, imag} */,
  {32'hbfe0fabd, 32'h3f307440} /* (1, 18, 27) {real, imag} */,
  {32'hbf025edb, 32'hbfbf652f} /* (1, 18, 26) {real, imag} */,
  {32'hbfa2f7e4, 32'hbfe8b479} /* (1, 18, 25) {real, imag} */,
  {32'hbe8f17ba, 32'h3f4cf01b} /* (1, 18, 24) {real, imag} */,
  {32'h40211688, 32'hbd5cf583} /* (1, 18, 23) {real, imag} */,
  {32'hbfd71641, 32'h3c69f29b} /* (1, 18, 22) {real, imag} */,
  {32'hbe9401dd, 32'h40171320} /* (1, 18, 21) {real, imag} */,
  {32'hbfd51c94, 32'hbe95d55b} /* (1, 18, 20) {real, imag} */,
  {32'h3faf9b77, 32'hbf14bd06} /* (1, 18, 19) {real, imag} */,
  {32'hbfa46a65, 32'h40046b4a} /* (1, 18, 18) {real, imag} */,
  {32'hbeb253d9, 32'hbf8c1b00} /* (1, 18, 17) {real, imag} */,
  {32'h3f68e0b7, 32'h3fc29364} /* (1, 18, 16) {real, imag} */,
  {32'hc0083aae, 32'h3e2d26a8} /* (1, 18, 15) {real, imag} */,
  {32'h3e0fab20, 32'h3dbc912d} /* (1, 18, 14) {real, imag} */,
  {32'h3fe8829c, 32'hbed19077} /* (1, 18, 13) {real, imag} */,
  {32'h3b47e049, 32'h3fd21971} /* (1, 18, 12) {real, imag} */,
  {32'h3e8298a4, 32'hc00b21af} /* (1, 18, 11) {real, imag} */,
  {32'h3da57182, 32'h3eb2b789} /* (1, 18, 10) {real, imag} */,
  {32'hc02a21f9, 32'h3f8d07e0} /* (1, 18, 9) {real, imag} */,
  {32'h3ff71bce, 32'hc04948d8} /* (1, 18, 8) {real, imag} */,
  {32'h3f86b93e, 32'hbe6473d6} /* (1, 18, 7) {real, imag} */,
  {32'hbfb78726, 32'h3dbb57e1} /* (1, 18, 6) {real, imag} */,
  {32'hbf6727ff, 32'hbe5e2dc6} /* (1, 18, 5) {real, imag} */,
  {32'hbe4d7cf6, 32'h3fe78d14} /* (1, 18, 4) {real, imag} */,
  {32'hbef711bf, 32'h40033f55} /* (1, 18, 3) {real, imag} */,
  {32'hbf669dd1, 32'hbf955736} /* (1, 18, 2) {real, imag} */,
  {32'h402cbae6, 32'h40014c0f} /* (1, 18, 1) {real, imag} */,
  {32'h4015d953, 32'h3f9cc1a7} /* (1, 18, 0) {real, imag} */,
  {32'hbec3162a, 32'hbf08169a} /* (1, 17, 31) {real, imag} */,
  {32'hbe8d62db, 32'hbebbc0cb} /* (1, 17, 30) {real, imag} */,
  {32'hbf3bcaa4, 32'hbeb76db7} /* (1, 17, 29) {real, imag} */,
  {32'h3f3e935e, 32'h3f0466b2} /* (1, 17, 28) {real, imag} */,
  {32'hbfdd1932, 32'h3e9c9b8e} /* (1, 17, 27) {real, imag} */,
  {32'h3dd490f4, 32'hbf672149} /* (1, 17, 26) {real, imag} */,
  {32'h3ee012ab, 32'h3f7c804b} /* (1, 17, 25) {real, imag} */,
  {32'hbfd179ef, 32'h40203834} /* (1, 17, 24) {real, imag} */,
  {32'hbf19ccfc, 32'hbfb9f420} /* (1, 17, 23) {real, imag} */,
  {32'h3f213c95, 32'h3e94319a} /* (1, 17, 22) {real, imag} */,
  {32'h3f8ce65b, 32'h3fbc80e1} /* (1, 17, 21) {real, imag} */,
  {32'hbf9b9b8d, 32'hbeba8858} /* (1, 17, 20) {real, imag} */,
  {32'h3e05868a, 32'hbf986e1d} /* (1, 17, 19) {real, imag} */,
  {32'hbfeae86e, 32'hbf8c8087} /* (1, 17, 18) {real, imag} */,
  {32'hbe4b9c02, 32'hbe97d001} /* (1, 17, 17) {real, imag} */,
  {32'hbeb0d866, 32'h3f3c11a3} /* (1, 17, 16) {real, imag} */,
  {32'hbd02e3f1, 32'hbe217ad9} /* (1, 17, 15) {real, imag} */,
  {32'hbf2a57ec, 32'h3f73b83f} /* (1, 17, 14) {real, imag} */,
  {32'h3f68760e, 32'h3fbccfa3} /* (1, 17, 13) {real, imag} */,
  {32'h3de5b477, 32'hbf81fe94} /* (1, 17, 12) {real, imag} */,
  {32'h3f068662, 32'h3f8d4ded} /* (1, 17, 11) {real, imag} */,
  {32'h3fef9670, 32'hbf907e41} /* (1, 17, 10) {real, imag} */,
  {32'hbf31f466, 32'h401a7d58} /* (1, 17, 9) {real, imag} */,
  {32'h401b9d7d, 32'hbdd138f0} /* (1, 17, 8) {real, imag} */,
  {32'hbf1f985c, 32'h3f61908e} /* (1, 17, 7) {real, imag} */,
  {32'h40422c14, 32'hbf80769a} /* (1, 17, 6) {real, imag} */,
  {32'h3f75a701, 32'h3ec1e93a} /* (1, 17, 5) {real, imag} */,
  {32'hbfd64d13, 32'hbf2d804b} /* (1, 17, 4) {real, imag} */,
  {32'h3f4e7403, 32'h3cf6c35b} /* (1, 17, 3) {real, imag} */,
  {32'h3f1c99b3, 32'h3e98287c} /* (1, 17, 2) {real, imag} */,
  {32'hbffdbb20, 32'h3fbd54aa} /* (1, 17, 1) {real, imag} */,
  {32'hc01b169f, 32'h3ec713ee} /* (1, 17, 0) {real, imag} */,
  {32'h3f818d20, 32'h3ef86f0a} /* (1, 16, 31) {real, imag} */,
  {32'h3f475e26, 32'h40258797} /* (1, 16, 30) {real, imag} */,
  {32'h3fd80838, 32'h3f2d16d4} /* (1, 16, 29) {real, imag} */,
  {32'h3eaa0ed8, 32'h3e027f0b} /* (1, 16, 28) {real, imag} */,
  {32'h3e21a2fe, 32'hbe96422e} /* (1, 16, 27) {real, imag} */,
  {32'h3fd937b4, 32'h3f7fef36} /* (1, 16, 26) {real, imag} */,
  {32'hbf2b9441, 32'hbfa1184c} /* (1, 16, 25) {real, imag} */,
  {32'hbe519ca3, 32'h3ff58a40} /* (1, 16, 24) {real, imag} */,
  {32'hbfb42fb1, 32'h3daac685} /* (1, 16, 23) {real, imag} */,
  {32'h3b61ff91, 32'hbfaddc8c} /* (1, 16, 22) {real, imag} */,
  {32'hbfa36618, 32'h3f730f3b} /* (1, 16, 21) {real, imag} */,
  {32'h3fafd41b, 32'h3d11291e} /* (1, 16, 20) {real, imag} */,
  {32'hbfbd17c6, 32'hbf4ef2ed} /* (1, 16, 19) {real, imag} */,
  {32'hbf6de832, 32'h3fee736c} /* (1, 16, 18) {real, imag} */,
  {32'hbd87c77d, 32'hbf8c80bb} /* (1, 16, 17) {real, imag} */,
  {32'h3f1392e1, 32'hbed7fdcd} /* (1, 16, 16) {real, imag} */,
  {32'hc007b5ae, 32'hbff2fa12} /* (1, 16, 15) {real, imag} */,
  {32'h3f8bcd92, 32'h3e9ef901} /* (1, 16, 14) {real, imag} */,
  {32'h3f95b8b3, 32'hbf68c66b} /* (1, 16, 13) {real, imag} */,
  {32'hbf1695d1, 32'hbfa75c2e} /* (1, 16, 12) {real, imag} */,
  {32'h3fc3a467, 32'hbf74089e} /* (1, 16, 11) {real, imag} */,
  {32'hbc9c7f25, 32'h3efbf6f1} /* (1, 16, 10) {real, imag} */,
  {32'h3fd406f6, 32'h3dda1ae2} /* (1, 16, 9) {real, imag} */,
  {32'h3fad19c6, 32'hbf92073d} /* (1, 16, 8) {real, imag} */,
  {32'hbe4d37c2, 32'hbf2e36cf} /* (1, 16, 7) {real, imag} */,
  {32'hbf890f30, 32'hbde5e854} /* (1, 16, 6) {real, imag} */,
  {32'hbf5b1f2b, 32'hbecfbc1b} /* (1, 16, 5) {real, imag} */,
  {32'hbf1512c6, 32'h3f3b1cea} /* (1, 16, 4) {real, imag} */,
  {32'hbf6da3c7, 32'h3eb481a6} /* (1, 16, 3) {real, imag} */,
  {32'hbf307ae3, 32'hbf11e38a} /* (1, 16, 2) {real, imag} */,
  {32'h3f9085fe, 32'h3ed3b0e6} /* (1, 16, 1) {real, imag} */,
  {32'hbe79f132, 32'hbea9a70e} /* (1, 16, 0) {real, imag} */,
  {32'h3e412b34, 32'hbf56f2fc} /* (1, 15, 31) {real, imag} */,
  {32'hbf3ab295, 32'hbdb1cbce} /* (1, 15, 30) {real, imag} */,
  {32'hbe83e5a8, 32'hbfad6794} /* (1, 15, 29) {real, imag} */,
  {32'h3f2636eb, 32'hbffe5f3e} /* (1, 15, 28) {real, imag} */,
  {32'h3fc23fef, 32'hc0014e71} /* (1, 15, 27) {real, imag} */,
  {32'h3fb615ab, 32'hbe08fa40} /* (1, 15, 26) {real, imag} */,
  {32'h3db0f2fd, 32'h400e383e} /* (1, 15, 25) {real, imag} */,
  {32'hbe3afc1b, 32'h3de7e8a3} /* (1, 15, 24) {real, imag} */,
  {32'hbdebb25d, 32'h3ed0b2ea} /* (1, 15, 23) {real, imag} */,
  {32'hbfd73cc1, 32'h4051650b} /* (1, 15, 22) {real, imag} */,
  {32'h402c9471, 32'h40350bed} /* (1, 15, 21) {real, imag} */,
  {32'h3f015bae, 32'h3ff5b649} /* (1, 15, 20) {real, imag} */,
  {32'hbf8c6498, 32'hbf9a2591} /* (1, 15, 19) {real, imag} */,
  {32'h3e5514cf, 32'hbf0a4226} /* (1, 15, 18) {real, imag} */,
  {32'hbec5f17f, 32'h3e11d6ab} /* (1, 15, 17) {real, imag} */,
  {32'h3fc1cdec, 32'hbf45b93d} /* (1, 15, 16) {real, imag} */,
  {32'hbddd7fd4, 32'h3f69ced5} /* (1, 15, 15) {real, imag} */,
  {32'hbea8d9f1, 32'h3eef1dc6} /* (1, 15, 14) {real, imag} */,
  {32'hbfcbe16a, 32'hbf94b9ff} /* (1, 15, 13) {real, imag} */,
  {32'hbda750aa, 32'hbf03a6ab} /* (1, 15, 12) {real, imag} */,
  {32'h3d6426e1, 32'hbe94d071} /* (1, 15, 11) {real, imag} */,
  {32'hbc85630a, 32'hbf95419f} /* (1, 15, 10) {real, imag} */,
  {32'hbfb2d781, 32'hbf488efb} /* (1, 15, 9) {real, imag} */,
  {32'hbfcecff6, 32'hbfa30fbb} /* (1, 15, 8) {real, imag} */,
  {32'h3f0e39d7, 32'h3f7a8231} /* (1, 15, 7) {real, imag} */,
  {32'h3f3acfa1, 32'h3f0814ce} /* (1, 15, 6) {real, imag} */,
  {32'hbf1fc5b7, 32'h3f40de12} /* (1, 15, 5) {real, imag} */,
  {32'h3f6f33c2, 32'h3eeb684a} /* (1, 15, 4) {real, imag} */,
  {32'hbf513254, 32'hc002e7cb} /* (1, 15, 3) {real, imag} */,
  {32'hbfcd813e, 32'h3f933277} /* (1, 15, 2) {real, imag} */,
  {32'h40113d7b, 32'h3e6c9b0d} /* (1, 15, 1) {real, imag} */,
  {32'h3f100cee, 32'hbf8016d5} /* (1, 15, 0) {real, imag} */,
  {32'hc08be964, 32'hbfb1996a} /* (1, 14, 31) {real, imag} */,
  {32'h3d992927, 32'hbfa37dca} /* (1, 14, 30) {real, imag} */,
  {32'h3f3dfc67, 32'hbe90c3c5} /* (1, 14, 29) {real, imag} */,
  {32'h3f2b2b68, 32'h3fbd7477} /* (1, 14, 28) {real, imag} */,
  {32'h3f835cbe, 32'h3fc09175} /* (1, 14, 27) {real, imag} */,
  {32'hbebe1b96, 32'hbf7e3aa6} /* (1, 14, 26) {real, imag} */,
  {32'hbf706505, 32'h3e05660d} /* (1, 14, 25) {real, imag} */,
  {32'h3d34b848, 32'hbf37f462} /* (1, 14, 24) {real, imag} */,
  {32'hbfd2dc28, 32'h3f926134} /* (1, 14, 23) {real, imag} */,
  {32'h3e45186e, 32'h3e99809b} /* (1, 14, 22) {real, imag} */,
  {32'h3f5ebc46, 32'hbfd11bc5} /* (1, 14, 21) {real, imag} */,
  {32'hbd98c70f, 32'hc0113816} /* (1, 14, 20) {real, imag} */,
  {32'hbf6d719b, 32'hbf87c7bf} /* (1, 14, 19) {real, imag} */,
  {32'hbf4d13da, 32'h3f9d1270} /* (1, 14, 18) {real, imag} */,
  {32'hbe831669, 32'h3ee3ac8e} /* (1, 14, 17) {real, imag} */,
  {32'h3f11de77, 32'h3e7237cc} /* (1, 14, 16) {real, imag} */,
  {32'h3fa800cd, 32'hbd83b4f4} /* (1, 14, 15) {real, imag} */,
  {32'h400ef1e0, 32'hbe57b842} /* (1, 14, 14) {real, imag} */,
  {32'hbfa59bd5, 32'h3ebac522} /* (1, 14, 13) {real, imag} */,
  {32'h3e9112c0, 32'h3f5aa8a4} /* (1, 14, 12) {real, imag} */,
  {32'h3eb88052, 32'h3fb3d030} /* (1, 14, 11) {real, imag} */,
  {32'hbfe7c218, 32'h3ee777cd} /* (1, 14, 10) {real, imag} */,
  {32'h3e15e754, 32'h3f33df29} /* (1, 14, 9) {real, imag} */,
  {32'hbf3dc827, 32'h3e88e968} /* (1, 14, 8) {real, imag} */,
  {32'hc0175c19, 32'h3f5ad9bd} /* (1, 14, 7) {real, imag} */,
  {32'h4015912a, 32'h401af90c} /* (1, 14, 6) {real, imag} */,
  {32'h40565eb0, 32'hbddf41ba} /* (1, 14, 5) {real, imag} */,
  {32'hbfce6a82, 32'h3f44bc23} /* (1, 14, 4) {real, imag} */,
  {32'hbf10b1c4, 32'h4002c461} /* (1, 14, 3) {real, imag} */,
  {32'h3f5f58fe, 32'hbecbeb24} /* (1, 14, 2) {real, imag} */,
  {32'hc076de31, 32'hbff22aa6} /* (1, 14, 1) {real, imag} */,
  {32'hc0228f13, 32'hc032571e} /* (1, 14, 0) {real, imag} */,
  {32'hc095af5f, 32'hbffb872f} /* (1, 13, 31) {real, imag} */,
  {32'h4063bfe1, 32'hc0155108} /* (1, 13, 30) {real, imag} */,
  {32'h3fbccd12, 32'h3e596391} /* (1, 13, 29) {real, imag} */,
  {32'h3feb8fbe, 32'hbf0c2d0e} /* (1, 13, 28) {real, imag} */,
  {32'hbfa0e682, 32'h40448c96} /* (1, 13, 27) {real, imag} */,
  {32'h40438ab0, 32'hbf945489} /* (1, 13, 26) {real, imag} */,
  {32'hbfe0116e, 32'hbf22d718} /* (1, 13, 25) {real, imag} */,
  {32'h3f29cf4f, 32'hbd9045fe} /* (1, 13, 24) {real, imag} */,
  {32'hbf008dea, 32'h405baede} /* (1, 13, 23) {real, imag} */,
  {32'hbfa0868a, 32'hbfcb0574} /* (1, 13, 22) {real, imag} */,
  {32'hbfc37fdc, 32'h3eadc67a} /* (1, 13, 21) {real, imag} */,
  {32'hbfe70951, 32'h40264706} /* (1, 13, 20) {real, imag} */,
  {32'hbf844687, 32'hbf654d37} /* (1, 13, 19) {real, imag} */,
  {32'h3eaede22, 32'h3e35d315} /* (1, 13, 18) {real, imag} */,
  {32'hbee31729, 32'hbf58676c} /* (1, 13, 17) {real, imag} */,
  {32'h3d573b05, 32'h3fc8c1ed} /* (1, 13, 16) {real, imag} */,
  {32'hbfc5d692, 32'hbfd0a0e1} /* (1, 13, 15) {real, imag} */,
  {32'h400b426b, 32'h400093c4} /* (1, 13, 14) {real, imag} */,
  {32'h401d2eff, 32'hbfc5e022} /* (1, 13, 13) {real, imag} */,
  {32'h3ef6d26f, 32'h3f4c55f8} /* (1, 13, 12) {real, imag} */,
  {32'h3f0b9ea0, 32'h3edcabef} /* (1, 13, 11) {real, imag} */,
  {32'hbf74ef1e, 32'h3f1b483e} /* (1, 13, 10) {real, imag} */,
  {32'hbfa36183, 32'h3e19e99d} /* (1, 13, 9) {real, imag} */,
  {32'hc04aee14, 32'h4004d974} /* (1, 13, 8) {real, imag} */,
  {32'hbead4c9a, 32'h3fee9c78} /* (1, 13, 7) {real, imag} */,
  {32'hc0390e8f, 32'hc006f539} /* (1, 13, 6) {real, imag} */,
  {32'hbe1d7700, 32'h3ea377a5} /* (1, 13, 5) {real, imag} */,
  {32'hbe97d612, 32'h3dc89d0d} /* (1, 13, 4) {real, imag} */,
  {32'h3f7b1889, 32'h3fcedea3} /* (1, 13, 3) {real, imag} */,
  {32'hbedc0e59, 32'hc00635d4} /* (1, 13, 2) {real, imag} */,
  {32'h40844eaa, 32'hc00205b5} /* (1, 13, 1) {real, imag} */,
  {32'h3fd5a783, 32'h3f70286c} /* (1, 13, 0) {real, imag} */,
  {32'h402be7f6, 32'hc05be44d} /* (1, 12, 31) {real, imag} */,
  {32'hbdcf253f, 32'h3ef2144c} /* (1, 12, 30) {real, imag} */,
  {32'h3ec55d64, 32'hc0069a28} /* (1, 12, 29) {real, imag} */,
  {32'h3ddcfd07, 32'h3f75bbb1} /* (1, 12, 28) {real, imag} */,
  {32'h3faa9b83, 32'h3fbf59ae} /* (1, 12, 27) {real, imag} */,
  {32'hbf3edac1, 32'h3ddf9a73} /* (1, 12, 26) {real, imag} */,
  {32'hc03c82a4, 32'hc04243f2} /* (1, 12, 25) {real, imag} */,
  {32'hc02e5013, 32'hbf6dba1f} /* (1, 12, 24) {real, imag} */,
  {32'h3f2dc7ec, 32'h403b4397} /* (1, 12, 23) {real, imag} */,
  {32'h40060663, 32'hbe97fe70} /* (1, 12, 22) {real, imag} */,
  {32'h3fcf6b8a, 32'h3e8e3d54} /* (1, 12, 21) {real, imag} */,
  {32'hbfcabdf1, 32'h3f221f17} /* (1, 12, 20) {real, imag} */,
  {32'hbef14f25, 32'h3f29a2af} /* (1, 12, 19) {real, imag} */,
  {32'h3f318f27, 32'hbf7f0be5} /* (1, 12, 18) {real, imag} */,
  {32'hbf804afc, 32'h3fd67960} /* (1, 12, 17) {real, imag} */,
  {32'hbf312fc1, 32'hbceb4557} /* (1, 12, 16) {real, imag} */,
  {32'hbf1f00aa, 32'h3fb4b894} /* (1, 12, 15) {real, imag} */,
  {32'h3e4ecdc5, 32'h3f0c97af} /* (1, 12, 14) {real, imag} */,
  {32'hbe385614, 32'h3fd9d3b7} /* (1, 12, 13) {real, imag} */,
  {32'hbf0e85d5, 32'h3f242ca9} /* (1, 12, 12) {real, imag} */,
  {32'hc00d171c, 32'hbfa6fcf1} /* (1, 12, 11) {real, imag} */,
  {32'hbebd38b6, 32'hc049d19e} /* (1, 12, 10) {real, imag} */,
  {32'h401b1a7b, 32'hc087fdda} /* (1, 12, 9) {real, imag} */,
  {32'hc01b1edf, 32'h3d126bdd} /* (1, 12, 8) {real, imag} */,
  {32'hbf518937, 32'h3fe428e3} /* (1, 12, 7) {real, imag} */,
  {32'h3f8c940c, 32'h3d18770e} /* (1, 12, 6) {real, imag} */,
  {32'hbd708314, 32'hc01bec0c} /* (1, 12, 5) {real, imag} */,
  {32'hbf6a199e, 32'h3ea85265} /* (1, 12, 4) {real, imag} */,
  {32'h3ea80f8a, 32'h40210cde} /* (1, 12, 3) {real, imag} */,
  {32'h3f5c0785, 32'hbf8aff8b} /* (1, 12, 2) {real, imag} */,
  {32'hc0281452, 32'hbfc841a0} /* (1, 12, 1) {real, imag} */,
  {32'h3fe85382, 32'h3f21c761} /* (1, 12, 0) {real, imag} */,
  {32'hbf2f07d3, 32'h40a56eac} /* (1, 11, 31) {real, imag} */,
  {32'h4072ac32, 32'hc06711e1} /* (1, 11, 30) {real, imag} */,
  {32'h3e581771, 32'h4021ad13} /* (1, 11, 29) {real, imag} */,
  {32'h3f67b5b8, 32'hbeb3606f} /* (1, 11, 28) {real, imag} */,
  {32'hbe3154de, 32'hc05a8b84} /* (1, 11, 27) {real, imag} */,
  {32'h3f710ad3, 32'h3ea186ca} /* (1, 11, 26) {real, imag} */,
  {32'hbf177472, 32'h407d9559} /* (1, 11, 25) {real, imag} */,
  {32'hbec17e94, 32'hbeafcf2c} /* (1, 11, 24) {real, imag} */,
  {32'hbe377a29, 32'h4003977a} /* (1, 11, 23) {real, imag} */,
  {32'hc016e5a9, 32'h3f920683} /* (1, 11, 22) {real, imag} */,
  {32'h3f835bfe, 32'hc0008c23} /* (1, 11, 21) {real, imag} */,
  {32'h3f7d20e4, 32'hbf5834bb} /* (1, 11, 20) {real, imag} */,
  {32'hbf34e7ff, 32'h3e8b16fc} /* (1, 11, 19) {real, imag} */,
  {32'hbf1397f7, 32'hbd01140d} /* (1, 11, 18) {real, imag} */,
  {32'h3efc86d5, 32'hbf74eb7a} /* (1, 11, 17) {real, imag} */,
  {32'h3f852f3a, 32'hbd0b5d9d} /* (1, 11, 16) {real, imag} */,
  {32'hbf4d43cd, 32'hbfb6c910} /* (1, 11, 15) {real, imag} */,
  {32'h3f565db2, 32'hbf0d8b98} /* (1, 11, 14) {real, imag} */,
  {32'hbfcd8d40, 32'hbeca8e77} /* (1, 11, 13) {real, imag} */,
  {32'hbde2ca78, 32'hbdc8e9d0} /* (1, 11, 12) {real, imag} */,
  {32'hbf3dd551, 32'h401c7065} /* (1, 11, 11) {real, imag} */,
  {32'hbfa4ffdc, 32'h403a709f} /* (1, 11, 10) {real, imag} */,
  {32'hbf8f6823, 32'hbf292a38} /* (1, 11, 9) {real, imag} */,
  {32'h3e81d1f1, 32'hbfd3d129} /* (1, 11, 8) {real, imag} */,
  {32'hbd9e9074, 32'hbf607380} /* (1, 11, 7) {real, imag} */,
  {32'hbf8dfe58, 32'hbff32a04} /* (1, 11, 6) {real, imag} */,
  {32'h3fb04ea7, 32'h3f4cbff6} /* (1, 11, 5) {real, imag} */,
  {32'hc0037859, 32'hbf834568} /* (1, 11, 4) {real, imag} */,
  {32'h3f8fc082, 32'h3f832640} /* (1, 11, 3) {real, imag} */,
  {32'h40419d4e, 32'h4012050c} /* (1, 11, 2) {real, imag} */,
  {32'hc09ad55e, 32'h3fecabb5} /* (1, 11, 1) {real, imag} */,
  {32'hc081f377, 32'h3e83a5ce} /* (1, 11, 0) {real, imag} */,
  {32'h40383bde, 32'hbff3419e} /* (1, 10, 31) {real, imag} */,
  {32'hc0780fa5, 32'h40748377} /* (1, 10, 30) {real, imag} */,
  {32'h3fb9257a, 32'h403af9b5} /* (1, 10, 29) {real, imag} */,
  {32'h4007395e, 32'hc029f354} /* (1, 10, 28) {real, imag} */,
  {32'h40841d70, 32'hbee6d711} /* (1, 10, 27) {real, imag} */,
  {32'h4004154f, 32'hc02d5da7} /* (1, 10, 26) {real, imag} */,
  {32'h3f711ce8, 32'hbef4d81f} /* (1, 10, 25) {real, imag} */,
  {32'h3f02d428, 32'hbf6cc8aa} /* (1, 10, 24) {real, imag} */,
  {32'hc01da3a3, 32'hc004b322} /* (1, 10, 23) {real, imag} */,
  {32'h3fe9afc7, 32'h3e80e91a} /* (1, 10, 22) {real, imag} */,
  {32'hc046052b, 32'hbfff85a5} /* (1, 10, 21) {real, imag} */,
  {32'hbeeee40b, 32'h40568f1c} /* (1, 10, 20) {real, imag} */,
  {32'h402fa7b5, 32'h3fa22842} /* (1, 10, 19) {real, imag} */,
  {32'hbf2817bf, 32'h3f0571a1} /* (1, 10, 18) {real, imag} */,
  {32'hbf90b800, 32'hbfccbb57} /* (1, 10, 17) {real, imag} */,
  {32'h3f6e457a, 32'h3f36445a} /* (1, 10, 16) {real, imag} */,
  {32'h4022017d, 32'hbf291cf3} /* (1, 10, 15) {real, imag} */,
  {32'h3ed4fd4f, 32'h3f17a100} /* (1, 10, 14) {real, imag} */,
  {32'h3e4be579, 32'h3ef33953} /* (1, 10, 13) {real, imag} */,
  {32'h3dfbe87a, 32'hbff78e78} /* (1, 10, 12) {real, imag} */,
  {32'hbff06e71, 32'hc023b567} /* (1, 10, 11) {real, imag} */,
  {32'hbfadaef9, 32'h400ca718} /* (1, 10, 10) {real, imag} */,
  {32'h3f5d4a88, 32'h3aeefa4e} /* (1, 10, 9) {real, imag} */,
  {32'h3e47a747, 32'hc00b7553} /* (1, 10, 8) {real, imag} */,
  {32'h401f594c, 32'h3d71f007} /* (1, 10, 7) {real, imag} */,
  {32'h3fe3c034, 32'hbf9cbbe1} /* (1, 10, 6) {real, imag} */,
  {32'hc06f0cb9, 32'hc05dc255} /* (1, 10, 5) {real, imag} */,
  {32'h40483d5b, 32'h3f837128} /* (1, 10, 4) {real, imag} */,
  {32'h3fe8f4e2, 32'h3c188db3} /* (1, 10, 3) {real, imag} */,
  {32'hc08b10db, 32'hbf146348} /* (1, 10, 2) {real, imag} */,
  {32'h3ff86b9c, 32'hc053ba7a} /* (1, 10, 1) {real, imag} */,
  {32'h3f87df4f, 32'hbf76ce24} /* (1, 10, 0) {real, imag} */,
  {32'h3feab4c5, 32'h40557dc7} /* (1, 9, 31) {real, imag} */,
  {32'hbf5e64ef, 32'hbe077887} /* (1, 9, 30) {real, imag} */,
  {32'hc049536b, 32'hbe28a974} /* (1, 9, 29) {real, imag} */,
  {32'hbf1e17e8, 32'hbf83740a} /* (1, 9, 28) {real, imag} */,
  {32'h3fa00ff2, 32'h40673690} /* (1, 9, 27) {real, imag} */,
  {32'hbf92ea80, 32'hc0876faa} /* (1, 9, 26) {real, imag} */,
  {32'hbefc61ea, 32'h3e572340} /* (1, 9, 25) {real, imag} */,
  {32'hbfe0cbdc, 32'hbfbbc197} /* (1, 9, 24) {real, imag} */,
  {32'hbf9eda83, 32'hc010208c} /* (1, 9, 23) {real, imag} */,
  {32'hbf834740, 32'hbf5fbddf} /* (1, 9, 22) {real, imag} */,
  {32'h3e66ccf0, 32'hbfa36655} /* (1, 9, 21) {real, imag} */,
  {32'h3fdaef10, 32'hbf3ac462} /* (1, 9, 20) {real, imag} */,
  {32'hc01e491d, 32'h3faeccc7} /* (1, 9, 19) {real, imag} */,
  {32'hbe9410e9, 32'h3fcf9d71} /* (1, 9, 18) {real, imag} */,
  {32'h402397ad, 32'hbfaf1e95} /* (1, 9, 17) {real, imag} */,
  {32'h404788e9, 32'hbe7b48b1} /* (1, 9, 16) {real, imag} */,
  {32'hbef96ccc, 32'h40403b1d} /* (1, 9, 15) {real, imag} */,
  {32'hc011ea36, 32'h3f87a171} /* (1, 9, 14) {real, imag} */,
  {32'hbc2360d4, 32'hbf875a84} /* (1, 9, 13) {real, imag} */,
  {32'h3f0eb261, 32'h3f8a9177} /* (1, 9, 12) {real, imag} */,
  {32'hc00f7c54, 32'hbf1ba66b} /* (1, 9, 11) {real, imag} */,
  {32'hbf504fe9, 32'hbf93e724} /* (1, 9, 10) {real, imag} */,
  {32'h3ed54fad, 32'h3ef0398b} /* (1, 9, 9) {real, imag} */,
  {32'h3f99e880, 32'h3dc7827d} /* (1, 9, 8) {real, imag} */,
  {32'h404177b4, 32'hbf626274} /* (1, 9, 7) {real, imag} */,
  {32'h3e7bb245, 32'h40728afd} /* (1, 9, 6) {real, imag} */,
  {32'hc0641535, 32'h4045ab8a} /* (1, 9, 5) {real, imag} */,
  {32'h403e0bdb, 32'h3f6a0a8b} /* (1, 9, 4) {real, imag} */,
  {32'h3eb8022d, 32'hbf81821c} /* (1, 9, 3) {real, imag} */,
  {32'hc022b7ec, 32'hc08af764} /* (1, 9, 2) {real, imag} */,
  {32'h40927803, 32'hc007e91f} /* (1, 9, 1) {real, imag} */,
  {32'hc0e05343, 32'h402f6bc9} /* (1, 9, 0) {real, imag} */,
  {32'hc0e4bf63, 32'h412190c1} /* (1, 8, 31) {real, imag} */,
  {32'h3fcfe120, 32'hc0ad4816} /* (1, 8, 30) {real, imag} */,
  {32'h3f8a314a, 32'h3fca0f8c} /* (1, 8, 29) {real, imag} */,
  {32'h3fc812ed, 32'hbfc6c3b7} /* (1, 8, 28) {real, imag} */,
  {32'hc00b83e8, 32'hc1267ab1} /* (1, 8, 27) {real, imag} */,
  {32'h401eef85, 32'hbf94e423} /* (1, 8, 26) {real, imag} */,
  {32'h4014936d, 32'h403044c4} /* (1, 8, 25) {real, imag} */,
  {32'hbf0d9b54, 32'h405627f4} /* (1, 8, 24) {real, imag} */,
  {32'hbf122d7e, 32'hbfbf6728} /* (1, 8, 23) {real, imag} */,
  {32'h3fca3d71, 32'hbfec697e} /* (1, 8, 22) {real, imag} */,
  {32'h3fae5eae, 32'hbef80a72} /* (1, 8, 21) {real, imag} */,
  {32'h3e20c76a, 32'hbfc6a66a} /* (1, 8, 20) {real, imag} */,
  {32'h3e86e151, 32'h3f5c5204} /* (1, 8, 19) {real, imag} */,
  {32'hbdb58dd1, 32'hc043946a} /* (1, 8, 18) {real, imag} */,
  {32'h3f5efda2, 32'h4008c90d} /* (1, 8, 17) {real, imag} */,
  {32'h3f932648, 32'hbfba007e} /* (1, 8, 16) {real, imag} */,
  {32'h3f8f3828, 32'h3fc6edc1} /* (1, 8, 15) {real, imag} */,
  {32'hbe8ad6a5, 32'h3db78bc7} /* (1, 8, 14) {real, imag} */,
  {32'h4020f0d6, 32'h3f5a1f2e} /* (1, 8, 13) {real, imag} */,
  {32'hbf2f5895, 32'hbfd5f43c} /* (1, 8, 12) {real, imag} */,
  {32'hbfdf5dd4, 32'h3fcac007} /* (1, 8, 11) {real, imag} */,
  {32'h3f7a487e, 32'hbfebe1b4} /* (1, 8, 10) {real, imag} */,
  {32'h3ff8efe3, 32'h3faaf990} /* (1, 8, 9) {real, imag} */,
  {32'h405ccb28, 32'hc04c7dae} /* (1, 8, 8) {real, imag} */,
  {32'h40416878, 32'h3fbafdc3} /* (1, 8, 7) {real, imag} */,
  {32'hc086f6f7, 32'h3fcb36d0} /* (1, 8, 6) {real, imag} */,
  {32'h40629544, 32'hbf90bb22} /* (1, 8, 5) {real, imag} */,
  {32'hc09cc120, 32'h40cde85c} /* (1, 8, 4) {real, imag} */,
  {32'hbedec9e5, 32'h3e8e00d5} /* (1, 8, 3) {real, imag} */,
  {32'h40367e84, 32'hc1037261} /* (1, 8, 2) {real, imag} */,
  {32'hc0aa3801, 32'h40a0fa9c} /* (1, 8, 1) {real, imag} */,
  {32'hc08b7462, 32'h408cebb7} /* (1, 8, 0) {real, imag} */,
  {32'h3f5195d5, 32'hc09dc796} /* (1, 7, 31) {real, imag} */,
  {32'hc0c410b0, 32'h40c58bb1} /* (1, 7, 30) {real, imag} */,
  {32'h3f8b6e18, 32'h4069308f} /* (1, 7, 29) {real, imag} */,
  {32'hc045ff83, 32'h3f530ac8} /* (1, 7, 28) {real, imag} */,
  {32'h3eb11e4c, 32'hbee2d6f3} /* (1, 7, 27) {real, imag} */,
  {32'h3fe99f3a, 32'h3ecd0f71} /* (1, 7, 26) {real, imag} */,
  {32'hbf8bb162, 32'hbf82daaf} /* (1, 7, 25) {real, imag} */,
  {32'hbf5f8b88, 32'h3f8ea523} /* (1, 7, 24) {real, imag} */,
  {32'hc037a0b8, 32'h40aef25e} /* (1, 7, 23) {real, imag} */,
  {32'h3fb78b39, 32'hbfe88e17} /* (1, 7, 22) {real, imag} */,
  {32'h3f06a278, 32'h3f798add} /* (1, 7, 21) {real, imag} */,
  {32'hbf850c4c, 32'hbf9f8f57} /* (1, 7, 20) {real, imag} */,
  {32'h3f764e5a, 32'hbeb4b5f8} /* (1, 7, 19) {real, imag} */,
  {32'hbf8bcba3, 32'hbf903ad9} /* (1, 7, 18) {real, imag} */,
  {32'h3f4d2ac3, 32'h3f154163} /* (1, 7, 17) {real, imag} */,
  {32'h3fa09cf0, 32'h3f0139c8} /* (1, 7, 16) {real, imag} */,
  {32'h3e4a8f08, 32'h3ddee26a} /* (1, 7, 15) {real, imag} */,
  {32'hbf0f9621, 32'hbfc535a3} /* (1, 7, 14) {real, imag} */,
  {32'hbe6a14c2, 32'h4049cdcb} /* (1, 7, 13) {real, imag} */,
  {32'hc00b14c1, 32'h3efae141} /* (1, 7, 12) {real, imag} */,
  {32'hbf7bca81, 32'hc02363fa} /* (1, 7, 11) {real, imag} */,
  {32'h3ff546cb, 32'hc07459a1} /* (1, 7, 10) {real, imag} */,
  {32'h40b6da70, 32'h3fa0b8ae} /* (1, 7, 9) {real, imag} */,
  {32'h3f6c39bc, 32'h3fcd7291} /* (1, 7, 8) {real, imag} */,
  {32'h401528b8, 32'hbfe6a6ea} /* (1, 7, 7) {real, imag} */,
  {32'hbfd6aba3, 32'h3fe7b85e} /* (1, 7, 6) {real, imag} */,
  {32'h4079b545, 32'hbf858ecf} /* (1, 7, 5) {real, imag} */,
  {32'h400e8ee2, 32'hbdeb0e5d} /* (1, 7, 4) {real, imag} */,
  {32'hbf9ea797, 32'h40314e01} /* (1, 7, 3) {real, imag} */,
  {32'hc0e0ad80, 32'h406fde6f} /* (1, 7, 2) {real, imag} */,
  {32'h4130aa83, 32'hc061b55e} /* (1, 7, 1) {real, imag} */,
  {32'h40fd9587, 32'hc01b2a8b} /* (1, 7, 0) {real, imag} */,
  {32'hc05d0c51, 32'h40662491} /* (1, 6, 31) {real, imag} */,
  {32'hc0c015f3, 32'hbdb64700} /* (1, 6, 30) {real, imag} */,
  {32'h40754371, 32'hbf7e4ab9} /* (1, 6, 29) {real, imag} */,
  {32'hc07015b6, 32'h3f030fa1} /* (1, 6, 28) {real, imag} */,
  {32'h404727b2, 32'hc06e5f86} /* (1, 6, 27) {real, imag} */,
  {32'h3f5503d7, 32'hc02df677} /* (1, 6, 26) {real, imag} */,
  {32'h3f96787c, 32'h3fa0b8e5} /* (1, 6, 25) {real, imag} */,
  {32'h401080e0, 32'h406530d6} /* (1, 6, 24) {real, imag} */,
  {32'hbfeec62b, 32'hc0768424} /* (1, 6, 23) {real, imag} */,
  {32'hbdc43537, 32'hbf12d3af} /* (1, 6, 22) {real, imag} */,
  {32'hbf469b5f, 32'hc03f9ce4} /* (1, 6, 21) {real, imag} */,
  {32'hbe1af801, 32'h402634e2} /* (1, 6, 20) {real, imag} */,
  {32'h4006202b, 32'hc01f55a8} /* (1, 6, 19) {real, imag} */,
  {32'h3ee36f8d, 32'h3f5e414f} /* (1, 6, 18) {real, imag} */,
  {32'hbfcb168a, 32'h3f9cc199} /* (1, 6, 17) {real, imag} */,
  {32'h3f89e255, 32'h3ee28903} /* (1, 6, 16) {real, imag} */,
  {32'hbff8022d, 32'hbf1a4bf9} /* (1, 6, 15) {real, imag} */,
  {32'hbfa0d9be, 32'h3e52ab43} /* (1, 6, 14) {real, imag} */,
  {32'h3d68b3ec, 32'h3f7315c3} /* (1, 6, 13) {real, imag} */,
  {32'hbfff588c, 32'h3d0f3424} /* (1, 6, 12) {real, imag} */,
  {32'h3edb90a8, 32'hc03eca24} /* (1, 6, 11) {real, imag} */,
  {32'h3f4ffa8e, 32'hc0473037} /* (1, 6, 10) {real, imag} */,
  {32'h407ccc96, 32'h407fee99} /* (1, 6, 9) {real, imag} */,
  {32'h3d6a9425, 32'hbf15ac45} /* (1, 6, 8) {real, imag} */,
  {32'h404c5ec8, 32'hbfb7a113} /* (1, 6, 7) {real, imag} */,
  {32'h3dce4676, 32'h406078bd} /* (1, 6, 6) {real, imag} */,
  {32'hbde99d7e, 32'h4030e0d1} /* (1, 6, 5) {real, imag} */,
  {32'h401ff486, 32'hc0083027} /* (1, 6, 4) {real, imag} */,
  {32'h4002a5e3, 32'h40a02d2b} /* (1, 6, 3) {real, imag} */,
  {32'hc0de9241, 32'h40218deb} /* (1, 6, 2) {real, imag} */,
  {32'hc058cc7e, 32'hbfec3245} /* (1, 6, 1) {real, imag} */,
  {32'h40e9f4dd, 32'hc0526f8b} /* (1, 6, 0) {real, imag} */,
  {32'hbfc6fcba, 32'h41ba6d4e} /* (1, 5, 31) {real, imag} */,
  {32'h407f630c, 32'hc17451df} /* (1, 5, 30) {real, imag} */,
  {32'hbff953b3, 32'hbf5f9430} /* (1, 5, 29) {real, imag} */,
  {32'h404c158b, 32'hbfabf1b0} /* (1, 5, 28) {real, imag} */,
  {32'h405feff4, 32'hc0c76489} /* (1, 5, 27) {real, imag} */,
  {32'h40524e1d, 32'hc01f3e23} /* (1, 5, 26) {real, imag} */,
  {32'h3fe81a00, 32'h4001856e} /* (1, 5, 25) {real, imag} */,
  {32'hc071ed45, 32'h3fb8235a} /* (1, 5, 24) {real, imag} */,
  {32'h3bfcc686, 32'hbf8532a3} /* (1, 5, 23) {real, imag} */,
  {32'hbf9a132b, 32'h3bed0b6e} /* (1, 5, 22) {real, imag} */,
  {32'hbff60355, 32'hbeeb03bd} /* (1, 5, 21) {real, imag} */,
  {32'h3e2f5e7b, 32'h3fd05a73} /* (1, 5, 20) {real, imag} */,
  {32'h3fab88fd, 32'h3f938f3b} /* (1, 5, 19) {real, imag} */,
  {32'hc057bda1, 32'h4014a430} /* (1, 5, 18) {real, imag} */,
  {32'hbfa7cd4e, 32'hbe797c2a} /* (1, 5, 17) {real, imag} */,
  {32'hbece53ad, 32'hbf4c4bed} /* (1, 5, 16) {real, imag} */,
  {32'hbfe9e9cd, 32'hbfb7fca5} /* (1, 5, 15) {real, imag} */,
  {32'h400a9a3f, 32'hbf11baf4} /* (1, 5, 14) {real, imag} */,
  {32'h3f87685c, 32'hbf25df9a} /* (1, 5, 13) {real, imag} */,
  {32'hbfbbf870, 32'h3edf1e7d} /* (1, 5, 12) {real, imag} */,
  {32'h3cdb3c01, 32'hbffe8f55} /* (1, 5, 11) {real, imag} */,
  {32'h405915a5, 32'h3ea3be6f} /* (1, 5, 10) {real, imag} */,
  {32'h4001d0c2, 32'h3fb513d3} /* (1, 5, 9) {real, imag} */,
  {32'hbf568f22, 32'hbf9faa39} /* (1, 5, 8) {real, imag} */,
  {32'hc086d206, 32'h407bd098} /* (1, 5, 7) {real, imag} */,
  {32'h3fbce8f7, 32'h3fa8fd41} /* (1, 5, 6) {real, imag} */,
  {32'h4015c1ba, 32'hc0d4716e} /* (1, 5, 5) {real, imag} */,
  {32'hc12c9a50, 32'h3f5efea8} /* (1, 5, 4) {real, imag} */,
  {32'h3ff1725d, 32'hbef9ddc5} /* (1, 5, 3) {real, imag} */,
  {32'h41ccb713, 32'hc06f4438} /* (1, 5, 2) {real, imag} */,
  {32'hc1b22a28, 32'h40e42970} /* (1, 5, 1) {real, imag} */,
  {32'hc13ae3c2, 32'h410a3851} /* (1, 5, 0) {real, imag} */,
  {32'h41d5ed1b, 32'h4078323f} /* (1, 4, 31) {real, imag} */,
  {32'hc1dca5de, 32'h42071833} /* (1, 4, 30) {real, imag} */,
  {32'hc03af72a, 32'h40ba6b24} /* (1, 4, 29) {real, imag} */,
  {32'h41158831, 32'hc15843e9} /* (1, 4, 28) {real, imag} */,
  {32'hbf435fcb, 32'h40c3a4d3} /* (1, 4, 27) {real, imag} */,
  {32'h4091d70c, 32'h3f82f947} /* (1, 4, 26) {real, imag} */,
  {32'hbfb7549b, 32'hc0cffe0b} /* (1, 4, 25) {real, imag} */,
  {32'hc110cfd6, 32'h40921bb5} /* (1, 4, 24) {real, imag} */,
  {32'hc0270a20, 32'hbfe80d2c} /* (1, 4, 23) {real, imag} */,
  {32'hbf8e6661, 32'hbe064ef6} /* (1, 4, 22) {real, imag} */,
  {32'h3f8b48ef, 32'hc023b76e} /* (1, 4, 21) {real, imag} */,
  {32'h3ff17d6c, 32'h3e3875cf} /* (1, 4, 20) {real, imag} */,
  {32'hbee64a2a, 32'h401c2c42} /* (1, 4, 19) {real, imag} */,
  {32'hbfaa514c, 32'h3fcf95ad} /* (1, 4, 18) {real, imag} */,
  {32'h3fa1ed52, 32'hbf3c3b56} /* (1, 4, 17) {real, imag} */,
  {32'h3f2985d7, 32'hbfae77c2} /* (1, 4, 16) {real, imag} */,
  {32'hbe8a24b0, 32'h3f2e7925} /* (1, 4, 15) {real, imag} */,
  {32'hc04d7a1c, 32'h3f433794} /* (1, 4, 14) {real, imag} */,
  {32'h3f899e70, 32'hbecb4847} /* (1, 4, 13) {real, imag} */,
  {32'h409ec28c, 32'hbfc3262d} /* (1, 4, 12) {real, imag} */,
  {32'hc083f46a, 32'h3fa28daf} /* (1, 4, 11) {real, imag} */,
  {32'hbfd289a8, 32'h3eceed64} /* (1, 4, 10) {real, imag} */,
  {32'h3f3cc9e2, 32'hbf9f90e3} /* (1, 4, 9) {real, imag} */,
  {32'hc0aaeb2a, 32'h40b1e5bd} /* (1, 4, 8) {real, imag} */,
  {32'hbe2ffc5f, 32'h3e487aaf} /* (1, 4, 7) {real, imag} */,
  {32'h403efcff, 32'hc0c3cbde} /* (1, 4, 6) {real, imag} */,
  {32'hc07946bc, 32'hbfba3d84} /* (1, 4, 5) {real, imag} */,
  {32'h41612e92, 32'h4095cb99} /* (1, 4, 4) {real, imag} */,
  {32'h41814fcb, 32'h41321ad2} /* (1, 4, 3) {real, imag} */,
  {32'hc1be648c, 32'h41d76d83} /* (1, 4, 2) {real, imag} */,
  {32'h4080ba3c, 32'hc1e55f98} /* (1, 4, 1) {real, imag} */,
  {32'h4146a760, 32'hc1422e5c} /* (1, 4, 0) {real, imag} */,
  {32'h418db6d8, 32'h423baebc} /* (1, 3, 31) {real, imag} */,
  {32'hc22dba90, 32'hc208b6ca} /* (1, 3, 30) {real, imag} */,
  {32'h40c34e79, 32'hbeda147a} /* (1, 3, 29) {real, imag} */,
  {32'h410533e4, 32'hc135567c} /* (1, 3, 28) {real, imag} */,
  {32'h409238b9, 32'h40b11d43} /* (1, 3, 27) {real, imag} */,
  {32'h400a7054, 32'h405d7f5a} /* (1, 3, 26) {real, imag} */,
  {32'h405b3196, 32'hbf994a0c} /* (1, 3, 25) {real, imag} */,
  {32'hc0a4e06e, 32'h401438d0} /* (1, 3, 24) {real, imag} */,
  {32'h3f879b70, 32'hbf8273ce} /* (1, 3, 23) {real, imag} */,
  {32'h405e795d, 32'h4043bee8} /* (1, 3, 22) {real, imag} */,
  {32'hc005c1be, 32'hbf37f442} /* (1, 3, 21) {real, imag} */,
  {32'h3ec92e59, 32'h3eebc76e} /* (1, 3, 20) {real, imag} */,
  {32'h3f0ba43b, 32'h3f1c3423} /* (1, 3, 19) {real, imag} */,
  {32'hbff14442, 32'h3f64b853} /* (1, 3, 18) {real, imag} */,
  {32'h3fdc1770, 32'hc02996f7} /* (1, 3, 17) {real, imag} */,
  {32'hbfaaa570, 32'hbda43bd3} /* (1, 3, 16) {real, imag} */,
  {32'h3f8964d2, 32'hbec77069} /* (1, 3, 15) {real, imag} */,
  {32'hbfd66753, 32'hbec6802d} /* (1, 3, 14) {real, imag} */,
  {32'hbe5fccb7, 32'hbf90e310} /* (1, 3, 13) {real, imag} */,
  {32'h3fe3ca16, 32'hbefb83dd} /* (1, 3, 12) {real, imag} */,
  {32'hbfe3bb99, 32'hc00fb292} /* (1, 3, 11) {real, imag} */,
  {32'hbf863e64, 32'hc0172f33} /* (1, 3, 10) {real, imag} */,
  {32'h40824be9, 32'h3fcf494b} /* (1, 3, 9) {real, imag} */,
  {32'h3f4a695e, 32'h3e2fd4c2} /* (1, 3, 8) {real, imag} */,
  {32'hc0147cab, 32'h3fcce75d} /* (1, 3, 7) {real, imag} */,
  {32'hc1099b50, 32'hc0e2976f} /* (1, 3, 6) {real, imag} */,
  {32'h3fdcc3eb, 32'hc06cdbed} /* (1, 3, 5) {real, imag} */,
  {32'h409e1d60, 32'h4166a721} /* (1, 3, 4) {real, imag} */,
  {32'hc05815b0, 32'h40e3d64c} /* (1, 3, 3) {real, imag} */,
  {32'hc20a3ff3, 32'h4058c6da} /* (1, 3, 2) {real, imag} */,
  {32'h41f56310, 32'hc1bafaa6} /* (1, 3, 1) {real, imag} */,
  {32'h3ffed618, 32'h41415cf9} /* (1, 3, 0) {real, imag} */,
  {32'hc2618a05, 32'h43cb743e} /* (1, 2, 31) {real, imag} */,
  {32'hc1c404b4, 32'hc33dfba2} /* (1, 2, 30) {real, imag} */,
  {32'h40e0cf33, 32'h3f9726d0} /* (1, 2, 29) {real, imag} */,
  {32'h41722c3e, 32'h415751c0} /* (1, 2, 28) {real, imag} */,
  {32'hc0acfcf4, 32'hc11da220} /* (1, 2, 27) {real, imag} */,
  {32'hc07de68f, 32'hbfd86a91} /* (1, 2, 26) {real, imag} */,
  {32'hc08b6286, 32'h40ba04e2} /* (1, 2, 25) {real, imag} */,
  {32'hbfd155e6, 32'hbf5399b3} /* (1, 2, 24) {real, imag} */,
  {32'h404b9db5, 32'h4015a8b2} /* (1, 2, 23) {real, imag} */,
  {32'h400da93a, 32'hc030d079} /* (1, 2, 22) {real, imag} */,
  {32'hc01c90d5, 32'hbf90f220} /* (1, 2, 21) {real, imag} */,
  {32'hbf1fc917, 32'h3fc8fc65} /* (1, 2, 20) {real, imag} */,
  {32'h3f172da3, 32'hc0408e89} /* (1, 2, 19) {real, imag} */,
  {32'hc05871bf, 32'hbbed09ec} /* (1, 2, 18) {real, imag} */,
  {32'h40250f7a, 32'h3f697eca} /* (1, 2, 17) {real, imag} */,
  {32'hbf0477ea, 32'hbf8195ac} /* (1, 2, 16) {real, imag} */,
  {32'hbe3828e9, 32'h3eff18f5} /* (1, 2, 15) {real, imag} */,
  {32'h3f19226c, 32'hbfac12e0} /* (1, 2, 14) {real, imag} */,
  {32'h3e79231f, 32'hbf2d7d20} /* (1, 2, 13) {real, imag} */,
  {32'h3fc1d77e, 32'hbfcc5434} /* (1, 2, 12) {real, imag} */,
  {32'h40d15181, 32'h3ed00a88} /* (1, 2, 11) {real, imag} */,
  {32'h3f379520, 32'h3fa4baac} /* (1, 2, 10) {real, imag} */,
  {32'h4068d29d, 32'hbdac41c5} /* (1, 2, 9) {real, imag} */,
  {32'hc0136634, 32'h3e963717} /* (1, 2, 8) {real, imag} */,
  {32'hbfe4fe7e, 32'h40974ea7} /* (1, 2, 7) {real, imag} */,
  {32'h3f8d126f, 32'hc08d7d53} /* (1, 2, 6) {real, imag} */,
  {32'h41c99a66, 32'hc1bcfbd2} /* (1, 2, 5) {real, imag} */,
  {32'hc153100e, 32'h4221904a} /* (1, 2, 4) {real, imag} */,
  {32'hc0590731, 32'hc02281a9} /* (1, 2, 3) {real, imag} */,
  {32'h3fab070e, 32'hc2dd3cea} /* (1, 2, 2) {real, imag} */,
  {32'hc0a50780, 32'h4375fbf4} /* (1, 2, 1) {real, imag} */,
  {32'hc285841e, 32'h434aebe0} /* (1, 2, 0) {real, imag} */,
  {32'hc2a80409, 32'hc416d8d6} /* (1, 1, 31) {real, imag} */,
  {32'hc1ce3b51, 32'h4302df7d} /* (1, 1, 30) {real, imag} */,
  {32'h41621cac, 32'hc10224ae} /* (1, 1, 29) {real, imag} */,
  {32'h418f91a2, 32'hc1a2b5a5} /* (1, 1, 28) {real, imag} */,
  {32'hc0f80d9d, 32'h41fc83b1} /* (1, 1, 27) {real, imag} */,
  {32'hc0845430, 32'hbdc1e6dc} /* (1, 1, 26) {real, imag} */,
  {32'hc017d079, 32'hc111a736} /* (1, 1, 25) {real, imag} */,
  {32'h40ea77af, 32'h40ea43b7} /* (1, 1, 24) {real, imag} */,
  {32'h402bc7f7, 32'h4007357b} /* (1, 1, 23) {real, imag} */,
  {32'hbf8ff761, 32'hc03afb85} /* (1, 1, 22) {real, imag} */,
  {32'h40d1d4ce, 32'h409a7b37} /* (1, 1, 21) {real, imag} */,
  {32'hbd427d46, 32'h3f6f415f} /* (1, 1, 20) {real, imag} */,
  {32'hbf28da14, 32'hbed6d99b} /* (1, 1, 19) {real, imag} */,
  {32'h3fcd27ac, 32'h3f22c772} /* (1, 1, 18) {real, imag} */,
  {32'h3ea6d04a, 32'hbe9b3261} /* (1, 1, 17) {real, imag} */,
  {32'hbf012c87, 32'hbeb0fd6e} /* (1, 1, 16) {real, imag} */,
  {32'h400e7989, 32'hbe8dc66d} /* (1, 1, 15) {real, imag} */,
  {32'hc03ac907, 32'hbfd2971e} /* (1, 1, 14) {real, imag} */,
  {32'h3f2e034e, 32'h3f172bc6} /* (1, 1, 13) {real, imag} */,
  {32'hc0621ccf, 32'h3f87948f} /* (1, 1, 12) {real, imag} */,
  {32'hc0d14041, 32'hbf5e3097} /* (1, 1, 11) {real, imag} */,
  {32'hc0a174a0, 32'h4004d2cd} /* (1, 1, 10) {real, imag} */,
  {32'hbe7b0c50, 32'h3fa6cd93} /* (1, 1, 9) {real, imag} */,
  {32'hc10c0492, 32'h3e293e34} /* (1, 1, 8) {real, imag} */,
  {32'hbf46adf7, 32'hc0b7705d} /* (1, 1, 7) {real, imag} */,
  {32'hc0a6d9e8, 32'h414434ac} /* (1, 1, 6) {real, imag} */,
  {32'hc16f8cb4, 32'h419a5db1} /* (1, 1, 5) {real, imag} */,
  {32'h41e97e4d, 32'hc179d236} /* (1, 1, 4) {real, imag} */,
  {32'hc059f50f, 32'h411e006d} /* (1, 1, 3) {real, imag} */,
  {32'hc33947d5, 32'h43070542} /* (1, 1, 2) {real, imag} */,
  {32'h4405adb8, 32'hc44bf626} /* (1, 1, 1) {real, imag} */,
  {32'h432eb4b6, 32'hc4392af1} /* (1, 1, 0) {real, imag} */,
  {32'hc3b5ba3a, 32'hc41220bc} /* (1, 0, 31) {real, imag} */,
  {32'h42a5062c, 32'h42aaf1e8} /* (1, 0, 30) {real, imag} */,
  {32'h40e92c10, 32'hc0b1590d} /* (1, 0, 29) {real, imag} */,
  {32'h4119f0b6, 32'h40984cf1} /* (1, 0, 28) {real, imag} */,
  {32'h40766113, 32'h41647cd2} /* (1, 0, 27) {real, imag} */,
  {32'h40282af0, 32'h3f1f976d} /* (1, 0, 26) {real, imag} */,
  {32'hc0a4ec6a, 32'h3f407311} /* (1, 0, 25) {real, imag} */,
  {32'h4086b665, 32'hc0009ca8} /* (1, 0, 24) {real, imag} */,
  {32'h3f56a504, 32'hbeaf3d27} /* (1, 0, 23) {real, imag} */,
  {32'h40542e0e, 32'h40163344} /* (1, 0, 22) {real, imag} */,
  {32'h3e720b74, 32'h40afa305} /* (1, 0, 21) {real, imag} */,
  {32'hbf8195f2, 32'hbf41d5af} /* (1, 0, 20) {real, imag} */,
  {32'hbf05cd0b, 32'hbfc0526f} /* (1, 0, 19) {real, imag} */,
  {32'h40829427, 32'h3ec200ee} /* (1, 0, 18) {real, imag} */,
  {32'hbed34cd7, 32'h3c1599da} /* (1, 0, 17) {real, imag} */,
  {32'hbf1bb697, 32'h402b344d} /* (1, 0, 16) {real, imag} */,
  {32'h3f7c92f4, 32'h4018ee15} /* (1, 0, 15) {real, imag} */,
  {32'hbf9c77e3, 32'h3fab8ca8} /* (1, 0, 14) {real, imag} */,
  {32'h3eba03a0, 32'hbf9207e4} /* (1, 0, 13) {real, imag} */,
  {32'hbfaf02d5, 32'hbeed8bee} /* (1, 0, 12) {real, imag} */,
  {32'hbf40ada2, 32'h400bc104} /* (1, 0, 11) {real, imag} */,
  {32'h3ef0d534, 32'hbf4db9d7} /* (1, 0, 10) {real, imag} */,
  {32'hbfb50995, 32'h3d9071fb} /* (1, 0, 9) {real, imag} */,
  {32'hc122d2b2, 32'h3f5f2e60} /* (1, 0, 8) {real, imag} */,
  {32'hbe5e227a, 32'h3f6ba998} /* (1, 0, 7) {real, imag} */,
  {32'hbe569a77, 32'hc0900d4c} /* (1, 0, 6) {real, imag} */,
  {32'h3eb178f7, 32'h41b2c9b5} /* (1, 0, 5) {real, imag} */,
  {32'hc10f78d7, 32'h4134bfd9} /* (1, 0, 4) {real, imag} */,
  {32'h40b9f1d8, 32'h410688cd} /* (1, 0, 3) {real, imag} */,
  {32'hc2c83a22, 32'h41b9a883} /* (1, 0, 2) {real, imag} */,
  {32'h43f8eeaf, 32'hc3f2ee9e} /* (1, 0, 1) {real, imag} */,
  {32'h42ad3089, 32'hc470e74f} /* (1, 0, 0) {real, imag} */,
  {32'hbf1c2969, 32'h41e3fcc8} /* (0, 31, 31) {real, imag} */,
  {32'hc1e94968, 32'h417f7ea1} /* (0, 31, 30) {real, imag} */,
  {32'hbfb5a27e, 32'h40c8f4d8} /* (0, 31, 29) {real, imag} */,
  {32'hc01f6fcb, 32'h4151fd65} /* (0, 31, 28) {real, imag} */,
  {32'hc051e10c, 32'hc1185483} /* (0, 31, 27) {real, imag} */,
  {32'hc08ea0b3, 32'h40dbd6e2} /* (0, 31, 26) {real, imag} */,
  {32'h3ea2be01, 32'h3f1469fb} /* (0, 31, 25) {real, imag} */,
  {32'h4036e20e, 32'h3c0fbf62} /* (0, 31, 24) {real, imag} */,
  {32'hbfa35ee5, 32'hc01853ed} /* (0, 31, 23) {real, imag} */,
  {32'hc085851e, 32'h3fe73478} /* (0, 31, 22) {real, imag} */,
  {32'hbf6c8f54, 32'hc02e4445} /* (0, 31, 21) {real, imag} */,
  {32'h40477e0c, 32'h402e3b03} /* (0, 31, 20) {real, imag} */,
  {32'h40110526, 32'h3fc5db6c} /* (0, 31, 19) {real, imag} */,
  {32'hbf74ca53, 32'hbe330d28} /* (0, 31, 18) {real, imag} */,
  {32'h3e0e6ee2, 32'hc01a93ea} /* (0, 31, 17) {real, imag} */,
  {32'hbec6804d, 32'h3fa99050} /* (0, 31, 16) {real, imag} */,
  {32'h3f92ab7d, 32'hbf561cd7} /* (0, 31, 15) {real, imag} */,
  {32'hbe7e0fd8, 32'hbffc46e8} /* (0, 31, 14) {real, imag} */,
  {32'h3fa4d3f9, 32'h40089e38} /* (0, 31, 13) {real, imag} */,
  {32'h3f9ef6ad, 32'hc04da3b2} /* (0, 31, 12) {real, imag} */,
  {32'hbed485b5, 32'hc019ed58} /* (0, 31, 11) {real, imag} */,
  {32'h4076bb1e, 32'hbc18b4b6} /* (0, 31, 10) {real, imag} */,
  {32'hbc5394ad, 32'h406aa4f6} /* (0, 31, 9) {real, imag} */,
  {32'hbfcf8fbb, 32'h40519c4b} /* (0, 31, 8) {real, imag} */,
  {32'hc09545cf, 32'hbe0d2728} /* (0, 31, 7) {real, imag} */,
  {32'h40eb03e5, 32'h40b8ee8b} /* (0, 31, 6) {real, imag} */,
  {32'h4146551a, 32'hbfb9149b} /* (0, 31, 5) {real, imag} */,
  {32'hc11d6710, 32'h408aafcf} /* (0, 31, 4) {real, imag} */,
  {32'h411d4350, 32'h40f80886} /* (0, 31, 3) {real, imag} */,
  {32'h40536963, 32'hc1de1c21} /* (0, 31, 2) {real, imag} */,
  {32'h416ccc3d, 32'h418231f0} /* (0, 31, 1) {real, imag} */,
  {32'h42236899, 32'h41aebe41} /* (0, 31, 0) {real, imag} */,
  {32'h3f780f3f, 32'hc1de58d0} /* (0, 30, 31) {real, imag} */,
  {32'h409bf46b, 32'hc117ac3b} /* (0, 30, 30) {real, imag} */,
  {32'hbffaf8f0, 32'h40d78ddf} /* (0, 30, 29) {real, imag} */,
  {32'h410b9216, 32'h416a84f5} /* (0, 30, 28) {real, imag} */,
  {32'hc11a353a, 32'h40cb3c23} /* (0, 30, 27) {real, imag} */,
  {32'h408a892a, 32'hc11189ab} /* (0, 30, 26) {real, imag} */,
  {32'h402736e8, 32'h408d88c5} /* (0, 30, 25) {real, imag} */,
  {32'hbfc8ebef, 32'h4025d3aa} /* (0, 30, 24) {real, imag} */,
  {32'h40348a5f, 32'hc09adb9c} /* (0, 30, 23) {real, imag} */,
  {32'hbcf02d69, 32'hc009faf2} /* (0, 30, 22) {real, imag} */,
  {32'hbee27faf, 32'hbe5a3195} /* (0, 30, 21) {real, imag} */,
  {32'h3f1054dd, 32'hbf67eb75} /* (0, 30, 20) {real, imag} */,
  {32'hbfd55052, 32'h3f194618} /* (0, 30, 19) {real, imag} */,
  {32'h3f988b6e, 32'h3f85249c} /* (0, 30, 18) {real, imag} */,
  {32'h3e903620, 32'h3ecdcb53} /* (0, 30, 17) {real, imag} */,
  {32'h3e9c3dd5, 32'h3dda7130} /* (0, 30, 16) {real, imag} */,
  {32'h3f14efa5, 32'h3fdf9b70} /* (0, 30, 15) {real, imag} */,
  {32'h3e5404d0, 32'h3fd43f95} /* (0, 30, 14) {real, imag} */,
  {32'hc05ac888, 32'hbfaf0628} /* (0, 30, 13) {real, imag} */,
  {32'h400c1d80, 32'h3fc36d79} /* (0, 30, 12) {real, imag} */,
  {32'h3fb36295, 32'hbf4fa318} /* (0, 30, 11) {real, imag} */,
  {32'hbfbca171, 32'h3f6c98dd} /* (0, 30, 10) {real, imag} */,
  {32'hc0649519, 32'hbefe7e3b} /* (0, 30, 9) {real, imag} */,
  {32'h400ba9a9, 32'hc0ba1e35} /* (0, 30, 8) {real, imag} */,
  {32'h403ae9ef, 32'hbe308a76} /* (0, 30, 7) {real, imag} */,
  {32'h400914be, 32'hc089e71d} /* (0, 30, 6) {real, imag} */,
  {32'h3ff1d8e1, 32'h4086a9e2} /* (0, 30, 5) {real, imag} */,
  {32'h40508a90, 32'hc0b5dca2} /* (0, 30, 4) {real, imag} */,
  {32'h417cd738, 32'hc13698b5} /* (0, 30, 3) {real, imag} */,
  {32'h415baadd, 32'h4183e558} /* (0, 30, 2) {real, imag} */,
  {32'hc0ad06dc, 32'h3e417e0b} /* (0, 30, 1) {real, imag} */,
  {32'hc181149b, 32'h40ba5814} /* (0, 30, 0) {real, imag} */,
  {32'h3f99f6f1, 32'hc141bda1} /* (0, 29, 31) {real, imag} */,
  {32'h4034ff38, 32'hc1a94125} /* (0, 29, 30) {real, imag} */,
  {32'h3f2e21c0, 32'h40d6951a} /* (0, 29, 29) {real, imag} */,
  {32'h408e1dab, 32'hc109525c} /* (0, 29, 28) {real, imag} */,
  {32'hc1094b83, 32'hc0e72d4c} /* (0, 29, 27) {real, imag} */,
  {32'hc09869e4, 32'h3f2fd050} /* (0, 29, 26) {real, imag} */,
  {32'hbf3374ff, 32'h40802a5a} /* (0, 29, 25) {real, imag} */,
  {32'hc0835cf6, 32'hc014c529} /* (0, 29, 24) {real, imag} */,
  {32'hbe89a660, 32'h400308a9} /* (0, 29, 23) {real, imag} */,
  {32'hbe016f07, 32'hbfd5821a} /* (0, 29, 22) {real, imag} */,
  {32'h3e5b8bf5, 32'h4016bc03} /* (0, 29, 21) {real, imag} */,
  {32'h40676594, 32'h408215a3} /* (0, 29, 20) {real, imag} */,
  {32'hbec62251, 32'h3f3acd5e} /* (0, 29, 19) {real, imag} */,
  {32'h3fec7d9d, 32'hc004c096} /* (0, 29, 18) {real, imag} */,
  {32'h3ecde21b, 32'h3eb38a09} /* (0, 29, 17) {real, imag} */,
  {32'h3e8e3bc6, 32'h3fa3c5c5} /* (0, 29, 16) {real, imag} */,
  {32'h3fe849ed, 32'h3e2c35f5} /* (0, 29, 15) {real, imag} */,
  {32'hbe04cbf9, 32'h401117a1} /* (0, 29, 14) {real, imag} */,
  {32'h3f8a01cd, 32'hbf9789de} /* (0, 29, 13) {real, imag} */,
  {32'hbd26a81f, 32'hbf99fb7c} /* (0, 29, 12) {real, imag} */,
  {32'hc03cf7f0, 32'h3f0a6aa1} /* (0, 29, 11) {real, imag} */,
  {32'hbec554c6, 32'hbec3e2cb} /* (0, 29, 10) {real, imag} */,
  {32'hbff85d0c, 32'h407380eb} /* (0, 29, 9) {real, imag} */,
  {32'h3fab2fad, 32'h3fd35c0c} /* (0, 29, 8) {real, imag} */,
  {32'hc0f00ed0, 32'hc09acc3f} /* (0, 29, 7) {real, imag} */,
  {32'hc0a8e599, 32'hc0201276} /* (0, 29, 6) {real, imag} */,
  {32'h3fc6fc69, 32'h40d88869} /* (0, 29, 5) {real, imag} */,
  {32'h3f2d5c7e, 32'hc04a6c80} /* (0, 29, 4) {real, imag} */,
  {32'hc0d124dd, 32'hc0d0f0ec} /* (0, 29, 3) {real, imag} */,
  {32'h4093cf3b, 32'h400bce0e} /* (0, 29, 2) {real, imag} */,
  {32'h3f2037ef, 32'h417210ea} /* (0, 29, 1) {real, imag} */,
  {32'h41c41208, 32'hc1095396} /* (0, 29, 0) {real, imag} */,
  {32'h40274864, 32'hc0c7bd15} /* (0, 28, 31) {real, imag} */,
  {32'h4180ec4d, 32'h3ed93dd8} /* (0, 28, 30) {real, imag} */,
  {32'hc0ab5f44, 32'hc08da032} /* (0, 28, 29) {real, imag} */,
  {32'h41367738, 32'h401b29f8} /* (0, 28, 28) {real, imag} */,
  {32'h4021381e, 32'h40e4bb03} /* (0, 28, 27) {real, imag} */,
  {32'hc0be6d33, 32'hc0fd5d1f} /* (0, 28, 26) {real, imag} */,
  {32'hc0be99d3, 32'h3f759371} /* (0, 28, 25) {real, imag} */,
  {32'h3f905208, 32'h3f6a05bf} /* (0, 28, 24) {real, imag} */,
  {32'h405c582f, 32'h3fde0cea} /* (0, 28, 23) {real, imag} */,
  {32'h3fd78dc5, 32'hbe7cb19c} /* (0, 28, 22) {real, imag} */,
  {32'h40521539, 32'hc03df432} /* (0, 28, 21) {real, imag} */,
  {32'hc03d8214, 32'h3fc19829} /* (0, 28, 20) {real, imag} */,
  {32'h40237b6c, 32'hbff02f88} /* (0, 28, 19) {real, imag} */,
  {32'hbd16685e, 32'hbf0ee4e9} /* (0, 28, 18) {real, imag} */,
  {32'hbfe33f35, 32'h3f5908ce} /* (0, 28, 17) {real, imag} */,
  {32'hbfb4279f, 32'hbf71540b} /* (0, 28, 16) {real, imag} */,
  {32'h3f76d61d, 32'hbf8878a2} /* (0, 28, 15) {real, imag} */,
  {32'hbf1bc6cd, 32'h3fbc6aaa} /* (0, 28, 14) {real, imag} */,
  {32'hbfd02fca, 32'h3f88b862} /* (0, 28, 13) {real, imag} */,
  {32'h40573fe8, 32'hbfd50a08} /* (0, 28, 12) {real, imag} */,
  {32'h3f330768, 32'hbffdbbd6} /* (0, 28, 11) {real, imag} */,
  {32'hbf5908b1, 32'hbee0e833} /* (0, 28, 10) {real, imag} */,
  {32'hbfee3f4e, 32'h40550856} /* (0, 28, 9) {real, imag} */,
  {32'h40b54d14, 32'h40cfd3ac} /* (0, 28, 8) {real, imag} */,
  {32'h3fca95c4, 32'hc0cc5e62} /* (0, 28, 7) {real, imag} */,
  {32'hc0d543af, 32'h40608da2} /* (0, 28, 6) {real, imag} */,
  {32'h3f59c75a, 32'h40edbcdb} /* (0, 28, 5) {real, imag} */,
  {32'hc015b0d0, 32'h3f73a440} /* (0, 28, 4) {real, imag} */,
  {32'hc0e912d9, 32'h405d6cd3} /* (0, 28, 3) {real, imag} */,
  {32'hc167492f, 32'hc108c3ce} /* (0, 28, 2) {real, imag} */,
  {32'hbf902fe7, 32'h41383efd} /* (0, 28, 1) {real, imag} */,
  {32'hc1349101, 32'h40aaa0c3} /* (0, 28, 0) {real, imag} */,
  {32'h3f4eceb3, 32'hc131b135} /* (0, 27, 31) {real, imag} */,
  {32'h40bddc69, 32'h401afe34} /* (0, 27, 30) {real, imag} */,
  {32'hc02141eb, 32'h4088ba7f} /* (0, 27, 29) {real, imag} */,
  {32'hbf84c375, 32'hc03579ac} /* (0, 27, 28) {real, imag} */,
  {32'h3ff541dc, 32'hc02beb55} /* (0, 27, 27) {real, imag} */,
  {32'hbf475c54, 32'hbf9b86bd} /* (0, 27, 26) {real, imag} */,
  {32'h40477e0e, 32'hbff7d3f3} /* (0, 27, 25) {real, imag} */,
  {32'h4063f0fa, 32'hc031a8e2} /* (0, 27, 24) {real, imag} */,
  {32'h3f912700, 32'h3fa51f0c} /* (0, 27, 23) {real, imag} */,
  {32'h3e230203, 32'hbfdab27f} /* (0, 27, 22) {real, imag} */,
  {32'hbf977e36, 32'h4090550a} /* (0, 27, 21) {real, imag} */,
  {32'h3fa0b29f, 32'h4031cf5b} /* (0, 27, 20) {real, imag} */,
  {32'h3fe2501d, 32'hbfa9306a} /* (0, 27, 19) {real, imag} */,
  {32'hbf807abb, 32'hbfe8a724} /* (0, 27, 18) {real, imag} */,
  {32'hbf992a27, 32'hbed9ce83} /* (0, 27, 17) {real, imag} */,
  {32'hbf9a452c, 32'h3e3922eb} /* (0, 27, 16) {real, imag} */,
  {32'hbf8666a0, 32'h3fbfe5da} /* (0, 27, 15) {real, imag} */,
  {32'hbf8cc1cb, 32'hbf91a24f} /* (0, 27, 14) {real, imag} */,
  {32'hbea3c10f, 32'hbfa89c17} /* (0, 27, 13) {real, imag} */,
  {32'h3f2fde6d, 32'h405598d2} /* (0, 27, 12) {real, imag} */,
  {32'h3dcb499f, 32'h403d36d7} /* (0, 27, 11) {real, imag} */,
  {32'hc05ed478, 32'h3e71db53} /* (0, 27, 10) {real, imag} */,
  {32'hbf010320, 32'hc01ae8cb} /* (0, 27, 9) {real, imag} */,
  {32'hc057cdc8, 32'h3fe4b142} /* (0, 27, 8) {real, imag} */,
  {32'hbfacfc53, 32'hc047aa9f} /* (0, 27, 7) {real, imag} */,
  {32'h3f5c8a67, 32'hc030f554} /* (0, 27, 6) {real, imag} */,
  {32'hbf5a4c16, 32'hc0957f79} /* (0, 27, 5) {real, imag} */,
  {32'hc0977a69, 32'hc08791ea} /* (0, 27, 4) {real, imag} */,
  {32'h403be311, 32'hc012f43f} /* (0, 27, 3) {real, imag} */,
  {32'hc128ceb0, 32'h40e635ad} /* (0, 27, 2) {real, imag} */,
  {32'h3f326234, 32'hc0881df2} /* (0, 27, 1) {real, imag} */,
  {32'hc0ca53d9, 32'hc0e552a7} /* (0, 27, 0) {real, imag} */,
  {32'hc041104c, 32'hbf92e5d8} /* (0, 26, 31) {real, imag} */,
  {32'h3eb0490e, 32'h4048cdb4} /* (0, 26, 30) {real, imag} */,
  {32'h40012bc6, 32'h3fc83499} /* (0, 26, 29) {real, imag} */,
  {32'h402f246c, 32'hbe8e8801} /* (0, 26, 28) {real, imag} */,
  {32'hbe8ff9e5, 32'hbd73742e} /* (0, 26, 27) {real, imag} */,
  {32'hc019fe20, 32'h4002589e} /* (0, 26, 26) {real, imag} */,
  {32'h407805ef, 32'hc0b108f9} /* (0, 26, 25) {real, imag} */,
  {32'hbfdf3f5a, 32'h40580e54} /* (0, 26, 24) {real, imag} */,
  {32'hbf1d1340, 32'hc034fcd8} /* (0, 26, 23) {real, imag} */,
  {32'hbfeabb08, 32'hbf64afd8} /* (0, 26, 22) {real, imag} */,
  {32'hbe0d73dc, 32'hbf03fd4b} /* (0, 26, 21) {real, imag} */,
  {32'h3eeb1e92, 32'hbeec9967} /* (0, 26, 20) {real, imag} */,
  {32'h4014a7f3, 32'h3fba3aca} /* (0, 26, 19) {real, imag} */,
  {32'hbe9959d4, 32'hbf267d93} /* (0, 26, 18) {real, imag} */,
  {32'h3e13548b, 32'h3e303161} /* (0, 26, 17) {real, imag} */,
  {32'hbf101065, 32'h3f70a0d1} /* (0, 26, 16) {real, imag} */,
  {32'h3cc341ee, 32'h402f0de9} /* (0, 26, 15) {real, imag} */,
  {32'h4018c91c, 32'hbf8bc7f9} /* (0, 26, 14) {real, imag} */,
  {32'hbea1ff68, 32'h3fe5f628} /* (0, 26, 13) {real, imag} */,
  {32'hbe6ed7cc, 32'h3f15b311} /* (0, 26, 12) {real, imag} */,
  {32'hbffb7cda, 32'h3f5fb73c} /* (0, 26, 11) {real, imag} */,
  {32'h4049b156, 32'h3db69013} /* (0, 26, 10) {real, imag} */,
  {32'h3ff88905, 32'hc0136e17} /* (0, 26, 9) {real, imag} */,
  {32'hc01f4568, 32'hbe893062} /* (0, 26, 8) {real, imag} */,
  {32'hbf9d3804, 32'hbecea8be} /* (0, 26, 7) {real, imag} */,
  {32'h3fe67c28, 32'hc05dd231} /* (0, 26, 6) {real, imag} */,
  {32'hbf4c4dd2, 32'h3f2604ed} /* (0, 26, 5) {real, imag} */,
  {32'h3f8fe3bf, 32'h4093c62b} /* (0, 26, 4) {real, imag} */,
  {32'h3f2fbc5b, 32'h40abc257} /* (0, 26, 3) {real, imag} */,
  {32'hc047f3b0, 32'h3f98a75f} /* (0, 26, 2) {real, imag} */,
  {32'h4019db63, 32'hc0aa3711} /* (0, 26, 1) {real, imag} */,
  {32'h406f10b5, 32'h3deea6e3} /* (0, 26, 0) {real, imag} */,
  {32'h3fcf3406, 32'hbfd669e7} /* (0, 25, 31) {real, imag} */,
  {32'hbe6586ec, 32'h3f812cc5} /* (0, 25, 30) {real, imag} */,
  {32'hbeb195c9, 32'hc0c86e82} /* (0, 25, 29) {real, imag} */,
  {32'h407014ac, 32'hbed1aa06} /* (0, 25, 28) {real, imag} */,
  {32'h405babba, 32'hbff65751} /* (0, 25, 27) {real, imag} */,
  {32'h409b5a64, 32'h4027fbd2} /* (0, 25, 26) {real, imag} */,
  {32'hc020d1e5, 32'h3fb4e2e7} /* (0, 25, 25) {real, imag} */,
  {32'hbdfd6182, 32'h4052c8af} /* (0, 25, 24) {real, imag} */,
  {32'h4035d1b3, 32'hc03c9236} /* (0, 25, 23) {real, imag} */,
  {32'hbf8ca5f1, 32'hc05be771} /* (0, 25, 22) {real, imag} */,
  {32'hbf2aeeb6, 32'hbf757ad9} /* (0, 25, 21) {real, imag} */,
  {32'hc009b319, 32'h3eb1b2ad} /* (0, 25, 20) {real, imag} */,
  {32'hbfb4fdb1, 32'hbfacf7a3} /* (0, 25, 19) {real, imag} */,
  {32'hc014188c, 32'hbdda7ec1} /* (0, 25, 18) {real, imag} */,
  {32'hbf84df0d, 32'hbfa43aa5} /* (0, 25, 17) {real, imag} */,
  {32'h3f5c5cae, 32'hbee8d40f} /* (0, 25, 16) {real, imag} */,
  {32'h3ec237b4, 32'h3e8e9d07} /* (0, 25, 15) {real, imag} */,
  {32'hbeca7955, 32'h3f89a9fa} /* (0, 25, 14) {real, imag} */,
  {32'h3cd5ce75, 32'hc03d7f0e} /* (0, 25, 13) {real, imag} */,
  {32'h3fc57e48, 32'h3ff13d57} /* (0, 25, 12) {real, imag} */,
  {32'h401deedf, 32'hbfed02e2} /* (0, 25, 11) {real, imag} */,
  {32'hbdc5b9dd, 32'hc0470058} /* (0, 25, 10) {real, imag} */,
  {32'hc0377d9c, 32'hc0ad1d62} /* (0, 25, 9) {real, imag} */,
  {32'hbff0e9f0, 32'h4042bf12} /* (0, 25, 8) {real, imag} */,
  {32'hbeb2c180, 32'hbf7ec762} /* (0, 25, 7) {real, imag} */,
  {32'hc01d4b3c, 32'hbf2fd070} /* (0, 25, 6) {real, imag} */,
  {32'hc04f4c18, 32'hc0bc1989} /* (0, 25, 5) {real, imag} */,
  {32'hc0d7acd5, 32'hbe84aa25} /* (0, 25, 4) {real, imag} */,
  {32'hc08603bb, 32'hbe4e791b} /* (0, 25, 3) {real, imag} */,
  {32'h3ed78b1a, 32'h40ae77da} /* (0, 25, 2) {real, imag} */,
  {32'hc072cf9d, 32'hbea550e2} /* (0, 25, 1) {real, imag} */,
  {32'h3e858e63, 32'h4074f16f} /* (0, 25, 0) {real, imag} */,
  {32'hc05321a3, 32'h3ef83046} /* (0, 24, 31) {real, imag} */,
  {32'hbf0a2c66, 32'h3fe2c54f} /* (0, 24, 30) {real, imag} */,
  {32'hc00b6a96, 32'hc09693bf} /* (0, 24, 29) {real, imag} */,
  {32'hc065630b, 32'h3f9e75a0} /* (0, 24, 28) {real, imag} */,
  {32'hbe9b5129, 32'h4000c3b7} /* (0, 24, 27) {real, imag} */,
  {32'hbdb79fef, 32'h40414117} /* (0, 24, 26) {real, imag} */,
  {32'hbfc08261, 32'hbf47815a} /* (0, 24, 25) {real, imag} */,
  {32'hc03ebe8c, 32'h40231263} /* (0, 24, 24) {real, imag} */,
  {32'hc0212afe, 32'hc06e35f7} /* (0, 24, 23) {real, imag} */,
  {32'h3f85ac19, 32'hc091a21b} /* (0, 24, 22) {real, imag} */,
  {32'h40c987e3, 32'h3f83dc3b} /* (0, 24, 21) {real, imag} */,
  {32'h3eb40050, 32'hbf8e99e0} /* (0, 24, 20) {real, imag} */,
  {32'hbffa7b2d, 32'h401a5ba6} /* (0, 24, 19) {real, imag} */,
  {32'h3f445a0a, 32'h3d9938a2} /* (0, 24, 18) {real, imag} */,
  {32'h3e95d038, 32'hc0209094} /* (0, 24, 17) {real, imag} */,
  {32'h3f4ca77d, 32'hbf838dca} /* (0, 24, 16) {real, imag} */,
  {32'hbf1e0646, 32'hbf183e8c} /* (0, 24, 15) {real, imag} */,
  {32'h4003f3e6, 32'hbff2d2f9} /* (0, 24, 14) {real, imag} */,
  {32'hbf834d50, 32'h3f69c7d4} /* (0, 24, 13) {real, imag} */,
  {32'hbf29548b, 32'hbfbd112b} /* (0, 24, 12) {real, imag} */,
  {32'h3f8049d4, 32'hc0505ac4} /* (0, 24, 11) {real, imag} */,
  {32'hc045a64c, 32'h3ff2ebed} /* (0, 24, 10) {real, imag} */,
  {32'h3ffe88de, 32'h3fee2780} /* (0, 24, 9) {real, imag} */,
  {32'hc0043f27, 32'h4026ae6b} /* (0, 24, 8) {real, imag} */,
  {32'h40b5cdc7, 32'h407102a2} /* (0, 24, 7) {real, imag} */,
  {32'h400392e8, 32'hbf889ee9} /* (0, 24, 6) {real, imag} */,
  {32'hc02d788f, 32'h4018fbbb} /* (0, 24, 5) {real, imag} */,
  {32'h403d12b3, 32'hc09fb151} /* (0, 24, 4) {real, imag} */,
  {32'h3fe593e0, 32'h40a1580a} /* (0, 24, 3) {real, imag} */,
  {32'hbf7398f4, 32'hc04ee22f} /* (0, 24, 2) {real, imag} */,
  {32'hc04ff26a, 32'h3f47dbde} /* (0, 24, 1) {real, imag} */,
  {32'hbfd6bf8b, 32'hbebec07b} /* (0, 24, 0) {real, imag} */,
  {32'hc003ed0c, 32'h40b1ba40} /* (0, 23, 31) {real, imag} */,
  {32'hc005b236, 32'h40a47f26} /* (0, 23, 30) {real, imag} */,
  {32'hbf3f8c36, 32'h3fa85006} /* (0, 23, 29) {real, imag} */,
  {32'hbfd04065, 32'h3f2e878d} /* (0, 23, 28) {real, imag} */,
  {32'hbfafbc16, 32'hc0827f1d} /* (0, 23, 27) {real, imag} */,
  {32'hbf9a1077, 32'h3e9dc093} /* (0, 23, 26) {real, imag} */,
  {32'h3f431a89, 32'hc035299e} /* (0, 23, 25) {real, imag} */,
  {32'hbeb41ff5, 32'h3ef88a63} /* (0, 23, 24) {real, imag} */,
  {32'h40193f5d, 32'hc05be6e7} /* (0, 23, 23) {real, imag} */,
  {32'hbf8a827d, 32'h3fc560eb} /* (0, 23, 22) {real, imag} */,
  {32'hc0460cee, 32'hbfd85cfc} /* (0, 23, 21) {real, imag} */,
  {32'hbf0d276d, 32'h3fdf2773} /* (0, 23, 20) {real, imag} */,
  {32'hbfb0f85c, 32'hbf34b9a0} /* (0, 23, 19) {real, imag} */,
  {32'hbf64b5cf, 32'hbf682133} /* (0, 23, 18) {real, imag} */,
  {32'hbe3fb274, 32'h3f3700b1} /* (0, 23, 17) {real, imag} */,
  {32'h40161c5f, 32'hbfe5ae67} /* (0, 23, 16) {real, imag} */,
  {32'hbfc4ef44, 32'hbfcc8ef1} /* (0, 23, 15) {real, imag} */,
  {32'h3f919bed, 32'h3f69823a} /* (0, 23, 14) {real, imag} */,
  {32'h3f50d1c0, 32'hbfa80900} /* (0, 23, 13) {real, imag} */,
  {32'h405b4e5c, 32'h3ce41195} /* (0, 23, 12) {real, imag} */,
  {32'hbff08fa0, 32'h3f0cdabf} /* (0, 23, 11) {real, imag} */,
  {32'hbfc83c59, 32'h3f29009f} /* (0, 23, 10) {real, imag} */,
  {32'hc01ff6ed, 32'hc02dbab1} /* (0, 23, 9) {real, imag} */,
  {32'hbe623b24, 32'h3e5d5f8c} /* (0, 23, 8) {real, imag} */,
  {32'hbef488b8, 32'hbefdf04e} /* (0, 23, 7) {real, imag} */,
  {32'h3eb312d7, 32'hbf0a5446} /* (0, 23, 6) {real, imag} */,
  {32'h3f1acfda, 32'hbf2b7612} /* (0, 23, 5) {real, imag} */,
  {32'hbfc1a8dc, 32'hbebb1841} /* (0, 23, 4) {real, imag} */,
  {32'h3ff211ed, 32'h4005f2e8} /* (0, 23, 3) {real, imag} */,
  {32'h40b83d29, 32'hc0570189} /* (0, 23, 2) {real, imag} */,
  {32'hc098a70f, 32'hc104147b} /* (0, 23, 1) {real, imag} */,
  {32'hc02e824f, 32'h3f530b9a} /* (0, 23, 0) {real, imag} */,
  {32'hbfbca121, 32'h4066ccda} /* (0, 22, 31) {real, imag} */,
  {32'h3fa21564, 32'hbf22c4fa} /* (0, 22, 30) {real, imag} */,
  {32'h3f943743, 32'hbf0b484d} /* (0, 22, 29) {real, imag} */,
  {32'h3f95a3a7, 32'h4005d7c6} /* (0, 22, 28) {real, imag} */,
  {32'hbf9b4551, 32'h3f89926b} /* (0, 22, 27) {real, imag} */,
  {32'hbf6cece4, 32'hbd578750} /* (0, 22, 26) {real, imag} */,
  {32'h40a3fc5f, 32'hbf158b80} /* (0, 22, 25) {real, imag} */,
  {32'hbf0db571, 32'hc0028806} /* (0, 22, 24) {real, imag} */,
  {32'h40094b84, 32'h3fa8268e} /* (0, 22, 23) {real, imag} */,
  {32'hc0004648, 32'hc040c514} /* (0, 22, 22) {real, imag} */,
  {32'h4026b7eb, 32'hbee6da32} /* (0, 22, 21) {real, imag} */,
  {32'hc0ab5ede, 32'hbeea9c86} /* (0, 22, 20) {real, imag} */,
  {32'h3fb6b47b, 32'h40289a2f} /* (0, 22, 19) {real, imag} */,
  {32'h3f848f68, 32'h3f8d6620} /* (0, 22, 18) {real, imag} */,
  {32'hbfaec0fc, 32'hbf6c6bc1} /* (0, 22, 17) {real, imag} */,
  {32'hbf99cf2a, 32'h3e41b7c5} /* (0, 22, 16) {real, imag} */,
  {32'h3f9ffc55, 32'h3e2fa5c9} /* (0, 22, 15) {real, imag} */,
  {32'hbf7172fb, 32'hbf422cfd} /* (0, 22, 14) {real, imag} */,
  {32'h4030bf0f, 32'h3eaa1a2b} /* (0, 22, 13) {real, imag} */,
  {32'h3f30a5b2, 32'hbed00b23} /* (0, 22, 12) {real, imag} */,
  {32'hbd65ee0e, 32'h40985ba8} /* (0, 22, 11) {real, imag} */,
  {32'h3ebcdfd3, 32'hbc834b36} /* (0, 22, 10) {real, imag} */,
  {32'h3f812456, 32'hbf579c25} /* (0, 22, 9) {real, imag} */,
  {32'hbfa66a4a, 32'h3f6e9a72} /* (0, 22, 8) {real, imag} */,
  {32'hc01d3e0c, 32'h3f866038} /* (0, 22, 7) {real, imag} */,
  {32'h3f7adab1, 32'h3dfda713} /* (0, 22, 6) {real, imag} */,
  {32'h40001132, 32'h3f5ccb1d} /* (0, 22, 5) {real, imag} */,
  {32'hc05610c3, 32'h4081acda} /* (0, 22, 4) {real, imag} */,
  {32'hc0ca2bfa, 32'h3fb04689} /* (0, 22, 3) {real, imag} */,
  {32'h3f9448d4, 32'hbedf2370} /* (0, 22, 2) {real, imag} */,
  {32'h3f79417b, 32'hbead3437} /* (0, 22, 1) {real, imag} */,
  {32'hbf7572a3, 32'hbf3a5d2e} /* (0, 22, 0) {real, imag} */,
  {32'hbf0b5aa5, 32'h3ef9e287} /* (0, 21, 31) {real, imag} */,
  {32'hbfcc366b, 32'hbfe81f94} /* (0, 21, 30) {real, imag} */,
  {32'h3fa02f97, 32'h3f931b26} /* (0, 21, 29) {real, imag} */,
  {32'hbfeaf23d, 32'h3fb9f058} /* (0, 21, 28) {real, imag} */,
  {32'hc00a2060, 32'h3d525387} /* (0, 21, 27) {real, imag} */,
  {32'hbfddf3d9, 32'hc0082772} /* (0, 21, 26) {real, imag} */,
  {32'hbfd881f7, 32'hbfebc6da} /* (0, 21, 25) {real, imag} */,
  {32'h3f088186, 32'hbdaa0945} /* (0, 21, 24) {real, imag} */,
  {32'h3fbd3a25, 32'h3fb0085d} /* (0, 21, 23) {real, imag} */,
  {32'hc0278a7f, 32'hbce1fb83} /* (0, 21, 22) {real, imag} */,
  {32'h3fa6a163, 32'h3f151b14} /* (0, 21, 21) {real, imag} */,
  {32'hbf505f2f, 32'h3f9c2a7d} /* (0, 21, 20) {real, imag} */,
  {32'hc0168847, 32'hbe895d89} /* (0, 21, 19) {real, imag} */,
  {32'h3f6c942b, 32'h403756c5} /* (0, 21, 18) {real, imag} */,
  {32'hbddfacd6, 32'hbff501bd} /* (0, 21, 17) {real, imag} */,
  {32'hbfa76150, 32'hc0062393} /* (0, 21, 16) {real, imag} */,
  {32'hbd898143, 32'hbf9b4b9d} /* (0, 21, 15) {real, imag} */,
  {32'hbf350062, 32'h3e1b963c} /* (0, 21, 14) {real, imag} */,
  {32'h3e5c91e9, 32'h3fd98671} /* (0, 21, 13) {real, imag} */,
  {32'h3e99483d, 32'hbf60dda7} /* (0, 21, 12) {real, imag} */,
  {32'h3f369baa, 32'hc069f11b} /* (0, 21, 11) {real, imag} */,
  {32'hbfd475df, 32'hbe41ce8e} /* (0, 21, 10) {real, imag} */,
  {32'h3f2712ab, 32'h40679b98} /* (0, 21, 9) {real, imag} */,
  {32'h3feda6bd, 32'h3f5f2c0e} /* (0, 21, 8) {real, imag} */,
  {32'hbd19b26c, 32'h40074476} /* (0, 21, 7) {real, imag} */,
  {32'h3f31236c, 32'h3fe931af} /* (0, 21, 6) {real, imag} */,
  {32'h3fb072d8, 32'hbdddb78d} /* (0, 21, 5) {real, imag} */,
  {32'hbf64bc80, 32'hbfe03ba0} /* (0, 21, 4) {real, imag} */,
  {32'h3e73ed86, 32'hbf62f11b} /* (0, 21, 3) {real, imag} */,
  {32'h3f5fc23f, 32'h3fbee8ad} /* (0, 21, 2) {real, imag} */,
  {32'h3fa21663, 32'h3e57bfcf} /* (0, 21, 1) {real, imag} */,
  {32'h3e39381c, 32'h40053d4c} /* (0, 21, 0) {real, imag} */,
  {32'h403d375d, 32'hc00968c9} /* (0, 20, 31) {real, imag} */,
  {32'hbf165b68, 32'hbfdf7537} /* (0, 20, 30) {real, imag} */,
  {32'hc0410416, 32'h3fdcdd05} /* (0, 20, 29) {real, imag} */,
  {32'h3ee9789c, 32'h3f98d00f} /* (0, 20, 28) {real, imag} */,
  {32'h3eb5465d, 32'h3f82ea0b} /* (0, 20, 27) {real, imag} */,
  {32'h3e13595c, 32'h3f14a507} /* (0, 20, 26) {real, imag} */,
  {32'hbc5a2faa, 32'h3f7e8aef} /* (0, 20, 25) {real, imag} */,
  {32'h3fa47be7, 32'h3b8fedf2} /* (0, 20, 24) {real, imag} */,
  {32'hbe0fe454, 32'h3fce3528} /* (0, 20, 23) {real, imag} */,
  {32'hbec0d323, 32'hbfb2b7b6} /* (0, 20, 22) {real, imag} */,
  {32'hbeaf5868, 32'hbdeb3cab} /* (0, 20, 21) {real, imag} */,
  {32'h3fbd5b29, 32'hbf81ca87} /* (0, 20, 20) {real, imag} */,
  {32'hc0241bca, 32'h3f3f0201} /* (0, 20, 19) {real, imag} */,
  {32'hbf494fee, 32'h3f5ce554} /* (0, 20, 18) {real, imag} */,
  {32'h3f652aeb, 32'hbfb6c01e} /* (0, 20, 17) {real, imag} */,
  {32'hbf708bfc, 32'h3cdd0eab} /* (0, 20, 16) {real, imag} */,
  {32'h3f7c7665, 32'hbfc2dad2} /* (0, 20, 15) {real, imag} */,
  {32'hc00daf55, 32'hbdfbf8ae} /* (0, 20, 14) {real, imag} */,
  {32'h3fecfb24, 32'hbebeaaa5} /* (0, 20, 13) {real, imag} */,
  {32'h3f9a73b0, 32'hbfadaf78} /* (0, 20, 12) {real, imag} */,
  {32'hc0242d05, 32'hc02c8d32} /* (0, 20, 11) {real, imag} */,
  {32'h40145427, 32'hbe90b128} /* (0, 20, 10) {real, imag} */,
  {32'h3f5dd6fc, 32'h3f1eefbe} /* (0, 20, 9) {real, imag} */,
  {32'hc01e9e8a, 32'hbffa395a} /* (0, 20, 8) {real, imag} */,
  {32'h4015b848, 32'h3f49e1bc} /* (0, 20, 7) {real, imag} */,
  {32'hc0239a1d, 32'h3e3944f1} /* (0, 20, 6) {real, imag} */,
  {32'h3f34d18d, 32'h3f9a7dea} /* (0, 20, 5) {real, imag} */,
  {32'hbf703537, 32'h3faff773} /* (0, 20, 4) {real, imag} */,
  {32'h3ed8f54d, 32'h4008df4e} /* (0, 20, 3) {real, imag} */,
  {32'hbf880b39, 32'hbf1c7d17} /* (0, 20, 2) {real, imag} */,
  {32'h3f0f23d7, 32'hbf66a489} /* (0, 20, 1) {real, imag} */,
  {32'h40730a5b, 32'h402b9cda} /* (0, 20, 0) {real, imag} */,
  {32'h3f09f247, 32'hc04cb612} /* (0, 19, 31) {real, imag} */,
  {32'h401401fe, 32'h3f988bc7} /* (0, 19, 30) {real, imag} */,
  {32'h3f93b1b5, 32'hbffc2a1e} /* (0, 19, 29) {real, imag} */,
  {32'hc03172da, 32'hbe3d10bb} /* (0, 19, 28) {real, imag} */,
  {32'h3e0d4bc7, 32'h3e6168a6} /* (0, 19, 27) {real, imag} */,
  {32'h40194963, 32'h3eba0aff} /* (0, 19, 26) {real, imag} */,
  {32'hbfe4eecc, 32'h3ccde7ff} /* (0, 19, 25) {real, imag} */,
  {32'h4014e6c2, 32'hbf65a74e} /* (0, 19, 24) {real, imag} */,
  {32'hc063256d, 32'hbf70e953} /* (0, 19, 23) {real, imag} */,
  {32'h3f04b8a4, 32'hbfae0993} /* (0, 19, 22) {real, imag} */,
  {32'hc05e18de, 32'h3d863d72} /* (0, 19, 21) {real, imag} */,
  {32'h3f4b6ea0, 32'hbf309075} /* (0, 19, 20) {real, imag} */,
  {32'h3ed7260b, 32'h3f3780b0} /* (0, 19, 19) {real, imag} */,
  {32'h3f4cad3f, 32'h3fc012b8} /* (0, 19, 18) {real, imag} */,
  {32'h3ef3b3c6, 32'h3f823d26} /* (0, 19, 17) {real, imag} */,
  {32'hbf86157c, 32'h3f025429} /* (0, 19, 16) {real, imag} */,
  {32'hbf2ce7c9, 32'h3f2ba610} /* (0, 19, 15) {real, imag} */,
  {32'hbfe1cdd6, 32'h3f927666} /* (0, 19, 14) {real, imag} */,
  {32'h3fdf8b2c, 32'hbff7b0ae} /* (0, 19, 13) {real, imag} */,
  {32'hc018a4ee, 32'h400fe41a} /* (0, 19, 12) {real, imag} */,
  {32'h3ddebfb3, 32'h3f093c3b} /* (0, 19, 11) {real, imag} */,
  {32'h3fc29204, 32'hbffdaa03} /* (0, 19, 10) {real, imag} */,
  {32'h3e8dd9af, 32'hbf3a9b58} /* (0, 19, 9) {real, imag} */,
  {32'h3fa6eb80, 32'h3fec63c4} /* (0, 19, 8) {real, imag} */,
  {32'h4021636b, 32'hbfe1f2c1} /* (0, 19, 7) {real, imag} */,
  {32'hc0197c9b, 32'h400a1869} /* (0, 19, 6) {real, imag} */,
  {32'h3e63244f, 32'h401aa16e} /* (0, 19, 5) {real, imag} */,
  {32'hbf6f83cb, 32'hbea4bad4} /* (0, 19, 4) {real, imag} */,
  {32'hbd5ecd84, 32'hbf2407dc} /* (0, 19, 3) {real, imag} */,
  {32'hc01ad8fc, 32'hbf735fef} /* (0, 19, 2) {real, imag} */,
  {32'hbfb29d87, 32'h40511fc3} /* (0, 19, 1) {real, imag} */,
  {32'hbff10ed4, 32'h3e6911a1} /* (0, 19, 0) {real, imag} */,
  {32'hc063f975, 32'h3fc80936} /* (0, 18, 31) {real, imag} */,
  {32'hbf5636c5, 32'hbde0eb89} /* (0, 18, 30) {real, imag} */,
  {32'h3fcf6106, 32'h3ed84a24} /* (0, 18, 29) {real, imag} */,
  {32'hbfc69bed, 32'h3e94c645} /* (0, 18, 28) {real, imag} */,
  {32'hbf96ed35, 32'hbf018b86} /* (0, 18, 27) {real, imag} */,
  {32'hbea51d2d, 32'hbf87fefa} /* (0, 18, 26) {real, imag} */,
  {32'hc04de13c, 32'h3d17c48e} /* (0, 18, 25) {real, imag} */,
  {32'h40450c57, 32'h3f82daeb} /* (0, 18, 24) {real, imag} */,
  {32'h3fceeadd, 32'hbf7cd1e3} /* (0, 18, 23) {real, imag} */,
  {32'hbece1c1e, 32'h3ca1c7ab} /* (0, 18, 22) {real, imag} */,
  {32'hbe35f0e4, 32'hbf46bfcf} /* (0, 18, 21) {real, imag} */,
  {32'h3f014735, 32'h3f5f4e5b} /* (0, 18, 20) {real, imag} */,
  {32'h3f1f21e0, 32'h4029f1f2} /* (0, 18, 19) {real, imag} */,
  {32'h3ecd0e06, 32'hbf8d60d5} /* (0, 18, 18) {real, imag} */,
  {32'h3f87ee7f, 32'h3eae5016} /* (0, 18, 17) {real, imag} */,
  {32'hbef029f6, 32'h3f8d71d0} /* (0, 18, 16) {real, imag} */,
  {32'h3de4ebf2, 32'hbf8d6cc9} /* (0, 18, 15) {real, imag} */,
  {32'h3f1388a6, 32'hbfcfb9fb} /* (0, 18, 14) {real, imag} */,
  {32'hbf65b450, 32'hbf517e55} /* (0, 18, 13) {real, imag} */,
  {32'h3f68a137, 32'hbef2afc3} /* (0, 18, 12) {real, imag} */,
  {32'h3fb6b84c, 32'h3f50c257} /* (0, 18, 11) {real, imag} */,
  {32'h3ec3b956, 32'h3fa08f88} /* (0, 18, 10) {real, imag} */,
  {32'hbf20609f, 32'h3fd993c1} /* (0, 18, 9) {real, imag} */,
  {32'h3f0c1c0d, 32'h3fbceb62} /* (0, 18, 8) {real, imag} */,
  {32'h3e8d5eba, 32'h3f1f30fe} /* (0, 18, 7) {real, imag} */,
  {32'h3f076b1d, 32'h3bffbb64} /* (0, 18, 6) {real, imag} */,
  {32'hbee1878f, 32'h3eaede0b} /* (0, 18, 5) {real, imag} */,
  {32'h3fc0b120, 32'h3f84ec5b} /* (0, 18, 4) {real, imag} */,
  {32'h400df282, 32'h3f80d782} /* (0, 18, 3) {real, imag} */,
  {32'hbfc43525, 32'hbe6272d9} /* (0, 18, 2) {real, imag} */,
  {32'hbe981b0d, 32'hbfc5f5f9} /* (0, 18, 1) {real, imag} */,
  {32'h3e48acda, 32'hc011c60b} /* (0, 18, 0) {real, imag} */,
  {32'h3f2549eb, 32'h3f0e92ce} /* (0, 17, 31) {real, imag} */,
  {32'h3fdb84cc, 32'h3ed10c0f} /* (0, 17, 30) {real, imag} */,
  {32'h3edad649, 32'h3ee3d909} /* (0, 17, 29) {real, imag} */,
  {32'hbfb8d4f8, 32'h3e931271} /* (0, 17, 28) {real, imag} */,
  {32'hbfd72be9, 32'hbf13e3a9} /* (0, 17, 27) {real, imag} */,
  {32'h3f297a8f, 32'hc00d65f9} /* (0, 17, 26) {real, imag} */,
  {32'h3fa4f360, 32'hbf753992} /* (0, 17, 25) {real, imag} */,
  {32'hbd4243db, 32'hbf9c6287} /* (0, 17, 24) {real, imag} */,
  {32'hbf916ce9, 32'h401ba22f} /* (0, 17, 23) {real, imag} */,
  {32'hbff69fa0, 32'hbf61613a} /* (0, 17, 22) {real, imag} */,
  {32'h3fd779fe, 32'h3fac3c34} /* (0, 17, 21) {real, imag} */,
  {32'h40011151, 32'h3f8e75aa} /* (0, 17, 20) {real, imag} */,
  {32'hbda150a3, 32'h3edc8c0a} /* (0, 17, 19) {real, imag} */,
  {32'h3f422860, 32'h3fad9eea} /* (0, 17, 18) {real, imag} */,
  {32'h3ebe28b1, 32'hbe731591} /* (0, 17, 17) {real, imag} */,
  {32'h3ea0a6e8, 32'h3f8a878a} /* (0, 17, 16) {real, imag} */,
  {32'hbf4b8e93, 32'hbfd59479} /* (0, 17, 15) {real, imag} */,
  {32'h3f143f68, 32'h3f7fffcc} /* (0, 17, 14) {real, imag} */,
  {32'hbee1a008, 32'hbf359e62} /* (0, 17, 13) {real, imag} */,
  {32'hbeffb0d0, 32'hbf3571b5} /* (0, 17, 12) {real, imag} */,
  {32'hbe5adb10, 32'hbef614ec} /* (0, 17, 11) {real, imag} */,
  {32'hbfe85129, 32'hbeeb6165} /* (0, 17, 10) {real, imag} */,
  {32'h3f1332b2, 32'h3f9736b1} /* (0, 17, 9) {real, imag} */,
  {32'h3f037def, 32'hbf01c0a2} /* (0, 17, 8) {real, imag} */,
  {32'hbea1dc9c, 32'h3e7322ec} /* (0, 17, 7) {real, imag} */,
  {32'h3f683f28, 32'hbf93dfd4} /* (0, 17, 6) {real, imag} */,
  {32'hbfbd4e79, 32'hbf1a9a50} /* (0, 17, 5) {real, imag} */,
  {32'h3fd68fb1, 32'h3e3116e1} /* (0, 17, 4) {real, imag} */,
  {32'hbfa222fa, 32'hbfb4d4aa} /* (0, 17, 3) {real, imag} */,
  {32'hbf849b85, 32'hbf485fc3} /* (0, 17, 2) {real, imag} */,
  {32'hbfe3a9f1, 32'h40015baf} /* (0, 17, 1) {real, imag} */,
  {32'h3eac929a, 32'h3e1d2e2e} /* (0, 17, 0) {real, imag} */,
  {32'h3f4b06d3, 32'h3f97c0d6} /* (0, 16, 31) {real, imag} */,
  {32'hbf86ee1b, 32'h3f3fdd68} /* (0, 16, 30) {real, imag} */,
  {32'hbf700f91, 32'h3f7e8f07} /* (0, 16, 29) {real, imag} */,
  {32'h3f54021d, 32'h3d9ac7c1} /* (0, 16, 28) {real, imag} */,
  {32'hbf39f096, 32'hbfd37b22} /* (0, 16, 27) {real, imag} */,
  {32'h3ec69069, 32'hbd6649ec} /* (0, 16, 26) {real, imag} */,
  {32'hbf2022bd, 32'hbec299e7} /* (0, 16, 25) {real, imag} */,
  {32'hbf9642cb, 32'h3f9c73c0} /* (0, 16, 24) {real, imag} */,
  {32'hc00d0417, 32'hbd7279c0} /* (0, 16, 23) {real, imag} */,
  {32'h3e10342c, 32'hbd169681} /* (0, 16, 22) {real, imag} */,
  {32'hbe2d9359, 32'hbf029712} /* (0, 16, 21) {real, imag} */,
  {32'h3f606fd1, 32'hbdef4881} /* (0, 16, 20) {real, imag} */,
  {32'h3e93799c, 32'h3e809cd2} /* (0, 16, 19) {real, imag} */,
  {32'h3fb41f44, 32'hbf8f1398} /* (0, 16, 18) {real, imag} */,
  {32'hbef002b9, 32'hbf5ad715} /* (0, 16, 17) {real, imag} */,
  {32'h3e6c87d2, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hbef002b9, 32'h3f5ad715} /* (0, 16, 15) {real, imag} */,
  {32'h3fb41f44, 32'h3f8f1398} /* (0, 16, 14) {real, imag} */,
  {32'h3e93799c, 32'hbe809cd2} /* (0, 16, 13) {real, imag} */,
  {32'h3f606fd1, 32'h3def4881} /* (0, 16, 12) {real, imag} */,
  {32'hbe2d9359, 32'h3f029712} /* (0, 16, 11) {real, imag} */,
  {32'h3e10342c, 32'h3d169681} /* (0, 16, 10) {real, imag} */,
  {32'hc00d0417, 32'h3d7279c0} /* (0, 16, 9) {real, imag} */,
  {32'hbf9642cb, 32'hbf9c73c0} /* (0, 16, 8) {real, imag} */,
  {32'hbf2022bd, 32'h3ec299e7} /* (0, 16, 7) {real, imag} */,
  {32'h3ec69069, 32'h3d6649ec} /* (0, 16, 6) {real, imag} */,
  {32'hbf39f096, 32'h3fd37b22} /* (0, 16, 5) {real, imag} */,
  {32'h3f54021d, 32'hbd9ac7c1} /* (0, 16, 4) {real, imag} */,
  {32'hbf700f91, 32'hbf7e8f07} /* (0, 16, 3) {real, imag} */,
  {32'hbf86ee1b, 32'hbf3fdd68} /* (0, 16, 2) {real, imag} */,
  {32'h3f4b06d3, 32'hbf97c0d6} /* (0, 16, 1) {real, imag} */,
  {32'h3ff24080, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'hbfe3a9f1, 32'hc0015baf} /* (0, 15, 31) {real, imag} */,
  {32'hbf849b85, 32'h3f485fc3} /* (0, 15, 30) {real, imag} */,
  {32'hbfa222fa, 32'h3fb4d4aa} /* (0, 15, 29) {real, imag} */,
  {32'h3fd68fb1, 32'hbe3116e1} /* (0, 15, 28) {real, imag} */,
  {32'hbfbd4e79, 32'h3f1a9a50} /* (0, 15, 27) {real, imag} */,
  {32'h3f683f28, 32'h3f93dfd4} /* (0, 15, 26) {real, imag} */,
  {32'hbea1dc9c, 32'hbe7322ec} /* (0, 15, 25) {real, imag} */,
  {32'h3f037def, 32'h3f01c0a2} /* (0, 15, 24) {real, imag} */,
  {32'h3f1332b2, 32'hbf9736b1} /* (0, 15, 23) {real, imag} */,
  {32'hbfe85129, 32'h3eeb6165} /* (0, 15, 22) {real, imag} */,
  {32'hbe5adb10, 32'h3ef614ec} /* (0, 15, 21) {real, imag} */,
  {32'hbeffb0d0, 32'h3f3571b5} /* (0, 15, 20) {real, imag} */,
  {32'hbee1a008, 32'h3f359e62} /* (0, 15, 19) {real, imag} */,
  {32'h3f143f68, 32'hbf7fffcc} /* (0, 15, 18) {real, imag} */,
  {32'hbf4b8e93, 32'h3fd59479} /* (0, 15, 17) {real, imag} */,
  {32'h3ea0a6e8, 32'hbf8a878a} /* (0, 15, 16) {real, imag} */,
  {32'h3ebe28b1, 32'h3e731591} /* (0, 15, 15) {real, imag} */,
  {32'h3f422860, 32'hbfad9eea} /* (0, 15, 14) {real, imag} */,
  {32'hbda150a3, 32'hbedc8c0a} /* (0, 15, 13) {real, imag} */,
  {32'h40011151, 32'hbf8e75aa} /* (0, 15, 12) {real, imag} */,
  {32'h3fd779fe, 32'hbfac3c34} /* (0, 15, 11) {real, imag} */,
  {32'hbff69fa0, 32'h3f61613a} /* (0, 15, 10) {real, imag} */,
  {32'hbf916ce9, 32'hc01ba22f} /* (0, 15, 9) {real, imag} */,
  {32'hbd4243db, 32'h3f9c6287} /* (0, 15, 8) {real, imag} */,
  {32'h3fa4f360, 32'h3f753992} /* (0, 15, 7) {real, imag} */,
  {32'h3f297a8f, 32'h400d65f9} /* (0, 15, 6) {real, imag} */,
  {32'hbfd72be9, 32'h3f13e3a9} /* (0, 15, 5) {real, imag} */,
  {32'hbfb8d4f8, 32'hbe931271} /* (0, 15, 4) {real, imag} */,
  {32'h3edad649, 32'hbee3d909} /* (0, 15, 3) {real, imag} */,
  {32'h3fdb84cc, 32'hbed10c0f} /* (0, 15, 2) {real, imag} */,
  {32'h3f2549eb, 32'hbf0e92ce} /* (0, 15, 1) {real, imag} */,
  {32'h3eac929a, 32'hbe1d2e2e} /* (0, 15, 0) {real, imag} */,
  {32'hbe981b0d, 32'h3fc5f5f9} /* (0, 14, 31) {real, imag} */,
  {32'hbfc43525, 32'h3e6272d9} /* (0, 14, 30) {real, imag} */,
  {32'h400df282, 32'hbf80d782} /* (0, 14, 29) {real, imag} */,
  {32'h3fc0b120, 32'hbf84ec5b} /* (0, 14, 28) {real, imag} */,
  {32'hbee1878f, 32'hbeaede0b} /* (0, 14, 27) {real, imag} */,
  {32'h3f076b1d, 32'hbbffbb64} /* (0, 14, 26) {real, imag} */,
  {32'h3e8d5eba, 32'hbf1f30fe} /* (0, 14, 25) {real, imag} */,
  {32'h3f0c1c0d, 32'hbfbceb62} /* (0, 14, 24) {real, imag} */,
  {32'hbf20609f, 32'hbfd993c1} /* (0, 14, 23) {real, imag} */,
  {32'h3ec3b956, 32'hbfa08f88} /* (0, 14, 22) {real, imag} */,
  {32'h3fb6b84c, 32'hbf50c257} /* (0, 14, 21) {real, imag} */,
  {32'h3f68a137, 32'h3ef2afc3} /* (0, 14, 20) {real, imag} */,
  {32'hbf65b450, 32'h3f517e55} /* (0, 14, 19) {real, imag} */,
  {32'h3f1388a6, 32'h3fcfb9fb} /* (0, 14, 18) {real, imag} */,
  {32'h3de4ebf2, 32'h3f8d6cc9} /* (0, 14, 17) {real, imag} */,
  {32'hbef029f6, 32'hbf8d71d0} /* (0, 14, 16) {real, imag} */,
  {32'h3f87ee7f, 32'hbeae5016} /* (0, 14, 15) {real, imag} */,
  {32'h3ecd0e06, 32'h3f8d60d5} /* (0, 14, 14) {real, imag} */,
  {32'h3f1f21e0, 32'hc029f1f2} /* (0, 14, 13) {real, imag} */,
  {32'h3f014735, 32'hbf5f4e5b} /* (0, 14, 12) {real, imag} */,
  {32'hbe35f0e4, 32'h3f46bfcf} /* (0, 14, 11) {real, imag} */,
  {32'hbece1c1e, 32'hbca1c7ab} /* (0, 14, 10) {real, imag} */,
  {32'h3fceeadd, 32'h3f7cd1e3} /* (0, 14, 9) {real, imag} */,
  {32'h40450c57, 32'hbf82daeb} /* (0, 14, 8) {real, imag} */,
  {32'hc04de13c, 32'hbd17c48e} /* (0, 14, 7) {real, imag} */,
  {32'hbea51d2d, 32'h3f87fefa} /* (0, 14, 6) {real, imag} */,
  {32'hbf96ed35, 32'h3f018b86} /* (0, 14, 5) {real, imag} */,
  {32'hbfc69bed, 32'hbe94c645} /* (0, 14, 4) {real, imag} */,
  {32'h3fcf6106, 32'hbed84a24} /* (0, 14, 3) {real, imag} */,
  {32'hbf5636c5, 32'h3de0eb89} /* (0, 14, 2) {real, imag} */,
  {32'hc063f975, 32'hbfc80936} /* (0, 14, 1) {real, imag} */,
  {32'h3e48acda, 32'h4011c60b} /* (0, 14, 0) {real, imag} */,
  {32'hbfb29d87, 32'hc0511fc3} /* (0, 13, 31) {real, imag} */,
  {32'hc01ad8fc, 32'h3f735fef} /* (0, 13, 30) {real, imag} */,
  {32'hbd5ecd84, 32'h3f2407dc} /* (0, 13, 29) {real, imag} */,
  {32'hbf6f83cb, 32'h3ea4bad4} /* (0, 13, 28) {real, imag} */,
  {32'h3e63244f, 32'hc01aa16e} /* (0, 13, 27) {real, imag} */,
  {32'hc0197c9b, 32'hc00a1869} /* (0, 13, 26) {real, imag} */,
  {32'h4021636b, 32'h3fe1f2c1} /* (0, 13, 25) {real, imag} */,
  {32'h3fa6eb80, 32'hbfec63c4} /* (0, 13, 24) {real, imag} */,
  {32'h3e8dd9af, 32'h3f3a9b58} /* (0, 13, 23) {real, imag} */,
  {32'h3fc29204, 32'h3ffdaa03} /* (0, 13, 22) {real, imag} */,
  {32'h3ddebfb3, 32'hbf093c3b} /* (0, 13, 21) {real, imag} */,
  {32'hc018a4ee, 32'hc00fe41a} /* (0, 13, 20) {real, imag} */,
  {32'h3fdf8b2c, 32'h3ff7b0ae} /* (0, 13, 19) {real, imag} */,
  {32'hbfe1cdd6, 32'hbf927666} /* (0, 13, 18) {real, imag} */,
  {32'hbf2ce7c9, 32'hbf2ba610} /* (0, 13, 17) {real, imag} */,
  {32'hbf86157c, 32'hbf025429} /* (0, 13, 16) {real, imag} */,
  {32'h3ef3b3c6, 32'hbf823d26} /* (0, 13, 15) {real, imag} */,
  {32'h3f4cad3f, 32'hbfc012b8} /* (0, 13, 14) {real, imag} */,
  {32'h3ed7260b, 32'hbf3780b0} /* (0, 13, 13) {real, imag} */,
  {32'h3f4b6ea0, 32'h3f309075} /* (0, 13, 12) {real, imag} */,
  {32'hc05e18de, 32'hbd863d72} /* (0, 13, 11) {real, imag} */,
  {32'h3f04b8a4, 32'h3fae0993} /* (0, 13, 10) {real, imag} */,
  {32'hc063256d, 32'h3f70e953} /* (0, 13, 9) {real, imag} */,
  {32'h4014e6c2, 32'h3f65a74e} /* (0, 13, 8) {real, imag} */,
  {32'hbfe4eecc, 32'hbccde7ff} /* (0, 13, 7) {real, imag} */,
  {32'h40194963, 32'hbeba0aff} /* (0, 13, 6) {real, imag} */,
  {32'h3e0d4bc7, 32'hbe6168a6} /* (0, 13, 5) {real, imag} */,
  {32'hc03172da, 32'h3e3d10bb} /* (0, 13, 4) {real, imag} */,
  {32'h3f93b1b5, 32'h3ffc2a1e} /* (0, 13, 3) {real, imag} */,
  {32'h401401fe, 32'hbf988bc7} /* (0, 13, 2) {real, imag} */,
  {32'h3f09f247, 32'h404cb612} /* (0, 13, 1) {real, imag} */,
  {32'hbff10ed4, 32'hbe6911a1} /* (0, 13, 0) {real, imag} */,
  {32'h3f0f23d7, 32'h3f66a489} /* (0, 12, 31) {real, imag} */,
  {32'hbf880b39, 32'h3f1c7d17} /* (0, 12, 30) {real, imag} */,
  {32'h3ed8f54d, 32'hc008df4e} /* (0, 12, 29) {real, imag} */,
  {32'hbf703537, 32'hbfaff773} /* (0, 12, 28) {real, imag} */,
  {32'h3f34d18d, 32'hbf9a7dea} /* (0, 12, 27) {real, imag} */,
  {32'hc0239a1d, 32'hbe3944f1} /* (0, 12, 26) {real, imag} */,
  {32'h4015b848, 32'hbf49e1bc} /* (0, 12, 25) {real, imag} */,
  {32'hc01e9e8a, 32'h3ffa395a} /* (0, 12, 24) {real, imag} */,
  {32'h3f5dd6fc, 32'hbf1eefbe} /* (0, 12, 23) {real, imag} */,
  {32'h40145427, 32'h3e90b128} /* (0, 12, 22) {real, imag} */,
  {32'hc0242d05, 32'h402c8d32} /* (0, 12, 21) {real, imag} */,
  {32'h3f9a73b0, 32'h3fadaf78} /* (0, 12, 20) {real, imag} */,
  {32'h3fecfb24, 32'h3ebeaaa5} /* (0, 12, 19) {real, imag} */,
  {32'hc00daf55, 32'h3dfbf8ae} /* (0, 12, 18) {real, imag} */,
  {32'h3f7c7665, 32'h3fc2dad2} /* (0, 12, 17) {real, imag} */,
  {32'hbf708bfc, 32'hbcdd0eab} /* (0, 12, 16) {real, imag} */,
  {32'h3f652aeb, 32'h3fb6c01e} /* (0, 12, 15) {real, imag} */,
  {32'hbf494fee, 32'hbf5ce554} /* (0, 12, 14) {real, imag} */,
  {32'hc0241bca, 32'hbf3f0201} /* (0, 12, 13) {real, imag} */,
  {32'h3fbd5b29, 32'h3f81ca87} /* (0, 12, 12) {real, imag} */,
  {32'hbeaf5868, 32'h3deb3cab} /* (0, 12, 11) {real, imag} */,
  {32'hbec0d323, 32'h3fb2b7b6} /* (0, 12, 10) {real, imag} */,
  {32'hbe0fe454, 32'hbfce3528} /* (0, 12, 9) {real, imag} */,
  {32'h3fa47be7, 32'hbb8fedf2} /* (0, 12, 8) {real, imag} */,
  {32'hbc5a2faa, 32'hbf7e8aef} /* (0, 12, 7) {real, imag} */,
  {32'h3e13595c, 32'hbf14a507} /* (0, 12, 6) {real, imag} */,
  {32'h3eb5465d, 32'hbf82ea0b} /* (0, 12, 5) {real, imag} */,
  {32'h3ee9789c, 32'hbf98d00f} /* (0, 12, 4) {real, imag} */,
  {32'hc0410416, 32'hbfdcdd05} /* (0, 12, 3) {real, imag} */,
  {32'hbf165b68, 32'h3fdf7537} /* (0, 12, 2) {real, imag} */,
  {32'h403d375d, 32'h400968c9} /* (0, 12, 1) {real, imag} */,
  {32'h40730a5b, 32'hc02b9cda} /* (0, 12, 0) {real, imag} */,
  {32'h3fa21663, 32'hbe57bfcf} /* (0, 11, 31) {real, imag} */,
  {32'h3f5fc23f, 32'hbfbee8ad} /* (0, 11, 30) {real, imag} */,
  {32'h3e73ed86, 32'h3f62f11b} /* (0, 11, 29) {real, imag} */,
  {32'hbf64bc80, 32'h3fe03ba0} /* (0, 11, 28) {real, imag} */,
  {32'h3fb072d8, 32'h3dddb78d} /* (0, 11, 27) {real, imag} */,
  {32'h3f31236c, 32'hbfe931af} /* (0, 11, 26) {real, imag} */,
  {32'hbd19b26c, 32'hc0074476} /* (0, 11, 25) {real, imag} */,
  {32'h3feda6bd, 32'hbf5f2c0e} /* (0, 11, 24) {real, imag} */,
  {32'h3f2712ab, 32'hc0679b98} /* (0, 11, 23) {real, imag} */,
  {32'hbfd475df, 32'h3e41ce8e} /* (0, 11, 22) {real, imag} */,
  {32'h3f369baa, 32'h4069f11b} /* (0, 11, 21) {real, imag} */,
  {32'h3e99483d, 32'h3f60dda7} /* (0, 11, 20) {real, imag} */,
  {32'h3e5c91e9, 32'hbfd98671} /* (0, 11, 19) {real, imag} */,
  {32'hbf350062, 32'hbe1b963c} /* (0, 11, 18) {real, imag} */,
  {32'hbd898143, 32'h3f9b4b9d} /* (0, 11, 17) {real, imag} */,
  {32'hbfa76150, 32'h40062393} /* (0, 11, 16) {real, imag} */,
  {32'hbddfacd6, 32'h3ff501bd} /* (0, 11, 15) {real, imag} */,
  {32'h3f6c942b, 32'hc03756c5} /* (0, 11, 14) {real, imag} */,
  {32'hc0168847, 32'h3e895d89} /* (0, 11, 13) {real, imag} */,
  {32'hbf505f2f, 32'hbf9c2a7d} /* (0, 11, 12) {real, imag} */,
  {32'h3fa6a163, 32'hbf151b14} /* (0, 11, 11) {real, imag} */,
  {32'hc0278a7f, 32'h3ce1fb83} /* (0, 11, 10) {real, imag} */,
  {32'h3fbd3a25, 32'hbfb0085d} /* (0, 11, 9) {real, imag} */,
  {32'h3f088186, 32'h3daa0945} /* (0, 11, 8) {real, imag} */,
  {32'hbfd881f7, 32'h3febc6da} /* (0, 11, 7) {real, imag} */,
  {32'hbfddf3d9, 32'h40082772} /* (0, 11, 6) {real, imag} */,
  {32'hc00a2060, 32'hbd525387} /* (0, 11, 5) {real, imag} */,
  {32'hbfeaf23d, 32'hbfb9f058} /* (0, 11, 4) {real, imag} */,
  {32'h3fa02f97, 32'hbf931b26} /* (0, 11, 3) {real, imag} */,
  {32'hbfcc366b, 32'h3fe81f94} /* (0, 11, 2) {real, imag} */,
  {32'hbf0b5aa5, 32'hbef9e287} /* (0, 11, 1) {real, imag} */,
  {32'h3e39381c, 32'hc0053d4c} /* (0, 11, 0) {real, imag} */,
  {32'h3f79417b, 32'h3ead3437} /* (0, 10, 31) {real, imag} */,
  {32'h3f9448d4, 32'h3edf2370} /* (0, 10, 30) {real, imag} */,
  {32'hc0ca2bfa, 32'hbfb04689} /* (0, 10, 29) {real, imag} */,
  {32'hc05610c3, 32'hc081acda} /* (0, 10, 28) {real, imag} */,
  {32'h40001132, 32'hbf5ccb1d} /* (0, 10, 27) {real, imag} */,
  {32'h3f7adab1, 32'hbdfda713} /* (0, 10, 26) {real, imag} */,
  {32'hc01d3e0c, 32'hbf866038} /* (0, 10, 25) {real, imag} */,
  {32'hbfa66a4a, 32'hbf6e9a72} /* (0, 10, 24) {real, imag} */,
  {32'h3f812456, 32'h3f579c25} /* (0, 10, 23) {real, imag} */,
  {32'h3ebcdfd3, 32'h3c834b36} /* (0, 10, 22) {real, imag} */,
  {32'hbd65ee0e, 32'hc0985ba8} /* (0, 10, 21) {real, imag} */,
  {32'h3f30a5b2, 32'h3ed00b23} /* (0, 10, 20) {real, imag} */,
  {32'h4030bf0f, 32'hbeaa1a2b} /* (0, 10, 19) {real, imag} */,
  {32'hbf7172fb, 32'h3f422cfd} /* (0, 10, 18) {real, imag} */,
  {32'h3f9ffc55, 32'hbe2fa5c9} /* (0, 10, 17) {real, imag} */,
  {32'hbf99cf2a, 32'hbe41b7c5} /* (0, 10, 16) {real, imag} */,
  {32'hbfaec0fc, 32'h3f6c6bc1} /* (0, 10, 15) {real, imag} */,
  {32'h3f848f68, 32'hbf8d6620} /* (0, 10, 14) {real, imag} */,
  {32'h3fb6b47b, 32'hc0289a2f} /* (0, 10, 13) {real, imag} */,
  {32'hc0ab5ede, 32'h3eea9c86} /* (0, 10, 12) {real, imag} */,
  {32'h4026b7eb, 32'h3ee6da32} /* (0, 10, 11) {real, imag} */,
  {32'hc0004648, 32'h4040c514} /* (0, 10, 10) {real, imag} */,
  {32'h40094b84, 32'hbfa8268e} /* (0, 10, 9) {real, imag} */,
  {32'hbf0db571, 32'h40028806} /* (0, 10, 8) {real, imag} */,
  {32'h40a3fc5f, 32'h3f158b80} /* (0, 10, 7) {real, imag} */,
  {32'hbf6cece4, 32'h3d578750} /* (0, 10, 6) {real, imag} */,
  {32'hbf9b4551, 32'hbf89926b} /* (0, 10, 5) {real, imag} */,
  {32'h3f95a3a7, 32'hc005d7c6} /* (0, 10, 4) {real, imag} */,
  {32'h3f943743, 32'h3f0b484d} /* (0, 10, 3) {real, imag} */,
  {32'h3fa21564, 32'h3f22c4fa} /* (0, 10, 2) {real, imag} */,
  {32'hbfbca121, 32'hc066ccda} /* (0, 10, 1) {real, imag} */,
  {32'hbf7572a3, 32'h3f3a5d2e} /* (0, 10, 0) {real, imag} */,
  {32'hc098a70f, 32'h4104147b} /* (0, 9, 31) {real, imag} */,
  {32'h40b83d29, 32'h40570189} /* (0, 9, 30) {real, imag} */,
  {32'h3ff211ed, 32'hc005f2e8} /* (0, 9, 29) {real, imag} */,
  {32'hbfc1a8dc, 32'h3ebb1841} /* (0, 9, 28) {real, imag} */,
  {32'h3f1acfda, 32'h3f2b7612} /* (0, 9, 27) {real, imag} */,
  {32'h3eb312d7, 32'h3f0a5446} /* (0, 9, 26) {real, imag} */,
  {32'hbef488b8, 32'h3efdf04e} /* (0, 9, 25) {real, imag} */,
  {32'hbe623b24, 32'hbe5d5f8c} /* (0, 9, 24) {real, imag} */,
  {32'hc01ff6ed, 32'h402dbab1} /* (0, 9, 23) {real, imag} */,
  {32'hbfc83c59, 32'hbf29009f} /* (0, 9, 22) {real, imag} */,
  {32'hbff08fa0, 32'hbf0cdabf} /* (0, 9, 21) {real, imag} */,
  {32'h405b4e5c, 32'hbce41195} /* (0, 9, 20) {real, imag} */,
  {32'h3f50d1c0, 32'h3fa80900} /* (0, 9, 19) {real, imag} */,
  {32'h3f919bed, 32'hbf69823a} /* (0, 9, 18) {real, imag} */,
  {32'hbfc4ef44, 32'h3fcc8ef1} /* (0, 9, 17) {real, imag} */,
  {32'h40161c5f, 32'h3fe5ae67} /* (0, 9, 16) {real, imag} */,
  {32'hbe3fb274, 32'hbf3700b1} /* (0, 9, 15) {real, imag} */,
  {32'hbf64b5cf, 32'h3f682133} /* (0, 9, 14) {real, imag} */,
  {32'hbfb0f85c, 32'h3f34b9a0} /* (0, 9, 13) {real, imag} */,
  {32'hbf0d276d, 32'hbfdf2773} /* (0, 9, 12) {real, imag} */,
  {32'hc0460cee, 32'h3fd85cfc} /* (0, 9, 11) {real, imag} */,
  {32'hbf8a827d, 32'hbfc560eb} /* (0, 9, 10) {real, imag} */,
  {32'h40193f5d, 32'h405be6e7} /* (0, 9, 9) {real, imag} */,
  {32'hbeb41ff5, 32'hbef88a63} /* (0, 9, 8) {real, imag} */,
  {32'h3f431a89, 32'h4035299e} /* (0, 9, 7) {real, imag} */,
  {32'hbf9a1077, 32'hbe9dc093} /* (0, 9, 6) {real, imag} */,
  {32'hbfafbc16, 32'h40827f1d} /* (0, 9, 5) {real, imag} */,
  {32'hbfd04065, 32'hbf2e878d} /* (0, 9, 4) {real, imag} */,
  {32'hbf3f8c36, 32'hbfa85006} /* (0, 9, 3) {real, imag} */,
  {32'hc005b236, 32'hc0a47f26} /* (0, 9, 2) {real, imag} */,
  {32'hc003ed0c, 32'hc0b1ba40} /* (0, 9, 1) {real, imag} */,
  {32'hc02e824f, 32'hbf530b9a} /* (0, 9, 0) {real, imag} */,
  {32'hc04ff26a, 32'hbf47dbde} /* (0, 8, 31) {real, imag} */,
  {32'hbf7398f4, 32'h404ee22f} /* (0, 8, 30) {real, imag} */,
  {32'h3fe593e0, 32'hc0a1580a} /* (0, 8, 29) {real, imag} */,
  {32'h403d12b3, 32'h409fb151} /* (0, 8, 28) {real, imag} */,
  {32'hc02d788f, 32'hc018fbbb} /* (0, 8, 27) {real, imag} */,
  {32'h400392e8, 32'h3f889ee9} /* (0, 8, 26) {real, imag} */,
  {32'h40b5cdc7, 32'hc07102a2} /* (0, 8, 25) {real, imag} */,
  {32'hc0043f27, 32'hc026ae6b} /* (0, 8, 24) {real, imag} */,
  {32'h3ffe88de, 32'hbfee2780} /* (0, 8, 23) {real, imag} */,
  {32'hc045a64c, 32'hbff2ebed} /* (0, 8, 22) {real, imag} */,
  {32'h3f8049d4, 32'h40505ac4} /* (0, 8, 21) {real, imag} */,
  {32'hbf29548b, 32'h3fbd112b} /* (0, 8, 20) {real, imag} */,
  {32'hbf834d50, 32'hbf69c7d4} /* (0, 8, 19) {real, imag} */,
  {32'h4003f3e6, 32'h3ff2d2f9} /* (0, 8, 18) {real, imag} */,
  {32'hbf1e0646, 32'h3f183e8c} /* (0, 8, 17) {real, imag} */,
  {32'h3f4ca77d, 32'h3f838dca} /* (0, 8, 16) {real, imag} */,
  {32'h3e95d038, 32'h40209094} /* (0, 8, 15) {real, imag} */,
  {32'h3f445a0a, 32'hbd9938a2} /* (0, 8, 14) {real, imag} */,
  {32'hbffa7b2d, 32'hc01a5ba6} /* (0, 8, 13) {real, imag} */,
  {32'h3eb40050, 32'h3f8e99e0} /* (0, 8, 12) {real, imag} */,
  {32'h40c987e3, 32'hbf83dc3b} /* (0, 8, 11) {real, imag} */,
  {32'h3f85ac19, 32'h4091a21b} /* (0, 8, 10) {real, imag} */,
  {32'hc0212afe, 32'h406e35f7} /* (0, 8, 9) {real, imag} */,
  {32'hc03ebe8c, 32'hc0231263} /* (0, 8, 8) {real, imag} */,
  {32'hbfc08261, 32'h3f47815a} /* (0, 8, 7) {real, imag} */,
  {32'hbdb79fef, 32'hc0414117} /* (0, 8, 6) {real, imag} */,
  {32'hbe9b5129, 32'hc000c3b7} /* (0, 8, 5) {real, imag} */,
  {32'hc065630b, 32'hbf9e75a0} /* (0, 8, 4) {real, imag} */,
  {32'hc00b6a96, 32'h409693bf} /* (0, 8, 3) {real, imag} */,
  {32'hbf0a2c66, 32'hbfe2c54f} /* (0, 8, 2) {real, imag} */,
  {32'hc05321a3, 32'hbef83046} /* (0, 8, 1) {real, imag} */,
  {32'hbfd6bf8b, 32'h3ebec07b} /* (0, 8, 0) {real, imag} */,
  {32'hc072cf9d, 32'h3ea550e2} /* (0, 7, 31) {real, imag} */,
  {32'h3ed78b1a, 32'hc0ae77da} /* (0, 7, 30) {real, imag} */,
  {32'hc08603bb, 32'h3e4e791b} /* (0, 7, 29) {real, imag} */,
  {32'hc0d7acd5, 32'h3e84aa25} /* (0, 7, 28) {real, imag} */,
  {32'hc04f4c18, 32'h40bc1989} /* (0, 7, 27) {real, imag} */,
  {32'hc01d4b3c, 32'h3f2fd070} /* (0, 7, 26) {real, imag} */,
  {32'hbeb2c180, 32'h3f7ec762} /* (0, 7, 25) {real, imag} */,
  {32'hbff0e9f0, 32'hc042bf12} /* (0, 7, 24) {real, imag} */,
  {32'hc0377d9c, 32'h40ad1d62} /* (0, 7, 23) {real, imag} */,
  {32'hbdc5b9dd, 32'h40470058} /* (0, 7, 22) {real, imag} */,
  {32'h401deedf, 32'h3fed02e2} /* (0, 7, 21) {real, imag} */,
  {32'h3fc57e48, 32'hbff13d57} /* (0, 7, 20) {real, imag} */,
  {32'h3cd5ce75, 32'h403d7f0e} /* (0, 7, 19) {real, imag} */,
  {32'hbeca7955, 32'hbf89a9fa} /* (0, 7, 18) {real, imag} */,
  {32'h3ec237b4, 32'hbe8e9d07} /* (0, 7, 17) {real, imag} */,
  {32'h3f5c5cae, 32'h3ee8d40f} /* (0, 7, 16) {real, imag} */,
  {32'hbf84df0d, 32'h3fa43aa5} /* (0, 7, 15) {real, imag} */,
  {32'hc014188c, 32'h3dda7ec1} /* (0, 7, 14) {real, imag} */,
  {32'hbfb4fdb1, 32'h3facf7a3} /* (0, 7, 13) {real, imag} */,
  {32'hc009b319, 32'hbeb1b2ad} /* (0, 7, 12) {real, imag} */,
  {32'hbf2aeeb6, 32'h3f757ad9} /* (0, 7, 11) {real, imag} */,
  {32'hbf8ca5f1, 32'h405be771} /* (0, 7, 10) {real, imag} */,
  {32'h4035d1b3, 32'h403c9236} /* (0, 7, 9) {real, imag} */,
  {32'hbdfd6182, 32'hc052c8af} /* (0, 7, 8) {real, imag} */,
  {32'hc020d1e5, 32'hbfb4e2e7} /* (0, 7, 7) {real, imag} */,
  {32'h409b5a64, 32'hc027fbd2} /* (0, 7, 6) {real, imag} */,
  {32'h405babba, 32'h3ff65751} /* (0, 7, 5) {real, imag} */,
  {32'h407014ac, 32'h3ed1aa06} /* (0, 7, 4) {real, imag} */,
  {32'hbeb195c9, 32'h40c86e82} /* (0, 7, 3) {real, imag} */,
  {32'hbe6586ec, 32'hbf812cc5} /* (0, 7, 2) {real, imag} */,
  {32'h3fcf3406, 32'h3fd669e7} /* (0, 7, 1) {real, imag} */,
  {32'h3e858e63, 32'hc074f16f} /* (0, 7, 0) {real, imag} */,
  {32'h4019db63, 32'h40aa3711} /* (0, 6, 31) {real, imag} */,
  {32'hc047f3b0, 32'hbf98a75f} /* (0, 6, 30) {real, imag} */,
  {32'h3f2fbc5b, 32'hc0abc257} /* (0, 6, 29) {real, imag} */,
  {32'h3f8fe3bf, 32'hc093c62b} /* (0, 6, 28) {real, imag} */,
  {32'hbf4c4dd2, 32'hbf2604ed} /* (0, 6, 27) {real, imag} */,
  {32'h3fe67c28, 32'h405dd231} /* (0, 6, 26) {real, imag} */,
  {32'hbf9d3804, 32'h3ecea8be} /* (0, 6, 25) {real, imag} */,
  {32'hc01f4568, 32'h3e893062} /* (0, 6, 24) {real, imag} */,
  {32'h3ff88905, 32'h40136e17} /* (0, 6, 23) {real, imag} */,
  {32'h4049b156, 32'hbdb69013} /* (0, 6, 22) {real, imag} */,
  {32'hbffb7cda, 32'hbf5fb73c} /* (0, 6, 21) {real, imag} */,
  {32'hbe6ed7cc, 32'hbf15b311} /* (0, 6, 20) {real, imag} */,
  {32'hbea1ff68, 32'hbfe5f628} /* (0, 6, 19) {real, imag} */,
  {32'h4018c91c, 32'h3f8bc7f9} /* (0, 6, 18) {real, imag} */,
  {32'h3cc341ee, 32'hc02f0de9} /* (0, 6, 17) {real, imag} */,
  {32'hbf101065, 32'hbf70a0d1} /* (0, 6, 16) {real, imag} */,
  {32'h3e13548b, 32'hbe303161} /* (0, 6, 15) {real, imag} */,
  {32'hbe9959d4, 32'h3f267d93} /* (0, 6, 14) {real, imag} */,
  {32'h4014a7f3, 32'hbfba3aca} /* (0, 6, 13) {real, imag} */,
  {32'h3eeb1e92, 32'h3eec9967} /* (0, 6, 12) {real, imag} */,
  {32'hbe0d73dc, 32'h3f03fd4b} /* (0, 6, 11) {real, imag} */,
  {32'hbfeabb08, 32'h3f64afd8} /* (0, 6, 10) {real, imag} */,
  {32'hbf1d1340, 32'h4034fcd8} /* (0, 6, 9) {real, imag} */,
  {32'hbfdf3f5a, 32'hc0580e54} /* (0, 6, 8) {real, imag} */,
  {32'h407805ef, 32'h40b108f9} /* (0, 6, 7) {real, imag} */,
  {32'hc019fe20, 32'hc002589e} /* (0, 6, 6) {real, imag} */,
  {32'hbe8ff9e5, 32'h3d73742e} /* (0, 6, 5) {real, imag} */,
  {32'h402f246c, 32'h3e8e8801} /* (0, 6, 4) {real, imag} */,
  {32'h40012bc6, 32'hbfc83499} /* (0, 6, 3) {real, imag} */,
  {32'h3eb0490e, 32'hc048cdb4} /* (0, 6, 2) {real, imag} */,
  {32'hc041104c, 32'h3f92e5d8} /* (0, 6, 1) {real, imag} */,
  {32'h406f10b5, 32'hbdeea6e3} /* (0, 6, 0) {real, imag} */,
  {32'h3f326234, 32'h40881df2} /* (0, 5, 31) {real, imag} */,
  {32'hc128ceb0, 32'hc0e635ad} /* (0, 5, 30) {real, imag} */,
  {32'h403be311, 32'h4012f43f} /* (0, 5, 29) {real, imag} */,
  {32'hc0977a69, 32'h408791ea} /* (0, 5, 28) {real, imag} */,
  {32'hbf5a4c16, 32'h40957f79} /* (0, 5, 27) {real, imag} */,
  {32'h3f5c8a67, 32'h4030f554} /* (0, 5, 26) {real, imag} */,
  {32'hbfacfc53, 32'h4047aa9f} /* (0, 5, 25) {real, imag} */,
  {32'hc057cdc8, 32'hbfe4b142} /* (0, 5, 24) {real, imag} */,
  {32'hbf010320, 32'h401ae8cb} /* (0, 5, 23) {real, imag} */,
  {32'hc05ed478, 32'hbe71db53} /* (0, 5, 22) {real, imag} */,
  {32'h3dcb499f, 32'hc03d36d7} /* (0, 5, 21) {real, imag} */,
  {32'h3f2fde6d, 32'hc05598d2} /* (0, 5, 20) {real, imag} */,
  {32'hbea3c10f, 32'h3fa89c17} /* (0, 5, 19) {real, imag} */,
  {32'hbf8cc1cb, 32'h3f91a24f} /* (0, 5, 18) {real, imag} */,
  {32'hbf8666a0, 32'hbfbfe5da} /* (0, 5, 17) {real, imag} */,
  {32'hbf9a452c, 32'hbe3922eb} /* (0, 5, 16) {real, imag} */,
  {32'hbf992a27, 32'h3ed9ce83} /* (0, 5, 15) {real, imag} */,
  {32'hbf807abb, 32'h3fe8a724} /* (0, 5, 14) {real, imag} */,
  {32'h3fe2501d, 32'h3fa9306a} /* (0, 5, 13) {real, imag} */,
  {32'h3fa0b29f, 32'hc031cf5b} /* (0, 5, 12) {real, imag} */,
  {32'hbf977e36, 32'hc090550a} /* (0, 5, 11) {real, imag} */,
  {32'h3e230203, 32'h3fdab27f} /* (0, 5, 10) {real, imag} */,
  {32'h3f912700, 32'hbfa51f0c} /* (0, 5, 9) {real, imag} */,
  {32'h4063f0fa, 32'h4031a8e2} /* (0, 5, 8) {real, imag} */,
  {32'h40477e0e, 32'h3ff7d3f3} /* (0, 5, 7) {real, imag} */,
  {32'hbf475c54, 32'h3f9b86bd} /* (0, 5, 6) {real, imag} */,
  {32'h3ff541dc, 32'h402beb55} /* (0, 5, 5) {real, imag} */,
  {32'hbf84c375, 32'h403579ac} /* (0, 5, 4) {real, imag} */,
  {32'hc02141eb, 32'hc088ba7f} /* (0, 5, 3) {real, imag} */,
  {32'h40bddc69, 32'hc01afe34} /* (0, 5, 2) {real, imag} */,
  {32'h3f4eceb3, 32'h4131b135} /* (0, 5, 1) {real, imag} */,
  {32'hc0ca53d9, 32'h40e552a7} /* (0, 5, 0) {real, imag} */,
  {32'hbf902fe7, 32'hc1383efd} /* (0, 4, 31) {real, imag} */,
  {32'hc167492f, 32'h4108c3ce} /* (0, 4, 30) {real, imag} */,
  {32'hc0e912d9, 32'hc05d6cd3} /* (0, 4, 29) {real, imag} */,
  {32'hc015b0d0, 32'hbf73a440} /* (0, 4, 28) {real, imag} */,
  {32'h3f59c75a, 32'hc0edbcdb} /* (0, 4, 27) {real, imag} */,
  {32'hc0d543af, 32'hc0608da2} /* (0, 4, 26) {real, imag} */,
  {32'h3fca95c4, 32'h40cc5e62} /* (0, 4, 25) {real, imag} */,
  {32'h40b54d14, 32'hc0cfd3ac} /* (0, 4, 24) {real, imag} */,
  {32'hbfee3f4e, 32'hc0550856} /* (0, 4, 23) {real, imag} */,
  {32'hbf5908b1, 32'h3ee0e833} /* (0, 4, 22) {real, imag} */,
  {32'h3f330768, 32'h3ffdbbd6} /* (0, 4, 21) {real, imag} */,
  {32'h40573fe8, 32'h3fd50a08} /* (0, 4, 20) {real, imag} */,
  {32'hbfd02fca, 32'hbf88b862} /* (0, 4, 19) {real, imag} */,
  {32'hbf1bc6cd, 32'hbfbc6aaa} /* (0, 4, 18) {real, imag} */,
  {32'h3f76d61d, 32'h3f8878a2} /* (0, 4, 17) {real, imag} */,
  {32'hbfb4279f, 32'h3f71540b} /* (0, 4, 16) {real, imag} */,
  {32'hbfe33f35, 32'hbf5908ce} /* (0, 4, 15) {real, imag} */,
  {32'hbd16685e, 32'h3f0ee4e9} /* (0, 4, 14) {real, imag} */,
  {32'h40237b6c, 32'h3ff02f88} /* (0, 4, 13) {real, imag} */,
  {32'hc03d8214, 32'hbfc19829} /* (0, 4, 12) {real, imag} */,
  {32'h40521539, 32'h403df432} /* (0, 4, 11) {real, imag} */,
  {32'h3fd78dc5, 32'h3e7cb19c} /* (0, 4, 10) {real, imag} */,
  {32'h405c582f, 32'hbfde0cea} /* (0, 4, 9) {real, imag} */,
  {32'h3f905208, 32'hbf6a05bf} /* (0, 4, 8) {real, imag} */,
  {32'hc0be99d3, 32'hbf759371} /* (0, 4, 7) {real, imag} */,
  {32'hc0be6d33, 32'h40fd5d1f} /* (0, 4, 6) {real, imag} */,
  {32'h4021381e, 32'hc0e4bb03} /* (0, 4, 5) {real, imag} */,
  {32'h41367738, 32'hc01b29f8} /* (0, 4, 4) {real, imag} */,
  {32'hc0ab5f44, 32'h408da032} /* (0, 4, 3) {real, imag} */,
  {32'h4180ec4d, 32'hbed93dd8} /* (0, 4, 2) {real, imag} */,
  {32'h40274864, 32'h40c7bd15} /* (0, 4, 1) {real, imag} */,
  {32'hc1349101, 32'hc0aaa0c3} /* (0, 4, 0) {real, imag} */,
  {32'h3f2037ef, 32'hc17210ea} /* (0, 3, 31) {real, imag} */,
  {32'h4093cf3b, 32'hc00bce0e} /* (0, 3, 30) {real, imag} */,
  {32'hc0d124dd, 32'h40d0f0ec} /* (0, 3, 29) {real, imag} */,
  {32'h3f2d5c7e, 32'h404a6c80} /* (0, 3, 28) {real, imag} */,
  {32'h3fc6fc69, 32'hc0d88869} /* (0, 3, 27) {real, imag} */,
  {32'hc0a8e599, 32'h40201276} /* (0, 3, 26) {real, imag} */,
  {32'hc0f00ed0, 32'h409acc3f} /* (0, 3, 25) {real, imag} */,
  {32'h3fab2fad, 32'hbfd35c0c} /* (0, 3, 24) {real, imag} */,
  {32'hbff85d0c, 32'hc07380eb} /* (0, 3, 23) {real, imag} */,
  {32'hbec554c6, 32'h3ec3e2cb} /* (0, 3, 22) {real, imag} */,
  {32'hc03cf7f0, 32'hbf0a6aa1} /* (0, 3, 21) {real, imag} */,
  {32'hbd26a81f, 32'h3f99fb7c} /* (0, 3, 20) {real, imag} */,
  {32'h3f8a01cd, 32'h3f9789de} /* (0, 3, 19) {real, imag} */,
  {32'hbe04cbf9, 32'hc01117a1} /* (0, 3, 18) {real, imag} */,
  {32'h3fe849ed, 32'hbe2c35f5} /* (0, 3, 17) {real, imag} */,
  {32'h3e8e3bc6, 32'hbfa3c5c5} /* (0, 3, 16) {real, imag} */,
  {32'h3ecde21b, 32'hbeb38a09} /* (0, 3, 15) {real, imag} */,
  {32'h3fec7d9d, 32'h4004c096} /* (0, 3, 14) {real, imag} */,
  {32'hbec62251, 32'hbf3acd5e} /* (0, 3, 13) {real, imag} */,
  {32'h40676594, 32'hc08215a3} /* (0, 3, 12) {real, imag} */,
  {32'h3e5b8bf5, 32'hc016bc03} /* (0, 3, 11) {real, imag} */,
  {32'hbe016f07, 32'h3fd5821a} /* (0, 3, 10) {real, imag} */,
  {32'hbe89a660, 32'hc00308a9} /* (0, 3, 9) {real, imag} */,
  {32'hc0835cf6, 32'h4014c529} /* (0, 3, 8) {real, imag} */,
  {32'hbf3374ff, 32'hc0802a5a} /* (0, 3, 7) {real, imag} */,
  {32'hc09869e4, 32'hbf2fd050} /* (0, 3, 6) {real, imag} */,
  {32'hc1094b83, 32'h40e72d4c} /* (0, 3, 5) {real, imag} */,
  {32'h408e1dab, 32'h4109525c} /* (0, 3, 4) {real, imag} */,
  {32'h3f2e21c0, 32'hc0d6951a} /* (0, 3, 3) {real, imag} */,
  {32'h4034ff38, 32'h41a94125} /* (0, 3, 2) {real, imag} */,
  {32'h3f99f6f1, 32'h4141bda1} /* (0, 3, 1) {real, imag} */,
  {32'h41c41208, 32'h41095396} /* (0, 3, 0) {real, imag} */,
  {32'hc0ad06dc, 32'hbe417e0b} /* (0, 2, 31) {real, imag} */,
  {32'h415baadd, 32'hc183e558} /* (0, 2, 30) {real, imag} */,
  {32'h417cd738, 32'h413698b5} /* (0, 2, 29) {real, imag} */,
  {32'h40508a90, 32'h40b5dca2} /* (0, 2, 28) {real, imag} */,
  {32'h3ff1d8e1, 32'hc086a9e2} /* (0, 2, 27) {real, imag} */,
  {32'h400914be, 32'h4089e71d} /* (0, 2, 26) {real, imag} */,
  {32'h403ae9ef, 32'h3e308a76} /* (0, 2, 25) {real, imag} */,
  {32'h400ba9a9, 32'h40ba1e35} /* (0, 2, 24) {real, imag} */,
  {32'hc0649519, 32'h3efe7e3b} /* (0, 2, 23) {real, imag} */,
  {32'hbfbca171, 32'hbf6c98dd} /* (0, 2, 22) {real, imag} */,
  {32'h3fb36295, 32'h3f4fa318} /* (0, 2, 21) {real, imag} */,
  {32'h400c1d80, 32'hbfc36d79} /* (0, 2, 20) {real, imag} */,
  {32'hc05ac888, 32'h3faf0628} /* (0, 2, 19) {real, imag} */,
  {32'h3e5404d0, 32'hbfd43f95} /* (0, 2, 18) {real, imag} */,
  {32'h3f14efa5, 32'hbfdf9b70} /* (0, 2, 17) {real, imag} */,
  {32'h3e9c3dd5, 32'hbdda7130} /* (0, 2, 16) {real, imag} */,
  {32'h3e903620, 32'hbecdcb53} /* (0, 2, 15) {real, imag} */,
  {32'h3f988b6e, 32'hbf85249c} /* (0, 2, 14) {real, imag} */,
  {32'hbfd55052, 32'hbf194618} /* (0, 2, 13) {real, imag} */,
  {32'h3f1054dd, 32'h3f67eb75} /* (0, 2, 12) {real, imag} */,
  {32'hbee27faf, 32'h3e5a3195} /* (0, 2, 11) {real, imag} */,
  {32'hbcf02d69, 32'h4009faf2} /* (0, 2, 10) {real, imag} */,
  {32'h40348a5f, 32'h409adb9c} /* (0, 2, 9) {real, imag} */,
  {32'hbfc8ebef, 32'hc025d3aa} /* (0, 2, 8) {real, imag} */,
  {32'h402736e8, 32'hc08d88c5} /* (0, 2, 7) {real, imag} */,
  {32'h408a892a, 32'h411189ab} /* (0, 2, 6) {real, imag} */,
  {32'hc11a353a, 32'hc0cb3c23} /* (0, 2, 5) {real, imag} */,
  {32'h410b9216, 32'hc16a84f5} /* (0, 2, 4) {real, imag} */,
  {32'hbffaf8f0, 32'hc0d78ddf} /* (0, 2, 3) {real, imag} */,
  {32'h409bf46b, 32'h4117ac3b} /* (0, 2, 2) {real, imag} */,
  {32'h3f780f3f, 32'h41de58d0} /* (0, 2, 1) {real, imag} */,
  {32'hc181149b, 32'hc0ba5814} /* (0, 2, 0) {real, imag} */,
  {32'h416ccc3d, 32'hc18231f0} /* (0, 1, 31) {real, imag} */,
  {32'h40536963, 32'h41de1c21} /* (0, 1, 30) {real, imag} */,
  {32'h411d4350, 32'hc0f80886} /* (0, 1, 29) {real, imag} */,
  {32'hc11d6710, 32'hc08aafcf} /* (0, 1, 28) {real, imag} */,
  {32'h4146551a, 32'h3fb9149b} /* (0, 1, 27) {real, imag} */,
  {32'h40eb03e5, 32'hc0b8ee8b} /* (0, 1, 26) {real, imag} */,
  {32'hc09545cf, 32'h3e0d2728} /* (0, 1, 25) {real, imag} */,
  {32'hbfcf8fbb, 32'hc0519c4b} /* (0, 1, 24) {real, imag} */,
  {32'hbc5394ad, 32'hc06aa4f6} /* (0, 1, 23) {real, imag} */,
  {32'h4076bb1e, 32'h3c18b4b6} /* (0, 1, 22) {real, imag} */,
  {32'hbed485b5, 32'h4019ed58} /* (0, 1, 21) {real, imag} */,
  {32'h3f9ef6ad, 32'h404da3b2} /* (0, 1, 20) {real, imag} */,
  {32'h3fa4d3f9, 32'hc0089e38} /* (0, 1, 19) {real, imag} */,
  {32'hbe7e0fd8, 32'h3ffc46e8} /* (0, 1, 18) {real, imag} */,
  {32'h3f92ab7d, 32'h3f561cd7} /* (0, 1, 17) {real, imag} */,
  {32'hbec6804d, 32'hbfa99050} /* (0, 1, 16) {real, imag} */,
  {32'h3e0e6ee2, 32'h401a93ea} /* (0, 1, 15) {real, imag} */,
  {32'hbf74ca53, 32'h3e330d28} /* (0, 1, 14) {real, imag} */,
  {32'h40110526, 32'hbfc5db6c} /* (0, 1, 13) {real, imag} */,
  {32'h40477e0c, 32'hc02e3b03} /* (0, 1, 12) {real, imag} */,
  {32'hbf6c8f54, 32'h402e4445} /* (0, 1, 11) {real, imag} */,
  {32'hc085851e, 32'hbfe73478} /* (0, 1, 10) {real, imag} */,
  {32'hbfa35ee5, 32'h401853ed} /* (0, 1, 9) {real, imag} */,
  {32'h4036e20e, 32'hbc0fbf62} /* (0, 1, 8) {real, imag} */,
  {32'h3ea2be01, 32'hbf1469fb} /* (0, 1, 7) {real, imag} */,
  {32'hc08ea0b3, 32'hc0dbd6e2} /* (0, 1, 6) {real, imag} */,
  {32'hc051e10c, 32'h41185483} /* (0, 1, 5) {real, imag} */,
  {32'hc01f6fcb, 32'hc151fd65} /* (0, 1, 4) {real, imag} */,
  {32'hbfb5a27e, 32'hc0c8f4d8} /* (0, 1, 3) {real, imag} */,
  {32'hc1e94968, 32'hc17f7ea1} /* (0, 1, 2) {real, imag} */,
  {32'hbf1c2969, 32'hc1e3fcc8} /* (0, 1, 1) {real, imag} */,
  {32'h42236899, 32'hc1aebe41} /* (0, 1, 0) {real, imag} */,
  {32'hc2a50613, 32'h41cb788f} /* (0, 0, 31) {real, imag} */,
  {32'hc122dca1, 32'h421cb3b1} /* (0, 0, 30) {real, imag} */,
  {32'h411a45e2, 32'hc1306e5f} /* (0, 0, 29) {real, imag} */,
  {32'h3eb6698c, 32'hc1b03b8e} /* (0, 0, 28) {real, imag} */,
  {32'h3fbb167b, 32'h40afa535} /* (0, 0, 27) {real, imag} */,
  {32'h40af4759, 32'hc0392aa8} /* (0, 0, 26) {real, imag} */,
  {32'h402e8f82, 32'hc0b8469f} /* (0, 0, 25) {real, imag} */,
  {32'h40330a06, 32'hbf84a823} /* (0, 0, 24) {real, imag} */,
  {32'h3f7b6fdd, 32'h3ffff6be} /* (0, 0, 23) {real, imag} */,
  {32'hc02da1db, 32'h3c6d5b8d} /* (0, 0, 22) {real, imag} */,
  {32'hc00ef2d8, 32'h3f8226e3} /* (0, 0, 21) {real, imag} */,
  {32'hbf9289d5, 32'hc01216f1} /* (0, 0, 20) {real, imag} */,
  {32'h3f815be9, 32'hc00c5699} /* (0, 0, 19) {real, imag} */,
  {32'h3f8a941c, 32'h3f435b19} /* (0, 0, 18) {real, imag} */,
  {32'hbeea427d, 32'h3f5dd4b6} /* (0, 0, 17) {real, imag} */,
  {32'h3f57d8af, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'hbeea427d, 32'hbf5dd4b6} /* (0, 0, 15) {real, imag} */,
  {32'h3f8a941c, 32'hbf435b19} /* (0, 0, 14) {real, imag} */,
  {32'h3f815be9, 32'h400c5699} /* (0, 0, 13) {real, imag} */,
  {32'hbf9289d5, 32'h401216f1} /* (0, 0, 12) {real, imag} */,
  {32'hc00ef2d8, 32'hbf8226e3} /* (0, 0, 11) {real, imag} */,
  {32'hc02da1db, 32'hbc6d5b8d} /* (0, 0, 10) {real, imag} */,
  {32'h3f7b6fdd, 32'hbffff6be} /* (0, 0, 9) {real, imag} */,
  {32'h40330a06, 32'h3f84a823} /* (0, 0, 8) {real, imag} */,
  {32'h402e8f82, 32'h40b8469f} /* (0, 0, 7) {real, imag} */,
  {32'h40af4759, 32'h40392aa8} /* (0, 0, 6) {real, imag} */,
  {32'h3fbb167b, 32'hc0afa535} /* (0, 0, 5) {real, imag} */,
  {32'h3eb6698c, 32'h41b03b8e} /* (0, 0, 4) {real, imag} */,
  {32'h411a45e2, 32'h41306e5f} /* (0, 0, 3) {real, imag} */,
  {32'hc122dca1, 32'hc21cb3b1} /* (0, 0, 2) {real, imag} */,
  {32'hc2a50613, 32'hc1cb788f} /* (0, 0, 1) {real, imag} */,
  {32'hb7000000, 32'h00000000} /* (0, 0, 0) {real, imag} */};
