-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
oVT6hW1mr5hLYTkx6Zg2p40Q21+rkDwbT/DMboiHZDuH3UzV8x77a1116AHe/Xdl
W7i3Cbi9uiLM/tV4Iaeb++FaQSglDGSvJjgANEnETvuK6AbegsDgoxohO00ptoQY
BEnz9qunSSfwbB4z4nXfiAyvq7T7T3vGbShuB3MQ8C0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 21408)
`protect data_block
RrCgM1NH8pjC770M36H+gyX7IV4NbM+9oFUXMhx45aKowv6ch8FZGvmE1iB23nl+
uTK0wCImjdFsxqOyN/+RC44QXBk/rm7E0Sw9YQH3/qa2XpgNuOVH7hsDG4jbpREl
/AndJnH/8hJbdohD46DTnlWkBfd7Y3hr3WJ662MUTemz4JwYqi2FwUrUJhCofk48
65YJ7Wxl5aA6G4+fIekhAe2qLuHq6TkCBlOpSai4jinJUHHNnJLcZQdMHj1wk5Vs
0Yw8G3eP+S2MY3iF/XnlFPLnbTFrX/s1k7CrplFmEcio+opPrxQmLrVVFOS3pD7l
+yhuy8KgAwTxSwQRKFWrWPgfFEgMzXOTx6jVh+4eC7PGV94qoUSd9kybqHPgZWER
dD1nkYvjGdiyGb5RASc+DRmPLtE8kK8WEqjmpznCJKKy8cEZFerbJYytzissf6cc
sTkoaJjg4o5R7+28Od5RadIVbKD9SrV3Zgac7CYqV2LBYkq+Yi/eBr0FtWjoys4K
NbrjpBrJWkdoqUpK2xSLWBV8QfY4VDT5BrA+Zg8Uj9MlwaiEccWC+9cUgA3MyPX2
W+AEe/ReK7pmcro28l+YPTmmeRIvaxTpEXPM90mnLKCh6qYgcV7dyzIsF+yS8IcA
HKqBLmYaSlN/FwcGBE6vW1qg/1dZMvKawZZvdVauHa8vwUOk01sCHlS0I2d4BSim
VfmMxRH/IfAVZ8HviEZkZEZane7llXVYR7dy28zjnFWDqrRvOx4y7AmP0ZSO/sox
vXb71ooaX3Yub4LivYv/X4YvCRTX0qWUcVrrGJatCmpxYdnrs0+6SGRXKdPdcWNN
9kosC8jdB9xpQHBUmWcFpY1op7Pn4Yvk4gDeKQ3JF5hh+dU9+umzezLiZr55wPFe
+5tABe2jLKcqHzRap2bnfjGTSBhDQLphSMwKBn7w51o9eBlGWTzNnQB4eBP1irw5
lJ49n/ZDWW9fG4K7PdjHisa5BXxM2K0XI3HPm9IMUSHm7KPql3kixg+MMlasS4WE
8B/XrAof4NAI0lySlFVZ+WwsW2fBZ/Bh/7sQj4XNnNn8lWOD+jhk3D9pD2cAH25H
slA9j44djUHEsS09M3hWwF+M9r5XMRled+eanRHOWrerl333WzRKSgwPjywchHRY
34rOFMvzEjl/46GbVv1LyLfMLNqo3dy9D0tqn44/s04xgMhTUTIiZiRqR2tYZBMn
ruTCNOXJ8tx9y+8ND5ggEY00LgkmKRSodxXnLI7QQqVSiztpRy7PKH59RGMTjX8+
X3kMsaHqp0RRyMm9KE3OxDtBQGgOBeengIrzlotE6sp21vtnKw4Vna9s9APxj+yo
8rLAkdaHq/1jlHPXFL8Gjfz9D0r9+xSvTFrPyS9iNTZxTZZt7HZEhNGRle6YMI++
W7pJpdn/93BEiNoa0EIPCvf2+L00BNT2OusqgOk41I6VAE4X8d1E9dQJh24ZkBk1
AaNnEgOHU5WfeJukeLk/vKLnSsS5XSkbPFGinapMdMTuPLyS1AmGg3gyeMgcUdO8
OiimK3Z4GgXOj1DNgUQ6OckMfEVNg2Q4TSZ1aynCdCp1fv2p4WbzAq/S5CjHZ2qQ
DMp2cnFtZEnEDnqhdJ7qbxfMXKAQs1x+6Vi6RfKEIZl/P0HrFDXiAhwzU426q/nA
3JBVJj58IemQWoHdplHFlg6tWCLpeAhK/BmQCCNSs1IWtaOQcW/FGTQebMkD87Hx
KjZcW9RL43iQ87Ftk5jGfpU3+TerTXuH4Tfk/IFBBMtPXlGM8P5ZXJdWBzpjibMq
8lN/0r+FDKoifE9hd6ELAg7IxSsK/PNHkR9xnvbMxcREQeMirKDUXW92tlBCetY1
cIm8gqfC+Ct6VWY0qtV2LtBBNbhCwfcN+xxNCQJzKzAyfsjKEF/OSKsasCW9OO6i
QMhi80cnaAn1EoteLK8Mjig4qjh+g5rp/AgLWDNnQe+a7K+ARUwsSlvSSx6Qv9qj
acwygpvLTHPMbqtFsfXgMWfa24nD3RJfZYPds6plsNOWyTmb0Ut+v1CnX8k3jQ0t
ag7o0MnMz5sazsDB1fF0YwFOx8ITVpO89Sv3lIvTS1kS3vddgQktibxjZOXmqzgy
pFUGfa79suDK3Y5wNXCpB24OT2glLCYjQrthbnx4f8Xo74J6Mr9ZfWYSynJgLTeA
7GN6X04w8Vvlm7+g/8CRNKjC9Zs76CrJf3MvLUvz3TefVEcW0qTBTqQLDuog7vA0
fyGsrxtSLTzOUCAOmX/J9JAXYG8zW7VZuWzHOxY39d5FtO8sUiz9IZNLE2NzA4da
H6b4jeFY5GVcIUiy7eAWx4b8g1yBB5tvKHU4Um0ddCoj6UstEDsxF26KlPLaVVXq
njoimRbPpJtpqAorxYjf3nw0Iku7iRc9vq14V3nt0Cy5pUS7eZZi3uJJ7pz7GFB7
uALqIEXP1HuTphs9uBA1gevelWs2835d09r15F2vVH428iBAtXUGEuhLE6rs/MP4
ug1tenonDrEHXQxi1X9e3crA6AUH/sy1IeO7WHzSWbLZQkmYCEKDwX3xhw+jVzLW
c4t+qJ59eRjIb3Pwotbgp4PcNjWx3n+cjy118XA/motmivy1GeavCad8JuRg0PSr
ZtK/Mnp20F9DSGiKQcZEe9E96SNOI76fJ/mgOTZORQ7qWVQ9jG4cRGtKx0FrRccy
qEmpS6B0LIcGvHFZ/rtORlxWFWAFbNattnlMAkHSQcydN9ss1uYrqGKDFpPMJq+f
odYvAb8UQpx1b1mdl/7lw/8HndmIOo9Fp5JQikBWh32pJZsoVyN12BvaaeNkNUov
pQeVEn5LEoZyUKTZrxT+PX/Z58t5gfFssfSGCh4PWMf+7dyhOdkN28m4QZQgSWw4
2CYNz90eQMN7nGxpgW+mlAeMTnQoQhncyEIeuMpCaqlSkrcUfKKRlmCA7O/nQo+d
FhtW5jpUVDyD1waMQXmV+Armzb5lPW4p1996kj27FHUn+2W/FuaS0p3y0ko8HVEK
QPLUMk8wutNkAf1HAz3U1S9O9rkrB4MF1yPZRol8U8gSrZsS6dAe4mcmba9KwlTu
mEAj+7H8SfbqWHRCRnlMFUhPX5tIN4YZX11Eqgogd7ToP0bHaYPDCHXGsPKDoh/o
l/Vqoyg4oZiEE5vatgxD1nx9JXzR6g+oy6xYtcicjVqDDEyTvP1imszEiBVkjr/f
+f8VqA2artoutThivWJ85X3a72lDG1okp10bmAnYZtOWbyHat5up2vg9lCL0lITk
5Nu1ITD8WjBXgNXl/pkqOV2t+Z1rIrNlJOvC1cfBrTKRgKoLxbv41CAQ6G2SGEiW
bh9B9fQI0lXpBgHFuYBJ4iNISa/t/WIHwxpXK/TT/is8T823InERZwZV+8E9aD9m
E8M/Blom9Z4OuOD46nW3hfy9Sc2+whGzcymJ7xpVUzX9n4Q492+sGUUaLSOc+3mS
eZCp79Aj1HZbV0jvFk22KGgN8V4NW4+AiUQiRBSdY/OrtQ91MHXmRXLu13GIVxmQ
74PecK6dBbSleqb0Q8xKHiuORcg2nz5DE6S+H5UH+7rcuI8pRsXSdgttV0AkDfE4
iNgoaH6xzPia0RSSkYmLrVb7vww7LmKlK4lDv3E7ynSCkG/9RBHbfPyZ6mWouD3V
1v2Rwqx0Jht3LHXLPlUNO8LdyWnIyqf17PUghm6lC3Kw+6WhabPYQnX+dY7IqTpa
VJCiSnXe01f63rt2iawkBSbKA/JL+98vJbvWQUKw51afaAjMwgEQZwUSeKbJ/F/w
fjuDC28Dx4JLqsj3LbHbCtgA+BcsZInmU5ywkWMxlCsIQqoSHgt2OMyBY26uXqNP
UZCRQkdAPPD+jHcE5wgnF8fjbnnjqVmmwYAkcH9jsl9/sfqhDVazKfjLMO05DCQj
1X0ki90BwsLOO5PuicrSB9ccDd+EQhHorX1Va0l6DKExARUzeS70q5/eUoKLyflh
VSkC0DAO00DV9DvVgiDB20gpTeaNcISk1J4HH+uvk7EJGRhiri17nWGS9ceLCIhd
JT/PAVA6brbSrznZoLxzTR+tfyPhNmR7GpfbSeovyU2c7BfE6OJMAzwZgx6WwovF
x2qr4g05H5cbqJXLbmhZ2nHUkdpN1TUvtcVqhSeoQeGwAW1WDIs4+Z9OqoqlX+vq
Wi27o8LDU8ZDseFiJp2AAKQUiqJv04JisB+4ftMZKYxKrlW5vK/GFmC+H+N6pUiM
h6R4YqPpC9sDgTJ3L8TYTN0iP+HBVjQ8KDfbiRUJw+t71FZJwxp5Kh7Exa009lU9
13OASeQ5Qk+QvcyRsCQOesmHNRvlaSJsFGxylaRtSMdQy+woS1+uJlfvcY0RVG1+
HNuhiwjAv+qyblH5LEnUxIRNFS5EkfLzzGhXczFIIj1iBsE5Pyq2zOjV7cJd5n+d
xVOKpb8Xk91+lHS7SZSjzHyBCFXqDfxz1bNW0ytiLQp/94msb93YNCk4h1jWQ02Y
wOEKZOWdMfilIKbPSPLUgNB4lXerhIUh0Ct5Sk4v3kEXiUQMZJuuGPPlRFG4B7Y7
hq93FPpg7K5EpUkoRmm8X5r7XljqMbk9lZ8jmYb2P3iaYp1vEEf/kGYNTNg7rBxe
AVjVfObJ4q65eiKtRBEcsDrLFQ9W5OFtDPqKUmbPTtb16/+zyv+p6k4kx4sGrWby
1vczTlsTOt9UYYkwPfEBu/r82kAbKrmDrpTlsygLtMxS5z//XT0c1rBVVel2MwD7
DldRHXPOsLmjV6WGb7JKAS/pD2Cv4ftcdvIhwhdI3+8Kc9REDK7XaoV7zXZL63Oi
2MF4mT62Ciw2GiUH1ujqUGWPwQCvd5WcXCYIvHs+B1SYj70cY+WKZNJn5QOQqMqQ
bqzGZ8ZyIhR/Tirw7/oJrDASPvSng0waFzMBGML9NfcXHtl1ITwEbGRHoyoD8wZy
HAEub3hHLOPchfr10XtxkkI2nkMtsAIyq2FJp5I0FpACRli0GdaMVJ89e0brDfV1
1ju+nBykrxWb1O/yh+NHyEhXJNNs6BWZRlpxbMGRwjJ+7tEqTj6qbiA2DdypcteR
HHuBgdHHoU6+Xfa/6YrpcW8JVSS+0M6wamPxKjeoabTE1BUzYsCC2MEapOz42xSy
ci90hpCbSMzmjMl3wkMgdNoVJ1mb14PHhPeOXGpd1xkQ5rNJDA+jrSI1cA13bR76
5HxWHzOjRlP1FXce3Y4q9AyGz9odXWX1+D+wsly1CLo6+CGH6S2eN5y8p9qBAJYw
tH3MuUWY8SEktMzsiXiVq9wO0VCGLgs8FPk9WYtzx7fBJUFcTQdUz2LkvQJn9+/7
DGKJwiw/RT7Bl8TpVXiR4cH1wU5KYlFJClFeXb7OIRuI9yuv3CQEvusJamAh+IkC
dmcpv7cVSigHDWNo9BXIFTklljVEYdnSAHQYnWKsTpCRxdvsH9hvpndD+5XNrurW
CRUSIIM8ZPFdnU9m/zxIhx9kr7IoHgATviGG5Vq5Ux8y4ZMw5sFAGsdeLwqyrD0e
PcxDkmBiLtaRKmekXG0uZlMryYf3YbqiazYRYJbyiUXPUBWPucgyuNBXJH1iz6VP
h+e38tAUql2C22Up5ToK1wkDKSnt46Ho/fo1vDDacPtY34HJGn1742ZL9SA4pGYP
762gMd2CkcDTG8jqJRw1IJoGejwcU8FLBg/5AEMFc+rOUerst+gTf001h8Fq//gf
WMYUnZRJcbGUItE7LLHrm2csyn+LZm3cD9YEYrtyjJEU/Zle975NMVXSgsvdJTkm
5uFy34jXGwyp/aZSNLK5W5CK8Sz3VeQJZCJFcvdTPGZVgQuCJLDIZFL8i0cjl8E4
mqde+WHSe+HBkdSxF9d4wDOmUFBuKTMiAbmv8t4CkvKXuRbnpSEhoZmw/2I3DB62
U0mIqmHgok2T5Q8uuwDromRvljJ0NgJzKYB1vEwfGo0f5u+42S3GUm2WhnRbkaYk
IEMy1ww1cXYLnIB7VvuY+aU+Z4vDPTGI6sHFAVyk13ychcIEkMGBvs9J2EMs+1Zb
I/cTn/3el8kIr+w9q5KnMziyv4r6OL3AI6isXKNO1fq6kvfz5182hH0iA2Hq7CeZ
anX0ZPE4zg2wTZ+JFOINTbdEOv/kGurajiwc8AzKvSe7UBIV/VNmsaK9SknG0uVM
SldbSvb+r1TYatZRQ++7cWcbcAFFPBkyXkQNDWLPO8tKjcWNTEGKpuJqunL5rgbu
8ev0hZU1gRf4+/ZECtzeEBns4LIr+O5xpBafw+j1+1GTgoTc9gU7hdfrjsvWD96R
y8ZrMMrV7jueGNL+RBWBhr7ZCSdzNjs5WtYaJ+VMalQriw5cOFYHzRhVm9dnmLDZ
4cBvBxAs7X2m2pDldFUpaWBYyDMePXbk4CwnLH/61p2pTtMrRWHzsBB55YU03bJ6
5bIFn8YnYQS5YkDVMz7RNKzKYTodwcu7xYd9yhKaOWpeZhDvNuj/7YrN5e1th9FJ
RBUpHYCqx6jYXKGlsbjYHX6c/lh8efqrdZs+6BmtVSOuW6x4tLVOJydX2ioy8cP7
bkiiRNnKewGpQkrdWoyRayvQal+oBhIT3rWO+4DB+BfwY4fVW4YZutQ+zxotosf2
kv77TLKRN3hKs+/exA63HXaUWtxXgouxbfrB3SaBDYp7PcdEaVM5i1D0EfB3XwLP
Dx7YjQutfz84bMHz0jEd9rvM++O85L8qeKzpi0CgrP03CLr8V/gKnzSCVjotGJYI
qNQD/x2WaHpUu4TB97Gekla4Sxrht9B7PDWr+HJMtVXmaOrNUDq/g9h4y7FQ79Z6
8GhS6QEUJi0Y9f0e3Tf+oJo2uvxGyYmIPVB6+NvtNaYraa084o+rdwvSvsZzKffS
aX4Cyfq2FcF+wX4CFX7VFwrug5RTvRV43uEuUEltpE3IyiKKEgQ86Yf5DdO2lhPi
dW3oXxefWpQuO5eidTibIy/sPccVkEpg7XXRzSPM7d+6mu4yYRx4B6uY7QMxEqtL
iy3tDIZb9I7HBOhbMPLR0KoOB4Etf5o+CB8FAGO+Ghqa13U+TJ1nOV/0o68Cbg/s
BRTKZwhcBA74/PnxllGAWtXYUiE+oBp76cSm+pC3OllIbgmYxbfEqncUsBK9wIsj
OOpY1oHG+g4GHnLwZIphoN1SyI3ROtKGKQTMIn3lGI0Bfd6S70ql/y6r+biLfuiG
NiZLV9smBObWD1CyW6VCUUmrMg6sAoqbLQoVcmYVkNu2lTJS85uo8sU7J/X7Z3+H
XIghtCc0HG6g+vedAfxHOcm+B/yLcuhDg/zv9KbIAeVc7oyKVo0+WRoDZg+YRr3L
a4N7nf8YX2FLfmiTekDGPVCgGHmTt7hwx66oNeRPMTHOyUiu0zF8f3xjhYjm1WA8
bmb0Wrm2FRA7z71JwJ/pS5D7OtmfL3WpL/ceUzKgPAd30y3SVwHUHbgMQgCkMHFQ
b4wva16xCcoSMJIFyIelAsEQ8qHqhVXuASlIBEUsqoflhDu0bE3D2+3Gy3dks/8d
f0OT8grXxdmdNj/PJh6ywO9F47JWJhAd/HuengqY3ia6U81FRj0uRLk8EkIztSvP
kHFU6zwKGZ4KJ77yTvks4HLoYTfMtKQYSgnPEWPzTpzS13qAk/F2AhQFjv9wBT5u
yDSRXyNEzBzkzfKszhUwLB/1Cj8R89HtGgBBG+Ke/mZIu/eE44ODIbXptOLj7/FF
1nz4zUtHMiKuCrsAy6g7XhMcwR0ThpIokZmfuxVse5VRcj9UIU+QbgApYiRmL9w9
CyfM3QfmhhS8zjnGHSgm2d+a2ETwqhq5vacB94PyniA9VWLfzl4vvYF//cTkBrYt
zW6JhniCLx7oidPjVDpSBHH+//rQhjOWXWvdyZ2THsXisgDiRoyTTMZgxVF457mB
9lTj0NPkVn6hHYWiKuGDxNbQR8psv/uiXBO8axmgbu0MQJyP61jy5E70IIB/hYRI
dNQ+B8uBHE5jZm90BVCvYuOw4EMdmIPJeW6ZlD6+YNBdR/WdfG4b0R1v/8jwOshP
Ym6svO1CWyfRnlgrKF5PEZU85lL7sKGh9cA4xx+FB+/hikAyc73EymQl7EPU+jVB
ifQBnm1Qp00tIX+vnC3apzuivy72xyUHIvYg42Co5GnMIlnbYn1b1X23xhYgWrO3
7DJAqqKwZY4dL/zr5FtlDs9Sp8CMf3LVBgwMqfEBwrvTCUAwfgnK79vsvAiGr+PZ
EfYoE2tblWgf0yq8S9sjFvxsB6mC3g4MRTDW8vyHKfNVitHIpgONtl3r+PU1z2b4
ykRT7X780fhkaXgmvDi/YwCUVXs4gwN0StL5tNw4n8fYDi2ZBc+kvD570pTq8U2P
GrvdQalX7+rkB0t/Dmr4ELHo9QCqcWttCqztSMzZGtANWElHZ0UFbPADZ7IcLj1g
Vv34FHr7gkPbdjYwMmSLROE9alWUZTet3YIFpj20cB5gEv7lzzPBJrrCg8IbLdBE
mPiE73oB6oJrny4duwMqqu2LS9Iaa2d6tIxcOX7t849N/qC0lXJsuwbAfCnUgT5B
8LxLlf+NUTF16DNAnF2wERflc1IT+IvRmJ3GfOon9318U4fANjyW0gap3EhzBGRj
fBcrtCFqwEyVs8qSBAVOgr4XUz2ofeGNQ/ckK2LtYo/eTt0yRGsUi2HepxJsYLGL
A9aP6p2uF4HKU/hjr/qhrfNKK2LEUZPIGLC/xNZ/oh1sHJ++Jab18fB+8/xH/PJF
nmS1FPlCAewNS3LpNwCR5H07FXprsoc1C6V3aZdTHUu3g2z2UzmEXm8vWVA1bM8Z
D1Ax0ypkPgO+jsBoouG2/eWFULHhbDeLDC/PMPzFbEqQ2xwPUMlfMFJtH9f5vAUt
ySzz3RtyH+UNway55qDHobqU3pkWcGRk3HwWhJXqNYgfFoCCRAAmKOmKCQ/dq8kh
rwr0ZAr1Uq4xr+9icliOWMgf0+VSPujzgdQ9zwWFv1NwJqQmeIkZDpxCq8AhV/XG
UVIVVUnBxMtnyjrqNSV+KvK0HIJvftZNKZY9nK3gs/rnh2jVvH7AePewGURV6gEQ
4NjtYawqemh1ZrRna+vkU8Vy8lMSOO8ktcuu3HRVz9nxxeIJqP2jkWT3OEUIH40d
xcQal3X68o9FVvjWN1cS1SJrdzRja4hiHg3uxftX+mZQo1jXRwI5VkBeb8IFeBjP
uXjtGSRUYxCaBBRjA89eLyUlR13YVSZ/qVzVOGilkJMF16ERWMeVpsqrfLpqxp1A
jtDmWGDOrF2XfUzUbfmWMk3PmVo+CdmTVWmM/k4bK8FEPa6ocKfe0Vt0Af2jdN3S
DnKqXVTelkHTcvpnTfQwGC6kEunLn2GJeuuKEHM2EDYXN0HX4ych8BK8KQcHhw7Q
LrdwygzvB1zps+DLbGZXPA8C2pcX2yYX/Yl5UWdexLznCfFhPwWexuuj0ISKx4ik
dNZN+bPIS6RY4D5ASFcJR6RYIwNbc6quEpqikzGLHi3sY9KCcCTwrR/O7qZ09oqY
UAJtq0aj5iVADrTI0QfGclFvEofqrBbgA8Vuq3KtnWZwxtYLbTnnzRHIom7Ry+M6
/VHsKbq3Zs4DVdXm9mkTWf2/1muEelw28u4TTEStTFaw+i98w2AUvZRsG+6kBSwq
0iGElSEq8bMPTDw46PSK8xVNCMuXbzgjmvf5NOaXL5T3/s49tVDT5kERJ7bw9i+b
NFntzRMtvE3qZZOeaIxdoNqCo8mCluZaRHPffDbzamc6B/b6aELeqoBSHT6Urnlo
dXrhWudgMNzvFew9vFKItt3qZGk0N+PLYCAqdaXNhwIKXweZjIBnRSe3YzTymTsW
4q8o2XP8uTNjP/V9Ppg5xDlWsdRaSCE6SJNSUzticqyyn8LQaV7CQQ8PquXhbAqs
48QFhqlJ/gIqXIScFSQs0nqKmBQv8NzQjnbPWbNrtsxqExvhZ6ZWIowNzz8QyTJJ
QhJsW6liFRoV+uPO+QSxC85hC+hViCJ0MnWE8p5bBFlCzrVjIhahxQB5tv37uR+V
uvBpgm5DSfu1CBcb+jC3cvhox3v5sUrSIPrA8BWhr/IW05zy9OnDebDFHYn/QstN
dZZqVoxc3yf8P+SATgWIXCaztkovwpxajFdVnUoM79P3MC1h/scuKLmPX3MKyyJW
WRicN3EeiGlVH3UNMcC2HJDK0Svc0J4jfaYZHNnunYN3LhnUWVXtods8htMuwAhv
bXr2aB9DLnu4/VpScNup94pxsY6CEHqDXxgZ/RYwxb6IbxD6/ddyoJuJlsIdTzUz
GuxOS5tVjH/h2T1F1j1EZAha541BgHeZPItDORta8n1MKzly01yNPihNwoOrfau6
ieM7TAvdCqUjf1u9ErHPI6AzBzrD7rZAxNN/TEf9iY8hVBBjmT/9bDECKtbMoZju
CLhw8VzO65ljInNc5qkGdKAibjZrckT+Ht3mStEtGyucax0aaCu1ENfRDUS/lrvj
sWriPyQ7L0UvSZcex3jkq6qFJklA1/hTVd2OiHDTcQQ+72nlogrAjcurUa5Y5xZG
r4YnjT/IEU3VJOVGg2ia9wJ0crdbYvHYUrC/Hu9Fm2wzVlNhAwqZgOiX4krDj01r
XH7Wj4S5K7EyNU4LLuZ+orSof8Po6bfv+N7ED6bJ+gQojIbvvcHRFqcEgnsEwt3b
qTYRT3VU65tJbjYw0VySPVqDzzEN6JclUVanWB8DEBk5HSYrsYnWX8QwtzTusrZ7
1mWW2hKqNmo11Of4Hnlza61ba+DHOdB8HDQosQ3iIngeTGYA23Tu9aCnxkzeBBsx
WqCau/6xSw8KlZ34tCsBfcgZ03WBi/NM4weTt+n4041iTI9NNJQJzfUwO1ZLDByy
nKo2G7LiQSJ0eBVwTTwNyMq50cU9DfJpo18wuOYOsLEhNb9/sEZuBepKlCGyxXHg
ZCmKy3nimwlHaRITAUujtjrjWZK5yUrlNYUj7sAeoLf4f7CtFPRRe7CLgKT23yDz
nD1awtDpW1Fuk73W+CIyjpR+62nDOkV/yHh48D6ek0UsRlN3cf4HcpX6x/KZdJjZ
jbCJja70NhMVmVaiNAIzScA0Ct2/UumCdUaOVnhUo9E08sqVIf3hvknYUUhRYpeI
Exi8g09kAnTGZ3hPfKmPbAJ+fpBnHV4lqwElaD5yxjU6n0KSD6AQfMCWgoYfMyli
jGKhzI6GpMXUPWNyidN+xn9mYGT5xaOysj8aiNk2KnGfpFBNzjbk5yiWWA7UhvRU
puMbAcb+1tD8jC68TWUMdw6MW23fgiGFtBCtS8CCqc7PFGn9pfdHMDTEO5zyB/RP
4POqwJIE1uKKSNhvnTVN5jQtYoRIT6bmlg3HrCt87l8KfXOVVVBBUw0oGQ/j5GBc
bD47ZZ5mQ6VqlxFEQeKR387+MtqIiCka73j0tYY8iI3DjIpsZt7lSB4DiB3tZW+l
GIinKGQLDJZR64nkOdfiujajslf1w46JBJqrciHK3y8Q9n+7JwfKPK+DMWc0JIPg
/fRrhbCkWXop+kLZi9F0QlLc3dFCKUxEr8t2Q4/SXPvEV/O07EbHpdxjyAt4MhpK
gWwm1xCdLWwTFCJ1ii/4Cnyf1eT2WaJdqa9/jPisZNH4JGi0kzPmQJmTs5I7tzNZ
wcSaOFqfQuCNYNs05QgjjKavQaJl3jCUsXCDKpTK9fBq/s3eZv+sL/TT9PTKvtRX
YxQQL+1TW5E1Cw8fdjmXm4GcSW17wzEPJpBj1xcg3+1eWzA13fykrVMsnQvRv2cw
8FTok8rIQ0PoGi1z5uMTD2huaEqyHruQKGXegdbX80Z5C1S14XNYV3Z2bwHIWeZh
AgMulBUIfbXCsai8QlMxHcL8m/OcyzVuQwgPCrkfovX9T9ZKHDlgtuu+Zw1TK1mH
c7xm0iPc683W4CKvyF63R8IWagtGQqruMYvv/Q1hoTyxoeT6toNcSE4NjIhopHtu
EBYh5G+/Hm3w1IaIo9iKkPJbbEgSDQ0wTvtWHrJIZtYqx/YJjFmfh21g2avR30n1
9ejPSIBzeaMrFID1CjDeZlwzD8zDTnczKCDfvaDBEczhCrthULuKftmbPxXbkp1E
6risCAzlsyg4jWGwBgX20s+jJofzaHDiHMi6bKRHuT9AfSKxKhe8//t54xtPEOVq
UmYw2t5LGjKZKphCCp2XzIMXo1Z66sRj6hlIQm5QQMksdTDAlTzABt3mesnpGbdM
LpuQzXJcxFFpGecETKAXvNG85buxh1XZekcDBR4/weww36JITaxRNNEtmneOD2wM
wpTbodBLv63ihke6EctM2wsjCpewIRgVayV2tVaXF0hservAPDFPSoabUusJTO9r
0l4suh0LbSHjOGNnh/7Ujdvi1UMR70Rksp1R4Zhy1ZJYSJ2FowGWbcP2vnWhmEIh
X+Ww9Eiezz3sRZ0TCBqM7A1Bpv7QrMqnHigqon7R9uGcNM19UANrN+q31mnMLWEK
kCi90rTQ3osX/kbMC4X6StojuIDbEtltJL949OTmbZp1CNjPHfCvKNOHcZaHtTm3
+SO2tjs9FMPKG4WRrUXicBS9zdv9lkN8q05O2iLqcAcHhLixeYvNMFwI/GXWus/K
Xb1POgD9hoLKbrSLWlljB686CNymC1g1tOJNMG83wbawVoFC53kjSSyY0p23hORC
NEdFLkLlJ4RYxlxLhA5gA81XEmkmVtpRoA41A9Ajk2pFUqU+AfshHu1FgmP/m1s5
z+yhoKOl4xOSdriXL7ZnbIGgEmlWj/gWI2wwfQOmdUoIvKHAsWJVHICW5uwApI7o
O2ABHhWEzz1Qqokp2Mk/Be9IEt3zJEY7t6dE0OOt/V24ISUZnYx4auLvJRN7J729
zMYlpsr+l5iFzJ5CWzje1DPSgsgX6jxXskJ06f/9KRAnzLjFG+v1bOaq/lWJuLP+
q/nW3ragd6gba+5SNSrU51JvZJA+R/TSu4nnj6WhX1AqPK5X1/kH8CjQRP/cChPJ
UkDKGnV9NV+416c1Br7Kq/10K03qLr78rNklTks9J35tvM6x0BJhPzO3UZQImxWK
JGS9hwp7p7fwZ6KyYZzJ4NpzQGma5w7OehlTFk2b0CAy2NAcs8VQ2uy0BSVtc9ur
cxCCvSsU6oKM7vYOZ24MI93nqNp23ZSRMlOdwULgn934IDxaBDHTcFMkgYHO7Pw2
hC3QB8HFd8wlmdFMfVLrG9FgZWVVlhIReqwk6bS2IVazt0Ic0xLxdl14vF6grLky
Ixrov7foJw7TpRoxqS/qrg4ORz3HHzq/RsNpEyAoUXVYHCJrUxWwIzy6TvArDiqs
+aOiOFEO/ClM9nSro8TVIpS5zs5B4QASotOpl9I7W+EHYdq/oDLOsdcCRt3vYvCE
1SEjJOTyEcnOOeCDRL+tzBDa0NPLB70ACSbnkSdFwI4FR5SK9mSexlhLnfSLdN2i
7r4iThlxqJea/MYoajhQnhTad/QwN0Xtgk/SZ+iS811p6Ixk++F+xri81hF+dO5C
yg7wh2C9w7C2ji8VCRdQNRvQfCS4k9K3mt/1f5xCD05MzNNo4U2sw4Rl3dNaI6IX
XCV50LaaQrA/fGnxlyyIUsKWaqRFTdzY2SKIo/fIIJQhg5kIXZBILhq5bkFtkZ6y
/ZrtoWdxKxw4eFi1sM3jUmZHVIxa7lUmbmAdwXanZtb9Ar2U8D5qj4ExYyTt8dz5
q4gadqatAEE0aV1XAMIsrtoYk2ndpQQ0TKJewg/PG5LZGh+p96ZiDlOjrVnchE36
UYjy04hvV7KZg8qhF6JrwB3W0rerNxvXP2GSVhlxUrR175YXh6wln49wabRU1WtB
cWw3vtKm3vq3B5teHA1lfro+yBwxD7oGsHR4Sso3RwQuhui4bu90FNstirGUNz2H
RUlbkZGT/mNi9ZMK2kDyR6rfG+81YE3oSlkKWrNcznk4MnSlqK8fA8YNVJHoik0Q
Td1MWBGd2K5NQ44Pvu26JF5LAkm9AOiReRBrJlQ8LLkDJbtu2B2JsVoK+XWnemyW
mDcAiOV79XwaXJmVlfuChhpYu3bD//6kLtQ1GpSC0jyMBm5jk/o/g8KblqR1E0r9
rmBHCLK6l4rF/1AVPbRNU+nky1gbXaNCw73+oQLkfrh/G6DhYEmgA06B0wVfxeFn
KKnZ1bz7JLKpGZofjWBdUI/OAOnvmez6oZZCcaeABkBxkXfK7juv7J969/TvzC9j
XoNstDpDt8rePRAzP7CgAK+yCVNPmUf9fBHyeDo6elFl4QFATHEMiwbLXdcPLgGe
DLVsRza/1pQlq1qxUkDkVIZL00f0/MvdBsOsG+aMs4UP4UEg83ammG4vuEtc1fap
5gt8gAKGXJfLk6GNpAkjfYm4G7kAjnwo0zcQRibID7IJKQxBPpL9vExukZY2v5+a
1ygpbe4vCojWnO7osDxGb0E5l1g62yF93f4Wmjw2AKtlGaucqE5nUCinLIWNOszq
m72pXwsdxqo3VUZZUcHPpNVWfWtkz4qe20WRUBAktIDZLwiDepCwwd95K3PwYEST
9Jc4ptN5vqFMQrnpl/L3AgsseFyUSM2geaY5sfh04wFSlcGm3InwlI8AoxwQGnZM
1gOK5nlPOpDCKaJmOOFoH5+ZRwUCBiNNX25R5XJ6It7nem3bWriBHk185J5xs3tj
RoFGNUytsl+G2BzCw73TMI4/dwPwgzEsrFl/DDHvL+97Khkzb7l4Sx1WY592sjXW
2XdrW0RjRG6Ifjn+9ZhD3a8IypNNCl7KOxVuReMowLxca+2Y5KYOdPPCW9gNaQ2y
E/CMdwbWzL8nNbhcvqzS+fvTqLXUUMplpmzLK/pJUxBHWPcFUlDOrxsIxwsI0F49
R6ONuNlk2eWIiuh5mo/qVYMFVbZm8t9NZgM8gh/OXWdNDJ6o++s6/mse7p9SKpOS
37Zu/eyauUZNVbM/cBhWVH9VGFn/cHjk/k5P6AF4FVvMj6HBNHmTRdl0bNoTf5ys
fvuxBNP0gWJWYGuViO7hnAsIsRttTQm52bgHo7mqCPEfJgS4xIZiQec6OkPVHB/4
+AqCJEge87C4n+ET3nCMggAsHsxW7HOCamhHMtsm+5/q6emspX3ZfYeMn9ISM5oE
V76g5I6eOqKvjj3Y4SljeS7bHHvGuHc1oNsw7fsUjAHWYmVUYca3cBGGVfONVbPK
d2kHxKxnkDxJTdSblunu56FhvlwsNJmdk7JR8XROQx/78y2QGu3ZfY8B3cl+wu3E
qJkyr0oTKHkf3F9SYqTqMNenp2yZRI9uCb9foywrllWCeu5z/ou774U+7RsbkZPC
eWVHGC8jT5R2MGIJ64ZKzb/UAVRgg/NBsu6UZ4YthD/UhakHZs06NvZ6oqKDpCHv
8yJDwc42LRN6Yc+z6DdNzXPrUcMS8DE9tCfu9WGa05oHng9pK7P4+XkVN2B2KUBu
FwQKe4j1csJdIWSSz1gtDxhAGHlaU09GnnlhJ8tzOsPRkCJD88cCDJjlfd+0wiio
V0FXof1+9Iruu9i7/PyUKU0KWgWlCCF6/wrNamCLDYW3z9nJPT469+R6EMr0G1rx
HIaVO+iHy+iSH+EHjp/2Si46lApQxvY1eFbElk/CO4d6G9UMjn9KozKE/jvxO2G/
opdi8eJoxoIPg48IqUe6xCY8LyAFPUBPWu86aZtb1lSMZMCncJnwu03AHaUbWLpQ
MySHkfCw/sROyYwU6AjoH8V5Y7VuO/K4RGe9jxq0SIBzMJ3pTIQeuhW1fYJ2/6t4
uP8AFZqgF4cKP2/PBevi+Apsjl8y2AWTuwL0ZpCQFYb7G9sYTJyxnSnGOB/I/dJF
BHDGo87RPJOGuo3xg0JSi5NjNebtH+EBf7HQti5f3oLKF5qV1AY9VWunGCs1CV4u
Vq8/Yw19EdM/zihLnHSFIZKbbBcul70OtPBhCKnVd7Mehu5BnjBG25EfZF2fArtM
BEeqzneb7Fr4HeiizvKB/TE0JsCcftgrwwTDQYGcTJgqu2jvrLQJlyPokGLPeYjh
ns4EwdNjUhDMfPIHDeoAvGijWq0m1jn1MBBK/9x7II549Ahf3opuZGi5LQVtbA/L
cZ/KBP+hV7byAP7tmXOE4CIGjBxnWmPYVOseW8T3yofgPQDny7N3OOJ3Ir7KBFvl
085JVSj7Fqmiv+BS0OC2hlg2bxj8IIOwXg87r0bCS9nL7948We6hyPYlJDv+yutI
MuFUJGwVqYXHzcdGrLyyKOC8bx/Foq3Z0THRAY2du1XOyefziucEn9MAvZqOdwhy
3hpp7F0WCtvfC8PgkxNHkQQhUDCbMyI66CIq/PpvxpyF1nRsn86C4q2fISf82ORf
nbcsmx/TxhHgfOq/E+oUQPxcrizrea1QJubIbrLiFYi9YdSZICOGgr1Q+WWvUS3Q
XUvcA3Qtwfyyk8BZrLjYIcVDYKdEg72qgI585dKrs9jCRhu6sy/UlOXSjK2Oh99a
EmdnrGrgn9a8qoHf8Spagl1ODkZu42yEsokgJgu/p6wUNffICdEOcCzq42ayqpXi
q3vPq63DEv8G3rk4wA2rRNqJyTfQf13mnRoLAsMordirpfEms5hFQ9Gu0st4sxpg
ZY/pt/Yv0mawmWutlTHUXAbO2QLOLUw7kCVJCyHmfg+AyVBYb9mmj0a+PtLKVGx0
yfBJsRI4MFtbLIHFFisu1hNDmhH67ivMvNcm5Ps1aKwfnU+mi+36BXE+lK0OLJ+A
hFqi8Uvi+yRIN+HM/LbuBvcoa3a0N8KsH0fAaSCLrXVLLLz9TtRewMxhr14p0wXr
p4XiW/RiVSfUCshCXEI+/kFqLSZ65Ea5JeMenHQj9ZsOfRWFOf3pJBtx8vNDIPKf
IuuVXwaniwTMZNcKnRqLaGaj7hDlIQcqyKkgr+/3xi6cUZGAr9T85r/y00xnURgN
aQDAsfWfiPEKxjOnZ86G9jRapDoOHRJrXTRLKuAfAaAJMrC61tixyr619diKuCE1
Xk6nxmk3OZUumb0ROXZXGUcXrRIreLTPYrS/eEUXOz+XQm18P/d/0P4VsN3PFWsx
y8oDzsQwbhPtGxsGgDev576N3xuXaSLbxAluQgEgs56Zx46NzRCWmmf2/aaBcy7I
kVyeLMrPnMxQkBpc32GDxD5+VF7cuBsjQOs8x+ZsMCaejxk6c65U2rgRLzQXE5yi
+T9tmczUZRa6xmR6KkAlq0tiPTmFllH9DzD34eA0Zo0Az+JN1ygCiWQcPAT2I5fb
HV5pk7a99oaLDJQpT3q6yE+4Ex6CnZ/xYeSkhz3PeZkT8v5PBuPDplpcgYOsRvGZ
B7s4fVm0FOHSKazf43H38sFBHxsC+pkc/eXoIPLAYGfqYqSS5QnncPmCOpPVUIVn
Sd3kp+UhOcuvR8xpVTMnHKd2ONNpIoZPm3eoxLIxfmrj4B+NzvzV9k40wDPIhf/Q
LiY/QN6fqLcIQZe/aRmPq7xR/8JliXUpwT5XmNCegU/eclLjGlD6SbYy3LeGjTjq
lxMrKPwC3EDkIStvFsz7WTRrjwPAa1lW91hLC1wTyE8b/ZR8veykvvpPE5A8srJR
gp6Df3bo3J0R61ZJClP/TziiRNQUhcJ1txVDx3dQ79ipm5aEEr0RBiLdpf0umfrB
bzSjteMXByP15yimU5rNMmTXlvmwXHyzOfAQZ8ukatk+u+h735u0zsCC0MP1CJiS
arRBlxdDpm4r1rYZHcQpPsLTXPe00GzKAUESUe1TnqBamIYZXAEGuIyqKNsEIAu5
KAkfnzYwLBYYK0jbKnTILDj9clBz7ZAHTNM67Zuq10EHf3V97AsauyxdeaqQ74re
PhxlrspaXIUaQakOl8p0eOPJFAKH+c9Emi75Hotzuh/QzMhE26yeOwdNWuv2DUn2
zLfBGLpUhdIholhptzH/Br4uSyR3cOsHeyg/zK+LVxKavIeDPSglB7UzF+WOlCII
IO8gjIqTU3CngJNxLaSgMriLGcZtqIY4JRw0HK5QgHmnXkXRNjJTyPUhjP75YMlH
wMCskxE9SVH1CrEw+wCEqyVCdMV1f2yWZRJuzWtP8wjihwP9fHUgGKLQkjLlpyDv
/Xe+lJ0EjR7abEcnsulmnUOAt9j3NIqPI+TfDF6kmptiNAHFOZnDnO3xpDEGEUAu
Di11sz93KVN/I1QHEvc2jbB+LESrxTVgV201hsT+DFbeAuIorAY1WQtvZI332b0i
f98G6fhLr9Ld+c2Ri2AdIDQQvZ2KLOGdQocDLGvAvE0JhsZR2BotuW4/bvT13eiB
uExUvnzer0LWB9WJXDSFgLIkQ76VYkv8Z48V3R8CwYZN09BWR549hHfX2UUvVVrM
QvKHYpzp0HoxzBrTFh6xNefQm7Z0+FNFYkCor2+cjBJiNKpS80SYI8RVm+rdShPQ
Ah7xjL/1VxEG1GaAwm1O1u4583sxBwO/YUMJhZt8i1kq6SuNXahO5dvlUkcou1Yw
tiulV/4kcWaN+SMglY5ZRPIFB6Xx7Q2F258ta3KD6u3Je3F9GPvQgxT28WCzIr4d
GqqtCv2EEj7mr+PX46XN7yWsf4X666hdu9H5sHlZ9qilo9JZo2warGCpHA8SGDak
ha15DgHOMkCoUNGajujKX57sNob07vPT0zYUyD5LXWjPgCZUTd8WGzA8UOoV+h2k
aEk0ZFYN9jNzkJvVDrDWFcx8AJgjeA86n4KT2vCPz3TSx2w79/Hj77zZQANrVi48
aM8n2o9RIWFjGU43DhVDYHuaaAbyO1bRkSc7DeXyiq/PtbBMErTBFhb53edFRMG6
hgz+6er9OjXpsKCw+zCtkVdk1QowP8RzLXdcop1sRHAgK1+d5Cq6k/EVrmnfC4qO
tZDNE9mmLjTILOodtNTjBi7lvZ7WhCtS6vQlChN8qstvp9GnyE89xRv4N09+H74H
djn5aRSVYY0a3+09tEfkP27M5l3mCZtZlN7LJtWNMvDmgnVZ9AWQ8F0+cEW0oswx
ofByC0sXG0MMrCOXw8EJMjpPyD8blErx9Mvl3RE6aZau2OhuShjjVBwEUtcaJc+5
en+3rcFAuhHQo1kzXuG4dQwMGy+7gCczpfsIIKfNsB2EBl+hpOiCujx5nvq5CSCh
kMmMv5HwoEMX++m4+ww20zRZFqdxAiV0lcMLXBD0LbsUYfQ9vKWssIMxwLOkli65
buYv+2ftaD5FZmq645MSQnuq/IIje7vkNie7OUgs3sJUmsGtcjLaCqU+9I3gyoAH
CfCVQVpb4nHaXobkTTzZDJ78usu0ct40DyfBdhZJcPA6p5FL+DY/x9uOwYAqDKMN
/KhVvP0t5tV4HtPfIwQyJP1tozTuykBwmLWWudcASHf/URmoAxVrp/uaRIlxKnot
Dh/fP52Zml8S75EnlI5QeuvxJoNSHtH/Yfg6oFaK7CjvzJ0q172zpuKE9fVKVVEd
w2v9aCjKqnQhBcMuP3a8q0/Df9SWiS66Rqwby09OJvqZmGA4iu/stlix6AU+fRof
f+ooQ19+ee1Nu1ywT/InyFGzB8ovod25LgSBzPSlCaqERlvY/0Jmc4uJ663OJ70X
CcjZVGNu1QQHzd+IhQ1s2vvjiKMcGgv+l+1649Kn5Y7xeqgb5LbEcPdEbnmSjm5y
gW9MGFsTL7FnVsKS6azjkM1k+Ug3rROM2WljzMKhfn0nDyGP/5OHrUIRt4hGm1OY
sJ7l+cl0TIlsSgLmKalh40CJEmMnLI4OaUCo7QnZ/LtkLEQZVPsaltzkkX4yiDuw
nOYqcorWvy54FtTD2GkeOP4iR7pXaE28OxB/xnlK9iTrTWFjAQlST3ukf+EDAOtq
w+vF1rKmfE1HTzaJX1dgzo+7Fj6feXLLsAtQ8AicKTj7xvkowsHpcB6Kbv970gOo
EcUDZUFvytMk8qb7QO8+y3h6qGf+1DCXxj4nvd84gn/MAekb0rWRU7T3tvHpsFUe
9kEf37vqvl6FWioh32ITsqaWUpGvKid6EFbbZd4XJyJ5lPPGq76uM6M6Yg8b4EsV
WM5mxyjoF/1M1LuBmaD/FG+AyjYfOBsW60UCAShhwR/xwyJIAIVQ0LXLhNbM+cl5
y775fz1h2JxFrAXiOWVWmXjm0s55sch5KY34wnKNkcfFIBggdeBD90BzTNtltRZ/
9NoE37iXFaGePo+M753k/ojtiVPD+3i3/pNA8clwM/gqizms16byOyL+vrHA6Tcd
Qjt3wuSFcyFpTW7pNIwnnWYYh6eTinm0RnHMGtLNhclYJldZV8GhikgwY1g+D5hP
3V4PtiojNNXOZKEUr64PJO11JDUy/RFUBKmy/VFZfIqyD5CeuIb0hGhz2fGDCAfB
VQ1yUTibHdGR4wrJtVO77kr7HDySyB65O6ZDJPiqoIX7De66DhJAbhMbpxvnlolM
HZQPyFM8F6GXeoTWIjGmZBj6AdcPkDv3jwNKs+ONg52wmiLsX8+k78zZ7gtG/AHr
FWOrkw+XVbw6ufutGviwsUcu05CJFbfxvgpgEjU9OaSLn1JaABFp/+VtmISsZN6t
Om39CtmNzwMgmz0od0N0XsEU0RS+bN3aaY2OiNr2Y9Wd/h7oGtzCC0BE+ugtKiQF
h2l1l/ujvlzf9g0QZmTxOJMOUTuKkXmi1URbjkDel4He6TnOGqVTqBgqNWK6etoi
neP0IyyMGOCb1bSdShulXs5nXlpFXettRpVB8pwwt9AaePQXCMyK+nynanA9hcvu
nJktUK42Kf/LAEOzeYvVUK1Iqu9dmwQg90Dy2Fk22Yi9CyS3IwmIs+Hyb8Eh2Dbm
n1TgBPsCcIvidE6LvwNXGjqj+KeE9FpjxmXEozdqrjNICePk2G991p8YLSQhQW2L
tIh101fJhNZg6c2YPDslXCIKfxM3uF0p+v0tAYIUN5jUwlWgZdOkAPVU8kHMMJxp
SNTV7UZfQlDn8ZmJCqu33aCepVDKtajyhoQNwLgTWh6uev9IglMQQ89nJvVFxf1V
RAAM6MZqzGbxl1qIgT+Ml5Oe9MrgiMw1pC1TuC6rzpChYAlzEigstZVpISV2ITmV
9YgvoGeze0X5wvBZeAOG85Rl+5+wElUMx91jl6+7MX9mv+UAt6ar3sKoXcPGxedh
JJtsqIvtwPk3T1yHs0+1zAgUctiFa4qOWbfQhM67aZYEU1Wb259yVOzul9Fwzj/g
XHbH1UZMAbpYuSJBufNE8Rv6lpqDyXH9DAFsp9JN1N9z1MYY7YjPmQNc0ioe4ORJ
qpCsKFNu9qCf/43+CUITfXRmeFsuQCklNh1mIVKDcAIIjgliiBrn+z9JfYvWFaaA
zAVmOWkkVYZ6kw2IQWjqsi/87thgox3jbe1NRoF4cnXiluyFN8rjBxzRMU5NePSO
UumyIAy3oGJDftHvR9zGKYiu4uY48HuCdXITn/2ocJp3pc6eIVvJzR5Acr8k5x99
lVRXy2eB9ZBkGTuUmHrMetgXeg9LW2Ar/gn1Sqfn1ZwCyaasmXU8CtHfBF4MZ5WS
LUAkec7S6s2afFoQoeipuHkBQ5wFkMVZEWZIAE+o/pxGT09E9D8waDwScTDasHW9
Zk/6TxH9GMhxZkjxiudgqPw6Voli+/cjfdL+MnhUaQE7kc+fsBeVrrfirbQAzXcX
DXcZUFp+cgYSCYvSwOhjSPtiCrWIeSwVOoM7pKyd+uUeHd+gL94x5U/6QD5fbxNW
hPrjc8Kgw8zL0toKq8dhNN8/OL8//8yiDPZO1cgj64ZWyMt9IaSfOQKTqrqutwyn
DQ8SOlqFkEFddcs1nNZ3SQKXpe0Kar0jl7HB3WZZoAIJwUBw542/auJDisQIIKHU
T6DF1GGa9EVfWyEMBis+bHSQxIN5k16E8N3XWOiQSyq8niKCtVFXS4Eo/35Zf4Pp
EG7QPBshp6HNoS9gdcIR5M+njuRunOUuIu+0ez/pa9g6O4Fiv6iVazU65r/2nN1e
Bz3Q1Li58c67781zfXgjUIJibec5sBNFp9JO+rs/ebd6eJC12pQF8o8uSgaMOg68
q389WkyLd9hBtDEhBhIbP8Hno1vSdOcJmcAik2myJuZr09DTUxDiZNbfHkDf442l
TptCS1DWA0cFQl3Gn/ZtJa6mNHBPGzNGkJ/jts2yYouihGXcDtp1j+Sbd44y/wSW
qYwrPDj4ug3l6+47cCgRDhdIIa9zUSbcoPgECsSFVveQzomrfNDHI1Hdj8Tfaz+K
HNK/LkbIbTzgxJ8Ln6jb5dgbBou3XtuJ+wBlCHStDwfQPPAMZs4kH8Pvkg97SikE
irs8/7Xt8bCLqK0n5pIRZEhg1E9aX4/ogW5CPV+evwW3J9hGkSkf2jgrtzaZJkLK
l0QCL2YJXGqSKHcsMn3WgU1vmlWf6jshRLsDdLH/8N1B4/5OeaYPdGYEZ02UT81K
3QhnFNg9dHC/rbVgw0ighbA2TrI8EjRutQ6y3hT2vlFz0tGuppW+fYtHqjxjA+io
V3gTKzOANo7A/ThOb0W6HYffvHp9k7v4VQKaDfV26yKZOXFoiFEbxsKs/7EXlorp
ItX0uhNJ1kDJulgNWQccTPlaosd1L8wwWXkWUKoIjgwOxZDet+LwSLkfrIU55Alk
LRoNc9vkJ+/zmHfV6NGYljtLLgfINQ+r8IsyrNkU/kwkcfxE4gRl9Fv3PKPHB15P
VxvS1phaVZ2zGB+BLtQoyH3s6y/QWpJxSfh8SGVc1ZC81hzttzjPPzpS9nWQCdM2
O2HQMJlwcKOiXcJ29EXZfEKyNEAOLit7YJMwEJYONjMkxmca8Hfo8OjfBiWrHhNd
5jRCC+1KC8oEu+CbL/xeFvgZPhYhFWuZAUq6ewnJga0fSyPrQL0gl/icMSwqbMfS
2espPuWex7JrG8RsURllLfSL7HxBDiaWDp6sc85gQCnQL7Ix2V2FPI++3GDA3UwB
lJxRYp0dHXce1LXZOtHenoAw/IpGsL0XvGLGwER3f4c28pjIH5isExe5r6qH29Nj
kpw7gWn1NJSsFr9J0YNjJCefTpLR9AwxCm5IrRFvkeC2zC8TFath7LoPUV+Fk/g2
5B591F955CWDn4fxOjLob8VTIzkfdaFGQGLjL9ix7xCZXdQ/kCAYhgQkH7hzjdP5
dcc/5fuL8W+Q8fS5j7K1ECmACuDcpetPflgNvjGZ0VPf5uz21giseyHpHtojvYGZ
qU71Anx3zvV/BxOKGj8awKRJRfuuvbYJBaoBsFGuA9naMndL5T9bOoSsOqXdtspl
yn0dbffxd3DOdOgvZu3KLeifg9lwv240glypanZG/sxrjtUe125ZWIPYlJt3bstw
n9yqW8gW172rnnSXGfxA/bWLSrSjjAeTk1/UkcjcMowI0m72shWL9+y7AX3tIVn7
WfVvwpzoTnh7HSSy2mylBVbEkCILSfVqLG8c2Cg4QJoy8lYM5ZDgJNS966cocjg0
+YfodSktf6d6ou3cw4p9LL3kP6e7vgf2MtIBLNsRQmF8FuaLoL00LVDMGYdvgfin
2D6Mt9W05iCoWG4zD7fzH9W0MjLyRK2mQfTmB7ceue/hetaz/sJ/C7mYDos5n46M
KiW9RxCPQkPA9lD+f9poxYylBR8sZMjQazYqcfM7R88yZYchrF1YAib2BGkQmHe7
aBuMOe+YMK8n0shb6edU/8uh6B+cbxvbSZaYdVXrrZzrqhXvYmGn5LQ9gjbTpZU5
zILIy1PgeDhhIpy7Jw79c6Acz68UMSm/wWBqwrsCs+9o+0UOe8qUKOBnpzPrw3lF
tL3CFCvHAbABCStbFo0ybKKNkLo2/zBy5bzFS61s2p7MEvCRU6u5eidwlL2nmOLi
iZ1LkhXn5MNSz9WzX4f4cIR2NGnfFCeDZVBP4C5v1Pv3P9wYTZbYUqGBk2nvh+qf
Af0gTpxzzQOCp2Pa95C6U0PNX1wXuh3e2J9PZT4UDGqjKyrduWQCR43dl9mqoUYs
bponRMCahMvpRFjOf0vTfjgB6WolD8Jwiy953WTaxnSss2dwdS+c/iIBtagLlWlh
isYsQezbH618OmCEasuRRQZQsd34NruInKmhiuHCZBVH0J3SCckEoQzFpNyc1b7Y
XriZrVw1B1w7qwo8ep0OKab+gm11uiBo6HsXRbUyIFVPLYorVOwdsUUvwTnjUSg4
v4SwhU5ts0aRaGludsgQwjSh/I1ExQMm4PTYQm6eCL3DXdUDDlD9cpiaqCWCC3X9
fqCgL9223SoCYB9VeDCJLkfXq2fyk1POkxbutOWAIzXi626vL3i0H67lgOCAS4Ur
bOLc/T9zSMux20dlsQfwYJQIHMif6q+HldMt+JLo4AAYnbQSfDA78f3ghblQw4uF
FYxYJYBzAjxdyrhZ/u6bjOlfbcfTI/ZlKm/Uf0mTqBeKYeX16ltRBHqPMllRwItm
mAQismbUARCKYE+fwuZ+NnKPWqfVkbV+OV8GhgTYfI/tImGlEUiIUREQr+b5k9SZ
jVRqukntKBmsW6Wusv2/+Ql4D6UYY+k8rL8Rm7IRYN/2xr7nOwNH2aSt3dc8BKNO
qZxZeH4FwFBm1IF7nNiEs0CuN3DKzflQsT4idYkhySJq084aKIFVlUYLTX2VCYyK
BuTz/j7uUkrJ3Wf4s2AFl8R/PhMf/fXuQhA0kiDSYqSSbxvUYrIz0jshfP1cC8lI
Vs/xIOtYjP7Dq2C0t2YaJGZWhWUnRuE8ittNFe8DmE/mJwJgDO/bLAntrZrW8qke
kEayCfugvB6Oq0FjSjRLwUQxvc5slbN1fj6kjFj0qYNVvpGoqkWxnT4PT0vqQejL
cUoX5L8IhAoKM/DlpKN0bqoVyTXlG634n2vvg4ihgN2NUiQMOsx3/MgGVixk4z5f
FUGtW6b8krD631CWu1RMzcasZZA/qXna5erEAcyTDkDLoAbTWkhJ1Dh3n7Wdzc4Y
fMKPakr4x/9S2qO8aRQod347ewOa8y+KFvXwOoALFO/bJu8qQl7R5c9egMs3E4w1
wLXARl0ro3ZEjyQSs0ItsPmSOa78kLeJZ241MzgcOBU709rijaKzlNxVH4suVPk5
kxbAaBgnbTUgh/OA2Mun6KDZ9qINQkFJqyzcFi2+hXy4UB1v2Z3QX+Zt/IvvlQKw
by70cvrRanRVV4e+mxx/zZ8RyXyj1ZTOrTZ4wNGd8ON68UI8ieCRZDxhbbBc0yQu
Gx8+yqUFJid/UctJsAnRizhb0OMlNSwwcw/KnO+O0C+ZL+dO63hnDC3WvOmhO1SB
4vsFRRv7pXr8IgyGs/57Sf+FSEpkQQGls0uUg+l9Sw3PBsITDnMtObwwt2dHu/ko
xWQZ8XYT7np2h1PnXrlk2BwgVLBo2SRZVrsZ7+W+8AO3f7QTFLZUWloUL63G0pv3
aCMmbspBTJl6WnK/kDtXjdj5Zxj8WrA72VpXtJJ19+2jdBYtiRxZBdUUC/Z1KvfY
5NEROLNCEu/iKGuNRyWdk3GEsL9KLPOsAUoFFlcAmKiJXiqryQPCNze1cTRtRItG
orxfWVneORlRbrzgj+kNWF/Zui6z2WBYTg9HxsnIvK4Np20qUWNYruK+RzJDuVRj
gjdwvGoO2nXViyAilzx8Rtp8NqmoXFd2k2DIxXo6yL3e2OMykorVNfZsXZKjnopg
WcI5gShTu8qBp22JMvO1OOsPbKGdlTqF2h+eHdHr2gYk0efRI4jxvKDcQ0tCHxOb
XxuqEuKHtufBiRLo1Z3SjthBHys1Pox/AI0JII9B7VU9NhqHoWPlh25lNmE5IwZE
XKJiOjvNWXkem7/9BCwJrNS0w37NQK+p47Rw7uB+LB0IlDK6uZx9ERibrQPP2m4l
hWn9c/3mtQiqtOoaAhCU8OpjSZb2jKdmMTRh3ibR88DDpNj1BCaPclXx/wOoqRSp
/5sO2gjiByUdm9zhUu0eyBtIV/BEnNjBqkdfuraMzjEBgpL6h58pxqQwHffbc20u
JrhQr0PsAFXpiaskaW/gPE6r3eFh0S9c2WTwcGZQLsY36nTWY0z9J7Gjkw9SLGyZ
7ZRj++y1GBLAogKFPekCegWTtZhx9JaIXh/3X4kfFdaUkyO8Zcb4HCs9ZcHAEVjs
OIAgrcCMjQp7GY2rwnLmV8/zyUjI/p+9tLMZZ+mHRzMwXRteIKNxcydmaZTughXE
rDlljC7dvADK01B4R8F8614BZ4hh1SBGe6RItG1w+eumMr0RmT745r21n+f4qc2C
zm3UlHC4HY/7gWTP1rIDjrsruBduvyi/XvOHUrDfAmPvWeP5NujPw5fgAcQkNyXj
hWAPR2mEH+SsWVkJlRVLy92D5iSIenAyjoqJONKJdZt2rp3oWtro632YyJDgg620
1rlSVJc9ZKNuDRvHq7Wwt684mPJ+aEu54KGCQp87vo8VAdwgnsyDzj0W+TyJSE3g
Jc5FLe4kvKFjXnC74+lg9JmN+8VKEsbL+uQ/LNEUSjW36HDP0S0aqR18xoscvhd9
70kymZh9R6CIbXe6+dmJ+3CJ5O6Evfy8j/NoDiC0RJPzPHiUTk2gYvWQ681w5hWM
fXYlzKlPuPrjvxV+e7ZMwY4IkiY1u+cX7OY5TBvsPo6RSBDtnSJ5HB97jA5Mh+9h
v1/KwN5iSc7kxDMxC+4Vh7sQVW28dj2Ws6jsye69f+cwJ3+qcq2DhD+ut01u0tyx
ydq6CI3F4DttKPgt4NgtF3m/0k6gMhlocZkU2Y7mzpPgLo6P04XmoZsDSwUT7KuB
cP2EpudKfgAJ8YMjK4MfJJcSLIIckyFAsNB2GgnAfAXK8XG+CVtcw7Bnd2RTgcp3
C9C+BfhqXb+iUoLEUBmSQQY4yU6Qo7W/AXik+YErwImujE0ELOfrst6uI7UuzeAP
WLlTvH7q1faRgDzVLePfPaAZ1II3KZ18qTlMRYjfpP/wou2bIUI1S2TwNrBV/9jl
io4hd4rkrMO+l5KJLxUzYs9+RVLbjj8Oh5cX7Ha26r9EvZIRkbSLc7DzCZcN8ags
88TzX5uKaT/ucqk7VU6QULjSr6UNcurxFVjT9UcPrwe7aGBNhwvgYn1QV0lmYklE
puao1yTiEVElpxM7EUEc+mabB+leu1kxXUXcSpRfBUEgwW9uwedrnNnn4AxQLvIA
yCipwuE/uCsrncKyvUh+ogrKVaflz7WA/vT3avkPEEQsi+nFA21G92ajJOKkt2P7
JiMTddjjWSStTF0KTiXjw5tEHOgPPvShRXHQxVsVQZsQUwmumHFAAM7/Ag/zSKGe
uAtK1wMCWgXbaB2bXDnZnL9+dAcPEIEnzwvx3ol5BVxKNPw8UpjQ8aBsdynI1+mr
ZxLPLiMO6ek6/+8LdzXMihXs63zGSSyVazWvZ5x7TNY5tN1dVW2VmjUdnedrA1Sd
z/7ETCdMQJLDEAh1IiAAoukU3N8/1B1dIrboOz4u8MuA0K+Scn7Rr09YKloEJRIi
Ouwe20MSCn88HOZUV2tf1RBYqcSMLuYHmL+t9dQHnu02TGoXmbvvL2eC3DC4Z6vw
zIF2Mc7lJsfZ0bXK+mTLYOTB2rYXJ9LpLW8H2/vCBk3V4/9HLnWZiZLQkz/xNqVF
hV5t7qHU7Ph6GN2tUpA1d+ZkW3RkhIP0gnJ5irRneOQnd3hhVW7t6wjq3jWVE8Xk
L4wXPo+eM1HXbyvYZQHYkPfg36HTK9yzQFSM3Aj5oZLdQIJf6XNvl+/gUvIlc89j
irmuy9vDmVyN5VNwBaWwLRrW6D9VF6fw8B61jUNMCyOIOFaDkEy/OZrhkeKayAOa
hCYe5zRzKuQxb8t1ADlkF4VU1pZw6vacRYS05S4vdu7JJQkvZDMiXr0+yXOzgEAQ
gT+1yD1nB3fJL6o3lst4E0L6Effk+aFfcwCpudnR+gCv0gdAa6iRoNNAyd8jxwJD
Gq4A2gVeraDUoQLQI4scerU9ApKyvq4iw789d7xwjL7FIzd6YXrz6/I7LAP1pzQ8
cYzAyBo7znJpiWdrqotduOp7t4/mtkl9/hY9lmw2yjzEoPJhYPzMPlo+AZo776zM
fVmjPN+0bjEUXEnwSv4Vvrl+KB08LUH+GFoxdX2s3VGmT9wa5fFrJZYqhd7OeBtl
NIM0gDisiNAX6ESiL/IMLvuYkZPzAvcNu16lryzhfsRz2UHb1H+Rn307otGWhGvg
INNSTv6uE0/nypHq/Pk0NEZLXWdJDza84rbbGDBn4bAF/CHpFIF3G+fx1ceU5IAF
Il+NQboDRnkV1NIrYSsQ3XppEpjCLhJdegexLzqKg8D7z8zFKHKw5vp/bE67pm9f
HVPrHgoXnw7HMKdy3SR+/dsygkdxr06LyM2WiFtJxWeCzJ+/7WIegpvDAm7bahDF
mTR8naPrseB/DDaQ6HYjoLYVP7FWyxHwMbhhYyzz48c8wUlqFN+V6AZqbYY2yzrx
06KIdfkmkKVd/kzF8qibhaSUgqvV+nSwMpwFhHf2iX2/hiY8AR8WV5Z8Wg6ZkpqG
CC8QpMPdK03K0V4h7S644EuHKjVbaJS4A34APeGOBc5U2yDBcIcj50e+KGOUZzsb
+dLJINSQ6rV2JC9j6mHyEGecpKlLn0kLJHrc187z2VNyp49qlvkRMuUYz8wPk0v/
44ujdQp3jXVwLRab4E9lcGLDJVU7DFmU2ZcK6F4C9mZdHQNbtyH+tFEuV5ACK4To
L/zgi8MRjzxbMxn0CO8CzqqYDxO1sk3F37LtGGmG2OiaQ0LpxhQhuf9oX4Kqteot
`protect end_protected
