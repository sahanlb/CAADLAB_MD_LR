-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Yc4NcnjzwsuEkWS0g6Ms7SpnURrIC2Cm3UH/dRB6MTG8Lg1fs/qXx6fJ3b+gYK6T
As+qmHzgPXweC72PKKKrc38bTsYmsNbzHe4phKrxRWKxCrERIO/TBJT9HKfBup9i
WqZLxRgKhCC1VBGVWXEghvImv23xxcD6JyaO33eXAls=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10688)
`protect data_block
pfOQyQxlF0Iq97L0NJtVbw3j2MN67NMb/y7YYQu4314Y4rimf/WRDq50btjrEgps
3jYEfCzsJbAaIM1WHUwteSCcjF6nMaWPS0357AbGerDwEFHybZKnjuWwozqw/+kX
dFGNs6iI+7Iil9IGhC2DtZsa9oSbkRzB5bGeqFnVXFl+nRZdObUtP6f179byRl9F
Rj3rDyzmY/Oq+ntDNDGNjGSYFxMUiWxLSIDp/+4t4hy+RE0li0duveq/lQGdDUnq
ONpyHvdQFH2Q5SaxRiM/g04yFvi8q2jSxiGUMXgfvjgPWhhF0dVs3579jB2V03DF
JtZ0DddkTfGNKKiFsPkqkNi3s2iIW8/XrmYima+rxNI+MXwpni+v11R5j+u4IhHa
G/I5OmdJFzffIl9VGm1hC/HvNteb0N2EkqxEbk0bz/Pu12QDbDDsDA0sQDOzZZa1
IoHRWVSeUbtGdZHbt6vT034RAZKkvlLiwL4nObLUtDZgskC615ZA/Vvesi79U/c2
TVPThLF7Vgmz6vNstvj5akParWEUyG7ozW1qJR/CC/aVlJxENWQkCpReQfcz0Dho
GlUaWfw9MMAKHSxZsV1Yrdksj9CBq8K1xcJN4Q1UpQqgN6hK3FRLDQMR672QwFCD
QVm90ECFYJdYlzq+J9dfqoOnM06xrCqe1VJx7X8qRa0kk/Jq3d0cWjKynPXB7M4J
XBdJHGD8DLZKPNm/J9nz5x66Hog1suSEiu5iK0lhWWdeg8kz78E2aviqkc/SZFjW
LAbZtud0NDjUkaK3LQt/dLEYz4NWL9749bNCJXhOBAduEG/zP7qxBMojv30bZz5O
bEkTNf2T+I4uYuhvaQ7Xkv+Yzu4T2X1mBRCWmeWKBqbyBhqHxYzaB/Jg7AJVZSJ7
YBinN5S0DPaGAHnXBdREWUhddN0VAf69p2K9Zv5WdM1ccDjuQhk+bM1G4bPJM5li
G3saa9AYDOUpkasaDoPpUDlBrn9gHJXe1CQnm8kWqBtYyItJmbtG/wYy2SQI7TNE
A7OIwk4NfqNAa3YOQGOrTq8AWB6UIqN9QFowKUV3ZNtFTU58bqnu6I10HsgOkr1v
hWJd50nL++f5T540nwBwGkuS3wb7A68aM4AMQ4SXZ1TOlumE4SymTRNVsP5QYsMC
DvLRsixsgkHII1dSmJxs8FBWobxphOztWnWjrk3kyi+7rVN9uiOu4i+khIGuvUXC
W1hfJhBIOJUo/JfH9pBOD5CQN0uxE610+RzsUSaGxzUqEGpKxRa5bc3NTC97L6jF
lzPNKgviDOJ4Q+XYuLeG5MkKlTZSafgwy/EPmbUbDlKcilBCtZHqIj5eRTzizGWH
/PiTdMhikrPLr8PsQmxyKKALgoAmhBMMp070C5lFEi+ICVZV1hPyItm/p0dJIRQb
KvEwB+dFJ09e86nhNAxnC13Ou7ww5GnOuoW1QI8ODAWA5Q4fYF+sBiKIW+2yysSb
0JzbSeXUYgjjab2zD5TJZFcTjoKn+hqxz410S8Jxg+Ouj7/Hx+Vw17BsWRmmmG/7
oZPccXzcyeVK7VpI4DysTvjSNFS0nX+bKxYGuft0LbOXzQU5XpRRyjbd51WhInAN
rdalLzX0vdqljFCxHJS3BUJ9csfK9prOUSWV5G6iRVDnP5FTTft4N+p8xjpAbyXm
AFfJ+V2pyfsUeTSqy+J0qgBEnQox1oUYuecZP5PeY3YMffvN+Skhdvzq8MI2gcMv
bubHm5e//E2AgX6cvrkMCH4QsuQUlEVlTbJFXiX04BXMCcl2JXYJMIZ10jth0gJ4
15DaoZtLw643YGXkXM+FuR3ULAVH83BDJWr34T9kwDalKZZRW8IByT8u2n8LnmQ8
Dt7D59PrcVFSvRIMN1Xt3TUCWkKePloTlfz9CiT6Z+SAEx04+9zCHf/llBv0boka
jLpH6up3BdaavuRXFUr+sW1ay3OmysiZMwa3x4LfNK/15MfAaw5S2XadK6ikZ06i
axU8rXgf8FJpm1QYmKzKHiCAYr+hGYtJZ6dCn01796egLDJ3qG6CXqrU8oD26tqe
nnvjNACzqP0M7QDFhUOBbebD1iQ5bdx02xo51a0KVr1Q+ilvBeT6vgPkaWEA1OhL
NIZGky8UnngSW+wVaBgYBDQnZyeiQ5El0Nlk6AkLYTI9uJXbiUBYCph0xQVCiZ2w
rthhF/Jt8hxFLDtRj7ne5cP+s14Qcw7cHG9y1FVu8nYzZHxwQzeLUeAR3aNv2Wz3
YBKDp4rn2egfKMUXq7pZy99wjwhHcNPd6gPn+jioo+JSSNZFBNtaeFwH0wmhfqJx
CjZNQ+W6uhgWbHk2V9LLTlROPwmAjMFf/3S+rnlcWX/dpNbbGHEanvt+0o7vwUp0
zZtNJnNUkRLTOUs8YQWZSIf1bMZIUoupnOLqkK039P4+rK7tIBevbSag17Ea+Wta
MXPXyTYKR0vYErmTlTI7mcbiaqgbdxJqv/MlJg102exVn3eaFWFGIqTzrJ+REU7t
Un7WJRdyyrrmM+aB+UArui3pdKTt0dAYNgjmbQaq59hCunCFXC/jAot8XQtBhUGB
XMo83/njH+BZzuzAnBYeoPtpNX1RDNtTthycyTjKYVdIz6sVlJt+cW02cM09YThD
2Z0IUe7BSNhRNgAmYZiYCs/P/TSoY51i5TK+wcYwDj6Z4rTUwgSAOFx/hC9xngdi
aoatqJ2zLHGXG8sUFpCEnh4d5yWPEwmKFpRB+B86fPkgvyNamQ7tZ8V+/LVbV8KR
+ROr0dd+n8pvN32zoccJtN7SNS663oZduQwhpc3cR4lw7BR37bRqoAR8oE+B4ixj
WDi5sM6aLd8G0V7FHva0Q0ynZsyR+hiidDEAmqa/SKwHxOy1WLpY5e5gngOiFY+y
kNLk4sG7JJ1sLNPPoTZQOr9VN17rS/g7zksvYU0B8bOcP260gNE0i4S/JOdvKAG2
Mo3PXyCCC2Hd1Z36sQQXUpewiaINeZr0rJ58IH2v3Edq8LPOlI3aEq1Zzny3BhkL
7P90BYn/8RkDue/ZS+VfmEK3XmM8S72HV/LD4+vItwgV/dW4UTXNe+a+GBXufrNQ
VOyW4+zTJQRvKRA0ViGPpv+iaZi8MjJx62CmaiaH9cyyqOKYoT65rdvHFXKQu4xO
/YW42Vq/tmYnw8aF1/jAikTGWOpbtbE4321ylpN5fIaWagZ5z20QeMZzoG5+rncZ
0pY/lrWz50miPCL/C10NUW5lql0OSQIpwQ1+qzTVkauUA/Dxb5OzWdsvv8pdEzcr
dT4Ui8MrPBgkCd0u+zk3qWPvez9tVARuRz72ODNUiJCBNR3oFalKGv3ymYV5nbIi
Td/Ui7TYzPI1FQvZ8yxrVWXvEVXpzOosUwjSpbyN5BIyVnq83FvfZxIb1SmUVimu
jFWWNHr+vt1grmb944NdKZzB/Iur/FAByI+Zn2eBiZFK0GZJryw2p3ZCUUcbdWO0
92VH7E90Qp3IRpL0AVrO0xHx0/sXiJdGf2h7PFx8vKaPfOZKBRuxRJ8a4rB/JSQX
1rKj5eHJ2sqiJNA19SLlUhJwfyOc96qo2s/QBfMvDg2/BGcWtYRu/XlFmzYYZoXu
m9dE8csCM/0vzkws6ROeDnufeai9iKZJY4WNnvw929X+BQdtT7mwEkietN2+4b1m
xJ1EcGQd4PI5+eN7H/tjzUDv3kPOTUf7bva1zh1l4B68iT/ATw0ZcLgLLB4Vpbi4
QraZ8296Dieat6euPGZdwm9zn28z4+09gHQ201rZrnk0VzoWIOpJY9MIJR3R9cFI
HMSX83CSJhdgf6+CXa2A6AhbMcygeVfI84Zcoc+RqcVbr0h1uMPARFM1aPFgX2qz
zyc1LIYSTNgwNVfVs6JoPZ9QRuctsQYJHNfSv5VOKGDvHgvDwkbZX5u7MJyl7sr7
oicLhQBE8ON2PWh1POLI8ebbayxLkgQ0MwsVesH/1XN4PJYBn9dHDdpSxlxgEDx/
0eQlBe/C9+K/XTeO/QE5SL/hjIgbqsWChcQEyn6yb+GHvYqTQZFjKCHjZwVPDXFm
cKLPZfbUeeeEkoRroTHXWkS5/6KMMsKeMlasWFZQlNN4yT9USPU2tZAh9ICXhR2U
/Ftg599Ji41Q+7zSNlopaAfd6RWaN784yv1hzt5t0xqCDVtE/exnOzKF67ieS9oe
cYYg/6Zw11r4O3AYhoj4m6bC4kdlVUXlWF6YKRs21K3IxdRIbbO9tK8mc9sB/yrD
9Gj14yxjVWNRbS80cEPy4OL+AsEy4P/gCc4LD3GXUfaROodt2NyU/39TjTBIW37I
7LfhXfi0QfPuY4bejh+o1dHnT3Q9Xo25fiNMh9XB7K6yAxl6bFnNdOnsj0NeahkQ
F8R1hs8sSCBnvb9OuE/NbHCjG39vLzpa7gZTdT1vo/w7i9EdhTaMknEmSevx1epG
7dmwUxG4KLrIiiQpuzlZceiypYlGmGnm0Rzkyt6iB8bIIoUkoPErMqesmpZalR4I
YXzFm0ZSjKZo9J5JFvOp8aydlea6+C1ROoIJ7ldSJ6KVOr/EkmPddX9qd/Oh4koo
GiH9+y/TmhFxa8XaWLy81mLqdc6HdIMDGsAmWKosLey7IBfHDEbXjEh+tPefL3Oa
/WvMftYcC2MtPYjPlcTBtyVdttmmeOnnFM3b3Q8oFosj1Ul4XhEkmZrB5SGni78d
iy0zLrNwZXxwp9IlrKAlPpaOT53GtNvXOcbTM/CIzM4ViNHKnEAtZamNUwsp100Y
pVQpbA1DPVOKS5YejZFLpmjb4RbNY+dKpQtafIzlzGWfPjad4IVTXD3Fx6Papi88
GhUWGLy4io2t+0VZ2b//JI3NcGisV9ymcN6v+XE9rDzk2gOTgmi+SUD8XGdMAxuG
fEYK3eI9VeEDKVh4Wvi25s0JsJZk0Au71l2cj54VnbpKNR2GsHCnNKGYK9Db5gmd
sHZ0mFaAdDPha3XDmSuJq96GAURXwCAPzuMlCKkv/hkPQCk+PufnYCkvUHTdCRXM
m2c5qAnZFaPe8FL7lvF9sq+Rxnky7R0ZiShmxq4POQyFWGHBZqrcGM2KfL5PwO5U
IoVo6F4zRuA6b4arf9xGDlQzvtFuYxQ96cWomK85pnRkpzNMkUgrANiClxi4WOWa
qXXdrAfSKaBy/2M84AKV8JQj/47D+iqykQMR9tbj7/W7lcEjzT/Vwdd25m8unNgG
2T79TN3r5s4IYAOOCCzvOTof5TOfUi5UVuypfl+ZpzsLgokJxoREBbXxDAzV17n1
C+rtdvzkn1XvHJoN2tAiqiJyg84e42HJBu2TFDjLHCv922Qqpf1mUvAPYBwA5cNr
RqwAY3NE2Je7OQ/KeW6gjz7tV1vbtXlPixeC3FyNghcdl4bj7aZgXeg5WksHGUkk
bPMbuzyqSufx//L9Rf1uYaRGi4SRdKKK3lny0YsfVZz4GCUvwQ4uQtTPW75GWAAr
3vqu6/IhBkOYyiKREYaqXzip+7m6565wegYXX+dzHNBeoP9hAmQlTdKP1zzFJZXf
6z++OztZ9SezDQN1yLMa2q+oIh2RAmoq0CR8DXkkdfYCoZeIkBe9OQJ1v8jBbXsR
SV+p6h93KEPiV6ZEM+XrJGkif29ZPpvUDmjqHJwWpSgfy9ToqB3I2fyOcbkgOvLs
Fj9RpdBUKcysqZC2uZ2QU7hHk3Cu51mVm6bdjd3SRa1UAknB6EUbgce77NuWDbDO
FdyHNStrO8hgtBH9AZbRzQ/w3x9amC45ORJ3U+exaqUp6tAMXOmpvVBB5MYxWTrf
1uYByNzH68eOE3EDLxSatsPCVyftOlpy4buyZ4vkCIF9fg1CitTzXTWVA5nrZf7H
wKno6XmCV63AtOBRrr0PQlKdDTGZWVVNKJIECOexDfQHmsYcw7S3lL/0YHhDoMjB
ktYf6eO3J7JtPJvo8ZLBqVNOvZzCcaUgg2fs5kkNX93VsUxiSE+1uAXuK3DIrj4D
V1LvzAWXooYaf4fqQEDnPETlBzCS805nLnq1ywOJN7WOBzneWDbJoz8gU6eBdy2K
87MBxDGKz9Pc8Jdxqz2JAzIFd6dLYjbpeNQ7pNWkDmxl+O4d4DcfB/0Kej81FlJT
8auf5IW/6q7vjCDyW+wuFQVFs33BlUL8jj8qFNBGC0AKc4Q8FNknGXD2VkSlmxzR
e2tik21RdQTrfn01NV8ZbzrKbRauvpkk495Tc6P/K0rXByPm7GpbUKjlvBMFd/yr
2HGq6ggfxuf9sQIAwUlmxlOr/6k+s4DpOeui2YTVkqLgr+tNiMcO8jw9RfMdsMsN
Jmxf0a+0x/yF1uA6W92rxYC7Gor6sRhKigYCybZ6eR+29P0BVtUgBfJa72fvtGXN
dZboxhqn0VMW6wqswyMcf5Toirld+5QGp8vXvNVgqdaMEpNM5EwIlfuDQvZzyl4W
lJIhzStLxPPtPyMX6qOcne+biJXS1hOfBoGwyl7+lRsrgVNVbYnbWGUPHJIskhhW
+spNhXx4azt667D4SA5FTRbbm0LGEQeZ721alGEiUydoq2kEd2Ob2LFyS18WTo9R
4NlLeZALXAEMiQtxMcuiWijRPiHX2JrTEWxYSMwfIc/G6/V2JsxEVNXVwL+cw/yS
9IFPoSfCo5VhDAqJU2qoC0dE9V2u15OvW4q5RkuddIl5ENfKPO23KzeSg17pKo0N
VUC47yHhlYC6tfZCJelC19ovUodFbMAwQAHTxz5xbRUaRyQ5MVJLUfwsZk0xF9QF
FdX1u6Gy7ahjkda8swHDcyB916IVJtVBGJtbbpWtw7GkNftJOUOkyc7KDGOtYf3d
XwwPrnNisMlZZWjj90Jdzr8aaAR87zujPNpzThJX21t4htmzHBfnMLmJIXbH+NKa
6TlZELRKTFWiFLyYVDoohBM8+bmptFJ4WNArNpkbvb8qnhM/ISypDD4pba5ai+zK
u7TLuDwfKukPy5PTtryco8iqK7G5t3lZzGdR6tTARie+YL5pG7NcGVxmsH+Zu9d2
LHpbVeb6cQUmBtdneIHzXFqovqR88bFGMywFe8POTKOYgybHVeNnX78HZRR3ULe1
Vu+RONkD+MN+E2CDBmmWfy1/rXydw9gykGb0uaNo9ktrfp9gBm+sd34cARUFLnfb
PruD4I2h66i1PO6PpqpbRyzn9KtsCPt99FpibEV9mXFWWdLqM16zP4liaYwX98rP
lVyo1alCIPzRiD/X/sVUhsVrSYOhKQQyo6K5ubG7yJucjnuJjWCxEX3vIPke/XFU
cjdWqJoyhCIiqaxW9rpRIXKiEitxIUXXxsRmSPs7WvQCFkgp17ZYBEjhE2Yk78SS
CYt+HYdoqQz+05IAEJykUd1J2kD/CYOf5rDTffiQf5PUfUo5XcwHQbNbXFpLElvP
mnHa9AMYgdmUVJQJsXnf95ArjeT+EhUUjf4DPR2vLFidjoblgJUTIqHxVAVw51Fc
Yp3s6o+jPvd3PC/fDehMi+3AW5OYqRh5IAO6ooXI+RbkrxJMrPcoj/ibYsvwQC9l
Xt4wW988FiNT5A2pjY9PDdpXBAxqZZ7EylbIbrdpx/GV3p7raeDK5ohuq4GLLw2K
+scOo7iu3WxO0itaGyshhqF17sA+LdsK3z8qQdTZHrHpalyDmLuTLn4niHgrVhUL
oKnLkJAK+4HC2avtCR7t8nSOs8fk9+7fnDY33w8LVPdVO2lsGKpuZh1ZfgX4QD3l
FfjkNvwONrODl851W8T4EKKBYXIhs7/vlFCIx2onczuLp/Lv8b+u3IJNCrOtTU+z
6h00dyOzJySs5ltLyaH/Smoso/CiWE4GCrh7AUdfnQ3iXthO16Hj4S+EdoXbOPZ/
mSnJCGaNeXvAvqKcfYrzpwDUmcaV/PeUu5gOt4kmhnqiAfcy4kI5hAYNFgJad16t
/5Xqr1RtijszJkvKR9miwKfeexnstIGOr5cKwZV4aOmSsAVAfywzG/X3u9E87XpA
KAzYoWKsae4bylZ7dJY7+BaDSq3WimXL80Fs8mtAI3VSPZ6ppK4RBQkHpuHC9//1
tY58qBR3w4G/ZTBXdYAqLRWpjrcmUmAH5ZHV5DkL9WCHZq/iSwCSoqILSzOVlbQK
Ihi4ZugDZwOrGRKUTk7gZk/T8FQP+5BPi5hipBGDwmkhKX1TuPTVQEAYg3A799qU
30Hf7Fg4VWQ8mTdBl0zI8/Z7mF2hfLSkqBHs4i2YfR3PvuqaBo5UVwgSRY4SCSn7
C0cwybR+Y1qG5bz218KutspVwPxSg9LD3O3MjvL7FwEymXLz6E/nBVS6oCaqwCK7
ZEg0qsOrBWa+f2scas52B4oQUT1qdU5qGiXf5tzimMgC1Xu9IfjDmfp11gJZUn1V
CzAEqAQ6jnmKbRo3huYpeMzloMn54QeId3SQtgXhYrr4l1feMQC16XZpWflc4Uae
xM06W1XHJgz3EaU+FcFIZ9/tymUcIdJz0AGLx21xADSmsCQQlTBILjNVrlK9E6ws
D6sAAXiWEZaeFvuEMwNDq0oIkMsXqbHiBlh+sQbzirYv/EEzlFo1fhns6AaSXxhN
5vmqIrk4vgIfi+q2MNAwBroIon0T2DsB8li07clHciEq+rY+07VPHIcdFBSPLM69
REvMpQF77G0Cs8UC1IClzYs354udg8z8BsztVbq0yBOw1C1R775kz0NHtquNcUcK
pJvoHPLdPIV8xaXscwrySTFJ0Y9PwKPtE2rN1N7g7cx+adrlYF+yILs1+XOtMQ9G
3xMiXm8ZukKPJTF0I0qyufUsPmCRn6QXf0W89Ke7WSpNZaGAHlSyZfwy15fn671V
94+eNqgZVvUYUKbsMwICRgVrpO+YMryYNrGpUjvDojfyQJtPUg8jL6in1b1XBQ9Z
YhISycZYkaNnfhLgRMPamXv0Ww8tHEPrS9k9tvjW4rh3/8cQriIjKsI5iKTeciAQ
i4lOzklxWC3ztrW65PNvtLMvXzIgqkK6T42O6/anZ0dZAL7CaQ5wuNHXWiMoZFhW
dAvBPjsCOhdjsKQknFmFFWp/UaEsb4epA5S5fRi6pzMEEUMqh+KC5mDd0YElktaJ
fB4np1SuubuhTdr0OU0NlY6EyjwBiHCIyDCAyw6sTq+3uj8c6slAYK620YNbikWM
rv9TGk2DxCLtk4tQhqnWeP4CYdHd8sW0q5U3GkXHeKTt2GQuBoB/dVLj4gsLD/BN
wv7MdGZcVvAt3ZA5NgFRbMV2OB8nWY9672cSraF/7COrTFWllq00wvvsuXH9vtym
hRULrl8Km5DtEyWiP6T/qJVpMirSnlw0K7BvZP/GQzs75efU9hOzQYdC2iQvWy9M
ZbDrPL02Vah2dO9fNHPxBcsLlzuh2kw/kvYFbCVj8duNa9c9cy+5t3zbJMAnuqB6
H8OPgHGj6GQrtRYWGjo6nuXSuANlBEKt09FUSDFmMHuvLUrwoUDRlWWJIUCjfxTZ
m8zKVkDfPsLxVknO1cF3X6GP6TtWNiCbH67g1MqcwLU3f3w1EaNbQA4ud0t9oqCA
JGqqczuJPZRVfsy6AAzDQe3VArQuxYVCprCtbKYNXFEHDjDOv03UlhIkyHDskYzx
JG6QIM6KU3XrFA6cNmscm+nCnhmLWzqSMLKcIMap+7JoEGiECGdLA0YXJMYURuNJ
c3axZtpBXWY6WTwqvCMXYLNLsJF2HbcsLaMJpuakrbxyRdXNOrj0Gk13FbmL9V4o
w8N5LIpcOlcRpgkcUbP6yIWGP4bC55kTryrPw+XeC2si8q+qPeKKKgmusyz7EWWO
EcpYU+Oc/4x3VQLJnWBvAf1aXmw33uUg0UDVwtOv3D4uyuX5MiMdnXrblHdrqoPu
jzWTEDrHrcQwuSd1thiFqJJzfkz12a2Dk8ewEwTYmnV7oov94RT0Bh+EKX0iOWpt
8/nzXVgerK9+tyipL2eAvAZkfi1LPFc4vlJzBHgiMW1UxVc68cPqOYJvSdBSG2Kg
aNic2eZCu9c7M4VZnA2tclrc1IPaVN4Dk31ST20ZdSi1x12sk14A7HevJFAlT3H0
iwEmNYEqT+uOb3YhedOCmuj4npCHhxzPwPl6IfcHTn5M2P2RpforYUCUXipNarrZ
h5MvxJBH0e0kpmCQmH0J44DlxUPTRefWVIyGT4Tf50SmktCqCFxGMQMWPQSIl585
2e/18HjImIbXuRzflE5aHZ4O7JJqLS8wpW6539IhalrjAauAdrAzwhYcwjEpZsUm
hB0BKO6ocE5iA7tSyeaD//92IOdaAyF6zOZ4s0dmE2OD3Y9fD+6LxCofZXhLOcP9
Kc1oZPgWvvosopK8+MHyWHIVQuoquSOg7O7Fy5y2S2HWom19MHYVGws7f94Y5bH+
DzaZZaFcjWrXQ65HshNF0f2kMKiGqPeSS36c1IpsgT1eMnBtQoBY6hYU5fBYPEbV
GBpP+qxmSQMcH6umG4RE9JkZZMTmlZx93CO/y3euMyqY25k/VqvJ6FoJbvUpgpkR
PQ6fECv9t0s91jw9CRnWPkTIvgjof6vUfZj2uXSkJ7UNYz2wAEheN3VSoqk0oakM
Pq2LgVU1fQKWaG6cO5gOokgKdz1mpbpnfV/Ecfb5NN/paY4scg41L4DUUdycdR3y
II8hahrFCW0QIG1jGcLVOKgUNnxsw3R5PsXxjnFJh/a2AW+B9YIFwVn3tPEayRls
mCxB+7tUwmsCvxpoJ5et9wbH7q0UkNTCKKftLuz3dIP/jyqtPjCwPuLy8yHtcG0x
FOn2D5IrneDB6M2YqnVAvuyHGFBHo8LdBAIB3okt/7vxkM9+Cy41En/s/kQCumUZ
e4A2bNlqzunUFCjseE5hE0aHuG92oWKQe7VL/TXVrgDYHfG1Fyk8wOIJ4/Sq5y6Y
kDvSR5kCu+tDm0CNj//88RuXM0WiwkEbdofx6v2Nl21i/kYvjDh1yJEvNtvEsBOb
atswN/7Hy0/jDPQf39n5nzHCdSnd8p8C3MUL6PT84datV5z5jXm3tIDWD/skV72K
x7eapht5ykZjaesu7SVQuRbbHOlZKE19IRZwP9jsPXK71ROaxmHT+NVZ/WrDER/N
FPrue6g9+CCVd4tzQaLjORyKDEecIaEyzUKiMi9HBtAkT+3JH74D9nHEk2neE20m
Limgp4upLEDyz8DZQ8J357lqdM5i2Z126f2u+4Uqdqz3wmQeIhpf8Yxl5mcd9ufJ
ZINbwYXmQsuSMWy0j0k+O4IUO/pI83zFEEfvsnzEhH5NSnVWDwEXLmB5X1Cpzl48
erkAI6cnff39yzIlI0pU+LWv9TSnvhNqHIz5IM5/CuaFV+X6yJXjKOoh17YmaYEn
/Bed/3+3CmptS0bAjOhfHStCaxhuQ2cyJOF/7kyyz33+fc/fUI9PKk56QU+g9tGo
La/ZWTt49Ce/fkTVABM2Ycor1yTGlIv/moN0TgeOV9GRiSkgxtOWF8GZsLKNFbYp
P0j0jdcUoUaJw3memC/tazQnwIycVv6fUvxnMRSi2X3uEaKcwVVAEPV94uy3WTE5
IvjJlCTIda7vZF1r3ZElbSMLp+BCgFf1gtE2zOGturQJDyvgYhvlmz6r8pe7YM0K
YKigJOU6ktS5js63Z7UIv8qourekZhYOvs6sfeLjlkEom4JoJ0U+5mmjUuWUj0Dr
w6tLKaUAkxh62g9ef9Six7hk12EZj1sJmh337W8j+DplErCrgwg/rDU+fdZPP5rq
mZv22+LaNSdeyD8a8c6V+VS5tlHUvU/nH6Rwre+pZ1MayHtRgQ5M5vP30g68ikRB
ebo99YCGT+6ElM8j/lCYRdzgiiMQY+eiSuw838B5Rztts5ANQFd1OUb5sC7stZts
YywreHImxCHaKVG/kow+aDjPgSzzk/J3V3Ne5pzhnDPFExpAN3bXT0j3Beg9WhrX
DtAbGWgff7vXMENRd/Q7hHKawo/gxqgIUtXqb8G2IEn4iLw2YmDm5lK+agZ7A07n
oRq05q/9JDyIjYM/cm1qhNUYMLAOKXuJc4oCTd8q4vJryURFeoSzCJNlwoBmktIf
brYY3iOUG///+M4zgb9KOqmPdUwq+28R5xqzunQEsu/53PgeAx1yu9PurljPYUxE
PrQ0HHQ2I4/kdpgtNgztFmU7ao2HROSdxNfkCs1ivmwJpiW+rpwpJAThcAqkImYg
A3dyojiZEOLs8uuUox4cEXpQRfomxlkb2hU5NNH3HHwkAR1hZdN7bRJGnmyhm2AL
sR6xmKIRTxjxYyKf2/HnueGfQ7IH+l8QeKLVpyNMN+UVEm1lxAPNHqZ5hvdqMDvc
h8qXEoFzwL9Ww9EHqdKZInSo1bbm38uoewgVx87WFQdalBzt7MDziJ9JH4hmYS4i
D5ndrSIR6KlnR8g0SnCKPTYTRXNSLgkk4ezqwmtBIaIS67SJ12fSmXnBnT1ZqsPs
LK2r87eXyjVkw0MnmmkjIDJJtYHGnJROU7roDbEAzdeqYtuixZlSwNlOKIEUGji3
Y1cFie7JW++N8BnGSp8tSUsoKjf/pvJdrv0W2LJYOnuSVKhgw8zujYiy6jTCW4x3
F0jQuVDJOYKIFVDs7pv0iOXaBKC8JzxnCTyPiONpbeP5M8XzRSC4KLDKRT0dwVJ4
QiMkd20MuZrXqrWdpq0PegowwIRkTu9r8tJBPvsYx/ArKaIl4AFGyjicQmc6xUSS
r9+Gdm0Z6m/Un3M4Sf57MES46nkHjKgc9Y6hdAXtgp6PEarVMHZmP11dk3ZL8eZp
ZdNQ3k7ssuNB6KOwdiyfARr83gqDYbjxSdin6jdMNNXlG2Wn2p9phPQzz8521Ydx
5l5pWEMQd3sl0dN/HsJM5wJzVsAg3Vu8abuB3FpS5Kcjg3jkPA0nHaCYvlXv+RKC
Ox01YWM+8gfEKf/IHdNyBOvvTz4g3ppTH6LjGUN3obvQEiMwESpo9hl73Crcrwou
E3FLJuQzwlXmjAiBAdvYQk3oDanZWWyGno+blACTC/5XhbRmcLviU6fPwnNvv/Pd
5yS2xpMYtkewul/KaeF8QXoaeHr6IAsXjz5FQ/Sw7xE7gXslMaAa+XJgGOrTT0pp
2T9Sz2h6U3HQk450kCsmH76vaJxfApVSBXBAoAA5j3a7al/BXPV4JiBCaliw1qBd
Ih3/hGJLzQnSgUOMEy1C3QYJiWiloxEZkvV5LxvFfini0G8uVwNRVp1SF7z58bP+
p6mEanl9lcWADOJes8EbiQ50RTpdEZKH36AF52CbY/Yr6p9K3CKHGdOb4B5SpayX
dv80fCFjK7yuBxK9wNTfOQsVQQH2n2FBxaMLMf//MRVDiC1K7jncqXcuG0ffDmdD
Y0x4wQG4+LopEBoGzlFsIBpRM7PSL75lb/DCwemvMdbFRyvO1320ZcPUGIYTNz0/
cRJhXzHrQoIOtm534epWN5CzWHpRbmsxmVEwMSzpxlF7TTnWFw4EmPLRHgtr54aW
sfPIiVPPm8lGeAObx1RNjGm2CEi+a0CAa2c5NXzvDZv5+myf1uQKzZqJA8REMyfk
Ik5q24qpxPWr38wRuw/czOEDQo29uMj04bMBrxIvMgqQP7veyc/9QwJ5XYOricnT
e0IwSi/utOlvXvmb1YdPXGebS78wNZcpN4RAYux+Zti6CdfVM4+yfrpTuh9vdLf8
2HXcUqeKq2D06+x7BKs3GYccWcGUix9UPtKEraFWOQZMSyuk641Uiak8X81hp/Gb
cEPB4gOUAfCGNdv8e55aQuCaNQTjk4ZEDRAzk0WaVBfYiMZ4gpCnVoQyD8HhcxBF
uJc0s4bemOBT3OBrZyVq2U4GOy9xOYa3juBDHob5U7WNnyNkDmO+xjxWydAKJNVj
7KX8KlFuCFhw3tqUA6iMJsad00+/VMTchSdzorRRKQD5rPST3TM1AhVQM3phWISi
gE2ZKNU7jyx6f5zjkwK9QeX74KbcM1d869h0Ha7yXJUukAzNDYmdwNJgWnBWhIfx
24fP1/Cat21jyDk4ivLVn97iJ4eSDqd++ZM04dyOZHxoOn9/xAjH5VVnkCCFeED4
eEXRJCUOpGA1Y5h51Y7g0M8pST6eY5piJ03J/mDimoX+/IvFM+wMP0pnvrPzjwQ9
lUkd2wk72sYFjHtf99vGg+ROcn3qn8xo3y4hzeHiG3AdFnVX2pm8mRCiPzJKu8S7
/vEkfqm7wqYSwU4A3VSEAqB4n3WeT4uu5EminEQLu+hxcqRd+vB7TYrmHWquXUcl
y3GZIVa9dZDxYdFpmeBKOYvi48fJWDTJdKyxhz08iLFXBOFtSDpJkkxkZ4p1az7+
JRexY8rA4t6yHt6FOqDgljWAZ50YMjpnhoo+z0j82G8=
`protect end_protected
