localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_CMAP_CHK = {
  {32'hbce46269, 32'h00000000} /* (15, 15, 15) {real, imag} */,
  {32'hbdfb6981, 32'h00000000} /* (15, 15, 14) {real, imag} */,
  {32'hbb861256, 32'h00000000} /* (15, 15, 13) {real, imag} */,
  {32'h3d807083, 32'h00000000} /* (15, 15, 12) {real, imag} */,
  {32'h3dd4b771, 32'h00000000} /* (15, 15, 11) {real, imag} */,
  {32'h3dfd286a, 32'h00000000} /* (15, 15, 10) {real, imag} */,
  {32'hbcb8f23e, 32'h00000000} /* (15, 15, 9) {real, imag} */,
  {32'hbe0b4707, 32'h00000000} /* (15, 15, 8) {real, imag} */,
  {32'hbd0b3b94, 32'h00000000} /* (15, 15, 7) {real, imag} */,
  {32'hbd9b5eb7, 32'h00000000} /* (15, 15, 6) {real, imag} */,
  {32'hbeaa401f, 32'h00000000} /* (15, 15, 5) {real, imag} */,
  {32'hbe8b4706, 32'h00000000} /* (15, 15, 4) {real, imag} */,
  {32'hbe8e6eff, 32'h00000000} /* (15, 15, 3) {real, imag} */,
  {32'hbea6f2dc, 32'h00000000} /* (15, 15, 2) {real, imag} */,
  {32'hbe7d0728, 32'h00000000} /* (15, 15, 1) {real, imag} */,
  {32'hbe095a14, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hbded86a8, 32'h00000000} /* (15, 14, 15) {real, imag} */,
  {32'hbeb3fc5c, 32'h00000000} /* (15, 14, 14) {real, imag} */,
  {32'hbe165327, 32'h00000000} /* (15, 14, 13) {real, imag} */,
  {32'h3cadd258, 32'h00000000} /* (15, 14, 12) {real, imag} */,
  {32'h3e4b9e78, 32'h00000000} /* (15, 14, 11) {real, imag} */,
  {32'h3e3954b3, 32'h00000000} /* (15, 14, 10) {real, imag} */,
  {32'h3d9414d9, 32'h00000000} /* (15, 14, 9) {real, imag} */,
  {32'h3df13ada, 32'h00000000} /* (15, 14, 8) {real, imag} */,
  {32'h3d8b5772, 32'h00000000} /* (15, 14, 7) {real, imag} */,
  {32'hbd70fe3d, 32'h00000000} /* (15, 14, 6) {real, imag} */,
  {32'hbee006ab, 32'h00000000} /* (15, 14, 5) {real, imag} */,
  {32'hbe1dc603, 32'h00000000} /* (15, 14, 4) {real, imag} */,
  {32'hbe4671a7, 32'h00000000} /* (15, 14, 3) {real, imag} */,
  {32'hbe369692, 32'h00000000} /* (15, 14, 2) {real, imag} */,
  {32'hbdc84929, 32'h00000000} /* (15, 14, 1) {real, imag} */,
  {32'hbe096e58, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'h3deebc4b, 32'h00000000} /* (15, 13, 15) {real, imag} */,
  {32'h3d695cd6, 32'h00000000} /* (15, 13, 14) {real, imag} */,
  {32'hbe59e528, 32'h00000000} /* (15, 13, 13) {real, imag} */,
  {32'hbea7a4ed, 32'h00000000} /* (15, 13, 12) {real, imag} */,
  {32'hbde6acb2, 32'h00000000} /* (15, 13, 11) {real, imag} */,
  {32'hbda7038e, 32'h00000000} /* (15, 13, 10) {real, imag} */,
  {32'hbe192a92, 32'h00000000} /* (15, 13, 9) {real, imag} */,
  {32'h3e796c7d, 32'h00000000} /* (15, 13, 8) {real, imag} */,
  {32'h3e14be1b, 32'h00000000} /* (15, 13, 7) {real, imag} */,
  {32'h3eb0183e, 32'h00000000} /* (15, 13, 6) {real, imag} */,
  {32'h3dd8e9e8, 32'h00000000} /* (15, 13, 5) {real, imag} */,
  {32'hbd424dee, 32'h00000000} /* (15, 13, 4) {real, imag} */,
  {32'hbe34c92f, 32'h00000000} /* (15, 13, 3) {real, imag} */,
  {32'hbd3317f6, 32'h00000000} /* (15, 13, 2) {real, imag} */,
  {32'h3eca78b1, 32'h00000000} /* (15, 13, 1) {real, imag} */,
  {32'h3ea6edc8, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'h3e49ee2b, 32'h00000000} /* (15, 12, 15) {real, imag} */,
  {32'h3e985631, 32'h00000000} /* (15, 12, 14) {real, imag} */,
  {32'hbd766624, 32'h00000000} /* (15, 12, 13) {real, imag} */,
  {32'hbe68ca24, 32'h00000000} /* (15, 12, 12) {real, imag} */,
  {32'hbec9952f, 32'h00000000} /* (15, 12, 11) {real, imag} */,
  {32'hbe79f831, 32'h00000000} /* (15, 12, 10) {real, imag} */,
  {32'hbe13623d, 32'h00000000} /* (15, 12, 9) {real, imag} */,
  {32'hbcc9e37e, 32'h00000000} /* (15, 12, 8) {real, imag} */,
  {32'h3b06d365, 32'h00000000} /* (15, 12, 7) {real, imag} */,
  {32'h3e69496a, 32'h00000000} /* (15, 12, 6) {real, imag} */,
  {32'h3e55b2a3, 32'h00000000} /* (15, 12, 5) {real, imag} */,
  {32'hbe0dabe8, 32'h00000000} /* (15, 12, 4) {real, imag} */,
  {32'hbe715020, 32'h00000000} /* (15, 12, 3) {real, imag} */,
  {32'hbca9a87e, 32'h00000000} /* (15, 12, 2) {real, imag} */,
  {32'h3e79aa57, 32'h00000000} /* (15, 12, 1) {real, imag} */,
  {32'h3dd1a431, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'h3e9a72ff, 32'h00000000} /* (15, 11, 15) {real, imag} */,
  {32'h3ec00c67, 32'h00000000} /* (15, 11, 14) {real, imag} */,
  {32'h3c2f592b, 32'h00000000} /* (15, 11, 13) {real, imag} */,
  {32'hbbe3e1e8, 32'h00000000} /* (15, 11, 12) {real, imag} */,
  {32'hbe681f0e, 32'h00000000} /* (15, 11, 11) {real, imag} */,
  {32'hbe8525f1, 32'h00000000} /* (15, 11, 10) {real, imag} */,
  {32'hbdc24d66, 32'h00000000} /* (15, 11, 9) {real, imag} */,
  {32'h3b70342d, 32'h00000000} /* (15, 11, 8) {real, imag} */,
  {32'h3d98d837, 32'h00000000} /* (15, 11, 7) {real, imag} */,
  {32'h3e65178c, 32'h00000000} /* (15, 11, 6) {real, imag} */,
  {32'h3d5c7be8, 32'h00000000} /* (15, 11, 5) {real, imag} */,
  {32'hbd861ad9, 32'h00000000} /* (15, 11, 4) {real, imag} */,
  {32'hbe0ef347, 32'h00000000} /* (15, 11, 3) {real, imag} */,
  {32'h3d4fb720, 32'h00000000} /* (15, 11, 2) {real, imag} */,
  {32'h3d1402fb, 32'h00000000} /* (15, 11, 1) {real, imag} */,
  {32'hbdb8ca7f, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h3e113cff, 32'h00000000} /* (15, 10, 15) {real, imag} */,
  {32'h3e6a6ee5, 32'h00000000} /* (15, 10, 14) {real, imag} */,
  {32'hbe24aec2, 32'h00000000} /* (15, 10, 13) {real, imag} */,
  {32'hbe22085f, 32'h00000000} /* (15, 10, 12) {real, imag} */,
  {32'h3e363838, 32'h00000000} /* (15, 10, 11) {real, imag} */,
  {32'h3d90a0be, 32'h00000000} /* (15, 10, 10) {real, imag} */,
  {32'hbecd0037, 32'h00000000} /* (15, 10, 9) {real, imag} */,
  {32'hbea0c5e8, 32'h00000000} /* (15, 10, 8) {real, imag} */,
  {32'h3dbb420e, 32'h00000000} /* (15, 10, 7) {real, imag} */,
  {32'h3de1d07f, 32'h00000000} /* (15, 10, 6) {real, imag} */,
  {32'hbe0b564f, 32'h00000000} /* (15, 10, 5) {real, imag} */,
  {32'h3a3141cd, 32'h00000000} /* (15, 10, 4) {real, imag} */,
  {32'hbcf08c53, 32'h00000000} /* (15, 10, 3) {real, imag} */,
  {32'h3d690d0a, 32'h00000000} /* (15, 10, 2) {real, imag} */,
  {32'h3da0b139, 32'h00000000} /* (15, 10, 1) {real, imag} */,
  {32'h3d494b19, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'hbe48a40c, 32'h00000000} /* (15, 9, 15) {real, imag} */,
  {32'hbf087e47, 32'h00000000} /* (15, 9, 14) {real, imag} */,
  {32'hbe402a01, 32'h00000000} /* (15, 9, 13) {real, imag} */,
  {32'hbd381444, 32'h00000000} /* (15, 9, 12) {real, imag} */,
  {32'h3e25da1d, 32'h00000000} /* (15, 9, 11) {real, imag} */,
  {32'h3e04379b, 32'h00000000} /* (15, 9, 10) {real, imag} */,
  {32'hbf28f123, 32'h00000000} /* (15, 9, 9) {real, imag} */,
  {32'hbf06efa4, 32'h00000000} /* (15, 9, 8) {real, imag} */,
  {32'hbdb28e34, 32'h00000000} /* (15, 9, 7) {real, imag} */,
  {32'hbe0bf314, 32'h00000000} /* (15, 9, 6) {real, imag} */,
  {32'hbea0923f, 32'h00000000} /* (15, 9, 5) {real, imag} */,
  {32'hbdf8eefc, 32'h00000000} /* (15, 9, 4) {real, imag} */,
  {32'h3d95d3c5, 32'h00000000} /* (15, 9, 3) {real, imag} */,
  {32'h3da8355f, 32'h00000000} /* (15, 9, 2) {real, imag} */,
  {32'h3d6c7114, 32'h00000000} /* (15, 9, 1) {real, imag} */,
  {32'h3de0aff7, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'hbe294563, 32'h00000000} /* (15, 8, 15) {real, imag} */,
  {32'hbf076196, 32'h00000000} /* (15, 8, 14) {real, imag} */,
  {32'hbe75524d, 32'h00000000} /* (15, 8, 13) {real, imag} */,
  {32'hbe7c895b, 32'h00000000} /* (15, 8, 12) {real, imag} */,
  {32'hbdfc93e3, 32'h00000000} /* (15, 8, 11) {real, imag} */,
  {32'h3dcb8d16, 32'h00000000} /* (15, 8, 10) {real, imag} */,
  {32'hbe7f2f2b, 32'h00000000} /* (15, 8, 9) {real, imag} */,
  {32'hbf148a77, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'hbead3ef4, 32'h00000000} /* (15, 8, 7) {real, imag} */,
  {32'hbe57a645, 32'h00000000} /* (15, 8, 6) {real, imag} */,
  {32'hbe0beffd, 32'h00000000} /* (15, 8, 5) {real, imag} */,
  {32'h3df762fa, 32'h00000000} /* (15, 8, 4) {real, imag} */,
  {32'h3e4233c9, 32'h00000000} /* (15, 8, 3) {real, imag} */,
  {32'h3dd168f8, 32'h00000000} /* (15, 8, 2) {real, imag} */,
  {32'h3d0f79cd, 32'h00000000} /* (15, 8, 1) {real, imag} */,
  {32'hbd3a7299, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h3d7ed8c7, 32'h00000000} /* (15, 7, 15) {real, imag} */,
  {32'hbd2e9c41, 32'h00000000} /* (15, 7, 14) {real, imag} */,
  {32'hbe8b48ce, 32'h00000000} /* (15, 7, 13) {real, imag} */,
  {32'hbef84f68, 32'h00000000} /* (15, 7, 12) {real, imag} */,
  {32'hbef83438, 32'h00000000} /* (15, 7, 11) {real, imag} */,
  {32'hbdb3064f, 32'h00000000} /* (15, 7, 10) {real, imag} */,
  {32'hbce6b2f5, 32'h00000000} /* (15, 7, 9) {real, imag} */,
  {32'hbe8eb982, 32'h00000000} /* (15, 7, 8) {real, imag} */,
  {32'hbc8c9ff8, 32'h00000000} /* (15, 7, 7) {real, imag} */,
  {32'h3e591e09, 32'h00000000} /* (15, 7, 6) {real, imag} */,
  {32'h3da4aa93, 32'h00000000} /* (15, 7, 5) {real, imag} */,
  {32'h3e1e0e2d, 32'h00000000} /* (15, 7, 4) {real, imag} */,
  {32'hbcd9136b, 32'h00000000} /* (15, 7, 3) {real, imag} */,
  {32'hbe841f96, 32'h00000000} /* (15, 7, 2) {real, imag} */,
  {32'hbe8196b0, 32'h00000000} /* (15, 7, 1) {real, imag} */,
  {32'hbd60ce36, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'hbd741e97, 32'h00000000} /* (15, 6, 15) {real, imag} */,
  {32'hbd3af67a, 32'h00000000} /* (15, 6, 14) {real, imag} */,
  {32'hbea6a143, 32'h00000000} /* (15, 6, 13) {real, imag} */,
  {32'hbd88d71b, 32'h00000000} /* (15, 6, 12) {real, imag} */,
  {32'hbdcfc947, 32'h00000000} /* (15, 6, 11) {real, imag} */,
  {32'h3d49bf31, 32'h00000000} /* (15, 6, 10) {real, imag} */,
  {32'h3e47e2ab, 32'h00000000} /* (15, 6, 9) {real, imag} */,
  {32'h3d091f66, 32'h00000000} /* (15, 6, 8) {real, imag} */,
  {32'h3e6804ab, 32'h00000000} /* (15, 6, 7) {real, imag} */,
  {32'h3e7f4b3a, 32'h00000000} /* (15, 6, 6) {real, imag} */,
  {32'hbd02696c, 32'h00000000} /* (15, 6, 5) {real, imag} */,
  {32'h3cf4675d, 32'h00000000} /* (15, 6, 4) {real, imag} */,
  {32'hbdbe893c, 32'h00000000} /* (15, 6, 3) {real, imag} */,
  {32'hbef37f9e, 32'h00000000} /* (15, 6, 2) {real, imag} */,
  {32'hbeae9a6a, 32'h00000000} /* (15, 6, 1) {real, imag} */,
  {32'hbd480751, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h3da9cfce, 32'h00000000} /* (15, 5, 15) {real, imag} */,
  {32'h3e252081, 32'h00000000} /* (15, 5, 14) {real, imag} */,
  {32'hbe2fe318, 32'h00000000} /* (15, 5, 13) {real, imag} */,
  {32'h3d0543d3, 32'h00000000} /* (15, 5, 12) {real, imag} */,
  {32'hbd84cfe8, 32'h00000000} /* (15, 5, 11) {real, imag} */,
  {32'hbd9e5547, 32'h00000000} /* (15, 5, 10) {real, imag} */,
  {32'hbd10b8b7, 32'h00000000} /* (15, 5, 9) {real, imag} */,
  {32'hbd67b18e, 32'h00000000} /* (15, 5, 8) {real, imag} */,
  {32'hbc951ae0, 32'h00000000} /* (15, 5, 7) {real, imag} */,
  {32'hbc5682a7, 32'h00000000} /* (15, 5, 6) {real, imag} */,
  {32'hbe58df6f, 32'h00000000} /* (15, 5, 5) {real, imag} */,
  {32'hbdda123d, 32'h00000000} /* (15, 5, 4) {real, imag} */,
  {32'h3b63c4f3, 32'h00000000} /* (15, 5, 3) {real, imag} */,
  {32'h3e7d5dda, 32'h00000000} /* (15, 5, 2) {real, imag} */,
  {32'h3e513715, 32'h00000000} /* (15, 5, 1) {real, imag} */,
  {32'hbd06bba0, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'hbcddc748, 32'h00000000} /* (15, 4, 15) {real, imag} */,
  {32'hbd5be1e3, 32'h00000000} /* (15, 4, 14) {real, imag} */,
  {32'hbec295e0, 32'h00000000} /* (15, 4, 13) {real, imag} */,
  {32'hbdbe0c1c, 32'h00000000} /* (15, 4, 12) {real, imag} */,
  {32'hbe789549, 32'h00000000} /* (15, 4, 11) {real, imag} */,
  {32'hbc718703, 32'h00000000} /* (15, 4, 10) {real, imag} */,
  {32'hbe434932, 32'h00000000} /* (15, 4, 9) {real, imag} */,
  {32'hbd4d414c, 32'h00000000} /* (15, 4, 8) {real, imag} */,
  {32'hbd59ad26, 32'h00000000} /* (15, 4, 7) {real, imag} */,
  {32'h3c59c0a0, 32'h00000000} /* (15, 4, 6) {real, imag} */,
  {32'hbe80fd57, 32'h00000000} /* (15, 4, 5) {real, imag} */,
  {32'h3de97580, 32'h00000000} /* (15, 4, 4) {real, imag} */,
  {32'h3e1fd470, 32'h00000000} /* (15, 4, 3) {real, imag} */,
  {32'h3e2f89c8, 32'h00000000} /* (15, 4, 2) {real, imag} */,
  {32'hbd9c1d4b, 32'h00000000} /* (15, 4, 1) {real, imag} */,
  {32'hbe2cd5de, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'hbdcb29be, 32'h00000000} /* (15, 3, 15) {real, imag} */,
  {32'h3c0095b8, 32'h00000000} /* (15, 3, 14) {real, imag} */,
  {32'h3c91d6fc, 32'h00000000} /* (15, 3, 13) {real, imag} */,
  {32'h3d4f9272, 32'h00000000} /* (15, 3, 12) {real, imag} */,
  {32'hbd276a5e, 32'h00000000} /* (15, 3, 11) {real, imag} */,
  {32'h3e66024d, 32'h00000000} /* (15, 3, 10) {real, imag} */,
  {32'hbc12f276, 32'h00000000} /* (15, 3, 9) {real, imag} */,
  {32'hbd010bad, 32'h00000000} /* (15, 3, 8) {real, imag} */,
  {32'hbdb9ea9c, 32'h00000000} /* (15, 3, 7) {real, imag} */,
  {32'h3e162d81, 32'h00000000} /* (15, 3, 6) {real, imag} */,
  {32'hbe11e93c, 32'h00000000} /* (15, 3, 5) {real, imag} */,
  {32'hbad268a8, 32'h00000000} /* (15, 3, 4) {real, imag} */,
  {32'h3e305326, 32'h00000000} /* (15, 3, 3) {real, imag} */,
  {32'hbe085116, 32'h00000000} /* (15, 3, 2) {real, imag} */,
  {32'hbe150ce7, 32'h00000000} /* (15, 3, 1) {real, imag} */,
  {32'h3e889ca1, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'h3d1aa218, 32'h00000000} /* (15, 2, 15) {real, imag} */,
  {32'h3c0e5808, 32'h00000000} /* (15, 2, 14) {real, imag} */,
  {32'h3e98ebbc, 32'h00000000} /* (15, 2, 13) {real, imag} */,
  {32'h3e236938, 32'h00000000} /* (15, 2, 12) {real, imag} */,
  {32'hbe02171e, 32'h00000000} /* (15, 2, 11) {real, imag} */,
  {32'h3e359276, 32'h00000000} /* (15, 2, 10) {real, imag} */,
  {32'h3e383959, 32'h00000000} /* (15, 2, 9) {real, imag} */,
  {32'h3e18b597, 32'h00000000} /* (15, 2, 8) {real, imag} */,
  {32'hbe26ec46, 32'h00000000} /* (15, 2, 7) {real, imag} */,
  {32'hbedcc37b, 32'h00000000} /* (15, 2, 6) {real, imag} */,
  {32'hbe9d151e, 32'h00000000} /* (15, 2, 5) {real, imag} */,
  {32'hbe2a01eb, 32'h00000000} /* (15, 2, 4) {real, imag} */,
  {32'hbe131115, 32'h00000000} /* (15, 2, 3) {real, imag} */,
  {32'hbebab336, 32'h00000000} /* (15, 2, 2) {real, imag} */,
  {32'hbeb38fd3, 32'h00000000} /* (15, 2, 1) {real, imag} */,
  {32'h3e5c737b, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'hbd7de194, 32'h00000000} /* (15, 1, 15) {real, imag} */,
  {32'hbe6b4093, 32'h00000000} /* (15, 1, 14) {real, imag} */,
  {32'hbe0e5da0, 32'h00000000} /* (15, 1, 13) {real, imag} */,
  {32'h3da56838, 32'h00000000} /* (15, 1, 12) {real, imag} */,
  {32'hbd566d40, 32'h00000000} /* (15, 1, 11) {real, imag} */,
  {32'h3dbfe2ab, 32'h00000000} /* (15, 1, 10) {real, imag} */,
  {32'h3ecb5130, 32'h00000000} /* (15, 1, 9) {real, imag} */,
  {32'h3e3e27ac, 32'h00000000} /* (15, 1, 8) {real, imag} */,
  {32'hbea1aa72, 32'h00000000} /* (15, 1, 7) {real, imag} */,
  {32'hbf22cb5e, 32'h00000000} /* (15, 1, 6) {real, imag} */,
  {32'hbf27d8d8, 32'h00000000} /* (15, 1, 5) {real, imag} */,
  {32'hbea86ca3, 32'h00000000} /* (15, 1, 4) {real, imag} */,
  {32'hbe378011, 32'h00000000} /* (15, 1, 3) {real, imag} */,
  {32'hbdc85e5a, 32'h00000000} /* (15, 1, 2) {real, imag} */,
  {32'hbe849e56, 32'h00000000} /* (15, 1, 1) {real, imag} */,
  {32'hbdf1a715, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'hbc1185ee, 32'h00000000} /* (15, 0, 15) {real, imag} */,
  {32'hbcf6b707, 32'h00000000} /* (15, 0, 14) {real, imag} */,
  {32'hbe32a237, 32'h00000000} /* (15, 0, 13) {real, imag} */,
  {32'h3ba7ca13, 32'h00000000} /* (15, 0, 12) {real, imag} */,
  {32'h3c288227, 32'h00000000} /* (15, 0, 11) {real, imag} */,
  {32'hbddae4a6, 32'h00000000} /* (15, 0, 10) {real, imag} */,
  {32'h3bb2658d, 32'h00000000} /* (15, 0, 9) {real, imag} */,
  {32'hbc625fda, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'hbe26e1b7, 32'h00000000} /* (15, 0, 7) {real, imag} */,
  {32'hbe1073a8, 32'h00000000} /* (15, 0, 6) {real, imag} */,
  {32'hbe5ec9b3, 32'h00000000} /* (15, 0, 5) {real, imag} */,
  {32'hbd8b7b04, 32'h00000000} /* (15, 0, 4) {real, imag} */,
  {32'h39afa704, 32'h00000000} /* (15, 0, 3) {real, imag} */,
  {32'h3b7c0699, 32'h00000000} /* (15, 0, 2) {real, imag} */,
  {32'hbd4a9fb6, 32'h00000000} /* (15, 0, 1) {real, imag} */,
  {32'hbcc0e65a, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h3dc8d762, 32'h00000000} /* (14, 15, 15) {real, imag} */,
  {32'hbe7a11bf, 32'h00000000} /* (14, 15, 14) {real, imag} */,
  {32'hbc8e6ac9, 32'h00000000} /* (14, 15, 13) {real, imag} */,
  {32'h3dcf93e5, 32'h00000000} /* (14, 15, 12) {real, imag} */,
  {32'h3de17fbb, 32'h00000000} /* (14, 15, 11) {real, imag} */,
  {32'hbe9dee7a, 32'h00000000} /* (14, 15, 10) {real, imag} */,
  {32'hbee65715, 32'h00000000} /* (14, 15, 9) {real, imag} */,
  {32'hbe8794b8, 32'h00000000} /* (14, 15, 8) {real, imag} */,
  {32'hbda6ff6d, 32'h00000000} /* (14, 15, 7) {real, imag} */,
  {32'h3d484b7c, 32'h00000000} /* (14, 15, 6) {real, imag} */,
  {32'h3e305122, 32'h00000000} /* (14, 15, 5) {real, imag} */,
  {32'hbd8e5ea5, 32'h00000000} /* (14, 15, 4) {real, imag} */,
  {32'hbe39eacb, 32'h00000000} /* (14, 15, 3) {real, imag} */,
  {32'hbe4ea1e0, 32'h00000000} /* (14, 15, 2) {real, imag} */,
  {32'hbefe9520, 32'h00000000} /* (14, 15, 1) {real, imag} */,
  {32'hbd91d48a, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'h3d0059f8, 32'h00000000} /* (14, 14, 15) {real, imag} */,
  {32'hbecee0fa, 32'h00000000} /* (14, 14, 14) {real, imag} */,
  {32'hbe358731, 32'h00000000} /* (14, 14, 13) {real, imag} */,
  {32'hbe13cdb2, 32'h00000000} /* (14, 14, 12) {real, imag} */,
  {32'h3e6fc42e, 32'h00000000} /* (14, 14, 11) {real, imag} */,
  {32'h3dea1845, 32'h00000000} /* (14, 14, 10) {real, imag} */,
  {32'hbe8732bc, 32'h00000000} /* (14, 14, 9) {real, imag} */,
  {32'hbe453b31, 32'h00000000} /* (14, 14, 8) {real, imag} */,
  {32'h3e2a66a9, 32'h00000000} /* (14, 14, 7) {real, imag} */,
  {32'h3d73b144, 32'h00000000} /* (14, 14, 6) {real, imag} */,
  {32'hbe65099a, 32'h00000000} /* (14, 14, 5) {real, imag} */,
  {32'hbdaa20cb, 32'h00000000} /* (14, 14, 4) {real, imag} */,
  {32'hbe823d2a, 32'h00000000} /* (14, 14, 3) {real, imag} */,
  {32'hbefb05d8, 32'h00000000} /* (14, 14, 2) {real, imag} */,
  {32'hbf09e590, 32'h00000000} /* (14, 14, 1) {real, imag} */,
  {32'hbd148964, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'h3e928be6, 32'h00000000} /* (14, 13, 15) {real, imag} */,
  {32'h3cf92483, 32'h00000000} /* (14, 13, 14) {real, imag} */,
  {32'hbe95253a, 32'h00000000} /* (14, 13, 13) {real, imag} */,
  {32'hbf29bfd9, 32'h00000000} /* (14, 13, 12) {real, imag} */,
  {32'hbeaf6e99, 32'h00000000} /* (14, 13, 11) {real, imag} */,
  {32'h3dc0203d, 32'h00000000} /* (14, 13, 10) {real, imag} */,
  {32'h3ded4dee, 32'h00000000} /* (14, 13, 9) {real, imag} */,
  {32'hbd372dc0, 32'h00000000} /* (14, 13, 8) {real, imag} */,
  {32'hbe2015f8, 32'h00000000} /* (14, 13, 7) {real, imag} */,
  {32'h3e9be68e, 32'h00000000} /* (14, 13, 6) {real, imag} */,
  {32'hbd285edb, 32'h00000000} /* (14, 13, 5) {real, imag} */,
  {32'h3c9fc901, 32'h00000000} /* (14, 13, 4) {real, imag} */,
  {32'hbe4eeabc, 32'h00000000} /* (14, 13, 3) {real, imag} */,
  {32'hbeaaad80, 32'h00000000} /* (14, 13, 2) {real, imag} */,
  {32'h3d7cae76, 32'h00000000} /* (14, 13, 1) {real, imag} */,
  {32'h3ea2d57b, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'h3e22ea8f, 32'h00000000} /* (14, 12, 15) {real, imag} */,
  {32'h3dc3a15c, 32'h00000000} /* (14, 12, 14) {real, imag} */,
  {32'hbd5348d5, 32'h00000000} /* (14, 12, 13) {real, imag} */,
  {32'hbeacd419, 32'h00000000} /* (14, 12, 12) {real, imag} */,
  {32'hbf44172c, 32'h00000000} /* (14, 12, 11) {real, imag} */,
  {32'hbe66dce2, 32'h00000000} /* (14, 12, 10) {real, imag} */,
  {32'hbd7ce55e, 32'h00000000} /* (14, 12, 9) {real, imag} */,
  {32'hbe450668, 32'h00000000} /* (14, 12, 8) {real, imag} */,
  {32'hbedaf207, 32'h00000000} /* (14, 12, 7) {real, imag} */,
  {32'hbe76fb5c, 32'h00000000} /* (14, 12, 6) {real, imag} */,
  {32'hbe06d9bc, 32'h00000000} /* (14, 12, 5) {real, imag} */,
  {32'hbe344380, 32'h00000000} /* (14, 12, 4) {real, imag} */,
  {32'hbe84ea84, 32'h00000000} /* (14, 12, 3) {real, imag} */,
  {32'hbea78323, 32'h00000000} /* (14, 12, 2) {real, imag} */,
  {32'h3e9ede29, 32'h00000000} /* (14, 12, 1) {real, imag} */,
  {32'h3dc5ecc7, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'h3dbd04fe, 32'h00000000} /* (14, 11, 15) {real, imag} */,
  {32'h3eb2a655, 32'h00000000} /* (14, 11, 14) {real, imag} */,
  {32'h3e182e80, 32'h00000000} /* (14, 11, 13) {real, imag} */,
  {32'h3d217b8a, 32'h00000000} /* (14, 11, 12) {real, imag} */,
  {32'hbdd1ee25, 32'h00000000} /* (14, 11, 11) {real, imag} */,
  {32'hbf089bb2, 32'h00000000} /* (14, 11, 10) {real, imag} */,
  {32'hbd9f02df, 32'h00000000} /* (14, 11, 9) {real, imag} */,
  {32'h3e95d17d, 32'h00000000} /* (14, 11, 8) {real, imag} */,
  {32'hbdabd352, 32'h00000000} /* (14, 11, 7) {real, imag} */,
  {32'hbeb166fe, 32'h00000000} /* (14, 11, 6) {real, imag} */,
  {32'hbd65f6e3, 32'h00000000} /* (14, 11, 5) {real, imag} */,
  {32'h3ef0eafa, 32'h00000000} /* (14, 11, 4) {real, imag} */,
  {32'h3e36fe10, 32'h00000000} /* (14, 11, 3) {real, imag} */,
  {32'hbe6ae0ca, 32'h00000000} /* (14, 11, 2) {real, imag} */,
  {32'h3db9fe2a, 32'h00000000} /* (14, 11, 1) {real, imag} */,
  {32'hbe077dd5, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h3d116adc, 32'h00000000} /* (14, 10, 15) {real, imag} */,
  {32'h3ea6c795, 32'h00000000} /* (14, 10, 14) {real, imag} */,
  {32'hbdddbd94, 32'h00000000} /* (14, 10, 13) {real, imag} */,
  {32'hbde90819, 32'h00000000} /* (14, 10, 12) {real, imag} */,
  {32'h3dbae2fb, 32'h00000000} /* (14, 10, 11) {real, imag} */,
  {32'hbeae994e, 32'h00000000} /* (14, 10, 10) {real, imag} */,
  {32'hbede8ed9, 32'h00000000} /* (14, 10, 9) {real, imag} */,
  {32'h3dabf133, 32'h00000000} /* (14, 10, 8) {real, imag} */,
  {32'h3e9544be, 32'h00000000} /* (14, 10, 7) {real, imag} */,
  {32'hbcaa141e, 32'h00000000} /* (14, 10, 6) {real, imag} */,
  {32'h3cdb4a99, 32'h00000000} /* (14, 10, 5) {real, imag} */,
  {32'h3ec25962, 32'h00000000} /* (14, 10, 4) {real, imag} */,
  {32'h3e7068dd, 32'h00000000} /* (14, 10, 3) {real, imag} */,
  {32'hbea1f9bb, 32'h00000000} /* (14, 10, 2) {real, imag} */,
  {32'h3d6a5268, 32'h00000000} /* (14, 10, 1) {real, imag} */,
  {32'h3e8d79b6, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h3bf92921, 32'h00000000} /* (14, 9, 15) {real, imag} */,
  {32'hbe3a0d46, 32'h00000000} /* (14, 9, 14) {real, imag} */,
  {32'hbe5072d6, 32'h00000000} /* (14, 9, 13) {real, imag} */,
  {32'h3eb0442d, 32'h00000000} /* (14, 9, 12) {real, imag} */,
  {32'h3f15885f, 32'h00000000} /* (14, 9, 11) {real, imag} */,
  {32'h3e314f7c, 32'h00000000} /* (14, 9, 10) {real, imag} */,
  {32'hbf6cd44d, 32'h00000000} /* (14, 9, 9) {real, imag} */,
  {32'hbe83ebe5, 32'h00000000} /* (14, 9, 8) {real, imag} */,
  {32'hbe07f4ea, 32'h00000000} /* (14, 9, 7) {real, imag} */,
  {32'hbed419dd, 32'h00000000} /* (14, 9, 6) {real, imag} */,
  {32'h3d5cdd22, 32'h00000000} /* (14, 9, 5) {real, imag} */,
  {32'hbc59ff3d, 32'h00000000} /* (14, 9, 4) {real, imag} */,
  {32'h3d65d8d7, 32'h00000000} /* (14, 9, 3) {real, imag} */,
  {32'hbe77521e, 32'h00000000} /* (14, 9, 2) {real, imag} */,
  {32'hbe6d33d4, 32'h00000000} /* (14, 9, 1) {real, imag} */,
  {32'h3ece2531, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'hbe7a5dbe, 32'h00000000} /* (14, 8, 15) {real, imag} */,
  {32'hbf193cee, 32'h00000000} /* (14, 8, 14) {real, imag} */,
  {32'hbe9b6f0d, 32'h00000000} /* (14, 8, 13) {real, imag} */,
  {32'hbe9c18e0, 32'h00000000} /* (14, 8, 12) {real, imag} */,
  {32'h3ea0bd9a, 32'h00000000} /* (14, 8, 11) {real, imag} */,
  {32'h3ef13759, 32'h00000000} /* (14, 8, 10) {real, imag} */,
  {32'hbe06f704, 32'h00000000} /* (14, 8, 9) {real, imag} */,
  {32'h3d0e3422, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'hbe92cbcf, 32'h00000000} /* (14, 8, 7) {real, imag} */,
  {32'hbeffe8f7, 32'h00000000} /* (14, 8, 6) {real, imag} */,
  {32'h3d80ebe4, 32'h00000000} /* (14, 8, 5) {real, imag} */,
  {32'h3eb69416, 32'h00000000} /* (14, 8, 4) {real, imag} */,
  {32'h3d76e65d, 32'h00000000} /* (14, 8, 3) {real, imag} */,
  {32'hbcd86fa6, 32'h00000000} /* (14, 8, 2) {real, imag} */,
  {32'hbdac8bf7, 32'h00000000} /* (14, 8, 1) {real, imag} */,
  {32'hbdc76d2b, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'hbdb474ed, 32'h00000000} /* (14, 7, 15) {real, imag} */,
  {32'hbeeec781, 32'h00000000} /* (14, 7, 14) {real, imag} */,
  {32'hbf2c1832, 32'h00000000} /* (14, 7, 13) {real, imag} */,
  {32'hbf2e60e0, 32'h00000000} /* (14, 7, 12) {real, imag} */,
  {32'h3dfe74bb, 32'h00000000} /* (14, 7, 11) {real, imag} */,
  {32'h3ecfeb33, 32'h00000000} /* (14, 7, 10) {real, imag} */,
  {32'h3ee81b31, 32'h00000000} /* (14, 7, 9) {real, imag} */,
  {32'h3dafafb5, 32'h00000000} /* (14, 7, 8) {real, imag} */,
  {32'hbde0bbda, 32'h00000000} /* (14, 7, 7) {real, imag} */,
  {32'h3e034fad, 32'h00000000} /* (14, 7, 6) {real, imag} */,
  {32'h3e105ee6, 32'h00000000} /* (14, 7, 5) {real, imag} */,
  {32'hbbfbeefe, 32'h00000000} /* (14, 7, 4) {real, imag} */,
  {32'hbe408b7e, 32'h00000000} /* (14, 7, 3) {real, imag} */,
  {32'hbe58d76c, 32'h00000000} /* (14, 7, 2) {real, imag} */,
  {32'hbdbb6d3c, 32'h00000000} /* (14, 7, 1) {real, imag} */,
  {32'hbe22c186, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'h3d2c1852, 32'h00000000} /* (14, 6, 15) {real, imag} */,
  {32'h3d69d962, 32'h00000000} /* (14, 6, 14) {real, imag} */,
  {32'hbeb4271c, 32'h00000000} /* (14, 6, 13) {real, imag} */,
  {32'h3cad72d9, 32'h00000000} /* (14, 6, 12) {real, imag} */,
  {32'h3f06c84b, 32'h00000000} /* (14, 6, 11) {real, imag} */,
  {32'h3ee9e97a, 32'h00000000} /* (14, 6, 10) {real, imag} */,
  {32'h3f3a9568, 32'h00000000} /* (14, 6, 9) {real, imag} */,
  {32'h3daa758e, 32'h00000000} /* (14, 6, 8) {real, imag} */,
  {32'h3e8090f4, 32'h00000000} /* (14, 6, 7) {real, imag} */,
  {32'h3d3f8771, 32'h00000000} /* (14, 6, 6) {real, imag} */,
  {32'hbeae2427, 32'h00000000} /* (14, 6, 5) {real, imag} */,
  {32'hbe3ac87b, 32'h00000000} /* (14, 6, 4) {real, imag} */,
  {32'h3ded253a, 32'h00000000} /* (14, 6, 3) {real, imag} */,
  {32'hbeadfb83, 32'h00000000} /* (14, 6, 2) {real, imag} */,
  {32'hbd86b22f, 32'h00000000} /* (14, 6, 1) {real, imag} */,
  {32'h3e292b42, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h3df02f43, 32'h00000000} /* (14, 5, 15) {real, imag} */,
  {32'h3ed515b1, 32'h00000000} /* (14, 5, 14) {real, imag} */,
  {32'hbee2afc1, 32'h00000000} /* (14, 5, 13) {real, imag} */,
  {32'hbebda036, 32'h00000000} /* (14, 5, 12) {real, imag} */,
  {32'h3df630e2, 32'h00000000} /* (14, 5, 11) {real, imag} */,
  {32'h3e28558f, 32'h00000000} /* (14, 5, 10) {real, imag} */,
  {32'h3e691651, 32'h00000000} /* (14, 5, 9) {real, imag} */,
  {32'hbdfee465, 32'h00000000} /* (14, 5, 8) {real, imag} */,
  {32'hbdc43a94, 32'h00000000} /* (14, 5, 7) {real, imag} */,
  {32'hbe8a6cc5, 32'h00000000} /* (14, 5, 6) {real, imag} */,
  {32'hbf15a107, 32'h00000000} /* (14, 5, 5) {real, imag} */,
  {32'hbcd71eb2, 32'h00000000} /* (14, 5, 4) {real, imag} */,
  {32'h3e94c3ad, 32'h00000000} /* (14, 5, 3) {real, imag} */,
  {32'h3e048a25, 32'h00000000} /* (14, 5, 2) {real, imag} */,
  {32'h3ef47b5b, 32'h00000000} /* (14, 5, 1) {real, imag} */,
  {32'h3de2fda2, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'hbd4c2fb7, 32'h00000000} /* (14, 4, 15) {real, imag} */,
  {32'hbcf8a124, 32'h00000000} /* (14, 4, 14) {real, imag} */,
  {32'hbeffd8cb, 32'h00000000} /* (14, 4, 13) {real, imag} */,
  {32'hbc8b68b3, 32'h00000000} /* (14, 4, 12) {real, imag} */,
  {32'hbb0cf820, 32'h00000000} /* (14, 4, 11) {real, imag} */,
  {32'h3c54a00a, 32'h00000000} /* (14, 4, 10) {real, imag} */,
  {32'hbb74b384, 32'h00000000} /* (14, 4, 9) {real, imag} */,
  {32'h3e82c7ee, 32'h00000000} /* (14, 4, 8) {real, imag} */,
  {32'hbc1ca770, 32'h00000000} /* (14, 4, 7) {real, imag} */,
  {32'hbe894d09, 32'h00000000} /* (14, 4, 6) {real, imag} */,
  {32'hbf4c5e8b, 32'h00000000} /* (14, 4, 5) {real, imag} */,
  {32'hbe5c0953, 32'h00000000} /* (14, 4, 4) {real, imag} */,
  {32'h3d0212d2, 32'h00000000} /* (14, 4, 3) {real, imag} */,
  {32'hbe2fdd99, 32'h00000000} /* (14, 4, 2) {real, imag} */,
  {32'h3e770289, 32'h00000000} /* (14, 4, 1) {real, imag} */,
  {32'h3e3f9c65, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'hbbcca100, 32'h00000000} /* (14, 3, 15) {real, imag} */,
  {32'h3dca7354, 32'h00000000} /* (14, 3, 14) {real, imag} */,
  {32'h3ebfc5e4, 32'h00000000} /* (14, 3, 13) {real, imag} */,
  {32'h3f401c41, 32'h00000000} /* (14, 3, 12) {real, imag} */,
  {32'h3eb3d948, 32'h00000000} /* (14, 3, 11) {real, imag} */,
  {32'h3db32831, 32'h00000000} /* (14, 3, 10) {real, imag} */,
  {32'hbdbe4914, 32'h00000000} /* (14, 3, 9) {real, imag} */,
  {32'hbda68f47, 32'h00000000} /* (14, 3, 8) {real, imag} */,
  {32'hbeb793f4, 32'h00000000} /* (14, 3, 7) {real, imag} */,
  {32'hbe81be46, 32'h00000000} /* (14, 3, 6) {real, imag} */,
  {32'hbf16fc10, 32'h00000000} /* (14, 3, 5) {real, imag} */,
  {32'hbf2636dc, 32'h00000000} /* (14, 3, 4) {real, imag} */,
  {32'h3e7008e0, 32'h00000000} /* (14, 3, 3) {real, imag} */,
  {32'h3db0530b, 32'h00000000} /* (14, 3, 2) {real, imag} */,
  {32'h3dd20508, 32'h00000000} /* (14, 3, 1) {real, imag} */,
  {32'h3f34d5a8, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h3ee83ace, 32'h00000000} /* (14, 2, 15) {real, imag} */,
  {32'h3f0bd215, 32'h00000000} /* (14, 2, 14) {real, imag} */,
  {32'h3f163733, 32'h00000000} /* (14, 2, 13) {real, imag} */,
  {32'h3f1b3be1, 32'h00000000} /* (14, 2, 12) {real, imag} */,
  {32'hbe44a0ef, 32'h00000000} /* (14, 2, 11) {real, imag} */,
  {32'h3eafab8e, 32'h00000000} /* (14, 2, 10) {real, imag} */,
  {32'hbcd61284, 32'h00000000} /* (14, 2, 9) {real, imag} */,
  {32'hbea08174, 32'h00000000} /* (14, 2, 8) {real, imag} */,
  {32'hbef84b8b, 32'h00000000} /* (14, 2, 7) {real, imag} */,
  {32'hbf269edd, 32'h00000000} /* (14, 2, 6) {real, imag} */,
  {32'hbf882fbe, 32'h00000000} /* (14, 2, 5) {real, imag} */,
  {32'hbf3e7b73, 32'h00000000} /* (14, 2, 4) {real, imag} */,
  {32'hbe3323e9, 32'h00000000} /* (14, 2, 3) {real, imag} */,
  {32'hbe3e6c51, 32'h00000000} /* (14, 2, 2) {real, imag} */,
  {32'hbebed993, 32'h00000000} /* (14, 2, 1) {real, imag} */,
  {32'h3e78432d, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h3e29ddc9, 32'h00000000} /* (14, 1, 15) {real, imag} */,
  {32'h3e66ca0f, 32'h00000000} /* (14, 1, 14) {real, imag} */,
  {32'h3e92cc92, 32'h00000000} /* (14, 1, 13) {real, imag} */,
  {32'h3ea9964a, 32'h00000000} /* (14, 1, 12) {real, imag} */,
  {32'hbedf46c3, 32'h00000000} /* (14, 1, 11) {real, imag} */,
  {32'h3da7be55, 32'h00000000} /* (14, 1, 10) {real, imag} */,
  {32'h3f3c110f, 32'h00000000} /* (14, 1, 9) {real, imag} */,
  {32'h3e28ff69, 32'h00000000} /* (14, 1, 8) {real, imag} */,
  {32'hbf53b1f7, 32'h00000000} /* (14, 1, 7) {real, imag} */,
  {32'hbf89596c, 32'h00000000} /* (14, 1, 6) {real, imag} */,
  {32'hbf8a5c81, 32'h00000000} /* (14, 1, 5) {real, imag} */,
  {32'hbf4b6092, 32'h00000000} /* (14, 1, 4) {real, imag} */,
  {32'hbec9af2b, 32'h00000000} /* (14, 1, 3) {real, imag} */,
  {32'hbe1ed7c9, 32'h00000000} /* (14, 1, 2) {real, imag} */,
  {32'hbf1de868, 32'h00000000} /* (14, 1, 1) {real, imag} */,
  {32'hbe941bc5, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h3d66e983, 32'h00000000} /* (14, 0, 15) {real, imag} */,
  {32'h3dcf7e5b, 32'h00000000} /* (14, 0, 14) {real, imag} */,
  {32'h3e8367a6, 32'h00000000} /* (14, 0, 13) {real, imag} */,
  {32'h3eb5f2bb, 32'h00000000} /* (14, 0, 12) {real, imag} */,
  {32'hbda88064, 32'h00000000} /* (14, 0, 11) {real, imag} */,
  {32'hbed3e6b4, 32'h00000000} /* (14, 0, 10) {real, imag} */,
  {32'h3df62907, 32'h00000000} /* (14, 0, 9) {real, imag} */,
  {32'h3e881b34, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hbf09d699, 32'h00000000} /* (14, 0, 7) {real, imag} */,
  {32'hbf0046df, 32'h00000000} /* (14, 0, 6) {real, imag} */,
  {32'hbe243e79, 32'h00000000} /* (14, 0, 5) {real, imag} */,
  {32'hbd110db0, 32'h00000000} /* (14, 0, 4) {real, imag} */,
  {32'h3d5e464b, 32'h00000000} /* (14, 0, 3) {real, imag} */,
  {32'h3dae4d7e, 32'h00000000} /* (14, 0, 2) {real, imag} */,
  {32'hbe277b65, 32'h00000000} /* (14, 0, 1) {real, imag} */,
  {32'hbd160d06, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h3e40c486, 32'h00000000} /* (13, 15, 15) {real, imag} */,
  {32'hbde9fe8c, 32'h00000000} /* (13, 15, 14) {real, imag} */,
  {32'hbe2a9a80, 32'h00000000} /* (13, 15, 13) {real, imag} */,
  {32'hbc363e64, 32'h00000000} /* (13, 15, 12) {real, imag} */,
  {32'h3c0a8e31, 32'h00000000} /* (13, 15, 11) {real, imag} */,
  {32'hbf3fe516, 32'h00000000} /* (13, 15, 10) {real, imag} */,
  {32'hbf0f0d95, 32'h00000000} /* (13, 15, 9) {real, imag} */,
  {32'hbe51a8b1, 32'h00000000} /* (13, 15, 8) {real, imag} */,
  {32'h3ded6091, 32'h00000000} /* (13, 15, 7) {real, imag} */,
  {32'hbded4989, 32'h00000000} /* (13, 15, 6) {real, imag} */,
  {32'h3c6e86f7, 32'h00000000} /* (13, 15, 5) {real, imag} */,
  {32'h3e07773b, 32'h00000000} /* (13, 15, 4) {real, imag} */,
  {32'h3e67c740, 32'h00000000} /* (13, 15, 3) {real, imag} */,
  {32'h3e3ba1e1, 32'h00000000} /* (13, 15, 2) {real, imag} */,
  {32'h3e7eb06c, 32'h00000000} /* (13, 15, 1) {real, imag} */,
  {32'h3f1651d5, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'h3e503efc, 32'h00000000} /* (13, 14, 15) {real, imag} */,
  {32'hbeb46bb7, 32'h00000000} /* (13, 14, 14) {real, imag} */,
  {32'hbefc6151, 32'h00000000} /* (13, 14, 13) {real, imag} */,
  {32'hbe8e9813, 32'h00000000} /* (13, 14, 12) {real, imag} */,
  {32'hbda094fd, 32'h00000000} /* (13, 14, 11) {real, imag} */,
  {32'hbf6fb568, 32'h00000000} /* (13, 14, 10) {real, imag} */,
  {32'hbf35dff7, 32'h00000000} /* (13, 14, 9) {real, imag} */,
  {32'hbec4df5f, 32'h00000000} /* (13, 14, 8) {real, imag} */,
  {32'h3e80614f, 32'h00000000} /* (13, 14, 7) {real, imag} */,
  {32'h3de2b435, 32'h00000000} /* (13, 14, 6) {real, imag} */,
  {32'hbe98f292, 32'h00000000} /* (13, 14, 5) {real, imag} */,
  {32'hbe2378f6, 32'h00000000} /* (13, 14, 4) {real, imag} */,
  {32'hbe56e0b1, 32'h00000000} /* (13, 14, 3) {real, imag} */,
  {32'hbefe759c, 32'h00000000} /* (13, 14, 2) {real, imag} */,
  {32'hbe971154, 32'h00000000} /* (13, 14, 1) {real, imag} */,
  {32'h3eb35b7e, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'h3dd9e3cc, 32'h00000000} /* (13, 13, 15) {real, imag} */,
  {32'hbeb06473, 32'h00000000} /* (13, 13, 14) {real, imag} */,
  {32'hbec2a3ac, 32'h00000000} /* (13, 13, 13) {real, imag} */,
  {32'hbec174b0, 32'h00000000} /* (13, 13, 12) {real, imag} */,
  {32'hbdf805b0, 32'h00000000} /* (13, 13, 11) {real, imag} */,
  {32'hbe154060, 32'h00000000} /* (13, 13, 10) {real, imag} */,
  {32'h3e19485a, 32'h00000000} /* (13, 13, 9) {real, imag} */,
  {32'hbe96a319, 32'h00000000} /* (13, 13, 8) {real, imag} */,
  {32'hbebfef7d, 32'h00000000} /* (13, 13, 7) {real, imag} */,
  {32'h3e4fafcf, 32'h00000000} /* (13, 13, 6) {real, imag} */,
  {32'hbe44f8af, 32'h00000000} /* (13, 13, 5) {real, imag} */,
  {32'hbe1490fb, 32'h00000000} /* (13, 13, 4) {real, imag} */,
  {32'hbe7bacf8, 32'h00000000} /* (13, 13, 3) {real, imag} */,
  {32'hbe9f8156, 32'h00000000} /* (13, 13, 2) {real, imag} */,
  {32'hbecc7ae8, 32'h00000000} /* (13, 13, 1) {real, imag} */,
  {32'hbe0490ce, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'h3d75f958, 32'h00000000} /* (13, 12, 15) {real, imag} */,
  {32'hbe076b23, 32'h00000000} /* (13, 12, 14) {real, imag} */,
  {32'hbc94886c, 32'h00000000} /* (13, 12, 13) {real, imag} */,
  {32'h3dbaf941, 32'h00000000} /* (13, 12, 12) {real, imag} */,
  {32'hbdf0e0a4, 32'h00000000} /* (13, 12, 11) {real, imag} */,
  {32'h3de4c380, 32'h00000000} /* (13, 12, 10) {real, imag} */,
  {32'h3f2a6ea6, 32'h00000000} /* (13, 12, 9) {real, imag} */,
  {32'h3d2021e3, 32'h00000000} /* (13, 12, 8) {real, imag} */,
  {32'hbf2f8bb9, 32'h00000000} /* (13, 12, 7) {real, imag} */,
  {32'hbf035451, 32'h00000000} /* (13, 12, 6) {real, imag} */,
  {32'hbd9ecf58, 32'h00000000} /* (13, 12, 5) {real, imag} */,
  {32'hbd33dc0e, 32'h00000000} /* (13, 12, 4) {real, imag} */,
  {32'hbe9d1eef, 32'h00000000} /* (13, 12, 3) {real, imag} */,
  {32'hbf419372, 32'h00000000} /* (13, 12, 2) {real, imag} */,
  {32'hbe6c8504, 32'h00000000} /* (13, 12, 1) {real, imag} */,
  {32'hbe969b84, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hbe3caed4, 32'h00000000} /* (13, 11, 15) {real, imag} */,
  {32'hbe763f13, 32'h00000000} /* (13, 11, 14) {real, imag} */,
  {32'h3d0254cc, 32'h00000000} /* (13, 11, 13) {real, imag} */,
  {32'h3e36b89d, 32'h00000000} /* (13, 11, 12) {real, imag} */,
  {32'h3e94d811, 32'h00000000} /* (13, 11, 11) {real, imag} */,
  {32'hbe47b230, 32'h00000000} /* (13, 11, 10) {real, imag} */,
  {32'h3ebd1761, 32'h00000000} /* (13, 11, 9) {real, imag} */,
  {32'h3efb13dd, 32'h00000000} /* (13, 11, 8) {real, imag} */,
  {32'hbe431546, 32'h00000000} /* (13, 11, 7) {real, imag} */,
  {32'hbf4c67a1, 32'h00000000} /* (13, 11, 6) {real, imag} */,
  {32'hbed4e710, 32'h00000000} /* (13, 11, 5) {real, imag} */,
  {32'hbbbb9f9d, 32'h00000000} /* (13, 11, 4) {real, imag} */,
  {32'hbe2b4bcd, 32'h00000000} /* (13, 11, 3) {real, imag} */,
  {32'hbf2f5c88, 32'h00000000} /* (13, 11, 2) {real, imag} */,
  {32'hbe4579db, 32'h00000000} /* (13, 11, 1) {real, imag} */,
  {32'hbe610f40, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'hbda3347b, 32'h00000000} /* (13, 10, 15) {real, imag} */,
  {32'hbe3d54b6, 32'h00000000} /* (13, 10, 14) {real, imag} */,
  {32'h3dc09bf9, 32'h00000000} /* (13, 10, 13) {real, imag} */,
  {32'h3ee90056, 32'h00000000} /* (13, 10, 12) {real, imag} */,
  {32'h3ea33dc7, 32'h00000000} /* (13, 10, 11) {real, imag} */,
  {32'hbe8fdcbb, 32'h00000000} /* (13, 10, 10) {real, imag} */,
  {32'hbda11876, 32'h00000000} /* (13, 10, 9) {real, imag} */,
  {32'hbdad988c, 32'h00000000} /* (13, 10, 8) {real, imag} */,
  {32'h3e06e947, 32'h00000000} /* (13, 10, 7) {real, imag} */,
  {32'h3d6fa310, 32'h00000000} /* (13, 10, 6) {real, imag} */,
  {32'hbe9c2704, 32'h00000000} /* (13, 10, 5) {real, imag} */,
  {32'hbdaffdf8, 32'h00000000} /* (13, 10, 4) {real, imag} */,
  {32'h3e68cd2f, 32'h00000000} /* (13, 10, 3) {real, imag} */,
  {32'hbeb7e1f4, 32'h00000000} /* (13, 10, 2) {real, imag} */,
  {32'hbdda2d68, 32'h00000000} /* (13, 10, 1) {real, imag} */,
  {32'h3e44dc2d, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h3f037755, 32'h00000000} /* (13, 9, 15) {real, imag} */,
  {32'h3f21c17c, 32'h00000000} /* (13, 9, 14) {real, imag} */,
  {32'h3e0fb234, 32'h00000000} /* (13, 9, 13) {real, imag} */,
  {32'h3ed4e09e, 32'h00000000} /* (13, 9, 12) {real, imag} */,
  {32'h3e8e583f, 32'h00000000} /* (13, 9, 11) {real, imag} */,
  {32'h3d18dc2c, 32'h00000000} /* (13, 9, 10) {real, imag} */,
  {32'hbedf3ef0, 32'h00000000} /* (13, 9, 9) {real, imag} */,
  {32'hbef5c762, 32'h00000000} /* (13, 9, 8) {real, imag} */,
  {32'hbe7d3490, 32'h00000000} /* (13, 9, 7) {real, imag} */,
  {32'hbe1a4053, 32'h00000000} /* (13, 9, 6) {real, imag} */,
  {32'h3dd13341, 32'h00000000} /* (13, 9, 5) {real, imag} */,
  {32'hbda79763, 32'h00000000} /* (13, 9, 4) {real, imag} */,
  {32'hbc4b2881, 32'h00000000} /* (13, 9, 3) {real, imag} */,
  {32'h3d4de570, 32'h00000000} /* (13, 9, 2) {real, imag} */,
  {32'hbe4ea840, 32'h00000000} /* (13, 9, 1) {real, imag} */,
  {32'h3dcc525e, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'hbe2ae800, 32'h00000000} /* (13, 8, 15) {real, imag} */,
  {32'h3d00dd77, 32'h00000000} /* (13, 8, 14) {real, imag} */,
  {32'h3d1672ca, 32'h00000000} /* (13, 8, 13) {real, imag} */,
  {32'h3e2a392e, 32'h00000000} /* (13, 8, 12) {real, imag} */,
  {32'h3e6ed48d, 32'h00000000} /* (13, 8, 11) {real, imag} */,
  {32'h3bea8ca1, 32'h00000000} /* (13, 8, 10) {real, imag} */,
  {32'hbd270b64, 32'h00000000} /* (13, 8, 9) {real, imag} */,
  {32'h3dbeae5d, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'hbe5b3fc0, 32'h00000000} /* (13, 8, 7) {real, imag} */,
  {32'hbed7979a, 32'h00000000} /* (13, 8, 6) {real, imag} */,
  {32'hbe79c69d, 32'h00000000} /* (13, 8, 5) {real, imag} */,
  {32'hbdf59804, 32'h00000000} /* (13, 8, 4) {real, imag} */,
  {32'hbe8dfe67, 32'h00000000} /* (13, 8, 3) {real, imag} */,
  {32'h3e0c26f5, 32'h00000000} /* (13, 8, 2) {real, imag} */,
  {32'hbe224e1c, 32'h00000000} /* (13, 8, 1) {real, imag} */,
  {32'hbf0459c9, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'hbf121200, 32'h00000000} /* (13, 7, 15) {real, imag} */,
  {32'hbf1dd1dd, 32'h00000000} /* (13, 7, 14) {real, imag} */,
  {32'hbea2c532, 32'h00000000} /* (13, 7, 13) {real, imag} */,
  {32'h3ed00e28, 32'h00000000} /* (13, 7, 12) {real, imag} */,
  {32'h3f04c7c7, 32'h00000000} /* (13, 7, 11) {real, imag} */,
  {32'h3e5abe21, 32'h00000000} /* (13, 7, 10) {real, imag} */,
  {32'h3ea46bff, 32'h00000000} /* (13, 7, 9) {real, imag} */,
  {32'h3e698555, 32'h00000000} /* (13, 7, 8) {real, imag} */,
  {32'h3db6b18a, 32'h00000000} /* (13, 7, 7) {real, imag} */,
  {32'h3e6bb367, 32'h00000000} /* (13, 7, 6) {real, imag} */,
  {32'hbd8a0576, 32'h00000000} /* (13, 7, 5) {real, imag} */,
  {32'hbd8e5b49, 32'h00000000} /* (13, 7, 4) {real, imag} */,
  {32'h3ea35bb6, 32'h00000000} /* (13, 7, 3) {real, imag} */,
  {32'h3eef2cb3, 32'h00000000} /* (13, 7, 2) {real, imag} */,
  {32'h3e1bd6a4, 32'h00000000} /* (13, 7, 1) {real, imag} */,
  {32'hbf07777e, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'hbe6cb5ed, 32'h00000000} /* (13, 6, 15) {real, imag} */,
  {32'hbe58b18f, 32'h00000000} /* (13, 6, 14) {real, imag} */,
  {32'hbe36d139, 32'h00000000} /* (13, 6, 13) {real, imag} */,
  {32'h3dc212da, 32'h00000000} /* (13, 6, 12) {real, imag} */,
  {32'h3e05ba56, 32'h00000000} /* (13, 6, 11) {real, imag} */,
  {32'h3f1fe056, 32'h00000000} /* (13, 6, 10) {real, imag} */,
  {32'h3f3228e5, 32'h00000000} /* (13, 6, 9) {real, imag} */,
  {32'hbd7bb129, 32'h00000000} /* (13, 6, 8) {real, imag} */,
  {32'h3f3b64f2, 32'h00000000} /* (13, 6, 7) {real, imag} */,
  {32'h3ec8d95d, 32'h00000000} /* (13, 6, 6) {real, imag} */,
  {32'h3dda3dfa, 32'h00000000} /* (13, 6, 5) {real, imag} */,
  {32'hbe453a97, 32'h00000000} /* (13, 6, 4) {real, imag} */,
  {32'h3e2220d3, 32'h00000000} /* (13, 6, 3) {real, imag} */,
  {32'h3dfba06c, 32'h00000000} /* (13, 6, 2) {real, imag} */,
  {32'hbe26d726, 32'h00000000} /* (13, 6, 1) {real, imag} */,
  {32'h3d456484, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h3db066e9, 32'h00000000} /* (13, 5, 15) {real, imag} */,
  {32'h3e2d4f5b, 32'h00000000} /* (13, 5, 14) {real, imag} */,
  {32'hbdf8538a, 32'h00000000} /* (13, 5, 13) {real, imag} */,
  {32'hbe4637cd, 32'h00000000} /* (13, 5, 12) {real, imag} */,
  {32'hbe676609, 32'h00000000} /* (13, 5, 11) {real, imag} */,
  {32'h3ddadcc9, 32'h00000000} /* (13, 5, 10) {real, imag} */,
  {32'h3e518bf9, 32'h00000000} /* (13, 5, 9) {real, imag} */,
  {32'hbe8b8f14, 32'h00000000} /* (13, 5, 8) {real, imag} */,
  {32'h3e79d9ac, 32'h00000000} /* (13, 5, 7) {real, imag} */,
  {32'h3eb13354, 32'h00000000} /* (13, 5, 6) {real, imag} */,
  {32'h3d4ce235, 32'h00000000} /* (13, 5, 5) {real, imag} */,
  {32'h3ed91999, 32'h00000000} /* (13, 5, 4) {real, imag} */,
  {32'h3f1cb988, 32'h00000000} /* (13, 5, 3) {real, imag} */,
  {32'h3e9da6bb, 32'h00000000} /* (13, 5, 2) {real, imag} */,
  {32'h3d4ee66f, 32'h00000000} /* (13, 5, 1) {real, imag} */,
  {32'h3cc54e6d, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h3e096d9e, 32'h00000000} /* (13, 4, 15) {real, imag} */,
  {32'h3dafde0f, 32'h00000000} /* (13, 4, 14) {real, imag} */,
  {32'h3e3c7340, 32'h00000000} /* (13, 4, 13) {real, imag} */,
  {32'h3f000d56, 32'h00000000} /* (13, 4, 12) {real, imag} */,
  {32'hbe805303, 32'h00000000} /* (13, 4, 11) {real, imag} */,
  {32'hbe6889f5, 32'h00000000} /* (13, 4, 10) {real, imag} */,
  {32'h3d4aa257, 32'h00000000} /* (13, 4, 9) {real, imag} */,
  {32'h3efd1df7, 32'h00000000} /* (13, 4, 8) {real, imag} */,
  {32'h3e9beac6, 32'h00000000} /* (13, 4, 7) {real, imag} */,
  {32'hbcfb5e49, 32'h00000000} /* (13, 4, 6) {real, imag} */,
  {32'hbf0b7869, 32'h00000000} /* (13, 4, 5) {real, imag} */,
  {32'hbe5f05db, 32'h00000000} /* (13, 4, 4) {real, imag} */,
  {32'h3edc5a43, 32'h00000000} /* (13, 4, 3) {real, imag} */,
  {32'hbc764a7a, 32'h00000000} /* (13, 4, 2) {real, imag} */,
  {32'h3e2dc4ef, 32'h00000000} /* (13, 4, 1) {real, imag} */,
  {32'h3e408b76, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'hbe261f56, 32'h00000000} /* (13, 3, 15) {real, imag} */,
  {32'hbe6b780c, 32'h00000000} /* (13, 3, 14) {real, imag} */,
  {32'h3f71eeea, 32'h00000000} /* (13, 3, 13) {real, imag} */,
  {32'h3faa95f7, 32'h00000000} /* (13, 3, 12) {real, imag} */,
  {32'h3eb5c9c8, 32'h00000000} /* (13, 3, 11) {real, imag} */,
  {32'hbe975c3f, 32'h00000000} /* (13, 3, 10) {real, imag} */,
  {32'hba9d387e, 32'h00000000} /* (13, 3, 9) {real, imag} */,
  {32'h3f3bd31e, 32'h00000000} /* (13, 3, 8) {real, imag} */,
  {32'h3ef968d4, 32'h00000000} /* (13, 3, 7) {real, imag} */,
  {32'hbeb5b14f, 32'h00000000} /* (13, 3, 6) {real, imag} */,
  {32'hbf0ac358, 32'h00000000} /* (13, 3, 5) {real, imag} */,
  {32'hbe9e0ffc, 32'h00000000} /* (13, 3, 4) {real, imag} */,
  {32'h3f08f4b9, 32'h00000000} /* (13, 3, 3) {real, imag} */,
  {32'h3da94169, 32'h00000000} /* (13, 3, 2) {real, imag} */,
  {32'hbd15158d, 32'h00000000} /* (13, 3, 1) {real, imag} */,
  {32'h3e87c54c, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h3ea4544a, 32'h00000000} /* (13, 2, 15) {real, imag} */,
  {32'h3ec3c710, 32'h00000000} /* (13, 2, 14) {real, imag} */,
  {32'h3f4c7102, 32'h00000000} /* (13, 2, 13) {real, imag} */,
  {32'h3f412c5a, 32'h00000000} /* (13, 2, 12) {real, imag} */,
  {32'hbe31b8fd, 32'h00000000} /* (13, 2, 11) {real, imag} */,
  {32'hbf1328f6, 32'h00000000} /* (13, 2, 10) {real, imag} */,
  {32'hbe91de12, 32'h00000000} /* (13, 2, 9) {real, imag} */,
  {32'hbe0d16c8, 32'h00000000} /* (13, 2, 8) {real, imag} */,
  {32'h3e4de79d, 32'h00000000} /* (13, 2, 7) {real, imag} */,
  {32'hbe9cfd16, 32'h00000000} /* (13, 2, 6) {real, imag} */,
  {32'hbf1361d9, 32'h00000000} /* (13, 2, 5) {real, imag} */,
  {32'hbe77d1fc, 32'h00000000} /* (13, 2, 4) {real, imag} */,
  {32'h3e6840c6, 32'h00000000} /* (13, 2, 3) {real, imag} */,
  {32'h3e16b045, 32'h00000000} /* (13, 2, 2) {real, imag} */,
  {32'h3d96349b, 32'h00000000} /* (13, 2, 1) {real, imag} */,
  {32'h3de636b1, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h3e748f00, 32'h00000000} /* (13, 1, 15) {real, imag} */,
  {32'h3ea42b27, 32'h00000000} /* (13, 1, 14) {real, imag} */,
  {32'h3f5883ce, 32'h00000000} /* (13, 1, 13) {real, imag} */,
  {32'h3ee98b75, 32'h00000000} /* (13, 1, 12) {real, imag} */,
  {32'hbf0e81fc, 32'h00000000} /* (13, 1, 11) {real, imag} */,
  {32'hbeb851bb, 32'h00000000} /* (13, 1, 10) {real, imag} */,
  {32'h3edab030, 32'h00000000} /* (13, 1, 9) {real, imag} */,
  {32'h3df5767e, 32'h00000000} /* (13, 1, 8) {real, imag} */,
  {32'hbee1753e, 32'h00000000} /* (13, 1, 7) {real, imag} */,
  {32'hbeaf9421, 32'h00000000} /* (13, 1, 6) {real, imag} */,
  {32'hbd5dd825, 32'h00000000} /* (13, 1, 5) {real, imag} */,
  {32'hbed7aa63, 32'h00000000} /* (13, 1, 4) {real, imag} */,
  {32'hbee61ec7, 32'h00000000} /* (13, 1, 3) {real, imag} */,
  {32'hbceb79fc, 32'h00000000} /* (13, 1, 2) {real, imag} */,
  {32'hbd7e330b, 32'h00000000} /* (13, 1, 1) {real, imag} */,
  {32'hbd0da717, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h3d48ccf0, 32'h00000000} /* (13, 0, 15) {real, imag} */,
  {32'h3d9682db, 32'h00000000} /* (13, 0, 14) {real, imag} */,
  {32'h3f17dfd4, 32'h00000000} /* (13, 0, 13) {real, imag} */,
  {32'h3ec1b868, 32'h00000000} /* (13, 0, 12) {real, imag} */,
  {32'hbe8a4660, 32'h00000000} /* (13, 0, 11) {real, imag} */,
  {32'hbe9caf11, 32'h00000000} /* (13, 0, 10) {real, imag} */,
  {32'h3e9c9c98, 32'h00000000} /* (13, 0, 9) {real, imag} */,
  {32'h3eed3440, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'hbe1e8cba, 32'h00000000} /* (13, 0, 7) {real, imag} */,
  {32'hbe17a88f, 32'h00000000} /* (13, 0, 6) {real, imag} */,
  {32'h3e91d7a9, 32'h00000000} /* (13, 0, 5) {real, imag} */,
  {32'h3e49ff5a, 32'h00000000} /* (13, 0, 4) {real, imag} */,
  {32'h3e1e5e54, 32'h00000000} /* (13, 0, 3) {real, imag} */,
  {32'h3e03c86d, 32'h00000000} /* (13, 0, 2) {real, imag} */,
  {32'h3dfef2a8, 32'h00000000} /* (13, 0, 1) {real, imag} */,
  {32'h3e4f6290, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h3e30d7a4, 32'h00000000} /* (12, 15, 15) {real, imag} */,
  {32'hbd856b7d, 32'h00000000} /* (12, 15, 14) {real, imag} */,
  {32'hbeb89aa6, 32'h00000000} /* (12, 15, 13) {real, imag} */,
  {32'h3add9fa2, 32'h00000000} /* (12, 15, 12) {real, imag} */,
  {32'h3da54a21, 32'h00000000} /* (12, 15, 11) {real, imag} */,
  {32'hbf257174, 32'h00000000} /* (12, 15, 10) {real, imag} */,
  {32'hbec02650, 32'h00000000} /* (12, 15, 9) {real, imag} */,
  {32'hbee71efe, 32'h00000000} /* (12, 15, 8) {real, imag} */,
  {32'hbdf8ef55, 32'h00000000} /* (12, 15, 7) {real, imag} */,
  {32'hbd576c8b, 32'h00000000} /* (12, 15, 6) {real, imag} */,
  {32'hbdf77f5b, 32'h00000000} /* (12, 15, 5) {real, imag} */,
  {32'h3ece922a, 32'h00000000} /* (12, 15, 4) {real, imag} */,
  {32'h3f25404e, 32'h00000000} /* (12, 15, 3) {real, imag} */,
  {32'h3e64013e, 32'h00000000} /* (12, 15, 2) {real, imag} */,
  {32'hbcaa3313, 32'h00000000} /* (12, 15, 1) {real, imag} */,
  {32'h3cb1685b, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'h3e894356, 32'h00000000} /* (12, 14, 15) {real, imag} */,
  {32'hbe493140, 32'h00000000} /* (12, 14, 14) {real, imag} */,
  {32'hbf1215a9, 32'h00000000} /* (12, 14, 13) {real, imag} */,
  {32'hbf0b044c, 32'h00000000} /* (12, 14, 12) {real, imag} */,
  {32'hbe4accc6, 32'h00000000} /* (12, 14, 11) {real, imag} */,
  {32'hbf9072f4, 32'h00000000} /* (12, 14, 10) {real, imag} */,
  {32'hbeeb0685, 32'h00000000} /* (12, 14, 9) {real, imag} */,
  {32'hbedb59b3, 32'h00000000} /* (12, 14, 8) {real, imag} */,
  {32'h3e856137, 32'h00000000} /* (12, 14, 7) {real, imag} */,
  {32'h3eb3e339, 32'h00000000} /* (12, 14, 6) {real, imag} */,
  {32'hbd71a56c, 32'h00000000} /* (12, 14, 5) {real, imag} */,
  {32'h3ea5b4ac, 32'h00000000} /* (12, 14, 4) {real, imag} */,
  {32'h3ede66ac, 32'h00000000} /* (12, 14, 3) {real, imag} */,
  {32'h3d977586, 32'h00000000} /* (12, 14, 2) {real, imag} */,
  {32'hbd9f6d4d, 32'h00000000} /* (12, 14, 1) {real, imag} */,
  {32'hbe0e609c, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'h3e7656cb, 32'h00000000} /* (12, 13, 15) {real, imag} */,
  {32'h3e051188, 32'h00000000} /* (12, 13, 14) {real, imag} */,
  {32'hbe243951, 32'h00000000} /* (12, 13, 13) {real, imag} */,
  {32'hbf06e09c, 32'h00000000} /* (12, 13, 12) {real, imag} */,
  {32'hbdd6fdce, 32'h00000000} /* (12, 13, 11) {real, imag} */,
  {32'hbd62ca97, 32'h00000000} /* (12, 13, 10) {real, imag} */,
  {32'h3deb8659, 32'h00000000} /* (12, 13, 9) {real, imag} */,
  {32'hbe6b5451, 32'h00000000} /* (12, 13, 8) {real, imag} */,
  {32'hbdca7173, 32'h00000000} /* (12, 13, 7) {real, imag} */,
  {32'h3d9a90a6, 32'h00000000} /* (12, 13, 6) {real, imag} */,
  {32'h3e266a98, 32'h00000000} /* (12, 13, 5) {real, imag} */,
  {32'h3ec1528d, 32'h00000000} /* (12, 13, 4) {real, imag} */,
  {32'hbd865f26, 32'h00000000} /* (12, 13, 3) {real, imag} */,
  {32'hbe94713b, 32'h00000000} /* (12, 13, 2) {real, imag} */,
  {32'hbe0b8342, 32'h00000000} /* (12, 13, 1) {real, imag} */,
  {32'hbdade333, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'h3eae8d57, 32'h00000000} /* (12, 12, 15) {real, imag} */,
  {32'h3e829ed5, 32'h00000000} /* (12, 12, 14) {real, imag} */,
  {32'hbe3088d8, 32'h00000000} /* (12, 12, 13) {real, imag} */,
  {32'h3e2b12f6, 32'h00000000} /* (12, 12, 12) {real, imag} */,
  {32'h3e22667b, 32'h00000000} /* (12, 12, 11) {real, imag} */,
  {32'h3e53262e, 32'h00000000} /* (12, 12, 10) {real, imag} */,
  {32'h3ea5cb92, 32'h00000000} /* (12, 12, 9) {real, imag} */,
  {32'hbe3d1ce9, 32'h00000000} /* (12, 12, 8) {real, imag} */,
  {32'hbef3af08, 32'h00000000} /* (12, 12, 7) {real, imag} */,
  {32'hbed5df30, 32'h00000000} /* (12, 12, 6) {real, imag} */,
  {32'h3e0258e3, 32'h00000000} /* (12, 12, 5) {real, imag} */,
  {32'h3df5423b, 32'h00000000} /* (12, 12, 4) {real, imag} */,
  {32'hbe5ef1d5, 32'h00000000} /* (12, 12, 3) {real, imag} */,
  {32'hbf34cf28, 32'h00000000} /* (12, 12, 2) {real, imag} */,
  {32'hbe6039ff, 32'h00000000} /* (12, 12, 1) {real, imag} */,
  {32'h3df2e78c, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'h3bd12324, 32'h00000000} /* (12, 11, 15) {real, imag} */,
  {32'hbe8985bb, 32'h00000000} /* (12, 11, 14) {real, imag} */,
  {32'hbceded31, 32'h00000000} /* (12, 11, 13) {real, imag} */,
  {32'h3ef2728e, 32'h00000000} /* (12, 11, 12) {real, imag} */,
  {32'h3f015fda, 32'h00000000} /* (12, 11, 11) {real, imag} */,
  {32'h3d8f79aa, 32'h00000000} /* (12, 11, 10) {real, imag} */,
  {32'h3eb55781, 32'h00000000} /* (12, 11, 9) {real, imag} */,
  {32'h3ecee7a0, 32'h00000000} /* (12, 11, 8) {real, imag} */,
  {32'h3eb55830, 32'h00000000} /* (12, 11, 7) {real, imag} */,
  {32'hbe2852c2, 32'h00000000} /* (12, 11, 6) {real, imag} */,
  {32'hbe70834c, 32'h00000000} /* (12, 11, 5) {real, imag} */,
  {32'hbec93fcb, 32'h00000000} /* (12, 11, 4) {real, imag} */,
  {32'hbe53ed75, 32'h00000000} /* (12, 11, 3) {real, imag} */,
  {32'hbcdc1a6e, 32'h00000000} /* (12, 11, 2) {real, imag} */,
  {32'h3d8eccb6, 32'h00000000} /* (12, 11, 1) {real, imag} */,
  {32'h3dab503d, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h3c95f6b8, 32'h00000000} /* (12, 10, 15) {real, imag} */,
  {32'hbeba43dc, 32'h00000000} /* (12, 10, 14) {real, imag} */,
  {32'hbd44b538, 32'h00000000} /* (12, 10, 13) {real, imag} */,
  {32'h3efb8203, 32'h00000000} /* (12, 10, 12) {real, imag} */,
  {32'h3f12df00, 32'h00000000} /* (12, 10, 11) {real, imag} */,
  {32'h3e8c8ba6, 32'h00000000} /* (12, 10, 10) {real, imag} */,
  {32'h3e1b9f8c, 32'h00000000} /* (12, 10, 9) {real, imag} */,
  {32'h3d1cd1d2, 32'h00000000} /* (12, 10, 8) {real, imag} */,
  {32'h3ec08db9, 32'h00000000} /* (12, 10, 7) {real, imag} */,
  {32'h3dab81dd, 32'h00000000} /* (12, 10, 6) {real, imag} */,
  {32'hbf19e030, 32'h00000000} /* (12, 10, 5) {real, imag} */,
  {32'hbebf0b9c, 32'h00000000} /* (12, 10, 4) {real, imag} */,
  {32'hbe182b97, 32'h00000000} /* (12, 10, 3) {real, imag} */,
  {32'h3d20ebf9, 32'h00000000} /* (12, 10, 2) {real, imag} */,
  {32'h3e4a3337, 32'h00000000} /* (12, 10, 1) {real, imag} */,
  {32'h3da6417f, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h3dedad8c, 32'h00000000} /* (12, 9, 15) {real, imag} */,
  {32'hbd2259f9, 32'h00000000} /* (12, 9, 14) {real, imag} */,
  {32'hbd5d5c37, 32'h00000000} /* (12, 9, 13) {real, imag} */,
  {32'h3ea9b0e1, 32'h00000000} /* (12, 9, 12) {real, imag} */,
  {32'h3f13db11, 32'h00000000} /* (12, 9, 11) {real, imag} */,
  {32'h3e6c0617, 32'h00000000} /* (12, 9, 10) {real, imag} */,
  {32'hbdfaed60, 32'h00000000} /* (12, 9, 9) {real, imag} */,
  {32'hbf2c7183, 32'h00000000} /* (12, 9, 8) {real, imag} */,
  {32'hbdd76ad6, 32'h00000000} /* (12, 9, 7) {real, imag} */,
  {32'hbe964c61, 32'h00000000} /* (12, 9, 6) {real, imag} */,
  {32'hbf5376e7, 32'h00000000} /* (12, 9, 5) {real, imag} */,
  {32'hbf14a02f, 32'h00000000} /* (12, 9, 4) {real, imag} */,
  {32'hbee734bc, 32'h00000000} /* (12, 9, 3) {real, imag} */,
  {32'h3d9e349b, 32'h00000000} /* (12, 9, 2) {real, imag} */,
  {32'h3eed7d70, 32'h00000000} /* (12, 9, 1) {real, imag} */,
  {32'h3db5c292, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'hbd8a6cfc, 32'h00000000} /* (12, 8, 15) {real, imag} */,
  {32'h3de2f582, 32'h00000000} /* (12, 8, 14) {real, imag} */,
  {32'hbdb99bda, 32'h00000000} /* (12, 8, 13) {real, imag} */,
  {32'hbea50af0, 32'h00000000} /* (12, 8, 12) {real, imag} */,
  {32'h3ca7015d, 32'h00000000} /* (12, 8, 11) {real, imag} */,
  {32'hbe22afb9, 32'h00000000} /* (12, 8, 10) {real, imag} */,
  {32'h3d020350, 32'h00000000} /* (12, 8, 9) {real, imag} */,
  {32'hbd91310b, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'hbe4e3f07, 32'h00000000} /* (12, 8, 7) {real, imag} */,
  {32'hbeb6c461, 32'h00000000} /* (12, 8, 6) {real, imag} */,
  {32'hbf68a8cc, 32'h00000000} /* (12, 8, 5) {real, imag} */,
  {32'hbf42a017, 32'h00000000} /* (12, 8, 4) {real, imag} */,
  {32'hbf3d1508, 32'h00000000} /* (12, 8, 3) {real, imag} */,
  {32'hbe9278f4, 32'h00000000} /* (12, 8, 2) {real, imag} */,
  {32'h3e2f63c0, 32'h00000000} /* (12, 8, 1) {real, imag} */,
  {32'hbd92958f, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'hbf55784e, 32'h00000000} /* (12, 7, 15) {real, imag} */,
  {32'hbf34dba4, 32'h00000000} /* (12, 7, 14) {real, imag} */,
  {32'hbf00ff89, 32'h00000000} /* (12, 7, 13) {real, imag} */,
  {32'hbdfc7dc0, 32'h00000000} /* (12, 7, 12) {real, imag} */,
  {32'h3ece6f12, 32'h00000000} /* (12, 7, 11) {real, imag} */,
  {32'h3ca8d2b5, 32'h00000000} /* (12, 7, 10) {real, imag} */,
  {32'h3e0813b3, 32'h00000000} /* (12, 7, 9) {real, imag} */,
  {32'h3e71bf70, 32'h00000000} /* (12, 7, 8) {real, imag} */,
  {32'h3dcb153b, 32'h00000000} /* (12, 7, 7) {real, imag} */,
  {32'h3dcd4b53, 32'h00000000} /* (12, 7, 6) {real, imag} */,
  {32'hbe8fd898, 32'h00000000} /* (12, 7, 5) {real, imag} */,
  {32'hbeadf416, 32'h00000000} /* (12, 7, 4) {real, imag} */,
  {32'hbd34ea42, 32'h00000000} /* (12, 7, 3) {real, imag} */,
  {32'hbd04ae82, 32'h00000000} /* (12, 7, 2) {real, imag} */,
  {32'hbe672073, 32'h00000000} /* (12, 7, 1) {real, imag} */,
  {32'hbe98a865, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'hbf3e1f75, 32'h00000000} /* (12, 6, 15) {real, imag} */,
  {32'hbeefd364, 32'h00000000} /* (12, 6, 14) {real, imag} */,
  {32'hbe337c72, 32'h00000000} /* (12, 6, 13) {real, imag} */,
  {32'hbe3ce753, 32'h00000000} /* (12, 6, 12) {real, imag} */,
  {32'h3e007b55, 32'h00000000} /* (12, 6, 11) {real, imag} */,
  {32'hbcada07e, 32'h00000000} /* (12, 6, 10) {real, imag} */,
  {32'h3ecb36e6, 32'h00000000} /* (12, 6, 9) {real, imag} */,
  {32'h3d9720e5, 32'h00000000} /* (12, 6, 8) {real, imag} */,
  {32'h3f397502, 32'h00000000} /* (12, 6, 7) {real, imag} */,
  {32'h3f0c326c, 32'h00000000} /* (12, 6, 6) {real, imag} */,
  {32'h3f36463f, 32'h00000000} /* (12, 6, 5) {real, imag} */,
  {32'h3ed62482, 32'h00000000} /* (12, 6, 4) {real, imag} */,
  {32'h3e11eb72, 32'h00000000} /* (12, 6, 3) {real, imag} */,
  {32'hbec2aab9, 32'h00000000} /* (12, 6, 2) {real, imag} */,
  {32'hbf6de0d8, 32'h00000000} /* (12, 6, 1) {real, imag} */,
  {32'hbe61ca88, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'hbd1c3d7c, 32'h00000000} /* (12, 5, 15) {real, imag} */,
  {32'h3e1f2786, 32'h00000000} /* (12, 5, 14) {real, imag} */,
  {32'h3c01b2c0, 32'h00000000} /* (12, 5, 13) {real, imag} */,
  {32'hbd9f5682, 32'h00000000} /* (12, 5, 12) {real, imag} */,
  {32'hbef00beb, 32'h00000000} /* (12, 5, 11) {real, imag} */,
  {32'hbeae862f, 32'h00000000} /* (12, 5, 10) {real, imag} */,
  {32'h3e3d1032, 32'h00000000} /* (12, 5, 9) {real, imag} */,
  {32'hbeefef37, 32'h00000000} /* (12, 5, 8) {real, imag} */,
  {32'h3f0716bc, 32'h00000000} /* (12, 5, 7) {real, imag} */,
  {32'h3f1052f5, 32'h00000000} /* (12, 5, 6) {real, imag} */,
  {32'h3e94431d, 32'h00000000} /* (12, 5, 5) {real, imag} */,
  {32'h3f09e79d, 32'h00000000} /* (12, 5, 4) {real, imag} */,
  {32'h3eed957b, 32'h00000000} /* (12, 5, 3) {real, imag} */,
  {32'h3e2d7ea3, 32'h00000000} /* (12, 5, 2) {real, imag} */,
  {32'hbe778a91, 32'h00000000} /* (12, 5, 1) {real, imag} */,
  {32'hbd9eb4ce, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h3e3ecd75, 32'h00000000} /* (12, 4, 15) {real, imag} */,
  {32'h3e3eaf86, 32'h00000000} /* (12, 4, 14) {real, imag} */,
  {32'h3e414fb0, 32'h00000000} /* (12, 4, 13) {real, imag} */,
  {32'h3f212afe, 32'h00000000} /* (12, 4, 12) {real, imag} */,
  {32'hbe6bf1a8, 32'h00000000} /* (12, 4, 11) {real, imag} */,
  {32'hbeadaedf, 32'h00000000} /* (12, 4, 10) {real, imag} */,
  {32'hbe202f03, 32'h00000000} /* (12, 4, 9) {real, imag} */,
  {32'h3d17b584, 32'h00000000} /* (12, 4, 8) {real, imag} */,
  {32'h3ee7fa5b, 32'h00000000} /* (12, 4, 7) {real, imag} */,
  {32'h3eacc647, 32'h00000000} /* (12, 4, 6) {real, imag} */,
  {32'h3e936389, 32'h00000000} /* (12, 4, 5) {real, imag} */,
  {32'h3ec46698, 32'h00000000} /* (12, 4, 4) {real, imag} */,
  {32'h3ee4794c, 32'h00000000} /* (12, 4, 3) {real, imag} */,
  {32'h3dfc0a4b, 32'h00000000} /* (12, 4, 2) {real, imag} */,
  {32'h3e08e0b5, 32'h00000000} /* (12, 4, 1) {real, imag} */,
  {32'hbbbc0f1d, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h3d9f6f4b, 32'h00000000} /* (12, 3, 15) {real, imag} */,
  {32'hbcc1005a, 32'h00000000} /* (12, 3, 14) {real, imag} */,
  {32'h3eb2d24d, 32'h00000000} /* (12, 3, 13) {real, imag} */,
  {32'h3f384709, 32'h00000000} /* (12, 3, 12) {real, imag} */,
  {32'h3e5b6bcf, 32'h00000000} /* (12, 3, 11) {real, imag} */,
  {32'h3d55424d, 32'h00000000} /* (12, 3, 10) {real, imag} */,
  {32'hbe21ef0a, 32'h00000000} /* (12, 3, 9) {real, imag} */,
  {32'h3e0388c8, 32'h00000000} /* (12, 3, 8) {real, imag} */,
  {32'h3f03cca0, 32'h00000000} /* (12, 3, 7) {real, imag} */,
  {32'h3ed39380, 32'h00000000} /* (12, 3, 6) {real, imag} */,
  {32'hbd7d5378, 32'h00000000} /* (12, 3, 5) {real, imag} */,
  {32'h3def3d16, 32'h00000000} /* (12, 3, 4) {real, imag} */,
  {32'h3e8aed3d, 32'h00000000} /* (12, 3, 3) {real, imag} */,
  {32'hbeab9399, 32'h00000000} /* (12, 3, 2) {real, imag} */,
  {32'hbaee7988, 32'h00000000} /* (12, 3, 1) {real, imag} */,
  {32'hbdbf98c7, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'hbcdb6a8b, 32'h00000000} /* (12, 2, 15) {real, imag} */,
  {32'hbe943d42, 32'h00000000} /* (12, 2, 14) {real, imag} */,
  {32'h3e26a82c, 32'h00000000} /* (12, 2, 13) {real, imag} */,
  {32'h3e33506b, 32'h00000000} /* (12, 2, 12) {real, imag} */,
  {32'h3e360e7f, 32'h00000000} /* (12, 2, 11) {real, imag} */,
  {32'h3d05e401, 32'h00000000} /* (12, 2, 10) {real, imag} */,
  {32'hbe62b734, 32'h00000000} /* (12, 2, 9) {real, imag} */,
  {32'hbe68f00d, 32'h00000000} /* (12, 2, 8) {real, imag} */,
  {32'h3e8ffdcb, 32'h00000000} /* (12, 2, 7) {real, imag} */,
  {32'hbc9fb323, 32'h00000000} /* (12, 2, 6) {real, imag} */,
  {32'hbf1e5b00, 32'h00000000} /* (12, 2, 5) {real, imag} */,
  {32'hbe641154, 32'h00000000} /* (12, 2, 4) {real, imag} */,
  {32'h3d985d34, 32'h00000000} /* (12, 2, 3) {real, imag} */,
  {32'hbe5e0fee, 32'h00000000} /* (12, 2, 2) {real, imag} */,
  {32'h3e3a0679, 32'h00000000} /* (12, 2, 1) {real, imag} */,
  {32'hbd2c0081, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'hbe35d51f, 32'h00000000} /* (12, 1, 15) {real, imag} */,
  {32'hbe999cd7, 32'h00000000} /* (12, 1, 14) {real, imag} */,
  {32'h3ea44330, 32'h00000000} /* (12, 1, 13) {real, imag} */,
  {32'h3db86706, 32'h00000000} /* (12, 1, 12) {real, imag} */,
  {32'h3e9fb8f3, 32'h00000000} /* (12, 1, 11) {real, imag} */,
  {32'h3e90bcaf, 32'h00000000} /* (12, 1, 10) {real, imag} */,
  {32'h3e256e91, 32'h00000000} /* (12, 1, 9) {real, imag} */,
  {32'h3e7d8a69, 32'h00000000} /* (12, 1, 8) {real, imag} */,
  {32'h3e449b96, 32'h00000000} /* (12, 1, 7) {real, imag} */,
  {32'hbe23087a, 32'h00000000} /* (12, 1, 6) {real, imag} */,
  {32'hbe22ef83, 32'h00000000} /* (12, 1, 5) {real, imag} */,
  {32'h3d5f4b20, 32'h00000000} /* (12, 1, 4) {real, imag} */,
  {32'hbe2025a3, 32'h00000000} /* (12, 1, 3) {real, imag} */,
  {32'hbdb1891a, 32'h00000000} /* (12, 1, 2) {real, imag} */,
  {32'hbd861767, 32'h00000000} /* (12, 1, 1) {real, imag} */,
  {32'hbc3cbebf, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'hbd1ad007, 32'h00000000} /* (12, 0, 15) {real, imag} */,
  {32'hbe073464, 32'h00000000} /* (12, 0, 14) {real, imag} */,
  {32'h3cf42678, 32'h00000000} /* (12, 0, 13) {real, imag} */,
  {32'hbbcf2c6c, 32'h00000000} /* (12, 0, 12) {real, imag} */,
  {32'hba86057f, 32'h00000000} /* (12, 0, 11) {real, imag} */,
  {32'h3d1c4466, 32'h00000000} /* (12, 0, 10) {real, imag} */,
  {32'h3e613307, 32'h00000000} /* (12, 0, 9) {real, imag} */,
  {32'h3e91a71b, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'h3c832a70, 32'h00000000} /* (12, 0, 7) {real, imag} */,
  {32'hbe66c764, 32'h00000000} /* (12, 0, 6) {real, imag} */,
  {32'hbd85690e, 32'h00000000} /* (12, 0, 5) {real, imag} */,
  {32'h3ea1b6a6, 32'h00000000} /* (12, 0, 4) {real, imag} */,
  {32'h3e8fa480, 32'h00000000} /* (12, 0, 3) {real, imag} */,
  {32'h3e802b55, 32'h00000000} /* (12, 0, 2) {real, imag} */,
  {32'h3da6bd24, 32'h00000000} /* (12, 0, 1) {real, imag} */,
  {32'h3e1de1a6, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h3e6bca48, 32'h00000000} /* (11, 15, 15) {real, imag} */,
  {32'h3dccc0b9, 32'h00000000} /* (11, 15, 14) {real, imag} */,
  {32'hbd95f6cf, 32'h00000000} /* (11, 15, 13) {real, imag} */,
  {32'h3db4be47, 32'h00000000} /* (11, 15, 12) {real, imag} */,
  {32'h3e47287e, 32'h00000000} /* (11, 15, 11) {real, imag} */,
  {32'hbd5e33cd, 32'h00000000} /* (11, 15, 10) {real, imag} */,
  {32'hbe8ad0d9, 32'h00000000} /* (11, 15, 9) {real, imag} */,
  {32'hbf52bf4e, 32'h00000000} /* (11, 15, 8) {real, imag} */,
  {32'hbe111e5e, 32'h00000000} /* (11, 15, 7) {real, imag} */,
  {32'h3e1e3fd7, 32'h00000000} /* (11, 15, 6) {real, imag} */,
  {32'h3dd04f1c, 32'h00000000} /* (11, 15, 5) {real, imag} */,
  {32'h3f066b8a, 32'h00000000} /* (11, 15, 4) {real, imag} */,
  {32'h3e9d0071, 32'h00000000} /* (11, 15, 3) {real, imag} */,
  {32'hbe6352f6, 32'h00000000} /* (11, 15, 2) {real, imag} */,
  {32'h3c528578, 32'h00000000} /* (11, 15, 1) {real, imag} */,
  {32'hbc14b343, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'h3ece9120, 32'h00000000} /* (11, 14, 15) {real, imag} */,
  {32'h3ec839bc, 32'h00000000} /* (11, 14, 14) {real, imag} */,
  {32'h3e37e102, 32'h00000000} /* (11, 14, 13) {real, imag} */,
  {32'hbe451ff4, 32'h00000000} /* (11, 14, 12) {real, imag} */,
  {32'h3e97224f, 32'h00000000} /* (11, 14, 11) {real, imag} */,
  {32'h3bbb9050, 32'h00000000} /* (11, 14, 10) {real, imag} */,
  {32'h3c09c41c, 32'h00000000} /* (11, 14, 9) {real, imag} */,
  {32'hbf008e1d, 32'h00000000} /* (11, 14, 8) {real, imag} */,
  {32'h3ee7da59, 32'h00000000} /* (11, 14, 7) {real, imag} */,
  {32'h3f061802, 32'h00000000} /* (11, 14, 6) {real, imag} */,
  {32'h3eebd47d, 32'h00000000} /* (11, 14, 5) {real, imag} */,
  {32'h3f11e8ff, 32'h00000000} /* (11, 14, 4) {real, imag} */,
  {32'h3eca0697, 32'h00000000} /* (11, 14, 3) {real, imag} */,
  {32'hbe73b46f, 32'h00000000} /* (11, 14, 2) {real, imag} */,
  {32'hbe330401, 32'h00000000} /* (11, 14, 1) {real, imag} */,
  {32'hbde48f2d, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'h3d89935c, 32'h00000000} /* (11, 13, 15) {real, imag} */,
  {32'h3f25dd02, 32'h00000000} /* (11, 13, 14) {real, imag} */,
  {32'h3e05c694, 32'h00000000} /* (11, 13, 13) {real, imag} */,
  {32'hbeadaad6, 32'h00000000} /* (11, 13, 12) {real, imag} */,
  {32'h3e0074b5, 32'h00000000} /* (11, 13, 11) {real, imag} */,
  {32'h3e541223, 32'h00000000} /* (11, 13, 10) {real, imag} */,
  {32'h3ea59bfd, 32'h00000000} /* (11, 13, 9) {real, imag} */,
  {32'h3e64e2d5, 32'h00000000} /* (11, 13, 8) {real, imag} */,
  {32'h3f7c8e9f, 32'h00000000} /* (11, 13, 7) {real, imag} */,
  {32'h3e7749c5, 32'h00000000} /* (11, 13, 6) {real, imag} */,
  {32'h3ddba8cd, 32'h00000000} /* (11, 13, 5) {real, imag} */,
  {32'h3f26ce66, 32'h00000000} /* (11, 13, 4) {real, imag} */,
  {32'h3e17f6d8, 32'h00000000} /* (11, 13, 3) {real, imag} */,
  {32'hbe78051f, 32'h00000000} /* (11, 13, 2) {real, imag} */,
  {32'h3e9ed536, 32'h00000000} /* (11, 13, 1) {real, imag} */,
  {32'h3da7c60c, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'hbcbbfa74, 32'h00000000} /* (11, 12, 15) {real, imag} */,
  {32'hbeae700e, 32'h00000000} /* (11, 12, 14) {real, imag} */,
  {32'hbeb48f9f, 32'h00000000} /* (11, 12, 13) {real, imag} */,
  {32'h3e9f4c63, 32'h00000000} /* (11, 12, 12) {real, imag} */,
  {32'h3f01e420, 32'h00000000} /* (11, 12, 11) {real, imag} */,
  {32'h3e17da66, 32'h00000000} /* (11, 12, 10) {real, imag} */,
  {32'hbddb0c30, 32'h00000000} /* (11, 12, 9) {real, imag} */,
  {32'hbe1add82, 32'h00000000} /* (11, 12, 8) {real, imag} */,
  {32'h3ea47019, 32'h00000000} /* (11, 12, 7) {real, imag} */,
  {32'hbd2651fa, 32'h00000000} /* (11, 12, 6) {real, imag} */,
  {32'hbda38f4c, 32'h00000000} /* (11, 12, 5) {real, imag} */,
  {32'h3f09a45f, 32'h00000000} /* (11, 12, 4) {real, imag} */,
  {32'h3e2dcb14, 32'h00000000} /* (11, 12, 3) {real, imag} */,
  {32'hbdfd7482, 32'h00000000} /* (11, 12, 2) {real, imag} */,
  {32'h3f0dd42b, 32'h00000000} /* (11, 12, 1) {real, imag} */,
  {32'h3f0bcd36, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'hbdc1a017, 32'h00000000} /* (11, 11, 15) {real, imag} */,
  {32'hbe9278fb, 32'h00000000} /* (11, 11, 14) {real, imag} */,
  {32'hbd3f7e70, 32'h00000000} /* (11, 11, 13) {real, imag} */,
  {32'h3e9fb8dc, 32'h00000000} /* (11, 11, 12) {real, imag} */,
  {32'h3ed09f5a, 32'h00000000} /* (11, 11, 11) {real, imag} */,
  {32'hbd6ad01e, 32'h00000000} /* (11, 11, 10) {real, imag} */,
  {32'hbd8288ec, 32'h00000000} /* (11, 11, 9) {real, imag} */,
  {32'hbe19c02c, 32'h00000000} /* (11, 11, 8) {real, imag} */,
  {32'h3eda3e23, 32'h00000000} /* (11, 11, 7) {real, imag} */,
  {32'h3ed99d04, 32'h00000000} /* (11, 11, 6) {real, imag} */,
  {32'h3ee7ec8d, 32'h00000000} /* (11, 11, 5) {real, imag} */,
  {32'h3ea1b0e0, 32'h00000000} /* (11, 11, 4) {real, imag} */,
  {32'h3dbca7e4, 32'h00000000} /* (11, 11, 3) {real, imag} */,
  {32'h3ea5a8b4, 32'h00000000} /* (11, 11, 2) {real, imag} */,
  {32'h3f1e60a2, 32'h00000000} /* (11, 11, 1) {real, imag} */,
  {32'h3ede8d92, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h3d4d5ae4, 32'h00000000} /* (11, 10, 15) {real, imag} */,
  {32'h3e100376, 32'h00000000} /* (11, 10, 14) {real, imag} */,
  {32'hbddc8874, 32'h00000000} /* (11, 10, 13) {real, imag} */,
  {32'h3e624d12, 32'h00000000} /* (11, 10, 12) {real, imag} */,
  {32'h3e023ef4, 32'h00000000} /* (11, 10, 11) {real, imag} */,
  {32'hbc2f456c, 32'h00000000} /* (11, 10, 10) {real, imag} */,
  {32'hbc1d4e6b, 32'h00000000} /* (11, 10, 9) {real, imag} */,
  {32'h3e456415, 32'h00000000} /* (11, 10, 8) {real, imag} */,
  {32'h3f83c1f1, 32'h00000000} /* (11, 10, 7) {real, imag} */,
  {32'h3eb3c349, 32'h00000000} /* (11, 10, 6) {real, imag} */,
  {32'h3f0a91f3, 32'h00000000} /* (11, 10, 5) {real, imag} */,
  {32'h3f2397f6, 32'h00000000} /* (11, 10, 4) {real, imag} */,
  {32'h3e50194e, 32'h00000000} /* (11, 10, 3) {real, imag} */,
  {32'h3ef68560, 32'h00000000} /* (11, 10, 2) {real, imag} */,
  {32'h3f3bc0c6, 32'h00000000} /* (11, 10, 1) {real, imag} */,
  {32'h3e354b62, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h3df5fe85, 32'h00000000} /* (11, 9, 15) {real, imag} */,
  {32'hbaebef55, 32'h00000000} /* (11, 9, 14) {real, imag} */,
  {32'hbe840eef, 32'h00000000} /* (11, 9, 13) {real, imag} */,
  {32'h3db9bd17, 32'h00000000} /* (11, 9, 12) {real, imag} */,
  {32'h3f0918c2, 32'h00000000} /* (11, 9, 11) {real, imag} */,
  {32'h3e8fba42, 32'h00000000} /* (11, 9, 10) {real, imag} */,
  {32'h3d020aa1, 32'h00000000} /* (11, 9, 9) {real, imag} */,
  {32'hbd16008c, 32'h00000000} /* (11, 9, 8) {real, imag} */,
  {32'h3f00649a, 32'h00000000} /* (11, 9, 7) {real, imag} */,
  {32'hbee3b772, 32'h00000000} /* (11, 9, 6) {real, imag} */,
  {32'hbf04fc4e, 32'h00000000} /* (11, 9, 5) {real, imag} */,
  {32'hbb3ac587, 32'h00000000} /* (11, 9, 4) {real, imag} */,
  {32'hbdd9fac1, 32'h00000000} /* (11, 9, 3) {real, imag} */,
  {32'h3de97bdf, 32'h00000000} /* (11, 9, 2) {real, imag} */,
  {32'h3f3e01f9, 32'h00000000} /* (11, 9, 1) {real, imag} */,
  {32'h3e0d84db, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h3eeb29a0, 32'h00000000} /* (11, 8, 15) {real, imag} */,
  {32'h3eed7920, 32'h00000000} /* (11, 8, 14) {real, imag} */,
  {32'hbe5fed74, 32'h00000000} /* (11, 8, 13) {real, imag} */,
  {32'hbf1f5bbc, 32'h00000000} /* (11, 8, 12) {real, imag} */,
  {32'h3e56996e, 32'h00000000} /* (11, 8, 11) {real, imag} */,
  {32'h3ce42837, 32'h00000000} /* (11, 8, 10) {real, imag} */,
  {32'h3e0df4a7, 32'h00000000} /* (11, 8, 9) {real, imag} */,
  {32'hbe7755c4, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'hbe5c7af5, 32'h00000000} /* (11, 8, 7) {real, imag} */,
  {32'hbf163780, 32'h00000000} /* (11, 8, 6) {real, imag} */,
  {32'hbee6cba1, 32'h00000000} /* (11, 8, 5) {real, imag} */,
  {32'hbe817bf3, 32'h00000000} /* (11, 8, 4) {real, imag} */,
  {32'hbf1f9d7d, 32'h00000000} /* (11, 8, 3) {real, imag} */,
  {32'hbedd5dbe, 32'h00000000} /* (11, 8, 2) {real, imag} */,
  {32'h3e2a0879, 32'h00000000} /* (11, 8, 1) {real, imag} */,
  {32'h3bae8f68, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h3e54af9b, 32'h00000000} /* (11, 7, 15) {real, imag} */,
  {32'h3e5278c8, 32'h00000000} /* (11, 7, 14) {real, imag} */,
  {32'hbf46bd16, 32'h00000000} /* (11, 7, 13) {real, imag} */,
  {32'hbec56559, 32'h00000000} /* (11, 7, 12) {real, imag} */,
  {32'h3ed7d14a, 32'h00000000} /* (11, 7, 11) {real, imag} */,
  {32'hbda780db, 32'h00000000} /* (11, 7, 10) {real, imag} */,
  {32'hbd5a8f1a, 32'h00000000} /* (11, 7, 9) {real, imag} */,
  {32'hbe16d298, 32'h00000000} /* (11, 7, 8) {real, imag} */,
  {32'h3db801b9, 32'h00000000} /* (11, 7, 7) {real, imag} */,
  {32'hbe7fd3c3, 32'h00000000} /* (11, 7, 6) {real, imag} */,
  {32'hbef18476, 32'h00000000} /* (11, 7, 5) {real, imag} */,
  {32'hbe50caf2, 32'h00000000} /* (11, 7, 4) {real, imag} */,
  {32'h3e7e6b76, 32'h00000000} /* (11, 7, 3) {real, imag} */,
  {32'h3dd081ca, 32'h00000000} /* (11, 7, 2) {real, imag} */,
  {32'hbe6242e8, 32'h00000000} /* (11, 7, 1) {real, imag} */,
  {32'h3c5b724a, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'hbd98ae69, 32'h00000000} /* (11, 6, 15) {real, imag} */,
  {32'h3d2923be, 32'h00000000} /* (11, 6, 14) {real, imag} */,
  {32'h3db87237, 32'h00000000} /* (11, 6, 13) {real, imag} */,
  {32'h3e130467, 32'h00000000} /* (11, 6, 12) {real, imag} */,
  {32'h3e3feb06, 32'h00000000} /* (11, 6, 11) {real, imag} */,
  {32'hbe7f7971, 32'h00000000} /* (11, 6, 10) {real, imag} */,
  {32'h3f316c64, 32'h00000000} /* (11, 6, 9) {real, imag} */,
  {32'h3ef4a8d4, 32'h00000000} /* (11, 6, 8) {real, imag} */,
  {32'h3f6cab7d, 32'h00000000} /* (11, 6, 7) {real, imag} */,
  {32'h3eb304a4, 32'h00000000} /* (11, 6, 6) {real, imag} */,
  {32'hbe952af8, 32'h00000000} /* (11, 6, 5) {real, imag} */,
  {32'hbe7449e4, 32'h00000000} /* (11, 6, 4) {real, imag} */,
  {32'h3eb3dd20, 32'h00000000} /* (11, 6, 3) {real, imag} */,
  {32'hbe1dc838, 32'h00000000} /* (11, 6, 2) {real, imag} */,
  {32'hbf30b6fc, 32'h00000000} /* (11, 6, 1) {real, imag} */,
  {32'h3d5e400e, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h3e2efa93, 32'h00000000} /* (11, 5, 15) {real, imag} */,
  {32'h3e4f1c07, 32'h00000000} /* (11, 5, 14) {real, imag} */,
  {32'hbdb555e5, 32'h00000000} /* (11, 5, 13) {real, imag} */,
  {32'hbe8a74a9, 32'h00000000} /* (11, 5, 12) {real, imag} */,
  {32'hbed44bde, 32'h00000000} /* (11, 5, 11) {real, imag} */,
  {32'hbee1b6ca, 32'h00000000} /* (11, 5, 10) {real, imag} */,
  {32'h3f3bda3f, 32'h00000000} /* (11, 5, 9) {real, imag} */,
  {32'h3ef8e7ca, 32'h00000000} /* (11, 5, 8) {real, imag} */,
  {32'h3f6c8ce2, 32'h00000000} /* (11, 5, 7) {real, imag} */,
  {32'h3e82de9e, 32'h00000000} /* (11, 5, 6) {real, imag} */,
  {32'hbe0ba919, 32'h00000000} /* (11, 5, 5) {real, imag} */,
  {32'h3edd30fb, 32'h00000000} /* (11, 5, 4) {real, imag} */,
  {32'h3eeddb2a, 32'h00000000} /* (11, 5, 3) {real, imag} */,
  {32'h3e8e9351, 32'h00000000} /* (11, 5, 2) {real, imag} */,
  {32'h3d2eeab8, 32'h00000000} /* (11, 5, 1) {real, imag} */,
  {32'h3e466ffa, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h3ec2b81f, 32'h00000000} /* (11, 4, 15) {real, imag} */,
  {32'h3e9ed267, 32'h00000000} /* (11, 4, 14) {real, imag} */,
  {32'hbeb6aa96, 32'h00000000} /* (11, 4, 13) {real, imag} */,
  {32'hbefb32d0, 32'h00000000} /* (11, 4, 12) {real, imag} */,
  {32'hbec4547c, 32'h00000000} /* (11, 4, 11) {real, imag} */,
  {32'hbeda940e, 32'h00000000} /* (11, 4, 10) {real, imag} */,
  {32'hbb80d18a, 32'h00000000} /* (11, 4, 9) {real, imag} */,
  {32'h3e530c86, 32'h00000000} /* (11, 4, 8) {real, imag} */,
  {32'h3eb92778, 32'h00000000} /* (11, 4, 7) {real, imag} */,
  {32'h3d01476d, 32'h00000000} /* (11, 4, 6) {real, imag} */,
  {32'hbe1b98fd, 32'h00000000} /* (11, 4, 5) {real, imag} */,
  {32'h3ec0b97b, 32'h00000000} /* (11, 4, 4) {real, imag} */,
  {32'h3f459f0c, 32'h00000000} /* (11, 4, 3) {real, imag} */,
  {32'h3ef1ca6c, 32'h00000000} /* (11, 4, 2) {real, imag} */,
  {32'h3ec14077, 32'h00000000} /* (11, 4, 1) {real, imag} */,
  {32'h3e9d7a0a, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h3d1b7c19, 32'h00000000} /* (11, 3, 15) {real, imag} */,
  {32'hbe8b12fd, 32'h00000000} /* (11, 3, 14) {real, imag} */,
  {32'hbed491f1, 32'h00000000} /* (11, 3, 13) {real, imag} */,
  {32'hbed0292d, 32'h00000000} /* (11, 3, 12) {real, imag} */,
  {32'hbbb30685, 32'h00000000} /* (11, 3, 11) {real, imag} */,
  {32'hbe624f2e, 32'h00000000} /* (11, 3, 10) {real, imag} */,
  {32'hbf049a2c, 32'h00000000} /* (11, 3, 9) {real, imag} */,
  {32'hbdf1a2af, 32'h00000000} /* (11, 3, 8) {real, imag} */,
  {32'h3bd74b70, 32'h00000000} /* (11, 3, 7) {real, imag} */,
  {32'hbd0a4174, 32'h00000000} /* (11, 3, 6) {real, imag} */,
  {32'hbec48aa0, 32'h00000000} /* (11, 3, 5) {real, imag} */,
  {32'hbe445314, 32'h00000000} /* (11, 3, 4) {real, imag} */,
  {32'h3f32b6ee, 32'h00000000} /* (11, 3, 3) {real, imag} */,
  {32'h3e379c58, 32'h00000000} /* (11, 3, 2) {real, imag} */,
  {32'hbda7f09e, 32'h00000000} /* (11, 3, 1) {real, imag} */,
  {32'hbb72d44c, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'hbe485d41, 32'h00000000} /* (11, 2, 15) {real, imag} */,
  {32'hbf35ce91, 32'h00000000} /* (11, 2, 14) {real, imag} */,
  {32'hbe843298, 32'h00000000} /* (11, 2, 13) {real, imag} */,
  {32'hbe112e0b, 32'h00000000} /* (11, 2, 12) {real, imag} */,
  {32'h3ef544a0, 32'h00000000} /* (11, 2, 11) {real, imag} */,
  {32'h3e3e50a3, 32'h00000000} /* (11, 2, 10) {real, imag} */,
  {32'hbec93d47, 32'h00000000} /* (11, 2, 9) {real, imag} */,
  {32'hbe076acb, 32'h00000000} /* (11, 2, 8) {real, imag} */,
  {32'h3e29878d, 32'h00000000} /* (11, 2, 7) {real, imag} */,
  {32'hbc9e2612, 32'h00000000} /* (11, 2, 6) {real, imag} */,
  {32'hbf1f57bd, 32'h00000000} /* (11, 2, 5) {real, imag} */,
  {32'hbeb499a7, 32'h00000000} /* (11, 2, 4) {real, imag} */,
  {32'hbe0d8ab8, 32'h00000000} /* (11, 2, 3) {real, imag} */,
  {32'hbf1b764e, 32'h00000000} /* (11, 2, 2) {real, imag} */,
  {32'hbebe5d30, 32'h00000000} /* (11, 2, 1) {real, imag} */,
  {32'hbdc17d85, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h3db31231, 32'h00000000} /* (11, 1, 15) {real, imag} */,
  {32'hbd3bd474, 32'h00000000} /* (11, 1, 14) {real, imag} */,
  {32'h3e0c7164, 32'h00000000} /* (11, 1, 13) {real, imag} */,
  {32'hbe56b5e6, 32'h00000000} /* (11, 1, 12) {real, imag} */,
  {32'h3e38d1bd, 32'h00000000} /* (11, 1, 11) {real, imag} */,
  {32'h3ef8ba29, 32'h00000000} /* (11, 1, 10) {real, imag} */,
  {32'h3d6f5dec, 32'h00000000} /* (11, 1, 9) {real, imag} */,
  {32'h3e184c60, 32'h00000000} /* (11, 1, 8) {real, imag} */,
  {32'h3effbe59, 32'h00000000} /* (11, 1, 7) {real, imag} */,
  {32'h3df37637, 32'h00000000} /* (11, 1, 6) {real, imag} */,
  {32'hbd77a68a, 32'h00000000} /* (11, 1, 5) {real, imag} */,
  {32'h3f0b6da4, 32'h00000000} /* (11, 1, 4) {real, imag} */,
  {32'h3c17d72c, 32'h00000000} /* (11, 1, 3) {real, imag} */,
  {32'hbe9ed469, 32'h00000000} /* (11, 1, 2) {real, imag} */,
  {32'hbcb99e6a, 32'h00000000} /* (11, 1, 1) {real, imag} */,
  {32'h3e5f7521, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h3d9f35cb, 32'h00000000} /* (11, 0, 15) {real, imag} */,
  {32'hbc2a7d6c, 32'h00000000} /* (11, 0, 14) {real, imag} */,
  {32'hbdbb78fa, 32'h00000000} /* (11, 0, 13) {real, imag} */,
  {32'hbe96c157, 32'h00000000} /* (11, 0, 12) {real, imag} */,
  {32'hbe3a015f, 32'h00000000} /* (11, 0, 11) {real, imag} */,
  {32'h3e19f5f5, 32'h00000000} /* (11, 0, 10) {real, imag} */,
  {32'hbc516194, 32'h00000000} /* (11, 0, 9) {real, imag} */,
  {32'hbde33724, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'h3e5b9ec1, 32'h00000000} /* (11, 0, 7) {real, imag} */,
  {32'hbe474c44, 32'h00000000} /* (11, 0, 6) {real, imag} */,
  {32'hbe808ecc, 32'h00000000} /* (11, 0, 5) {real, imag} */,
  {32'h3eed701f, 32'h00000000} /* (11, 0, 4) {real, imag} */,
  {32'h3e4cf990, 32'h00000000} /* (11, 0, 3) {real, imag} */,
  {32'h3e391cf5, 32'h00000000} /* (11, 0, 2) {real, imag} */,
  {32'h3e4d8d79, 32'h00000000} /* (11, 0, 1) {real, imag} */,
  {32'h3e943ba5, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h3e1d9d72, 32'h00000000} /* (10, 15, 15) {real, imag} */,
  {32'h3e1fcf32, 32'h00000000} /* (10, 15, 14) {real, imag} */,
  {32'h3e24b155, 32'h00000000} /* (10, 15, 13) {real, imag} */,
  {32'h3e5fa56a, 32'h00000000} /* (10, 15, 12) {real, imag} */,
  {32'h3e64315c, 32'h00000000} /* (10, 15, 11) {real, imag} */,
  {32'h3dd2770c, 32'h00000000} /* (10, 15, 10) {real, imag} */,
  {32'hbebd92ce, 32'h00000000} /* (10, 15, 9) {real, imag} */,
  {32'hbf188025, 32'h00000000} /* (10, 15, 8) {real, imag} */,
  {32'h3e095aea, 32'h00000000} /* (10, 15, 7) {real, imag} */,
  {32'h3e52eec6, 32'h00000000} /* (10, 15, 6) {real, imag} */,
  {32'h3e2d0bdd, 32'h00000000} /* (10, 15, 5) {real, imag} */,
  {32'hbca4b047, 32'h00000000} /* (10, 15, 4) {real, imag} */,
  {32'hbecbab46, 32'h00000000} /* (10, 15, 3) {real, imag} */,
  {32'hbdaf0c9f, 32'h00000000} /* (10, 15, 2) {real, imag} */,
  {32'h3e38c770, 32'h00000000} /* (10, 15, 1) {real, imag} */,
  {32'h3d55cd97, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'h3ed4a073, 32'h00000000} /* (10, 14, 15) {real, imag} */,
  {32'h3f621d52, 32'h00000000} /* (10, 14, 14) {real, imag} */,
  {32'h3f56925d, 32'h00000000} /* (10, 14, 13) {real, imag} */,
  {32'h3f04b19d, 32'h00000000} /* (10, 14, 12) {real, imag} */,
  {32'h3e964867, 32'h00000000} /* (10, 14, 11) {real, imag} */,
  {32'hbd63154a, 32'h00000000} /* (10, 14, 10) {real, imag} */,
  {32'hbf02b0f4, 32'h00000000} /* (10, 14, 9) {real, imag} */,
  {32'hbf13514e, 32'h00000000} /* (10, 14, 8) {real, imag} */,
  {32'h3e97b790, 32'h00000000} /* (10, 14, 7) {real, imag} */,
  {32'h3f016dfd, 32'h00000000} /* (10, 14, 6) {real, imag} */,
  {32'h3f24dda8, 32'h00000000} /* (10, 14, 5) {real, imag} */,
  {32'h3ca067e8, 32'h00000000} /* (10, 14, 4) {real, imag} */,
  {32'hbf1a4867, 32'h00000000} /* (10, 14, 3) {real, imag} */,
  {32'hbf22cd92, 32'h00000000} /* (10, 14, 2) {real, imag} */,
  {32'h3aa9f320, 32'h00000000} /* (10, 14, 1) {real, imag} */,
  {32'h3cd83800, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'h3e084e6f, 32'h00000000} /* (10, 13, 15) {real, imag} */,
  {32'h3f477853, 32'h00000000} /* (10, 13, 14) {real, imag} */,
  {32'h3ebd87e8, 32'h00000000} /* (10, 13, 13) {real, imag} */,
  {32'h3e543af3, 32'h00000000} /* (10, 13, 12) {real, imag} */,
  {32'h3ec46e5b, 32'h00000000} /* (10, 13, 11) {real, imag} */,
  {32'h3c5dd136, 32'h00000000} /* (10, 13, 10) {real, imag} */,
  {32'hbe26b698, 32'h00000000} /* (10, 13, 9) {real, imag} */,
  {32'hbd9070c8, 32'h00000000} /* (10, 13, 8) {real, imag} */,
  {32'h3f187f51, 32'h00000000} /* (10, 13, 7) {real, imag} */,
  {32'h3f2112c1, 32'h00000000} /* (10, 13, 6) {real, imag} */,
  {32'h3e1ca4d9, 32'h00000000} /* (10, 13, 5) {real, imag} */,
  {32'hbd00684d, 32'h00000000} /* (10, 13, 4) {real, imag} */,
  {32'hbd9fbaec, 32'h00000000} /* (10, 13, 3) {real, imag} */,
  {32'hbe6c39ee, 32'h00000000} /* (10, 13, 2) {real, imag} */,
  {32'h3efccbe0, 32'h00000000} /* (10, 13, 1) {real, imag} */,
  {32'h3e526632, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hbe11bcc6, 32'h00000000} /* (10, 12, 15) {real, imag} */,
  {32'hbea7761e, 32'h00000000} /* (10, 12, 14) {real, imag} */,
  {32'hbf154511, 32'h00000000} /* (10, 12, 13) {real, imag} */,
  {32'hbead18c4, 32'h00000000} /* (10, 12, 12) {real, imag} */,
  {32'hbd4197fc, 32'h00000000} /* (10, 12, 11) {real, imag} */,
  {32'hbe458197, 32'h00000000} /* (10, 12, 10) {real, imag} */,
  {32'h3ef05161, 32'h00000000} /* (10, 12, 9) {real, imag} */,
  {32'h3ef30c38, 32'h00000000} /* (10, 12, 8) {real, imag} */,
  {32'h3f2eb45e, 32'h00000000} /* (10, 12, 7) {real, imag} */,
  {32'h3f396a5f, 32'h00000000} /* (10, 12, 6) {real, imag} */,
  {32'h3e42a706, 32'h00000000} /* (10, 12, 5) {real, imag} */,
  {32'h3e5a51c5, 32'h00000000} /* (10, 12, 4) {real, imag} */,
  {32'hbdccd479, 32'h00000000} /* (10, 12, 3) {real, imag} */,
  {32'hbe2d6b4c, 32'h00000000} /* (10, 12, 2) {real, imag} */,
  {32'h3ed7239a, 32'h00000000} /* (10, 12, 1) {real, imag} */,
  {32'h3e86a6d0, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hbeaa47f1, 32'h00000000} /* (10, 11, 15) {real, imag} */,
  {32'hbdc391d1, 32'h00000000} /* (10, 11, 14) {real, imag} */,
  {32'hbe52f18e, 32'h00000000} /* (10, 11, 13) {real, imag} */,
  {32'hbe13e2a4, 32'h00000000} /* (10, 11, 12) {real, imag} */,
  {32'hbe03d1ef, 32'h00000000} /* (10, 11, 11) {real, imag} */,
  {32'h3d5aaeac, 32'h00000000} /* (10, 11, 10) {real, imag} */,
  {32'h3f7fd080, 32'h00000000} /* (10, 11, 9) {real, imag} */,
  {32'h3ef3db87, 32'h00000000} /* (10, 11, 8) {real, imag} */,
  {32'h3ee3985b, 32'h00000000} /* (10, 11, 7) {real, imag} */,
  {32'h3f291f1c, 32'h00000000} /* (10, 11, 6) {real, imag} */,
  {32'h3f4a14e1, 32'h00000000} /* (10, 11, 5) {real, imag} */,
  {32'h3f4a99df, 32'h00000000} /* (10, 11, 4) {real, imag} */,
  {32'h3e2ae5b9, 32'h00000000} /* (10, 11, 3) {real, imag} */,
  {32'h3ce6d550, 32'h00000000} /* (10, 11, 2) {real, imag} */,
  {32'h3d443450, 32'h00000000} /* (10, 11, 1) {real, imag} */,
  {32'hbd4085d0, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h3e01dd33, 32'h00000000} /* (10, 10, 15) {real, imag} */,
  {32'h3f03dd13, 32'h00000000} /* (10, 10, 14) {real, imag} */,
  {32'hbd6317f0, 32'h00000000} /* (10, 10, 13) {real, imag} */,
  {32'h3d64d882, 32'h00000000} /* (10, 10, 12) {real, imag} */,
  {32'hbea50310, 32'h00000000} /* (10, 10, 11) {real, imag} */,
  {32'hbeaa853c, 32'h00000000} /* (10, 10, 10) {real, imag} */,
  {32'h3ed83dee, 32'h00000000} /* (10, 10, 9) {real, imag} */,
  {32'h3f020f49, 32'h00000000} /* (10, 10, 8) {real, imag} */,
  {32'h3f3f8dea, 32'h00000000} /* (10, 10, 7) {real, imag} */,
  {32'h3e861390, 32'h00000000} /* (10, 10, 6) {real, imag} */,
  {32'h3edbd7ac, 32'h00000000} /* (10, 10, 5) {real, imag} */,
  {32'h3f2f711b, 32'h00000000} /* (10, 10, 4) {real, imag} */,
  {32'h3e9f404a, 32'h00000000} /* (10, 10, 3) {real, imag} */,
  {32'h3f229992, 32'h00000000} /* (10, 10, 2) {real, imag} */,
  {32'h3f034500, 32'h00000000} /* (10, 10, 1) {real, imag} */,
  {32'h3dc73eb2, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h3e9e82c5, 32'h00000000} /* (10, 9, 15) {real, imag} */,
  {32'h3f0a133b, 32'h00000000} /* (10, 9, 14) {real, imag} */,
  {32'h3d898e52, 32'h00000000} /* (10, 9, 13) {real, imag} */,
  {32'hbe46e7ba, 32'h00000000} /* (10, 9, 12) {real, imag} */,
  {32'h3d44a9ab, 32'h00000000} /* (10, 9, 11) {real, imag} */,
  {32'hbb838434, 32'h00000000} /* (10, 9, 10) {real, imag} */,
  {32'h3e958b1e, 32'h00000000} /* (10, 9, 9) {real, imag} */,
  {32'h3ec0d887, 32'h00000000} /* (10, 9, 8) {real, imag} */,
  {32'h3ef76980, 32'h00000000} /* (10, 9, 7) {real, imag} */,
  {32'hbf2681c9, 32'h00000000} /* (10, 9, 6) {real, imag} */,
  {32'hbf33e87f, 32'h00000000} /* (10, 9, 5) {real, imag} */,
  {32'hbe374a62, 32'h00000000} /* (10, 9, 4) {real, imag} */,
  {32'h3e30e75e, 32'h00000000} /* (10, 9, 3) {real, imag} */,
  {32'h3f06100e, 32'h00000000} /* (10, 9, 2) {real, imag} */,
  {32'h3f35af66, 32'h00000000} /* (10, 9, 1) {real, imag} */,
  {32'h3ee35b54, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h3f051b28, 32'h00000000} /* (10, 8, 15) {real, imag} */,
  {32'h3f4bfb89, 32'h00000000} /* (10, 8, 14) {real, imag} */,
  {32'h3ee2ee28, 32'h00000000} /* (10, 8, 13) {real, imag} */,
  {32'hbe3da0d7, 32'h00000000} /* (10, 8, 12) {real, imag} */,
  {32'h3e5b391f, 32'h00000000} /* (10, 8, 11) {real, imag} */,
  {32'h3db97955, 32'h00000000} /* (10, 8, 10) {real, imag} */,
  {32'h3edbb2f6, 32'h00000000} /* (10, 8, 9) {real, imag} */,
  {32'h3ebd16b8, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'h3eaf130a, 32'h00000000} /* (10, 8, 7) {real, imag} */,
  {32'hbf42d835, 32'h00000000} /* (10, 8, 6) {real, imag} */,
  {32'hbf144f33, 32'h00000000} /* (10, 8, 5) {real, imag} */,
  {32'hbe73add8, 32'h00000000} /* (10, 8, 4) {real, imag} */,
  {32'hbe99f355, 32'h00000000} /* (10, 8, 3) {real, imag} */,
  {32'hbdeb484a, 32'h00000000} /* (10, 8, 2) {real, imag} */,
  {32'hbd0a1d99, 32'h00000000} /* (10, 8, 1) {real, imag} */,
  {32'hbe4e58e1, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h3f273cb9, 32'h00000000} /* (10, 7, 15) {real, imag} */,
  {32'h3f80c47f, 32'h00000000} /* (10, 7, 14) {real, imag} */,
  {32'h3ec560c2, 32'h00000000} /* (10, 7, 13) {real, imag} */,
  {32'h3c00cdba, 32'h00000000} /* (10, 7, 12) {real, imag} */,
  {32'h3be87888, 32'h00000000} /* (10, 7, 11) {real, imag} */,
  {32'hbe9fcf9c, 32'h00000000} /* (10, 7, 10) {real, imag} */,
  {32'hbe475412, 32'h00000000} /* (10, 7, 9) {real, imag} */,
  {32'hbdcedec7, 32'h00000000} /* (10, 7, 8) {real, imag} */,
  {32'h3e475431, 32'h00000000} /* (10, 7, 7) {real, imag} */,
  {32'hbf024248, 32'h00000000} /* (10, 7, 6) {real, imag} */,
  {32'hbe7d2322, 32'h00000000} /* (10, 7, 5) {real, imag} */,
  {32'h3eaa6fd6, 32'h00000000} /* (10, 7, 4) {real, imag} */,
  {32'h3ef57000, 32'h00000000} /* (10, 7, 3) {real, imag} */,
  {32'h3e66ab74, 32'h00000000} /* (10, 7, 2) {real, imag} */,
  {32'hbeeb4741, 32'h00000000} /* (10, 7, 1) {real, imag} */,
  {32'hbe19aebc, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h3ec27e37, 32'h00000000} /* (10, 6, 15) {real, imag} */,
  {32'h3ea0f033, 32'h00000000} /* (10, 6, 14) {real, imag} */,
  {32'h3e9a5860, 32'h00000000} /* (10, 6, 13) {real, imag} */,
  {32'h3ee70c1b, 32'h00000000} /* (10, 6, 12) {real, imag} */,
  {32'hbddbab9c, 32'h00000000} /* (10, 6, 11) {real, imag} */,
  {32'hbea0aaa0, 32'h00000000} /* (10, 6, 10) {real, imag} */,
  {32'h3e72cd95, 32'h00000000} /* (10, 6, 9) {real, imag} */,
  {32'hbe7aa0cf, 32'h00000000} /* (10, 6, 8) {real, imag} */,
  {32'hbe1af8ad, 32'h00000000} /* (10, 6, 7) {real, imag} */,
  {32'h3db49e3d, 32'h00000000} /* (10, 6, 6) {real, imag} */,
  {32'h3e56fd9b, 32'h00000000} /* (10, 6, 5) {real, imag} */,
  {32'h3ed810e8, 32'h00000000} /* (10, 6, 4) {real, imag} */,
  {32'h3e048c7c, 32'h00000000} /* (10, 6, 3) {real, imag} */,
  {32'hbed813b4, 32'h00000000} /* (10, 6, 2) {real, imag} */,
  {32'hbf0ee6b5, 32'h00000000} /* (10, 6, 1) {real, imag} */,
  {32'h3e2a4749, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h3e3f77a5, 32'h00000000} /* (10, 5, 15) {real, imag} */,
  {32'h3e012278, 32'h00000000} /* (10, 5, 14) {real, imag} */,
  {32'hbe3e875a, 32'h00000000} /* (10, 5, 13) {real, imag} */,
  {32'hbe235e0a, 32'h00000000} /* (10, 5, 12) {real, imag} */,
  {32'hbe1c3054, 32'h00000000} /* (10, 5, 11) {real, imag} */,
  {32'hbf0f832a, 32'h00000000} /* (10, 5, 10) {real, imag} */,
  {32'h3dbb112b, 32'h00000000} /* (10, 5, 9) {real, imag} */,
  {32'hbdb6921f, 32'h00000000} /* (10, 5, 8) {real, imag} */,
  {32'hbb9bba1e, 32'h00000000} /* (10, 5, 7) {real, imag} */,
  {32'h3ea418fb, 32'h00000000} /* (10, 5, 6) {real, imag} */,
  {32'h3f296169, 32'h00000000} /* (10, 5, 5) {real, imag} */,
  {32'h3ec497e4, 32'h00000000} /* (10, 5, 4) {real, imag} */,
  {32'hbe8bf156, 32'h00000000} /* (10, 5, 3) {real, imag} */,
  {32'hbeea2315, 32'h00000000} /* (10, 5, 2) {real, imag} */,
  {32'hbecb4569, 32'h00000000} /* (10, 5, 1) {real, imag} */,
  {32'h3d969e42, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h3d7b7437, 32'h00000000} /* (10, 4, 15) {real, imag} */,
  {32'h3d99de34, 32'h00000000} /* (10, 4, 14) {real, imag} */,
  {32'hbe226125, 32'h00000000} /* (10, 4, 13) {real, imag} */,
  {32'hbf161d82, 32'h00000000} /* (10, 4, 12) {real, imag} */,
  {32'hbe25aec3, 32'h00000000} /* (10, 4, 11) {real, imag} */,
  {32'hbf0bbdd3, 32'h00000000} /* (10, 4, 10) {real, imag} */,
  {32'hbea1ba90, 32'h00000000} /* (10, 4, 9) {real, imag} */,
  {32'hbe064166, 32'h00000000} /* (10, 4, 8) {real, imag} */,
  {32'hbe963051, 32'h00000000} /* (10, 4, 7) {real, imag} */,
  {32'h3e4f387b, 32'h00000000} /* (10, 4, 6) {real, imag} */,
  {32'h3e3a247e, 32'h00000000} /* (10, 4, 5) {real, imag} */,
  {32'h3e41803b, 32'h00000000} /* (10, 4, 4) {real, imag} */,
  {32'h3ec551c3, 32'h00000000} /* (10, 4, 3) {real, imag} */,
  {32'h3eb1db81, 32'h00000000} /* (10, 4, 2) {real, imag} */,
  {32'h3e64ee9b, 32'h00000000} /* (10, 4, 1) {real, imag} */,
  {32'h3ec0a3f7, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'hbedd366c, 32'h00000000} /* (10, 3, 15) {real, imag} */,
  {32'hbef9fb21, 32'h00000000} /* (10, 3, 14) {real, imag} */,
  {32'hbe9154cb, 32'h00000000} /* (10, 3, 13) {real, imag} */,
  {32'hbf235893, 32'h00000000} /* (10, 3, 12) {real, imag} */,
  {32'hbe18430b, 32'h00000000} /* (10, 3, 11) {real, imag} */,
  {32'hbd63b2bd, 32'h00000000} /* (10, 3, 10) {real, imag} */,
  {32'hbd53d825, 32'h00000000} /* (10, 3, 9) {real, imag} */,
  {32'h3ea73d7f, 32'h00000000} /* (10, 3, 8) {real, imag} */,
  {32'h3b8c9958, 32'h00000000} /* (10, 3, 7) {real, imag} */,
  {32'h3dca5ee9, 32'h00000000} /* (10, 3, 6) {real, imag} */,
  {32'hbcfcfce0, 32'h00000000} /* (10, 3, 5) {real, imag} */,
  {32'h3d66e3f9, 32'h00000000} /* (10, 3, 4) {real, imag} */,
  {32'h3ebeba2b, 32'h00000000} /* (10, 3, 3) {real, imag} */,
  {32'h3e5e50d4, 32'h00000000} /* (10, 3, 2) {real, imag} */,
  {32'h3e47c063, 32'h00000000} /* (10, 3, 1) {real, imag} */,
  {32'h3e49c8a9, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'hbed70f24, 32'h00000000} /* (10, 2, 15) {real, imag} */,
  {32'hbf3322db, 32'h00000000} /* (10, 2, 14) {real, imag} */,
  {32'hbe9c1c5c, 32'h00000000} /* (10, 2, 13) {real, imag} */,
  {32'hbe91cb5c, 32'h00000000} /* (10, 2, 12) {real, imag} */,
  {32'h3e899844, 32'h00000000} /* (10, 2, 11) {real, imag} */,
  {32'h3e7d7191, 32'h00000000} /* (10, 2, 10) {real, imag} */,
  {32'hbe7daf0a, 32'h00000000} /* (10, 2, 9) {real, imag} */,
  {32'h3ec98d6b, 32'h00000000} /* (10, 2, 8) {real, imag} */,
  {32'h3f1aad66, 32'h00000000} /* (10, 2, 7) {real, imag} */,
  {32'h3e377617, 32'h00000000} /* (10, 2, 6) {real, imag} */,
  {32'hbd67ced4, 32'h00000000} /* (10, 2, 5) {real, imag} */,
  {32'h3e2fdb5b, 32'h00000000} /* (10, 2, 4) {real, imag} */,
  {32'hbd33b520, 32'h00000000} /* (10, 2, 3) {real, imag} */,
  {32'hbeb1fec4, 32'h00000000} /* (10, 2, 2) {real, imag} */,
  {32'hbe7091f3, 32'h00000000} /* (10, 2, 1) {real, imag} */,
  {32'h3da2306b, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h3d971daa, 32'h00000000} /* (10, 1, 15) {real, imag} */,
  {32'hbdef8eff, 32'h00000000} /* (10, 1, 14) {real, imag} */,
  {32'hbd382803, 32'h00000000} /* (10, 1, 13) {real, imag} */,
  {32'hbd3a277d, 32'h00000000} /* (10, 1, 12) {real, imag} */,
  {32'h3f126bda, 32'h00000000} /* (10, 1, 11) {real, imag} */,
  {32'h3ef477f7, 32'h00000000} /* (10, 1, 10) {real, imag} */,
  {32'hbdb75030, 32'h00000000} /* (10, 1, 9) {real, imag} */,
  {32'h3dd25f46, 32'h00000000} /* (10, 1, 8) {real, imag} */,
  {32'h3ec9e806, 32'h00000000} /* (10, 1, 7) {real, imag} */,
  {32'h3e221cf2, 32'h00000000} /* (10, 1, 6) {real, imag} */,
  {32'hbe15e905, 32'h00000000} /* (10, 1, 5) {real, imag} */,
  {32'h3f5623ad, 32'h00000000} /* (10, 1, 4) {real, imag} */,
  {32'h3eaa3a48, 32'h00000000} /* (10, 1, 3) {real, imag} */,
  {32'hbec34501, 32'h00000000} /* (10, 1, 2) {real, imag} */,
  {32'h3e9a2dea, 32'h00000000} /* (10, 1, 1) {real, imag} */,
  {32'h3f1548ed, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h3e8d4635, 32'h00000000} /* (10, 0, 15) {real, imag} */,
  {32'h3dd14b9b, 32'h00000000} /* (10, 0, 14) {real, imag} */,
  {32'h3de97696, 32'h00000000} /* (10, 0, 13) {real, imag} */,
  {32'h3e30e455, 32'h00000000} /* (10, 0, 12) {real, imag} */,
  {32'h3eeed216, 32'h00000000} /* (10, 0, 11) {real, imag} */,
  {32'h3ed11526, 32'h00000000} /* (10, 0, 10) {real, imag} */,
  {32'hbe44bcd4, 32'h00000000} /* (10, 0, 9) {real, imag} */,
  {32'hbeb3834a, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'h3dc610e1, 32'h00000000} /* (10, 0, 7) {real, imag} */,
  {32'hbe30a35e, 32'h00000000} /* (10, 0, 6) {real, imag} */,
  {32'hbea6c019, 32'h00000000} /* (10, 0, 5) {real, imag} */,
  {32'h3e98f525, 32'h00000000} /* (10, 0, 4) {real, imag} */,
  {32'h3dcfa055, 32'h00000000} /* (10, 0, 3) {real, imag} */,
  {32'hbe3bf6ea, 32'h00000000} /* (10, 0, 2) {real, imag} */,
  {32'h3e825a45, 32'h00000000} /* (10, 0, 1) {real, imag} */,
  {32'h3ee3f79d, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h3d916460, 32'h00000000} /* (9, 15, 15) {real, imag} */,
  {32'h3dec735c, 32'h00000000} /* (9, 15, 14) {real, imag} */,
  {32'h3deb6b60, 32'h00000000} /* (9, 15, 13) {real, imag} */,
  {32'h3ecb23dd, 32'h00000000} /* (9, 15, 12) {real, imag} */,
  {32'h3e5e2bee, 32'h00000000} /* (9, 15, 11) {real, imag} */,
  {32'h3c0082dc, 32'h00000000} /* (9, 15, 10) {real, imag} */,
  {32'hbe62e1aa, 32'h00000000} /* (9, 15, 9) {real, imag} */,
  {32'hbecc48a1, 32'h00000000} /* (9, 15, 8) {real, imag} */,
  {32'hbd2c2136, 32'h00000000} /* (9, 15, 7) {real, imag} */,
  {32'h3d22816e, 32'h00000000} /* (9, 15, 6) {real, imag} */,
  {32'h3e135513, 32'h00000000} /* (9, 15, 5) {real, imag} */,
  {32'hbdccc528, 32'h00000000} /* (9, 15, 4) {real, imag} */,
  {32'hbd93e0bc, 32'h00000000} /* (9, 15, 3) {real, imag} */,
  {32'h3e95ff2c, 32'h00000000} /* (9, 15, 2) {real, imag} */,
  {32'h3e17aed9, 32'h00000000} /* (9, 15, 1) {real, imag} */,
  {32'h38dbd427, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'h3cf8575c, 32'h00000000} /* (9, 14, 15) {real, imag} */,
  {32'h3f228072, 32'h00000000} /* (9, 14, 14) {real, imag} */,
  {32'h3f5a0dc1, 32'h00000000} /* (9, 14, 13) {real, imag} */,
  {32'h3f5d8e4d, 32'h00000000} /* (9, 14, 12) {real, imag} */,
  {32'h3e014a0e, 32'h00000000} /* (9, 14, 11) {real, imag} */,
  {32'hbdcc865a, 32'h00000000} /* (9, 14, 10) {real, imag} */,
  {32'h3ddf2aea, 32'h00000000} /* (9, 14, 9) {real, imag} */,
  {32'hbea568ed, 32'h00000000} /* (9, 14, 8) {real, imag} */,
  {32'hbda23242, 32'h00000000} /* (9, 14, 7) {real, imag} */,
  {32'h3eedfaf2, 32'h00000000} /* (9, 14, 6) {real, imag} */,
  {32'h3f811565, 32'h00000000} /* (9, 14, 5) {real, imag} */,
  {32'hbe69afaf, 32'h00000000} /* (9, 14, 4) {real, imag} */,
  {32'hbf3c4ee7, 32'h00000000} /* (9, 14, 3) {real, imag} */,
  {32'hbee14713, 32'h00000000} /* (9, 14, 2) {real, imag} */,
  {32'hbddc13d5, 32'h00000000} /* (9, 14, 1) {real, imag} */,
  {32'hbd535437, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hbeda3974, 32'h00000000} /* (9, 13, 15) {real, imag} */,
  {32'h3e1e67b1, 32'h00000000} /* (9, 13, 14) {real, imag} */,
  {32'h3ebf3794, 32'h00000000} /* (9, 13, 13) {real, imag} */,
  {32'h3e80ed05, 32'h00000000} /* (9, 13, 12) {real, imag} */,
  {32'hbe1114b7, 32'h00000000} /* (9, 13, 11) {real, imag} */,
  {32'hbe30eaeb, 32'h00000000} /* (9, 13, 10) {real, imag} */,
  {32'h3e83b9ea, 32'h00000000} /* (9, 13, 9) {real, imag} */,
  {32'h3d5064e6, 32'h00000000} /* (9, 13, 8) {real, imag} */,
  {32'hbd2af3af, 32'h00000000} /* (9, 13, 7) {real, imag} */,
  {32'h3eab3678, 32'h00000000} /* (9, 13, 6) {real, imag} */,
  {32'h3f17834f, 32'h00000000} /* (9, 13, 5) {real, imag} */,
  {32'hbdcb1eeb, 32'h00000000} /* (9, 13, 4) {real, imag} */,
  {32'hbf449e31, 32'h00000000} /* (9, 13, 3) {real, imag} */,
  {32'hbebd39d6, 32'h00000000} /* (9, 13, 2) {real, imag} */,
  {32'h3e2bccb5, 32'h00000000} /* (9, 13, 1) {real, imag} */,
  {32'h3dc35015, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hbde4a1ea, 32'h00000000} /* (9, 12, 15) {real, imag} */,
  {32'hbe11b59a, 32'h00000000} /* (9, 12, 14) {real, imag} */,
  {32'hbec3b6b7, 32'h00000000} /* (9, 12, 13) {real, imag} */,
  {32'hbe59bd79, 32'h00000000} /* (9, 12, 12) {real, imag} */,
  {32'h3db2d4e0, 32'h00000000} /* (9, 12, 11) {real, imag} */,
  {32'h3e732302, 32'h00000000} /* (9, 12, 10) {real, imag} */,
  {32'h3f1bd818, 32'h00000000} /* (9, 12, 9) {real, imag} */,
  {32'h3ec641c2, 32'h00000000} /* (9, 12, 8) {real, imag} */,
  {32'h3dca9ef3, 32'h00000000} /* (9, 12, 7) {real, imag} */,
  {32'hbcd2baba, 32'h00000000} /* (9, 12, 6) {real, imag} */,
  {32'h3df653e5, 32'h00000000} /* (9, 12, 5) {real, imag} */,
  {32'h3e854507, 32'h00000000} /* (9, 12, 4) {real, imag} */,
  {32'hbeac4167, 32'h00000000} /* (9, 12, 3) {real, imag} */,
  {32'hbedba76a, 32'h00000000} /* (9, 12, 2) {real, imag} */,
  {32'h3e33fdb9, 32'h00000000} /* (9, 12, 1) {real, imag} */,
  {32'h3e177cf9, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'h3e59c0c7, 32'h00000000} /* (9, 11, 15) {real, imag} */,
  {32'h3e9955a6, 32'h00000000} /* (9, 11, 14) {real, imag} */,
  {32'hbe05f26e, 32'h00000000} /* (9, 11, 13) {real, imag} */,
  {32'hbf2899f8, 32'h00000000} /* (9, 11, 12) {real, imag} */,
  {32'hbe9f504e, 32'h00000000} /* (9, 11, 11) {real, imag} */,
  {32'h3e9dab9a, 32'h00000000} /* (9, 11, 10) {real, imag} */,
  {32'h3f418a80, 32'h00000000} /* (9, 11, 9) {real, imag} */,
  {32'hbda2433c, 32'h00000000} /* (9, 11, 8) {real, imag} */,
  {32'hbe657716, 32'h00000000} /* (9, 11, 7) {real, imag} */,
  {32'h3e17ad85, 32'h00000000} /* (9, 11, 6) {real, imag} */,
  {32'h3edbaf77, 32'h00000000} /* (9, 11, 5) {real, imag} */,
  {32'h3f21ebf1, 32'h00000000} /* (9, 11, 4) {real, imag} */,
  {32'h3e14c306, 32'h00000000} /* (9, 11, 3) {real, imag} */,
  {32'h3e4ef044, 32'h00000000} /* (9, 11, 2) {real, imag} */,
  {32'h3ee63ae4, 32'h00000000} /* (9, 11, 1) {real, imag} */,
  {32'h3d96f7d0, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h3d0feb17, 32'h00000000} /* (9, 10, 15) {real, imag} */,
  {32'h3eb65dc6, 32'h00000000} /* (9, 10, 14) {real, imag} */,
  {32'hbe155929, 32'h00000000} /* (9, 10, 13) {real, imag} */,
  {32'hbf097e60, 32'h00000000} /* (9, 10, 12) {real, imag} */,
  {32'hbed5322d, 32'h00000000} /* (9, 10, 11) {real, imag} */,
  {32'hbefaba87, 32'h00000000} /* (9, 10, 10) {real, imag} */,
  {32'h3f23bf12, 32'h00000000} /* (9, 10, 9) {real, imag} */,
  {32'h3ebcca83, 32'h00000000} /* (9, 10, 8) {real, imag} */,
  {32'h3e12e5e2, 32'h00000000} /* (9, 10, 7) {real, imag} */,
  {32'h3d56e3b2, 32'h00000000} /* (9, 10, 6) {real, imag} */,
  {32'hbe89cd39, 32'h00000000} /* (9, 10, 5) {real, imag} */,
  {32'h3e83a1a0, 32'h00000000} /* (9, 10, 4) {real, imag} */,
  {32'h3e8663a7, 32'h00000000} /* (9, 10, 3) {real, imag} */,
  {32'h3f0e30eb, 32'h00000000} /* (9, 10, 2) {real, imag} */,
  {32'h3f0143d9, 32'h00000000} /* (9, 10, 1) {real, imag} */,
  {32'hbcc1d02a, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'hbdb07952, 32'h00000000} /* (9, 9, 15) {real, imag} */,
  {32'h3e61c20d, 32'h00000000} /* (9, 9, 14) {real, imag} */,
  {32'hbe8de32a, 32'h00000000} /* (9, 9, 13) {real, imag} */,
  {32'hbf37e9a6, 32'h00000000} /* (9, 9, 12) {real, imag} */,
  {32'hbe0d7244, 32'h00000000} /* (9, 9, 11) {real, imag} */,
  {32'hbf2b1a28, 32'h00000000} /* (9, 9, 10) {real, imag} */,
  {32'hbda1efa3, 32'h00000000} /* (9, 9, 9) {real, imag} */,
  {32'h3ea2cf19, 32'h00000000} /* (9, 9, 8) {real, imag} */,
  {32'h3ecfbfb5, 32'h00000000} /* (9, 9, 7) {real, imag} */,
  {32'h3d351220, 32'h00000000} /* (9, 9, 6) {real, imag} */,
  {32'hbdc802af, 32'h00000000} /* (9, 9, 5) {real, imag} */,
  {32'h3e257be9, 32'h00000000} /* (9, 9, 4) {real, imag} */,
  {32'h3ec64ba5, 32'h00000000} /* (9, 9, 3) {real, imag} */,
  {32'h3ebfe940, 32'h00000000} /* (9, 9, 2) {real, imag} */,
  {32'h3f22513f, 32'h00000000} /* (9, 9, 1) {real, imag} */,
  {32'h3eb676cb, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h3ce2c2c4, 32'h00000000} /* (9, 8, 15) {real, imag} */,
  {32'h3e94f583, 32'h00000000} /* (9, 8, 14) {real, imag} */,
  {32'h3e02c24f, 32'h00000000} /* (9, 8, 13) {real, imag} */,
  {32'hbd307ef2, 32'h00000000} /* (9, 8, 12) {real, imag} */,
  {32'hbdbb1e02, 32'h00000000} /* (9, 8, 11) {real, imag} */,
  {32'hbf0a9327, 32'h00000000} /* (9, 8, 10) {real, imag} */,
  {32'hbed062de, 32'h00000000} /* (9, 8, 9) {real, imag} */,
  {32'hbdddc83c, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'h3ecb0857, 32'h00000000} /* (9, 8, 7) {real, imag} */,
  {32'h3e3bc6fe, 32'h00000000} /* (9, 8, 6) {real, imag} */,
  {32'h3da9f8a3, 32'h00000000} /* (9, 8, 5) {real, imag} */,
  {32'hbee09878, 32'h00000000} /* (9, 8, 4) {real, imag} */,
  {32'hbe5fecb1, 32'h00000000} /* (9, 8, 3) {real, imag} */,
  {32'h3aca097a, 32'h00000000} /* (9, 8, 2) {real, imag} */,
  {32'h3e92d1ad, 32'h00000000} /* (9, 8, 1) {real, imag} */,
  {32'h3de8c062, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h3e418936, 32'h00000000} /* (9, 7, 15) {real, imag} */,
  {32'h3efe73fa, 32'h00000000} /* (9, 7, 14) {real, imag} */,
  {32'h3f1e3124, 32'h00000000} /* (9, 7, 13) {real, imag} */,
  {32'h3f46bb1e, 32'h00000000} /* (9, 7, 12) {real, imag} */,
  {32'hbe6c78aa, 32'h00000000} /* (9, 7, 11) {real, imag} */,
  {32'hbf488ca9, 32'h00000000} /* (9, 7, 10) {real, imag} */,
  {32'hbe67ac94, 32'h00000000} /* (9, 7, 9) {real, imag} */,
  {32'hbe2677ab, 32'h00000000} /* (9, 7, 8) {real, imag} */,
  {32'h3e0989dc, 32'h00000000} /* (9, 7, 7) {real, imag} */,
  {32'h3e5d1bea, 32'h00000000} /* (9, 7, 6) {real, imag} */,
  {32'h3d7f87a0, 32'h00000000} /* (9, 7, 5) {real, imag} */,
  {32'hbe5a3f2e, 32'h00000000} /* (9, 7, 4) {real, imag} */,
  {32'hbd2626e4, 32'h00000000} /* (9, 7, 3) {real, imag} */,
  {32'hbcd42846, 32'h00000000} /* (9, 7, 2) {real, imag} */,
  {32'hbe5ba1be, 32'h00000000} /* (9, 7, 1) {real, imag} */,
  {32'hbdb86c5c, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h3eb75057, 32'h00000000} /* (9, 6, 15) {real, imag} */,
  {32'h3eaebfcf, 32'h00000000} /* (9, 6, 14) {real, imag} */,
  {32'h3edb6b9f, 32'h00000000} /* (9, 6, 13) {real, imag} */,
  {32'h3f169751, 32'h00000000} /* (9, 6, 12) {real, imag} */,
  {32'hbe04686b, 32'h00000000} /* (9, 6, 11) {real, imag} */,
  {32'hbef4c0e0, 32'h00000000} /* (9, 6, 10) {real, imag} */,
  {32'h3e13f380, 32'h00000000} /* (9, 6, 9) {real, imag} */,
  {32'hbf216cdb, 32'h00000000} /* (9, 6, 8) {real, imag} */,
  {32'hbef424d7, 32'h00000000} /* (9, 6, 7) {real, imag} */,
  {32'h3ee06557, 32'h00000000} /* (9, 6, 6) {real, imag} */,
  {32'h3ef6e570, 32'h00000000} /* (9, 6, 5) {real, imag} */,
  {32'h3ddce34a, 32'h00000000} /* (9, 6, 4) {real, imag} */,
  {32'hbeefec1d, 32'h00000000} /* (9, 6, 3) {real, imag} */,
  {32'hbef9d59e, 32'h00000000} /* (9, 6, 2) {real, imag} */,
  {32'h3d1328fb, 32'h00000000} /* (9, 6, 1) {real, imag} */,
  {32'h3dc41ea2, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h3eaa0da9, 32'h00000000} /* (9, 5, 15) {real, imag} */,
  {32'h3ead07c6, 32'h00000000} /* (9, 5, 14) {real, imag} */,
  {32'h3dd6243e, 32'h00000000} /* (9, 5, 13) {real, imag} */,
  {32'h3eb6e88f, 32'h00000000} /* (9, 5, 12) {real, imag} */,
  {32'h3d439eda, 32'h00000000} /* (9, 5, 11) {real, imag} */,
  {32'hbe2db3fe, 32'h00000000} /* (9, 5, 10) {real, imag} */,
  {32'h3d16a5da, 32'h00000000} /* (9, 5, 9) {real, imag} */,
  {32'hbf0f1aa7, 32'h00000000} /* (9, 5, 8) {real, imag} */,
  {32'hbe3f56dd, 32'h00000000} /* (9, 5, 7) {real, imag} */,
  {32'h3f62951e, 32'h00000000} /* (9, 5, 6) {real, imag} */,
  {32'h3f61217c, 32'h00000000} /* (9, 5, 5) {real, imag} */,
  {32'h3e866a82, 32'h00000000} /* (9, 5, 4) {real, imag} */,
  {32'hbe950416, 32'h00000000} /* (9, 5, 3) {real, imag} */,
  {32'hbe9d61bc, 32'h00000000} /* (9, 5, 2) {real, imag} */,
  {32'hbeb81b95, 32'h00000000} /* (9, 5, 1) {real, imag} */,
  {32'h3c108cfa, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'hbd574e6a, 32'h00000000} /* (9, 4, 15) {real, imag} */,
  {32'h3e692c97, 32'h00000000} /* (9, 4, 14) {real, imag} */,
  {32'h3ead880d, 32'h00000000} /* (9, 4, 13) {real, imag} */,
  {32'h3e682f7c, 32'h00000000} /* (9, 4, 12) {real, imag} */,
  {32'hbddf992a, 32'h00000000} /* (9, 4, 11) {real, imag} */,
  {32'hbf62911f, 32'h00000000} /* (9, 4, 10) {real, imag} */,
  {32'hbf15f214, 32'h00000000} /* (9, 4, 9) {real, imag} */,
  {32'hbf263d33, 32'h00000000} /* (9, 4, 8) {real, imag} */,
  {32'hbe9b5984, 32'h00000000} /* (9, 4, 7) {real, imag} */,
  {32'h3efd55d0, 32'h00000000} /* (9, 4, 6) {real, imag} */,
  {32'h3e73ffb7, 32'h00000000} /* (9, 4, 5) {real, imag} */,
  {32'h3ebac0a5, 32'h00000000} /* (9, 4, 4) {real, imag} */,
  {32'h3e7e5873, 32'h00000000} /* (9, 4, 3) {real, imag} */,
  {32'hbdde7cf7, 32'h00000000} /* (9, 4, 2) {real, imag} */,
  {32'hbebd0ada, 32'h00000000} /* (9, 4, 1) {real, imag} */,
  {32'hbc34992e, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'hbe5a329d, 32'h00000000} /* (9, 3, 15) {real, imag} */,
  {32'hbe4407c1, 32'h00000000} /* (9, 3, 14) {real, imag} */,
  {32'hbf088839, 32'h00000000} /* (9, 3, 13) {real, imag} */,
  {32'hbe883f90, 32'h00000000} /* (9, 3, 12) {real, imag} */,
  {32'hbe1a03f8, 32'h00000000} /* (9, 3, 11) {real, imag} */,
  {32'hbf3e1f2e, 32'h00000000} /* (9, 3, 10) {real, imag} */,
  {32'hbc860a6c, 32'h00000000} /* (9, 3, 9) {real, imag} */,
  {32'hbd184b59, 32'h00000000} /* (9, 3, 8) {real, imag} */,
  {32'hbe297f6b, 32'h00000000} /* (9, 3, 7) {real, imag} */,
  {32'hbe3a10f8, 32'h00000000} /* (9, 3, 6) {real, imag} */,
  {32'hbe79076f, 32'h00000000} /* (9, 3, 5) {real, imag} */,
  {32'hbe59cede, 32'h00000000} /* (9, 3, 4) {real, imag} */,
  {32'hbe75dc22, 32'h00000000} /* (9, 3, 3) {real, imag} */,
  {32'h3c04fd9c, 32'h00000000} /* (9, 3, 2) {real, imag} */,
  {32'h3eef6f34, 32'h00000000} /* (9, 3, 1) {real, imag} */,
  {32'h3e3e2fb8, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'hbd327e04, 32'h00000000} /* (9, 2, 15) {real, imag} */,
  {32'hbe57cd45, 32'h00000000} /* (9, 2, 14) {real, imag} */,
  {32'hbf524d94, 32'h00000000} /* (9, 2, 13) {real, imag} */,
  {32'hbf1419bf, 32'h00000000} /* (9, 2, 12) {real, imag} */,
  {32'hbc5742f7, 32'h00000000} /* (9, 2, 11) {real, imag} */,
  {32'hbb9c574c, 32'h00000000} /* (9, 2, 10) {real, imag} */,
  {32'hbec60feb, 32'h00000000} /* (9, 2, 9) {real, imag} */,
  {32'h3d0dba1a, 32'h00000000} /* (9, 2, 8) {real, imag} */,
  {32'h3db83779, 32'h00000000} /* (9, 2, 7) {real, imag} */,
  {32'hbd21928d, 32'h00000000} /* (9, 2, 6) {real, imag} */,
  {32'hbe5ab2b0, 32'h00000000} /* (9, 2, 5) {real, imag} */,
  {32'h3dcb0565, 32'h00000000} /* (9, 2, 4) {real, imag} */,
  {32'hbdd30ed3, 32'h00000000} /* (9, 2, 3) {real, imag} */,
  {32'hbce497d0, 32'h00000000} /* (9, 2, 2) {real, imag} */,
  {32'h3f15085f, 32'h00000000} /* (9, 2, 1) {real, imag} */,
  {32'h3e87e640, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'hbd99fd0e, 32'h00000000} /* (9, 1, 15) {real, imag} */,
  {32'hbda33bfb, 32'h00000000} /* (9, 1, 14) {real, imag} */,
  {32'hbe4888a6, 32'h00000000} /* (9, 1, 13) {real, imag} */,
  {32'h3d632666, 32'h00000000} /* (9, 1, 12) {real, imag} */,
  {32'h3ee0e5f3, 32'h00000000} /* (9, 1, 11) {real, imag} */,
  {32'h3da8767f, 32'h00000000} /* (9, 1, 10) {real, imag} */,
  {32'hbb4ea475, 32'h00000000} /* (9, 1, 9) {real, imag} */,
  {32'h3ea02055, 32'h00000000} /* (9, 1, 8) {real, imag} */,
  {32'h3e9cb71e, 32'h00000000} /* (9, 1, 7) {real, imag} */,
  {32'h3cafd64c, 32'h00000000} /* (9, 1, 6) {real, imag} */,
  {32'hbebf7e0a, 32'h00000000} /* (9, 1, 5) {real, imag} */,
  {32'h3f39fe11, 32'h00000000} /* (9, 1, 4) {real, imag} */,
  {32'h3ea77d21, 32'h00000000} /* (9, 1, 3) {real, imag} */,
  {32'hbefd1068, 32'h00000000} /* (9, 1, 2) {real, imag} */,
  {32'h3daf9302, 32'h00000000} /* (9, 1, 1) {real, imag} */,
  {32'h3e133951, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h3e0089a2, 32'h00000000} /* (9, 0, 15) {real, imag} */,
  {32'hbd8ea50a, 32'h00000000} /* (9, 0, 14) {real, imag} */,
  {32'hbd6e9ba3, 32'h00000000} /* (9, 0, 13) {real, imag} */,
  {32'h3e40cd95, 32'h00000000} /* (9, 0, 12) {real, imag} */,
  {32'h3e68f382, 32'h00000000} /* (9, 0, 11) {real, imag} */,
  {32'h3dd2d97f, 32'h00000000} /* (9, 0, 10) {real, imag} */,
  {32'hbdd7d35d, 32'h00000000} /* (9, 0, 9) {real, imag} */,
  {32'hbd15d6cb, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'h3e3d7925, 32'h00000000} /* (9, 0, 7) {real, imag} */,
  {32'hbd51dbcf, 32'h00000000} /* (9, 0, 6) {real, imag} */,
  {32'hbe8d4684, 32'h00000000} /* (9, 0, 5) {real, imag} */,
  {32'h3de29332, 32'h00000000} /* (9, 0, 4) {real, imag} */,
  {32'h3d6d3b97, 32'h00000000} /* (9, 0, 3) {real, imag} */,
  {32'hbdc8ee1c, 32'h00000000} /* (9, 0, 2) {real, imag} */,
  {32'hbdae9635, 32'h00000000} /* (9, 0, 1) {real, imag} */,
  {32'hbd1c86bf, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h3dfc2765, 32'h00000000} /* (8, 15, 15) {real, imag} */,
  {32'h3d9c011e, 32'h00000000} /* (8, 15, 14) {real, imag} */,
  {32'h3d7ee2c6, 32'h00000000} /* (8, 15, 13) {real, imag} */,
  {32'h3df23bfe, 32'h00000000} /* (8, 15, 12) {real, imag} */,
  {32'h3ed355f6, 32'h00000000} /* (8, 15, 11) {real, imag} */,
  {32'h3e4188a2, 32'h00000000} /* (8, 15, 10) {real, imag} */,
  {32'h3ccc0520, 32'h00000000} /* (8, 15, 9) {real, imag} */,
  {32'hbec34382, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hbec2bf9e, 32'h00000000} /* (8, 15, 7) {real, imag} */,
  {32'hbdd72b6a, 32'h00000000} /* (8, 15, 6) {real, imag} */,
  {32'hbd8288ab, 32'h00000000} /* (8, 15, 5) {real, imag} */,
  {32'hbeb10e26, 32'h00000000} /* (8, 15, 4) {real, imag} */,
  {32'hbe8325cb, 32'h00000000} /* (8, 15, 3) {real, imag} */,
  {32'hbdf006fe, 32'h00000000} /* (8, 15, 2) {real, imag} */,
  {32'h3d801c65, 32'h00000000} /* (8, 15, 1) {real, imag} */,
  {32'h3d1b60b4, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'h3e817ee6, 32'h00000000} /* (8, 14, 15) {real, imag} */,
  {32'h3e8449c4, 32'h00000000} /* (8, 14, 14) {real, imag} */,
  {32'hbd0c2cfe, 32'h00000000} /* (8, 14, 13) {real, imag} */,
  {32'h3e6ed69d, 32'h00000000} /* (8, 14, 12) {real, imag} */,
  {32'h3eab892b, 32'h00000000} /* (8, 14, 11) {real, imag} */,
  {32'hbe987fc5, 32'h00000000} /* (8, 14, 10) {real, imag} */,
  {32'hbe10faf3, 32'h00000000} /* (8, 14, 9) {real, imag} */,
  {32'hbe90d907, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'hbefe92d2, 32'h00000000} /* (8, 14, 7) {real, imag} */,
  {32'h3dc231bd, 32'h00000000} /* (8, 14, 6) {real, imag} */,
  {32'h3e744f42, 32'h00000000} /* (8, 14, 5) {real, imag} */,
  {32'hbf20cd5d, 32'h00000000} /* (8, 14, 4) {real, imag} */,
  {32'hbe9a6236, 32'h00000000} /* (8, 14, 3) {real, imag} */,
  {32'hbdf75a54, 32'h00000000} /* (8, 14, 2) {real, imag} */,
  {32'hbe7d3279, 32'h00000000} /* (8, 14, 1) {real, imag} */,
  {32'hbc741f09, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hbe3a9545, 32'h00000000} /* (8, 13, 15) {real, imag} */,
  {32'hbed128bf, 32'h00000000} /* (8, 13, 14) {real, imag} */,
  {32'hbe5101c6, 32'h00000000} /* (8, 13, 13) {real, imag} */,
  {32'h3eb03c69, 32'h00000000} /* (8, 13, 12) {real, imag} */,
  {32'hbc08831c, 32'h00000000} /* (8, 13, 11) {real, imag} */,
  {32'hbe2d44ca, 32'h00000000} /* (8, 13, 10) {real, imag} */,
  {32'h3f051d87, 32'h00000000} /* (8, 13, 9) {real, imag} */,
  {32'h3cdfd0fa, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'hbedff107, 32'h00000000} /* (8, 13, 7) {real, imag} */,
  {32'h3ec74d83, 32'h00000000} /* (8, 13, 6) {real, imag} */,
  {32'h3efeda93, 32'h00000000} /* (8, 13, 5) {real, imag} */,
  {32'hbc2a534a, 32'h00000000} /* (8, 13, 4) {real, imag} */,
  {32'hbf09c0f7, 32'h00000000} /* (8, 13, 3) {real, imag} */,
  {32'hbdec7aaf, 32'h00000000} /* (8, 13, 2) {real, imag} */,
  {32'hbd0a9c38, 32'h00000000} /* (8, 13, 1) {real, imag} */,
  {32'h3df3239d, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'hbda77e98, 32'h00000000} /* (8, 12, 15) {real, imag} */,
  {32'hbdacc94b, 32'h00000000} /* (8, 12, 14) {real, imag} */,
  {32'h3d7decaa, 32'h00000000} /* (8, 12, 13) {real, imag} */,
  {32'hbd61c21c, 32'h00000000} /* (8, 12, 12) {real, imag} */,
  {32'hbe48a856, 32'h00000000} /* (8, 12, 11) {real, imag} */,
  {32'h3e4f9d20, 32'h00000000} /* (8, 12, 10) {real, imag} */,
  {32'h3f12c6aa, 32'h00000000} /* (8, 12, 9) {real, imag} */,
  {32'hbdb1a9bc, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'hbe8e5339, 32'h00000000} /* (8, 12, 7) {real, imag} */,
  {32'hbecfc05e, 32'h00000000} /* (8, 12, 6) {real, imag} */,
  {32'hbf007ad3, 32'h00000000} /* (8, 12, 5) {real, imag} */,
  {32'hbdc674bf, 32'h00000000} /* (8, 12, 4) {real, imag} */,
  {32'hbb62eea8, 32'h00000000} /* (8, 12, 3) {real, imag} */,
  {32'h3c5b13ef, 32'h00000000} /* (8, 12, 2) {real, imag} */,
  {32'hbca31da4, 32'h00000000} /* (8, 12, 1) {real, imag} */,
  {32'h3d0c8e08, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'h3e3e05b8, 32'h00000000} /* (8, 11, 15) {real, imag} */,
  {32'h3e541aea, 32'h00000000} /* (8, 11, 14) {real, imag} */,
  {32'hbb1fcae0, 32'h00000000} /* (8, 11, 13) {real, imag} */,
  {32'hbf53525a, 32'h00000000} /* (8, 11, 12) {real, imag} */,
  {32'hbf072baa, 32'h00000000} /* (8, 11, 11) {real, imag} */,
  {32'h3e4415c1, 32'h00000000} /* (8, 11, 10) {real, imag} */,
  {32'h3f0efacd, 32'h00000000} /* (8, 11, 9) {real, imag} */,
  {32'hbdf3edcf, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'hbe7ca4c3, 32'h00000000} /* (8, 11, 7) {real, imag} */,
  {32'hbef227ae, 32'h00000000} /* (8, 11, 6) {real, imag} */,
  {32'hbefd8e99, 32'h00000000} /* (8, 11, 5) {real, imag} */,
  {32'hbd6f329d, 32'h00000000} /* (8, 11, 4) {real, imag} */,
  {32'h3e2a2626, 32'h00000000} /* (8, 11, 3) {real, imag} */,
  {32'hbd30402e, 32'h00000000} /* (8, 11, 2) {real, imag} */,
  {32'hbd21c682, 32'h00000000} /* (8, 11, 1) {real, imag} */,
  {32'hbdb8ccc0, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'hbdec14c0, 32'h00000000} /* (8, 10, 15) {real, imag} */,
  {32'hbe1cc6fa, 32'h00000000} /* (8, 10, 14) {real, imag} */,
  {32'h3dd9e749, 32'h00000000} /* (8, 10, 13) {real, imag} */,
  {32'hbef9f2c5, 32'h00000000} /* (8, 10, 12) {real, imag} */,
  {32'hbeab93a2, 32'h00000000} /* (8, 10, 11) {real, imag} */,
  {32'hbd6e69e2, 32'h00000000} /* (8, 10, 10) {real, imag} */,
  {32'h3f082606, 32'h00000000} /* (8, 10, 9) {real, imag} */,
  {32'h3eaa2b1c, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'hbe3b6b2c, 32'h00000000} /* (8, 10, 7) {real, imag} */,
  {32'h3e3b7db0, 32'h00000000} /* (8, 10, 6) {real, imag} */,
  {32'hbd1a91ee, 32'h00000000} /* (8, 10, 5) {real, imag} */,
  {32'h3d467602, 32'h00000000} /* (8, 10, 4) {real, imag} */,
  {32'h3e8f51a0, 32'h00000000} /* (8, 10, 3) {real, imag} */,
  {32'h3eca848b, 32'h00000000} /* (8, 10, 2) {real, imag} */,
  {32'h3e9077d9, 32'h00000000} /* (8, 10, 1) {real, imag} */,
  {32'hbdf25283, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'hbe8beb36, 32'h00000000} /* (8, 9, 15) {real, imag} */,
  {32'hbe1f2ebd, 32'h00000000} /* (8, 9, 14) {real, imag} */,
  {32'h3dab79ef, 32'h00000000} /* (8, 9, 13) {real, imag} */,
  {32'hbde4d4a6, 32'h00000000} /* (8, 9, 12) {real, imag} */,
  {32'h3de1ad22, 32'h00000000} /* (8, 9, 11) {real, imag} */,
  {32'hbe20da10, 32'h00000000} /* (8, 9, 10) {real, imag} */,
  {32'hbe64aa7e, 32'h00000000} /* (8, 9, 9) {real, imag} */,
  {32'hbda6ebd8, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'hbe15fb5e, 32'h00000000} /* (8, 9, 7) {real, imag} */,
  {32'h3e8f65d7, 32'h00000000} /* (8, 9, 6) {real, imag} */,
  {32'h3eac5fd0, 32'h00000000} /* (8, 9, 5) {real, imag} */,
  {32'h3e64688e, 32'h00000000} /* (8, 9, 4) {real, imag} */,
  {32'hbbf13ff0, 32'h00000000} /* (8, 9, 3) {real, imag} */,
  {32'hbd82cc00, 32'h00000000} /* (8, 9, 2) {real, imag} */,
  {32'h3eca05ad, 32'h00000000} /* (8, 9, 1) {real, imag} */,
  {32'hbd77097f, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'hbe2af45c, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'h3c44d514, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'h3eff78a3, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'h3effeaef, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'h3de0f7cd, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'hbec2491c, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'hbf4c9931, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'hbe775cf7, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'h3dc8b82e, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'h3e0b70e4, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'h3db5a73f, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'hbf130921, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'hbf30cb75, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'hbed30b12, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'h3e95a4f4, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h3dfa443b, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h3db96cb4, 32'h00000000} /* (8, 7, 15) {real, imag} */,
  {32'h3e30470c, 32'h00000000} /* (8, 7, 14) {real, imag} */,
  {32'h3ecb529e, 32'h00000000} /* (8, 7, 13) {real, imag} */,
  {32'h3f80a1ff, 32'h00000000} /* (8, 7, 12) {real, imag} */,
  {32'h3edad61e, 32'h00000000} /* (8, 7, 11) {real, imag} */,
  {32'hbccfd054, 32'h00000000} /* (8, 7, 10) {real, imag} */,
  {32'hbe1e1534, 32'h00000000} /* (8, 7, 9) {real, imag} */,
  {32'h3d5a4f97, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h3e513936, 32'h00000000} /* (8, 7, 7) {real, imag} */,
  {32'h3e8fdc67, 32'h00000000} /* (8, 7, 6) {real, imag} */,
  {32'hbe3752d6, 32'h00000000} /* (8, 7, 5) {real, imag} */,
  {32'hbf006690, 32'h00000000} /* (8, 7, 4) {real, imag} */,
  {32'hbf007007, 32'h00000000} /* (8, 7, 3) {real, imag} */,
  {32'hbed3ecc2, 32'h00000000} /* (8, 7, 2) {real, imag} */,
  {32'hbeab62e7, 32'h00000000} /* (8, 7, 1) {real, imag} */,
  {32'hbd50412c, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h3d53221e, 32'h00000000} /* (8, 6, 15) {real, imag} */,
  {32'h3de2030e, 32'h00000000} /* (8, 6, 14) {real, imag} */,
  {32'hbd067b7c, 32'h00000000} /* (8, 6, 13) {real, imag} */,
  {32'h3e9492e4, 32'h00000000} /* (8, 6, 12) {real, imag} */,
  {32'h3ea61a98, 32'h00000000} /* (8, 6, 11) {real, imag} */,
  {32'hbed1eb59, 32'h00000000} /* (8, 6, 10) {real, imag} */,
  {32'hbe165f9b, 32'h00000000} /* (8, 6, 9) {real, imag} */,
  {32'hbe252206, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'hbefa2565, 32'h00000000} /* (8, 6, 7) {real, imag} */,
  {32'h3e942487, 32'h00000000} /* (8, 6, 6) {real, imag} */,
  {32'h3f053913, 32'h00000000} /* (8, 6, 5) {real, imag} */,
  {32'h3e180304, 32'h00000000} /* (8, 6, 4) {real, imag} */,
  {32'hbf090848, 32'h00000000} /* (8, 6, 3) {real, imag} */,
  {32'hbea7411e, 32'h00000000} /* (8, 6, 2) {real, imag} */,
  {32'h3e0635bc, 32'h00000000} /* (8, 6, 1) {real, imag} */,
  {32'hbd9c7051, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'h3d4715c3, 32'h00000000} /* (8, 5, 15) {real, imag} */,
  {32'h3ed70482, 32'h00000000} /* (8, 5, 14) {real, imag} */,
  {32'h3e75ba31, 32'h00000000} /* (8, 5, 13) {real, imag} */,
  {32'h3e8484ea, 32'h00000000} /* (8, 5, 12) {real, imag} */,
  {32'h3cdb3d94, 32'h00000000} /* (8, 5, 11) {real, imag} */,
  {32'hbe9b8758, 32'h00000000} /* (8, 5, 10) {real, imag} */,
  {32'hbd9c900f, 32'h00000000} /* (8, 5, 9) {real, imag} */,
  {32'hbef1f775, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'hbe368e75, 32'h00000000} /* (8, 5, 7) {real, imag} */,
  {32'h3f06aad9, 32'h00000000} /* (8, 5, 6) {real, imag} */,
  {32'h3f21d2f4, 32'h00000000} /* (8, 5, 5) {real, imag} */,
  {32'h3f0aff0a, 32'h00000000} /* (8, 5, 4) {real, imag} */,
  {32'hbcca585e, 32'h00000000} /* (8, 5, 3) {real, imag} */,
  {32'hbe166d4e, 32'h00000000} /* (8, 5, 2) {real, imag} */,
  {32'hbd156840, 32'h00000000} /* (8, 5, 1) {real, imag} */,
  {32'hbbc7eafd, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'hbe3ff53d, 32'h00000000} /* (8, 4, 15) {real, imag} */,
  {32'h3f315f58, 32'h00000000} /* (8, 4, 14) {real, imag} */,
  {32'h3f24478a, 32'h00000000} /* (8, 4, 13) {real, imag} */,
  {32'h3e76a54e, 32'h00000000} /* (8, 4, 12) {real, imag} */,
  {32'hbe344106, 32'h00000000} /* (8, 4, 11) {real, imag} */,
  {32'hbed18530, 32'h00000000} /* (8, 4, 10) {real, imag} */,
  {32'h3e12717f, 32'h00000000} /* (8, 4, 9) {real, imag} */,
  {32'hbe2c176f, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'h3e7f1e3f, 32'h00000000} /* (8, 4, 7) {real, imag} */,
  {32'h3efb88ca, 32'h00000000} /* (8, 4, 6) {real, imag} */,
  {32'h3e1780f9, 32'h00000000} /* (8, 4, 5) {real, imag} */,
  {32'h3f0b95ba, 32'h00000000} /* (8, 4, 4) {real, imag} */,
  {32'h3ed0c727, 32'h00000000} /* (8, 4, 3) {real, imag} */,
  {32'hbe871ec9, 32'h00000000} /* (8, 4, 2) {real, imag} */,
  {32'hbe7a5058, 32'h00000000} /* (8, 4, 1) {real, imag} */,
  {32'hbd147b09, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'hbd7dcef8, 32'h00000000} /* (8, 3, 15) {real, imag} */,
  {32'h3daaf962, 32'h00000000} /* (8, 3, 14) {real, imag} */,
  {32'hbeb67808, 32'h00000000} /* (8, 3, 13) {real, imag} */,
  {32'h3e20c1b8, 32'h00000000} /* (8, 3, 12) {real, imag} */,
  {32'h3db82823, 32'h00000000} /* (8, 3, 11) {real, imag} */,
  {32'hbef04bb5, 32'h00000000} /* (8, 3, 10) {real, imag} */,
  {32'hbdc101d5, 32'h00000000} /* (8, 3, 9) {real, imag} */,
  {32'h3d1b29d2, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'h3ebc2efe, 32'h00000000} /* (8, 3, 7) {real, imag} */,
  {32'h3f1856b4, 32'h00000000} /* (8, 3, 6) {real, imag} */,
  {32'h3e956f7c, 32'h00000000} /* (8, 3, 5) {real, imag} */,
  {32'hba8ffca6, 32'h00000000} /* (8, 3, 4) {real, imag} */,
  {32'h3c82ab9a, 32'h00000000} /* (8, 3, 3) {real, imag} */,
  {32'h3d9eceaf, 32'h00000000} /* (8, 3, 2) {real, imag} */,
  {32'h3c541ce3, 32'h00000000} /* (8, 3, 1) {real, imag} */,
  {32'hbc8190d8, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'h3d938744, 32'h00000000} /* (8, 2, 15) {real, imag} */,
  {32'hbeaf314b, 32'h00000000} /* (8, 2, 14) {real, imag} */,
  {32'hbf8260fe, 32'h00000000} /* (8, 2, 13) {real, imag} */,
  {32'hbeb5099a, 32'h00000000} /* (8, 2, 12) {real, imag} */,
  {32'hbe2ac1cd, 32'h00000000} /* (8, 2, 11) {real, imag} */,
  {32'hbe5124d7, 32'h00000000} /* (8, 2, 10) {real, imag} */,
  {32'hbdc44f2d, 32'h00000000} /* (8, 2, 9) {real, imag} */,
  {32'hbe95f56b, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'hbe28a8bf, 32'h00000000} /* (8, 2, 7) {real, imag} */,
  {32'h3f279d31, 32'h00000000} /* (8, 2, 6) {real, imag} */,
  {32'h3ee9276b, 32'h00000000} /* (8, 2, 5) {real, imag} */,
  {32'h3e8dd3cf, 32'h00000000} /* (8, 2, 4) {real, imag} */,
  {32'h3d7cb9e4, 32'h00000000} /* (8, 2, 3) {real, imag} */,
  {32'h3d041fa4, 32'h00000000} /* (8, 2, 2) {real, imag} */,
  {32'hbe45126b, 32'h00000000} /* (8, 2, 1) {real, imag} */,
  {32'hbe10b6e0, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'hbddf30dd, 32'h00000000} /* (8, 1, 15) {real, imag} */,
  {32'hbebfb29c, 32'h00000000} /* (8, 1, 14) {real, imag} */,
  {32'hbed48fe2, 32'h00000000} /* (8, 1, 13) {real, imag} */,
  {32'h3e778455, 32'h00000000} /* (8, 1, 12) {real, imag} */,
  {32'hbea6886a, 32'h00000000} /* (8, 1, 11) {real, imag} */,
  {32'hbe667600, 32'h00000000} /* (8, 1, 10) {real, imag} */,
  {32'h3f15e9e6, 32'h00000000} /* (8, 1, 9) {real, imag} */,
  {32'h3d91a861, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'h3e0db675, 32'h00000000} /* (8, 1, 7) {real, imag} */,
  {32'h3f05c399, 32'h00000000} /* (8, 1, 6) {real, imag} */,
  {32'h3e827944, 32'h00000000} /* (8, 1, 5) {real, imag} */,
  {32'h3e61f3e7, 32'h00000000} /* (8, 1, 4) {real, imag} */,
  {32'hbd601b37, 32'h00000000} /* (8, 1, 3) {real, imag} */,
  {32'hbe5cf2cf, 32'h00000000} /* (8, 1, 2) {real, imag} */,
  {32'hbec41300, 32'h00000000} /* (8, 1, 1) {real, imag} */,
  {32'hbe8509b3, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'hbe4e17c3, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'hbe19b963, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'h3e2481e8, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'h3e872bf1, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'hbddb29b5, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'hbd40914f, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'h3ed072b7, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'h3e9e39db, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'h3e81113e, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'h3e885c4a, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'h3e4a482e, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'h3bc6361b, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'hbda67cd9, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'hbc92d78a, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'hbe5f0bf0, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'hbe3c0837, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h3e37e089, 32'h00000000} /* (7, 15, 15) {real, imag} */,
  {32'h3e10ed87, 32'h00000000} /* (7, 15, 14) {real, imag} */,
  {32'hbe2198d4, 32'h00000000} /* (7, 15, 13) {real, imag} */,
  {32'hbe9eb237, 32'h00000000} /* (7, 15, 12) {real, imag} */,
  {32'h3de439c3, 32'h00000000} /* (7, 15, 11) {real, imag} */,
  {32'hbe167141, 32'h00000000} /* (7, 15, 10) {real, imag} */,
  {32'hbe414bc8, 32'h00000000} /* (7, 15, 9) {real, imag} */,
  {32'hbe13f284, 32'h00000000} /* (7, 15, 8) {real, imag} */,
  {32'h3e0d969a, 32'h00000000} /* (7, 15, 7) {real, imag} */,
  {32'h3ec4659e, 32'h00000000} /* (7, 15, 6) {real, imag} */,
  {32'h3d87fb0e, 32'h00000000} /* (7, 15, 5) {real, imag} */,
  {32'hbf29f975, 32'h00000000} /* (7, 15, 4) {real, imag} */,
  {32'hbed9a302, 32'h00000000} /* (7, 15, 3) {real, imag} */,
  {32'hbe585369, 32'h00000000} /* (7, 15, 2) {real, imag} */,
  {32'h3deaf2f5, 32'h00000000} /* (7, 15, 1) {real, imag} */,
  {32'h3dbf9fc9, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'h3ea0b1e6, 32'h00000000} /* (7, 14, 15) {real, imag} */,
  {32'h3dcad83d, 32'h00000000} /* (7, 14, 14) {real, imag} */,
  {32'hbef3c4c0, 32'h00000000} /* (7, 14, 13) {real, imag} */,
  {32'hbed3b32a, 32'h00000000} /* (7, 14, 12) {real, imag} */,
  {32'hbcb97dd8, 32'h00000000} /* (7, 14, 11) {real, imag} */,
  {32'hbf20e097, 32'h00000000} /* (7, 14, 10) {real, imag} */,
  {32'hbecacd26, 32'h00000000} /* (7, 14, 9) {real, imag} */,
  {32'h3cb9c2e5, 32'h00000000} /* (7, 14, 8) {real, imag} */,
  {32'hbcecbc96, 32'h00000000} /* (7, 14, 7) {real, imag} */,
  {32'h3eebf23a, 32'h00000000} /* (7, 14, 6) {real, imag} */,
  {32'h3e7eb6cb, 32'h00000000} /* (7, 14, 5) {real, imag} */,
  {32'hbf223192, 32'h00000000} /* (7, 14, 4) {real, imag} */,
  {32'hbe530a80, 32'h00000000} /* (7, 14, 3) {real, imag} */,
  {32'h3cd03c02, 32'h00000000} /* (7, 14, 2) {real, imag} */,
  {32'h3e08cf0a, 32'h00000000} /* (7, 14, 1) {real, imag} */,
  {32'h3e1e7c9a, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hbdcf053f, 32'h00000000} /* (7, 13, 15) {real, imag} */,
  {32'hbe05981b, 32'h00000000} /* (7, 13, 14) {real, imag} */,
  {32'hbe2d0395, 32'h00000000} /* (7, 13, 13) {real, imag} */,
  {32'h3e8d4fbc, 32'h00000000} /* (7, 13, 12) {real, imag} */,
  {32'h3ddba40e, 32'h00000000} /* (7, 13, 11) {real, imag} */,
  {32'hbddfed87, 32'h00000000} /* (7, 13, 10) {real, imag} */,
  {32'h3f20662d, 32'h00000000} /* (7, 13, 9) {real, imag} */,
  {32'h3ea44a9e, 32'h00000000} /* (7, 13, 8) {real, imag} */,
  {32'hbdf5b8ac, 32'h00000000} /* (7, 13, 7) {real, imag} */,
  {32'h3f5e8768, 32'h00000000} /* (7, 13, 6) {real, imag} */,
  {32'h3ea98063, 32'h00000000} /* (7, 13, 5) {real, imag} */,
  {32'hbdd3c806, 32'h00000000} /* (7, 13, 4) {real, imag} */,
  {32'hbdb6098b, 32'h00000000} /* (7, 13, 3) {real, imag} */,
  {32'h3e3eb352, 32'h00000000} /* (7, 13, 2) {real, imag} */,
  {32'h3e58408b, 32'h00000000} /* (7, 13, 1) {real, imag} */,
  {32'h3d25b7be, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'hbc274723, 32'h00000000} /* (7, 12, 15) {real, imag} */,
  {32'h3d6952bf, 32'h00000000} /* (7, 12, 14) {real, imag} */,
  {32'h3e7a419c, 32'h00000000} /* (7, 12, 13) {real, imag} */,
  {32'hbd2c5ea5, 32'h00000000} /* (7, 12, 12) {real, imag} */,
  {32'hbea96618, 32'h00000000} /* (7, 12, 11) {real, imag} */,
  {32'hbe4d6dc1, 32'h00000000} /* (7, 12, 10) {real, imag} */,
  {32'h3efea5ff, 32'h00000000} /* (7, 12, 9) {real, imag} */,
  {32'h3d1cef1a, 32'h00000000} /* (7, 12, 8) {real, imag} */,
  {32'hbe67f0b5, 32'h00000000} /* (7, 12, 7) {real, imag} */,
  {32'hbe19e89a, 32'h00000000} /* (7, 12, 6) {real, imag} */,
  {32'hbe93a7df, 32'h00000000} /* (7, 12, 5) {real, imag} */,
  {32'hbd802e78, 32'h00000000} /* (7, 12, 4) {real, imag} */,
  {32'h3e16ab83, 32'h00000000} /* (7, 12, 3) {real, imag} */,
  {32'h3df949a2, 32'h00000000} /* (7, 12, 2) {real, imag} */,
  {32'hbe0b45bf, 32'h00000000} /* (7, 12, 1) {real, imag} */,
  {32'h3db54eef, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'h3e1fb5af, 32'h00000000} /* (7, 11, 15) {real, imag} */,
  {32'h3ec33552, 32'h00000000} /* (7, 11, 14) {real, imag} */,
  {32'h3e430fe0, 32'h00000000} /* (7, 11, 13) {real, imag} */,
  {32'hbeb0144a, 32'h00000000} /* (7, 11, 12) {real, imag} */,
  {32'hbede3c45, 32'h00000000} /* (7, 11, 11) {real, imag} */,
  {32'hbdddd284, 32'h00000000} /* (7, 11, 10) {real, imag} */,
  {32'h3d9afb50, 32'h00000000} /* (7, 11, 9) {real, imag} */,
  {32'hbd82e03f, 32'h00000000} /* (7, 11, 8) {real, imag} */,
  {32'hbd13bfc1, 32'h00000000} /* (7, 11, 7) {real, imag} */,
  {32'hbeb120b9, 32'h00000000} /* (7, 11, 6) {real, imag} */,
  {32'h3c3ab236, 32'h00000000} /* (7, 11, 5) {real, imag} */,
  {32'h3ea6c79f, 32'h00000000} /* (7, 11, 4) {real, imag} */,
  {32'h3ebec9f1, 32'h00000000} /* (7, 11, 3) {real, imag} */,
  {32'hbdd2ded4, 32'h00000000} /* (7, 11, 2) {real, imag} */,
  {32'hbea3afb8, 32'h00000000} /* (7, 11, 1) {real, imag} */,
  {32'hbdfeb295, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'hbddfcf67, 32'h00000000} /* (7, 10, 15) {real, imag} */,
  {32'hbc24d877, 32'h00000000} /* (7, 10, 14) {real, imag} */,
  {32'h3ea50e1e, 32'h00000000} /* (7, 10, 13) {real, imag} */,
  {32'hbd2d6255, 32'h00000000} /* (7, 10, 12) {real, imag} */,
  {32'hbcc7937a, 32'h00000000} /* (7, 10, 11) {real, imag} */,
  {32'h3ec686a2, 32'h00000000} /* (7, 10, 10) {real, imag} */,
  {32'h3ef95851, 32'h00000000} /* (7, 10, 9) {real, imag} */,
  {32'h3e4eb438, 32'h00000000} /* (7, 10, 8) {real, imag} */,
  {32'hbb18a62d, 32'h00000000} /* (7, 10, 7) {real, imag} */,
  {32'hbc979eaf, 32'h00000000} /* (7, 10, 6) {real, imag} */,
  {32'h3f05e2be, 32'h00000000} /* (7, 10, 5) {real, imag} */,
  {32'h3f48a66f, 32'h00000000} /* (7, 10, 4) {real, imag} */,
  {32'h3f35ffbb, 32'h00000000} /* (7, 10, 3) {real, imag} */,
  {32'h3eb4ae24, 32'h00000000} /* (7, 10, 2) {real, imag} */,
  {32'hbd544b98, 32'h00000000} /* (7, 10, 1) {real, imag} */,
  {32'hbe881f59, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'hbd258eb8, 32'h00000000} /* (7, 9, 15) {real, imag} */,
  {32'hbe4d140f, 32'h00000000} /* (7, 9, 14) {real, imag} */,
  {32'hbd23ec09, 32'h00000000} /* (7, 9, 13) {real, imag} */,
  {32'h3e715e22, 32'h00000000} /* (7, 9, 12) {real, imag} */,
  {32'h3ee7b3bf, 32'h00000000} /* (7, 9, 11) {real, imag} */,
  {32'h3dc3cf54, 32'h00000000} /* (7, 9, 10) {real, imag} */,
  {32'h3e4d9cf2, 32'h00000000} /* (7, 9, 9) {real, imag} */,
  {32'hbc4886ce, 32'h00000000} /* (7, 9, 8) {real, imag} */,
  {32'hbed58bda, 32'h00000000} /* (7, 9, 7) {real, imag} */,
  {32'h3d16b840, 32'h00000000} /* (7, 9, 6) {real, imag} */,
  {32'h3f1b7c9b, 32'h00000000} /* (7, 9, 5) {real, imag} */,
  {32'h3e847c2f, 32'h00000000} /* (7, 9, 4) {real, imag} */,
  {32'h3d959f39, 32'h00000000} /* (7, 9, 3) {real, imag} */,
  {32'h3d9edb90, 32'h00000000} /* (7, 9, 2) {real, imag} */,
  {32'h3ec85ac9, 32'h00000000} /* (7, 9, 1) {real, imag} */,
  {32'hbe0cff73, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'hbc586972, 32'h00000000} /* (7, 8, 15) {real, imag} */,
  {32'hbe30a707, 32'h00000000} /* (7, 8, 14) {real, imag} */,
  {32'h3d8bbae9, 32'h00000000} /* (7, 8, 13) {real, imag} */,
  {32'h3e85cfcc, 32'h00000000} /* (7, 8, 12) {real, imag} */,
  {32'h3e15eec4, 32'h00000000} /* (7, 8, 11) {real, imag} */,
  {32'h3cedf16a, 32'h00000000} /* (7, 8, 10) {real, imag} */,
  {32'h3d8de02f, 32'h00000000} /* (7, 8, 9) {real, imag} */,
  {32'h3c2265d5, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'h3d50a649, 32'h00000000} /* (7, 8, 7) {real, imag} */,
  {32'h3e2c4a5c, 32'h00000000} /* (7, 8, 6) {real, imag} */,
  {32'h3e856ee3, 32'h00000000} /* (7, 8, 5) {real, imag} */,
  {32'hbe1d3fde, 32'h00000000} /* (7, 8, 4) {real, imag} */,
  {32'h3e1c21c5, 32'h00000000} /* (7, 8, 3) {real, imag} */,
  {32'hbd37cd9f, 32'h00000000} /* (7, 8, 2) {real, imag} */,
  {32'h3dc8fb17, 32'h00000000} /* (7, 8, 1) {real, imag} */,
  {32'hbd4c6e48, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'hbe290aa9, 32'h00000000} /* (7, 7, 15) {real, imag} */,
  {32'hbeefc18e, 32'h00000000} /* (7, 7, 14) {real, imag} */,
  {32'hbe1e016b, 32'h00000000} /* (7, 7, 13) {real, imag} */,
  {32'h3d6e0bbc, 32'h00000000} /* (7, 7, 12) {real, imag} */,
  {32'h3e929dac, 32'h00000000} /* (7, 7, 11) {real, imag} */,
  {32'h3ec33222, 32'h00000000} /* (7, 7, 10) {real, imag} */,
  {32'h3cc6a47c, 32'h00000000} /* (7, 7, 9) {real, imag} */,
  {32'hbe842e72, 32'h00000000} /* (7, 7, 8) {real, imag} */,
  {32'hbdcdcb60, 32'h00000000} /* (7, 7, 7) {real, imag} */,
  {32'h3db94944, 32'h00000000} /* (7, 7, 6) {real, imag} */,
  {32'hbe92dd49, 32'h00000000} /* (7, 7, 5) {real, imag} */,
  {32'hbec6dda4, 32'h00000000} /* (7, 7, 4) {real, imag} */,
  {32'h3d2978e9, 32'h00000000} /* (7, 7, 3) {real, imag} */,
  {32'hbd2df8ea, 32'h00000000} /* (7, 7, 2) {real, imag} */,
  {32'hbf0a2165, 32'h00000000} /* (7, 7, 1) {real, imag} */,
  {32'hbea3583e, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'hbec27d3a, 32'h00000000} /* (7, 6, 15) {real, imag} */,
  {32'hbf0f2949, 32'h00000000} /* (7, 6, 14) {real, imag} */,
  {32'hbef025bc, 32'h00000000} /* (7, 6, 13) {real, imag} */,
  {32'hbee55618, 32'h00000000} /* (7, 6, 12) {real, imag} */,
  {32'h3e3be562, 32'h00000000} /* (7, 6, 11) {real, imag} */,
  {32'h3d5a1d68, 32'h00000000} /* (7, 6, 10) {real, imag} */,
  {32'h3eaac678, 32'h00000000} /* (7, 6, 9) {real, imag} */,
  {32'h3e842733, 32'h00000000} /* (7, 6, 8) {real, imag} */,
  {32'hbeac5e00, 32'h00000000} /* (7, 6, 7) {real, imag} */,
  {32'h3d061e6c, 32'h00000000} /* (7, 6, 6) {real, imag} */,
  {32'hbd00d68c, 32'h00000000} /* (7, 6, 5) {real, imag} */,
  {32'h3d2b8e70, 32'h00000000} /* (7, 6, 4) {real, imag} */,
  {32'hbed45b42, 32'h00000000} /* (7, 6, 3) {real, imag} */,
  {32'hbea17362, 32'h00000000} /* (7, 6, 2) {real, imag} */,
  {32'h3e0a273f, 32'h00000000} /* (7, 6, 1) {real, imag} */,
  {32'h3d681c5b, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'hbe91ba0f, 32'h00000000} /* (7, 5, 15) {real, imag} */,
  {32'hbe861a79, 32'h00000000} /* (7, 5, 14) {real, imag} */,
  {32'hbe383fef, 32'h00000000} /* (7, 5, 13) {real, imag} */,
  {32'hbea41097, 32'h00000000} /* (7, 5, 12) {real, imag} */,
  {32'hbd67fdd7, 32'h00000000} /* (7, 5, 11) {real, imag} */,
  {32'hbea0c618, 32'h00000000} /* (7, 5, 10) {real, imag} */,
  {32'h3f0084fe, 32'h00000000} /* (7, 5, 9) {real, imag} */,
  {32'h3e0e3540, 32'h00000000} /* (7, 5, 8) {real, imag} */,
  {32'h3dc1b851, 32'h00000000} /* (7, 5, 7) {real, imag} */,
  {32'h3eddf2c3, 32'h00000000} /* (7, 5, 6) {real, imag} */,
  {32'h3f02382c, 32'h00000000} /* (7, 5, 5) {real, imag} */,
  {32'h3f2a6d73, 32'h00000000} /* (7, 5, 4) {real, imag} */,
  {32'hbe8c5139, 32'h00000000} /* (7, 5, 3) {real, imag} */,
  {32'hbee258bf, 32'h00000000} /* (7, 5, 2) {real, imag} */,
  {32'h3c4ff3fc, 32'h00000000} /* (7, 5, 1) {real, imag} */,
  {32'h3d2c4a66, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'hbea7b773, 32'h00000000} /* (7, 4, 15) {real, imag} */,
  {32'h3e92b366, 32'h00000000} /* (7, 4, 14) {real, imag} */,
  {32'h3ee2b1c1, 32'h00000000} /* (7, 4, 13) {real, imag} */,
  {32'h3e59c470, 32'h00000000} /* (7, 4, 12) {real, imag} */,
  {32'h3e8ba3ab, 32'h00000000} /* (7, 4, 11) {real, imag} */,
  {32'hbe3f60ff, 32'h00000000} /* (7, 4, 10) {real, imag} */,
  {32'h3f4eff82, 32'h00000000} /* (7, 4, 9) {real, imag} */,
  {32'h3dfec397, 32'h00000000} /* (7, 4, 8) {real, imag} */,
  {32'hbd1db7c8, 32'h00000000} /* (7, 4, 7) {real, imag} */,
  {32'h3f1b8118, 32'h00000000} /* (7, 4, 6) {real, imag} */,
  {32'h3f438d60, 32'h00000000} /* (7, 4, 5) {real, imag} */,
  {32'h3f3f80b4, 32'h00000000} /* (7, 4, 4) {real, imag} */,
  {32'hbdc143f0, 32'h00000000} /* (7, 4, 3) {real, imag} */,
  {32'hbf24ea36, 32'h00000000} /* (7, 4, 2) {real, imag} */,
  {32'hbe3cd518, 32'h00000000} /* (7, 4, 1) {real, imag} */,
  {32'h3ce79640, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'hbe1d67f2, 32'h00000000} /* (7, 3, 15) {real, imag} */,
  {32'h3f2c2962, 32'h00000000} /* (7, 3, 14) {real, imag} */,
  {32'h3f4eaf27, 32'h00000000} /* (7, 3, 13) {real, imag} */,
  {32'h3e88efc8, 32'h00000000} /* (7, 3, 12) {real, imag} */,
  {32'h3f0acb20, 32'h00000000} /* (7, 3, 11) {real, imag} */,
  {32'hbcf3838d, 32'h00000000} /* (7, 3, 10) {real, imag} */,
  {32'hbd7a2bd8, 32'h00000000} /* (7, 3, 9) {real, imag} */,
  {32'hbc20be64, 32'h00000000} /* (7, 3, 8) {real, imag} */,
  {32'h3dab258e, 32'h00000000} /* (7, 3, 7) {real, imag} */,
  {32'h3efa37e0, 32'h00000000} /* (7, 3, 6) {real, imag} */,
  {32'h3f395bc6, 32'h00000000} /* (7, 3, 5) {real, imag} */,
  {32'h3ccb5857, 32'h00000000} /* (7, 3, 4) {real, imag} */,
  {32'hbe7aace8, 32'h00000000} /* (7, 3, 3) {real, imag} */,
  {32'hbe8a1ab1, 32'h00000000} /* (7, 3, 2) {real, imag} */,
  {32'hbecf7d3f, 32'h00000000} /* (7, 3, 1) {real, imag} */,
  {32'hbe1d8e9b, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'h3df22405, 32'h00000000} /* (7, 2, 15) {real, imag} */,
  {32'h3d62f54e, 32'h00000000} /* (7, 2, 14) {real, imag} */,
  {32'h3e7166ea, 32'h00000000} /* (7, 2, 13) {real, imag} */,
  {32'h3eb1de2d, 32'h00000000} /* (7, 2, 12) {real, imag} */,
  {32'hbe144c31, 32'h00000000} /* (7, 2, 11) {real, imag} */,
  {32'hbed93c33, 32'h00000000} /* (7, 2, 10) {real, imag} */,
  {32'hbec99ac7, 32'h00000000} /* (7, 2, 9) {real, imag} */,
  {32'hbf03c3d3, 32'h00000000} /* (7, 2, 8) {real, imag} */,
  {32'hbd80ba6f, 32'h00000000} /* (7, 2, 7) {real, imag} */,
  {32'h3ef4a84c, 32'h00000000} /* (7, 2, 6) {real, imag} */,
  {32'h3ed13080, 32'h00000000} /* (7, 2, 5) {real, imag} */,
  {32'h3e090d19, 32'h00000000} /* (7, 2, 4) {real, imag} */,
  {32'hbd9fdaeb, 32'h00000000} /* (7, 2, 3) {real, imag} */,
  {32'hbedec0f1, 32'h00000000} /* (7, 2, 2) {real, imag} */,
  {32'hbf649d8b, 32'h00000000} /* (7, 2, 1) {real, imag} */,
  {32'hbea4fd7c, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h3e6c1e25, 32'h00000000} /* (7, 1, 15) {real, imag} */,
  {32'hbdb99a81, 32'h00000000} /* (7, 1, 14) {real, imag} */,
  {32'hbe0ef177, 32'h00000000} /* (7, 1, 13) {real, imag} */,
  {32'h3e9dbd30, 32'h00000000} /* (7, 1, 12) {real, imag} */,
  {32'hbeea907c, 32'h00000000} /* (7, 1, 11) {real, imag} */,
  {32'hbe9572d5, 32'h00000000} /* (7, 1, 10) {real, imag} */,
  {32'hbcfd456e, 32'h00000000} /* (7, 1, 9) {real, imag} */,
  {32'hbee4b400, 32'h00000000} /* (7, 1, 8) {real, imag} */,
  {32'h3dd19c94, 32'h00000000} /* (7, 1, 7) {real, imag} */,
  {32'h3ec534ac, 32'h00000000} /* (7, 1, 6) {real, imag} */,
  {32'h3eb46960, 32'h00000000} /* (7, 1, 5) {real, imag} */,
  {32'h3f25103e, 32'h00000000} /* (7, 1, 4) {real, imag} */,
  {32'h3e8580f9, 32'h00000000} /* (7, 1, 3) {real, imag} */,
  {32'hbebadbd4, 32'h00000000} /* (7, 1, 2) {real, imag} */,
  {32'hbf35d63c, 32'h00000000} /* (7, 1, 1) {real, imag} */,
  {32'hbd5a6496, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'hbd621877, 32'h00000000} /* (7, 0, 15) {real, imag} */,
  {32'hbe20039c, 32'h00000000} /* (7, 0, 14) {real, imag} */,
  {32'hbddf4d2c, 32'h00000000} /* (7, 0, 13) {real, imag} */,
  {32'h3dcc7c3b, 32'h00000000} /* (7, 0, 12) {real, imag} */,
  {32'h3ca02ef4, 32'h00000000} /* (7, 0, 11) {real, imag} */,
  {32'h3d1706bd, 32'h00000000} /* (7, 0, 10) {real, imag} */,
  {32'h3ea847ad, 32'h00000000} /* (7, 0, 9) {real, imag} */,
  {32'h3dd4cee8, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'h3d38c910, 32'h00000000} /* (7, 0, 7) {real, imag} */,
  {32'h3e6e0472, 32'h00000000} /* (7, 0, 6) {real, imag} */,
  {32'h3ebabad6, 32'h00000000} /* (7, 0, 5) {real, imag} */,
  {32'h3e510c45, 32'h00000000} /* (7, 0, 4) {real, imag} */,
  {32'h3c9827bd, 32'h00000000} /* (7, 0, 3) {real, imag} */,
  {32'h3c04f2b0, 32'h00000000} /* (7, 0, 2) {real, imag} */,
  {32'h3d6f62fb, 32'h00000000} /* (7, 0, 1) {real, imag} */,
  {32'h3e8f4c22, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'hbcc9038b, 32'h00000000} /* (6, 15, 15) {real, imag} */,
  {32'h3c7546e4, 32'h00000000} /* (6, 15, 14) {real, imag} */,
  {32'hbe4609b7, 32'h00000000} /* (6, 15, 13) {real, imag} */,
  {32'hbe3ed581, 32'h00000000} /* (6, 15, 12) {real, imag} */,
  {32'hbd90e3b2, 32'h00000000} /* (6, 15, 11) {real, imag} */,
  {32'hbdc41f5b, 32'h00000000} /* (6, 15, 10) {real, imag} */,
  {32'h3d525d47, 32'h00000000} /* (6, 15, 9) {real, imag} */,
  {32'h3e59c180, 32'h00000000} /* (6, 15, 8) {real, imag} */,
  {32'h3c799537, 32'h00000000} /* (6, 15, 7) {real, imag} */,
  {32'hbd03b689, 32'h00000000} /* (6, 15, 6) {real, imag} */,
  {32'hbe32d45c, 32'h00000000} /* (6, 15, 5) {real, imag} */,
  {32'hbeccfd7d, 32'h00000000} /* (6, 15, 4) {real, imag} */,
  {32'hbe161ac0, 32'h00000000} /* (6, 15, 3) {real, imag} */,
  {32'hbe655574, 32'h00000000} /* (6, 15, 2) {real, imag} */,
  {32'h3d2e3384, 32'h00000000} /* (6, 15, 1) {real, imag} */,
  {32'h3e5bec84, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'h3c34cc35, 32'h00000000} /* (6, 14, 15) {real, imag} */,
  {32'hbe810ade, 32'h00000000} /* (6, 14, 14) {real, imag} */,
  {32'hbee87d7a, 32'h00000000} /* (6, 14, 13) {real, imag} */,
  {32'hbe831e08, 32'h00000000} /* (6, 14, 12) {real, imag} */,
  {32'h3b3e2cc9, 32'h00000000} /* (6, 14, 11) {real, imag} */,
  {32'hbde85d30, 32'h00000000} /* (6, 14, 10) {real, imag} */,
  {32'h3c984989, 32'h00000000} /* (6, 14, 9) {real, imag} */,
  {32'h3dd5f023, 32'h00000000} /* (6, 14, 8) {real, imag} */,
  {32'hba8853ba, 32'h00000000} /* (6, 14, 7) {real, imag} */,
  {32'h3dd97b50, 32'h00000000} /* (6, 14, 6) {real, imag} */,
  {32'hbe6514ab, 32'h00000000} /* (6, 14, 5) {real, imag} */,
  {32'hbeb9f42a, 32'h00000000} /* (6, 14, 4) {real, imag} */,
  {32'hbe333b99, 32'h00000000} /* (6, 14, 3) {real, imag} */,
  {32'hbe8e98b1, 32'h00000000} /* (6, 14, 2) {real, imag} */,
  {32'h3e0d07ca, 32'h00000000} /* (6, 14, 1) {real, imag} */,
  {32'h3ea7eb87, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hbe48d5ae, 32'h00000000} /* (6, 13, 15) {real, imag} */,
  {32'hbe468680, 32'h00000000} /* (6, 13, 14) {real, imag} */,
  {32'hbe9532e8, 32'h00000000} /* (6, 13, 13) {real, imag} */,
  {32'hbebe75e0, 32'h00000000} /* (6, 13, 12) {real, imag} */,
  {32'h3d81b33e, 32'h00000000} /* (6, 13, 11) {real, imag} */,
  {32'h3edaf08b, 32'h00000000} /* (6, 13, 10) {real, imag} */,
  {32'h3de22575, 32'h00000000} /* (6, 13, 9) {real, imag} */,
  {32'hbe0e525e, 32'h00000000} /* (6, 13, 8) {real, imag} */,
  {32'h3d0b6513, 32'h00000000} /* (6, 13, 7) {real, imag} */,
  {32'h3e564fd7, 32'h00000000} /* (6, 13, 6) {real, imag} */,
  {32'hbe999a45, 32'h00000000} /* (6, 13, 5) {real, imag} */,
  {32'hbf013e53, 32'h00000000} /* (6, 13, 4) {real, imag} */,
  {32'hbe5e5d41, 32'h00000000} /* (6, 13, 3) {real, imag} */,
  {32'hbcf4d620, 32'h00000000} /* (6, 13, 2) {real, imag} */,
  {32'hbdadef96, 32'h00000000} /* (6, 13, 1) {real, imag} */,
  {32'hbe55be48, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'h3ca04648, 32'h00000000} /* (6, 12, 15) {real, imag} */,
  {32'h3d0073b7, 32'h00000000} /* (6, 12, 14) {real, imag} */,
  {32'h3d80d3d4, 32'h00000000} /* (6, 12, 13) {real, imag} */,
  {32'hbea42ffa, 32'h00000000} /* (6, 12, 12) {real, imag} */,
  {32'h3c556938, 32'h00000000} /* (6, 12, 11) {real, imag} */,
  {32'hbda2ecf5, 32'h00000000} /* (6, 12, 10) {real, imag} */,
  {32'hbe0b93a4, 32'h00000000} /* (6, 12, 9) {real, imag} */,
  {32'h3e0f70e8, 32'h00000000} /* (6, 12, 8) {real, imag} */,
  {32'hbd83839e, 32'h00000000} /* (6, 12, 7) {real, imag} */,
  {32'h3c3ae31a, 32'h00000000} /* (6, 12, 6) {real, imag} */,
  {32'hbe324e6d, 32'h00000000} /* (6, 12, 5) {real, imag} */,
  {32'h3d088972, 32'h00000000} /* (6, 12, 4) {real, imag} */,
  {32'h3e715317, 32'h00000000} /* (6, 12, 3) {real, imag} */,
  {32'hbd91d8fd, 32'h00000000} /* (6, 12, 2) {real, imag} */,
  {32'hbe890e44, 32'h00000000} /* (6, 12, 1) {real, imag} */,
  {32'hbe0e9842, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'h3f359573, 32'h00000000} /* (6, 11, 15) {real, imag} */,
  {32'h3f2345b6, 32'h00000000} /* (6, 11, 14) {real, imag} */,
  {32'hbe62fb70, 32'h00000000} /* (6, 11, 13) {real, imag} */,
  {32'hbdda892f, 32'h00000000} /* (6, 11, 12) {real, imag} */,
  {32'hbea204db, 32'h00000000} /* (6, 11, 11) {real, imag} */,
  {32'hbf17aa22, 32'h00000000} /* (6, 11, 10) {real, imag} */,
  {32'hbed34ad4, 32'h00000000} /* (6, 11, 9) {real, imag} */,
  {32'hbdf154b0, 32'h00000000} /* (6, 11, 8) {real, imag} */,
  {32'hbe861818, 32'h00000000} /* (6, 11, 7) {real, imag} */,
  {32'hbb1217a3, 32'h00000000} /* (6, 11, 6) {real, imag} */,
  {32'h3e2ba49e, 32'h00000000} /* (6, 11, 5) {real, imag} */,
  {32'h3ec726f5, 32'h00000000} /* (6, 11, 4) {real, imag} */,
  {32'h3f249f8b, 32'h00000000} /* (6, 11, 3) {real, imag} */,
  {32'hbd001614, 32'h00000000} /* (6, 11, 2) {real, imag} */,
  {32'h3dd8684b, 32'h00000000} /* (6, 11, 1) {real, imag} */,
  {32'h3d934239, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h3ef3e06c, 32'h00000000} /* (6, 10, 15) {real, imag} */,
  {32'h3d2ea6b7, 32'h00000000} /* (6, 10, 14) {real, imag} */,
  {32'hbf09f7e1, 32'h00000000} /* (6, 10, 13) {real, imag} */,
  {32'hbe1eaf0b, 32'h00000000} /* (6, 10, 12) {real, imag} */,
  {32'hbd7cee54, 32'h00000000} /* (6, 10, 11) {real, imag} */,
  {32'hbe16dffe, 32'h00000000} /* (6, 10, 10) {real, imag} */,
  {32'h3e2a2e4f, 32'h00000000} /* (6, 10, 9) {real, imag} */,
  {32'h3d64ef31, 32'h00000000} /* (6, 10, 8) {real, imag} */,
  {32'hbe0a9b99, 32'h00000000} /* (6, 10, 7) {real, imag} */,
  {32'hbb1eea27, 32'h00000000} /* (6, 10, 6) {real, imag} */,
  {32'h3eba27d3, 32'h00000000} /* (6, 10, 5) {real, imag} */,
  {32'h3f7635f3, 32'h00000000} /* (6, 10, 4) {real, imag} */,
  {32'h3f90bbaa, 32'h00000000} /* (6, 10, 3) {real, imag} */,
  {32'h3ee4c70c, 32'h00000000} /* (6, 10, 2) {real, imag} */,
  {32'h3ed247d5, 32'h00000000} /* (6, 10, 1) {real, imag} */,
  {32'h3e003bc8, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h3f0e72f7, 32'h00000000} /* (6, 9, 15) {real, imag} */,
  {32'hbe402fe2, 32'h00000000} /* (6, 9, 14) {real, imag} */,
  {32'hbf16d236, 32'h00000000} /* (6, 9, 13) {real, imag} */,
  {32'hbc61da10, 32'h00000000} /* (6, 9, 12) {real, imag} */,
  {32'h3f06cb92, 32'h00000000} /* (6, 9, 11) {real, imag} */,
  {32'h3e8b326c, 32'h00000000} /* (6, 9, 10) {real, imag} */,
  {32'h3f272569, 32'h00000000} /* (6, 9, 9) {real, imag} */,
  {32'h3f1d2000, 32'h00000000} /* (6, 9, 8) {real, imag} */,
  {32'h3eac3d0d, 32'h00000000} /* (6, 9, 7) {real, imag} */,
  {32'h3de5a40c, 32'h00000000} /* (6, 9, 6) {real, imag} */,
  {32'h3ec0738e, 32'h00000000} /* (6, 9, 5) {real, imag} */,
  {32'h3ed0b822, 32'h00000000} /* (6, 9, 4) {real, imag} */,
  {32'h3e810fc8, 32'h00000000} /* (6, 9, 3) {real, imag} */,
  {32'h3e9561f4, 32'h00000000} /* (6, 9, 2) {real, imag} */,
  {32'h3e97047e, 32'h00000000} /* (6, 9, 1) {real, imag} */,
  {32'hbdefda37, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h3f129f22, 32'h00000000} /* (6, 8, 15) {real, imag} */,
  {32'hbdff0c88, 32'h00000000} /* (6, 8, 14) {real, imag} */,
  {32'hbf2a21a1, 32'h00000000} /* (6, 8, 13) {real, imag} */,
  {32'hbe96a32f, 32'h00000000} /* (6, 8, 12) {real, imag} */,
  {32'hbcac065a, 32'h00000000} /* (6, 8, 11) {real, imag} */,
  {32'h3dd76d13, 32'h00000000} /* (6, 8, 10) {real, imag} */,
  {32'h3e80f4bc, 32'h00000000} /* (6, 8, 9) {real, imag} */,
  {32'h3ddf620b, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'h3ed4a521, 32'h00000000} /* (6, 8, 7) {real, imag} */,
  {32'h3e5975aa, 32'h00000000} /* (6, 8, 6) {real, imag} */,
  {32'h3e4a36a8, 32'h00000000} /* (6, 8, 5) {real, imag} */,
  {32'hbd348772, 32'h00000000} /* (6, 8, 4) {real, imag} */,
  {32'h3e4c1f01, 32'h00000000} /* (6, 8, 3) {real, imag} */,
  {32'h3d2aa448, 32'h00000000} /* (6, 8, 2) {real, imag} */,
  {32'hbe119765, 32'h00000000} /* (6, 8, 1) {real, imag} */,
  {32'hbcfb2d46, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h3dd3921c, 32'h00000000} /* (6, 7, 15) {real, imag} */,
  {32'hbebe994d, 32'h00000000} /* (6, 7, 14) {real, imag} */,
  {32'hbf334c9a, 32'h00000000} /* (6, 7, 13) {real, imag} */,
  {32'hbf6707b3, 32'h00000000} /* (6, 7, 12) {real, imag} */,
  {32'hbee958f9, 32'h00000000} /* (6, 7, 11) {real, imag} */,
  {32'hbb43f47c, 32'h00000000} /* (6, 7, 10) {real, imag} */,
  {32'hbea43068, 32'h00000000} /* (6, 7, 9) {real, imag} */,
  {32'hbf0dc554, 32'h00000000} /* (6, 7, 8) {real, imag} */,
  {32'hbdcb407d, 32'h00000000} /* (6, 7, 7) {real, imag} */,
  {32'h3dba9de6, 32'h00000000} /* (6, 7, 6) {real, imag} */,
  {32'hbeb2cbbf, 32'h00000000} /* (6, 7, 5) {real, imag} */,
  {32'hbe951adb, 32'h00000000} /* (6, 7, 4) {real, imag} */,
  {32'h3ef15973, 32'h00000000} /* (6, 7, 3) {real, imag} */,
  {32'h3ed0f37f, 32'h00000000} /* (6, 7, 2) {real, imag} */,
  {32'h3eb0d71c, 32'h00000000} /* (6, 7, 1) {real, imag} */,
  {32'h3e7ce46c, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'hbd8b737e, 32'h00000000} /* (6, 6, 15) {real, imag} */,
  {32'hbe8881c8, 32'h00000000} /* (6, 6, 14) {real, imag} */,
  {32'hbefd30aa, 32'h00000000} /* (6, 6, 13) {real, imag} */,
  {32'hbf462c0c, 32'h00000000} /* (6, 6, 12) {real, imag} */,
  {32'h3dac0906, 32'h00000000} /* (6, 6, 11) {real, imag} */,
  {32'h3e4b1839, 32'h00000000} /* (6, 6, 10) {real, imag} */,
  {32'hbe8e021c, 32'h00000000} /* (6, 6, 9) {real, imag} */,
  {32'hbe80b250, 32'h00000000} /* (6, 6, 8) {real, imag} */,
  {32'hbdc6eff7, 32'h00000000} /* (6, 6, 7) {real, imag} */,
  {32'h3e184725, 32'h00000000} /* (6, 6, 6) {real, imag} */,
  {32'hbe6fcbc7, 32'h00000000} /* (6, 6, 5) {real, imag} */,
  {32'hbe6cdbf8, 32'h00000000} /* (6, 6, 4) {real, imag} */,
  {32'hbd829b07, 32'h00000000} /* (6, 6, 3) {real, imag} */,
  {32'h3df0acfe, 32'h00000000} /* (6, 6, 2) {real, imag} */,
  {32'h3e75fbeb, 32'h00000000} /* (6, 6, 1) {real, imag} */,
  {32'h3e9e2757, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'hbea05cfb, 32'h00000000} /* (6, 5, 15) {real, imag} */,
  {32'hbe51d628, 32'h00000000} /* (6, 5, 14) {real, imag} */,
  {32'hbe08c20a, 32'h00000000} /* (6, 5, 13) {real, imag} */,
  {32'hbf008ab6, 32'h00000000} /* (6, 5, 12) {real, imag} */,
  {32'hbe6e9da0, 32'h00000000} /* (6, 5, 11) {real, imag} */,
  {32'hbe950884, 32'h00000000} /* (6, 5, 10) {real, imag} */,
  {32'h3d5a753a, 32'h00000000} /* (6, 5, 9) {real, imag} */,
  {32'h3d8980d5, 32'h00000000} /* (6, 5, 8) {real, imag} */,
  {32'h3e6c99ee, 32'h00000000} /* (6, 5, 7) {real, imag} */,
  {32'h3eb98070, 32'h00000000} /* (6, 5, 6) {real, imag} */,
  {32'h3dbdb099, 32'h00000000} /* (6, 5, 5) {real, imag} */,
  {32'h3abfc3c4, 32'h00000000} /* (6, 5, 4) {real, imag} */,
  {32'hbf114879, 32'h00000000} /* (6, 5, 3) {real, imag} */,
  {32'hbee43656, 32'h00000000} /* (6, 5, 2) {real, imag} */,
  {32'hbec94b9e, 32'h00000000} /* (6, 5, 1) {real, imag} */,
  {32'hbab552d6, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'hbd2fec84, 32'h00000000} /* (6, 4, 15) {real, imag} */,
  {32'h3ec23336, 32'h00000000} /* (6, 4, 14) {real, imag} */,
  {32'h3e84e940, 32'h00000000} /* (6, 4, 13) {real, imag} */,
  {32'hbcd09b2c, 32'h00000000} /* (6, 4, 12) {real, imag} */,
  {32'hbd9e9b15, 32'h00000000} /* (6, 4, 11) {real, imag} */,
  {32'hbd653965, 32'h00000000} /* (6, 4, 10) {real, imag} */,
  {32'h3eee5e1e, 32'h00000000} /* (6, 4, 9) {real, imag} */,
  {32'hb8337430, 32'h00000000} /* (6, 4, 8) {real, imag} */,
  {32'hbe754fca, 32'h00000000} /* (6, 4, 7) {real, imag} */,
  {32'h3e7a06ff, 32'h00000000} /* (6, 4, 6) {real, imag} */,
  {32'h3f0d6f82, 32'h00000000} /* (6, 4, 5) {real, imag} */,
  {32'h3e0b4c48, 32'h00000000} /* (6, 4, 4) {real, imag} */,
  {32'hbf5f25c0, 32'h00000000} /* (6, 4, 3) {real, imag} */,
  {32'hbed25452, 32'h00000000} /* (6, 4, 2) {real, imag} */,
  {32'hbbaf2fb6, 32'h00000000} /* (6, 4, 1) {real, imag} */,
  {32'hbb9a835f, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'hbe49155a, 32'h00000000} /* (6, 3, 15) {real, imag} */,
  {32'h3efb774c, 32'h00000000} /* (6, 3, 14) {real, imag} */,
  {32'h3f4394d3, 32'h00000000} /* (6, 3, 13) {real, imag} */,
  {32'hbdbe5c7a, 32'h00000000} /* (6, 3, 12) {real, imag} */,
  {32'h3f0ec032, 32'h00000000} /* (6, 3, 11) {real, imag} */,
  {32'h3d928a4b, 32'h00000000} /* (6, 3, 10) {real, imag} */,
  {32'hbe1ca11c, 32'h00000000} /* (6, 3, 9) {real, imag} */,
  {32'hbe80a9de, 32'h00000000} /* (6, 3, 8) {real, imag} */,
  {32'hbecbea93, 32'h00000000} /* (6, 3, 7) {real, imag} */,
  {32'hbe0a5bda, 32'h00000000} /* (6, 3, 6) {real, imag} */,
  {32'h3e42300a, 32'h00000000} /* (6, 3, 5) {real, imag} */,
  {32'hbf0731ee, 32'h00000000} /* (6, 3, 4) {real, imag} */,
  {32'hbf12ff0c, 32'h00000000} /* (6, 3, 3) {real, imag} */,
  {32'h3de6d968, 32'h00000000} /* (6, 3, 2) {real, imag} */,
  {32'h3e0d4f78, 32'h00000000} /* (6, 3, 1) {real, imag} */,
  {32'hbd194662, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'hbede1c52, 32'h00000000} /* (6, 2, 15) {real, imag} */,
  {32'hbe212282, 32'h00000000} /* (6, 2, 14) {real, imag} */,
  {32'h3eb0ff98, 32'h00000000} /* (6, 2, 13) {real, imag} */,
  {32'hbe4c4be5, 32'h00000000} /* (6, 2, 12) {real, imag} */,
  {32'hbe49be42, 32'h00000000} /* (6, 2, 11) {real, imag} */,
  {32'hbf2d311f, 32'h00000000} /* (6, 2, 10) {real, imag} */,
  {32'hbea8b042, 32'h00000000} /* (6, 2, 9) {real, imag} */,
  {32'hbec76300, 32'h00000000} /* (6, 2, 8) {real, imag} */,
  {32'h3d30f39e, 32'h00000000} /* (6, 2, 7) {real, imag} */,
  {32'h3e397e35, 32'h00000000} /* (6, 2, 6) {real, imag} */,
  {32'hbe2c46d2, 32'h00000000} /* (6, 2, 5) {real, imag} */,
  {32'h3e1632f7, 32'h00000000} /* (6, 2, 4) {real, imag} */,
  {32'h3e9b8ba6, 32'h00000000} /* (6, 2, 3) {real, imag} */,
  {32'hbd4e070a, 32'h00000000} /* (6, 2, 2) {real, imag} */,
  {32'hbeeeef67, 32'h00000000} /* (6, 2, 1) {real, imag} */,
  {32'hbea6866e, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'hbe852708, 32'h00000000} /* (6, 1, 15) {real, imag} */,
  {32'h3e22ff63, 32'h00000000} /* (6, 1, 14) {real, imag} */,
  {32'h3e9c0cce, 32'h00000000} /* (6, 1, 13) {real, imag} */,
  {32'hbe0c963e, 32'h00000000} /* (6, 1, 12) {real, imag} */,
  {32'hbf530306, 32'h00000000} /* (6, 1, 11) {real, imag} */,
  {32'hbedeb70e, 32'h00000000} /* (6, 1, 10) {real, imag} */,
  {32'h3e725096, 32'h00000000} /* (6, 1, 9) {real, imag} */,
  {32'hbe21b5f0, 32'h00000000} /* (6, 1, 8) {real, imag} */,
  {32'hbeebe081, 32'h00000000} /* (6, 1, 7) {real, imag} */,
  {32'hbe36d943, 32'h00000000} /* (6, 1, 6) {real, imag} */,
  {32'h3ec01fdc, 32'h00000000} /* (6, 1, 5) {real, imag} */,
  {32'h3f8b986b, 32'h00000000} /* (6, 1, 4) {real, imag} */,
  {32'h3f00ceeb, 32'h00000000} /* (6, 1, 3) {real, imag} */,
  {32'hbe4c8b8c, 32'h00000000} /* (6, 1, 2) {real, imag} */,
  {32'hbf03d02a, 32'h00000000} /* (6, 1, 1) {real, imag} */,
  {32'hbeb3a7a6, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'hbcf10760, 32'h00000000} /* (6, 0, 15) {real, imag} */,
  {32'h3dc60dad, 32'h00000000} /* (6, 0, 14) {real, imag} */,
  {32'h3d7c9d55, 32'h00000000} /* (6, 0, 13) {real, imag} */,
  {32'hbd9a00d7, 32'h00000000} /* (6, 0, 12) {real, imag} */,
  {32'hbe7113cd, 32'h00000000} /* (6, 0, 11) {real, imag} */,
  {32'hbdb66f47, 32'h00000000} /* (6, 0, 10) {real, imag} */,
  {32'h3e40fdb5, 32'h00000000} /* (6, 0, 9) {real, imag} */,
  {32'h3df4382c, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'hbe8d2693, 32'h00000000} /* (6, 0, 7) {real, imag} */,
  {32'hbe50ffe1, 32'h00000000} /* (6, 0, 6) {real, imag} */,
  {32'h3ef32646, 32'h00000000} /* (6, 0, 5) {real, imag} */,
  {32'h3ebea95d, 32'h00000000} /* (6, 0, 4) {real, imag} */,
  {32'h3d36d1f1, 32'h00000000} /* (6, 0, 3) {real, imag} */,
  {32'hbd03e6f2, 32'h00000000} /* (6, 0, 2) {real, imag} */,
  {32'hbc68f02a, 32'h00000000} /* (6, 0, 1) {real, imag} */,
  {32'h3dec9e1e, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'hbf1164d2, 32'h00000000} /* (5, 15, 15) {real, imag} */,
  {32'hbea24b09, 32'h00000000} /* (5, 15, 14) {real, imag} */,
  {32'hbc94d28c, 32'h00000000} /* (5, 15, 13) {real, imag} */,
  {32'hbd3e1db2, 32'h00000000} /* (5, 15, 12) {real, imag} */,
  {32'hbe7ae64a, 32'h00000000} /* (5, 15, 11) {real, imag} */,
  {32'hbe23f88c, 32'h00000000} /* (5, 15, 10) {real, imag} */,
  {32'hbc22af71, 32'h00000000} /* (5, 15, 9) {real, imag} */,
  {32'hbd5b6a7c, 32'h00000000} /* (5, 15, 8) {real, imag} */,
  {32'hbe34822a, 32'h00000000} /* (5, 15, 7) {real, imag} */,
  {32'hbda588dc, 32'h00000000} /* (5, 15, 6) {real, imag} */,
  {32'h3e07db0e, 32'h00000000} /* (5, 15, 5) {real, imag} */,
  {32'h3ec3b0ad, 32'h00000000} /* (5, 15, 4) {real, imag} */,
  {32'h3d2a021a, 32'h00000000} /* (5, 15, 3) {real, imag} */,
  {32'hbecb91df, 32'h00000000} /* (5, 15, 2) {real, imag} */,
  {32'h3c1c1510, 32'h00000000} /* (5, 15, 1) {real, imag} */,
  {32'h3e80fce5, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hbeb3570f, 32'h00000000} /* (5, 14, 15) {real, imag} */,
  {32'hbea7ebbc, 32'h00000000} /* (5, 14, 14) {real, imag} */,
  {32'hbed90d72, 32'h00000000} /* (5, 14, 13) {real, imag} */,
  {32'hbece4ef9, 32'h00000000} /* (5, 14, 12) {real, imag} */,
  {32'hbe2174ba, 32'h00000000} /* (5, 14, 11) {real, imag} */,
  {32'hbe3b9f1b, 32'h00000000} /* (5, 14, 10) {real, imag} */,
  {32'hbdb387d9, 32'h00000000} /* (5, 14, 9) {real, imag} */,
  {32'hbe6d5d18, 32'h00000000} /* (5, 14, 8) {real, imag} */,
  {32'h3a0de628, 32'h00000000} /* (5, 14, 7) {real, imag} */,
  {32'h3d922312, 32'h00000000} /* (5, 14, 6) {real, imag} */,
  {32'hbe0c24a4, 32'h00000000} /* (5, 14, 5) {real, imag} */,
  {32'hbda47536, 32'h00000000} /* (5, 14, 4) {real, imag} */,
  {32'hbeaf0221, 32'h00000000} /* (5, 14, 3) {real, imag} */,
  {32'hbf437175, 32'h00000000} /* (5, 14, 2) {real, imag} */,
  {32'h3e3dee45, 32'h00000000} /* (5, 14, 1) {real, imag} */,
  {32'h3f28fa73, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hbe3906c9, 32'h00000000} /* (5, 13, 15) {real, imag} */,
  {32'hbde976ea, 32'h00000000} /* (5, 13, 14) {real, imag} */,
  {32'hbe91d685, 32'h00000000} /* (5, 13, 13) {real, imag} */,
  {32'hbf2ec472, 32'h00000000} /* (5, 13, 12) {real, imag} */,
  {32'hbea0dabe, 32'h00000000} /* (5, 13, 11) {real, imag} */,
  {32'hbbb5ca4a, 32'h00000000} /* (5, 13, 10) {real, imag} */,
  {32'hbedf63b2, 32'h00000000} /* (5, 13, 9) {real, imag} */,
  {32'hbe70a868, 32'h00000000} /* (5, 13, 8) {real, imag} */,
  {32'h3e355025, 32'h00000000} /* (5, 13, 7) {real, imag} */,
  {32'hbe005223, 32'h00000000} /* (5, 13, 6) {real, imag} */,
  {32'hbf195b90, 32'h00000000} /* (5, 13, 5) {real, imag} */,
  {32'hbf3f605e, 32'h00000000} /* (5, 13, 4) {real, imag} */,
  {32'hbe1299b9, 32'h00000000} /* (5, 13, 3) {real, imag} */,
  {32'hbe961449, 32'h00000000} /* (5, 13, 2) {real, imag} */,
  {32'hbeef1e1b, 32'h00000000} /* (5, 13, 1) {real, imag} */,
  {32'hbe546d64, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'hbe108666, 32'h00000000} /* (5, 12, 15) {real, imag} */,
  {32'h3e8bc9ea, 32'h00000000} /* (5, 12, 14) {real, imag} */,
  {32'h3e781604, 32'h00000000} /* (5, 12, 13) {real, imag} */,
  {32'hbf0ca32c, 32'h00000000} /* (5, 12, 12) {real, imag} */,
  {32'hbec08222, 32'h00000000} /* (5, 12, 11) {real, imag} */,
  {32'hbf0081eb, 32'h00000000} /* (5, 12, 10) {real, imag} */,
  {32'hbf4aecd9, 32'h00000000} /* (5, 12, 9) {real, imag} */,
  {32'hbea53a6a, 32'h00000000} /* (5, 12, 8) {real, imag} */,
  {32'hbbf1989b, 32'h00000000} /* (5, 12, 7) {real, imag} */,
  {32'hbea489d5, 32'h00000000} /* (5, 12, 6) {real, imag} */,
  {32'hbe9ff6eb, 32'h00000000} /* (5, 12, 5) {real, imag} */,
  {32'hbeb6a605, 32'h00000000} /* (5, 12, 4) {real, imag} */,
  {32'hbdaa646b, 32'h00000000} /* (5, 12, 3) {real, imag} */,
  {32'hbe166cd7, 32'h00000000} /* (5, 12, 2) {real, imag} */,
  {32'hbee4c621, 32'h00000000} /* (5, 12, 1) {real, imag} */,
  {32'hbed850e6, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h3e4686f6, 32'h00000000} /* (5, 11, 15) {real, imag} */,
  {32'hbe6ed078, 32'h00000000} /* (5, 11, 14) {real, imag} */,
  {32'hbf41fba4, 32'h00000000} /* (5, 11, 13) {real, imag} */,
  {32'hbe5370f1, 32'h00000000} /* (5, 11, 12) {real, imag} */,
  {32'hbd834ef0, 32'h00000000} /* (5, 11, 11) {real, imag} */,
  {32'hbf2fcb34, 32'h00000000} /* (5, 11, 10) {real, imag} */,
  {32'hbf4fa054, 32'h00000000} /* (5, 11, 9) {real, imag} */,
  {32'hbf2bdf78, 32'h00000000} /* (5, 11, 8) {real, imag} */,
  {32'hbe0dc2ce, 32'h00000000} /* (5, 11, 7) {real, imag} */,
  {32'h3e948e9a, 32'h00000000} /* (5, 11, 6) {real, imag} */,
  {32'h3e0dc3d3, 32'h00000000} /* (5, 11, 5) {real, imag} */,
  {32'hbdc85bad, 32'h00000000} /* (5, 11, 4) {real, imag} */,
  {32'h3da4a8f2, 32'h00000000} /* (5, 11, 3) {real, imag} */,
  {32'hbdf40346, 32'h00000000} /* (5, 11, 2) {real, imag} */,
  {32'hbe266c64, 32'h00000000} /* (5, 11, 1) {real, imag} */,
  {32'hbe3c0c5d, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'hbd52e4e8, 32'h00000000} /* (5, 10, 15) {real, imag} */,
  {32'hbef72502, 32'h00000000} /* (5, 10, 14) {real, imag} */,
  {32'hbf1d30b2, 32'h00000000} /* (5, 10, 13) {real, imag} */,
  {32'hbeaa4529, 32'h00000000} /* (5, 10, 12) {real, imag} */,
  {32'hbcc602b8, 32'h00000000} /* (5, 10, 11) {real, imag} */,
  {32'hbe00dae8, 32'h00000000} /* (5, 10, 10) {real, imag} */,
  {32'hbe4d4d05, 32'h00000000} /* (5, 10, 9) {real, imag} */,
  {32'hbe9ae406, 32'h00000000} /* (5, 10, 8) {real, imag} */,
  {32'hbe791286, 32'h00000000} /* (5, 10, 7) {real, imag} */,
  {32'h3e190422, 32'h00000000} /* (5, 10, 6) {real, imag} */,
  {32'h3ea4a0d8, 32'h00000000} /* (5, 10, 5) {real, imag} */,
  {32'h3ea3cb4a, 32'h00000000} /* (5, 10, 4) {real, imag} */,
  {32'h3e1d4c54, 32'h00000000} /* (5, 10, 3) {real, imag} */,
  {32'h3de20c9a, 32'h00000000} /* (5, 10, 2) {real, imag} */,
  {32'h3e43537a, 32'h00000000} /* (5, 10, 1) {real, imag} */,
  {32'hbc30f2e0, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'h3e023bee, 32'h00000000} /* (5, 9, 15) {real, imag} */,
  {32'h3d542b3b, 32'h00000000} /* (5, 9, 14) {real, imag} */,
  {32'h3e0b74af, 32'h00000000} /* (5, 9, 13) {real, imag} */,
  {32'hbf0ee813, 32'h00000000} /* (5, 9, 12) {real, imag} */,
  {32'hbba24990, 32'h00000000} /* (5, 9, 11) {real, imag} */,
  {32'h3efd3b36, 32'h00000000} /* (5, 9, 10) {real, imag} */,
  {32'h3e8e4ced, 32'h00000000} /* (5, 9, 9) {real, imag} */,
  {32'h3d6db1b2, 32'h00000000} /* (5, 9, 8) {real, imag} */,
  {32'h3e275093, 32'h00000000} /* (5, 9, 7) {real, imag} */,
  {32'hbedf03d7, 32'h00000000} /* (5, 9, 6) {real, imag} */,
  {32'hbd92b9dd, 32'h00000000} /* (5, 9, 5) {real, imag} */,
  {32'hbc3f79f5, 32'h00000000} /* (5, 9, 4) {real, imag} */,
  {32'hbe7aa07c, 32'h00000000} /* (5, 9, 3) {real, imag} */,
  {32'h3b2faee8, 32'h00000000} /* (5, 9, 2) {real, imag} */,
  {32'h3df28b55, 32'h00000000} /* (5, 9, 1) {real, imag} */,
  {32'hbd748e7e, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'h3f218784, 32'h00000000} /* (5, 8, 15) {real, imag} */,
  {32'h3e44c85a, 32'h00000000} /* (5, 8, 14) {real, imag} */,
  {32'hbefb9f4e, 32'h00000000} /* (5, 8, 13) {real, imag} */,
  {32'hbf598f8a, 32'h00000000} /* (5, 8, 12) {real, imag} */,
  {32'hbea29a80, 32'h00000000} /* (5, 8, 11) {real, imag} */,
  {32'h3ec7f2d3, 32'h00000000} /* (5, 8, 10) {real, imag} */,
  {32'h3e4a4796, 32'h00000000} /* (5, 8, 9) {real, imag} */,
  {32'hbbfe8f60, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h3ed1990c, 32'h00000000} /* (5, 8, 7) {real, imag} */,
  {32'hbd20131d, 32'h00000000} /* (5, 8, 6) {real, imag} */,
  {32'h3e80facd, 32'h00000000} /* (5, 8, 5) {real, imag} */,
  {32'h3e68773a, 32'h00000000} /* (5, 8, 4) {real, imag} */,
  {32'hbe38baac, 32'h00000000} /* (5, 8, 3) {real, imag} */,
  {32'h3c9c0a3a, 32'h00000000} /* (5, 8, 2) {real, imag} */,
  {32'h3e84e7c2, 32'h00000000} /* (5, 8, 1) {real, imag} */,
  {32'h3ea3416a, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h3ebd1c1c, 32'h00000000} /* (5, 7, 15) {real, imag} */,
  {32'h3e89e663, 32'h00000000} /* (5, 7, 14) {real, imag} */,
  {32'hbeeb6e9e, 32'h00000000} /* (5, 7, 13) {real, imag} */,
  {32'hbf7767d0, 32'h00000000} /* (5, 7, 12) {real, imag} */,
  {32'hbf77f09c, 32'h00000000} /* (5, 7, 11) {real, imag} */,
  {32'h3dabe1ae, 32'h00000000} /* (5, 7, 10) {real, imag} */,
  {32'h3e24e550, 32'h00000000} /* (5, 7, 9) {real, imag} */,
  {32'h3d46e272, 32'h00000000} /* (5, 7, 8) {real, imag} */,
  {32'h3dd3c8d4, 32'h00000000} /* (5, 7, 7) {real, imag} */,
  {32'h3e7d2943, 32'h00000000} /* (5, 7, 6) {real, imag} */,
  {32'h3ed8b958, 32'h00000000} /* (5, 7, 5) {real, imag} */,
  {32'h3d83b829, 32'h00000000} /* (5, 7, 4) {real, imag} */,
  {32'hbcd77846, 32'h00000000} /* (5, 7, 3) {real, imag} */,
  {32'hbd59d1b2, 32'h00000000} /* (5, 7, 2) {real, imag} */,
  {32'h3eba673c, 32'h00000000} /* (5, 7, 1) {real, imag} */,
  {32'h3e10530c, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'h3e23e1ce, 32'h00000000} /* (5, 6, 15) {real, imag} */,
  {32'h3e89cdd7, 32'h00000000} /* (5, 6, 14) {real, imag} */,
  {32'hbeba2b78, 32'h00000000} /* (5, 6, 13) {real, imag} */,
  {32'hbf2d9d28, 32'h00000000} /* (5, 6, 12) {real, imag} */,
  {32'hbed1672f, 32'h00000000} /* (5, 6, 11) {real, imag} */,
  {32'h3d90c88d, 32'h00000000} /* (5, 6, 10) {real, imag} */,
  {32'hbe2fa51a, 32'h00000000} /* (5, 6, 9) {real, imag} */,
  {32'hbd524e6b, 32'h00000000} /* (5, 6, 8) {real, imag} */,
  {32'hbcb9ef29, 32'h00000000} /* (5, 6, 7) {real, imag} */,
  {32'h3d66e0e4, 32'h00000000} /* (5, 6, 6) {real, imag} */,
  {32'h3e4deff0, 32'h00000000} /* (5, 6, 5) {real, imag} */,
  {32'hbdf4f921, 32'h00000000} /* (5, 6, 4) {real, imag} */,
  {32'hbed77782, 32'h00000000} /* (5, 6, 3) {real, imag} */,
  {32'hbf53992a, 32'h00000000} /* (5, 6, 2) {real, imag} */,
  {32'hbee81844, 32'h00000000} /* (5, 6, 1) {real, imag} */,
  {32'h3d6acd4a, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'hbd881c6b, 32'h00000000} /* (5, 5, 15) {real, imag} */,
  {32'h3e841221, 32'h00000000} /* (5, 5, 14) {real, imag} */,
  {32'hbe122281, 32'h00000000} /* (5, 5, 13) {real, imag} */,
  {32'hbe823c83, 32'h00000000} /* (5, 5, 12) {real, imag} */,
  {32'hbdbee9e6, 32'h00000000} /* (5, 5, 11) {real, imag} */,
  {32'hbde5aff6, 32'h00000000} /* (5, 5, 10) {real, imag} */,
  {32'hbe047171, 32'h00000000} /* (5, 5, 9) {real, imag} */,
  {32'h3c8e7b52, 32'h00000000} /* (5, 5, 8) {real, imag} */,
  {32'h3db8dce5, 32'h00000000} /* (5, 5, 7) {real, imag} */,
  {32'h3e661314, 32'h00000000} /* (5, 5, 6) {real, imag} */,
  {32'h3dae41a7, 32'h00000000} /* (5, 5, 5) {real, imag} */,
  {32'hbe20674e, 32'h00000000} /* (5, 5, 4) {real, imag} */,
  {32'hbeaf1a9b, 32'h00000000} /* (5, 5, 3) {real, imag} */,
  {32'hbf0ae6f3, 32'h00000000} /* (5, 5, 2) {real, imag} */,
  {32'hbf50b586, 32'h00000000} /* (5, 5, 1) {real, imag} */,
  {32'hbdc91c3f, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'h3ec29207, 32'h00000000} /* (5, 4, 15) {real, imag} */,
  {32'h3f07457d, 32'h00000000} /* (5, 4, 14) {real, imag} */,
  {32'hbe23f29d, 32'h00000000} /* (5, 4, 13) {real, imag} */,
  {32'hbe8b42c8, 32'h00000000} /* (5, 4, 12) {real, imag} */,
  {32'h3d2dde2d, 32'h00000000} /* (5, 4, 11) {real, imag} */,
  {32'h3eaf91e3, 32'h00000000} /* (5, 4, 10) {real, imag} */,
  {32'h3eaf46b0, 32'h00000000} /* (5, 4, 9) {real, imag} */,
  {32'hbe64b809, 32'h00000000} /* (5, 4, 8) {real, imag} */,
  {32'hbe8164ca, 32'h00000000} /* (5, 4, 7) {real, imag} */,
  {32'h3e42ff3c, 32'h00000000} /* (5, 4, 6) {real, imag} */,
  {32'h3f239386, 32'h00000000} /* (5, 4, 5) {real, imag} */,
  {32'hbe13266a, 32'h00000000} /* (5, 4, 4) {real, imag} */,
  {32'hbf38d10b, 32'h00000000} /* (5, 4, 3) {real, imag} */,
  {32'hbe80bef6, 32'h00000000} /* (5, 4, 2) {real, imag} */,
  {32'hbe1fddc6, 32'h00000000} /* (5, 4, 1) {real, imag} */,
  {32'hbd674b53, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'h3be0e05d, 32'h00000000} /* (5, 3, 15) {real, imag} */,
  {32'h3ebf9aaf, 32'h00000000} /* (5, 3, 14) {real, imag} */,
  {32'h3e9b2ec8, 32'h00000000} /* (5, 3, 13) {real, imag} */,
  {32'hbda05133, 32'h00000000} /* (5, 3, 12) {real, imag} */,
  {32'h3f215ef7, 32'h00000000} /* (5, 3, 11) {real, imag} */,
  {32'h3e8aa23a, 32'h00000000} /* (5, 3, 10) {real, imag} */,
  {32'hbcd33775, 32'h00000000} /* (5, 3, 9) {real, imag} */,
  {32'hbeb02507, 32'h00000000} /* (5, 3, 8) {real, imag} */,
  {32'hbe5771d3, 32'h00000000} /* (5, 3, 7) {real, imag} */,
  {32'hbe3c4d4d, 32'h00000000} /* (5, 3, 6) {real, imag} */,
  {32'h3c4c49c0, 32'h00000000} /* (5, 3, 5) {real, imag} */,
  {32'hbf743025, 32'h00000000} /* (5, 3, 4) {real, imag} */,
  {32'hbf1cb042, 32'h00000000} /* (5, 3, 3) {real, imag} */,
  {32'hbe4d5479, 32'h00000000} /* (5, 3, 2) {real, imag} */,
  {32'h3e120961, 32'h00000000} /* (5, 3, 1) {real, imag} */,
  {32'h3e23657f, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'hbf13d011, 32'h00000000} /* (5, 2, 15) {real, imag} */,
  {32'hbea89bb4, 32'h00000000} /* (5, 2, 14) {real, imag} */,
  {32'h3e9e99f2, 32'h00000000} /* (5, 2, 13) {real, imag} */,
  {32'hbcfdab30, 32'h00000000} /* (5, 2, 12) {real, imag} */,
  {32'h3d2ff7c0, 32'h00000000} /* (5, 2, 11) {real, imag} */,
  {32'hbf381c70, 32'h00000000} /* (5, 2, 10) {real, imag} */,
  {32'hbd85b158, 32'h00000000} /* (5, 2, 9) {real, imag} */,
  {32'h3e066280, 32'h00000000} /* (5, 2, 8) {real, imag} */,
  {32'h3e0e7cf7, 32'h00000000} /* (5, 2, 7) {real, imag} */,
  {32'h3c9ce96a, 32'h00000000} /* (5, 2, 6) {real, imag} */,
  {32'h3ec392a0, 32'h00000000} /* (5, 2, 5) {real, imag} */,
  {32'h3e83bebb, 32'h00000000} /* (5, 2, 4) {real, imag} */,
  {32'h3da91bf7, 32'h00000000} /* (5, 2, 3) {real, imag} */,
  {32'hbe430287, 32'h00000000} /* (5, 2, 2) {real, imag} */,
  {32'hbe5513bb, 32'h00000000} /* (5, 2, 1) {real, imag} */,
  {32'hbe74e4eb, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'hbedbe507, 32'h00000000} /* (5, 1, 15) {real, imag} */,
  {32'h3ddfebf0, 32'h00000000} /* (5, 1, 14) {real, imag} */,
  {32'h3ef7c29d, 32'h00000000} /* (5, 1, 13) {real, imag} */,
  {32'h3dcc56d6, 32'h00000000} /* (5, 1, 12) {real, imag} */,
  {32'hbe597511, 32'h00000000} /* (5, 1, 11) {real, imag} */,
  {32'h3e1894ad, 32'h00000000} /* (5, 1, 10) {real, imag} */,
  {32'h3eedbec1, 32'h00000000} /* (5, 1, 9) {real, imag} */,
  {32'h3df226fd, 32'h00000000} /* (5, 1, 8) {real, imag} */,
  {32'hbece131d, 32'h00000000} /* (5, 1, 7) {real, imag} */,
  {32'hbdb6d31b, 32'h00000000} /* (5, 1, 6) {real, imag} */,
  {32'h3ed6ee54, 32'h00000000} /* (5, 1, 5) {real, imag} */,
  {32'h3e8a86ab, 32'h00000000} /* (5, 1, 4) {real, imag} */,
  {32'hbe8e45e6, 32'h00000000} /* (5, 1, 3) {real, imag} */,
  {32'hbeb6e608, 32'h00000000} /* (5, 1, 2) {real, imag} */,
  {32'hbe87b0d4, 32'h00000000} /* (5, 1, 1) {real, imag} */,
  {32'hbebe06b3, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'hbe23ebf9, 32'h00000000} /* (5, 0, 15) {real, imag} */,
  {32'h3d851943, 32'h00000000} /* (5, 0, 14) {real, imag} */,
  {32'h3d72f67e, 32'h00000000} /* (5, 0, 13) {real, imag} */,
  {32'hbe9e908f, 32'h00000000} /* (5, 0, 12) {real, imag} */,
  {32'hbe9abb9f, 32'h00000000} /* (5, 0, 11) {real, imag} */,
  {32'hbe0dbb9a, 32'h00000000} /* (5, 0, 10) {real, imag} */,
  {32'h3bd2685a, 32'h00000000} /* (5, 0, 9) {real, imag} */,
  {32'h3eb1d732, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'hbd8ee4a6, 32'h00000000} /* (5, 0, 7) {real, imag} */,
  {32'hbd51aad3, 32'h00000000} /* (5, 0, 6) {real, imag} */,
  {32'h3e82ac7a, 32'h00000000} /* (5, 0, 5) {real, imag} */,
  {32'h3daa4954, 32'h00000000} /* (5, 0, 4) {real, imag} */,
  {32'h3d43af41, 32'h00000000} /* (5, 0, 3) {real, imag} */,
  {32'hbda405d9, 32'h00000000} /* (5, 0, 2) {real, imag} */,
  {32'hbe14d165, 32'h00000000} /* (5, 0, 1) {real, imag} */,
  {32'hbd26bb94, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hbe4e4819, 32'h00000000} /* (4, 15, 15) {real, imag} */,
  {32'hbe4d3f2b, 32'h00000000} /* (4, 15, 14) {real, imag} */,
  {32'h3e8ca39c, 32'h00000000} /* (4, 15, 13) {real, imag} */,
  {32'h3e745c7d, 32'h00000000} /* (4, 15, 12) {real, imag} */,
  {32'h3dc85f50, 32'h00000000} /* (4, 15, 11) {real, imag} */,
  {32'hbc6f5fe1, 32'h00000000} /* (4, 15, 10) {real, imag} */,
  {32'hbe099b04, 32'h00000000} /* (4, 15, 9) {real, imag} */,
  {32'hbdf24597, 32'h00000000} /* (4, 15, 8) {real, imag} */,
  {32'hbe02dbdd, 32'h00000000} /* (4, 15, 7) {real, imag} */,
  {32'h3e2de8b1, 32'h00000000} /* (4, 15, 6) {real, imag} */,
  {32'h3ece93c0, 32'h00000000} /* (4, 15, 5) {real, imag} */,
  {32'h3e86db7a, 32'h00000000} /* (4, 15, 4) {real, imag} */,
  {32'h3e1207dc, 32'h00000000} /* (4, 15, 3) {real, imag} */,
  {32'hbd8a9c12, 32'h00000000} /* (4, 15, 2) {real, imag} */,
  {32'h3c1b88a1, 32'h00000000} /* (4, 15, 1) {real, imag} */,
  {32'h3dbc25bc, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'hbe78d636, 32'h00000000} /* (4, 14, 15) {real, imag} */,
  {32'hbf3207b6, 32'h00000000} /* (4, 14, 14) {real, imag} */,
  {32'hbea2a575, 32'h00000000} /* (4, 14, 13) {real, imag} */,
  {32'h3d1381be, 32'h00000000} /* (4, 14, 12) {real, imag} */,
  {32'h3da03a9d, 32'h00000000} /* (4, 14, 11) {real, imag} */,
  {32'hbf142fbe, 32'h00000000} /* (4, 14, 10) {real, imag} */,
  {32'hbf52e26f, 32'h00000000} /* (4, 14, 9) {real, imag} */,
  {32'hbea2ae66, 32'h00000000} /* (4, 14, 8) {real, imag} */,
  {32'hbc841626, 32'h00000000} /* (4, 14, 7) {real, imag} */,
  {32'h3e18689f, 32'h00000000} /* (4, 14, 6) {real, imag} */,
  {32'h3db3c507, 32'h00000000} /* (4, 14, 5) {real, imag} */,
  {32'h3e28dde4, 32'h00000000} /* (4, 14, 4) {real, imag} */,
  {32'h3de10f24, 32'h00000000} /* (4, 14, 3) {real, imag} */,
  {32'hbe0dc7ec, 32'h00000000} /* (4, 14, 2) {real, imag} */,
  {32'h3ebae93d, 32'h00000000} /* (4, 14, 1) {real, imag} */,
  {32'h3f0e195b, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'hbe407002, 32'h00000000} /* (4, 13, 15) {real, imag} */,
  {32'hbf23e308, 32'h00000000} /* (4, 13, 14) {real, imag} */,
  {32'hbe6af644, 32'h00000000} /* (4, 13, 13) {real, imag} */,
  {32'h3ea3fe52, 32'h00000000} /* (4, 13, 12) {real, imag} */,
  {32'hbe9dfdae, 32'h00000000} /* (4, 13, 11) {real, imag} */,
  {32'hbf02feed, 32'h00000000} /* (4, 13, 10) {real, imag} */,
  {32'hbf2723fa, 32'h00000000} /* (4, 13, 9) {real, imag} */,
  {32'h3dec0760, 32'h00000000} /* (4, 13, 8) {real, imag} */,
  {32'h3ee96f57, 32'h00000000} /* (4, 13, 7) {real, imag} */,
  {32'h3ea1e938, 32'h00000000} /* (4, 13, 6) {real, imag} */,
  {32'h3dd3beee, 32'h00000000} /* (4, 13, 5) {real, imag} */,
  {32'h3d2722fe, 32'h00000000} /* (4, 13, 4) {real, imag} */,
  {32'h3ef449eb, 32'h00000000} /* (4, 13, 3) {real, imag} */,
  {32'hbc642ac7, 32'h00000000} /* (4, 13, 2) {real, imag} */,
  {32'hbc04aad2, 32'h00000000} /* (4, 13, 1) {real, imag} */,
  {32'h3e18c06a, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'hbec08784, 32'h00000000} /* (4, 12, 15) {real, imag} */,
  {32'hbe3106f2, 32'h00000000} /* (4, 12, 14) {real, imag} */,
  {32'h3f19ad09, 32'h00000000} /* (4, 12, 13) {real, imag} */,
  {32'h3e96c49e, 32'h00000000} /* (4, 12, 12) {real, imag} */,
  {32'hbeea23ae, 32'h00000000} /* (4, 12, 11) {real, imag} */,
  {32'hbeb59d9d, 32'h00000000} /* (4, 12, 10) {real, imag} */,
  {32'hbe6faedf, 32'h00000000} /* (4, 12, 9) {real, imag} */,
  {32'hbdb7a37b, 32'h00000000} /* (4, 12, 8) {real, imag} */,
  {32'hbc8b753a, 32'h00000000} /* (4, 12, 7) {real, imag} */,
  {32'h3eb52345, 32'h00000000} /* (4, 12, 6) {real, imag} */,
  {32'h3f507931, 32'h00000000} /* (4, 12, 5) {real, imag} */,
  {32'hbe19f6de, 32'h00000000} /* (4, 12, 4) {real, imag} */,
  {32'hbe145edc, 32'h00000000} /* (4, 12, 3) {real, imag} */,
  {32'hbe2251dc, 32'h00000000} /* (4, 12, 2) {real, imag} */,
  {32'h3df52040, 32'h00000000} /* (4, 12, 1) {real, imag} */,
  {32'hbd9b2458, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'hbe61f723, 32'h00000000} /* (4, 11, 15) {real, imag} */,
  {32'hbe99795b, 32'h00000000} /* (4, 11, 14) {real, imag} */,
  {32'h3e39d0d8, 32'h00000000} /* (4, 11, 13) {real, imag} */,
  {32'h3c1b172f, 32'h00000000} /* (4, 11, 12) {real, imag} */,
  {32'hbed6a431, 32'h00000000} /* (4, 11, 11) {real, imag} */,
  {32'hbebcaaa2, 32'h00000000} /* (4, 11, 10) {real, imag} */,
  {32'hbe852f76, 32'h00000000} /* (4, 11, 9) {real, imag} */,
  {32'hbea7d978, 32'h00000000} /* (4, 11, 8) {real, imag} */,
  {32'h3e9619d1, 32'h00000000} /* (4, 11, 7) {real, imag} */,
  {32'h3f3d35fe, 32'h00000000} /* (4, 11, 6) {real, imag} */,
  {32'h3f840682, 32'h00000000} /* (4, 11, 5) {real, imag} */,
  {32'h3e8d4ca7, 32'h00000000} /* (4, 11, 4) {real, imag} */,
  {32'hbd8d1e0f, 32'h00000000} /* (4, 11, 3) {real, imag} */,
  {32'hbda215c0, 32'h00000000} /* (4, 11, 2) {real, imag} */,
  {32'hbbe7c5b5, 32'h00000000} /* (4, 11, 1) {real, imag} */,
  {32'h3dd88f1d, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hbe183ad7, 32'h00000000} /* (4, 10, 15) {real, imag} */,
  {32'hbeb271d9, 32'h00000000} /* (4, 10, 14) {real, imag} */,
  {32'h3e0ed26b, 32'h00000000} /* (4, 10, 13) {real, imag} */,
  {32'h3e125556, 32'h00000000} /* (4, 10, 12) {real, imag} */,
  {32'hbdd5eb1e, 32'h00000000} /* (4, 10, 11) {real, imag} */,
  {32'h3cd31e47, 32'h00000000} /* (4, 10, 10) {real, imag} */,
  {32'hbe9c6b57, 32'h00000000} /* (4, 10, 9) {real, imag} */,
  {32'hbd9e0c46, 32'h00000000} /* (4, 10, 8) {real, imag} */,
  {32'h3d85ccc4, 32'h00000000} /* (4, 10, 7) {real, imag} */,
  {32'hbb83e1b7, 32'h00000000} /* (4, 10, 6) {real, imag} */,
  {32'h3eb2999a, 32'h00000000} /* (4, 10, 5) {real, imag} */,
  {32'h3e7be574, 32'h00000000} /* (4, 10, 4) {real, imag} */,
  {32'hbe2d1578, 32'h00000000} /* (4, 10, 3) {real, imag} */,
  {32'hbeb3c667, 32'h00000000} /* (4, 10, 2) {real, imag} */,
  {32'hbe06b8fc, 32'h00000000} /* (4, 10, 1) {real, imag} */,
  {32'h3e2ac351, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'hbde7e398, 32'h00000000} /* (4, 9, 15) {real, imag} */,
  {32'hbe32729e, 32'h00000000} /* (4, 9, 14) {real, imag} */,
  {32'h3e34659b, 32'h00000000} /* (4, 9, 13) {real, imag} */,
  {32'hbec75922, 32'h00000000} /* (4, 9, 12) {real, imag} */,
  {32'hbee200ab, 32'h00000000} /* (4, 9, 11) {real, imag} */,
  {32'hbb18accf, 32'h00000000} /* (4, 9, 10) {real, imag} */,
  {32'hbe8ab82e, 32'h00000000} /* (4, 9, 9) {real, imag} */,
  {32'hbcce5447, 32'h00000000} /* (4, 9, 8) {real, imag} */,
  {32'h3e6b92d7, 32'h00000000} /* (4, 9, 7) {real, imag} */,
  {32'hbee06c52, 32'h00000000} /* (4, 9, 6) {real, imag} */,
  {32'hbe89865a, 32'h00000000} /* (4, 9, 5) {real, imag} */,
  {32'hbecc539a, 32'h00000000} /* (4, 9, 4) {real, imag} */,
  {32'hbed3229f, 32'h00000000} /* (4, 9, 3) {real, imag} */,
  {32'hbeaeb5f0, 32'h00000000} /* (4, 9, 2) {real, imag} */,
  {32'h3de00bd6, 32'h00000000} /* (4, 9, 1) {real, imag} */,
  {32'h3e8171db, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'h3f1835e2, 32'h00000000} /* (4, 8, 15) {real, imag} */,
  {32'h3e79f84f, 32'h00000000} /* (4, 8, 14) {real, imag} */,
  {32'hbe1536e6, 32'h00000000} /* (4, 8, 13) {real, imag} */,
  {32'hbefbde37, 32'h00000000} /* (4, 8, 12) {real, imag} */,
  {32'hbede4942, 32'h00000000} /* (4, 8, 11) {real, imag} */,
  {32'hbbccc573, 32'h00000000} /* (4, 8, 10) {real, imag} */,
  {32'hbd62497c, 32'h00000000} /* (4, 8, 9) {real, imag} */,
  {32'hbf0862b6, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'hbb4a40e0, 32'h00000000} /* (4, 8, 7) {real, imag} */,
  {32'h3e93dbb1, 32'h00000000} /* (4, 8, 6) {real, imag} */,
  {32'h3eaeb807, 32'h00000000} /* (4, 8, 5) {real, imag} */,
  {32'hbe88a51a, 32'h00000000} /* (4, 8, 4) {real, imag} */,
  {32'hbf26a27c, 32'h00000000} /* (4, 8, 3) {real, imag} */,
  {32'hbec73186, 32'h00000000} /* (4, 8, 2) {real, imag} */,
  {32'h3e6b3665, 32'h00000000} /* (4, 8, 1) {real, imag} */,
  {32'h3ee3ec9b, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'h3ea041d1, 32'h00000000} /* (4, 7, 15) {real, imag} */,
  {32'h3e9ba329, 32'h00000000} /* (4, 7, 14) {real, imag} */,
  {32'hbe03a97d, 32'h00000000} /* (4, 7, 13) {real, imag} */,
  {32'hbeda651d, 32'h00000000} /* (4, 7, 12) {real, imag} */,
  {32'hbf244591, 32'h00000000} /* (4, 7, 11) {real, imag} */,
  {32'hbdbd16ba, 32'h00000000} /* (4, 7, 10) {real, imag} */,
  {32'h3f25983b, 32'h00000000} /* (4, 7, 9) {real, imag} */,
  {32'hbd3cf03a, 32'h00000000} /* (4, 7, 8) {real, imag} */,
  {32'hbdba8524, 32'h00000000} /* (4, 7, 7) {real, imag} */,
  {32'h3d098ce4, 32'h00000000} /* (4, 7, 6) {real, imag} */,
  {32'h3db80a4e, 32'h00000000} /* (4, 7, 5) {real, imag} */,
  {32'hbea08007, 32'h00000000} /* (4, 7, 4) {real, imag} */,
  {32'hbe83c7dc, 32'h00000000} /* (4, 7, 3) {real, imag} */,
  {32'hbe43504e, 32'h00000000} /* (4, 7, 2) {real, imag} */,
  {32'hbe8665fa, 32'h00000000} /* (4, 7, 1) {real, imag} */,
  {32'hbd506bd6, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'h3d534f5a, 32'h00000000} /* (4, 6, 15) {real, imag} */,
  {32'hbe81bc9c, 32'h00000000} /* (4, 6, 14) {real, imag} */,
  {32'hbf29a84d, 32'h00000000} /* (4, 6, 13) {real, imag} */,
  {32'hbf40057e, 32'h00000000} /* (4, 6, 12) {real, imag} */,
  {32'hbf217bed, 32'h00000000} /* (4, 6, 11) {real, imag} */,
  {32'hbe981cfd, 32'h00000000} /* (4, 6, 10) {real, imag} */,
  {32'h3e927b88, 32'h00000000} /* (4, 6, 9) {real, imag} */,
  {32'h3da3d721, 32'h00000000} /* (4, 6, 8) {real, imag} */,
  {32'h3dc16a74, 32'h00000000} /* (4, 6, 7) {real, imag} */,
  {32'h3ec3149e, 32'h00000000} /* (4, 6, 6) {real, imag} */,
  {32'hbda7769e, 32'h00000000} /* (4, 6, 5) {real, imag} */,
  {32'hbdf6dabf, 32'h00000000} /* (4, 6, 4) {real, imag} */,
  {32'hbe14c1cc, 32'h00000000} /* (4, 6, 3) {real, imag} */,
  {32'hbf1fd533, 32'h00000000} /* (4, 6, 2) {real, imag} */,
  {32'hbf0ae657, 32'h00000000} /* (4, 6, 1) {real, imag} */,
  {32'hbe76de03, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'hbdfe0455, 32'h00000000} /* (4, 5, 15) {real, imag} */,
  {32'hbe743823, 32'h00000000} /* (4, 5, 14) {real, imag} */,
  {32'hbed7b076, 32'h00000000} /* (4, 5, 13) {real, imag} */,
  {32'hbd986ffd, 32'h00000000} /* (4, 5, 12) {real, imag} */,
  {32'h3b449fe3, 32'h00000000} /* (4, 5, 11) {real, imag} */,
  {32'h3bff3e2a, 32'h00000000} /* (4, 5, 10) {real, imag} */,
  {32'h3e4c1e0b, 32'h00000000} /* (4, 5, 9) {real, imag} */,
  {32'h3e7c6515, 32'h00000000} /* (4, 5, 8) {real, imag} */,
  {32'h3eb262e3, 32'h00000000} /* (4, 5, 7) {real, imag} */,
  {32'h3f628076, 32'h00000000} /* (4, 5, 6) {real, imag} */,
  {32'h3e931b5a, 32'h00000000} /* (4, 5, 5) {real, imag} */,
  {32'h3e2838e8, 32'h00000000} /* (4, 5, 4) {real, imag} */,
  {32'h3e4a7efb, 32'h00000000} /* (4, 5, 3) {real, imag} */,
  {32'hbe482215, 32'h00000000} /* (4, 5, 2) {real, imag} */,
  {32'hbd082558, 32'h00000000} /* (4, 5, 1) {real, imag} */,
  {32'hbd665218, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hbe031325, 32'h00000000} /* (4, 4, 15) {real, imag} */,
  {32'hbe7c5c01, 32'h00000000} /* (4, 4, 14) {real, imag} */,
  {32'hbea5d1bb, 32'h00000000} /* (4, 4, 13) {real, imag} */,
  {32'h3e841cb9, 32'h00000000} /* (4, 4, 12) {real, imag} */,
  {32'h3f092ab3, 32'h00000000} /* (4, 4, 11) {real, imag} */,
  {32'h3eda16fa, 32'h00000000} /* (4, 4, 10) {real, imag} */,
  {32'h3e983394, 32'h00000000} /* (4, 4, 9) {real, imag} */,
  {32'hbe7f21cf, 32'h00000000} /* (4, 4, 8) {real, imag} */,
  {32'hbf04b97d, 32'h00000000} /* (4, 4, 7) {real, imag} */,
  {32'h3d1af311, 32'h00000000} /* (4, 4, 6) {real, imag} */,
  {32'h3eaf6018, 32'h00000000} /* (4, 4, 5) {real, imag} */,
  {32'hbdde1916, 32'h00000000} /* (4, 4, 4) {real, imag} */,
  {32'hbe862e70, 32'h00000000} /* (4, 4, 3) {real, imag} */,
  {32'hbe6c9a00, 32'h00000000} /* (4, 4, 2) {real, imag} */,
  {32'hbe1830e3, 32'h00000000} /* (4, 4, 1) {real, imag} */,
  {32'h3e00d24b, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hbe532b15, 32'h00000000} /* (4, 3, 15) {real, imag} */,
  {32'hbeb363dd, 32'h00000000} /* (4, 3, 14) {real, imag} */,
  {32'hbea05c25, 32'h00000000} /* (4, 3, 13) {real, imag} */,
  {32'h3ec6ecc4, 32'h00000000} /* (4, 3, 12) {real, imag} */,
  {32'h3f079c91, 32'h00000000} /* (4, 3, 11) {real, imag} */,
  {32'hbb90543e, 32'h00000000} /* (4, 3, 10) {real, imag} */,
  {32'h3e7b66af, 32'h00000000} /* (4, 3, 9) {real, imag} */,
  {32'hbe1efed6, 32'h00000000} /* (4, 3, 8) {real, imag} */,
  {32'hbdb6084e, 32'h00000000} /* (4, 3, 7) {real, imag} */,
  {32'hbe504f02, 32'h00000000} /* (4, 3, 6) {real, imag} */,
  {32'hbe8cd295, 32'h00000000} /* (4, 3, 5) {real, imag} */,
  {32'hbf349462, 32'h00000000} /* (4, 3, 4) {real, imag} */,
  {32'hbf0c53ab, 32'h00000000} /* (4, 3, 3) {real, imag} */,
  {32'hbee466f5, 32'h00000000} /* (4, 3, 2) {real, imag} */,
  {32'hbecf061c, 32'h00000000} /* (4, 3, 1) {real, imag} */,
  {32'h3e5d8ece, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hbedf5c77, 32'h00000000} /* (4, 2, 15) {real, imag} */,
  {32'hbed33d04, 32'h00000000} /* (4, 2, 14) {real, imag} */,
  {32'h3e38871f, 32'h00000000} /* (4, 2, 13) {real, imag} */,
  {32'h3f1239bc, 32'h00000000} /* (4, 2, 12) {real, imag} */,
  {32'h3e264962, 32'h00000000} /* (4, 2, 11) {real, imag} */,
  {32'hbeb4223c, 32'h00000000} /* (4, 2, 10) {real, imag} */,
  {32'hbdd7f0ca, 32'h00000000} /* (4, 2, 9) {real, imag} */,
  {32'h3a9cfbcb, 32'h00000000} /* (4, 2, 8) {real, imag} */,
  {32'h3d1fdd9a, 32'h00000000} /* (4, 2, 7) {real, imag} */,
  {32'hbe21c943, 32'h00000000} /* (4, 2, 6) {real, imag} */,
  {32'hbe242882, 32'h00000000} /* (4, 2, 5) {real, imag} */,
  {32'hbf12970e, 32'h00000000} /* (4, 2, 4) {real, imag} */,
  {32'hbf135860, 32'h00000000} /* (4, 2, 3) {real, imag} */,
  {32'hbed42f52, 32'h00000000} /* (4, 2, 2) {real, imag} */,
  {32'hbe557d4b, 32'h00000000} /* (4, 2, 1) {real, imag} */,
  {32'h3d50b2e7, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hbe38279e, 32'h00000000} /* (4, 1, 15) {real, imag} */,
  {32'h3da84578, 32'h00000000} /* (4, 1, 14) {real, imag} */,
  {32'h3f0e0b87, 32'h00000000} /* (4, 1, 13) {real, imag} */,
  {32'h3e382153, 32'h00000000} /* (4, 1, 12) {real, imag} */,
  {32'hbe339db8, 32'h00000000} /* (4, 1, 11) {real, imag} */,
  {32'h3e041334, 32'h00000000} /* (4, 1, 10) {real, imag} */,
  {32'h3dbedbf6, 32'h00000000} /* (4, 1, 9) {real, imag} */,
  {32'h3e005fcd, 32'h00000000} /* (4, 1, 8) {real, imag} */,
  {32'hbe1484ac, 32'h00000000} /* (4, 1, 7) {real, imag} */,
  {32'h3c21c760, 32'h00000000} /* (4, 1, 6) {real, imag} */,
  {32'h3e9bbe20, 32'h00000000} /* (4, 1, 5) {real, imag} */,
  {32'hbe5e003e, 32'h00000000} /* (4, 1, 4) {real, imag} */,
  {32'hbe68236a, 32'h00000000} /* (4, 1, 3) {real, imag} */,
  {32'hbe7df46e, 32'h00000000} /* (4, 1, 2) {real, imag} */,
  {32'hbebb6e80, 32'h00000000} /* (4, 1, 1) {real, imag} */,
  {32'hbd9efbfa, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hbdcc3b62, 32'h00000000} /* (4, 0, 15) {real, imag} */,
  {32'h3e098eb1, 32'h00000000} /* (4, 0, 14) {real, imag} */,
  {32'h3e7e0ade, 32'h00000000} /* (4, 0, 13) {real, imag} */,
  {32'hbed84770, 32'h00000000} /* (4, 0, 12) {real, imag} */,
  {32'hbf0d7a32, 32'h00000000} /* (4, 0, 11) {real, imag} */,
  {32'hbd8a9cd9, 32'h00000000} /* (4, 0, 10) {real, imag} */,
  {32'h3d12c78d, 32'h00000000} /* (4, 0, 9) {real, imag} */,
  {32'h3e9f58f8, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'hbd89091c, 32'h00000000} /* (4, 0, 7) {real, imag} */,
  {32'h3e112d68, 32'h00000000} /* (4, 0, 6) {real, imag} */,
  {32'h3ee91ff3, 32'h00000000} /* (4, 0, 5) {real, imag} */,
  {32'h3e52bf1d, 32'h00000000} /* (4, 0, 4) {real, imag} */,
  {32'hb9e6eb7e, 32'h00000000} /* (4, 0, 3) {real, imag} */,
  {32'hbe5eebae, 32'h00000000} /* (4, 0, 2) {real, imag} */,
  {32'hbe59fcd3, 32'h00000000} /* (4, 0, 1) {real, imag} */,
  {32'hbc6775d9, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hbe14d9a9, 32'h00000000} /* (3, 15, 15) {real, imag} */,
  {32'hbe8b9b5a, 32'h00000000} /* (3, 15, 14) {real, imag} */,
  {32'h3d58c449, 32'h00000000} /* (3, 15, 13) {real, imag} */,
  {32'h3e23f14c, 32'h00000000} /* (3, 15, 12) {real, imag} */,
  {32'h3ebc7874, 32'h00000000} /* (3, 15, 11) {real, imag} */,
  {32'h3e3ec425, 32'h00000000} /* (3, 15, 10) {real, imag} */,
  {32'h3dad6584, 32'h00000000} /* (3, 15, 9) {real, imag} */,
  {32'h3e9f1a7b, 32'h00000000} /* (3, 15, 8) {real, imag} */,
  {32'h3e288830, 32'h00000000} /* (3, 15, 7) {real, imag} */,
  {32'h3ba04b49, 32'h00000000} /* (3, 15, 6) {real, imag} */,
  {32'h3e1a8560, 32'h00000000} /* (3, 15, 5) {real, imag} */,
  {32'hbe6f17e0, 32'h00000000} /* (3, 15, 4) {real, imag} */,
  {32'hbdcb5208, 32'h00000000} /* (3, 15, 3) {real, imag} */,
  {32'h3dee2d2b, 32'h00000000} /* (3, 15, 2) {real, imag} */,
  {32'hbdf304e0, 32'h00000000} /* (3, 15, 1) {real, imag} */,
  {32'hbe474cec, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'h3dd2368a, 32'h00000000} /* (3, 14, 15) {real, imag} */,
  {32'hbef1922a, 32'h00000000} /* (3, 14, 14) {real, imag} */,
  {32'hbed8f243, 32'h00000000} /* (3, 14, 13) {real, imag} */,
  {32'h3e9d2ffa, 32'h00000000} /* (3, 14, 12) {real, imag} */,
  {32'h3f1c0855, 32'h00000000} /* (3, 14, 11) {real, imag} */,
  {32'hbe22c747, 32'h00000000} /* (3, 14, 10) {real, imag} */,
  {32'hbeb45f43, 32'h00000000} /* (3, 14, 9) {real, imag} */,
  {32'h3f029d16, 32'h00000000} /* (3, 14, 8) {real, imag} */,
  {32'h3c23d03a, 32'h00000000} /* (3, 14, 7) {real, imag} */,
  {32'hbe7cab26, 32'h00000000} /* (3, 14, 6) {real, imag} */,
  {32'h3e55f71a, 32'h00000000} /* (3, 14, 5) {real, imag} */,
  {32'h3e0449b9, 32'h00000000} /* (3, 14, 4) {real, imag} */,
  {32'h3d2932a7, 32'h00000000} /* (3, 14, 3) {real, imag} */,
  {32'hbdcd548a, 32'h00000000} /* (3, 14, 2) {real, imag} */,
  {32'hbe666150, 32'h00000000} /* (3, 14, 1) {real, imag} */,
  {32'h3e5768b0, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h3d6d635a, 32'h00000000} /* (3, 13, 15) {real, imag} */,
  {32'hbf18eb73, 32'h00000000} /* (3, 13, 14) {real, imag} */,
  {32'hbdde4277, 32'h00000000} /* (3, 13, 13) {real, imag} */,
  {32'h3f33793d, 32'h00000000} /* (3, 13, 12) {real, imag} */,
  {32'h3e3f6c68, 32'h00000000} /* (3, 13, 11) {real, imag} */,
  {32'hbe9f1d49, 32'h00000000} /* (3, 13, 10) {real, imag} */,
  {32'hbec33567, 32'h00000000} /* (3, 13, 9) {real, imag} */,
  {32'h3ea43834, 32'h00000000} /* (3, 13, 8) {real, imag} */,
  {32'h3db42468, 32'h00000000} /* (3, 13, 7) {real, imag} */,
  {32'h3e184671, 32'h00000000} /* (3, 13, 6) {real, imag} */,
  {32'h3eb144c4, 32'h00000000} /* (3, 13, 5) {real, imag} */,
  {32'h3e387d64, 32'h00000000} /* (3, 13, 4) {real, imag} */,
  {32'h3edfcd48, 32'h00000000} /* (3, 13, 3) {real, imag} */,
  {32'h3d4a0125, 32'h00000000} /* (3, 13, 2) {real, imag} */,
  {32'h3e27e3ea, 32'h00000000} /* (3, 13, 1) {real, imag} */,
  {32'h3eb85002, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'hbdb1918b, 32'h00000000} /* (3, 12, 15) {real, imag} */,
  {32'hbe5155f3, 32'h00000000} /* (3, 12, 14) {real, imag} */,
  {32'h3f260ace, 32'h00000000} /* (3, 12, 13) {real, imag} */,
  {32'h3f2eb8cc, 32'h00000000} /* (3, 12, 12) {real, imag} */,
  {32'hbe12778e, 32'h00000000} /* (3, 12, 11) {real, imag} */,
  {32'hbe60e74b, 32'h00000000} /* (3, 12, 10) {real, imag} */,
  {32'hbe0065b4, 32'h00000000} /* (3, 12, 9) {real, imag} */,
  {32'h3cdf0a38, 32'h00000000} /* (3, 12, 8) {real, imag} */,
  {32'h3d049990, 32'h00000000} /* (3, 12, 7) {real, imag} */,
  {32'h3f01b2b5, 32'h00000000} /* (3, 12, 6) {real, imag} */,
  {32'h3f46acfc, 32'h00000000} /* (3, 12, 5) {real, imag} */,
  {32'hbdad42d4, 32'h00000000} /* (3, 12, 4) {real, imag} */,
  {32'hbe20748b, 32'h00000000} /* (3, 12, 3) {real, imag} */,
  {32'hbe19b2f6, 32'h00000000} /* (3, 12, 2) {real, imag} */,
  {32'hba7e1065, 32'h00000000} /* (3, 12, 1) {real, imag} */,
  {32'h3d04f7ae, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'hbe002cfe, 32'h00000000} /* (3, 11, 15) {real, imag} */,
  {32'hbea16b26, 32'h00000000} /* (3, 11, 14) {real, imag} */,
  {32'h3eb71342, 32'h00000000} /* (3, 11, 13) {real, imag} */,
  {32'h3e7afc63, 32'h00000000} /* (3, 11, 12) {real, imag} */,
  {32'h3e7d40ce, 32'h00000000} /* (3, 11, 11) {real, imag} */,
  {32'h3ad04ab1, 32'h00000000} /* (3, 11, 10) {real, imag} */,
  {32'h3e1b847f, 32'h00000000} /* (3, 11, 9) {real, imag} */,
  {32'h3e2121f2, 32'h00000000} /* (3, 11, 8) {real, imag} */,
  {32'hbea6800b, 32'h00000000} /* (3, 11, 7) {real, imag} */,
  {32'hbe16db9c, 32'h00000000} /* (3, 11, 6) {real, imag} */,
  {32'h3f0fd08e, 32'h00000000} /* (3, 11, 5) {real, imag} */,
  {32'h3f0a1763, 32'h00000000} /* (3, 11, 4) {real, imag} */,
  {32'h3e412d7e, 32'h00000000} /* (3, 11, 3) {real, imag} */,
  {32'hbd9d426b, 32'h00000000} /* (3, 11, 2) {real, imag} */,
  {32'hbe63e862, 32'h00000000} /* (3, 11, 1) {real, imag} */,
  {32'h3e0ef36e, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'h3cd8d23d, 32'h00000000} /* (3, 10, 15) {real, imag} */,
  {32'hbf2efa64, 32'h00000000} /* (3, 10, 14) {real, imag} */,
  {32'hbed12868, 32'h00000000} /* (3, 10, 13) {real, imag} */,
  {32'h3e55613d, 32'h00000000} /* (3, 10, 12) {real, imag} */,
  {32'h3ea21547, 32'h00000000} /* (3, 10, 11) {real, imag} */,
  {32'h3ea1c80e, 32'h00000000} /* (3, 10, 10) {real, imag} */,
  {32'hbc359d28, 32'h00000000} /* (3, 10, 9) {real, imag} */,
  {32'hbebb3ed0, 32'h00000000} /* (3, 10, 8) {real, imag} */,
  {32'hbeb0b35b, 32'h00000000} /* (3, 10, 7) {real, imag} */,
  {32'hbeea1cc7, 32'h00000000} /* (3, 10, 6) {real, imag} */,
  {32'hbdab59ac, 32'h00000000} /* (3, 10, 5) {real, imag} */,
  {32'h3ed8236b, 32'h00000000} /* (3, 10, 4) {real, imag} */,
  {32'hbd6bfd80, 32'h00000000} /* (3, 10, 3) {real, imag} */,
  {32'hbe8303bc, 32'h00000000} /* (3, 10, 2) {real, imag} */,
  {32'hbc859df5, 32'h00000000} /* (3, 10, 1) {real, imag} */,
  {32'h3e5dba03, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'h3e288b3e, 32'h00000000} /* (3, 9, 15) {real, imag} */,
  {32'h3c5dc2c1, 32'h00000000} /* (3, 9, 14) {real, imag} */,
  {32'hbe290330, 32'h00000000} /* (3, 9, 13) {real, imag} */,
  {32'hbe53aa56, 32'h00000000} /* (3, 9, 12) {real, imag} */,
  {32'hbe871271, 32'h00000000} /* (3, 9, 11) {real, imag} */,
  {32'hbd5f6e03, 32'h00000000} /* (3, 9, 10) {real, imag} */,
  {32'hbd58454b, 32'h00000000} /* (3, 9, 9) {real, imag} */,
  {32'hbe1c5d52, 32'h00000000} /* (3, 9, 8) {real, imag} */,
  {32'h3e337ae9, 32'h00000000} /* (3, 9, 7) {real, imag} */,
  {32'h3c638def, 32'h00000000} /* (3, 9, 6) {real, imag} */,
  {32'hbce0ca68, 32'h00000000} /* (3, 9, 5) {real, imag} */,
  {32'h3e6e21c6, 32'h00000000} /* (3, 9, 4) {real, imag} */,
  {32'hbd88c459, 32'h00000000} /* (3, 9, 3) {real, imag} */,
  {32'hbef4cade, 32'h00000000} /* (3, 9, 2) {real, imag} */,
  {32'h3e310c2f, 32'h00000000} /* (3, 9, 1) {real, imag} */,
  {32'h3e6ee82d, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'h3ea93b90, 32'h00000000} /* (3, 8, 15) {real, imag} */,
  {32'h3f07d90c, 32'h00000000} /* (3, 8, 14) {real, imag} */,
  {32'h3d632d13, 32'h00000000} /* (3, 8, 13) {real, imag} */,
  {32'hbe95288d, 32'h00000000} /* (3, 8, 12) {real, imag} */,
  {32'hbe16f278, 32'h00000000} /* (3, 8, 11) {real, imag} */,
  {32'hbd09b402, 32'h00000000} /* (3, 8, 10) {real, imag} */,
  {32'h3e9e2b2b, 32'h00000000} /* (3, 8, 9) {real, imag} */,
  {32'h3dbcde2f, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'h3db6b564, 32'h00000000} /* (3, 8, 7) {real, imag} */,
  {32'h3f34918c, 32'h00000000} /* (3, 8, 6) {real, imag} */,
  {32'h3eca45d0, 32'h00000000} /* (3, 8, 5) {real, imag} */,
  {32'h3d6213c7, 32'h00000000} /* (3, 8, 4) {real, imag} */,
  {32'hbeaf0648, 32'h00000000} /* (3, 8, 3) {real, imag} */,
  {32'hbf7994e8, 32'h00000000} /* (3, 8, 2) {real, imag} */,
  {32'hbed3cbea, 32'h00000000} /* (3, 8, 1) {real, imag} */,
  {32'h3b883d4e, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'h3d8b207e, 32'h00000000} /* (3, 7, 15) {real, imag} */,
  {32'h3d6f8cbc, 32'h00000000} /* (3, 7, 14) {real, imag} */,
  {32'h3dd7591a, 32'h00000000} /* (3, 7, 13) {real, imag} */,
  {32'hbe8b3ccf, 32'h00000000} /* (3, 7, 12) {real, imag} */,
  {32'hbe79f387, 32'h00000000} /* (3, 7, 11) {real, imag} */,
  {32'h3e0037a7, 32'h00000000} /* (3, 7, 10) {real, imag} */,
  {32'h3f27479c, 32'h00000000} /* (3, 7, 9) {real, imag} */,
  {32'h3df29093, 32'h00000000} /* (3, 7, 8) {real, imag} */,
  {32'hbe8dfe4e, 32'h00000000} /* (3, 7, 7) {real, imag} */,
  {32'hbdf1fd03, 32'h00000000} /* (3, 7, 6) {real, imag} */,
  {32'hbe94e561, 32'h00000000} /* (3, 7, 5) {real, imag} */,
  {32'hbeceb46e, 32'h00000000} /* (3, 7, 4) {real, imag} */,
  {32'hbe70f67b, 32'h00000000} /* (3, 7, 3) {real, imag} */,
  {32'hbf258961, 32'h00000000} /* (3, 7, 2) {real, imag} */,
  {32'hbf1e3dc5, 32'h00000000} /* (3, 7, 1) {real, imag} */,
  {32'hbe8f8b61, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hbc3fe324, 32'h00000000} /* (3, 6, 15) {real, imag} */,
  {32'hbf37b4b4, 32'h00000000} /* (3, 6, 14) {real, imag} */,
  {32'hbee08595, 32'h00000000} /* (3, 6, 13) {real, imag} */,
  {32'hbd8d8145, 32'h00000000} /* (3, 6, 12) {real, imag} */,
  {32'hbe9db993, 32'h00000000} /* (3, 6, 11) {real, imag} */,
  {32'hbd5d8c04, 32'h00000000} /* (3, 6, 10) {real, imag} */,
  {32'h3da53951, 32'h00000000} /* (3, 6, 9) {real, imag} */,
  {32'hbe9059ca, 32'h00000000} /* (3, 6, 8) {real, imag} */,
  {32'hbdeee36b, 32'h00000000} /* (3, 6, 7) {real, imag} */,
  {32'h3e32b77f, 32'h00000000} /* (3, 6, 6) {real, imag} */,
  {32'hbea5c468, 32'h00000000} /* (3, 6, 5) {real, imag} */,
  {32'hbee0d1fa, 32'h00000000} /* (3, 6, 4) {real, imag} */,
  {32'hbdde8df6, 32'h00000000} /* (3, 6, 3) {real, imag} */,
  {32'hbf2808bc, 32'h00000000} /* (3, 6, 2) {real, imag} */,
  {32'hbe60a86b, 32'h00000000} /* (3, 6, 1) {real, imag} */,
  {32'hbe297b6a, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hbe5d4412, 32'h00000000} /* (3, 5, 15) {real, imag} */,
  {32'hbefff48d, 32'h00000000} /* (3, 5, 14) {real, imag} */,
  {32'hbe91f8e2, 32'h00000000} /* (3, 5, 13) {real, imag} */,
  {32'hbe0f9ecf, 32'h00000000} /* (3, 5, 12) {real, imag} */,
  {32'hbeaf635a, 32'h00000000} /* (3, 5, 11) {real, imag} */,
  {32'h3da562ca, 32'h00000000} /* (3, 5, 10) {real, imag} */,
  {32'h3e618a9b, 32'h00000000} /* (3, 5, 9) {real, imag} */,
  {32'h3de66cba, 32'h00000000} /* (3, 5, 8) {real, imag} */,
  {32'h3eac13ac, 32'h00000000} /* (3, 5, 7) {real, imag} */,
  {32'h3ea74db6, 32'h00000000} /* (3, 5, 6) {real, imag} */,
  {32'hbe9a186e, 32'h00000000} /* (3, 5, 5) {real, imag} */,
  {32'hbe1d735f, 32'h00000000} /* (3, 5, 4) {real, imag} */,
  {32'hbe21b3fe, 32'h00000000} /* (3, 5, 3) {real, imag} */,
  {32'hbee09e6d, 32'h00000000} /* (3, 5, 2) {real, imag} */,
  {32'h3ebc8086, 32'h00000000} /* (3, 5, 1) {real, imag} */,
  {32'h3e037405, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hbec755db, 32'h00000000} /* (3, 4, 15) {real, imag} */,
  {32'hbee79f50, 32'h00000000} /* (3, 4, 14) {real, imag} */,
  {32'hbe7b0a83, 32'h00000000} /* (3, 4, 13) {real, imag} */,
  {32'hbd1338b1, 32'h00000000} /* (3, 4, 12) {real, imag} */,
  {32'h3e81daa9, 32'h00000000} /* (3, 4, 11) {real, imag} */,
  {32'h3e896111, 32'h00000000} /* (3, 4, 10) {real, imag} */,
  {32'hbe7d10f7, 32'h00000000} /* (3, 4, 9) {real, imag} */,
  {32'h3e19c1f9, 32'h00000000} /* (3, 4, 8) {real, imag} */,
  {32'hbe57b9ee, 32'h00000000} /* (3, 4, 7) {real, imag} */,
  {32'hbefdebd5, 32'h00000000} /* (3, 4, 6) {real, imag} */,
  {32'hbda07906, 32'h00000000} /* (3, 4, 5) {real, imag} */,
  {32'hbe1551ef, 32'h00000000} /* (3, 4, 4) {real, imag} */,
  {32'hbe2738d6, 32'h00000000} /* (3, 4, 3) {real, imag} */,
  {32'hbecce9fc, 32'h00000000} /* (3, 4, 2) {real, imag} */,
  {32'hbe5afbb4, 32'h00000000} /* (3, 4, 1) {real, imag} */,
  {32'hbde36964, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hbe960291, 32'h00000000} /* (3, 3, 15) {real, imag} */,
  {32'hbf1d1aae, 32'h00000000} /* (3, 3, 14) {real, imag} */,
  {32'hbf091e70, 32'h00000000} /* (3, 3, 13) {real, imag} */,
  {32'hbd398250, 32'h00000000} /* (3, 3, 12) {real, imag} */,
  {32'h3e6e173c, 32'h00000000} /* (3, 3, 11) {real, imag} */,
  {32'hbe5934e1, 32'h00000000} /* (3, 3, 10) {real, imag} */,
  {32'hbe3ba1a5, 32'h00000000} /* (3, 3, 9) {real, imag} */,
  {32'h3d7c12cf, 32'h00000000} /* (3, 3, 8) {real, imag} */,
  {32'hbe12afb4, 32'h00000000} /* (3, 3, 7) {real, imag} */,
  {32'hbee6f33d, 32'h00000000} /* (3, 3, 6) {real, imag} */,
  {32'hbd1a0c09, 32'h00000000} /* (3, 3, 5) {real, imag} */,
  {32'hbe2eb6a5, 32'h00000000} /* (3, 3, 4) {real, imag} */,
  {32'hbe24ede5, 32'h00000000} /* (3, 3, 3) {real, imag} */,
  {32'h3d0de88a, 32'h00000000} /* (3, 3, 2) {real, imag} */,
  {32'h3d604a05, 32'h00000000} /* (3, 3, 1) {real, imag} */,
  {32'hbb8f14df, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hbea31a1a, 32'h00000000} /* (3, 2, 15) {real, imag} */,
  {32'hbeaad315, 32'h00000000} /* (3, 2, 14) {real, imag} */,
  {32'hbbbab1eb, 32'h00000000} /* (3, 2, 13) {real, imag} */,
  {32'h3e79661f, 32'h00000000} /* (3, 2, 12) {real, imag} */,
  {32'h3e0882c6, 32'h00000000} /* (3, 2, 11) {real, imag} */,
  {32'hbe1fa57c, 32'h00000000} /* (3, 2, 10) {real, imag} */,
  {32'hbe30c73f, 32'h00000000} /* (3, 2, 9) {real, imag} */,
  {32'hbdc9eae1, 32'h00000000} /* (3, 2, 8) {real, imag} */,
  {32'hbc96eb1a, 32'h00000000} /* (3, 2, 7) {real, imag} */,
  {32'h3d83b2a7, 32'h00000000} /* (3, 2, 6) {real, imag} */,
  {32'hbea19e55, 32'h00000000} /* (3, 2, 5) {real, imag} */,
  {32'hbf457d1a, 32'h00000000} /* (3, 2, 4) {real, imag} */,
  {32'hbf071470, 32'h00000000} /* (3, 2, 3) {real, imag} */,
  {32'hbe553e52, 32'h00000000} /* (3, 2, 2) {real, imag} */,
  {32'hbe4477f0, 32'h00000000} /* (3, 2, 1) {real, imag} */,
  {32'h3d7172ea, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hbe88adc3, 32'h00000000} /* (3, 1, 15) {real, imag} */,
  {32'hbe1f5eb8, 32'h00000000} /* (3, 1, 14) {real, imag} */,
  {32'h3f194ede, 32'h00000000} /* (3, 1, 13) {real, imag} */,
  {32'h3f04bc5f, 32'h00000000} /* (3, 1, 12) {real, imag} */,
  {32'h3e401bca, 32'h00000000} /* (3, 1, 11) {real, imag} */,
  {32'hbe14e540, 32'h00000000} /* (3, 1, 10) {real, imag} */,
  {32'hbeba8484, 32'h00000000} /* (3, 1, 9) {real, imag} */,
  {32'hbe8097c9, 32'h00000000} /* (3, 1, 8) {real, imag} */,
  {32'hbe6c5bc7, 32'h00000000} /* (3, 1, 7) {real, imag} */,
  {32'h3e43a9b5, 32'h00000000} /* (3, 1, 6) {real, imag} */,
  {32'hbd922ca6, 32'h00000000} /* (3, 1, 5) {real, imag} */,
  {32'hbeeaf5dd, 32'h00000000} /* (3, 1, 4) {real, imag} */,
  {32'h3dd7a32f, 32'h00000000} /* (3, 1, 3) {real, imag} */,
  {32'h3eee28d4, 32'h00000000} /* (3, 1, 2) {real, imag} */,
  {32'hbe334fdc, 32'h00000000} /* (3, 1, 1) {real, imag} */,
  {32'h3d0c82e7, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hbe7dd0c1, 32'h00000000} /* (3, 0, 15) {real, imag} */,
  {32'h3e0ac90b, 32'h00000000} /* (3, 0, 14) {real, imag} */,
  {32'h3f5694ad, 32'h00000000} /* (3, 0, 13) {real, imag} */,
  {32'h3ed002aa, 32'h00000000} /* (3, 0, 12) {real, imag} */,
  {32'hbc8db1d8, 32'h00000000} /* (3, 0, 11) {real, imag} */,
  {32'hbd51e76b, 32'h00000000} /* (3, 0, 10) {real, imag} */,
  {32'hbe252541, 32'h00000000} /* (3, 0, 9) {real, imag} */,
  {32'hbde8c7a2, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'hbee3225b, 32'h00000000} /* (3, 0, 7) {real, imag} */,
  {32'hbd940411, 32'h00000000} /* (3, 0, 6) {real, imag} */,
  {32'h3e944933, 32'h00000000} /* (3, 0, 5) {real, imag} */,
  {32'h3ea56d1d, 32'h00000000} /* (3, 0, 4) {real, imag} */,
  {32'h3daea814, 32'h00000000} /* (3, 0, 3) {real, imag} */,
  {32'h3ed940f3, 32'h00000000} /* (3, 0, 2) {real, imag} */,
  {32'h3eb72165, 32'h00000000} /* (3, 0, 1) {real, imag} */,
  {32'h3dc4cc02, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hbdf322f2, 32'h00000000} /* (2, 15, 15) {real, imag} */,
  {32'hbd8d0a9e, 32'h00000000} /* (2, 15, 14) {real, imag} */,
  {32'hbcbf1003, 32'h00000000} /* (2, 15, 13) {real, imag} */,
  {32'hbd446659, 32'h00000000} /* (2, 15, 12) {real, imag} */,
  {32'h3e4924ce, 32'h00000000} /* (2, 15, 11) {real, imag} */,
  {32'h3e97ccac, 32'h00000000} /* (2, 15, 10) {real, imag} */,
  {32'h3e56efca, 32'h00000000} /* (2, 15, 9) {real, imag} */,
  {32'h3eac6f81, 32'h00000000} /* (2, 15, 8) {real, imag} */,
  {32'h3f00ebaa, 32'h00000000} /* (2, 15, 7) {real, imag} */,
  {32'h3c92f36b, 32'h00000000} /* (2, 15, 6) {real, imag} */,
  {32'hbe961767, 32'h00000000} /* (2, 15, 5) {real, imag} */,
  {32'hbea06d86, 32'h00000000} /* (2, 15, 4) {real, imag} */,
  {32'hbee2a8ed, 32'h00000000} /* (2, 15, 3) {real, imag} */,
  {32'hbe6b7e03, 32'h00000000} /* (2, 15, 2) {real, imag} */,
  {32'hbe17a15f, 32'h00000000} /* (2, 15, 1) {real, imag} */,
  {32'hbea81f7b, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h3ea79ec7, 32'h00000000} /* (2, 14, 15) {real, imag} */,
  {32'h3dbbb4bf, 32'h00000000} /* (2, 14, 14) {real, imag} */,
  {32'hbea695c4, 32'h00000000} /* (2, 14, 13) {real, imag} */,
  {32'hbe3e5fcc, 32'h00000000} /* (2, 14, 12) {real, imag} */,
  {32'h3d230d32, 32'h00000000} /* (2, 14, 11) {real, imag} */,
  {32'hbd5c5688, 32'h00000000} /* (2, 14, 10) {real, imag} */,
  {32'hbe80cdfe, 32'h00000000} /* (2, 14, 9) {real, imag} */,
  {32'h3ece9a59, 32'h00000000} /* (2, 14, 8) {real, imag} */,
  {32'h3e9bdb07, 32'h00000000} /* (2, 14, 7) {real, imag} */,
  {32'hbca1223f, 32'h00000000} /* (2, 14, 6) {real, imag} */,
  {32'hbd9d1374, 32'h00000000} /* (2, 14, 5) {real, imag} */,
  {32'hbe46991e, 32'h00000000} /* (2, 14, 4) {real, imag} */,
  {32'hbe99f5ef, 32'h00000000} /* (2, 14, 3) {real, imag} */,
  {32'hbef1f2b7, 32'h00000000} /* (2, 14, 2) {real, imag} */,
  {32'hbe8bdee6, 32'h00000000} /* (2, 14, 1) {real, imag} */,
  {32'h3df3b49d, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h3eb78aaa, 32'h00000000} /* (2, 13, 15) {real, imag} */,
  {32'hbeed6a0f, 32'h00000000} /* (2, 13, 14) {real, imag} */,
  {32'hbed8058d, 32'h00000000} /* (2, 13, 13) {real, imag} */,
  {32'h3d37ce3f, 32'h00000000} /* (2, 13, 12) {real, imag} */,
  {32'hbdba8ef6, 32'h00000000} /* (2, 13, 11) {real, imag} */,
  {32'hbed4fd04, 32'h00000000} /* (2, 13, 10) {real, imag} */,
  {32'hbf257b77, 32'h00000000} /* (2, 13, 9) {real, imag} */,
  {32'h3e67ffeb, 32'h00000000} /* (2, 13, 8) {real, imag} */,
  {32'h3e95aebd, 32'h00000000} /* (2, 13, 7) {real, imag} */,
  {32'h3dc8883a, 32'h00000000} /* (2, 13, 6) {real, imag} */,
  {32'h3e69d047, 32'h00000000} /* (2, 13, 5) {real, imag} */,
  {32'h3c841ae2, 32'h00000000} /* (2, 13, 4) {real, imag} */,
  {32'hbe3c9fee, 32'h00000000} /* (2, 13, 3) {real, imag} */,
  {32'hbf19cad2, 32'h00000000} /* (2, 13, 2) {real, imag} */,
  {32'hbcaaf105, 32'h00000000} /* (2, 13, 1) {real, imag} */,
  {32'h3f16c84b, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h3cf6b635, 32'h00000000} /* (2, 12, 15) {real, imag} */,
  {32'hbe8f5fc1, 32'h00000000} /* (2, 12, 14) {real, imag} */,
  {32'h3e804137, 32'h00000000} /* (2, 12, 13) {real, imag} */,
  {32'h3e4e4495, 32'h00000000} /* (2, 12, 12) {real, imag} */,
  {32'hbec063c4, 32'h00000000} /* (2, 12, 11) {real, imag} */,
  {32'hbe97f080, 32'h00000000} /* (2, 12, 10) {real, imag} */,
  {32'hbda03aa6, 32'h00000000} /* (2, 12, 9) {real, imag} */,
  {32'h3e5a4e1f, 32'h00000000} /* (2, 12, 8) {real, imag} */,
  {32'h3e4e141a, 32'h00000000} /* (2, 12, 7) {real, imag} */,
  {32'h3e6b5924, 32'h00000000} /* (2, 12, 6) {real, imag} */,
  {32'h3f2817b5, 32'h00000000} /* (2, 12, 5) {real, imag} */,
  {32'h3e1eb8b1, 32'h00000000} /* (2, 12, 4) {real, imag} */,
  {32'hbe973006, 32'h00000000} /* (2, 12, 3) {real, imag} */,
  {32'hbec76f53, 32'h00000000} /* (2, 12, 2) {real, imag} */,
  {32'h3d740bf4, 32'h00000000} /* (2, 12, 1) {real, imag} */,
  {32'h3e0d1308, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h3dae0a71, 32'h00000000} /* (2, 11, 15) {real, imag} */,
  {32'h3e836e75, 32'h00000000} /* (2, 11, 14) {real, imag} */,
  {32'h3f4e9880, 32'h00000000} /* (2, 11, 13) {real, imag} */,
  {32'h3ec8caa8, 32'h00000000} /* (2, 11, 12) {real, imag} */,
  {32'h3d3631db, 32'h00000000} /* (2, 11, 11) {real, imag} */,
  {32'hbe939a68, 32'h00000000} /* (2, 11, 10) {real, imag} */,
  {32'hbca24699, 32'h00000000} /* (2, 11, 9) {real, imag} */,
  {32'h3e696558, 32'h00000000} /* (2, 11, 8) {real, imag} */,
  {32'hbeddf36f, 32'h00000000} /* (2, 11, 7) {real, imag} */,
  {32'hbed237d6, 32'h00000000} /* (2, 11, 6) {real, imag} */,
  {32'h3e744269, 32'h00000000} /* (2, 11, 5) {real, imag} */,
  {32'h3e103446, 32'h00000000} /* (2, 11, 4) {real, imag} */,
  {32'hbe6c2567, 32'h00000000} /* (2, 11, 3) {real, imag} */,
  {32'hbe4cce0c, 32'h00000000} /* (2, 11, 2) {real, imag} */,
  {32'hbd2ad03c, 32'h00000000} /* (2, 11, 1) {real, imag} */,
  {32'h3e1da49d, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'h3ed1088e, 32'h00000000} /* (2, 10, 15) {real, imag} */,
  {32'h3e766232, 32'h00000000} /* (2, 10, 14) {real, imag} */,
  {32'hbe0c7185, 32'h00000000} /* (2, 10, 13) {real, imag} */,
  {32'h3e0c2a92, 32'h00000000} /* (2, 10, 12) {real, imag} */,
  {32'h3ea2c133, 32'h00000000} /* (2, 10, 11) {real, imag} */,
  {32'h3db17901, 32'h00000000} /* (2, 10, 10) {real, imag} */,
  {32'hbea553a5, 32'h00000000} /* (2, 10, 9) {real, imag} */,
  {32'hbf10bc22, 32'h00000000} /* (2, 10, 8) {real, imag} */,
  {32'hbef73d6f, 32'h00000000} /* (2, 10, 7) {real, imag} */,
  {32'h3da3598c, 32'h00000000} /* (2, 10, 6) {real, imag} */,
  {32'h3c93ba12, 32'h00000000} /* (2, 10, 5) {real, imag} */,
  {32'hbdffe8dc, 32'h00000000} /* (2, 10, 4) {real, imag} */,
  {32'hbeed0972, 32'h00000000} /* (2, 10, 3) {real, imag} */,
  {32'hbe4cbefa, 32'h00000000} /* (2, 10, 2) {real, imag} */,
  {32'h3cf124cb, 32'h00000000} /* (2, 10, 1) {real, imag} */,
  {32'h3e482efc, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'h3ecf7b8a, 32'h00000000} /* (2, 9, 15) {real, imag} */,
  {32'h3f241ca1, 32'h00000000} /* (2, 9, 14) {real, imag} */,
  {32'h3ea08288, 32'h00000000} /* (2, 9, 13) {real, imag} */,
  {32'h3df8e510, 32'h00000000} /* (2, 9, 12) {real, imag} */,
  {32'h3e678537, 32'h00000000} /* (2, 9, 11) {real, imag} */,
  {32'h3ededbd8, 32'h00000000} /* (2, 9, 10) {real, imag} */,
  {32'h3e4d86f4, 32'h00000000} /* (2, 9, 9) {real, imag} */,
  {32'hbe0834b2, 32'h00000000} /* (2, 9, 8) {real, imag} */,
  {32'h3ed10689, 32'h00000000} /* (2, 9, 7) {real, imag} */,
  {32'h3e8dbb2b, 32'h00000000} /* (2, 9, 6) {real, imag} */,
  {32'h3ef15a0d, 32'h00000000} /* (2, 9, 5) {real, imag} */,
  {32'h3f0fc9a6, 32'h00000000} /* (2, 9, 4) {real, imag} */,
  {32'h3ef154eb, 32'h00000000} /* (2, 9, 3) {real, imag} */,
  {32'hbd0d679c, 32'h00000000} /* (2, 9, 2) {real, imag} */,
  {32'h3e89cbd5, 32'h00000000} /* (2, 9, 1) {real, imag} */,
  {32'h3e4e98f5, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'h3f1c2d78, 32'h00000000} /* (2, 8, 15) {real, imag} */,
  {32'h3f9e507c, 32'h00000000} /* (2, 8, 14) {real, imag} */,
  {32'h3f153a8e, 32'h00000000} /* (2, 8, 13) {real, imag} */,
  {32'h3cf0aed2, 32'h00000000} /* (2, 8, 12) {real, imag} */,
  {32'h3e8bddc2, 32'h00000000} /* (2, 8, 11) {real, imag} */,
  {32'h3e5e4972, 32'h00000000} /* (2, 8, 10) {real, imag} */,
  {32'h3eb04906, 32'h00000000} /* (2, 8, 9) {real, imag} */,
  {32'h3e6a8cc6, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'h3f182c62, 32'h00000000} /* (2, 8, 7) {real, imag} */,
  {32'h3dd97a9b, 32'h00000000} /* (2, 8, 6) {real, imag} */,
  {32'h3e064440, 32'h00000000} /* (2, 8, 5) {real, imag} */,
  {32'h3f0de0e1, 32'h00000000} /* (2, 8, 4) {real, imag} */,
  {32'h3ef43e80, 32'h00000000} /* (2, 8, 3) {real, imag} */,
  {32'hbeb4c020, 32'h00000000} /* (2, 8, 2) {real, imag} */,
  {32'hbee65494, 32'h00000000} /* (2, 8, 1) {real, imag} */,
  {32'h3d9ad0c8, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'h3e9be504, 32'h00000000} /* (2, 7, 15) {real, imag} */,
  {32'h3edf87c0, 32'h00000000} /* (2, 7, 14) {real, imag} */,
  {32'h3f3704b5, 32'h00000000} /* (2, 7, 13) {real, imag} */,
  {32'h3e86f589, 32'h00000000} /* (2, 7, 12) {real, imag} */,
  {32'h3e899a66, 32'h00000000} /* (2, 7, 11) {real, imag} */,
  {32'hbea370f3, 32'h00000000} /* (2, 7, 10) {real, imag} */,
  {32'hbd6c484a, 32'h00000000} /* (2, 7, 9) {real, imag} */,
  {32'h3eb0a180, 32'h00000000} /* (2, 7, 8) {real, imag} */,
  {32'h3e437879, 32'h00000000} /* (2, 7, 7) {real, imag} */,
  {32'hbf088964, 32'h00000000} /* (2, 7, 6) {real, imag} */,
  {32'hbf026e45, 32'h00000000} /* (2, 7, 5) {real, imag} */,
  {32'h3ceb2111, 32'h00000000} /* (2, 7, 4) {real, imag} */,
  {32'h3c5e19b3, 32'h00000000} /* (2, 7, 3) {real, imag} */,
  {32'hbeff133d, 32'h00000000} /* (2, 7, 2) {real, imag} */,
  {32'hbe5d1ad8, 32'h00000000} /* (2, 7, 1) {real, imag} */,
  {32'h3f089390, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'h3e2f33e8, 32'h00000000} /* (2, 6, 15) {real, imag} */,
  {32'hbe972dbd, 32'h00000000} /* (2, 6, 14) {real, imag} */,
  {32'h3e9c6b42, 32'h00000000} /* (2, 6, 13) {real, imag} */,
  {32'h3f481d82, 32'h00000000} /* (2, 6, 12) {real, imag} */,
  {32'h3c8ccf7c, 32'h00000000} /* (2, 6, 11) {real, imag} */,
  {32'hbea1212d, 32'h00000000} /* (2, 6, 10) {real, imag} */,
  {32'hbe3b832a, 32'h00000000} /* (2, 6, 9) {real, imag} */,
  {32'hbdbaf21c, 32'h00000000} /* (2, 6, 8) {real, imag} */,
  {32'hbce2f89e, 32'h00000000} /* (2, 6, 7) {real, imag} */,
  {32'hbe232ed8, 32'h00000000} /* (2, 6, 6) {real, imag} */,
  {32'hbec7b5c5, 32'h00000000} /* (2, 6, 5) {real, imag} */,
  {32'hbdd9bd4a, 32'h00000000} /* (2, 6, 4) {real, imag} */,
  {32'hbe84acc3, 32'h00000000} /* (2, 6, 3) {real, imag} */,
  {32'hbf371cf6, 32'h00000000} /* (2, 6, 2) {real, imag} */,
  {32'h3dd170e9, 32'h00000000} /* (2, 6, 1) {real, imag} */,
  {32'h3ed329a6, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hbe81573b, 32'h00000000} /* (2, 5, 15) {real, imag} */,
  {32'hbf07d761, 32'h00000000} /* (2, 5, 14) {real, imag} */,
  {32'hbbf0ae5f, 32'h00000000} /* (2, 5, 13) {real, imag} */,
  {32'h3e487c9e, 32'h00000000} /* (2, 5, 12) {real, imag} */,
  {32'hbda6b1fe, 32'h00000000} /* (2, 5, 11) {real, imag} */,
  {32'h3cba6e66, 32'h00000000} /* (2, 5, 10) {real, imag} */,
  {32'hbd6b9c1d, 32'h00000000} /* (2, 5, 9) {real, imag} */,
  {32'h3e1e070b, 32'h00000000} /* (2, 5, 8) {real, imag} */,
  {32'h3c3929b5, 32'h00000000} /* (2, 5, 7) {real, imag} */,
  {32'hbed12380, 32'h00000000} /* (2, 5, 6) {real, imag} */,
  {32'hbf1a12bc, 32'h00000000} /* (2, 5, 5) {real, imag} */,
  {32'hbe1f25a5, 32'h00000000} /* (2, 5, 4) {real, imag} */,
  {32'hbec2d7fb, 32'h00000000} /* (2, 5, 3) {real, imag} */,
  {32'hbe80a3b7, 32'h00000000} /* (2, 5, 2) {real, imag} */,
  {32'h3f4dfe58, 32'h00000000} /* (2, 5, 1) {real, imag} */,
  {32'h3e9567bf, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hbecf937c, 32'h00000000} /* (2, 4, 15) {real, imag} */,
  {32'hbed15b15, 32'h00000000} /* (2, 4, 14) {real, imag} */,
  {32'h3e0a80e2, 32'h00000000} /* (2, 4, 13) {real, imag} */,
  {32'hbe46b572, 32'h00000000} /* (2, 4, 12) {real, imag} */,
  {32'h3df316bc, 32'h00000000} /* (2, 4, 11) {real, imag} */,
  {32'h3ed48148, 32'h00000000} /* (2, 4, 10) {real, imag} */,
  {32'hbd7535a1, 32'h00000000} /* (2, 4, 9) {real, imag} */,
  {32'h3e92df3e, 32'h00000000} /* (2, 4, 8) {real, imag} */,
  {32'hbd20098d, 32'h00000000} /* (2, 4, 7) {real, imag} */,
  {32'hbeeaff5b, 32'h00000000} /* (2, 4, 6) {real, imag} */,
  {32'hbeb895b2, 32'h00000000} /* (2, 4, 5) {real, imag} */,
  {32'hbe894ee2, 32'h00000000} /* (2, 4, 4) {real, imag} */,
  {32'hbc0280b8, 32'h00000000} /* (2, 4, 3) {real, imag} */,
  {32'h3d0988b0, 32'h00000000} /* (2, 4, 2) {real, imag} */,
  {32'h3f06a834, 32'h00000000} /* (2, 4, 1) {real, imag} */,
  {32'h3ddbe57b, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hbeb0ec6a, 32'h00000000} /* (2, 3, 15) {real, imag} */,
  {32'hbe8c8b35, 32'h00000000} /* (2, 3, 14) {real, imag} */,
  {32'h3e943931, 32'h00000000} /* (2, 3, 13) {real, imag} */,
  {32'h3d33583a, 32'h00000000} /* (2, 3, 12) {real, imag} */,
  {32'h3e927c34, 32'h00000000} /* (2, 3, 11) {real, imag} */,
  {32'h3ea7907e, 32'h00000000} /* (2, 3, 10) {real, imag} */,
  {32'hbd95a37f, 32'h00000000} /* (2, 3, 9) {real, imag} */,
  {32'h3a708c6e, 32'h00000000} /* (2, 3, 8) {real, imag} */,
  {32'hbe89b205, 32'h00000000} /* (2, 3, 7) {real, imag} */,
  {32'hbeed80e7, 32'h00000000} /* (2, 3, 6) {real, imag} */,
  {32'hbea5baf4, 32'h00000000} /* (2, 3, 5) {real, imag} */,
  {32'h3cd8a6b8, 32'h00000000} /* (2, 3, 4) {real, imag} */,
  {32'h3e89fc8f, 32'h00000000} /* (2, 3, 3) {real, imag} */,
  {32'h3eba825b, 32'h00000000} /* (2, 3, 2) {real, imag} */,
  {32'h3ebba6d1, 32'h00000000} /* (2, 3, 1) {real, imag} */,
  {32'h3e80a798, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hbdb2a8a6, 32'h00000000} /* (2, 2, 15) {real, imag} */,
  {32'h3d3c596a, 32'h00000000} /* (2, 2, 14) {real, imag} */,
  {32'h3ddae4bd, 32'h00000000} /* (2, 2, 13) {real, imag} */,
  {32'h3e8a1b8c, 32'h00000000} /* (2, 2, 12) {real, imag} */,
  {32'h3ec486e6, 32'h00000000} /* (2, 2, 11) {real, imag} */,
  {32'hbd56ba13, 32'h00000000} /* (2, 2, 10) {real, imag} */,
  {32'hbeac2ce0, 32'h00000000} /* (2, 2, 9) {real, imag} */,
  {32'hbde4bac0, 32'h00000000} /* (2, 2, 8) {real, imag} */,
  {32'h3eabd73c, 32'h00000000} /* (2, 2, 7) {real, imag} */,
  {32'h3e7251a9, 32'h00000000} /* (2, 2, 6) {real, imag} */,
  {32'hbe575d5e, 32'h00000000} /* (2, 2, 5) {real, imag} */,
  {32'hbe673a30, 32'h00000000} /* (2, 2, 4) {real, imag} */,
  {32'hbbfc189e, 32'h00000000} /* (2, 2, 3) {real, imag} */,
  {32'hbe9a79e5, 32'h00000000} /* (2, 2, 2) {real, imag} */,
  {32'hbdfce111, 32'h00000000} /* (2, 2, 1) {real, imag} */,
  {32'h3e82dd93, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hbea4ac85, 32'h00000000} /* (2, 1, 15) {real, imag} */,
  {32'hbeeaac3c, 32'h00000000} /* (2, 1, 14) {real, imag} */,
  {32'h3cc3b8a3, 32'h00000000} /* (2, 1, 13) {real, imag} */,
  {32'h3eb59416, 32'h00000000} /* (2, 1, 12) {real, imag} */,
  {32'h3ee63f0e, 32'h00000000} /* (2, 1, 11) {real, imag} */,
  {32'h3d3047de, 32'h00000000} /* (2, 1, 10) {real, imag} */,
  {32'hbdbaef48, 32'h00000000} /* (2, 1, 9) {real, imag} */,
  {32'hbef81546, 32'h00000000} /* (2, 1, 8) {real, imag} */,
  {32'h3e76c2a6, 32'h00000000} /* (2, 1, 7) {real, imag} */,
  {32'h3f0e25f4, 32'h00000000} /* (2, 1, 6) {real, imag} */,
  {32'hbcbdf257, 32'h00000000} /* (2, 1, 5) {real, imag} */,
  {32'hbe801136, 32'h00000000} /* (2, 1, 4) {real, imag} */,
  {32'hbdd37d8c, 32'h00000000} /* (2, 1, 3) {real, imag} */,
  {32'hbdfc08bf, 32'h00000000} /* (2, 1, 2) {real, imag} */,
  {32'hbc1558e0, 32'h00000000} /* (2, 1, 1) {real, imag} */,
  {32'h3dd958bd, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hbe3d1b15, 32'h00000000} /* (2, 0, 15) {real, imag} */,
  {32'hbe8c6d4e, 32'h00000000} /* (2, 0, 14) {real, imag} */,
  {32'h3e3595b6, 32'h00000000} /* (2, 0, 13) {real, imag} */,
  {32'h3f0f8133, 32'h00000000} /* (2, 0, 12) {real, imag} */,
  {32'h3eaa31a2, 32'h00000000} /* (2, 0, 11) {real, imag} */,
  {32'h3d98a1d0, 32'h00000000} /* (2, 0, 10) {real, imag} */,
  {32'h3dd93618, 32'h00000000} /* (2, 0, 9) {real, imag} */,
  {32'hbe75b1b0, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'h3dc983c8, 32'h00000000} /* (2, 0, 7) {real, imag} */,
  {32'h3e8c5e7d, 32'h00000000} /* (2, 0, 6) {real, imag} */,
  {32'hbdbe2635, 32'h00000000} /* (2, 0, 5) {real, imag} */,
  {32'h3af76150, 32'h00000000} /* (2, 0, 4) {real, imag} */,
  {32'h3dea73ad, 32'h00000000} /* (2, 0, 3) {real, imag} */,
  {32'h3ebc8559, 32'h00000000} /* (2, 0, 2) {real, imag} */,
  {32'h3e83e7bc, 32'h00000000} /* (2, 0, 1) {real, imag} */,
  {32'hbc9f3b95, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'h3d58ff9e, 32'h00000000} /* (1, 15, 15) {real, imag} */,
  {32'h3c89e186, 32'h00000000} /* (1, 15, 14) {real, imag} */,
  {32'hbd621ade, 32'h00000000} /* (1, 15, 13) {real, imag} */,
  {32'hbd7414ef, 32'h00000000} /* (1, 15, 12) {real, imag} */,
  {32'h3e7d3a2e, 32'h00000000} /* (1, 15, 11) {real, imag} */,
  {32'h3e7d7215, 32'h00000000} /* (1, 15, 10) {real, imag} */,
  {32'hbdb0512a, 32'h00000000} /* (1, 15, 9) {real, imag} */,
  {32'h3e18fe06, 32'h00000000} /* (1, 15, 8) {real, imag} */,
  {32'h3e90c163, 32'h00000000} /* (1, 15, 7) {real, imag} */,
  {32'h3e0aab54, 32'h00000000} /* (1, 15, 6) {real, imag} */,
  {32'hbe9a955f, 32'h00000000} /* (1, 15, 5) {real, imag} */,
  {32'hbe82fa12, 32'h00000000} /* (1, 15, 4) {real, imag} */,
  {32'hbecae4ce, 32'h00000000} /* (1, 15, 3) {real, imag} */,
  {32'hbe91f055, 32'h00000000} /* (1, 15, 2) {real, imag} */,
  {32'hbd73862a, 32'h00000000} /* (1, 15, 1) {real, imag} */,
  {32'hbe39bb89, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'h3ddeeef1, 32'h00000000} /* (1, 14, 15) {real, imag} */,
  {32'h3d36af58, 32'h00000000} /* (1, 14, 14) {real, imag} */,
  {32'hbe33c83e, 32'h00000000} /* (1, 14, 13) {real, imag} */,
  {32'hbd4edc3c, 32'h00000000} /* (1, 14, 12) {real, imag} */,
  {32'h3ee95821, 32'h00000000} /* (1, 14, 11) {real, imag} */,
  {32'h3e8dd432, 32'h00000000} /* (1, 14, 10) {real, imag} */,
  {32'h3cedf555, 32'h00000000} /* (1, 14, 9) {real, imag} */,
  {32'h3e4cc073, 32'h00000000} /* (1, 14, 8) {real, imag} */,
  {32'h3e9dcc35, 32'h00000000} /* (1, 14, 7) {real, imag} */,
  {32'h3f108d0d, 32'h00000000} /* (1, 14, 6) {real, imag} */,
  {32'h3d100f88, 32'h00000000} /* (1, 14, 5) {real, imag} */,
  {32'hbca4c0d9, 32'h00000000} /* (1, 14, 4) {real, imag} */,
  {32'hbee423f0, 32'h00000000} /* (1, 14, 3) {real, imag} */,
  {32'hbf12e75a, 32'h00000000} /* (1, 14, 2) {real, imag} */,
  {32'h3d105651, 32'h00000000} /* (1, 14, 1) {real, imag} */,
  {32'h3d1ab27e, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h3d6523cd, 32'h00000000} /* (1, 13, 15) {real, imag} */,
  {32'hbe69acb7, 32'h00000000} /* (1, 13, 14) {real, imag} */,
  {32'hbea8a962, 32'h00000000} /* (1, 13, 13) {real, imag} */,
  {32'h3e3f64da, 32'h00000000} /* (1, 13, 12) {real, imag} */,
  {32'h3eaa3d87, 32'h00000000} /* (1, 13, 11) {real, imag} */,
  {32'h3b67d844, 32'h00000000} /* (1, 13, 10) {real, imag} */,
  {32'hbdb0bc47, 32'h00000000} /* (1, 13, 9) {real, imag} */,
  {32'h3e2bebe9, 32'h00000000} /* (1, 13, 8) {real, imag} */,
  {32'h3c6753bc, 32'h00000000} /* (1, 13, 7) {real, imag} */,
  {32'h3dfdea3d, 32'h00000000} /* (1, 13, 6) {real, imag} */,
  {32'h3de91f70, 32'h00000000} /* (1, 13, 5) {real, imag} */,
  {32'hba8b0b3b, 32'h00000000} /* (1, 13, 4) {real, imag} */,
  {32'h3cccb7ad, 32'h00000000} /* (1, 13, 3) {real, imag} */,
  {32'hbe88a515, 32'h00000000} /* (1, 13, 2) {real, imag} */,
  {32'h3dc2ebc6, 32'h00000000} /* (1, 13, 1) {real, imag} */,
  {32'h3ee9f471, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'hbe6d20a8, 32'h00000000} /* (1, 12, 15) {real, imag} */,
  {32'hbe9f730e, 32'h00000000} /* (1, 12, 14) {real, imag} */,
  {32'h3e9c1592, 32'h00000000} /* (1, 12, 13) {real, imag} */,
  {32'h3ebe83f6, 32'h00000000} /* (1, 12, 12) {real, imag} */,
  {32'hbde6010a, 32'h00000000} /* (1, 12, 11) {real, imag} */,
  {32'hbe4525e1, 32'h00000000} /* (1, 12, 10) {real, imag} */,
  {32'hbe8209e4, 32'h00000000} /* (1, 12, 9) {real, imag} */,
  {32'hbef58b2f, 32'h00000000} /* (1, 12, 8) {real, imag} */,
  {32'hbf3ab53f, 32'h00000000} /* (1, 12, 7) {real, imag} */,
  {32'hbf1d50b4, 32'h00000000} /* (1, 12, 6) {real, imag} */,
  {32'hbe35ae7d, 32'h00000000} /* (1, 12, 5) {real, imag} */,
  {32'hbc8b0ffd, 32'h00000000} /* (1, 12, 4) {real, imag} */,
  {32'h3ecd6508, 32'h00000000} /* (1, 12, 3) {real, imag} */,
  {32'h3e9f2ec3, 32'h00000000} /* (1, 12, 2) {real, imag} */,
  {32'h3edd3b1f, 32'h00000000} /* (1, 12, 1) {real, imag} */,
  {32'h3e81d074, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'hbd424093, 32'h00000000} /* (1, 11, 15) {real, imag} */,
  {32'h3ebd0a74, 32'h00000000} /* (1, 11, 14) {real, imag} */,
  {32'h3f89bcb0, 32'h00000000} /* (1, 11, 13) {real, imag} */,
  {32'h3f4b2d09, 32'h00000000} /* (1, 11, 12) {real, imag} */,
  {32'h3dbcc3ab, 32'h00000000} /* (1, 11, 11) {real, imag} */,
  {32'h3e1f04bd, 32'h00000000} /* (1, 11, 10) {real, imag} */,
  {32'h3eae33f0, 32'h00000000} /* (1, 11, 9) {real, imag} */,
  {32'h3e533a6f, 32'h00000000} /* (1, 11, 8) {real, imag} */,
  {32'hbe98a7a2, 32'h00000000} /* (1, 11, 7) {real, imag} */,
  {32'hbdfefd2a, 32'h00000000} /* (1, 11, 6) {real, imag} */,
  {32'h3e0e8b82, 32'h00000000} /* (1, 11, 5) {real, imag} */,
  {32'h3d92ff7d, 32'h00000000} /* (1, 11, 4) {real, imag} */,
  {32'hbe86ee39, 32'h00000000} /* (1, 11, 3) {real, imag} */,
  {32'hbedc195c, 32'h00000000} /* (1, 11, 2) {real, imag} */,
  {32'h3e1d85fd, 32'h00000000} /* (1, 11, 1) {real, imag} */,
  {32'h3d83cc8f, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'h3eb68228, 32'h00000000} /* (1, 10, 15) {real, imag} */,
  {32'h3f2ac95d, 32'h00000000} /* (1, 10, 14) {real, imag} */,
  {32'h3ec0407e, 32'h00000000} /* (1, 10, 13) {real, imag} */,
  {32'h3f12bf8a, 32'h00000000} /* (1, 10, 12) {real, imag} */,
  {32'h3ec6582f, 32'h00000000} /* (1, 10, 11) {real, imag} */,
  {32'h3ee6b0f5, 32'h00000000} /* (1, 10, 10) {real, imag} */,
  {32'h3f2df550, 32'h00000000} /* (1, 10, 9) {real, imag} */,
  {32'h3f06efd6, 32'h00000000} /* (1, 10, 8) {real, imag} */,
  {32'h3c968cbc, 32'h00000000} /* (1, 10, 7) {real, imag} */,
  {32'h3e1602db, 32'h00000000} /* (1, 10, 6) {real, imag} */,
  {32'hbe7025df, 32'h00000000} /* (1, 10, 5) {real, imag} */,
  {32'hbea76244, 32'h00000000} /* (1, 10, 4) {real, imag} */,
  {32'hbe4d4ef0, 32'h00000000} /* (1, 10, 3) {real, imag} */,
  {32'hbec7ad12, 32'h00000000} /* (1, 10, 2) {real, imag} */,
  {32'hbe8d6aec, 32'h00000000} /* (1, 10, 1) {real, imag} */,
  {32'hbe2a6256, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'h3ee8ccfa, 32'h00000000} /* (1, 9, 15) {real, imag} */,
  {32'h3e561a79, 32'h00000000} /* (1, 9, 14) {real, imag} */,
  {32'hbd31c86f, 32'h00000000} /* (1, 9, 13) {real, imag} */,
  {32'h3eba900d, 32'h00000000} /* (1, 9, 12) {real, imag} */,
  {32'h3e9211a2, 32'h00000000} /* (1, 9, 11) {real, imag} */,
  {32'h3f2fde60, 32'h00000000} /* (1, 9, 10) {real, imag} */,
  {32'h3ed8d6f8, 32'h00000000} /* (1, 9, 9) {real, imag} */,
  {32'hbc42759c, 32'h00000000} /* (1, 9, 8) {real, imag} */,
  {32'h3ec39908, 32'h00000000} /* (1, 9, 7) {real, imag} */,
  {32'h3e80b3ea, 32'h00000000} /* (1, 9, 6) {real, imag} */,
  {32'h3eb2c37d, 32'h00000000} /* (1, 9, 5) {real, imag} */,
  {32'h3ec022e2, 32'h00000000} /* (1, 9, 4) {real, imag} */,
  {32'h3eab87e5, 32'h00000000} /* (1, 9, 3) {real, imag} */,
  {32'h3daf3379, 32'h00000000} /* (1, 9, 2) {real, imag} */,
  {32'h3ea2da7a, 32'h00000000} /* (1, 9, 1) {real, imag} */,
  {32'h3edc18ed, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'h3e9ea46d, 32'h00000000} /* (1, 8, 15) {real, imag} */,
  {32'h3e9cfdeb, 32'h00000000} /* (1, 8, 14) {real, imag} */,
  {32'hbd4621fd, 32'h00000000} /* (1, 8, 13) {real, imag} */,
  {32'h3e016471, 32'h00000000} /* (1, 8, 12) {real, imag} */,
  {32'hbd276818, 32'h00000000} /* (1, 8, 11) {real, imag} */,
  {32'h3ea0adbc, 32'h00000000} /* (1, 8, 10) {real, imag} */,
  {32'h3cc45bc1, 32'h00000000} /* (1, 8, 9) {real, imag} */,
  {32'hbe8e2388, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'h3e577ee4, 32'h00000000} /* (1, 8, 7) {real, imag} */,
  {32'hbed6c777, 32'h00000000} /* (1, 8, 6) {real, imag} */,
  {32'h3e52743c, 32'h00000000} /* (1, 8, 5) {real, imag} */,
  {32'h3f23edbf, 32'h00000000} /* (1, 8, 4) {real, imag} */,
  {32'h3f0f2337, 32'h00000000} /* (1, 8, 3) {real, imag} */,
  {32'h3ea97b7e, 32'h00000000} /* (1, 8, 2) {real, imag} */,
  {32'h3dfe1d22, 32'h00000000} /* (1, 8, 1) {real, imag} */,
  {32'h3ee0e79b, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hbceb821c, 32'h00000000} /* (1, 7, 15) {real, imag} */,
  {32'hbd13cb59, 32'h00000000} /* (1, 7, 14) {real, imag} */,
  {32'h3e0e4070, 32'h00000000} /* (1, 7, 13) {real, imag} */,
  {32'h3e2d7945, 32'h00000000} /* (1, 7, 12) {real, imag} */,
  {32'hbdb62296, 32'h00000000} /* (1, 7, 11) {real, imag} */,
  {32'hbe40df52, 32'h00000000} /* (1, 7, 10) {real, imag} */,
  {32'hbed97c09, 32'h00000000} /* (1, 7, 9) {real, imag} */,
  {32'hbdadb652, 32'h00000000} /* (1, 7, 8) {real, imag} */,
  {32'h3e451463, 32'h00000000} /* (1, 7, 7) {real, imag} */,
  {32'hbf6cd7c0, 32'h00000000} /* (1, 7, 6) {real, imag} */,
  {32'hbefb65a6, 32'h00000000} /* (1, 7, 5) {real, imag} */,
  {32'h3e462db0, 32'h00000000} /* (1, 7, 4) {real, imag} */,
  {32'h3e4417fc, 32'h00000000} /* (1, 7, 3) {real, imag} */,
  {32'h3de782f4, 32'h00000000} /* (1, 7, 2) {real, imag} */,
  {32'h3f0b0c7e, 32'h00000000} /* (1, 7, 1) {real, imag} */,
  {32'h3f88bdd5, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hbce1441f, 32'h00000000} /* (1, 6, 15) {real, imag} */,
  {32'hbe6afcc0, 32'h00000000} /* (1, 6, 14) {real, imag} */,
  {32'h3e37f8d8, 32'h00000000} /* (1, 6, 13) {real, imag} */,
  {32'h3ee904cd, 32'h00000000} /* (1, 6, 12) {real, imag} */,
  {32'h3e3a07c1, 32'h00000000} /* (1, 6, 11) {real, imag} */,
  {32'h3d239fb0, 32'h00000000} /* (1, 6, 10) {real, imag} */,
  {32'hbe52a3ae, 32'h00000000} /* (1, 6, 9) {real, imag} */,
  {32'hbd38ad33, 32'h00000000} /* (1, 6, 8) {real, imag} */,
  {32'h3e83b95b, 32'h00000000} /* (1, 6, 7) {real, imag} */,
  {32'hbedff30e, 32'h00000000} /* (1, 6, 6) {real, imag} */,
  {32'hbf1d1776, 32'h00000000} /* (1, 6, 5) {real, imag} */,
  {32'h3ddd092c, 32'h00000000} /* (1, 6, 4) {real, imag} */,
  {32'hbebb67ac, 32'h00000000} /* (1, 6, 3) {real, imag} */,
  {32'hbf4a76b9, 32'h00000000} /* (1, 6, 2) {real, imag} */,
  {32'h3ecc1dda, 32'h00000000} /* (1, 6, 1) {real, imag} */,
  {32'h3f81c8db, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hbe8107ac, 32'h00000000} /* (1, 5, 15) {real, imag} */,
  {32'hbf025b46, 32'h00000000} /* (1, 5, 14) {real, imag} */,
  {32'h3e04cf5a, 32'h00000000} /* (1, 5, 13) {real, imag} */,
  {32'h3ed1203d, 32'h00000000} /* (1, 5, 12) {real, imag} */,
  {32'h3ecba304, 32'h00000000} /* (1, 5, 11) {real, imag} */,
  {32'h3d3ac230, 32'h00000000} /* (1, 5, 10) {real, imag} */,
  {32'hbefd70dc, 32'h00000000} /* (1, 5, 9) {real, imag} */,
  {32'h3df79b50, 32'h00000000} /* (1, 5, 8) {real, imag} */,
  {32'h3e6e10f2, 32'h00000000} /* (1, 5, 7) {real, imag} */,
  {32'hbd7453cd, 32'h00000000} /* (1, 5, 6) {real, imag} */,
  {32'hbeb2cc79, 32'h00000000} /* (1, 5, 5) {real, imag} */,
  {32'h3e3a7814, 32'h00000000} /* (1, 5, 4) {real, imag} */,
  {32'h3e407a00, 32'h00000000} /* (1, 5, 3) {real, imag} */,
  {32'h3e881ba2, 32'h00000000} /* (1, 5, 2) {real, imag} */,
  {32'h3f59b33a, 32'h00000000} /* (1, 5, 1) {real, imag} */,
  {32'h3f38ee34, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hbf1c1a13, 32'h00000000} /* (1, 4, 15) {real, imag} */,
  {32'hbec57fc5, 32'h00000000} /* (1, 4, 14) {real, imag} */,
  {32'h3ec576ae, 32'h00000000} /* (1, 4, 13) {real, imag} */,
  {32'h3c046126, 32'h00000000} /* (1, 4, 12) {real, imag} */,
  {32'h3dce5d87, 32'h00000000} /* (1, 4, 11) {real, imag} */,
  {32'h3e5d73b4, 32'h00000000} /* (1, 4, 10) {real, imag} */,
  {32'hbed6e80a, 32'h00000000} /* (1, 4, 9) {real, imag} */,
  {32'hbdf81c46, 32'h00000000} /* (1, 4, 8) {real, imag} */,
  {32'h3e94a555, 32'h00000000} /* (1, 4, 7) {real, imag} */,
  {32'hbe95878e, 32'h00000000} /* (1, 4, 6) {real, imag} */,
  {32'hbf0a1aa0, 32'h00000000} /* (1, 4, 5) {real, imag} */,
  {32'hbdc5e649, 32'h00000000} /* (1, 4, 4) {real, imag} */,
  {32'h3e719ea5, 32'h00000000} /* (1, 4, 3) {real, imag} */,
  {32'h3f171ca1, 32'h00000000} /* (1, 4, 2) {real, imag} */,
  {32'h3f263297, 32'h00000000} /* (1, 4, 1) {real, imag} */,
  {32'h3ea25634, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hbe4e586d, 32'h00000000} /* (1, 3, 15) {real, imag} */,
  {32'h3e9cfebe, 32'h00000000} /* (1, 3, 14) {real, imag} */,
  {32'h3effbdf6, 32'h00000000} /* (1, 3, 13) {real, imag} */,
  {32'h3da033da, 32'h00000000} /* (1, 3, 12) {real, imag} */,
  {32'h3eeb6e17, 32'h00000000} /* (1, 3, 11) {real, imag} */,
  {32'h3e9153d3, 32'h00000000} /* (1, 3, 10) {real, imag} */,
  {32'h3e737ea8, 32'h00000000} /* (1, 3, 9) {real, imag} */,
  {32'h3d5f8e5c, 32'h00000000} /* (1, 3, 8) {real, imag} */,
  {32'h3e3c6c07, 32'h00000000} /* (1, 3, 7) {real, imag} */,
  {32'hbf2f3f1d, 32'h00000000} /* (1, 3, 6) {real, imag} */,
  {32'hbf9d3f2c, 32'h00000000} /* (1, 3, 5) {real, imag} */,
  {32'hbecb4ada, 32'h00000000} /* (1, 3, 4) {real, imag} */,
  {32'hbd946ff6, 32'h00000000} /* (1, 3, 3) {real, imag} */,
  {32'h3d80868e, 32'h00000000} /* (1, 3, 2) {real, imag} */,
  {32'hbe1e50fc, 32'h00000000} /* (1, 3, 1) {real, imag} */,
  {32'h3e083ea8, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hbe9653db, 32'h00000000} /* (1, 2, 15) {real, imag} */,
  {32'hbe0ce49a, 32'h00000000} /* (1, 2, 14) {real, imag} */,
  {32'h3cadf150, 32'h00000000} /* (1, 2, 13) {real, imag} */,
  {32'h3e1cbc78, 32'h00000000} /* (1, 2, 12) {real, imag} */,
  {32'h3f1ebfee, 32'h00000000} /* (1, 2, 11) {real, imag} */,
  {32'h3e3208ca, 32'h00000000} /* (1, 2, 10) {real, imag} */,
  {32'h3d3f30b8, 32'h00000000} /* (1, 2, 9) {real, imag} */,
  {32'h3e6326e6, 32'h00000000} /* (1, 2, 8) {real, imag} */,
  {32'h3f1a6517, 32'h00000000} /* (1, 2, 7) {real, imag} */,
  {32'h39c18419, 32'h00000000} /* (1, 2, 6) {real, imag} */,
  {32'hbdd5a12b, 32'h00000000} /* (1, 2, 5) {real, imag} */,
  {32'h3ddb1a62, 32'h00000000} /* (1, 2, 4) {real, imag} */,
  {32'hbcf5c324, 32'h00000000} /* (1, 2, 3) {real, imag} */,
  {32'hbef9d9a3, 32'h00000000} /* (1, 2, 2) {real, imag} */,
  {32'hbf078b15, 32'h00000000} /* (1, 2, 1) {real, imag} */,
  {32'h3e0b2aad, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hbedcf3bc, 32'h00000000} /* (1, 1, 15) {real, imag} */,
  {32'hbf3fcbb5, 32'h00000000} /* (1, 1, 14) {real, imag} */,
  {32'hbd92592f, 32'h00000000} /* (1, 1, 13) {real, imag} */,
  {32'h3efcaf66, 32'h00000000} /* (1, 1, 12) {real, imag} */,
  {32'h3e8e5543, 32'h00000000} /* (1, 1, 11) {real, imag} */,
  {32'hbe42a9f5, 32'h00000000} /* (1, 1, 10) {real, imag} */,
  {32'hbe209d76, 32'h00000000} /* (1, 1, 9) {real, imag} */,
  {32'h3e22037f, 32'h00000000} /* (1, 1, 8) {real, imag} */,
  {32'h3ec7804f, 32'h00000000} /* (1, 1, 7) {real, imag} */,
  {32'h3ef4a136, 32'h00000000} /* (1, 1, 6) {real, imag} */,
  {32'h3f2e8d01, 32'h00000000} /* (1, 1, 5) {real, imag} */,
  {32'h3dcd933f, 32'h00000000} /* (1, 1, 4) {real, imag} */,
  {32'hbe4d632f, 32'h00000000} /* (1, 1, 3) {real, imag} */,
  {32'hbeb57b94, 32'h00000000} /* (1, 1, 2) {real, imag} */,
  {32'h3e84c88d, 32'h00000000} /* (1, 1, 1) {real, imag} */,
  {32'h3e45c80b, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hbd8262f0, 32'h00000000} /* (1, 0, 15) {real, imag} */,
  {32'hbddbd8f5, 32'h00000000} /* (1, 0, 14) {real, imag} */,
  {32'h3c027134, 32'h00000000} /* (1, 0, 13) {real, imag} */,
  {32'h3eb867f9, 32'h00000000} /* (1, 0, 12) {real, imag} */,
  {32'h3e07c629, 32'h00000000} /* (1, 0, 11) {real, imag} */,
  {32'hbe87a56c, 32'h00000000} /* (1, 0, 10) {real, imag} */,
  {32'hbea79af3, 32'h00000000} /* (1, 0, 9) {real, imag} */,
  {32'hbe0c852e, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'h3de7ff54, 32'h00000000} /* (1, 0, 7) {real, imag} */,
  {32'h3e839aed, 32'h00000000} /* (1, 0, 6) {real, imag} */,
  {32'h3d9b5b37, 32'h00000000} /* (1, 0, 5) {real, imag} */,
  {32'hbe1e1001, 32'h00000000} /* (1, 0, 4) {real, imag} */,
  {32'hbe721540, 32'h00000000} /* (1, 0, 3) {real, imag} */,
  {32'hbd5f8d6e, 32'h00000000} /* (1, 0, 2) {real, imag} */,
  {32'h3e0d23e3, 32'h00000000} /* (1, 0, 1) {real, imag} */,
  {32'hbd8b74f7, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'h3e3c6c46, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'h3d6d18d9, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hbdfb0e81, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'h3d979be5, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'h3e2670a3, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hbe7070c0, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'hbee899f5, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'hbce63286, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'h3dd43aa8, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'h3dd44049, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'hbd8d7d73, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'hbdbf4f0b, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'hbd742ff8, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'hbc295098, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'h3d9a9a58, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'hbd118633, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h3eadfdea, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'h3da541be, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hbe76c552, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'h3daf84ba, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'h3f234303, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'hba1d54f2, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'hbe982bf4, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'hbc6b7f8d, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'hbd158a38, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'h3e81aeaa, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'h3d7c90fe, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'hbd0992f5, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'hbe06c785, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'hbc48e6c9, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'h3eb80a80, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'h3e5e66a5, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h3d23018c, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'h3e1d702e, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'h3c79ce02, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'h3e9ab4af, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'h3ede5c90, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'h3cdcea52, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'hbd73bee4, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'hbcc72db4, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'hbe1608e7, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'hbcbbb971, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'h3d352869, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'hbd9cbb8a, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'h3d8d3af1, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'h3e8a4f32, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h3eee388f, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h3e914c29, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'hbdef9a9f, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'h3da9a9e8, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'h3e87fcdf, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'h3e58ed22, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'h3dbd148f, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'hbe858b49, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'hbee4c2c8, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'hbf379348, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'hbeee0a7b, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'hbe96f5b8, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'hbe1fa6e2, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'hbe02ee71, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'h3ed55518, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'h3f100c74, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h3f176704, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h3e9cac54, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'hbd9213e3, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'h3db4e277, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'h3e079299, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'hbc71304e, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'hbba2d8bb, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'h3d9f02d8, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'h3e14d94b, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'h3c9a8fca, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'h3cec8a11, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'h3c412521, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'hbd58cc0d, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'hba84307d, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'hbdf4d51b, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'hbe1e9f08, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h3e5a8227, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h3da91dab, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'hbc83e331, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'h3df663de, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'hbc7d1a5f, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'h3d990dc5, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'h3e7ce05e, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'h3e91b2de, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'h3ed16a85, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'h3e1c8b0a, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'h3d249b6d, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'h3d7f5314, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'hbeb9cd1f, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'hbd4734a0, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'h3abb51f1, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'hbe83bdd6, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'hbe1ea16a, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'hbd9bc15e, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'h3d820fcf, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'hbe8626a8, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'hbeac1cc8, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'h3ddc2ba8, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h3e846a08, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'h3ee4e726, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'h3d9c921b, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hbec5d207, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'h3c6e87d2, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'h3f049419, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'h3dcb2d6b, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'h3e1d9839, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'h3e5c6700, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'h3e53a5ee, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'h3ea0dbc2, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'h3ea301d9, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'h3d9f883a, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'hbd8fc538, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'hbeb464f3, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'h3b78184c, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'hbd2f3b37, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'h3e4a2a58, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hbe2f4373, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hbf020e0d, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hbe69da96, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hbe599214, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'hbc18f100, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'h3db23741, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'h3e938366, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'h3ef6c13d, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'h3e8b80dc, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'h3e8f8504, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h3cbf10f1, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'hbd3882ac, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'hbe3cfd43, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'hbd8f8b7a, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'hbe164680, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'h3e4942d8, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'h3d95a18e, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'hbe1fca1d, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'hbde0ff58, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hbec4e236, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hbe95145b, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'h3d95f0ea, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'h3e3dc651, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'h3e323506, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'h3e8e6aab, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'h3ed6623f, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hbc066c73, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'hbe86e6bb, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'hbe588e42, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'h3d5f09a6, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'h3b75e070, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'h3e66d20a, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'h3db831b1, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'hbdf6a1a2, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'hbcd64549, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'hbdd7655c, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'hbe846322, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'hbd8cbd20, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hbed6619e, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hbf179f9a, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'h3e11fcfc, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'h3ed67479, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hbccd2b4b, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'hbe7c5717, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'hbd98b880, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'h3e30d61f, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'h3e73a7d6, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'h3e56a60d, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'hbd3e53f4, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'h3e3c6af0, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'h3e09bb01, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'h3ea1bb4f, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'h3c5dea77, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'h3cedf16d, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hbcdb53aa, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'h3e419995, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'h3ea35cd4, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'h3e3e840b, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hbbbebefa, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h3dc72a84, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h3e36708d, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'h3d2e2b9b, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'hbde4a78f, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'h3e00db00, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'hbcd9a5e5, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h3dc65906, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'h3e2baaf7, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'hbcbeb45a, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'hbe4098d5, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'hbdf9a0b4, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'h3d295324, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'h3e8bdd34, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'h3d7387c3, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'hbdbafd4d, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hbc5ce727, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'h3eb93e90, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h3ee7220a, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'hbcecfc19, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h3df8e8cc, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'h3cfa7508, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'h3e564548, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h3e92b886, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h3f042f90, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'hbe2de2f1, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hbec4538d, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'h3da15f5f, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'hbceb932a, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hbe478e13, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hbefed79a, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'hbe8466ac, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hbe5ce018, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'hbd864a0e, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h3e827fd7, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'hbd63558e, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h3eac847b, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'h3e86c0ee, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'h3ebbb502, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'h3ebdb534, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h3eecd64a, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'hbe87ef26, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'h3e977264, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'h3f249028, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'h3d394446, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hbec2237a, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hbee065b0, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'hbd4059d6, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hbebf48f9, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'hbeeb5e12, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h3d2d4d87, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h3e97a2cb, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'h3a78f988, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'hbe3e1387, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'h3e51c3d1, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'h3e34a9e0, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'h3e1470d3, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'h3e158fe4, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'h3eeae4ec, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'h3e98e53b, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hbd120adb, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hbe823a80, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'h3ddcbbba, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'h3e08c215, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hbe65cb63, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'hbe09430a, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'h3c50155b, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h3e9f2f28, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h3d21d3e2, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'hbea35f77, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'hbed15f63, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'hbde9e484, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h3cf3d977, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'h3d894ab7, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h3d9799d7, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'h3d0c1dc3, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'h3d964894, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'h3d9d2168, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'h3d9aeaff, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'h3820d31b, 32'h00000000} /* (0, 0, 0) {real, imag} */};
