-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
zMy8+Q1nhWWlo6TmpjcIFMEhh6m7eJ1sd1+USfY269rbIA1uPtdIJVNrim6/O7q7
7CF7wTWXWlOMfz9OyZBmnRqZyQoWsH8WMigxdwrxqCKixQa6TB78hff6ujhfkc2I
YdPiqH832Rs3Kt9+vVdLEHRLiVKKzDItBCxR2lUsxX4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 20112)
`protect data_block
jKjtXNmZc2NgAw4PcmuF6XVM0JtWXv52/WPkDDgt2NSGzpQZ0iSPkxwE/21PcFDp
Y71wOGcKKfUjPH2+HPFBPQ5njQRE3/XmmhOf5T6ynMhmAeISNzYSpTpG1CiSpUlf
0HjLMK1lh9xdLv3ip3pvzbSwA/M7bzzc2Ys/Q6Pd9ttHm6M1bCTSG/f380X+RHbd
vGCU04Mm5k6snKCFQ1oJ28hQa6Sa0JtH3WCH5fDzAF3MGfcxmgJvUoLsvmAlDlK1
FcUv3e8A4z9R5j1SyJmLQCnjFwrMaciaQpUb6Qj3jHsUHsfS/EyCYFXKIrO30R+Q
K03vY5Q5k139S7tUl0i1oyS7EoP1JGWL14UPjSdk+PAuz+ETPBtqNpiLM42pqN2b
Hi7sqACAYUC3mVnaZw53ep1CHBLmo8VUptBgk5gG+t2R4Jp7L6H2dpoUSSAIK6iJ
17kFzCYnL/tx0NgLkm7VQMUHAWQddZ2oc1zSHUO4CnxsWhE4XH5iDubWWloU+mdB
9zoQcCXLbdodoPjc99nABAH2ZZVcVSeg2i3I/TVI8/sdkgg7pbgIZcv4tuFAQnr6
ov9A1lcwy3i5h8ZYwYz67hvJTo3mH2bb8SHiXJdC423p0kcCHBHamQA7fpVRVyPO
AV13lLshpO9zQuTLkHyL6difxlxCT7LxuMmHQztPCWc2ZBxiB3ZLnPVSoZA4OUxn
2z9Nq/XSwiwoy5vrNDEk132yuxaRxhNk3PVTzWMTiEf3ZPkVBfV2WcLV1kHFu5O+
oQWD2vu62kjOgzErJDwPINMbHrElVco98G4rJOPn8o5h5xMcCKsPRx5+5VIwGMxn
4sjBMd3K/bVPH7L83Zb/osuS0WwIXUmAg6VbMSv4q1pNtg6Llee4esM+SsWjA+id
Kjzj75Pi0QcrITKFIPnFwv6xEIoiRgf/qt88sm8XYzUnnLan3EK9p20QAuOkzI8h
dFkWREReI/cNWUHB4g+yw0jlcdbY2jyNqluE6ioHoTsgS9VINHmHlmqL6VWAi2lz
87/sPM4vJVoPlZow1v0QlPUd/Cvi9nwyzDBx7VJgexQ2+AbSggwTrDVmh+hItCC9
OZX8By/VQyoHP2ND6GV2LNQ+PutHX7wFjTSQ4QUCiwxiZV1dvxngfvIZZcDaS1bl
ls7hxQJUITKOGG4LYxc19djYnnUoQonUvu0Cq3dvzlfSfS4mHpmYuYzqbAwgZUH+
g/m/YryyCh3JzpWo1MbMAlFS1OicuqZDNkXqtPDZPglY61KbFeaky1iswmlMkjDu
7wApPUti+RBok1WM/TxFHXCbXLNwEFwe97xnk6cgzGFGci73NVzQ8FwS/qbL0zJH
FwGKofyh2INikVByfROuFRGF/6tEICDA1BrY+/9m5C7P/jS3D9Kjd7Cf8okad7Ut
HowtLqFlouXNyhoR30GRo3sfPcC21PHcWCo6j3BzzVxucv4Lt6y7HJRFhoDymW+5
pe4NZaP8+y0klue8wCB2T/svzKXBUWYzroDZmS42mMk4QYVNwribSfAv/ugdDRjy
E2A2LhCEU2bzOEdoVsnvwWoV3H3JfgM24E8giAFJEj0JE+pPrNfkH/S+yYoRx4WT
veLxPe1bE/AEcfWmpWhPdgyyzKF7Iipj3aIeT2VD35d5TcR5Dh6E2PGS5LOIrcMT
Ta6YEENMNNW0NwKiQlGkZLinwsAVK9QeKf2o9d+zfWEML7kKqxoy1pyYHM0lgbmC
td0s+/j6jBcRIyyRqCCnzJ6nasdjWgRJBLMY5dJZvVQ+0QIaIJBPGqX1ltK6hQ4s
3pnxBtkZyhpYVenSzgFQ8qXDIWHkSRWYQ4Y0begE42xZiW1kg/MleWoGBHbyyLu5
rUdxaeb4qsRqcHbj/INCj9LzOZtzf62U46KFKEk726KxI7uFLJ4WEw3DUNrHlnc1
ZWd6McQyLOBHT9KgxnSIPhYLgwYg1jHDYq5Uaw4/y3NOYQQ+X1xP70n3EBtI9shI
gascrthxWNdD8/BKW++M/NFhw3D+/COxiRRkRaTXt/iBqkTy4Y1bVtQpamLdwSk+
9qUSYux09hiI0Q9RQHyt7U5/DbOWgx6j/c9QuTHuhHQI/rsoulgBMGoViwT4Ou83
ZzV5yltUhzZ4JBiS/mfsgfVXhHh9FY2fjodyGc3xFFqYQi+qoDnFHe5jP4sXYo4a
OC7NeyPEvQ2N5WzU6Smg8lIt7yXlyAPRVXK9kkzfikzC0VoabK5uz1JXWBNsWeuN
jhb1AAnn+0s6o3jgY5DZtVUzWWE6uLOdpTubLSfVqPnFzLH480vEXXmDOmPd4tCg
N0NtA/JGoYFiT+gtHI0zFKRx4Z4Uf32ywI+0sZcmfy6Xg+kqodQg+54JZQpvZbB2
HwhseRSVOPi2V1v8qZJb7TzjAZi7ZuW1ew3+caspjt3Yd81NyUe0EdlepB60595f
hJKK+yXxIy1kYtlxCtgPIE9tCvPhtFiaPR0QaIT1D/4oxwHGUfyu8MvJv+HLd8PD
nXtwfIjlzby09KlOIL5tNGHspwaHUzvJsODraSPB+CTMRd74sbvH1XZfrdeuCna9
yS8wlKnPdsHzp1iepOcGmeT1ijpObSL4gqRBjCTMwqKM55NBtFDqFzKphjSZXqXi
q4DiHqZww23Jao2mJRQfyQ5R1/20IvfvW80zp4f5qDPq4bkF/FUvr3fmCsvAZ5Bm
Rw8JWZBZEtRd4TdPUvUDnPmJ1nxpVMyoyv2FbWaQMAAF6A5Qc/RjYgt8zpinmPGD
rc/bVHMWeHy8iEyAo4Btvqar0yPhp2kIolxWO8zfgUgkOw/EP6/1NLabWIgPUTl7
28sFDd0aBD8V6AEkez+Q5XCabXLlbQH9dtBZcDPnKWBuoB7KNfvAqD/h8XRNBP2P
bdpzKvASeIYGPPvUjgKTzUdczjsHj631AO27KoRGUB09Uhgj+g6nxUa2ZA+MVgiG
Qp9Yd5WA2EbJUp+95p85XOH7Ax8YS+lxsqMlYENCxtFRlAT7crQG1KxLgaWRWASh
1ni69fkIC0WGX26q1oPvjM5qEINZtwPvep3RdxGrLvzwvddxeTiGu6w4uD+fqw0r
1H9/7RLVSwWRFOUI77x6eVOMVKMaRox2Pxzb6/5CS1GrohmcteBsD303mAUS7tfF
+vmrDwQ35x3FcFF/NDKs7OBxnFDjw7KeF26JEa2WbA+tMHhwUsR6t1bf6ObZrl8o
1tLgoOZB4zFFzRjrBqNQctYltadpT7KoRIKaOnRiUfX/UozIoqng+xyPAfA+SjV7
QM4Vd1AplhSaWL09gBF8dndU2xnRP34fGZNOWE0hK4LoNKjkQqSRVVdtD1eusM7F
hfTHibtUzEO/adWlVxbpGFFQCTpFFbRFnbFDH0/Nly+PBvxNnAZzCRT7XYd8RSIf
mky1/uKw3EQm3QmURMV1O9+3pe+6k9AcwHEfgTWfH9kjKe1rzMa4oelrCkcXUg2S
yEtg0EdZgpfZ0S/FZQVwk3BqIuRa4TIe/9bDtRYy0H9yydOGnaAxxb7wu345CQ5B
EDeHEIYjQNq1Mwiobv+RMcfD4nipB3WK0a5zeXOJLI4VIQRKKlDE4l7KMAWgvw4N
mu/UkGhJ19QQG5etoiShnb/7u8YCL0r2O0XkvZCUHAQL+jyJ8MRZBZputkWeqJsO
BNwtwYtkfbJTuwSQ4YUzlvdL2ceQlEptGmW38FgC8sWM1TJz0MPLC8see3L/IzbW
WWWt5t7rU+/4BrSa67sLPbM5vIhg3YFyZgqu+a3WatI9ngrQfs+g0G1AOC4rkSKM
UQdLjIMN1e65VfW3crLN0hshayzdljAnNY/ZInW9yJ4LWkq4ajUXpKQDzXqpN0lA
+7NuCLase3SWnip+rV2CwnTiyLbfvdkPnF5dV2sxzckmtJZcbanfQwkq38acJyT7
GM2r1oWzawKdzk8efKUOLZ8kbClpT7FXSgIWrJrbjfMRvFliYea7gJ6yskQn83bN
/XI3CqkWfmdQ1z7ZFMPDX/+TsIYK4lCuXcSlgdwV8xrbnwCq3Nw9BQCCnmvQKGJI
UEQvtU6PxxymPxREDMhVRhr/CqhHTZ3az+ajs0lw8W9yzGkHPjSPo72nfkjazmHK
36y6sL0uGWteUno78afbHCWdIE/nYI/K2o5l3ENmGSr40/hAZxYud/c/7SSHDATc
/SstAmTywkFsFNxDTlnMAktutF5kM2DHetzPrPj3vMsGlhuDI7mQjyc3yfXzSQa9
NcGMOEfPXye+s2Isq9cjywBuhteiyZp9UBros7HsocUIHoo31XT8ekF9FCCWEzyV
xSFqNg5BQQyXjrSM2U647W85JtOqmoXVq4gGeMRC0jraCULAvhoPeFSkizYuukJm
JAIgpWCNO6GBsCAOyceqtnncyeM2s3beX4rFXHMevS6Vnasvg8eF7u6ev6DwBDJe
x6yolxsaNp4OrUaGFddt6aETyuEAjGY2g3ojQzvPUfpqR+EoOfKWjl7LwQBUTMRi
Nkb8sHfH/g/WGZPLCUjRkSuPbdAgbkyKQ9Or8hEySlExPIT9OCJ6L27uSmmYZS23
ubgoFwQ+T1BddF/Fg9QYNBVbwxQ55Y29FuJ1plrY9JU1gQyTKLrMxKB/Ty2oSKIR
tQzQZ7XKPuhHIja3/2CSkAra2pXFUxGh5BYPDqhwpD+Mk92VexXb4NVb9Kcq8tKl
DD0wRCe8lTen9+Cqs8KBWIcBRTEk1FcIXGxSs5yYQD+iH/7Aj62zOIMsWRttnTGi
3anFP5ghCUqyzhYwIMthhh023KHMdBydKxqXTkwy7mzBLkJA4tn/ALVN0z3sJazw
O4yMTDM+rHSWpyPyjIfGU/kEL2svZbTUAseFciz7Gc8HYj1WpGFTGacmy3uwAZ1T
bIFKm1sKPV7Z3QkVXAviQA25dZZSdY0XEk9bUd1Lx/eWV3NcF/nnAzI5aZagqF2k
/OaNyawVs7n1I9v61WDCYvdqApJQaKp9xjovWME03T+fP+9jsz02DmekDzJZ/loV
062GH1oBbf7x8atvBSfhwn3805uiLTG3HPDsrqcrgaAfSGgHrN6DfXXDcrv3iZSZ
xdkvsRtHGiU2l+40LWM8LR9B+yQFvMC9am+H+sCM+pcG/d6ohCzOksqw4UOS1FPq
lYKq6o2K9U59F19SfEbMVYEf5Zb3dwB1r4BmDty7jvX4jzLaqVlLMohH9YGrDpaT
GfATabQCTXF8IJ0Y2tGcF93J9540pKT7/oIUJjaN352oeY7DM1ND5W8lHb8KH2Pe
vRDW1X43ITceZ/O4mtciFzu/ok7hTdmIb1w8iX3bXL3Gp2J/3uCOIaGqymlsW6IY
RikwDx+mvxOpHfPnTkiwLqDjvYYFm0AV3QT8HgDnZPYin3Lt0KIsdQGLZfTRJqDK
3Hwfk72oO0TcmrxCn1x24dvkHF+/cp6LcGsGGYf2wBR6wtuaMPgcPuD1zCET0aX1
ZdaUA+76CQOj3+FtDhlzE6wAv7m9iFAmMWdtwpyM4yy+pCrP/Cs7fDxqIRUJS8I9
heyGkXIvsF3guNzvUcL3VLMIlweAiCiex5Kc4XlRj9UMbloU99vgb0N9r3W3pk4v
ds0eNQp7P4frgW1PAo9BC6p7lPGIR0TjFyoWnIW4dO3M9d1G8jn2MtKWXTnampHG
NzoOjX6/996cLXJjTFopDoxc4pQbNlXJ4g31k0xH+JJowhGPgEAtfejjghUq0oEZ
lSdljh4VSJHI0OhL8w6Emje7dIkvA75KT0jqHZEv1Jvpyy/CnjmCHQ2JYDH44q1w
+Pc7YLiXp24WiLRSYlDT6zPmLaJa9jkofn2rp3dOdPXVaSZV5FzxP7Zhp8sWuMdZ
fTHCCwx/DI+DiLcBqhP5cXPQzxNxMzypFpCLZovuA4Ch7xeiv4bpwesRdLV7lh5k
5dPSc0HiZXk52QppSY5rAaFkCZzoI6u8J4Dv3WBxNXUzjauj0jmDG0ReYREvQp2b
3UHW6Vo2v4XJ9+i/xo5lkEdDytZYBUVxNlalh53coOi0BU3a73pZ2I3oO3MS7Ys8
JpTTric5wP2b567ZPnuC7ZBj9OXBQPk4HGcjzvdD8edxiC9yo691aYEltlI63Xkg
cichJFQzgURQAf4wABwPxLdP2kZ14RZzFeu5ptG9OAnJXjq93I1Sq6Jm1lh+IweP
Gkd1xXy3p+8E2JIM34uwPhQzn4WM1F9q0AXx9k/DzVptVpePO+dvhW5W8RbRRLTY
Fk6oi30I0SPqe7KUXwg0sYR6eugXThnUXBY08bB/BP7aCjierc5wca7xuivu/5NL
MeqaXFuR3GP8oTKOS7qOI1/cpu/s9SZsAKbSR5IK7G2uHWGMzuSpJfDHOKegg/zk
MBIICdW44o7cW6QbbDoI1o9vVEwyKykfeUnJ9TUnRnBNDv0NDFaWraaCEQVWOwCi
VM2meb5rWfzR+sxi4822Qw+rPluFfjDbSpV0AbtgU68xrgk2cJDjkuyEJaicVLcY
hbv3dwN1ldz9CkqpqwLRUmSV90beruKZ7kA2xx/oN277Zt5uoQp259JEllKz+3CJ
tDj4P2ahqmpjipPP2IDcKsh6zKu4+4QPhVwEggjFruuS4GNry2S4QRF3o2MuEURq
JFh7HuAQq+0PIXmYCTZyKylQe0MiQSF3deH2eBMcIdx8ed1zbH4ata3HwMVE4oXL
DRAFGE01tdOLr57ueG6OvpVJ3DR4R7mRtSSl05WPhSACflYPvizrfyK0QQPb0r4v
GkdYspz/1Mok1M6dXi67yTVpomkcXTtcx5cOwqU57e2w5HvFE+2tara2ZIM/rUIq
IBPYXROPNzgEoJxpHtmpqnA1AhaUqWqFjjXqtgZ5vxKvpD9lWitB5arHnxVLa7v6
K4Nxft84ViS+pJ6pm2aT6iWd7t53HrnLdOMEGoJ1pbIQ5Nq8U2Kyoik46BtfH/va
VVa/beRJ43pSBnj+BA4sommBWKwmxyX1ZsmGFOAAgrRqH+dkRb+voMPOQotfpMIU
uZ6YTyZkWhrpZJ8XectLrv/t/wDAe4xnU/QY8FaNsL/wLXoHwsGElhTbFCs+mHHw
GEmyBWo+q6vpoVZ0Xs4GI6Z2xuca9psUynzl50EhwJmoVbHHJ55c8wG512H/xqAY
9KNSrMaaYWDbtfxNjlQnpsoKxuMTFF3PzyPq2QOjRh3koSZmmvfEyi7axqkVJPDd
5G2bkgCJjGgHHXun7rCdIDgGEWKHej5cepYS4bZIyGcrrB6IOCzTrR8Yj6ISXCsn
Xg9okVWStw/4c3/2Ur5CWQI6xIuJQj7vXzz7iQfjFrn7hRKNuvmbrlRM9m63DMCG
F1gCfAfH6Cdv+DsxuP48TzLcnLQfp8Rr7k+6IAYZede1ngV9XcwYkb+K9CsUX42y
VjReg9PFoYDjR3TUDTEzHINZXn4p86fXOZeRGJVXBjpheqB7eWS3XgELDY80yMp5
Ud5nsQ8k9M9hnwSA7egqazGIp+imdhvDpljBX3I7QTxWWISrdRlqBUy6+Skv8QyD
XFQn891c9LIm9nvR0RfrOujTtf8YBrMAckBwC/WxP1trOGNBakRtpaZNiROaRHTi
kvqs1HmKDFcYFuyHUBgoVZOi/o9rZqKRQvIbiOCgx1BngIioGxga+G9nX0L5kRzn
Zx5CKPLZKBY2PBM+rXP5jnnHU3st0Ald+IpsM8SvIsHqzM1q7uI9aKiMZtmTJea+
lWXd9fvHaNmgNldDHADsYNjh9ARNUF85CgDZbE2KHAEgRuGFOTiuzURj1OMW8Svd
SGnXIxt/EXfHuDHJYNdyfEf8sRneeNLvW6nnifZmQ/TPIcQ/EUqfwtodxUkK7ogD
AFgrbWVfNUMWXW2GPU6/ui373ZUF9MmfLhwUPbM91coftVHB4O9i2lw58Ddg72Xh
9IN9NLW/1h56197HrKygErE0JZVFblJV3REOZ2n7hGTBgu4wOadRDwrBIlXoipXs
LgeTxx42bB2issHltwoqMaAg6h8w8oM5pFLVZ3AnDkiWyebaSXoxH6n+ipuPAbHy
GxbDC69Bn0k6nTl3zlDDUu80MFphBSkuslnzogvJyoeStelVmvpmp3uSgudAkvlE
m6I69v6enzg1/mCu9mibrbnEtmKmj9/K3x/acmdHrqYLCdk0fnQvVTS3QNp9sBt5
i/OMoE0vZNzBF0wsKwgYSd1MyO2F+oMb64mM1fTTSrCpwAqo8f8sPUigx2gTpe/C
tXZhfF69/DoMYgbsMxY07kCgLrm4b4frAQ0MPtKyGIT7cWn2LmJXN56f6Wjf8FtT
BY24SSzz6wqgvtCACB84NhnubqlxBFyIomEQ8ec9yEVJcXWEx8atVYioAk6Df3ub
TZuOmU8UR+dP7iWmSu6iZsPdcvpT1VsBRnGyFDrzETnhu9hrtI03MER0pfxloBHq
P3qu3baZT62KZErhCl2/Dnh308KEAaoL8/UFUvK5O/xc3sht5xF5vNwl6Dj4AKpj
XLo4CrKVizbrPrxJ8OCd+qT/HnGHzg8UWZeEICcRcxsrDvLleo8iPKYSHGKzPan9
AYjajXc3KQsNxxsMLsQX3+nIFvPuSre1UfQ6Erud7jr8q7whrSoBBjj2BCNSb805
Yj4A1KcsXwFPWMkYQCKqsjnEedurDF/FNnvqFtGl+9QXt2kFbFElTexhWYPA9eA/
1y2cycEn9CoUBfpeAazgZck1MVENFdbh+6uSgjI2ENhEG6V81C/MnMiWHQ4p+7gk
9221AeVfxqtBDQToYsefts9VmW41s0Oc9YMRq4xcJ5ZuF7q3PATD0h+FxXzcZXWo
5xpPhTsr1iH8aNhTs8o0A9iRnp5l5ptHf3RGPr1Y4OKWK/SNMmDc9WVVlET9CPMU
RWdo4E1hLdT1BlTJOQ053m9kIpedMzbTxT/5OP6jIaLjdsf6grRb/RLN+ngTCd/o
LPyjpooRuvq97c4ULDroALTmVSERrPjPDgRxIjlQ05+8A9ueOWFVwBpG8woFhJLi
77irG1MpBghe10wOKbW4jo/GOdNm0OXCMQAUTk/QOapJODQpej5EzkzDMRSixfD2
t9ZMrpanrOs/tzNreyQT4YdFNeer4HpzkWck+TeEOqSXSPKKOKiszhDZ5bnirXHR
Nd6f6NSA6fZEozsf1v+cd42NXkrmud4Euf9MuvcpuBVj7aLyN1mG9Mdt8j/fMZOO
NvKmd6M7pHPNO6/JgwtHGM35HiE0BfR4l8e69AjA3N4axaWOZwyKor9dEUhpRbQZ
8v29ip1FgVPLHxNsneG5s4EBACXYhoTlxjKkXDfcrt21zS2z0YDfbZLwks5XclsZ
ede9Bkk+bPW+sOIb/7VY4PYvysDj6hCZfDuKoFe6SIwl3l1s4v4rYA2WSvBulOsk
ir1IL3xOGPWFwMrGY/QNC/ewwuMr3vM2al3XQnaNyjg4KcVqKpiCcNCyzY91jZAK
OGlxNxR+KyxeHKrpqwggtvwDT9DqUziUMZFzk0qLmAaMmGIh+K5N8OWulBpwGxw1
fjBIny80Er+/GHRjo3mbI4sgUM61bEs4ixK9sURLyUmIMDA0p0VLGlHW6Md95rM0
ioeS1kgEb4cMcQ0i/paJ9KVvrphxxe/mABk2Drp+WaGqfjkCvfZZ+yVQC+asb0ih
G6llxxkJMX16sp9H9gbQfbF+uRgfcCQvhaYuTnBt/YMmrfGtrbngqSjK8uMn2lHt
dHhZcqajAqvFmtpevWqONB88o6NMxZ8++piqLD1AKdNUOPlX7+eHHsW+FKdFvQI/
GiiyE1DsKnCrx6O0Rw3sVAOYmcw8ea4XLFXQ9MMM8tvkhAXga0g+r4w8hHA2rHwR
wMZR+O6B0Et/4+NmK/0zdsOV0CDmp3shhcU5/oqP7sC5jAatfuWoEmYVpLKGxTPk
LPXXMJXZ+GVrcKc1k9uderILh/9XM8eZLar0R3/k5PSR4uJNtJcFd3dGcCPucahM
DJPo55pgVGZHXs9ic9GCbWXoRbJzaXTKZaGeWeY8kItjjDNeCIdJ3li3owd0g8Ol
hLlV3r8Q7cy/bZsWP7K/CKDkS8XxqBvmnXCPo6cY/FyUY/p01EVBcpoiqrBvvIFJ
/5Cp6mu8w3k1WonSs3MwkI/WFM68e1SIufcNJbxTPs4Y0IeQHLjUkYViUSDkivHq
chZe/x3Wfb1uL+S67aEeu4jhnSJkMqm7dCHjqajXudnQc3x9uuMiP2rYTib+K5xX
MgiO817Ha6Kr2flCgtbW7iq+LfO7jBrIc4uOvPaE94+eDiZO5S7U+5pnufcP/6sH
7ymLZW0qJUW23P4TMkOjsZSFJYReMGugHPswp44EtfPR8A5CgR3HVo78UNfuZtis
1vBUd744sEYkB3YvmJ8xT6u8ofp2zcx+ERMNzGD9Oyjlt/vhER4RXtWrPcSHRPRt
epL7iuW16+IEN6BgdytAuwvcyG4v97RsU6zSnyvySHrUOwhd6DpnBmPRM/AOxyLY
EY0dcYIg4IYZFtqInjNaZOmRuGYVz+odfsfysg5rmoMqobmXjAtAsfnlMQGE98Pl
H5VisQmd/HYXxGTTEU2hLT4Lwjd+9GvW6ZqcnFtXxATNp1/Y8GMCstgZLWdg2O+o
K7/ORuMEnnOBjWFQ6fhL5WxDnxJkzmjSaHpMr2K7+PFedj88Dz8C6JhrHv4Ed/AJ
19b0QObgypdaT871/ZcFyYdQYS9LC9ZEGHIqdXavFKIlUB2TZ0Tc66aCBuL26zGa
GqGAHcfKXePM2PpAQWfqnAaeg0XhLvK6e5MxjTXcMnLMwGpGonJ82Krph/F6x1ji
0peziFT3i4cs/fVjiZMT2AuJPggaQ3MuCHXHv1mDmLtZbwxeLXvT6NCvy9wBShME
SQTANf4IXZFctk1kcTnXFtAUE6iE3n7BH2mL9vGb32/HXVpHV8Fa8j8YosMlWKVh
IDxOgx3JOfLcWqcwSLWU5OLfKegLua0Op0wxLS54LIyAcrApSYAnyg6P9fnZaRYT
pII4NYD7k4Ba89GcfF2iLSwfDZpoR+Yoo35lT26Lmd8/0EtOTFx1iY3NjfWjW9Wy
GhyNpAZfAYHlE7ypR4qKPNy/sIBCS85xfptRN+ErSUNusmSuEhvdTd6TWqTn/dkD
uOPEpfJAGlr++VlQ+gLvpMEt0N8YfQb4wWr4wEEoasHRI32oUPDBW4CVrZM40Xu2
dLRQO9ATS4yJbVAiZvoou8blZqsxOUy+15ePU6L6EHr6D+idAzOiXy11QTTQmmt0
Q4IFSX6ggZR9/JAgcH/iucYyf5gt7H2+9kiT2zUcsWZky1t/zDvUBRSS+Ohb0tVW
PxJvSc3CU/hKLBWWyj4PsobBCZYunvU/aA8wBulqtAdBvbhjNXh+CyRNkBdl/HjN
Onx9ohq3X1ZRfPZ94g5xNIrAPVKSyXhvikp2txNWd6qvCcqH7Di9aix89FxneZI6
K+ef6Hw1uBnl0EkEZnl8DSN4N71kFyCCatnGJCgxBAFET4gEAwK3Kk+Vjs0M7hv9
ZKIczfSZ/M7tSGhjw38Ma6MX/5WOOrTVSYoEzK8mYhwW/idc4+jxpPcHOKIwYMsO
vJ1A5gH0Sck+n/dnJYdEJL7PKAkucWndrnXfOtrvMO0ZukUU7AP6LUwi/OzD0x3X
V6KrqH9ZAIBoJuMV3cmyhJm28Bd17E0oVSTMluHi4w8P+JO80x22WBR8dPgo//SR
k0rMYmJQ8xdkXyMPNTCXLJQwMn+8o6so7psdh4Rjf5ALsrNBaugacf1dRtLMg9an
CymLCPVBFuEmgmcV7HGiRa2gl8jHsY+X+UezjEMQ33t56wuOrNk8RkEkLPA+jk4A
oBCMXltL0Y/VMSDCKRRQKXP5zc75dy+T5B315zcj7M2+A1plZFUPDA74AqGdEL+5
YEXfjnGIr4zax1NuQZw7ey11pT2kxzBp1+SPukTVd898mTrwPXlM4fS0/MIXvIhE
YIB83vmYXykv885tm4lFPEA2+3h8kvygNZ/fcsHM5GJ4zDintDBICdZyd9aHo0jm
qw9bbSSQ0iBAnlijPchETO7HpygY6UJxxKJC29Zxv7Fq/yYqwjfz4r8T3gtNFINV
Qu4VlN2EuMBuvFkMxtzKJwvi15pBd+zFwgtA5fBppAsEiEBiVMjH+B88aX4rMvrD
4r422BQ4LVyvYblAvBN2RBvxMyU8AyCh0ruhk/UiUKYH8HVF0SsdD43T2FiM3sne
ZPhvsLsChlLqrJ1i4znykFH+5vDSRaNW+9+oh9l0xLDXMBN6xrjWq76mtzJYkVE7
/YGLctCbJiyaqn0d76zEMYIGZmnDG9D71+lVHH5ZLlIHfrT7pAad6yDib41ZrzeB
gmwogNfM6eeZ0r4B298zNu6n7xluC9oTyMbXLsADL9kMcPj9UMUYgA9JfVM2d0wQ
f4Y3lKbSYOQahbvFwVLgBiEWcGCnYhhGKRJCs3t0oU8EeS+iBnp3lOMIv9Po/ucD
DheLE7dukVAiXk1buM1mn/poZ6NsGoaj7g30hV25koNLdplmXDKwMzh/AApBqoV/
fbpXmndXCxHSfTFJJ5Az9NdHnneaipP5KGzyIFegLbVIOJcf76EEYA0kLiq0J+e8
mf7erPuawoAEAja+Fld2dDvzViNDYORDXnFJt7iCTPRmP9kvba47h7pouhQ0GUK4
dCuHUQHUFjZd25sgrHCWoBEHP1oAyvs82aBAbj245vROHmwuivXCLeFbeT7xLZOp
bzY/MlpHT8TlnEniim+WvffQ7NZfp/UMMdVsdaBey+PHi6iocv94M9iqG5seTR2T
vXEM7fxjdFmlb4fS9amZkIGlkiWmV7+xwjGzosHoqklBI3QxCw3Fev3BEdeZwvY+
6DfdExsRDxd98qy9RoxJ1v/7D6qL5PM5eAr1w2tB4cCKH196fgWby7nmC1wPKesM
SSjT6iQVU+bm055pZAWtLjILHV7SsSSn0O2KMY7kc8rqTFk1iqWM1rNnVOqZcWSE
Vrte7ZT3I8bbqM8KKCCCTB9jkl/9Bq4pgAHKDZrW9xxl+ridnT3jRbjZTkF9AELg
CNeQnWEba0yy8IHJRb4AaThbRTJH2QghEZhbmJDr5eTQ8I/pYlSffVOYOlCpS06J
bRDbnaBpYa1upWz/KBWmwPoUCB7RFatwZW6ViZWZhJVXiMsRgBIdN4PSBgB/LmHu
jGUIuOQfu4eeIngnMFynCxhulQJZhudprq3NVqe45C2lylB8gzlSGeSYqcEn8kke
lDWKsq3w2g2Kg2Vgrs41NHNNhd1WwI4ODctX74rSmv88Tkf6baZ8HAywAcXLhtv8
0nIXO57Ip3yukJu3hNWThABwHZsCD4V2LHSV4sBnOVa574rC+U3ODgpbxIpeDyTW
nuRijPuj2g5LC0+wAUPdJGM0VKwJyj9RB4wWg9u8JY7SFhJk7U82qsBKhUL8Zt8C
evbLiuZTukFRrlODhjLkML4k6BuRV6O/rDUGB9GDaris4RbQ0jQEgl2bMQrZbxjk
K0k7CklSMYcPkuKTOY9nC9gupWBraMa+mE5Fiyr1K0LwrVcGIniHbEXVaih36Chf
vc65SvP04/SJW7tR027KC08KRbaC6AA1rdFBkKn/SoN6FuFlEJTaD7L/c8sk6rkU
mc9Aq0g+X3QahiSPoEf6JW3UUzjOWc7rfRK7OkiZ1MtTXDWS9CsqG/CvrVC5vH2w
Jpoanw2Ky4ecdJl3XXdTwLe5HWfcVHzNIWBEbb35aiEoxZjxhUG7hn/VJ1qj1wmU
IfpoGsc2OMr+YKeDjeh0wau8knpd7ASr39AzsV5jSl5UYwdDbIJ7h7JHRvw5MtwJ
KLA2ddXArg40g7bmYySwziOXAPGVgv7xiACShzPoEP6qGrGpH8ZACoWojHfgvsuC
TRNpdUfQi7V/a0nPQbrW26T0W+UYP1J52fV20y2UM4aQZoJUMe3D5wEJ173lDB2N
Qlp6mCJA71mc/rDaX5RcO/6A6OAo7ffpD7GEyPjz1ifXiNA4HnHad+iDrUtWA8zi
8RJCAc9ldQ1e+L3z/+2hMVKjuv6YgvVxTnoWegu7G8/2XgGMnhpJij8piovJi6w3
Z94YvI218hHj/HoqdfFIEumFu/5AEpmHYV6Xo8PF0shVETZB2GYESVQ3njdazb0+
6cCMlbJVlQWMppZdN2Sr715sZGNMIWJSuKkPbCuYzxLRXVEXRuGIGwAImssyW6h+
wCBrcb5w+Tu/7k9zkQ57xsRbrY610nLDGVJ0YgxNCLWLs/2V+CN526hw+Yns7aP+
CUXCT7ByHWBgKExGpLQf9hMLujTjgJzHE5JAlGQxNkqUIAvqThJot2XYuxMRLxBw
zru8dcaNOU2uQHpi4gAffpsfmEPwq8y3x/HxlijGI7TD5w7iHcgA+ZHEr9HKHTrV
/cwQHJZcbf/bR2KY0a1aRCNMlViQtaR+IJW5f8yUS5d8JmIRAukRLEPRYtYe8Dzf
24g86F7t4SBwPJcCIrl88uDGCNl47fB+wvATSIexCi7qLxWwP440BwEqkyZMlwh8
Hvl2DpwgNDu1aRk4yQqV2jq9+lTTBuaUNwT+uKY1zkYcKjPxknhzh8A3sZ3JlsW8
N0wQPtIu5PsGfF2HZ8CLhntkQOmQ2ZqVTlIa2IN7cbkmzwbV03oc+aFhF+GAVWjy
xhNQQOk4I1Ww4d/c2oRYOnjtJlNYD4M1lj1QTqU5/gR2kMSNLigD5P51pJ/F3S3a
OUEQnuicm3EeO3nNAe5Zo0aPIv2uwnH22du5E9awmTXCe0gkIM+Vm4Yxaj77DCVW
N+aPSLBcwpZT4HTm5II4hjSQOx2QHkIqrY4NVUq13LfzpPLPbCsRZrDB61ZgUPZz
9/FIiwqJQuPvxlDxEPxvYeB2DfD9EqXaUB+9qTTiJomPRRA3Yp+kv3d8dhRepqxj
uK1S9dbC7Ipa0Sdn3mvomGa8EXddjZTSAR+WlRN9mAHjhtGIWtm3QB6WGpnt8ZXj
qJARGaOldkylmIQBdI72mQP1E3/RL3vZIBb7/MW9j0mdZ9ESxmIfaP+qyPY4SgSk
VtNTVRBEr0w4u1Lmg7SEcOhCZZCzfP4SlSU6vutobqE13NrYpEVMnG3S4sc5xEfH
XDkute7bIKX4KStkSHR4KbZTC4w1U3GPFvuuLr0nSPWFKu8uPBM+E6s2JyHJTTvv
31UwlLukZdri4FlwDlTeBZxl4deW0l//vfQNOnXSgMeD1XUDrvsYB/FUkJBSVDPN
6bM77naWgmGJq0ckTEGgjWfcJk4/VcCKDbKnXhq/HBykO/dwoKJZCA/fcHvGg4bk
FREWMkXsJbKKPhlGLW4hSGgp6PpLQKyKbPMxNbU5OfrlUz+n63CMeq62BOBUROqO
CBcv5HLMb3OiDu7JgOpnKEF4SyJKjC9x0QvHrAKnNUtfZvYP6yZXZD3nStQPn9iX
g0CLgMiijH170JV1VlSSEFgEKq5vSw2+kODdzwtPqQQN3BkncCDiAxAe/IUfVSL/
jZQUEswN7BD/T9mwHrHevSosHTOXoRZcl0e6sOMHanRFJkfLmdLKG4Jejm0ZrO4V
g8ROvEQjbGqFmf8E4U5SdvKzV8Hozs6JHkiLZQMVkp6Zpy5U5G3mUHl0Uy0CvPSC
HZ7cQ4NxmNEJxl3kIilhx4NgsAu31xRaDtkq6OY610kl+D4xrZWDpF56T27/uuMk
g5lNr2ot4nT5coMelKItV8pORIU6HGPbwK42VmsIO03FrSd+qZVSAPiwLIRKGWPK
wDp5QPPebe8CqYVf0jH/LwAWdxYznNgjOAjZIjdBBn9gEVtQAyCzDHTN77LEb9Cx
DiooptZiuwTh042gFoKEQdPYt22t9YNnlsNhjPjUHez2cDFVVP8MK1N46rr322MK
eYSVW/j0NH0KXSNMPD/OGYCpHS+X6bhDzr+R8cOwwHg/dIeJNugk2KiS2JMrQjMp
mI1G7FCohVSO5Cx4Lyj1c1keFiOqdvk79/YqKAxvjTI1xcOjDv1rMi2pPA6RmndV
Audv5kpH1Jgm5cXYZMp0HfU+AwqronWtHiKpAL8JxYjOkXAqTHuIDW1FEtEerxAE
DMNZBsiT/x+BauHfRt0JzFm9jS5UYnCkoG2v47BQiD7W7joLAfrhBFzr2cKwDLME
DtC/EiJjfHZjPM0NyYcpttJAjzViEUJ4qgzUoyQecse4UOROgDWGtZPEfDsEpzVJ
7+oAdbtNwx1jFo1N0Q0IqAilkoXUiBUATAH/1+NQrj4c8g8oZt9yF2Q9Q96MHZhb
XZ6mizkxBtNc5L2UXHzFVWlxK9mdKeNy5eas3KniOu8sKvivcB1rXuyYBRaMGwI0
VZVB4Eo3sF3MS8b04tvCaNm8voH81izUDxmc7z5mB8Mol4agtEs14ob9WYizU0OG
h1u7dYvsa1WV3IVxln+Uvdql3fIiF/Hj1bafhSrLCinh9pGICyfrNMrXmk2xOitI
1Yqj+OKMHDT9r2qSVlU1MMh6V9f21GHCiqvZteUhqeyKQjEcCt4W+TFXAJcyLgy0
8ErPpMSToI8ZVmrhvSjCS5hcX/Y0cQJqKX0fZKlid6mMELHyV3jw3raLNpLabtzf
uPsIqrJpV2j6UpbzT4WBh/pFg8eSiu5rShmjVpc1/j+DJq9hBAMS4zkQvtKydy8p
DMJPrHK9eoEr1amBvXNvvL7rhnjHZHrORd5wQ435YD1MbJRDIBtHc8Hjni5vY+w2
7j/2YffISf3pVMUEnNk8JhsIf7RxGwKQOV6DwL7nJ3K8RRc9m2I/Mxb5222Io04Z
7big2rW9OBSZjIzJtesBS2qvUT3pQJFdP+Sr4g6dL3+zbOPYCLdYK5Oj0I2Y1e2c
xVkFzktAYRfRdvx5no39G+9K6zyw6Bs7QJ19sJ+2W51p/7TiGfs8gPz+KmVmj9n9
YL0Gs3IGBBP9j5MTsHI556alarbqCk1P8BnmkUQjBUsCtWZCSSjumNl/Ipa2G4SE
QAbGpJfbg7KWMpCmB98znUBFBXR6Q9P72/7DXzPzo9IQ5LkfFc52WXnQKqTrKIUm
X8B3mdkzBHeM6CRZVsYPibSY80Gbj2WjvM6wNh3yeKedS2Kq3GarZKUeoYhRZVrH
/dWZXXwhyb+Yk5QENyNfd8aQGfFbLFTZ9OftxI3q/0fPDPPcHn13G2A1gtByEg9x
9Xl/6RgCSaBz/+ZbtbQgU2tz+xvxfmRFVrbMUQPmQLK8nAOLIAvi01z36XjJVqP8
p2YTmhN9qiCflAaG6Nq92xVBG2VEMrduLx4zcmTTbJnpRPt1xPyRxcxddNoSzLUg
D7PPsIArE7CTKMCV1GFVquaS7+U+bfdy/PbL+ftsA45cUeca249HKTTH0nxnFKrI
z+G1oVSrwAbIYescp4J3BupztOuBuWCeeavV2EP61L/pvppljoTRzYpqBlh5W9Qo
tOcHy/tfdUDj+zYBDAlnL4BNne19gBbDxM0QIqTLLNMCFK4U9jiMYVCTyQs4CRBw
lmYiaPbL99MN6xiD+qAq7IppKcM1zd9MsmhFWSCKw56AAmNcpBEgKln97kjKsq0n
qP7jdfgHTbkTQPQtz2kBc1l2FVKOmrPFqlgubq4w6yjP1Qbht0y3r5E+M6LIsHDX
fGU0Ai5C6ZE0f+pJSo4vrITFwF6F72Cs3orqWyObWA4Gr8nv5BegEMeFbKSTXyvh
KUoFnpeAwRX7GAuTb7hu+LeiXnyaVtZ4XOQ47rMpH9KWPyu/yYyxCAocUzdPP5fn
yC5RPJrizi92ziBl11UVLJYa/Ib6fvCyHxjLCA5lFVw5js1q9hVcQFqFMdBzlmCn
MrkS6dMooi+pY1jl5AoTuA69jLDmz1GKbSrT0h613dkkd7U3woVEyX6ZvH7phHyb
HiLru208d2DstbmA6EEEIrfrvJuw2JrrZqUGoDknGR/48vsIuIFHi13SKuVzl6Lk
RNn3G+SS8qFv6yM3N6apTbUVpUGpvd7tLQqXuHU7N9VWYs+pRvQ5OERXqLu36KNt
DiviguktvYtMa/ZoZa4wiEyO+rCtaHfe+umC+JLcDpBwJYMCUpcZNFR9vtfKCOkE
PTtIDdyPcQFXVlCyrl76KMk9g1HxjKybRPvXX7w9u7zpBt5lgVLHJLNALkLUeiYG
ZPLMRwstcT0kunMszBPAd0hjqDTbV9s4hd8J5juUqkGSlW/5/ChNfG7kxZNhT3KE
e/2GfjDiftoPdkor0JPG1riW1xX3ajXye40WrxPWkSvpNIBqS3ThymIMg7H2BmHj
tlWGde/2gM2lVmJwPjp7SMxPb9bMkR0oPuWTZwMZYeCwVVC4SbBZAFOfU9wU9IOL
rrYBybNQx4Di7ZjR/NLNI3KUBKEiuCQ/0go/q04dClVIgkKxttVJzhBLtgLrezOJ
jdV8u7CRDZ7+HzulTvZDse+Qn03F8u5hjCYJpMyPYSxfLbWKcYBBwFbIGDveXh3A
NNOgmnz0iLgxqEMGXmD1+npP9S1yUSzPzh82WNX/gB+HKsPJRRpWYiVbUKxCFlIU
G/HmON9Oq5E5dIiEbcJji2+5mdUslGVyFCzGCRrupYBvaQYFkKGZ5xJCz4f3XdS8
aOylYT+OV29GdkPaHuGLPN+X2xH1piLEbANVySdYLk8iczceS4hSkplMVNAbiap/
rNmLezy7pHHUFhyAfMizGVA1kLijzb5Riojo/0NtRkldaPlWQyjrTFv6GW1xuXW/
2QEc3QlCh5nawVv4wKg3IsaNVSZcD76EdiUxwgKb/xHHoN+kBdrviBYLYo6cNPqt
Tt2Plce6tIrH3W9Xi3U+/DhDPEFYPGTNW4O9Rnnqvh5i3pw3ajIWxi7dYdavXlM2
sD4WU7MGBxuNLEueTeHlD0FVgBpaDOjxJH5UT85zPDDvunziaalSIUDKnPIZ2aad
AYXrZ8ymknkHe41OYSh9tpj0cMkkwbO1jvzCIt4GWmnXgB6BJu7z8yceAOYKhDOd
qFVAszffAmlvUaLerSkoPUMBC2jJXImHI981/tx6HIw6ohJXBARMLOYVjGlD3n+Y
px9bsMFvAqaGPDZH6/ZBwaKP81ggmdjX5bG61IR+ct2wZaUvhIOIV7NoXAwr4g9b
J+bc7alCP+megnFiqp/KeqveTCuk8JEA0FSn6wmuQeplLWh+qxb34rFF8L/MrDj4
gsimo3rk0gzDh49SCS+62rsE8qZZFTPtqNK4jN4YDYzyHoYTvpgRuwWTKFD2+x//
/LWaneKcwqq77I0E3wPr3ZDH1niABmzHXy4qrT0AMl3PAB1wminNc8VAzGEYk5v2
j7Z36UqSiEeKtVWMRf7O/1CWpopDpRFm1IBUfncC6xNaG5pWzE2PxlxcHG8GFBbS
VhhrUNDKq6M0igiC19NOl1pceFoeNBCKP094Fkt3x5mM7JZkkVISn0nhQPnZQKSf
2q52LVupFBQ99d4qyQd11lDivesr/SHZMl7ajXerJsec6oteerhZ50fUIZxIAgrl
ptWEE0kwRR+DBO3kqtIJOWfvfjjcjjBE2bzSfHlJnwCiWYPaHDgW38x4bJWTp4fH
r6FZwuFlIVVjhsibOu0NpyvO6FRRCiHuLN4mjuKEax0s185qV+er4SRzlKVhrkbA
sm1NHVXRfVma+SV9k/LXfAhWp2YtTsiLmJeHfqvv1k8+DZB69ENtalnJ2LPP0tl1
c4j/RPICbGm+/CElshYr1ZeHxjc4gGSnclUi6zy0fKG+FzPeLz3inTNhxW0w3BAR
w3F/Bj6T0IafuFqmxYQ4RqU/PVY7o9e1wglt6/T5jeEZTFSXbuz/fflD4JtW7qvq
LNbWGICKJj4/6dGK4gdoIQgApNWxfU+4Ysu8oDG1V3jtwzVCdZPLRSX0Og/U+Cgj
KyIeFT49EUbqPub3LxA4MsdICRkyKSIkU/str8Su3u05ha2RgVyit4uQljOaHodW
6wTp6iajSHvUNDNUcFrX4Q82X9SMyTXoNFSc4qN36LCGcs3lF8EiWAL8XYgZ6hHu
SN5oCYPv4s3YTz7JgKtbcTdhoIpof3irB/8pvReLK2Ua9EnMI6bnPr36DRffegfX
XzVy9EkKf+xnjRIo0hFnUz0uySGPqjC9zBGAZ6pmusSkNy88RrqFyQUXaRE7g3XO
LhYZhXB8Z5Cqw3CKAtgDOsohF/lEw614QV79mOkcZPTtuoXWne4oNtR42gUTv6AS
O3R/ZKLUCOScw0wpwJHnaiqTlY6NAOmkHYLVuzLXeHs93ltd54gMtsDamtO9Fw4B
UDs3Mwqp6LIjbigbpoIBbIM9MSsTJKOVA/wF91Drgv6V7i9EYTnU3he44gPDj4AK
wKlP5gwGLFpjkNUA5aiaZ7gfWxretfpiR2Yu/JX0tqULEwX8+HBpg6hSPmzahWeR
iChRGG8abfpUwy3KVAWINdGM3pTrZE52MJiCCrYmetzw1r7hw8EUI8rpk137+0Z7
YR88X4Sw9jAdFhMaPGRLDYtr6Vy98tVUXeRs0BNO+c1DeSQuv4aP0ReZz2C5EVjF
hPSOYhwBJP1SXDM14ERK9SWfTtRWEW0h+4u9HeiYv0KNjXYlIiAM3XqJ0PTe9TWM
ZUXmaHMoi+k4QR2CYDY8Jt2nfWsHqWVegOnce6FyW2YiXHAN829I3GoIHnSgFGX8
WJ+KRzR62/jvcOSj7kODuTB3D4/AfRS8dzUJ/w8MmcVIdsR2jvwaaAihvjDvNzev
TsnTb7RU8pa8jZv2+BBAouwfNCV/27lKmn3HYHbEvw5M54lh5cQbk963325228rr
b5zTs7IShILMIzi8vaoyQWRgRXe+GD+6ZGu5I5H41P1p9fW6PQjT7lgnoifzyF7r
IvTZa2aMZxkm00h35TIxgx/qeBsT4ggZqPukNzMZg/c7LMz0VToO1+9HfBde3b+8
ki9kjmT/TIhw+lVcuQAxE888bPOR6vecwLxtGjyxbAXakc26kHe5jJPoZVnMxbb4
M8avHC9NFwWh9IvVWfzmc5NHKZCjUYfQxSmZFZjjgGKeghmLHDVjIz0BpO/WHkus
0ggfz6pHqtcwE01T9U/ogsiWCcIzgIA+7sSE85yu1oIH76hCSYLFlpePSsjUQy1S
Qph3vzJtIPWTc6/PO6NRysnsqpXjwRNuV+I4keqV3f4Wqk3xoEZxMwri5MA466o4
+1p4AEoNRI6gOfJgGdGF6rIbCynxpMaWjiRtsy2sMfYv5SdenmFcXDarwkTlKqmG
+V4HU7cbOffcbVDIFlRa5lm+hNuTE+k1qfwtAKbjcgTai7P6E8zjra2K5htgoHmh
49oC51W43dQalQspMn6AqrpNyOD4SMCRQnB9LKxhZZRdtq5J/adcLfIy7bxCyM/q
WpIryOkS6y+r4CGPczUspLtoOcC2tpnwhmwSMLJ64f2A4mjZEMZtstUQPRZY4B1J
MpJPQtngeF1aIj0iPMj6t2N1WckDgftrTTO+g5AEk/m/TXJh/y4E6mdVKyvbB/3+
VIPCHGGVraWvemuJtLsrwPJFSViorO496egcq8nwbyuxJWw/tFi6OSB6+wlF3eBA
t55ZjNWE6iK03m6Zfxe2raGGnebRQ6nSo+ys0Un9RynXmbmD+ZghpUFhGPQOmsFw
XDkBSDaqjkZdFgzI07293CYiEVkSz2PTFB/VSn5dchEyYzBQYckIhQ17L5RSzrir
/6D0CCPEsMi3tsSfBzP+/6JqwA01lfGimXD8sOK+z5uDSKRy+c87oPu6mRBL1Tt+
x6rYiOuSx1D+jHwkJVC1M6bJmE006IwSs5IXVITs8ynFPI3M7SRufR+7McRWyc0L
NZHPn92LEgzWbf+Uwa3Xx/wFlpV0pl1KHJwBjszSzvpaWGgDva1Ek8PKmognatYG
DPvra5UioYWxrWEDTB7WhevbSppLxdLatzs0GqoN3rNQkGUHI5cLxPqBlNCJZmrS
yRjbIt/lqnCo48oRzRtvQQlpvAKTda1lRtAIOaWnvOmSIZwP/zjrennsxuAVi9+2
VQiDs9C3Gl6Uo9AbIy+hhpte9c50FhFLTCBqWPCB5JbMq2a7bo4j24LKYj7VmINJ
YZGKQ6z+E0qA/5FseJlZFGdnlK1u0zA4hbOE1DkTSfiiVILD2/lJ3d847fTaPzd5
ed56LgyXg2jVamWHWf2E5vKwEwYAP3F4ns08hnEoURR4Rr3WFszDHnl3fV1tR5/8
X14MDMJBGujNrYZfMroz90+4LQVtKSPXF50QK3LbwUKZ+drDCyWsey+Ytxa3GaT4
2Y5asrCqq6irmjwCoj+7dIjPLiAgtRRcXeT/Ju6ufzBGfF9VeQmdWhSHODA+5y6S
49X3Z6QiVKauL0NuXEFiQFRVPTESu7PDVDCm76OUanpR4ZyY6DspiPMQUBgHAQ6E
SZr9EifVn0JUmvcJP/wFPouDr2OyRMKez6iY0lDJELcZohz+0OgqcUE2PMp/Uuy+
n48liQBbwvOLND955NyDileofQXbpuFQyWgPVAS/Y2g8VvY+muSyZnBxplDOZ23X
u9a1Tl1NPJJ4qudIU/11UMmDIZN49U7Y10R5cYysSdtmlrGtf87uO5frjSlGf3a1
O8nGsU7ViopLQEzc/xV+sR2Jm2XX8Niyq0QUWP7CS1eh1ArEb4MUtCF1WLuInbbN
bo0F7xpC/wTpUdTejHCFT/EXvhSHMPJ8KPsnXjNnsonqgswWqx9E2KPbnM3XZJjF
xG7M7v7mS5dkIJia2iNqKU3yc+vPutDy7Ed0B7kV+wJZz5gBYMjmmHCnAixRzpsf
scngb5ylXoQZgi7YLq1SpTwOSlfQeEeT0JUSSmTaeXL8FuySGR875JBjIxP2Gjj6
oEVSWA7jc4sQILQaAr5WeBmdkoxi1/6ubd07ZOssk6d8JHlgNqwtEl+yvzuF1RMs
Q9R1ixKbPYF6l1fkNPsUcDfgpw77ecE/hx+iMx2fbJdtHNZ7G7CGt0bT04A2caCA
nr7fBGnj2OdbA5eFS3vREGgpeUmMcYM6hyg6oWvk074j90SpCgMZXI/OJfx2tBG2
S6bVOsMvK6wPm/R3Aqvf9ElKV8gKutTHzOZGitjbC2Zn1JyK3BDNAS8cpP3l9Fbj
sK1q9diyDcjK9WvZmvXBG7N/PqzPF3judm24wQK/B/fUzoFrMRk1nTyK+yqGDbF9
xMRoG4XMXLHhQv1jHXsm1zxglHfq6ZF6+crL9P33lK63fny51MEulOb16yUUkcN4
is4+hHu4QbNbpTdqcaE0CXSLuFdx9zzrPAgSlwMKlr+1j9Fs1MDXY6YKTbXKFn6S
HsLCiflq8+G75oCBNwYCvUy/ruNjanUEQJugs1MDD3t08Z/1Z8f77Tf6SM0ZSbiL
Hk87MYhH1E2f2ykZZ+4SBEVJEI1SamHX+kuM4mPKyDe/GBLc5djgOJc6L1jbnBfV
v0pjtEbeY8/54C1NJzB13VbmLoRIT5cDLtGDdsVm3g7PLWj5dx5hknvF+ErwwlM5
Dtxp3XWCy4Vsy31FDqrgPa5SNLCKaUYvrBeICzDC83T1x3qHErAsqsp80DTJJOk5
/JjorwTOjvPY2kMIgXIRL7VB14NlCoVJ14qRaX4BQViXVoGSd1WJr20K2iOOViLR
OFLLEbgrpbfenBM/FlySOxONT1tTuc6fgUvC/C95beckoKyygvcFsepqSzs52l1g
DOUjJQNReOHS6Ne/T1qSxcNpKHMbmXrJGAVKIyM89JP5K3fiSGnnWvV5mhfDTHrE
7/HX1rErGX6XJoluOHRvYzTnVYk0+c6lKVgdI0c8GEZLs8aQcq3NamvebdD6tI0b
UjE3RhomxAYDB+Q28p2HZ1ds4vh4Noqcku+JL2EItkgFsBcIXpX6n95nHCGvSsXO
DXC8xfGDpTXklboKEGX3Z9Q9/kunHX5OFPtdvZZ7Nt23DywpvTtrs0t5NyVOFjS7
YOac2C+Rs4r2pA5hoOY0HxDXWZra36BlMrqNUhbreOp6jXbw7FhASEOukkmBxUa3
O6z1U6d9ZxuCU4pg7irz/yM66XtgN7aGXziDAmeuikreTA3l2DaN+R5j4lIo7b2S
HImOUk1/UvqMMKVVYf42AepydhzxKAQiIS/VHxqrBwosoa/QG9WQA66lxgG/Ri7b
OaoG5Drf0e+nLziHTTDPYKIy6OcPIE7vAjwebdlxbvGo+fQCYl9bMFJ9RkYLUsiy
JEQN9q2/H7x26+QZMMF4ph6/p4sb8YcRN9fsw0Ct/zydyATU5F0sYQc+/HfiHtOF
BI0mBtdcT79bpNXdXYp6U7wMEi0dgEbwhJVZMcLwkDeJhq4mOVc/F5NBqpQd6lgi
BGTJxa/Mgo9cJ6lrW4H5STW6+6cU96JXNh2FiKazV351xXDxFeqE3KsGNqpBJ00t
z0FaTCzMV1Ls3FrL7IxeUvWX35FQYqObwWOxh6DkvUrAjaOLVdQ3s50O/IH42opA
1rbe38fpEyeZ3aKBkNfawQqwdU5wBcTu+n0uFo2jHLXf/L5N4TIS1BQf1Q59sReX
1Fb+OQ34b8GeARiVj8InG8YvM9VKeOYplwnmP0Lc4Tl7h2PSr3BK9g6OWOx6VGSj
ENm3U0BhkSPapOba3FZFLvjO/ckepHSrUonoEe9L+yQ5lxMP91+MCIUUEnXIjS4b
/0rm7eGVhm8pBMvqBy3XxAewQjP8JPlYMpNNTn7aVXMp00mECC1swkiQUCHxQGl7
y/XulAuVzY/y3yAan/W3R4vn+8OwXsCwgWAQ8GztV6ARuTJhvqKFBKe+CXdCeqNi
DYr5tpT2nt8YJSoKrN9ugdrWeFAdCi5/M04jKogkKXCuqK3DboiWG7KsrFJvaTww
KpLOMGi23Dfil/GOrTLpR/vY7t/njwgPeuVwrQxoboycN8IIMaLEglVEUQudfXsP
fZ5Bb37kAhWFhFLNlOnmnHHeo0kcpwKznW7g56VtfQwSlu6h99vi7UDx08jdxVDG
/HJVL+AApsw8KQVAkK5lWd6Wy+gULigAa/gNDXHs9UnwI5+lORaoyAcv6LFqaSfk
+CwPk/idQ73SIo88NqeoOGx1EfqcEbYEHL4+vhb+Eatu6Lhrmmsln/IF+oJXnNzq
NC1JAUv+NJCE0LDPSZVHJ9wY4nUkDupccXhf1DvWgzTZi2zAQAXBiVjl1A/0s5Pq
O5nktCOUbeLEIJrb+QY1SFvbXnhSrP7gyq0r6BMquMaAyyDet+0lGeDZC+wUwR7+
37nKlSNAsc/jv21b/zzXtPLKQ7R24IPCUq6etxF6OT6rTKx9x94hYiCtKbvzJ5/2
4gzJIDQqFAtPNJanGEKxshU6u0DpN0fqeEq0Bkb8HRGLNC5Qn3FboMue11hQloAf
PKEgCqxKJgevRJ9YNA6AXztD1sKj6NhHlKemwGwIeFbjS8z0qTIvDPnlRpFXWB/5
ndhexdWtrX1RWJBwvpgFbhQfNjJD8TnU86QSDHRiP1ZyS3pyzEFBd0YXV4m0AveB
pPNpU1aGcUQIb0cQFd+3xWGiL4cLfGj56owuYakWxTEIG8D99j2YoXVL+o8UJI21
+UgIaP/s3HFBaeD1QmtGcn6gSqRksqMW7l9SHcHIMOJISOIyWxK8gTSDanAFlmCV
+yzBExy3wgVGvujHMIMqNOI0lfGIoHIJfVcRyyF6HlRj1OALS2TylsvqnlS7dPwk
dNAj6nzXaoJ3XkAxPMRUDTPij9Ccy6cYzMzeZu/l2nqqInJJy4OqumrnDJoQaQlx
60HKA8aHUV/1abSr3eSvyXUzrpaR4dmrF2uARWYT29WQzvwzupebZXN2nWSmLDq8
XrrkJ59Ghj6+EMeuic3hXuwvc9rgzS6CfJZsaKT7zELRR/kHxA+TuU3mIYnmluyi
Rq9v03RCjkBVJ3vU+zlFNjhTpOgW07Q6pvn0BeHqFsYWboD1JWDOKg9E+dDMGSAc
Sr6vnp1sF1P40DGCWwQERZkYL+WX5/jX1Z+9OhuQtaeJXvURSIolN0btjWzBgZ3b
N6N7SKYF/mpP56CefVDsnQh03/8q2ns5LkQm4UKfk4+RKP7GfHIOyDc+6LKP9Slf
xI+abJm44AqL98hpagl9VVIRKGJoTEFYljV9jmtLw9PcYGT9LLfMBReKcbstdPbg
1PDuaQrlxb3PVl4O9inJ6UZKqAoKoqRGh0aVHjoyYpj8zEnTkwUAKSZyjK9eySzu
yTEOyy8nm9Y2giDoDYegiMfkMXeFshk/l4zOxrS8KOAqzEq3NkkLUohGxuqfznWs
niF4598VKs+Yl2O8uLnhuL+YrkU8HJzdo0JaeLvtodLqsHTQfdMIL09FLECP4/iJ
+nW0px/j6mlSH2TSRhmGav3Whcqo1AL3X3R0uSK2mVnkTmvHww5eB9S5tyJ5j9li
jZ+3JXt0jL0ls1U1va2yzH0iYzAS1fB47zp7OHoBEkS/w1Si0N7d2jG+o2Pv1mN8
gqicd4pLhp+bNu5Qtxlb1WdKlEXQTclJmsRqBPxWykMxSNa33B+nvUCoEh+L7RyZ
uOOqNvfcPtlIzWSuPpt07p7RxNWCrvFXkuxQkwgoO2zOlP1G+326ovWyj005NGbd
hiYQP6pqZ+AlJr7f14106nn7a1CPY3dj7p1tXw9PjW6jYBubG88/MPfw1E2aEXz3
3MJDCa4oLnTqhAY9NHfi7/HPyVRIHkc/AtTq7utuFzEwOLQPOfHi7sVFqfIwrIR7
TauHdKoW5+f29NmQgs/V6hLox56DEp+Vwh+DV5Q5J0SAwqj/Oq1S59Nqz6B/05AI
FXbybOScUMRC4E/IgAldaXhtc+QApVjUPQuqA2NBrh4SI2Q26Su9WSKOZjHnuTRh
suK74EHONGzIIbX4AcyzCjNGzqznxuhqp08+ZI93QLoYU12ncqvlAcocxvH8Ql2l
mW2ULEgbPLGuMGyVuBuEk7kkZbJJKIOH9+21qa5tBGFzKrvvfKW7Fz43IxmPJFKV
`protect end_protected
