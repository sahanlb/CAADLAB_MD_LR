-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Utqc+FW2+VZUMi3vy9HNLF+3yTi93PxRz7nSfUsF9WnVzM0pv/GDoHM3oal4ZJdW
ICzjSdGG7q9Im9KdVdmA7fRfhC9jD3wUD8NmU+qRvTxqoS4kjvUoXe3dm3WKtAez
7IvU5iWXeKV4PG30BcA0+Gk49pR/6fxUtP8tOoYUZ9r3tbxkdxCPzA==
--pragma protect end_key_block
--pragma protect digest_block
LWtrLfhoOCtjGT0JOccuN9ouA7c=
--pragma protect end_digest_block
--pragma protect data_block
SQ50lRghw8lQon+aSsL58eUzawBNiHA/9B6fYax4d0A//v4MTIdrjcHgoBD5IMpG
rX47zzuby1gni0MVltt/PNWRb9tAhvpIKiGFz6Jy8iihVZ3ZU30UtVx2zEjaR/mB
TqF9OoH3AxsMKxx75arR5CWSyvtir7YbdEWGKRgl20pVP2lfzMQw9LSOTOvi2vnb
pxU6vG58Fixd7hMOC54/vz4HeF6hJUAHN5bJPTGConzyD1rJwv/Yjpd3ybNUW6N6
RyWdmHiLFWev0u3G986K9cvuVMtIJ/+c4+d2UsvVj1RbcN9N1Sybc9AGxQ8yeKwt
UlpMybRpPwtL2x2I9XmCMEwizvCaoX2sVz8EEsXt2ElPYXvtmCKibjTjnO+sZ3GN
OD2qjL2BuIImw/o+ub1v8BeDbvkR74hcGQdNWDt982u1cZIf744L9O6v25Oh/aMu
i1LQUPhVlODgRgV/PpaIdnml7Lj6j355C80O49mjcn2KfMRescY8/lxRk1wqTA3g
ABcqaHzdolp1vYHji5t7a8pGSOWDaPthSAq9cwW2UJBE3ft8GT8uudYlw0LCVv1V
rf6l7NdBjQo+V/Sli7c1KJSHgDDGWfDLqUk/62bUvagtGeQNMtr5mb2Tt7hspl6W
2jjmNbglT71tsNh/14/b6uwJk/iyzlQtOXx1uTxa1MAQHns1WLIq5vKTWwzD1JXy
YdSb13NkoidQ5hqqP3jUT1bvzVCRqnLiWJxnlaZEuSEwkRUd6VFU7xyKKbYq7ub9
VpEXTV9F2fPI22ADYJxxIjd+STE1wiNN6xOi8fKHgX8aX8Zr9dx+vb3hNv/rxByi
hnhnMXip15sn0aTSUlzbgZ/IAkjHsU/t+VXBPmrWv76Nj7I7fpcl3ENKBAYtMP8R
q0zdeCrLJM+8YUvb3LXNsuP9bmAlNtDPAMod82bhXjxZEfoNZSdGjHYjDigVWboD
vlX98q9SCqQn6Ocgr/pMPGC/QPMA7ugFPBYeqAT1mOlaPdu2KD6SDAWX1LQrR435
yzHFlroE3J7Y88GJF1lveQuLDXmSoPEBhPRAUNSaW4GchhYOOx7tks15zV+UkRyE
QquNHWToiWZrJMpAJ0KX6py2jxTd6fSK/OWNBN73YSEeeKXSAbqpvBmeeILa0zW9
oN73ANEtWZap+ZgeqmoUqnewDYOzkSqwNo/Z9Nic6y49ZoJs4arLZ6u33gcHFYGp
4QZFFBD6E9eaW8SGcG3n+0XcrqjaToEBqqTQk4UPKfk6vEwwzWisqLNUuK1jaXEW
0r67GIygYIHLIaSEPIDbiOCwcFbZRjT8QbcGnKZXJ7o1PE/YSufDZdHHQFt4Pq78
DEfMTPNxwVZE0+AYBOYyrUBlbnQnb9auhyzcwPNeQVI5Fi5fxkxdTdmF0bgM8f8Y
8s22WQI7zpkwFyObnk4koPJLUL69VitNJA3jO5AgBqT03OX7m0GR+JGiWo5rs2YW
fzNUotHBlGVJ49rDaN8N5+SKawneAq1g0daIR5Fuy5uSZjuu7VvPtQZPNvgWjzop
VAuQ65hVd4Sogpqp8DO85Aqe0hJquV1oW6vWtzdMd+EUbUoseXP8ugUl3MGUmTcW
5qShzpPbllpswiPUTib83Txw/kxArFNQGHSzbERo4de9cKXb+5/lEG66QMcgfTPN
b/x4a2ikS8iXXbKIBHl6G2KS5gQvdsrsGL+d6tdh1PWbbcNlqQcTh1VlkVwa98ZU
PZ6K2f6KuRIjcmmha///Fk5mIeY4lJo0OGCIkqsv0/oiJ/JI4YIEmcsCjD271V65
+AomUGf/s5/SQa1ILRiKToD9pIGBcqhLixx/oBRBY1G3YkAoKcY7mukfsjA85jNA
6YfMOo1mSP/e0pMJuusOQZohQjLATfV0ZAjeZZ35Ty0Fy2OF9HtsiVZgj/jY3t3W
nuPefHO9W8W563lzTDZYvWrlHhYBedIjcKcKPrYYVO6/iwPJbQNIkJ1OaX1EDH1w
HrXRWkKEnY/IdY7ejrJs3EedFcuBZ/cPlf8fFDHQy8MNK81skiySr93QPGvenYYA
5qU+fByBRC+6/zCB9Yiw6pUTDw96K0efGZ++UBRZXVno5Ad6v1yf2Pf9OQ5NGs3v
DMkRYnHD36yN+6Ay6aaeCSLLb8YLREtPXCv7KMHOtItDfJck3F9VVypzkbpb6Ef6
8LkhI+8p4CfdeV6s8NnIvEi5Bu0Xo3a983T1SDhMFBonr+rkO1j/Qr9HXJHmwa2Q
8/tJc/lN5YSbpjOLwJ1RN9+SzCwgYALZkf/1UfhunQOt7aH8KXofLZPrggvv0JzH
TBacYSvQnPGTjbF3Q0tSchi2QwoB/xedG3gBszHVudc/wwmuz3LJpx49SZOk1WMc
vNFCexrh7tmLAP7PhUf0bagpaU6e5/DY9kleFd1AHqI4kfHjpiO8m1BOmXEMWw3t
Vlpb3zLXhdlDNzJb0nVFPE7PnbzXm963+ptg7xACC4DgktJoq4euyvEH1qub3yj/
/WIQtYHptT1bFeo/LRGLS4PZQK6yHNl2Tw1B77uCoLgCPgsKa7GlHC1AjYexhTfI
gPZO2YgYQORegIs1LpCLmHTTJalRhu41vWIzjKYw8lew82nOiwDzCa1YwqiqYRHJ
+AbhKZqjrQ5uPyf1EQ0YCBNPhTwEBQEUKX396husH5Oh6sZTe6Be8NtYZp4zYYxA
n8490FupcfFHrp31/cAeBRbc1vIQeyrp00KtrAQVVVCFqn/ZtdNhY0uvMqvQFB9q
8WqJ1R/JCgElY65XFhAAmvr+iaPrrKojWU3JTLWnFfMJKhu3SvF60N5q7rA5eDDx
OAI73ewktmHPkX+BX8BkDstp+AkhhQNmBHL0dOcdDynDcsMVQND9SsuD3n203DQa
twb3Gcr7p02ooqI2EcaZB2HO/ZGavdrZheUv/MQC/D4kyCqFw3SnbJe5QtvulKAO
ebrbJzEIM2nMEK1pdZrnY82oZgq9S4jfd895jDxRPJ2QPHshHP6qCOFts2oQnojM
V6NxeZpPI2OWuzkElyiu0aPjx1SyoF73w8bjZhv7zmef+16kILi8lsfyb9p3igZC
UajhKUKwZ16g4+6sSZtsttdgEEs9noxl9vU2Kiv9UwVxsLk2D4PcP2J5Hfqi+g7P
nj9N8KbfwSufG+k9zfc7bPmUM5asfFtF7zmY3oS8pIlhFWArI+/STajH5Id2zRhf
OftV3hAsnE1tLXHV0svhmFJS3aQE3kLepPr9G8Yzj4A2cL9ZhmABJVECvwWI+INx
53PLxppk2AD8MT3LFctmY3Mn47plfxDfD1BwOzeDVGCfaBbNkkxjc2M9FahFcChv
HnUhfLtNDs+qEP3plyaKlD11ycOGRrg+ngWURHvlcDBUicHmVAXNQ7Gb728Gp44h
xZWwSiYlhHYPMImFzsymJ6/RDm0WYfnDRQnmdgWFUfP4mwrNtu6Ct8LLOy3P7w3b
2+HCBbHSpHraTNeebrXHWFgmijRZJvMeDE4zrR3gi9mnUnW1guq0zFslLvLgwnWK
VfUWZV8B6FUKP0zHAzCSahdvQje4Gvifq/4196n7jtiksiftYwrcioDJv66OSQoK
GXPjag3DMgz1k4zKQSN3RlI9piv4DP+lqy/RxznQix8qQzyW2O7VvSTeVHWBcHr+
4kVIZrXuVJ7nvP5+eTF4oqI3sUKMe1v5D14M8X9loNJfyCZcilWUM1WRzP3tyA9r
k70WuxgVagbjlw7FT9/Ofn8rivL3RtFeBt5ec4r7LzZW65DLWaLDyYFIrgJcNKc3
HBeNcw2rHmGyZdsMqP+AS0qlshPqJ868Br8gif2FXQEZAyAGduMusr88ONX6iOa8
GL3t6eCLDNR0CUe4O5I8T2F8KClAerQcpQXhU1Ramtg4mrHy4+dD7fJRfU5pkwHv
MMyP+J6RMDG6sEJFMFWNTR/y7iitH4y+hh8fRxbqYkFyAhl1vNoB6JcKn26ULLI3
j5BNertIhb356UQYBnNUhLoesA0cd82W9RHI9+lcC9/zBHoIp2aXzNNQaakUuaEO
M309FWbLeqo0dS77Pyy59XjJzvzsPMAwhXzWszZe/YSLTX5ub1O9Nc9QelX7O18m
zJjPNP7vEoP42s1K1Zczo1eZzV6kjSf8HTrZLcSOQTI6x2JTwQKtntln4mtLWNr6
9eIPERigEzYwiHRdjQ0g2U9YTr7tghMtO7qHx1vfz3ywR9+8G4+//0mf82GvKzax
TnumErw02k4DWvHMrp31U3jU6kO85/pNeNw/EWF7mEJGnv/9bekKRo337oC6L+ak
Vr82OqE7W+yWD31J2qOfyxf0mfMSQGT5AV9QFnWlbcl54g2/1IJbqF8/fG1AnYRm
0R4pMD7rBEPAUOt7t14FqDngmFnsrFU1xZzbEHWPki56zGTp8R0X/4R0/btkA3/y
ut2w8AsFB96cM1BiOOcKpFrnc3cb8pcTaJCQviKD0Wb8rI2uMDwMTmwLJayX84Ph
VtQ9G66UHpdaHbQgL/RkcXv+Z6UNfx1Go2JuQH3DGYf8P5zjv+A1KjEKuW+QEcpA
M2b8QfILaA2jMX+WlOgWI9I6AtvRP2TCMiXF7VcL9Vxbrmee2umxoHJ5+JAKPrUF
X8FlJBl0BgCnYfuWH4RhLgHLQV056BHUp3Bu6bNWLvl7BfNJg7HFbkiEkodoJsYo
IjDW5nU2Tp9wxu7zGoMhHmMWpN6DC1SI2BVQMp01O6jueuv854Hpi0r6kAZ9ik/s
JrqZCu2i7ZMNUWbFrTOXMnbof/uHyXU5SfcgM6XSR1Z1O1BkS+kB9bKlsBwaZCAS
A+KnV1KRskYXFl9D2EQKrYxzbG3QJ7BgjVIhKQj5+Gbl/MfmtkNP7Z7ZGAGDM6eT
NiFhDuEeEjqslElSNn42miU8y1tTau8nalgiscvNKznFc/8Fub6LQ6V2tG86J2oD
Xm+Ddqp4o/IsOkHjh0zvjkm2IXN+u87xo7zvGldOP44UFTlNQwLSyBAC9B3Ls5p2
/dtfkQlZwz3rl36XQj2QtTzfuVdq44GAdsr3iHBzsCA6LhSYzyUjwhF3YyUI3ZJo
qwe34Tj1G9g1Ag+vGAeVSwahTlRzyKBeomA/9SmK8sNh/i8UU7q2ivXUIhXij4Jl
1zNIsAk52FDrQFR+x4yCo7FBULeQZpe+5B+Uw+5TKr6E4AOKX8X9LgZdZcQUtfiU
yJw6D0wJT0Kb07+oilX4b3DcFziVvtgcCkf0sGRc7APVg8TDpFvOvIhoxPyDRDa4
se+Kr7AtK3pz7dUIBqfzSQv0u1ooKJoMqDW8mshexFaPoWk/5Z5FLVLAxd6A7inv
WOJNhJ/k3bjvGTJZEV65w3pnEDL8IT4oqqfnoOmYjMD7liFS/Tpi6ObFAM6P+Lzy
pqXUCprL2bg8WOsKzBbjAFZ1Ae3i1XCsi9Mo8RUcKp7gCUQlLBlAnDfWqW4J7KUQ
edP32hN5DSVHfmx43EAGyKgcGsOAhTg5IVfOifL8h78hlTdP0SOETdq4jdvGpdwA
/NL73+K6x28ecNRQOXMrPE2ZI6AFJiQQPCRjeHx42HGXxRh9QG+H8X03pBcOt8qe
WadsxBxCPm4fhBpp2ob3aWHqv0Wx5S0wD3n7ipt3k0DDpOAxVS3FfZZ7AXA2iU/e
eLVT4xLDyPOhZK7CGtw5gbOvf0+S9Y35h+mVBA1ipkoHwcWcqF5887oAHCrOCbQV
fniPEFcMU4oT6AFs8ARgb+UL79CSaAQKIGmDuQUiU6s8q0r2dTWHc+z8dAEYuIuz
GUNgQfwXD3E6eLJ1CZTTZLwfH6Nm/GEzFKtCGmn+wgLswM8hlRSCqYLATO4cRk7f
KtBvDqTeknRNWKdF8rS3e4XfpE2JUyHOwanExmDB5jQ+a3LzmfDHR4QiUj/x6e7c
42bZYrNJgImCLKqkrW3akMlgdG7qLC9fiTq5Otju/K/9+ZMCaKmlClBp3w5mDCaY
A6dpJT5xIyLKE417K/ntA5gFNSia/2MKRz3Rq4//1bGzHoOIAUMdUri8JUefL9DJ
k9URd7v0ZGrM2B94kwT25Z4fSxdArhxQGNnu3ciHy5Mj2/i4Pl7wfGwkPKdRqFru
PkzRdDSMOLdKtI5WpzL6IHOj0HdpAIYxH0TTNfGPr01vUkT5t7Cl0dPFZ3+cli6k
9BYguAcYkTzT6E5ERw0+CMuTEOWqLXkzZ94KRJFTs4WOpHtN9IrnamOzbt6JsvCg
PTi6MiVIpNGIVd1l6vLcXWNGcxmox/q1HVHZZASiTEeOedR/7G0LaET/ZoN/0lqU
omR8poZ9c21GOZ6pmjcwN6ecxViblkWzEVZKcG9nEnUxx9MMU/JX4xxuqEBT7CaE
jWFtrpkcHPoEdR0BxkOGFyIEFYk8h+jV9RiBMwDVh44mhuf+z3GL2R3u4O25mPqp
zVnmQbldKG8//hl00NBixquVukQtwYbXto7RsGGFbB0tk1NkFTQ5SQrTbNkNmErA
9AY2CVwhhD7uTSlaFrV7sv+N4cPpnzg1plvku+xbYlPpEwgYuI+JTmsGfqZczLwi
fkv5GMvux++RZWXe1yxe7JGslX1qstK+UXrIgXl8GLjCMwV+zQjD12M1/aBdY6dL
uUQhR0Irn9ROvfKqCmUvOQS5nFRcDPw6s7OTgTTlUg/5/CEBWKF1xZtA0saDp5xq
1Gvao+9Pw4H06urqXThnp3NEX+HnZgoEP9ouyin7mLjeOrYiSgxevHhs+Y9/Albt
tA8oRPf8JfkJvjALU92IAECvI7oJ08zGsPEr5vq+KfQTWOXQK3qwfcfE52Hh3Mxe
wvYr6QoGwO6mh/poNGpig2IvhSAcGH8ICXMhj3bCr1r+ySN8lW4/noEEWZ6eEpIV
fvt1bkl8elUSOtQpZRTsz/t6ibgQJVgMZhJ1tFHO7w2e6zUQbR33T2IcZdIcG0jV
KSOdL/pLcOHt8eb+fRAcgKBgk4vstSb3I/1yydU7Qs02na7ck7ChYhvxoBzRw5uL
8QvRSf7Mf0u6Whvqr3EQDLIop9DixSv233B32Y1frDcod+D/8SA4PSpNA+lg8W0/
GwA9zQQmwYRljGyy0a5yZ67I4ZxrEM7vWqfkg6OM3eHVAr0xW1L7cKkO+2ltPwyN
b1VlVTf9mTMV+njYuDDHhgGS1gSgD4kwWgLVIE98+WGVJot9JqgVnTz5wo86Qm0g
I/e+uFTE1cqcNWm6hHxRz+BKoOySA5fxn3n7gMpDrzE5RqKX3cATzA15T5iBeUpq
9YhOdU9Sib50OVyvq8IbKVPu2my/tbY0I2CMfMRquRvFkEwBNPkQiintSR7jjxFT
WXZksiBmwWZKVVODMai3lQ20L7TxBavHLtDn5BTMXPbIkgdXLUhy8DwXoyzzfxCE
qA2U7Bgw15lkxtIasvvGL7S4hEGdiSo/IE3I74+o5r36YuoEm5dL5TDKQbheEwzo
dRfcKDz933ygdYrwb2i796iK/OgQQwdiwWVbFHLQu67grv5d9JZQiO67n1LevXn9
ZRMQ1vJfd+G9t2S2UftOE0SD4JRsr61aN99+uqtR3fPJCfl9cUK1IGasDW1OyhpI
oKZcuvw4hALBL5VyWvdT0Z6VIgep6kMOjtMbPBMaKYymhWX35qmZrOmO0J9ZRHE6
dVPVgp2EF3OBWCvCX8qSonKvYz26zRL+WZXb3eyT7aVsM9Rct1rd8oX5pvd+dY/+
/lfAdMbk6+pp+L3b8LoPB+Ca7dzXTJH9KjBwXGZ0Ea1aK/I/nJ8Z/SoCDuQCCGVU
Nu03byjVZbrxzdx/tPfOJgM0QIfL3wrPBfjVkVImpjCXBjhS4d0l+zPT1Oo6O8uZ
0LGrWwZf8DEkhF5FSZlW5xDC4QTCtdr2HwYzg9Cy4oc2HF5ob/wunvicEzrqZgE+
iTALTnTPcxNS1nnuCIE6sbEDg/acVXFwMtlQPdzWlY26iGdPsdPxVnJgfleiPQ6M
sq+bnHjfn+FVMAhyHoBPFQVBuDyByisG/n9d0VGZMAkj/v75h2zcXNkDJd+fKc5K
KV3lmVuI3QVr4Yw7Df+cR/R4XBs3ZBXxRpEJ+Rg9B9xXF/9a2kDmYqLwmW/hHxjA
sR9qeH2xgwe5AKohyP/yt3aZZ96lD0JgobORvJ6kMzQbq51kSkgFhi0TcyLyWqeM
B69nZPUqgFlwBDUlYNxCp2952DKM4eEklm2RwMCLGXOAt2R1zsJnyuRcVnHplRFP
P0kK1S/6TS/KUvVFBuqx0iVJIN73JGyks1BhFcz8qftV7EwVm4vdR+IIvvIzCH7x
AzoAV22HOexHdbQNRT3F9vzHbD0wbsK+jz4Tzf5qezdUYxgyrygG2QvWsQ+lW+Zg
lVC5SoKLSz4zfR0/IAQowp9IVD/7dfxKq1NR2SpUA41bRgnW4meBgApEDf5P4t4r
H7TY61jArLy68fnCvnn21erGDHm5fb7uw0XQeHwk0G/KylSIB4cHpLFP4RFQk0G9
ogbuW8yDQg5ZLAmaGkcLNwXkcSr6fj5hBfhg9paTjiwveegKNdexNmNQiq8/dxdi
ZIKjoAdvLCRutyoXLZYzN07mbY/NwZnmcza5ZhZ+hwAhCQpTn3UHZNzSKqcdbdAr
3jpLVR2viEankKWFFMEwAY+Eg0ILKOAyWzhPVa9bAVn88NPafqz3O9sh3WNsB6KJ
HJSbrrh7eVB3KQBAs84dkayuvzbci4SqW2fcKeMO12L3FLrj4MlAZMr54aSQKhzP
wyAlcBp1L9n3MzP5ghqljDp/vZ4PsxYO44gYUPaXNReej8DmomhpV8VQgrAq0Brz
veaBpW9RPGerVUnjV65sMbuZC0Qm1qte0rdk73BBV41VsqCccaaxOXXI/thA2Wep
b5uI22KswDlUSqId2kKfZoIA0r4PYOLWhF/X9Jorzm9FLi3TrKFgW41z1syLeWbz
Txjs2IvIaIKjTlMC5GP0hBMCiPZmWkDGY92MtIg3h9J2xoBGUF8ZUYWiHxYHf5EW
cL4+DEEs+nrVJkAE3VpT9dneEvunqDZY1KiwNkO/ikodj8FOnmKfuWCmcyQK/O5X
+Cea85ZyonlXY76U5Rh2KU0iR/wEQHYO+uo4+ewp7ge0J9UVlL14Fe6jO8lU2K56
xO4MCk/xKdnIrzUXmfRjRPpHZLRaOL84DQhG8O9mCkFTMJB956+PSxG4zqF13KU+
Qi6geHL2Ky93zp9NtFSyb9/23YLLe/L/ECc95rdltXY9YpIUL0Gryj1gbWLVDpTO
LahqkF/17ATjHph+LoKGFqCSJ/Yibbkhr6nscaP7LJwi5SUDnB19IwJrmG7Z24hI
pjRJSeW9i02BGuaACPNEcmplC+CkRmbveqfvsDM0ckW4ahpyrbP7DQkJljw7BpUh
hOvewXwmagPgNZBwyQr1fDyGviPuSXABjns8CU+r0MNxAypQDeU7aKnUgWhWE4hc
waAiG3o7Z+aPJJYQak9dolbd4iXWMP2lF2NYOlbB6mUotUYRVfVB7qOeAaEeG1Lh
XmMs79BY94iQrrEa9Q7fY067/ZdMXS65wewZk0PULMPBu3+ZGzkwlabSuMs8wSP8
Cr+MqWS3HNGeKYFKfoRGss6IB/K+j82FwJbyyE5BiulNTNVRA0WySdIoEh7ITD3S
aMxE/7nwVHy7hAutritpwJfA+tgU8EF3C6lTKJhki0rUtnh/FGKjyrhTSatha65Q
65C1j4q5GuD0Mgkb1nIPUqBdiEhpA1i/OruOL2L+XAY0Se255qPcZbkbAjcXEmxh
8siqTgMPvU7uIaSBrCNq3mYXiwlVZ07sBtNQdNbnxd3kCBGDO1uxSW7JFtm6+P2G
vTBurrKQ1ZAurN8jA5XMgPppiIs23yjZicIKvDdTVSc/8Jyyif4i48ziR6vy1zRw
GW2cTasniES3V2jRth/5PTTL/1z8oUQqxQlM0DlLD1BQQleB103VaX23vihdqhB2
uP6bEOq97YId8g76iUlCgUnJ4ONnxvMVQomrAzEI/XYhKHW5cGgNYvn4Zm99CNkl
Hs6L2Ci+udIxdVRIIDvvhrD0RNYtI4XVJaLlBBtdnKInL6M1yXwp0jRWo6k4rba+
v5/+2FyoTpARdMG9RpWxgokHPSNHtAXu4vL4iKbEOWWcOlseRZTZBax8oJaA6Zcp
lDmHRKbjk/gKLBYzJPWdHaVRwIy1uKQ2v3O+R0jF1Iu0jZlnBHeUsAa8loy3xAoE
eIQO3f2wqANgVSu/Ik0FJ3uJ4fxovrk8RASliEyiqTvw47TaZJtg6BO5HFhnyL/F
By1RE1B7g/9DgaatOQ8EILnbwqvnRd1w5An7iZmSk9KNcNOl+CW08WDhPwOwJm6h
Ld7Gv/xaHjus0b2ZZQVJIjxD0MKDt2ctKLCyYr8q18+x/ygJU8CAJTH2oNi8P/Un
WirUqIsqwVGTNktfYP4mH8tNNwZlZb+1roIBcV4H3Nid7FMQMnQyzTuD9dg1oc9t
2s+Ep7arWndbYV6YA5z48pH7t2FqtNy8NzQM08cH2ItkJJfhSZA7H/pwwosIoBL6
hWoxm263PIzDjWGiDDyLjLfFYA4DW4dWVRUz0PFNBIgvqw4BVXvJrKPouyP6QLrE
INnrlRzEeOAnsKH836ELPAAc4t+faUyce04eUHCHxDR6HW1DwEGz9hPIYoWpeu5m
vWszKbmqoyWtRixzmmdYXDT8lST+0XNEOyDQMFbJwsUGIXDIcgwon4K+NK2wmEo4
c26fjqbXbttZZr+8Xy0zOx0nmza6x6swqz9tXI6yhCizjWXsJY+lpmamGszdMjSc
pSrKIXf81hBDvpmL1IdLaUmvB2cnEMHxo/dlRuNcPHdvQ4lnHGVr2io7HpttYfx3
5UXvV14ZbRLmHyiNM/LDAnUjPbvFvO1PnqHisurmwuBkX7D/chWAn2TMYSqOfPHd
cNzHJ9nN0q6u1dZ/PFBKFZ8ZxoAVA2g03YpG+35p6dpVp90MDfPZ/KEnx0P8Rwv1
HEcQswcD6dWysPXphbGxae0Gzxe3H8vsyY0nAhTYp+Kro6r2S7Y2snipz1nYfsgI
FnUt/oCChs3RZaLoCd4qCLMiMouKkwM/GeiolmFbJRhy9ZN6S1/IbWy5mP9UjUgh
blUMJSr5MHchDVeZkR7jKF1FDXPMBStUzU0F4dG1OMYWe7gCjNapjMwxmUywuJU6
vpsVrOPOFL3EOWpMIWMPOckRHx7jx0+Vh+NynXGr+3rSIROhGl4FoRtyWa7hu33C
Ofb75IBdyPYrpkFt9l1FrHdzOm35LSgt5XN59N7UqDdWxp9AcD0WeJ66t8YyI25T
GW1D5Z/sj84MhfLScEOlKAWcJoU0c4mEFWOmGvnxw3a38UtYchVtnC9nQ+Tu3MG6
WB9iaYtwvZFPhlDmuCKlJDEekfJ10UrNzqgL/p9T396FXQn98iWNtVcJIwsMgjUx
u8AhetqTDNaMOENmqF9ZsKe9G1jiyTfD+vosTVBTzoYj1IizZkr1BerulKuEOvmC
/64FPmLSp0lqRu9g0PUja2SNGe61EeQpYYqZE8hWY6JFzFgumaebaPvh0Y40os9w
Ik5rP/lKZX9aZIRkQ1dMyYpSwIwcH3MhgS9cAAcndK/z+lnV19OhRNuUTNb0lRGd
mXU4rSCnFXSPZldYGxvxzMsFlyhKZBBxgVF8nWtxA1Y0YfOtXQcDuoLhgEOB11DS
/wQIcqw8kTs16rfUPqAVhSDiyJ2xtZqLa4gsRKRdYA7/c4Zbxz42+14Z06y15YvV
mPNdySal4jNX+w95cbDMT109C9zN1iLPpvQbVNZ/dHs97YyghtT82r15ConaNGC0
yzn1PqQ6qNSLSdq8u3IMRk2Gk8S80kJGWZ9vPvES4D66O/WTyfKD2uXSjdkw5ZiX
BPUHGJ+Ntk8VUNmJOFhXPW6HH+bDgdCrAtX750Tadf2G/wuCKDhwTq4WaYcxRnxo
VHePhRPiDy62jYDfz7CyPqOL3TQKFq8s+hnpZ9FxslRuDCgqcy27W3Ymc56lo9YW
M7vWYfuhQ+xb3tZ1aNVZ3Iilwcogj5Cz2Ooes5+zI7nfARFYmEUgqMFB0UGCtu2I
wN6oEKqWVe9bhMrQGUSfmlHz8gRaJ3hxMraXFEqMyXJV272dd8Sl+/hgTqfKTamu
ocMXpmfqDpm+EjQKtA2k62J+sFjlIp6LY/Sq0X/UB2pd4haYi35YCegC7l6c1JGv
rQ4vE3VqxKI0yqh5900ZdovG/Pr91QSeNXJM2OryXWdo03qDaLTklTDqSrW6qtSi
2r32oSXLvjaM2eDmAWwitchzeSOlcqdCSSo+qz8k5f8K+o2XEyYfVop9x+LkWr2s
w9VPtRd6AGpg1cdnlMOc+QVZX9irvw2ON5IJmHAQsMn/3seGmuQDD0JiIJsteDcq
cpd+XifcVqTwVOQGO7CCRPCBGbIn7jX76Kv9pzCiHDn6yGORLRVgmox6vGXFi7tB
RSa9FgeRimP+OLhhs7oEOX8lMoqrKk8Mk7WgbNWyyNA8EXX6axMAbv0yVMjpoV3G
XV+DLU1kXHmtPr9aCiC/MG/ZJMe7C/XHghyFEfrGsiYqD/ucYa3P1VlGzceDtyMO
FvFu61ZkbwMbuXucMRit1Y1t1hg4RpnhHYnOA+xsmX4mY6XzZyGrkrZOdepPPtB1
4/HTNHt7TI4+4EfY9uuHqZjv4Hb0kFxj8RWAF8x+H2M+kMA2YcMrTYdPdJEex1X1
0F8sdCK0uEOfsfigm/SzTA==
--pragma protect end_data_block
--pragma protect digest_block
GCuDsSfs+2eRjhO8GGWER2RcYaE=
--pragma protect end_digest_block
--pragma protect end_protected
