-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hf+CwjpuFtUYBrtTH9T27MXZY05ExokIB0tdq0TbTACZU6rsL4QkVTgiEQXvEDWuf2m+U4u2rqXQ
JkeHQ0CCb8D5ZL25nKfLtp9qa61HBJnaiXoo42sa4a798GZ+P/EFPI0XNOVKsyEXrD7/8GmJobXA
6979MdjCCtLGBhtuIL8OGQ9ZaRPwNbDzE8To/5yCu2Z2YQ01LBn5zIyfAuVFLI68g1Kd0zd0SQXz
I2+Xr5Z4GAaTCiNm0ZQnQvXIKPWc1tIXaz3277EWVEq0TGO0qSp2TR6cdyQykjMkUV5ntPOr2n4n
D5c8UfuHiT5Iq/rD1m9fh5oBlQjLXBe10h3cZw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4832)
`protect data_block
sUGN15nd9IQy6qmcj6qvRzEl5VA9w5XZWg9Vof8miP5j1l2n86kjVWqw7S2PhtDKoEO9ZmMLiRFW
XyApsKujM8s9iuPyji/duSr+uruJGEnJn57zGF3RCgfbqBxayu1Va0mozwJBe9drfPrPF3sBivcZ
6vTwwvqnHZKdFPpOwzjeEtmhlcaIxYV0nJt/Ssfpmn0dv65mKAUlRv6ceiqqrSum+o5nz7SX38I7
UTrOSOoKcFPiDdrPWT9aRttsg6HLSYEYLdApIyd8wVQ1J15DR6zlSej/2ESUsoqcv7ID6q8TkiNT
WC3Xx/DOcfDf5p2XuoX+upmCC0G1dqd/M7GlW9CN0nskAzmVdm9uj5jMekH3I14SdkZfz6ykPDFU
7W+gMYcqQylj4IBwKQiyyVZJachECe6F8RZlqwVap/SEotNQqYM6evNdVT6hPBgXeRpCC67CFB6U
cPhMDnaXsLIkcwWhx8AxiUBGKTBFEgaHvUa+BrVCfEiU+rMF3JjDz9Wei7RNuaUBuszKoPHGVgAE
427oCjRMQSvY9oslxv9dQWE80Jz6//dpaUig6Bz6MY+u1djGvpm4g7Z8zMxxlT6H0Z0iwhgcBPzG
BsxM/37L8oS64pccnEgBWFXahORrff4AflB2NqjueUxbYb1RfDWFZRJoEKpcAcjl/Azkh0/UquJd
ekeQYUb76FwThJhBm2S769tBDvN9rN1BiPfD1cXmmauQsa+K0psIzRDnBR2QfyUHwvCoHp9RK5b3
CPUdSPY1iaS/UEtkTvDxdee1WSHU6dgdLPzWOYfLMgUB3oVVwhGWtTfFY0adIm9xkFgaVxSY/5gS
JFVsj8eDzzWjO3GdTOEUYONm499Nz7jpvkRlDjalsCDVYurG6MdDXj8aM37GH+IQ2oqlGuH160SI
nXdfXld2xDYBVBMSQHyr1yYNC57vgGwG1HwZnycCa0X1JLomzCpJBS4mGUD7N+9h11n/C7fCwan4
H7X0Kj6hfqtfnF4kgyVtVaDe7QVQlfzYi0nxuHGKm3Trszu/Cqt3LmhLH8NkCufnrLM0M82xJ3QL
7jDy/eD84LXID2iwZgrqJJCE7H1JguWzZHBHfnOwpb0vWlqOc10XkrT7/BBCr/YRkOGJRdDfy+OI
1L6kQPRFZRZWLXTztJFZtWqZVs6V4nD/1yBODGOGtIJHfPcSuU9WAZOQ1V3W1zXGKZbIo9A00SZV
4jsHi1g4w8CeVavYZvD3J0bEPTUqDKj4yHI4tlho+qonrr9DKpo0De4SP7M255lTDac3GJONE4oi
JCC1EvLhdNBmQ0Z6BBgikEjpCfiA4kXnvBgfpwbyojRXVZl13KpioBxQaPaU1L5SgDIOeK3sKmkB
MeUj8VzsZmnGbXcVNYJJBLVIYIimhI8JpJaq72Ra9A3gfHMGcDRaUC99F4IxTgOE72M4EPHQTzX1
75UMiYex6Y+sX6JdejAiClT9aEsipFCjTrFkghoeMqZGhuTzzQi7MwWcnbHHxK4AqHudFfyWXTU9
dChE4lVdrnIp/94tmnu5YXBZerr3Mi+avxo1az3R+Ld0L7eBEI/hlWP50LstwAWIUZdFL/tJj259
OoXWJ92nLUZOLzBbPTJ+QS4NffHLUQoZc/AoFDLM5b+gf3HZ0Q3kf91dFNMJv25f/PNX1lcxLLvI
hrdKLnCSzOJ834b19aR4cRJTtMRU+y/SQw4WMwWM/ZzbeUYH1Xugf3rGR5bs9RNU0LLhxHnuhk9c
nO/nVsjIFJp1veD09FIz2+LT0PsFO+JveMCYLL9XMu5XP6U9c0U62vu3pp0IpFcZ5eyE8nLDUgDJ
dncTWlWdGp/4cu90qqjwoSW+atffZzCjzKwY3MOaXQpuDtXWG7BfBd69O8CPmW02+vAJf0n5tUe1
zsaWH/XBq3lMlqu5f3BRQBKwZGSdnbNXA0qr7VH2kUPqr6VeVNPzG2rncPwL449qDDW7/GHSVdQW
cLAfgvUfCwcSOJknciVhpjdXl+zNFwx8dTPzxu6B7yItKTJlQnP4WgdO3bub4N6H2X3v/91T75AK
Opnbwkbln2xFyWcTkaB1ldEjGzZU9WtIdjr2ukbpaI2PtN3tvrnuxSU8H+2taJj0LZEmrR/txs8X
dP8HfnAUdoE83hyHpCb9yAzL94Kf4JGrNjr9aob1/ytMWlYVZQaaWr/UenYHx6vWjem9R1idNZBi
Of2GmHqqS2uE2VDJnfl1sLXwkTmm4QjQMztvYt7tIPlGSsEqdUX7xLIRBsv2eFg1BzXwhwEKAn7+
4UWIzrEZD8lmDhlthZZbzUdJ/9BEiKUSFNCA3jCYUgSpNDFiTIBIJ51IGz9+37XvSzCG0LsBwj+M
caKeTS+q2bQ3oE06byidTUck37yX+sPB/AnLHyikIDirCm3DcqVY1BirO+RtJJkdUQA+iX8UucSD
oNxwHUMG6uJGcV+pOq5sA1NycCRryWeU6X8YjqNqBH+YNgTjMfwpK9bvQPv0X8n+fDzry5b8czdv
fROtCCI+r6gKjLE99vD4pZzm1BTY+fSYV/2z7atWM0F2fceNck46y8xX8aZKOIElK9yMyJm37z+6
MUtKo18g2FSGJRblzBFWjwAbb1hoMZ4EV+XYClqaWVXeNOmdGM6sM2CpE5Ala9o5aWfbYis7S0SF
yJs+tlBVIZ0QwPb9w44sz4EwlyfFvKUMOsxxtTpJsdk05POJY88aCw9RLWI/7UqgqeWGI9e3xD2b
PpzlEnJwOe6KD4Otv9HLM14N8stFf6CXDLkrOGpoiSXY4YFD2Iz4nIVTLtVFUuH/L/PA2vDIn2fc
y6GfJ3KyIRWty+2gSODuz5/6k19rjrOSJnNgvNngX4LWukjyto0WVnsyOuRnXTNPrqQ4lRSDaO/y
6VIHYFUNwx/NgOZZny5IYlCxx+2IaL4dr7TO+dJIwOnMUILD7urEuJLx6zO9JQzKs9c0sAb1+pCY
OtYf9DcOegIa2zBlmyIFZqeJJXHMWe/kp3znlpXxp9748XoJ03M2w4VIVefyCrzNXQe4j6P6z9JZ
o7222ddkltJ4tnhi4Rm0croSiyJBNsjXNWXH6EM7yC3D2sW7io8d8U9MHZEAS1Lt9bQlOJ5LlsJL
K1DNek+Ux9YpSe+4yCv1R9RYCCVKkfwliAfV52HrIDC4sBaDUZ6t6j5rc1GUkNkU/W8xFIpvuFvj
5YOlA8e9ulxMVzoHwaKEE9KeqgNURS04yiSkauUsZrV5E7VwBa6MgzM6kjFgpzGVc5CKPtLDmRg9
IOMLI/bg10xXrk627jWqz34r4mo/BS4BjCJjsiIXEnlsZBo9mzkaeOpJtaMh2L0NhqxBg+JKyXH1
t0z3afadz2a7qX7Bv1bILjZtiufp8NyriNpldk6BI7ZeXv6hi/4NcK+S74gJvMo/KqrzA+JcL5js
glcybgMYh46ZXVXFc4gGYBt1pHYHGHOj26Qifpw7NIlfaGMOY3P9Q5T5Bu9Eyax/YvFHQ/Nswd83
XcPfQsxQKEALtDb583cuA/g5Sax+0DdOq8H08ZUP8A8meuf0AxEwOQy+mOK27OR6BvBwXSGGSXvP
GLkph4iRiEWInYp/aSvC7OLzaprZp+/BJ5nytNSgJOUeNfoFeZ2G/xMyy4iMQ79YE+lz2YXtOS7u
GXQPhTtQqISMXF/fuOtuyKZIhCjD+/1TccloTg0YyskYnlG1uTE1DEPrAulEyzZt3d3aA3bT/Wxh
rnYhxt77+baYSHPIG5SK9a7wA0AUNw9ustQ4ptPH3PcVYgbZIR1tb2XC9buhXmz2YaV+yhsqOK2j
QEVKBpG3TIbToVG4M1GQ4IYonCVtoPnJVflBq8nFwi7QYiX7xvIpBikBmt/qT64goRxrcWpcihPj
l6zC2ODRB/2y/kkt3hK5LJtxR4GXYRyhC3t4qVNOpYkK9xudSlE78CIjsUHx9ht6f8nzeuEZRtFj
1ewg2KqYXnkj+R2aUuZV/T48RHJrCgGhVUzY+aT8R3qPEbCziXyUGK2XDz8GsOTm3L6d8LI5Hb/7
YbyxxNDHJP+uA3Wbm0KDek9FWA3fMfF+QG4RHNtq9OgWRFJxJCUpkg8u02Mhrz3HXYI0YjT9aAXR
ez3EKHNVd9usRy4FavC82PI6XQjbNOGPal4GeuUlYXT1EJl+4wtRp3glr+kQ/ruh/TroS9rybTAJ
YvTj6ZtnxRAbnuP7wjwAaqqwuTb4w8sG8+xYJ3XU4oXP1S9v/TbFq4jp615CXDWDeesgfHIGnF4Z
e82/1KfO9ed6vQEgZvxtBBMXrB9T4vXQZz8iu7PHPJciiLnoKqQyNo4VKT4c1cdSULyZbMpUfTXS
kaNmqhCyeScskjDr85WepyS7dE/AleIJ9WuOtkHO3dWLJNsn9IYbBSXzjKZkUmtlNeVRDbII4B7b
rV+PfS5A1FsbVOWNHyodcY4o998YTSQKKDWlUTU5YE8ikwwAZNAH1B0nRRCTjuUkrptcYvv030F4
uYVC5nBzq5WqyNbo4XjR7K1/V1rS/1ToRRLTJJM5/n0jYOm/RIh7/SLWJfMtABfRRDCnl0ot+Tcc
jBU/rS5VldcRhjrMV2SQMs/FyJLD6wpmfO+KU3CDSUqqUC+GrN5U9vwZOyqelXrdBnQcrPCy2uDK
bF2EPfs9nw+CrAYSz9FMifa59sR8s7UQ6z9mDuPfv8Mj76+d90pkDLzUasFAjiZkwwW1GJdbEO1A
IyZu9o3BLDTnknYQtPzXT4LlaH2HAOPd95HuUwazoMnozwpX5dgZ3xyJdagrNfHiAEwkvv4CDQOy
5OZkKV5BlaVx4TMPTTPcsRTBZDY1pCi8jqBMwXP+Zt8DK8E/i9RFkAPKfWXtSvjML4f2yg4qa/4p
q3lGrwfye3bVW97e/OruFBHKn1ZuMPJC+cgJHD9ZFWdhP3J7/6UCvZYljgM72PT2EkFztHK0U197
vq1S0H4x/umNLuJe/gzeN4L3ABf3ZjYp93aPMHQduvz+b2LDTKU6mlpeYw6bCNH3YHX94/KexBRu
u32vJIZAeNJyCMEiZI0wItfvdO6Hkan3QOpgDf768QfxjnRw1aUxt6ZRBQMkW8IC0TkCRLP6pU8/
aHdzVbi0jljG+IYXQVFMks9CgmpwA8Mnj9DIZfWQqjGl5Qym3MQmzgI5VCh5YtF/gxCcGvRgxBf6
gdIxy2SWt27XqECo0MMuLiEl7b/gTYN4+PEatXceQ6zj0SH2Oun8aAYAmFt6BANh1jEcI7ZhSiGm
XQtYIFCisvB95pW+X4doj3hVY8DWbjE7BitKbiDG0ZBK8S2ve4OS11Maf/ujsa3QNsCKiuj0jWFx
S21lIQ1hAKTmSt7cYSc9dsdpi7tb6mwko1FYBEIUzFxJx6gJYeOmiYNigI8V/hLYI8HkDPnwbWD/
WuhWJn8ohjeXornshlH+vX/bG1tfkmhc8/GsbGsfTJExf9LjPZTZHDRGwGldotAosJDV4IdtBn7m
2j3wHDibGhleqGVK3/TXXX37+oze5u4NaEANobgROfwk7meF88/4prhl7x5trybAKGEx0ErbtkyL
LroQDhziYiApWyqfiy11jAWwSYU0Bw674nymNw7uBBwlwNrTvDayrHJC5Dq5pR99SjSGdxYs0VR7
EGirAG68Sl2q1pQhvX46P431KPmvnYTX4R8dKJ1zdF+nTSoFQCVapqjNF+MOLYQ/JHVoNuezBbxw
XkmvNgNsWFK38oLjoApDPW0Y9VjJRKShbLGdwGbq9VUF29SMm8x8OahTKN5PA13KMLvuzgcMctAI
WZUKP85EklZwq1bvKx0wg7GyR1WsJtIkEF8W3Og3cC5lsY0bpapv2h0xTXO9koGQliaTpjJBdkiA
pSUj50oK9X7+fV/dFze5/jIi0SvkcFkEtguCcBWHiz+Mn/CneVTjSKe/Um8A6m+lIs4qeKkK2z4n
SOuucz3FFof48tai6XZlKVro6NxWTbBz+Z2fGWyWluzWyXxguL7wqQFJmwpJhiYDGoL05rsMk26l
2EHDZHT6lKJuyRT1hoWX4oIM7xVdi2sef37JuxF9NyCSStVBRjlWnPBbrFsJxuPUl5YPZuB0i8uE
IBVp5xyxIppKpUekjPrah55LygpVRJ3PV8+pHGUvGYWui6Ecr1IGSPBTf3ksMqkU22jtGzFpAadt
EHCrislg1sPOxMPWGTglzLcgdH9I+m+2rnpnh52sJg5KJgFTXQBuv0qYCgUWApar0DgsAP/eBK1C
6MGqgIVbSXir18LVPg0l/HiTfrwrqZjz5vUF+mbE+n91FRaA1/Mcy0btFoZ1tCGtIZr+rJQb8x7m
RBeTVURoeuahDZXfHnr1KOiOO9LoWhBhnSWpMIG/f7iKBgTUvS27euwhJt2z4Clk7YGi5ABwlFGP
J60dyM5RxEzjB8iaWdplKSvMxOyYc9mnkTmYb0SE2t/PH1qziUOrBJOTVO0=
`protect end_protected
