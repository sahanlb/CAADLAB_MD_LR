-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
V+3VT1rtXmKJegc6VIIgOk4momY62J3uHz942E2UlLukXVXPB5GQJioh1SpFadi1
52jFFFx6hrP9aAN1SsX9MCEXyuWnVHchFbhP/1Y5caGVbGgzd9TKz5peOQU7XgXW
153XgrZl1Zmzb2FraNE+rgAkbCt7XeIvujd+ROt8iMQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5144)

`protect DATA_BLOCK
hO2cCl9oIPUZmJrpOIkQP72GmLIf9s/TBon5Xpu+L8cIAzwfC/YTHcq56okJDMvY
S6ckXPbEJ/iCTpdTo30cSnAZDQ0muiQnLEpuhjpmmprX7WmgxCZVTJJMMxbDlv1I
9TslNapy2jxxG9o56oXQLiEZn09+Px4ExtU0fMmO+w/Gz6wvInVog2EK1LV3LVcO
be+aTv7K2rrlzQoLRCKyaoE7AK9VgwqcVNKY2DsGA7ESIlT+KIa7fUbiETeE9KeU
d9LeCByrJ5VsiqgVHWa0+D4cwtH/W2/WhHRQTIlWx/6KzPmXDzCVMb8jGQT0Rbwn
ZRnhCXZjFxrzEDYmecPuMa/wPfS3yq5ekpTy8lqnHloNzandYdV7bbec3M8V1SK3
Ka5kB4AobORx7ejXyqID4X6cpOA5L+BsPJcO31fTTdXdlsIvVfFqvWa0CqOv/ujB
YiLZ7jKY47hHv92BOjySsRWLJOunAXGoHgC5TD6VrBh9A59pzxcqbIHwmK2Ix8qJ
U5n4SNn5E9bituu1o+cZC3t2JqOtIhf5sNUcRuoLHOyXBBpoBzZg9HFV+a0YbR2Y
SpWJZV83QghPJQbzTSj/EmgmlpO86PKTOzp6iLZQ5a3+TZZKTA2NA9GFGZ29roTK
IHeh40grA7rimCyJ25HeJhBuP5SaZQxNRp9HWQvFoIjZoOI0V5BjeeH+hg8Htcjk
3Qiy2y78jMAQdstlVPbQF1kDpSpKPNDzwQYp3Rxv0DpufmMpGS5yywE5SSgXItL9
PKxxLh6JQWQCktUv7l5GzbWQaSfRtpScBm+A3PzMMFRF60zI5LGiAeCEFl9XhNEV
M46YBRjbFfDldh4jXhKeQX9sFmTP/cLgJHAz1J8KBLFCPNsKl2bUPZ1HsDFN1Faw
CA2Vi2d7Z5rUB/yt7/ToRsgsG41Z/xXiqIgm+bCDrSmE9pQt/70HJeMBKjfHQSD+
KmEJwKLy4SmX7CXwgtw+QeWLeR8FaXHmlbK5CHfv5HaOIIiC4wDjRjiaqdIW8m3s
colTfctoaaISaB6sfIBIyNEM5DzuyidXWFoKPJLbE4P2YCrEXfzQTZSMEd0SINGe
AswRGFrag1x4c6Hj7VCQUUP34+KkajowLuq7OH+I96X1yoGVGmFRI1iaBIsavYRt
hfs/Cv79zZC3p8uJ7XYCCmDxWaLC3sf/mPQGfg+g0gnAHsy22t/aVKq+yYWf2iOV
7Qh8GdycjsF+XfXbXyTmigzZAeAU7XH13FyYmJ2FIhX1YxrTEO1I/i2wHU0ZE5c2
JBp95Q920zAmIypY1clKsfjkbIDtNaIWkuqg9fWWYrL0mIxJy0dRDwH+tyymcfsN
ZdTSWIlUjknDxr7tTzEuNxyr/30ODNg1JPOt5m19YJOvCli2AaUvntwIFO1GgITM
flNUCYRWo4+pgtLJqRX0BAIAuuPgUJ74FWcTvkerpbemsIQamnO0jQHCQebPT6bB
LTza4/Ui6c8YH1ww0j5x6nyLlSSPrU9LfRS5tGNzAxwVk2MZOHvQCxLcsYd43zVr
lrN52MpoVZtvmU13VaJeuVDDvt9jfDYZFxzYdhNItIuyrb+XNGRFsO3215dFkg+g
bJzfYmMXR9BH3dEuh6DmdTI3Y8Wtx/NMToN32um/iWCEKwcvVQ1GJ6HcCh1ScXuH
dgdlifvBj7IHA8SeqhDQU4zXh3qsQRTml2hodEN3RXl8rrhdG57YvektjeGdxgVQ
C7MEDlUYPrdt5O57hQ0oqOkuWnE+NH0YdPFE4EfFUdC4v1Q5nvYIisIHK87ATk5G
K37m2P1mOX2oMD8O01IPuFb3jSKnniPMgWp8Cv72c6VsATYujccQ4WdCCLp6Cyy5
UY45nkdszz17efyyU/ogLRTFKpPz0tGjCnt71XJfi5d9+bYMtRFn7qC/0Q5eidhz
B2DswDWAyFvvpx8FFn1a76w4HqC0HUHyNnK3/UGNlG0YyBmjGRM7uFt1STxGpwGm
AOpYGKKVgeKqjNfzCtV5LuOIY6tjvFqnctzxTcTtS5fvH8udysFGcoVhE4j6b9HK
KIKGip6VeqKD1iUBlBdwom0Kj25RJcmo689M6HPkQVGL/6nWJgKzywEeWVnC5aCy
Z93xI2a1Jr1xHYDwG1NPD0j1UiYubUDCmH4RwkTxBMcGthVj/9fJYvKMazlCNG+s
4Tr+7Xj3TrOSJZzABvSlXfi4NVdD6ZamgLlnfUMO0foB4DZQFB5hi9na236gnnsW
JhRH0+3EUeld1u9RsnxmQaCc+oHjXvtbGDj0WCT6zTQlnnxYfc8FeXkc9de0/udX
e5FaF+tw0LK18NIe3LyMdY6+F4GEGReEcnQSQb+hSzHLzD+Esj9RP2cpcrsMk2yP
BW2DZBY38fyhuLsW2M0dlX7ieIBkc9sMPpdnwYzXiKDyg2r14PQ+IBe+Pxv1NIOj
LUGM12CDZryNuZW2MG5sDbQxgRU0D4Ltrm5A7Y+sV7lTSl/aJxQ1LK/hf928o6+c
rg+O+QSWlu55nzRIvJ3y/P7aDg6u0wK6iSUXNlVkASq9fbZF27qKftrbM+t1aHLb
IJALS1/vrLQyXawNfJPDoqxrcJTYuH1DPMtTb5LshSwIgaOwu2pKVDVjzeGZb5+q
Ltq30gkXmRTfXFOMgdZiu7hCknZi3Hm+tYd5oGYflsHUTwXyh86bi3KRO/web02n
mAQ018ZTxsRa0N+C1BHDdOke3ZMK04POKYKT8aNmbE2WGa60rqhRV1FEm7LHveuD
1IbxXVa2hKSFsK3MOJR0ee9HjFIraAkkzOrm+4UwygoQKL7oRQvjTdUcIJ0t1HYb
t2DbSL0AolivSLZsLRGyQPpX/2g4yNLR0EbO/rvWJ+EP87ZLWPLpe4qm9+l68lz/
5Su/ffuJA+pDVyUYSjPB1PCb8nDrkGPN6gOVnX9w6jg/gqhPAMeKCN7eN1EuiylO
L2rKaHnJFvU2TF6W9vmslR9DwErXXw25wS2rf5YZ2WQBdCsDFsyT2tXZ/CNBTPMb
0DIZmjpqPSPUlSeAHCAGAQerSY7xtEz/k+oiY2mEfWGCm3yeJfdE7FYakbZoSuFm
nyRbnSY+cMt2ZyPKUvu1T8jqY4dd+GWqC0rZpSfymy+e2g0cwXKPJJfzZ/nzf2q8
+7HEdRi+xe5nEHe7iEG22XOlvmHUcTwlL0g9dOuHHfOejayy8jvKK5Im7OKRXDPH
ySJugEPic6qVXSa5AG3AU2KffIPC2B86UEJSNffIIsqKOOTS54Sw+p5WQ52f6BPy
e9DooC1udmnqWG4I8B/bkPt7URH/D1ogx1NQ5qfAYMM+43GGXFIJtb2kXvKUpdqz
ptW9hHlDg+g+pePANaQsVCBfsrcf1xxYZtQSZnjWCfhLV5k9JmyraqxT35brr2e7
wbP6c8ZbbWGxikkaTXvkBAY2dEPXL8H8RYDF49eU2x8PuMvDOuX9enUcUQjJChty
3gmgGU64F0CIh55ECcibplpjaMrG+Hf/mDUNOFD0wEDDEusWaq882H5L95H9ViJ5
URmYwGrdJx6D6boFrtRq9g2IqgfHXZjCYAbN8Pau5sX44nEMf6fA+XvEXhlruL6K
Nai5MWT8h4ODEJ/N+/EgR1xg0S+AgO29UdLuOu826o6buYYS7KPjr93lijON6Wew
Pov15yH4GndJKySebWT3iCyZa9X9npVNgFVQyeehK6JQBQ3IwrtjyJbKAY00FCBM
+0yhnvQiBHbo88dc87io650DBjdf/btWznH6KE0vcqAvGNA/OoKS1P566mBWDh7O
i6DRGyuAEbkgNC52IcIjP8nXaanAu15GahvNoZH0UzXDoJUGtHKqiYDlLixbWEii
tFUhwzUG9M92KI6IRH4AVPUNm9F/FsZRaQiVMoSpkk+kxYvqbT3NuS90GMBjij9B
Fi9FlUNfqKvYZUyyYplLreXJX9JYDaRcKPwrzaoDKj7KusR6WHeUZ6TIdBnQnv/K
7zSBxeEmdMNroP6hGmZKnt53aWs9aeLiBNPDDJfr1PVmxMRwJDVwR7ExAJVccHVg
6ok8Tw+2m6ixnfnIkMVi1OkmAaWlQbSLYcd7k+nvZsgD8xX1Q8VBlwuikEA2/AqC
hGtQr0E+iM9gqWI63T37jne8aKMADiWl7HhHSrLEx7nHvCBAvFnWnQUkQrJ4APOc
jwwhTJ59Kav9FTXGJtasi6NnHzjBei4I9Ch3dSEaofPLyh1TmGSRDvnRVylbhaOd
GXGbc6OV5hTAADiVjNWbM7Xs9KFXkQ96+8lb1PokdbA/KivlLa3OIeRK6odJobhs
sHbv4YznMCZTgOOBdEIjxPT8G1xr9toKhGYz0U20plS2EuVI/sMqUInS/2b95Q6d
WZj8KtGZ3ziTJ3QRRx8nD8tVlFD3aZtwKb1m2TZsoyOnVvCimzCbAjDLMWROHBCY
3bbttmmqciIZVU8nm7LwTabHI/6OrXgvaA3FkoU9xACAa92a5g2K94Nzq/CmIRSU
7twI4/6wHg3ZjVS35RzXSu098EAdcMh+POCM0EAKXHNqIeWujjpIr9vX/0Oz2rs7
S/1TO3I3C4Z4E/dCNOA7ikJDFAt6cLi2gpFG49+7ZqVrLPoqNxTox8oqyxSf2l1i
e7rgXmC+exlv1YKE53ypaULk/QhxVGnq6rRO9swFkww7ybnvM6Y+ENNHUCgULIGn
/u5YCk622UaDvC3L066jkoPfLabQca9yVtnEWz1ATxxhQILsNWmPqvNGaar8vCD9
72+aqvBJWpKonl9RpMYs5z4aduIn6ClenzoIO7qyU0iKuas0Fa8Ax9CNplVl3E6o
5XoVEw/8/CEX/5p2r6krOkF60NRWBChkPjgFn+Hr0cOEPaznTFdVQeMx47uhU1wG
lWINCZb8Ra73n/mgMK5erPUAySq/30LEDp0bEktb2xmEckXIu9UnSU2vULBqZcwQ
fhQmrpC/KW6rSlsr0mvreYL4AzHEqQampJ0fjItYYZH1aW4b0pdq9UtBNH+zIfso
TXjoPZSIWNKVySgXnVm4qLGmmx6YmtaC21RN8G7gbj5wQ2ag7m3dT2WhY2NZVigx
XaAs86ua3k55QecP1VYNYPKKJXLf8Efc6Dl4zFzOcnxZgKIRGV1GfUF41W4q3K64
qlRsCYfcZXIjQMtSDUCxPjsaFilvJ2YzDX4Dxo+9V/M24JTxzc5nSuL2MDSkkHzU
9INXGFcvuGMTnSOketPUQ31Wt6+HGNdaZpB3Fnrk7qaeanwlYo5juMOkkhFNvI1H
DOCG0EWcV4amaUTCbTirtor93fQlXASTFqoY6Vi1RQu9NcW0aZV1uIelElmDP6Iz
P9I7B0+BwGRYyydHqha37jp/pgz7PUNFAWF2vxQAOEoxluREB+SAWFweBVs6KL0n
VzDlizndbYMwAcgTfGJFKm4UeNrfQejOgXL8r62pPo2QgxGpXMUwb7FiCR0CEhA0
tfhAh7FU6y0CoP51/TQXfItUR0eAcnejY8bp0Htd/VZfGNwJAOn6nXM3YuWR0+sF
7s055cM68fmdv/pnrEL8/WVW9yxluuA9Fa74/6Fb0XsGylVnsqLau6KfzqerfpxW
ycTlKr0BfEhBoT3V/oBSzDzmvsSFZOUavD2b4GvXxDY8D8e8vbuTYHKjJcEgYW3j
75+njiPgTMzon5Pw3gQkL+AvgokGYJ95C1ckjOZqg051HELrqrn+LHa0/RY+J92a
2YyRbzUFy/Z9AsDJMF3YmqprkWxpQEMEWcBRJLp/XzckMs5E/k2JXwnw0Aym31ee
TqlptTGLJGuOxMZuzu8sszat/lpP633XFWDrYLac2lfg0wG69/3MrC90d8Le9HEU
kXEEptPlr714Vkctg4fsOqH5GWFaKDS2jEUOaHk6m/xoD5X9xDmP8RhiVcIN781i
3bDf/9LGSIfGgsgRybMLfjBi+xXzJAzN8RoKHyuoL98NpU8vtg+Q+nHYYSNaZVaZ
S3IA83nwoL/kapRtvEKR8lGmfeH2nZ+3zApv4PYf2smGFKLXifVX2Tz3ZDGUpfj+
fyAueZIyphFQLJNB0MaM4ZWsZR1LN4Z2mXFvjuL4ZXVODg8Ppm5IG1NF8K4GFZ5f
srOvOwzvXtOjGnO5C9f9+vT9W+YeyxLv9DYe2sOfnJFsKWogoOwFJm+CGFz1GsSO
JO7vnB3+0uJpU3vGtCAOuVMDU+NEYxpYZsYSGUL9H0hfuiD0tamBmHXlJgE9URbX
YV7PWsfrqkReYN1TVHAgfHhahn61ochMhCev1m+Yi/EVskuZthVqtEWEYA3HqDgz
UHw16U7KNJZ1f2pOW6Xs5ib6WEX6wF48NJJ7h1ZgVzCtbYwPA512SWSzuecrm+B6
3mzFzroBnqN+7jXW/dc7mPW3A2cDJ3A7CloM6FQRwjanVWKQkbNPSccNGAmyyAvO
FGHux/yyQiZZkPWBwruno18JwxEO4khSDIdnG9HwUaCjHQ/+xtxYRCrKb76G5HMN
gxKaeOEVFZIHEqcZzjysxj5mxIouYBSCv0Gl1gU8frTm8aPMrQWveUHyJXEUkqb5
qgi0bQc7SLRlFCAP63+L00rp/V7S7fKmUB19Y0JtR4VzjKL4bIVuSG+1VG8pT/i1
lxZwovcbb7tNk7jatJXvPR4wL/3d463y6EUYtR8eAKisqaqvCkzW1PKOS/q6BLae
3OzHqmStS+t34o+WJE/fgv2MDt5f0nVyID8h6LEJiCVvHkGi8+yY208OTs4YLwy0
HP1cgh5y1CSm0+4WElHA0Deu5w2pEj8oo/bq4AGDp+pWIjT8Yg8eyxp2Ahesdeqn
cVaJmNENSwyDe4HYCY01pKDZ/xhPfHU3F4kfVRfk4IcRTVOXXZ4lIIQQkybNBoyN
snrhYpwP3sFYzI2PzeQfslqPghFWCdaNN7KZ5rd3FbQ=
`protect END_PROTECTED