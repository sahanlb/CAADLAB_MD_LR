-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
asg3SVC2UinXOAwEs13fthxfKbBRAvnCdl4H/9fWJpR0ZWLvSCgGPyuJPsgr9L8N
GYkOpgNSfYQY04LXmN8dIHDguU0x7b8vxJYfdlD2TaXpFQdvoiUtrjfnAdQWDgzW
OWQG29CqGRMghEtXiCZ7UuzS2ISjvk+bgAejduCkllI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5984)
`protect data_block
X3+6zXx8xXSmy2+glT8AT6VOR8OeQvC+xlD1mjYDww4AkeTqEi2BY1iJl7BLrJ2T
P7FvdXSuMlvwDZRTXC8U5m7A2QgpWETLhxideaYmGJ5sfTLuYBOt1X533yv48GPw
3FE3xcCC5XZKHbql31m4YBRyucmCHacr6FHISaj+OsCCoQDs8U1CESJ36EeUT3kp
s8ocjEmjwlQd2nb5rKsMA0lWxd35+JBJ0Kt63jXR7nB458LQgBXN88BqLEXV+/Tr
1h4pBTGWatgUdm4jBY9iUqQubc95T2IfCp98V0ArukEGsxYCr7RTvRgwwBB0Bxn9
wgBFHcGqTvD6HqqUDB5olaCyGybdPsz5b8VYrbKDb2580696/PCXunsT6UJGiL54
Zk6q4FWXulEpwCL+U9WxKjPIcovVIJ2x7X8BwYgKkEeYwEuNvJFs3MxFz/CNW3yz
DMqRZVXG0b+08TNC7RBtW0+ZbbqpfPUvz/TsiT62XJkiLxKM3W2SI6ZnCpd8cJLh
Go15gF1R0JlfV1F1xcK61OVZ8ymhD9DusnXhctdqEODOhzUsAZg4MioRxB32LGcz
arHJ5bq+cOY+GhOGHBP4ogMJIifvsDjksOmDGt413+hGQrxn6xBT8anAPbNBLun2
D0YB60djKfEwKiAQmqSspAc4OpkwzqMzWnvmJgV01TjrLxBlLp871kAhvaPb5qJP
bxsULxcB4WY09p07RCdw9QEMTDq59Qt1yyho6nR+nDHv7L0cqcoPPmkjBF1LfH7S
OqNg38l4UpV5kPcVZYSic/oX5vfI+SeojTHdIU6WjSZZTz49SlYsgIT7EWZc6zKC
OBFHBG4kqDpiQalhmQ1xbF7sK+V18u8T06KQJgvk6K7+ngF2dHI1GQXEZifxgaYf
ppRGwgCtsDSK1AYqF3hEmc3LBHYpoeWORCgpAxJxYSXlKgny1Ng5GJw0UwwpNuTg
YfUC0yFdhTBmIsIFoKGHCROr79TBXMzjtVFUGUIc2lS+q6npiGxbtiIkb/FNSSyW
suwa5xcCAObQexPxBuOAAHOIW50Wcy3oJFcSEfQZa3gPYBolDUtZl9TGmeKmI/Ya
vZfSuQIt5YshNnWdwWLWuWlSLwbBcaY98OW/3nHD9v9KIlNI1h6BZtQRGJpn+U8E
0A/Rcnuqzu6ugPZXAaegga+/R4WkKimsRVdOlYOenmcAZZEKbl8nNCAVfaZnfRP9
pdR9h1GOKHWwl3fCmPbadJd/G16acwUR0xgpci+/MxdnAsfCFl3hbS2Cspd62lrx
M+cJ7afACnWJPiFnz6wp/peFA2JJFWvtGOWWLZc7x+fs/njHY5Y/OsaiunXZZHYp
1WCnU0/8pAyV4ZAv9wh8TtA31OD6F0EKEwcLZ5bwy/GYu46ZE+QHu25fYateBfiV
BEFniJoVFNv9E57FpLVwBP4SFm4CrBqS/8f2fmOnk1fbBRTYNJccL27906tg4/qi
G3dZU9kLnpH6WmrIwKECNyfqB1M4cZ2aMeNrCh7jx/2uy56POWtBktQ8+GMDbn/I
805i/yj3xExaWnfT7aV4vyBJsfP+iG4ScDwVqOL99V0sQRxQ8ewm4lo5ey08DNJg
m72MuIuJFTxxa0Q3GgLdC8ERpKztV9eSjjtfg36VO2UW042w9R4eFhALVZ3WmXTD
Zgielq7T+a166v+whNSRHXUVEhkWDSDV8l9ApzcpwRdkeL6YrvSu2nXXKxYogbM5
RLvR3ubG2dXK1JMmXncTVm4KGHhPsUdrQwL/oSDAW53PTtBGULRUW8607gjVWtdF
q5WRAvWRx9i9nM8zumaOPAlngwkZtjUqp+YeSgHvH/SCOk6RJUuBJyz1ZdhfgLtJ
3CmLzi80zBEBVD0YvfbGjT7rQ45JYmhzXD5Qo1+8arKhfI33/Nt6zxs/RPSOXL2p
s5YFviErdjxkSk2/i4FtnW347bLTPgySEAh36jLHhgIoeZccrDYRqBBaa16J6BvZ
kIIAjYKTsob6mJWa7BIfxmcd/CY4Kall07niphXzo4CrFS+ubF4DJeoT8fCk7QBP
g3YHNr1CiLGDF6KL6uoU2p2fBph0/m9hVc5FrKsPjvlp6H8okxi7uXwVH3Q7wB20
4/H/qzKwegDqnjHL038qO2INEP2BulxJn51y+gj1Th9CqP+6E8UBWxG6b35JuFZh
+qXH5ArN97qn2kzSk9lkWUp5XIoGIRtM0XxWZR/BCSlTSydj8E3B5bYVEut8nMhi
Z/agmuI87oFFyeUZwlo3grZSUz4DKsbTxmRuvEhEMeY72EXDBTphmCliZkszoZ0T
rwL0mWqTHVLUuG6e6PvuMw95XL5t9VH5wfQQ6fpxiILvggIIdWwIJPjSawK2XdHJ
v3qDblkbl+kwaH08F2k70q7JuKrXy94yDuM6gGh4cnfWNPhzjIhy3KX20/mlSNMD
t7N3GccLxKbD3i7HHuGTZeDCWKDKGjlwBYKGuCVPWmGPQ83Hqon7L0m5rclIFDy7
At1z4y6vbPntzUgbg0ZXzJUz6ycswQKbWGBPlVnWrRCqnjIYLDoYG19eeik0awdI
qmxgm8+bLu4GDZEKM+ECGE0GlVJaONbljGtXWH2QyT7dza8RZ7f8HFFGu4hIRw4o
IInvnUsRMUbrwvCWiTx9GaRHrduxOJ1NinUvKEVcDG3thQuhfLltpDjSfvGq05pH
qngXT+auA5jnYiTGh79I1Fc1O2Y/sxGCOhjof+VCKG5KgQNNrmpVgCCujqoU3YSR
0PemVGfmCJqkkeFY4SJPCo9Tzze3PrAcuEtQyupUYiOe55neQR+e9Zl1ZjOnVotq
tN6PtiyW2zVWv0teBAO9njfqcEyrtWenJykA7lf8hhCccM2b8ViRQyrWEmczotlq
8ZQZRys0nTGjHVyr1/azQR5Y9+BDI7PNtwosnMSC2Iqamwwh6CY6VNk6++FH2zEs
/xZJi9wb/Hjjz9j5Qmyw5bG8qEMI+FEl6xvCf12bSJudy0XB1UqWwx8ElK5a1Nn0
oGtK2CyTc0wM/BCU5lxEAG6KfmxBSEycE52ZpPp/iETJv4AECjcb1z4AmCABxOki
Q2nYvOy2XMjiElevGonHyvOrVApJldORvRVhU6qs8T20grnG0AuKjydlgy4/AxBw
Djb3c5ffkzPC6sxo1L2UOs+5f+4jBB1VT8b3ex9/+hy2EhIm7HpEa8+6hz9azJwh
Yo2e6x2vJtzzlqyslExJXVFCK/5HU1Un7tEK7NlE7BiWoZVP/mFacp+mSp1X/pIG
ZdjeDfMHxxEUtTYpLlwh+pnwPAMwyeHRcb0uzXjpgmsiJt7CmdwxjDrCr66I6itR
pREjwE9hhyKqdB6LTxFhbjdlQsG19XDBCK7lKHVxzoV1bOekkzQoWFtOAEK17A2B
VYYngLuiwvYS5yywMYVrLpUi7prVh1YiMFp3Kn81nzo1gu1UfxZBSovjhCFK9q/U
7g7F5cgTNNF+TT1N/Llh/cuttgs4+GF8mWhmkuDRBLrlOGzmNvxu3gaOBquEZhWq
Xtt8kqFkuAvNKGYGRV30AfcrtHp7utntDAmuR899zLf8agttOnl5mFYHlK/IWelu
2gRJ8lxRF3w8STPMMVcFEXJSzW5z4XeGvY98dApWdGU8C4EdaBl86VR1hwDzGfF5
fFF6GruC4J05PB1s/Gi90+Pbhib2LpbM24S/xyySkHqnVhT0lqrm70Mnuvj6e+u+
oCaUjz/rOiZqEUivSSmjijiHdLalH9b64Ucexe/FUGCfibokTl+wkipSJMkop/3r
aC3txd2m+hrRwGU31efx2I+xNQ0KyDX1JGWJqGvkSDA/aDwzg8Qzqw80Lq8XioYG
NuGMtP7TwEyCpXwHqvNK/mjLZZJTg1qfaE7gSV1bpcJaf5Vqj/8cxKLergxFSKIc
EwQ6qdMJxI8Pq+q4m1SLprC3XKNVNUCGvoYIH5qzyd6uqlAl0GC7Yk+ry6Vvc8gu
YIJhH19UL0xvpsyzoh0ZY6omjwh8zrfNzaRgUxUpPRJW/6NpcROZYjeVH3WGvI5Q
NfvfnBObboWCy6WLkjK54NhCXx269oqsoCepCugBQ3jD8sp4MInmj2oCIP8p8OLb
cwJlTRzR1XdTesV3tz5pbk9tbz4W57H6TJAbToufZWiUOcTU0EYWIBjzOkqOU3Nf
9YxW9FOCUghA2xrnI+3DS+9aTwYHBg4ZrhgkY3vaWSRpNFiJrPLlcz3+d2e/D0CF
vy+widWcWywV3ojDd7EHUbQZ8Ik/90u9xL6A/zUMErST8FvExYKuN5z+nIrvQ/2g
YqKzm3R54BbSnyw0X8SwZbxWwUl/DQy/AQLJd9Vmr6ayhm0x+77urfw4EnKZVJls
Rdm8HcdpdovdUxj/NJqUQyrkeMPUAtfeYmhLQwY4yPFksRgmGnME5kOkuNZtY+eF
KwhwqEAFuecTQKpN1MbWVfUJcLGwjkpyaG/df5n1rqT1P9uDAP71FXnnZm0ZB1Zh
40zs7h6MpsDXsUEPXkHmN8gyMTo5QzFjEspKRos6179JfTJT5CeFrNlv1hAVvDNW
VSQBPpulA8G5Rio3fildW4kpW91kBbQh9qzwh0/pQ8wGUGnrsLMO/9LCtUZEX6FQ
ufF0JtZ1aDhT+D9yzDEmLYq9fqxzfio8Bo2fMREmoILPzFfvoe0NS0TFeOP9o0f1
Ge8/tfwdgnT3KlPMbnk9XCtlUwnteRvFtzmYNgJLpW93smtwvKorEMFw0kPkOtT6
TA+O+Nl2JpiqScC8/DNNSB2gNfqkkiYzTcJGclGPftoh3OGdia0ZSDaUJ91X2732
r27vu/dRut/yUhFnw9q5cv4ODhs7aiB2ucYZbvGw6MCzK037MhqEV6+VwPPfpH7L
AmHybOGPg6Yg1Gwy775rsFfvwls7HfT3y0ehQHjtNC4Itol3JdZr+3gh1QvDw09d
5N/tisDqvMvxwmJe4zlb2kcHf7V7mbrcbwFE3jw1mCOvelub5RtA40//BmCATUSl
WSZ9N8+tbYNh9vo9xEbnpzktT0d7HKlJn0YFU+XztyHtxqCXusyaSFDxHY3qccRo
nxrfRoCR3mJbzTyzK9kpjtZkXQv9CG24c/pQlZrgRolZECMAsWRrih9XTy39ydy8
GF7N8LR4DsYExuqQ0GxNUud5EmaZfzDGlAs2N19Paw3j8OmB+w0AFvPkVcLnlPvQ
OnMpT42Rk59mQUwC2xVg046DYE5Sex/FN+9aasakkMD+BWp1L+Gir6wMuZlt3r3g
BqOl3HRFLdQ+6S2gNUwdkKFL2fP2Si2CHi4N8VE57ExCi1QUy+BQw+iKpDeCwgYG
RjbrdvdmlJCvDikBAjqFk32wMHatyQaz0ycU2ACVa1nbZUF3nqNh5fJ0wuB5ZTV8
cNivKJXetf7MN2T0OGM3bOOdqetplpC2vITSXjG6jKZJbKGD+FXiujEn9T1GAUSv
9pFowrOcgWOCAC2F4XaEoWXYLWV4pVC4jR1nTLjpize7JixMjn/QuH9VKI1L5cSP
H+wIG/bZ1Coah1hxAoVSQ9dG0PnDRZj1rnxtovcGLfxYrdIh6ok4FMpgL38+3RI4
o2+z1arPChxO5VHNAMy6dCLWfwgu3wVEN+BjgNzhhyliNFelDTrFSzSu8O3xc4w3
QFnotmyQ7/1XJEKn3CDuY6eySAo4zc7O9m+xJSutNSM8kdUxO+CIMICNFrCy0M1+
xY82xMNaKvGH2uKJtV/Mrj0S2bBF5rwjcHR2GRiuwBfy3+3cQI3Y7BtF5zMtt+AG
dd7CPOaGGOZ2a57o/08qf1AtJzvw7nae6RjHt1CjKn2wJvQndz3JxHZ4krHuJLmU
EiP0rbFbgEcwawwjCh6fZ6D41tyh20lH0H0IoLM3ZHvYk2AcC0xe+WtJXb/7qlAd
6qi1IMWFMxJBmwMGbFeyfqikepMLc4p/IH2FlvRHDCJETsHGe/eyu3sVQrvsE8s7
7V/uNdAcFFpBuF5+sEctYKlZ/1YWqbwEFazxAtTQYZxoo2HYBWUfxqJRk3dEcaH2
h/B0Ly6FZEm6O2hSxJ7AoiYyx2kSdy46p3ShaLYqrWdXjT8ohcpz3Jp43Y4/wmi/
WEuWat5b/4zclLv3hP7JzunF3/RVU7GtT+55H4alxONhaEjxytTX8wYWnPV8tL68
w/81MhX79swaI9XxYcJW4WZcjSmXgaMKJQbcsgCc9nnauL0k23w0acYvHxASzkzi
LIPO20US6NG9MHMlThqtY7+lMThvYoSlTUwLqlB2qtFRmElx0oa7u/Tqu877dPsW
4MpRefcjkacNCib7M7TTo7ZBboUM8Hx6QGckfjfoTuUAujBv7JANRFFRPjPhetEt
b7pYOYyqVUSq4piei73cn6308Do399xJASf/7c/gsX6BlAvMxiBvqeNz7LaL9VtS
H0zL0iPgt4/olBXRGWA/6JcI5YcmhXEU6OAvXzVLqw6/mzb8mV2h4x7DcljmvTx3
AOcQ9soxlVXSzy5xRVTgo1SkFp3uFpnP+7CH6THVj4/2/7p6+s44M4KK9WPlVgyH
Xr7SzMRSzZ/dGqGMG4dkguVXdYpn3gZo3pYpHl27rDZOqt6DnBdRapirQvs1CBWq
19+TvyPaCIvzZxv5cVpeMdnJL+pWQowA5sMfrVwg0P/KEzc1TB4vtCHY1dU9aO8s
WKNaHGLP3m5q8o54ywsVcAR8unQL/+OuIE46liZiHP0Qc+BRA+1xFdGQsc0g3put
RMCRNPFuQM0KsSLIV94tjs5E7sxg6KSzH0cuL1OowVgbkr16PlD//2rCzhIL3HTS
kDg58zc8gSMaRr6PGgPu9VtloKXwa8tjZq5YMXmofuPOQDT46lTyalh8bvjYIwET
K2hfsnE7o1QJBLEhUZOEDhT+dHkNhnTQyQimnGFt9JPTcXfZGLhBMgpTL+xV0CXI
nk5htRrFH4Gn701bD5LxYynpOQ99U0GtqWW356RWMkqhQuHFtX8ljJa4VM7RQhFc
l0jjQsm5WCu7qCBSnPyLSHtw5++RLdi8glQ84xMAARWNvvDWNKDHI3B6jYa3Q5JQ
tkeQ1xtwYCoOdO1ovlKRuqncJwanUqryF1bjbjZOtB2TnWM2lS/b3sAaMxfpvckU
iX1Dj8agNIMtOMO5cfzU8PswGPD8ucMtMUHfXk+g9Kg1VMly8XZR3XuymdgSu46A
TuwaQoJTjhvc/DGP9vmc0IPziUxqYDnk3KP1w8YAi41lMO5csE4sJSqHbVmcCHLU
i9bWAfkhWnOFDKMznCSLOrzdFqAm6YtkFB4kEPXmWkheGa6QW5nDiJVm01lJwPrC
yLUzTjSJNBW4umAOrRtdS8lJAAGmuFj9T/F7Kb8Y5qgazPtUk/TAr0k3B0T28/JE
RkEoPHqChHqjxXGSkHjldWE6Fik6q61kTdNrqTAHAyWryC6gJyj6dGcK7ixM2zsa
y2Nv7aCUO1lniybsYYI1C8R+WT61X7ZuUGscdjUcMlQxVvpVwZz7mjHaTcd1gRUY
Ifep8XvZlLnzAqzcPwFyFXyNaOmJeIGsURPGRpYTxTbvh5M8SQt/xiVrnD0y8tuY
fG4PYI7SDHLYAfe1vDS+kkmQLi/X57UeCwcvYKPpwN9f/n+0WJkLa3zBuhdKFr4O
dJW8s8KV0P3zl4C/vHUvQXNzfRCr6b0Ti8SOgkaAXi4P07WyP6CaL51m4CcMC1lN
wNljD0/ppWENVAx1TDTuDbh7d9nAyHBZaI3cjHcY3Yd4iVMgo9vK6XWGr8r46KTU
zofCJpCFLlNcyYO5my4vg7uwC5oz5U/aQ8NIkd15udRIK1Cq9eYgy+G+9OPC7h4x
sIUWACFJgs083WZhbnew4CfMeNdLiX9AkGU8PK/qDH1glYaHY/TWJS3tXoyLfcfs
gld6e8w1KnXvxaXt9nq3OxZFVzBEvZ/DWqBBVqgBEEYNGe44ss8r91zJa7uHRRxa
AA6tl3PUhViZVBCU4ZaLmeo3UpJUJV+/z3QMHpglunI=
`protect end_protected
