-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FnKGW0/pbvCyO8sKMHfreL6Gbs0xpwwrYwoZSSxpKHATSwahur2a+Bb8i3oTCxv+Y+zGrNrqQIXS
yFhAtJepYU493a9YHnbVUSZNCc4971B6o176mjJHMXXS5HGLHQOCAQCyqtnb5fAqdZ4uFmzlaw75
zUMRdnnUd8PDHskDR3DbpX3NAIzPZjTmUfXF1eIB+qnbqR8NnkzigkozMDW/uJayZBsI1LKQEoob
N3QdEERLn/63V63IQtJ+zfwaAtKUhRbVDxZnSol2/nXix4eNpkcbAqV6jlzrAPtcYC/NUyi6ZvqD
0G7aqRhpGQ8HP7fCsneqYOce3UZj5uhZAC6eJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1040)
`protect data_block
zVtaJwtcbuP7EjZtFrRNNlgJdlDQbBZtaBBw4DGe2HKnlKjeNf4kKltkUJx19HoAXqRg5yWrwr2Y
5bqx5YMwp1NddBPczwQ8jTgefqAi+UBzAoID04EaedC5YIT5XH0VXzTs7tuasauXy2e57V+lzD3V
dm3kwTQO8AmKohp3GOThM6/tXphpowrlzjOElqOL0+gkO7I90mXUp54C+15yOoWk670CpzcnqBaD
Ji8rkaCE6sHXzK3IbLqMPLTbcs9RqMnbaJTyjtC6wR2CgarcjRVIY2W54IG4nE3YXBiyap2w/SAD
GlCM8konMShGEenPqOhAZu8OAFCv+NKpzYupMTGUp0qXOyWQinY7CAiYmzE8N6QYDGgJM3B5Rc5T
xyPWRYA8TfriGiOEoA10jOR6ju27xxn4T6yoV/9a7mMyYUgztMGt7mjhZ9PVOZM5vkXuegXvfb05
GBx+K3HwLCadmjjfknM4CnaAbCoPES+11mxk/SirzD5j7xtmd5usqx+pWA4P7O/OcE9wX4aWG4ry
g88xZz3L1QBkqyjKG2FNLzsPLBICDnH4zjJ0/HkXxCnSlohAh8G7epIToG/8pTLheUYtmMK/yBXH
OGnXI/QiEXAXdAv3vZRqggqrvQDb0CFxeG3/VnQxMF9+jl3WFuKhjA41YmZD0mOA7GXFEp4qo4b1
gOa0gsTBlWfOTW7vrKLtZQH3FYqfBP/b7Z7oICr7g5Mu/apLWsGiy8QRQnIHlBhOnEQ2dDOGXsge
8blZgmc+1yKtMroR2Rw5rAFy/B03Oj1qK7CVA/86dHQDZQS3Ni4N8W05oZgkP46q6IH5CwQtQsM1
fef90JpO8WgAgZIGOPap+Qlku1i/Iiikhfqsb+a6WZQwPC18tmKHz6cnNmH+pG5C3i77ti3GZaZ9
0fDJo6w2Cy8pcDZPSlPXt/DyoNeFHRJfTVbv16AkFgypp9fOiZQlEwj688B3l7+aIVfwjAKrNXOt
6hH3fUZTtCmYHASMM3qVNw22u+bcwwTWZrpGlgKK8C2JL7Z3lzca4GBZI7SMmNnVYhfpLUTx4c/t
qtTC5BpXODPiCte06XSRgo2or09Jp76HQjvqykU265cwNxKVujHfpbuOS/tR/LonxMZjVHQ4UUHq
NKZaNNDf2MHugOy7OPYWOLVGv+IMG4gRxBGmBLP9Zz48a0whqD00vW6/DGuEBew5Rt4t9GPbwh4Q
S+kY3dme7biTTzOH7aYPZw+BQJJxsPSycmNPR9a0gxN40S9GEh70sMUb9zsv3+4X8nzrrRe9CMXB
rWQYe9LfQpU6KpfoN3922iqm5dPBludeb8ti4VlMOT7+1TrLpjnYaoXPaOMKt2NwA3t+AGi0Zv3t
mI6sUtkFSa8uJ3wHCVs=
`protect end_protected
