-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
UH+q6NBiT1avIhlBOwitKZFyQIqgr3E9bcYLDcrv/LanrGmD4XE25sBkzDCd1kmA
6JgbvbIP8uP2k+9Chj1+AqhKdJdDpcuncPxALmOIx2t/JR43c/0fw9AfGaESmj03
yN0SRIEytNt4gengQFaPwSDnWCD3wCslPTMOVvWUBOhFkoH1KNSrug==
--pragma protect end_key_block
--pragma protect digest_block
xn+xURQuj2bE6JN2+Q9nOnn8SzQ=
--pragma protect end_digest_block
--pragma protect data_block
uZJ+rFO9LiVr1FefRrnEov+2aZDfKbT3ZWdmPOqSmrpyT+IxCeVS2S7FHEkGUZtf
IvBbdE+h6xo/uA3U1fqEovvONF6Gtpug4ZZp980t5HxpXg+pAh8bEzc8IdmFmKVR
FNvVYf7WMeInt0ELnkG2YXHb1PCruHAKNJ6tZfPjWn/pj7uA0yBtrM7TvVzg4hKW
vlIoUdOQGlmgzA4epcK/4rwJ8S2NPivqYytwQmcQB5ZGM6saFTS8u0h7BSmVMAz3
nxtnuBGfqDWzMm2i8mGKlWiikaNzUw/ohRAmNNCmSf5cVPyZkmMC7CYUfjY7ilLH
abVDapa/AuOvWQPkUcrBQvT6Evo9ERVTJoJUwOVokweVMkoMR+Yl52nMtFGoCCQq
k9WsEBvkcn0MoEQkv2WDQlyUAQ/OMG+RL/k0Zfn4RTj39Tx/pqOzFObUWy2lbfTb
0xSz1APQrP5cMxa+uYf2j+tkso4zfPyRLTbrDKXsMW+2TcF7ldQYoD8fM10haMOP
/IKVw0Qw3Tctus+JcnUzV83B/0xyqLHpwWF+X0rLMQY0vAjM6gqG3bXWfJWBOg62
aaToS8xeliRngJ2nclg61HPAjb+KZoenz13FXsx9CGpQTFEjx9bLuBkma6+ZHCDP
5OMGEXq0U1Z5rnkibeSBa9YfOQoy+rJn/UP8tg28rkJJsC3kW02Wi3QcFfc1qYib
oMrWmInVN0XutD/TWaH+LuKmVZ8KCoxByBfHmRBGurSr/Eds5W1/zc0p/iYMDgtu
KJH6f2ZjcozwYwztSG7K4PqIGeIYBlEIr/9EejTXs/oYOf4lx0nbx9g38ojL9wyu
+yYSa7w/NMpbxVjTkiW0hUkW+PXJh7xmGVlkpTjEK4Njk0Qg9MkKZ24lucKOOkrM
WrQ0UwRBH58sn+KVNuCPnwlEjGO8OebG74UwvGnpPHolwOV9ibHsrdf0h331WyMO
ViO6jme+WqNtwS82WsCgVSilgUVNSSanl0m39fBCOfMvu8cYmEZhyVnzr+Id/I98
YOVRNjwuT7knB1qZneNwchfgZS+2Xt9t9Sl5eBpvAhUx55z1iPo0mXACKq1R7j7w
6qW4yMh/88gqR9dFXyHvvc4ly08RY+uO4ZXxzgzZJI528mH3RpyZqcN4jRMXAHAt
Q8QoqHGAMgFVBP+mXbpIBFs6gx60f0FcL4jThLT4y/8u015HZhr3biPLEaj8gdMx
Or5KsZCu6ReY53Ovxyg9UBc8xKYFYQ6O2gFg+nGcMlwadCASVSoIuRXATL7cjVmQ
sYGSQkofGcO+nxMkZm+rDq7aPsX2zbr6Z0E1iWxqFgfs3JKcy6XC0NpwS5V30+Iv
qpeXSFGj8yOe4nRI9cMnfv8yLYX8Kz6J04ScE5GZ4H3X/XCEhg6CjgDiftgvdh9/
F0npSgz8NVlylgVx2djRNN51BhoSDM0HHFlSBqNYqY/EjReRmIWzpRVOdEggT6cq
90HHTctcHU0ltETHGtoRMjbPQYPM0Bz7RkAOiT+1gn56EuwnU/ELsV8veQs0bXk9
gGpQu2Azr6+Z5InGOIgPLQomx0L97I3g8PGHI9gRV86s3rVZG9rtmyzDo0LcPSP4
l1DE/h6yZbR9ipeZYx8MllGXWkOdi776SAHk3KaerBB79+an4QxvnH1Qg0LYiZ8f
njunZgUSEMC+Ckl3zl6tRG8m7p8J+4hS0jNHO47LHGkDRRuV20N4EmiEEAgnuugu
MesKyKMYp20PUR+5BtZOmE2bR2MsgX7bCekYC8Za9D9Meq32IHo2u0ukm47G3627
9KyvbcgezQwxc6wwyaxaK5O5zkKQ/bTuo4b64+1z9et2Pgt9iq3WDNohhl+IZ2lm
1BjhOH0xdEOZKG0djGnI118GEwsJouWRu4WEtm+jIBx78IK9jlbhxUNTvSA9C2a8
QeiNdqi9I0wy/o1nuZZ4UDqBEsCvHycxaNKEihBBsszzrIho9dVuxWOyGiuRRcIA
ZuL/LG+C2cybAGJxv7R3t/92154ce18gtN8JQgNte77qJ2XKJpiSNAja4oBKmrSp
J7Zd6DUVUAr8v2P479z0T7NxqOn5k8EJywq60nWkrYoqBw0YUd9/QTwjqSXr/Qvj
8wo1fp9iW6KUnTSgDrl9ws5NTor8bRejW+mlbBokUtgU6L6M5tY8NGLZ1VYqWhlS
VziWXtuefmknotRDxrcK8rM2KXnaySp99J+KQ/Tp4CPaSl2viT9ALbQeVP0FvhIL
3zddW0mc8LdWCmESZulFirA/cKsAO0xYUcs+ISY8jP6V9IrC2BZue35Xihes+Tyu
XrI3nXDpwiqTJPpkQwlN51GfVJsnrMtasGQkE1W4lfh3EdK6lNi0vlq4x6SDV+G8
Z3gjMI2QVV3G9eQnnLWO5AHM+RfsEykvJhlpU+mB4t5pNPMoMoxk/PHBu9egPt8h
FuIB9NyRyxi5a58L+POIONinaB5pj+kAZ1FT2d9weSxpkQH/rMeWMnqqMGLbweOg
Am+SFYxxhacrlYTvO7cRW5sBFbwMWVv+Pbk8a6JXODCctp0PXtZlITHvbcx1gS2u
1cKlaTLyAUXQ5Y0/9rrCRJE3OmdqvsaFbaTA8V2+rk56/xHNtfChrUhusQV0MgXC
PEJnwSpF7KcYO4PMw4s3sJgccYp3xKGYdilb8hN1RF1zoQaASgyTjkuvrYaze3n4
8/SqpUHQXRpGUzo65OEBBO3Hm2ZeoTv8uPi3lTN4R10ATmnSM5Fpf98JK4rrYikC
kxfEJjlOoIuQY+R3mFP/Gz/tUrLrHObdkGq+SxSWOO/9maCYdA7b71zIjga/mQlZ
FL48cI48oLo2tCI9HjOngOrzTpEmVAy9+bxLAVd8FuMKyxAwpk0H50/BKHPV8I7i
hmW29gTPNjuLDueQKKo4WztY45yr29dddI65VCFohIIMQyRqaBhJFAZBa3BHWYIw
IV6FoEPsbJrCEFUn06pSA8G8UE03QwSFQh0y5o/BGJ/SVs9gVy7vOlzf4Rjq0ky6
fNWnqtYlNsjwJBxmT0l1xdi0Bp6oFP28Khsh2G4iHjXCU0rzRHSo6oxtOs1avM41
rAL4fQxD1n555TsZ402Dl9NhAUVVh/UsL8hDtXnTG8z7O3y1F8MPB/gq4uH0os5A
Ca09K9C6mwjH8s84gpJiGE/704H+YPqn0k6ySmD72ZwaEC72K4dH81gHT62fODcF
0cNipJtP6c/V61SXcWyAVGNSH8Moiw6SVAQC3accNs8Fd9hZz3PdyGrRTdOIYHnL
08um5lsL3tJS4dEZI1eXHal1wnN1BQKR6lb/Nfw6jHcXHWfaofrmIkChiKibkjfN
98Rff6ekJ4eXC5P9qEkLj8l5wJzRWa+nADr0nzJbIOrJR46UgVOJfWX17m7HpOYb
FONpW65XJcrCHmQkc6rlkkML0w217gq2xZc3wwT5NKeqjVy1o4jjPa5FmrbL8BBm
RbV7BDmLxXnzbZuq7vMoIQ85q8RQK7W3/6FZ6MYswWjymFYYbc3Pcwv7227FqT/5
y529DpS8CuMPv4XwTHwhbcljXWSVXnZ5v1vNQkRRwugInwvLQsL2vIIRXnAjQ6SX
xJLLAxLm+PR+bvuThIK/QythPpV+A+2VG+D2RwY2Max1XaxPUhCUQo7BSXqIx5G0
NIiSHePSlhC4tquumoTCc3BLkQjaOVku+GEsMGr7H0GN4E5p+/y6GKFR/YRHEzdK
yAskW0Slk04qJs6BJF9H+U7Cqcq2Lf+pCQOWrlRhA6puir8vJ+KHhdbqPIjrOmCf
Q8hGRphdddXOB0uDSDOpygS4/vCIwNStOSR/h0GQ7lyBoHvZeA9KLE1ksmau6EjQ
FykeAAYyJ1pqq3OPZ1lSgnFcg00P/YOAlt+wuSsMrnscVdeBPIONi3fPSprIrVEZ
qxkFJFuwmg+gnufynD2KvY2Vfrczm+B3j7BfCvS/MNyZdmOVcT4plwZvgEx03O2j
J9+bwiD8i8LtixUDc+uU5JU+EvXUUnSCT7HEIgXyPAilR6hcEbRt+CrsnZ8nJWNE
0Udc/HxdpsoqBHf1OmAdfOUomY1dHXEdbYzbzhz3ocpApDSXokKlMdLQyRUyvqtw
aDs5hbEnVE++jxg6Ny/omXyrQWXjLINi7kQy1bet2p2sfQ0/MjwRAUGJvBiXt4mC
QijrlKmlD2sWqRCEZc1XvqgGw1gydndcrd213Q+iNfHv+pQtG6CGbEUImz6xAAFz
WeNrGwkvaH6UgKC0M+gML5DtGCLkGnnmALXfZuijuRBVrPuSu8pTMD5dvCqtCeqX
0a8VJxtlNgvZI2cNy4X9usdXXbGsjt/OgSLB9icoyYfLy2F1jpg/ZxoC/zEF7qJh
EypWx2fEUekzsrJoc6JsGXqyWYo1gg+SYDAjGkNdsePQuEt5AJwqaqdGzt1GmtmM
AmLYGtjHIVHb0HI16b/A43ruOEcRoNKjfO5lEFWTmDu5nlSpDxxZlfHpmzgB6Gek
nnCQief07BJ+evZvLQ6RiXfN36nQI1yUkESkdp5/26W0uyWyoaMv/BtDkm5lEAOm
GlGq1X0u0oCznCQUnJ+78poOC1elMXcbo35YlKogm1STWH2C2ubenlcPxOsmpUv4
tfuZUEvw6uICLU4lnw01/4Jjcm+DEJJtnFfFwm8GdNs7CxSMAB5snc+3V11OzVeC
ujRgFiXVsZhRfqzEJlmyunqlan6ko4k+OG+m3mc2vfvF7+EdTA110ynHUcjNW6pi
YiZmsDYPQygRYuAtRL52Fvl4pXGueOi3flptUpS5lBqAmlRGsnb9tMRzJ/y+RUME
pg4BBLPHKDg3QG+Me/dRN1hMNYgS075DaBuTIuUzExiNFoJ8F2JiDmqklJoXa2AW
n+DbGmUgs4oRD7Uyu2fKUHu/PU6Z9P61TXXf86dcdszZg8EK+hl5jprGNyAKXbXl
ZMAxHuDkfhuIlYulIO0ccrwpjnt/JopkpbNghJzxTe1b7pihp0tXxZAm/brO+vhN
4dWlchI3+IZFLN3RVQ9G1uRMalgZmGGFctXpe4CT0OGIv1DqASAr7EV3GpDNvyer
/J4xoUTgZHKeNHNYpIF6twO8FzXXvPs6D9q/aoSGAA06FzoUJ5Io0ezElyqsBgqb
4Lc0VhfRzTx+yb5ti2vK01+HA8g8jVOHakC/02rA2DQ5zxXBCXa6ncdg6dllqU1U
ovwyNju6pJEMifyHPIhN4rNgf2u4w9h/V/zaevqOhH9vHS9zCqBIUuh9uNOr20VJ
zcjPrPFu9Hw99iPfQxq2OTBx06hQk5pVRJPgkAoWqoV8KW6yZbimeXzbPT4pDT/R
G9C7DkVbxSJXnCkPx5oXabNx7IN5RPtTB6roAxRaz006UXfSJiXpSI9O0S1byD+2
vYBNt0Ls3/ZrpW+je3xIhO4gzhf8jk0iIIGizjuIuHFQQl8AOEELSWUpExw0ajto
1uVqPZbfGAPhABZsWhfIdY7PjamFO0sKBxplZdZFo43sbCWlnwUawq8BC4SKzoL6
7OhRYvW+d0aSIVluNqOWwzFdqRXYCkSY/xXpT77RdhBixwj/Ij3lvVY3ySMKuH3I
mdGNMH3l4GHiyD3nbek3mxFtgQo1fF7atsKK+0e2fE6QW3wDrv1nyGyPKLcf+i5T
0OaaO362CaJZrYA5taRgzOGfMIOWoYv9SmkVnUw2YDvlJsWiHMB/+67uu7B9Yzg/
CEkP8ISEDtzrMDVk87L92nZF3Np5TJodwDxOeeePVvqfnFvoLRbRIri786OYYp/7
adLI/QiZG0PJEiEB2A8OrxmRfSV6aK3h7genYYV/TcEQ3/ocG0tyDGy3ADuHUyqF
wKNqyujJCIxdjV0FA7oaKA==
--pragma protect end_data_block
--pragma protect digest_block
CNjU+MDpfuPH0wCwoD6ozxmEZqg=
--pragma protect end_digest_block
--pragma protect end_protected
