-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
WalNz59YZpNAv9njzWmaXyOT8Pa5+H/SBnWm1NGu6WSt/3PhVckMG+Mmwbm/LHX8
sQEJHUK3V7NtkO9US1NUw4dBHygdKywIc+FLVYRUvd/oEujOEcxWumP6aj1vVaIw
1vk/b2POe9wICsbKOAdL7WgVXRfTZwxTshZjAabf/vA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13209)

`protect DATA_BLOCK
6ZTDwkX1dViD5AHO9QJZBWrO9f3m7Ltcw61nIgggsuVtLCj6GHtHSkS/81Jucp/c
qXaxFFP23BL3zbvVXnqp/Q/ztxmDmgSlO0MFoZWSDkkUkupPoikjhM39BybBwwR7
jmzq95rOxY+rfoG35IRSrWhN0s7O0RwKhRgchr+tW6NucIH20A27VfRbnDNVJXbK
Qq9lNwaj+MrPPjpRNwu/g47GK2ZRt5TBJEf3POg3exKVqD4iRPbRpbnrT9a/WeXT
ldaZUvockYI9w+lkunLKnmdBsp1ggRsMbWhP1sG2WnMq6jX6NeH2IbAnDQivvDII
4/qRO0sD/a4PgeVWMFLSuWP5vm7+T/Fh3wQJGs+pzDri2Hxtm3Yqb4PJs9+LSz5j
UCn612D2Cm7bpQ+97dDjPqecIbhi9qKSDq+bqleqjXEZ376qHz9B0qvVG+PQjdQ0
YHc1R/zO6doC0jSA1archTrGWrSC2eW9jQ8plrlm9BKhZwdJt8nDM8CC+TjghXL6
Kyx4pU9QRDbsxTqOu9QtB+j9VBZbBbrkRORSRFdMS3uyViXXVQrLPOtPdtIZEp4Q
uaLRkoFOBapbrxcf6eH5LpD8Xz8P/rR2Z33X/Whkc1/oNxEr/BmxwisEDllXBgis
3pk72SLin2ZZ2++m9krX+qjKcsNKnf/xMVa5O3WOWx7g0951mpPtyV6WYFOFO09w
6d92JZDiMo4qNdrtM2D490KQu/rTbpP2aovSQr+qOUjsQ9ZHx4Dr4uSP3F7kwqMJ
dKNiaMwBpc4aVkPnzd68EEbF3L64BEGTZlA1SHnNrKCO7ySGyYMF1GDbpO8aB6tb
oze/d8aXVUiNp/CYawowM2/24U299ZGaygrQIN/w7M2tLvET/wle9wL46MOvparK
kpS2gUAT36Ls2DEiLkT8GwcVUN6wyy+DdmTO8wFFqJuXVAiljIu/N9IuxryOnsmZ
BfN4ujKXQaS0j6xxh5Lc6mUB1tmyxnel9QNJItHXRABx7a4e61uGhU0DuP4Rqto7
Jdv/iJ76Uat1Beo2BcCA5Ldy9iaSEl9aQiH4+sXYSvUfrSuVwODE81iAnrquQTnm
0WYBZ23Zv1g8WjbUkWPPG/wd/d/btZKj+XX5me4UDbVfuy8OuOijdtGUx27VNlN/
OeztX4R5o+NseVmfAC69jC/vpe9a66qZnL7a6Tvv61MOfi+lEpHKuGDjNU80dnOM
vWYBSnxJz/JVhMrwVW42P7HjGvc4j7h4Xz4APbQ+geVW0YOqAhNzp5kojapQ4c6m
tpaPuwbsnjN++lTIvefhaR2tAQq3sqCcHPMiFDnTV6HgqkSWOjheao6qlznnrHCa
8utIPqCLRNfRmy2SS2J6FDuaushzP0W5s2Y4DdmBYvBUtWkwwNBpILiGYghy3041
N4+KWBIkM9OaKrQUjqr1MObXLd4PsxhRpirjOrizLWlCglzj+B3967q56I6wCIgR
bXk4KDhMPlqFWvGEQr685lgBJhyF5uLd5F1AVpc5qbR56LntqmaPvG0a5KiNZs0e
7GQBYfg6UImjS0caYfJcH02WCl7z2aOVGi5DFx41uDEq6FC0vmBkMpMJzRZfpwcN
R+g4V5s5y3sxjrzVWZplEqdEAFY4GJP+Q3p3RyIoftx/Gg1EockVhFlrPHsJ21/Q
k0/8cQdcquRuIlpZeZmsN0v4HtmV3JMflHjF1mgRQDC08iUpz9+AenLsGE1Xnp4R
4WhSTBVlPPJ5OZMTmP9GSDyGCVgFKK6mMstKiOWPJOMxa8npH3YFFOIqVkN541la
dbBWulicjzKNlm8WKDqiNLUEwTNq4mm2sKm/BbbewqQ695ZCggpJhQgXWKh/+2WR
ypttIne5wHBFgiHtZKX0hrifVQXteGcmZVTVu6SLVFfbp1EKulLSz7Tzl20Pe3d0
lqMbYf7dVhpYP/tgWJ8svkK80mTEpI/ZgkQvmUzKgmrMYP0/IgTAMi7noa3Q0Fo+
7IOwhAMDZ15v9Mcot02AQvvE5ifTh49mFWk9tg/6Sk11y6SrfkUfidPEcaf+ayoJ
yqVavq8fGuyzyZjIl90JZg9S7WvTb+deI1rPwC7gEqJyJ/zbR23YPzWJU5CPYYkN
21hHURxju+p/q7TuRJ9q5b2u1SII2nqR+sqC8nd7rRvr8p0LmshwLqLXwO2OcQSu
v5889yRw/hTyRnbnyM8Rc41RI7iO0owXFztO11rPJIWdHnpRTpQD84HJLa6hQ4Mq
3VSzlAl9GHxscmcCsudE+NyO9Eth1lTRvmYchPTfdP+pL4fp8kp1IQtY3fI29WGQ
uxcy7oDrPf5QLd3Q9cvOTmbQMNOJyiPOU4AxIe3kt+lo6ZlNoY2K5fChDgAU4Olv
hUP9ocUlL6o4mVHhLmnmZpDEdBL3QWpYLZu5AluLn32BsP65Yy48vrQM9mXfUyF1
d8vWlsChAyKwokq+cRsX9BOboZdtMuAGq+F85qALwI8vjFLtM12PvCaN/fy/WpIp
C8SUoWEs/Bca6jBsMbXPtqbXmZrYJ+e5Jz9zH80C47XRJrkjgKPYZrSrF/48P05t
V155dmt3rehgHR4Id2Ca/N/pA+qutOnUeDrLRGj12BTdq49dF5Fc+0tKpXO9ARCq
Tny6G6pRgywKe64aZ/Bfs3NXOrtyLnRTscuRPJN608DM5YQkbSQ8rgpFZOcrX21O
AD7PqC7q9vyw+dNBlN7aGPp6UXka6XPcYVK6Bsp92zVUcrwkWoNgdOLUbEKo3gxC
2zicBZpllCrkRGefR36OPSUEGb7IDj/m5OO1YRYifvGvjZpR00QUfMDlRw2ehQ02
ayAwnVAyLvzsHY9Q2Q6xvClhOajMpnBR0p/QWGIBQBZNj6PyiVpQVhhg/79dyLlX
Qs/rReGR+Kf80LRoCp6nRXmQ6K18/ax4RDTnkjC+aak4R7UwWFR7Kbqbf9ksZa4O
CDD4sAZHi6xHwjKuYFYtYo3084kAK3epXRaH4aQg5Rnt+Cqa1pKxtKpdZpGqXoMn
oO7ZhKaTgbVRYqFmLKYV/QVc1Rb+iyqtb6jhLwG+Plx5jJtkwaedg8n4Tp9fekm/
6se781f9JFtPf+T8TRsGBAc4RVOs/iyEycfif1yFSGzcpPbpqf9peoHwZCWxXCMm
/zfi4WLLb1zZIDjpYtu/lRRaHjbsdj5R8+pjHvHg7XJ4R63Jn+58t2ok2ou1wpSk
BLpvPK3K5hlSo2sY1WuHdaUT6MjyI0FR/gH/3FFzB0HY2iV34JjyDzHr2RuEs32e
obI9Ed5vmDVHdG+LqfOI86pMOBft51c8u3WV8X7dHwYHM3wNs+Gg0V24na82RQwb
ZWuOWlygh7s1PE6ON6SaTotDM8w0q60473NuWL2WY+RgGB5cbSueTfHD+AJ5FgN7
AXbqjuf0hQm4suDK+t6DQPf7VKsMBLSk9qbrQvpOLRKCeCmNp/DfHvzdOjaPGUYU
VQkLZn6lJF473dStP0Fs+mKMdOwoaUQiVZUKenu5iVfgni8kIF7PMCX44reMd2Bi
5vRdxP6AZQewnbFf21QEAjvfwWzbbZ8QDtuIE75riayGC8GtImWr8SJnP7kaE2iw
3wjjOtF6tp6YWwUI+PvJMYezMzHV04/dIvsUbjTQxjR7KTRz7L4brHJhBVAnKxzy
isVQgUKl1P36dua8hLP47f7KYNUen8xSn4iMt6wzbmNpcDnCojx47xcpT9TIuc9R
xX7UsaNpSRgotNcbiwzSyVns1rnPTNOd+GudEpkeXrmBe3oU1y1DZyG9HHMgPJmR
SnoTIV+RY0SYsyREsVL4kJpK0Yj+YuAC8+8VxDZMDowLx37q5mL49TrgRGa0fbyX
NrxBGJ5/0qnb8d2G6NTFQIjmwO6hvmhuDas0285hfDzhd24FIUXsstjMVQOyA9Pi
K8KEnprGoHl0qDBuVrO7+DsBlLXDgMbESEmJWCswiL7ctDswR6aq0KkfYxLE/IgX
ha+McdaAH2FvPTgymOd24c1jS3smExCOfSRCYSxAE8cFSC/MTA+r+pTo4JZQzzQd
Ml08QSoErogDb+njd8YjMg4ZpBPDpQKwiZ8adRdaWv+iAQGY7Na1EAEurolfeInK
m1Wwuq1G6JMPD+I5R1tQPWgb6kpG2EnbqLNX/nv2QVNyxzwUcnxYegCMGhhxqzgd
asboVRVA0AMIiEBNBoVBt4EvBhZWrbS0/HutCAz9eNetSMimWI4jnj+DCundXwKu
vV9LmHCh6PDd2WsSDdP9a8f3qfcR6PSUXQaJ0k8luq31tv9rrpN/QtAQk/SWgnqE
tCy4TlJC1gdqUAXfpVjxI/BcD4NKCCQonAbhK+QLej4vBE1FnM4o7NFt5732w/EQ
4xJhIM+D3rdmVXoMuhRTPY1QJJYyPdT1T11uXhWN12LHdh2sFGEVz3aXxDrlBZTW
hOw+JcUsQCaDBWRFavXCjdnqGKpYsEyKD7pmB/aib+lj5AAZ/oYQa+1sAR/f7k1b
TNGTmewTwAgaktvCRoQRVmAGrkFGJWRtNMaHL8z4ifokOEGPHP+5rRyfbKr4F2H3
9QC7CaP8vwExaGIY1rAiEtbcu3c5YulJD7cA+T5B41QrvfxpVUhlpF3oOBM6zBbN
w8lRFiKJXroFRNtotIY9wajw0FXNP2HirztjrJRzT/S47emkwU/5RaV+RUZJKy5i
riFe39CP6GEY3ViskhoN0P4I2ftD/QofWJ5/srLnmPCRmYnioBx3W5zyfMmB0tsX
yqSUUrf53yt/GxAWQfI25sJHlyl+KFqxRC4bwLXX5PRql2vgJtYdmwrtTNImTSdA
EzL+y8+ev+LS7cHrEVigfAjy9D8L3zC2j3U/C793g1B6w8aHt8Ra72oG8EtYKIeJ
x179WPe6DnMse98gDDvwSV7K9RIVUHGP/lBD74WSgz0hFAqTkhyPtS1uAxbXAImO
Nm0AMUkKhzWgZEc2kAMpCGJyKbeWLvutIAf54bFeSkaCXRPk6dfRIBKULyc4efEU
2rZCe/y6cxAVntGT3TR0x1YgcP9xgd6J+k/BZWOFhEUqOK0iyovrRhW7rqN6lMPw
0J/0P+KHz5Y5I7KhzoqdJo7YGjMWNWpeC3gtSjqqCfE6Zo4RQCuk4wU2icRNpSDX
QLcxyM04TvSjpDkxJATmV0ghMbgOeBZYuD3IOL0zQcsfboOgwIhkEYnf3jyaoggJ
E1SpSGz0v7uT4eMUrYuNgqhxLY0dlbyn+yB8OvNbKIXLFhSBje0/oxuvWT1zLyyS
u2DQIEvROa2dz1yyFIcgNJ86l8Im564AxtkGqfeoXZf1+OLupXm5qvTheN6nOmPi
LK9Mtg32YGhxtiLWYQOIiMsaYJ7HbaUIHHblnZty5cpsYe6eq1CRgcc8TpGqYXt9
dl1kH/gz0aq8KKPkf6/LWeW+klQRg9RA4W1utdCUAzyrbsEe915jWdSFe8A5dQTF
nR00F561PFWONESE+EbCKCDaHoz6cxqbNZZ3bOyooWe0fXYXym/D5lEjQtDDG3rS
Gevy2gbPSXFcGMRfpqJRjj5RbxZ3zi3r7Wr4sc6NufLTMqZO9GPyf+sgtLxnN6Gg
Md4BEPgSjUc+YRYrjq68vvHC1mpPsPRCKsPPPo6QDJiIXZ+jHmMnCmYsaU55KoGw
griiUjiOJGSY8fiTR1nT46zGVKD/g4iJd/HADGqTOiYgq4VkwqJcvGAvXEkUOUT+
U/g0/QHI7cpGXn+5XYgHIvFTF/4ufWLUjq9yrzIHwjxAPj/t4a55X7BL95sIuOzj
kjbxGjRpdRipcE6XQvKbE3qmr79tBEc79RW0m1M4kdC0co12Z7tVgaKbG57mrHch
mIhklZyIECTqZbG3DULJOsF0S6kuc8THErM2eCTl1FppfzNs78D8Kw5JygLYWo+c
MlBh/SNDgOQAt2KkU9PuOj0XV99d+sKqzMUQIHDmNwRuZzFG8yFoq9PztBZQ1PVe
btyWCQNs7DV8qOTp87Znp0IJWvU/ghsjuR9qUItW9TvXJHcoQgUIxl5vhgXBx9kb
koH/uBOFy85Yr5jPimD+9RNYKvL38UoynzcTfbSvjcbT8hI4X70jdvqWipudI5Cf
8QJesDVzOZjEbFjrkOz505/hFEo32UnVQFsyc1894yF4uuCFtnsmKS7kDuLDxYyj
aXMVnrZlfF4RRMkhrUe7aj5zXNTd5FVjzODcCXBK+lQ9jXyuR5AbXkziklDmG4Fc
59el2CP4nyc9MCfKM9LIpwrUMqFgQrGOMABqyIfAud8uouIikO/vTbRbYuD8u/K6
eSoxNt2EloDYoTt2UnDnaH6pKIEfBlcEjbFNmhMd4JA1LHZm/wL2ifB9oUxbX7z+
8n4xfqYQBvpcwC1pvWHM7j0vsDY0LFA4tzUzNkx6vxMmlbxhyBxFEyYZzw3HykWt
VWAXsSL0E5WEBZoe/v3+1KtUtUzkvZ+I3H2DAw5iML/L148X6WsfshTB8CYrZcfn
b+F8IOS/lRpJjqDwwPxipRqb9xjn2cjyy4q7i7jm+IMrgi+wYIop49heLRtf6s+t
ypTxOZklXM/HM3Wx2DwsBmh/I/FcmVNHSHyMqNoEJ00P9nhMMZUinmKTniyZD0vl
Zk3OxTkTlFkbpU3tIDiug4MeRJ2XoCkvYaFzFRqhu81eTsmtXt6BfYOOysYGcApY
8ALS3IUq/l2ffJrxGbDPzu/2188o025DwHxZ7rrPL5B0DG+6B36BRnJiZKuI0n+b
EkA3pCEzK/4P18gGYhDonyaPgqrM+dLP0p5QP0BJXPbumSHKTziW6ruq1XuZ4SDp
pI+eaqaQC+JKdblLKmS4P93BxpTWMvmDWiUi4lhXsn+Brav9TeZS/fJ4ucb7MNlX
PlrRBBWZkagFS+P6YfcnNXLUCOM/GTdB43CQUAMws0Uhjvqo/cxK9/3Zfx9IL5PA
b1/Benfll4VTRFJWvQsMQajW5g1CEsxP84I6KdZrSQGCKF7647LxwNgQfB/I2OaC
YPcHBC58FOgk1kaLhPGvyB3sDcWQ6VwRiaxJ7XBRKC7qEsg9MZG2f3oQZhNSC9KF
9P35cYWea4lLuKCZZG3Y3pZswZZwKwUmRKCBB5Mn8+I4Yp7M7baCBMOwPVMjJQUN
bWnsK15pznHM4It8WBGpLL1tK6Ca1wgbCspdN8KUQ7H1wYsUxM0L3BLPl/CZMc1U
RzfFv/+ZQ7T6/lMxtx1KhPn/K1TyTnxEocKsn/cAkEPeTJL8wGTaktRdd7DqdVs2
6YKo7P7HzSUrMTaLMgk8vSBbOv+JJjirPCmH+ck87Ittn0S0LrGNB5mb/pgzufmN
CWIPiDxPo54X0RRkxMbNqozv2UKUFOPysDa5aDWZYCVdZ9PmcBxMtg3+ps9WFdc8
rBZdrHw73MFfgrdtjc9DIHc5HGoNkmHgaPsoxCcsvwWRgAfd+wtMRSePlq+2LR6a
G9KpAQQ/IGLfx7sSXSRZIIRGG3i5w23f/mn85ZEssTDOhJ3/2fneuqUfmec1M5Ab
BvNp4+GJvVDcvi9WyfUBlhYp5tmLAGlDRNO6HvtHQZwnpjgRbQWlm/INyzuJCVAS
y5thnCqE2orpm6c+7AtbWdAD1OUsTpGolvy6RPE9Br2ZtQYAYQ7D8Qr/IoZnjly3
1DCEDo8aDVBsVtL+pwtxP74r01tVNyhJjdqHWTTja/1itlRHCoHg4bWwbvSFeIA7
787MpiJsbD5ds5iW+OEg6Mkyrdk1sbYpj/su3Fb3Qvq4Yu/sQACjywb9lOSfJUyG
LL5393v06UJg54VXwJyRds/YMsCbcoGBeCKAHugqOpl8zjVVEtYZalXjO/h+6Lwy
pUuITDxpzOVN42Q9B+Sg2ZruvBXx9P61EyyBZPbgKnGPVSMdS2lELE15YdUowuxp
0yGGQS8p8Y1iCGW2lb6zTgpxI4TRM0XbqS9WKjp9fi19++q/9YgsUucActNvwVii
iPE7tjVHlyyxGsNt2E7jxhrbEAJ4uPJlaYfl+mhkZ/V1xbLVxv+SqHm7pMgnU4uI
lmTFz35lEs0y1cMq5Wf2AwyZGxm8NnNcV9mr+SvlnCIHCb52dBo/xtR2RqJVvrUC
KdL+u7fGAohH8KE3dk+GgAF4k8v/pC3tfgR2XjjGlOZwvAoR2edunZNUWgSgBpGY
HNo+JIrkxbzelbE6LWq/jM9kdM6beLb4Q9r3b0D9nMV56d+ahFNQo/X8qs4bknz0
H1TS9LBFWzT8nF+4g74b7R8KKCo3lZ5NwZ+EFd4qyJo3ORiojqQ44aX25XMe3mLM
Fq/sVsuGSG7J/EeqKVKxAuMGeBgHv4NwJIcCDtlsq+vgNxZfqR4nDpwtK0LIAlmL
VE0iOXxlt9IKr0mAhTIbEFuKX5UPb3aVWhRwMpFzkRuAW+5TTyZF5QuxXQCuAePM
dr/HvJFyIsAd6Yp5FJ8IDpXyawW0Dk0UJFjkeWJup76X3QuIjmYpag+hQyQvPGJE
JItCqrO6ciZYgCC7SIoIblHzOaGFuDaLAmSyYMNU9W7J3W37ee5idSbRV1TSp/rD
z0EOlQe8mFrybtBUNeQz3qNiBER5Fr2AxeShaU7NfpGEO34g7RpqlIHyfiEVfL/k
RlK/uEiAPv7FLZoIA/fBGXNxV8NTc7z9ffiZMz+o2gVLXxhKeru3dXfyiJ/B8RHB
r18PidaQ6UREQw+4QkMvspn/fwJaxQPCOC/u8WOnNY9HBjLthMdSqJvtLaXQ7YQU
7oV0LvxpI09hzMfyJDdQ61+SgEZrQ46USQr02WMwHWbA3MQY99M+jx6ECUFjuukw
HrqxGe37UAiA0YrXnAtVPk/R2UmEahNbUKnJaIthwED1YoDFZ47SFxP1JQfhSvnM
hSVtfXJS1vQ9v6+IqXz7owxHnsJGAg7c3Cuk6OcezvcfBfJBussCsypZPbk0bg03
qPJRQ01O2NNdimOrZaGbPK1WbI/US6Weq49fspLHhjRFveh6VcxFpGO5Gjr8DeD1
f5rTvdeT5zTi1fAXz8sVNiCc1Bau6tZGknJtEKy2PDsV+mVxkrTgihvNzPSJ0KgM
DhrVd3hoILVMl8W6g4R41sht66dcIlYo9hCD0CU/pTxGb3miFdaFj8uzLaskCMKS
lE0ZYNE77/yEk8u2pw3fmwZjI/TSzkymdwQBYr2xqdZb6tKkgc5Ojqj67KtXdJHc
iee54dehPLHdB7HqbO6fvd+GF5sDMEzKNylqGggxiv24bzSdpm4xiuRw0iyW/Kub
tQsO0mKdcjaHf+8j8lLFb4mGHvJbCzsVrWFGZLoezvAYNrjP53aE4joZmVCPypc9
XoCO1d4vK7AtlbjTAtrvDsmw68vKO8AL+EapON7Uc1hiD7W3yqahxCdJgRX6b9w9
clMOoOsTRTvaXq4vVm/VOM10/Eaay3XG56MIZblYEn0+UiTjAGYojTdGvNufq+LU
xWjDfnxPOlYvI+rVcI/kXprwrH3DSPmm7ttIl+HAt+Wv8bJh6vpJBZDCMaalnOyM
ydqQtMlx8AX14A2X/YLSD51I7v2L9rSXuanspSbAqjlkosbX9xZNlk2suR10jTJa
FhuBwqmYrmtUyyAqEHDoCECxeZfjffFWNegbp4rJS62k18wMKneoWC4vumzxuGzj
jrgQebYj8u7jqLvphuca9pvrcEooLjknFlodvOWle1OXQRgsBpw3XDhFa9Tj4CpR
3ErBeQ3HClkAWETC5M/UlASc10fiIMdGVBoEcwQlJENrVEOGYd4eVqyVwfAiZ+kk
1a8r4wBaJb+X3k0P8mztg70UZMYypIt8bRnmkM6LaY0X9ZjxAgLXv53J2xCUj4+l
GtmfLITkaGdh21vcz9IiEHKaYTtxcD9rzrQ4BVHjxwiBC1z/ZDzvRMu/sQCei+Xn
H5wa7AgH1JzhbA4TQs9O0a5ybX5/S0QrgWKNRTy0o+/iHnitjGLsYOa5qKhvXj8X
C+VsECD0DtS67Gz3SplQqg1rcUcH/vtYIGd8Vv+VAT3gV8AjSpAk2G0tOvKYUlvr
n8ZoCkyFUYbexkfbDBb/fYlrN0oHAg8clLnvB7LxKFMLDtIKKb5VJrH9zX+IAk8W
EbAFqioyEuSbwrg/0GNVnN+0Y8HLECSnN7FiyM2hAtBt04/GDlZv2x3b71Fmb8xs
d5hM1oPiitboLRhUprWgCGmNP0Y3wDKzb9oCNmePIXWnIO8kjj7NqE2zaihHNu3l
otpvvzNfRVEf1+s6/lacognUhzS78e1Q//bDrAgMoNn/87gvHy7LowDYrSt5Txvy
BHC4hmcC32DGBsb478fXzzEWY4X2LPBTgZAXn3oUpK4wKjebXY6zffKWzSCVotlh
o1Pzdlik7sjS38HGRlFvjzvVxa7P5L7qIzz3HnSgEDO4tCBl8cTA6s0TmGgnVqYU
B4FIQu88ZeyZlSN9XcOcaJ5TJe6rgCb2uYATlTPFY9M2IduWEUup8dG++6xZijo3
n1wcwhu0jx5bg0iVBd8VCxFQbZIXCI6FLIbqbeGJr3iyPflKm+cli3egH2FMwkQa
n8AFN0NCbyOU4l4rMhNKjHnSo3yb6LfUoe6QNk8nw8r8TXqdKOMaRbG+W+l5rhRX
EAtuiCEJa6qrx//xpc4m906DbWx2p1lE6RxDihTglYxcgc+Gt6guasY5zjBKM8Mk
NmgZ+CNAvLXRZviwbOSy34qE2NkzYUtMkdbKpfpJVDf5DWNFCVdW9WGmROwF7RJG
2XJZd0ieiJGmrqX851mEbgCodJQ8Mzqp0estQtD+UmT0fGSeVNJc2L/ZgoANsX9B
cQDY35Lk1C0bIe7Dle4jAff0R9gHCXIELCkCS8sC5nno4X8UeG3YoUnZzleOfQx4
hTZ+NXsb2uislKUyTdUMn25huhp/72YAe1s0Dd9I1HWNBMTf8J6vdCGbvCi4tLu+
01fBcA/XOHu0sM0oVcZfRvrgl7HM+fw7126FxkzNI2e57Ph5PUaC2KXeApvmAJz5
dvhh3Yw0BZOM7spQQWz5DLr3w4/xmBnE7nYkfLmWxLO2ychxVRCCDXQX5fqKXAft
DFT7bSAHC3vDPA1BN9OsBzb0mwJGJR7Z7CtDrzYSqc/tJB9OlLUe9P9ISfaxsIJO
bJEi1/kgF0tYhagBMdaQ2PWTonNZxe/KjtGOSadjPDY2UikshiRaGsOPQTWych5x
hTw485jy0iiwgtKRxNKe9H849pXSCf1Vikz8I22ypLdMc1imKIFWWe0aO/IAerc1
68JxTuDHttkfj4Xh5c6CLtdEWX0k0gpnlonufHMqLs92QGYkofM2qnlMc6biVspb
bgkNrfdvhVJEkbgicmQwPWJ/nFgFOgjfUECdCI6dQJTAxkUuxMTqmuRR4q78gvZj
3lBeUcVdVBD00F12Z9IrRM2cbNqUYIz4OZ4JbW4Y94tWJ8ZY0pjkmziiEDLeEn5C
Uv0dY2HRRSFATcBCkhyG9CHbegehF5pBe6+HuREGQaZqcUr0e76/igHoon/dqDB0
bBv5xKFsPl+Et4GWDKwF2xMxIfY95EsC5UANytU/8c4ed4roN/G87XsaCrv3ioCi
PvEFiW0Izv628K9UwTyourFnDHKf6Gp/0Vccg7HUjDNlnVQvrD4bV4vqqOTMsesv
o0uoUxrXYRUFEh1SQEvvKkBLzhs7GPLF0IBWXI3dxVPRLV8K5vtq/yWPqzsFr6wr
5gu1CcDmyUNUf06VPYpH0Km4rTL2g9O2L0fSSgFRisy5ZWhh1/Q1iwuROd2qy/h6
QpaaNJNO8Dtzn8JnvZTksGbrd7dJQzkINY9T8c8EwLvdLAyLBt02rlIdvrhIxaym
hWpzyHbYHAfSl6Wok2XlPAwh0WxKjhePCnojxTk5/q6sz0vI3nIR6Y9ipa0Iq6Sv
2ZS7caGGcsUKn+p5ZlPK+EaUIar1jbFLot5289sy0T5/0i0k7T/nDE8I35hRdrUO
JNUJdUyeQVrm1gwbBwk1/61SPaKicbBdEhCPrKy0CkbaropEPxYGhZcXIenwmIYq
P1EEq00naJ8mv9ktBTubs4sbEPwYMUPozpj/d3IpvU6tfapdexRHQfCKi+tk2HdD
O2aerBmuIj4shLwu2VskHaF5z0EMDAy4BuuLzclQKsHGRPildXMPhDyhOa5ApVpC
Tv2mxcSq/lnmexXQHwMIlZm+75Ij4b7bFUwbLWAjT0g3/EdiPJ4dCK2/8XWeMLa6
bCtlkMUWI47wkJzxgUPg/Ad4Fj0jokY6cYrOrQOs2SL0cIumEjy4SezyA4cOxJLC
yBa8Dc3fTIxWJjOyiVB5TDFWXR6VM0LYdKM7VP//4+9j/r/Xwr/JRVouh28hDy4E
mEP4AVYkX35uvZZWwISVxLT5m5X/CnSzX8lLBylMtQu0RVTTQmKJxHgTUpb3VVTi
2cYnKgnF9i1Yuoimi0TLFXzuDMSSZUErDprHCME7xwjaZ654663xgB0asSYIk4Ul
8qAEhoz5Y6YqmkR+Y18gO1JWLiZaXogriVuIvuOlLhCvxCS2lOzpt0ESdpOnCZg+
RiaoZx0U1LlKj7tfa1aeF4aKpXi0Td1Hw2JhoOEseM64VVjcntAXtQTdnsmgvg1n
T+7Sushhg4H2kx+M/KOP3IrBmuFyyUO2f/VdbKgP0BTHlfChxmdJL7zTFjB9J+AI
4OY6SGKn40GMtIJJ/M+beQHx+L9OeFDVcRRcFeLAtk9asJbSMTP98jpbHoEdP/LX
uFSzLHd27FfXyAPm/xCfiNXn67JkFCdnU4c/8vh4i6jIUnvtWgSHFDB7UsAMCPmu
EpBqdBPSUA2adYVAwFoHNZ/14QXlvSeKzm/ZjlJQZ5D/HmmX39P8A2/zxdLkJjYh
ghdLvejP0YzGEBDo+WBiDNoyUQ/xDgD11t5MxkVzfu0MyPmvBgojwe/C5DU0jVjL
DOxyF7H5zICRaXqXce29gWfAPMYce377sHZq19Rc+Z6K7IlNecowSYPbxxmyyldb
yHDXLR4hi8xiynM+ivnF0efoTX9vabFQUkGBypmdElPGiGtkB1C5eUWVpiSC4BgS
I8dHN4Inm4X2O8gSaA1H0WY5jh+RP0JXXAit7Aozqx3D72XMWb4QU/v619EDM2Uf
NoKHr8NyeDQiT6eSfnyz/XjTGBs3ipEtVvaKzpjN6GbIj6U0yy5B9VUFrXxYd4LH
Ur9nBG2twjSvkQf+rnpjA8CzCGGb11ewh0HG2i6bemetM1CMeBFsHkkPJGRTMm12
WMdhnMRYMiRm0lUomxqxsM8kJ5iEdsJ32m/02+IFP/KQi1FuD/Nv83mR9RSC2vj0
bngFtC4/FDLSohs/vxINpd/2Wu9Lio0MZZYH942RF6AfAvVsNRbGTmPHeqx/s/lw
mE3ZP8UkP2pbYisZyO4K8hpbjys5MuIc/8a2bnyofw9C32W1Pz1KS7zEPlrhA388
LpTh9KM+RlbbhRSXlPBlmB8B+mxDBeOXdSY570XRmGZ3WTUJfSTFJdk8RmSj6Mh2
GXHhgxzkQKDrK/hBK02nR9rEZvODxNeuaUXS3NvKI1fRNQ3uTnqZcT0f+ZXDvzXU
WaJUpx5k9vF6mTpC0LgfP3PJlZKkkehiq0aXtjWlqELUbqNrwLuWGNbXpk3wNPDg
nSyDpX7FEgeLR+zwWULW+5BzY2HXE9m0+uIw/aTxDsoJT6dx8k7KKaaqznhsx5k7
rzxHDFf3KLsqqDCzzVaiVAgjGaakH8nQoUKIZpRq8iMjgdYrlFnDz0iAWNChbS4O
9aM6ZGkCx8UAwzPpLUrTtPzhXRzB8yMM6weZ6QDxBKgMmfXvfJD6SwOueKCk6vPS
TC2hloNcEADZtKvx9+6V+EMFIcDjr6Tz2o/ujMMAmuRRHga7ZJ54PG82ifWMHoTN
qVgKlyCrrMOtzuEx1wQtUsiZXtty4UvxeNgVRHVTlqZun3ySc6lVFkvx1MqX/SZD
wHA0r2NoeZGccCRgnYwt5sfyWplESVitnHI3FDyYchgKu7COEM5aTCdDJVv4HI4B
qnm3A1u2uerbFaTYoni7dLOlMYigNbo38yuDB3Pc+cW4XJKpuOWNRjvUJPbcEyMN
STEi8cAQilKhvK1f9FIGgdGVFP6N6GjQTDqCyjC8WPsjJEt/ZApFE5nWGoIkf2mQ
CAHbMeAW+M9SJcYf+YcM52w9K6MNI+fqrlMkCth7PwqttChGpl5QuTdm6odgN986
fuYBdOhrwvB6qwQEYBSOVuaEJX1iJN4BwpcUbfoYWfieINVraMlcnLYVqEwp69YR
JiEaMYt8mSdcKzClws8fTWNX1SW2uG3q9bSlEFh6YzPX0zvQP1piET80R6prgYJo
STcMjne1sUVhoQmcHR4TM6S4kOb7l1eL6F5sx1fNPbP5X2nnzZT4DocpT1O1N7vB
yytUiyzv7T8N+nAPReYrn35t6r8FXbmJrYQKQ/2e274tzdasZu2n2qkaLbVXtCvR
/0NigRGwRwiLVFJrjIUurGIx5yuVcbN1W1Y4Mnu2e7S6q/qHznt6rlYWHZYX2PS6
pI2CSkzoVqVbLEpGU46RoZZjPhmKa6Vkwv3A/Y/jDNfVnqGoGYH5cBPZ1okipIo8
uAzqmKjeR442tgmlKlBvzob4aPnMrYex5wFvCopatwg9+c+Q+QINT2tdQOy4svx3
lLktjO3k3NOq8O2cVivQCTIb584mr6CI4dLWsiwm0a5DhaRLiquZCto/i0XtBwud
SNwjwUxpVaYSyoa+VNhBTUOaBvVvW6/m9/ftbEYWM1yrN7GxA+91Ig1nvneBhcYJ
2LmwNh+RL6G689Uv1WkRLLqKtzqRy9+VoZVMYQzfKPNX9cu0MtwcBIMcxZi3ggnl
kazsCHwgXlxC/OqfHISeU5R/VfA4Qfr6kFPknQpaOzWDgdRjl2CcF4Au7GV1GMob
Gam5oWEM1yXA9uEAIi84xpQ781gcGeTALAmXka6yRXWjvggPAV6/tPYun/3f1Kxo
9lvkopcRLK9c5OQBTNTRBSYHaBWYOdo2ftGKUmeIf5HX4rmnYuMGkq9kF97T1aQe
W3Rw4AtovzSuoE8GwbjzJxyBfRFwsiwSZ1HuUX6yuF0mSlSSHHmQTnHN7KbbVz6V
G05IWTufPkcrpkc5mxZ3xfwSBETSiy+cZc2RTHxeojs2yjqZDv686dO7CE2n8v5g
NFBPZp5dEoW3Jjt3eO2C7eIL60jmE7k1pn/WxaX48Chai0TtAG5dY7We4YaZPW+a
OGhvXrCJPp7OeV9eQW/SsjqeX2yIr4ZvvZPNeTmpIWIX/fMcoYEgQDkEq8jU6Rn5
9lHvmSbFjQeXRUbkFGLntJekRoOcdBygsOlgd1M7NbhaQabg4/5cAzVeQe+vcBR/
gfxdrDCGpj50/azlXcowdYbI50oEJuCz7byacbW0bZvpT0ha77c9cPSWmeym09xJ
edIjUC1COpGBGnRxBGGD8eOM0uAySeIgjPlTn6T7JFDvzldUtp+Ac1uVj10+M+GG
TIcfAUOJQFF4yoO7i3e2699OSR5MM65GMXZyYqSsQhuwtb/1jP/1oUuH9ncCvH7r
iD1fzrbobVR9tc0PU716vp58rVbdvxr6NFGAsQE+PCBp31QOukuIc7SgQFnTz8H7
uuzgouN6t5svf7eq2Uor/Fi7Z23drxh1yeG1P4RjRVaOIcLW/8yWIMFt1Bs5ZP3C
gUPkBVEZVT5Kx/AIJ8hgpNtE72/azm3xd1JoYDze+ZfuugFBejYYLk8Ow1/plb90
82wDq9gYbFAOh/5+ilGkm5JZv2L8qRwV92xL1fCWaki7vXWbJ6aK3Y/Ft5+zGEM6
QrkVkjWTeqyOOl+E4ERNWVkOx7Cts5NoP0ZEBnzuI7lLOpyonsFRbLo3eAVVz7rP
U0XNyWyJ9tdWQLoJKKD04M/djxvgpY3nlS04zX0cfioCcLedf4NycXCVccf1mB2Y
q1+InCltSIRQtJXILwUFUNHKl+qkGhdNHYylchTwgGA5qGeyqEitBjyqk7MwoY8i
oo6BOyRLhWLNOhEZL1zDt/HaPcVceLxzL+TwG4oAZTr2KaZiHgL/bSCPdQRUjJb1
7akzh9qnT/s5P3K+KDtcAv31pMvNUSMK2dH18Wcc2kyhJ2wc2cZNvi70DEilxGVQ
05qjVbt2rg2+p89SUe3IvBO+Y+YIrWRYH59ND5w9phIZDSO0zCZfbVMbqRmV3rfk
yE3ourTUILxAFuoZBlGyT4O2VT2p0i1aiDALWUs1j1duryL8jpgO4LfTtvkCiTGK
TXIKztKCxSWMqcrEhW5Yofq9xDb9XrxOXni9Ow8NuLmnDZDVy/TDBoQBpP9bcQ6M
6B4HJVxp609RG1lXXWllbctUmg69v5qRE0+Ke+mCmA2Kkcuk9BiNBa9kL6aPTvBf
d6jncRfyCGlnrle8ZXIdkpJQbfpC4SQ//vZNytKKAECT8uPS8ACgeag1sREQDXJt
ozLHAbEX9g0FRDCoED7wjwMMeHwhjXTH10xC6l7G7IoncRoxlYBxMKZWr3JHJOYO
sJjnTN0I2VLpE5Dw+VDI4a48YYLcgNgzhFq0r0re+vzYdlRXEAsefh0YfXN6SL7s
Y1NLHpWh5G/h10sso+IM8YR/tZZv1IZV2aT+maL2TF5U7rzGILfCtna6wYZxLobM
EoCFZkgCq691Fm9P03MnFdBXfUY/btR2AzcuePMpEoH7bdOuWRVDiyMYpDYq6CQD
qZo5KUTtNNz5kRosSaGgWBUBRGkmAXxhGOP7fjdesLUSQKrdgerDsE+DMw5/YwSS
I1KREiYK4K1/WbPolEGeFW7zIbkndXbF6Lgo3esXzRmPt5S2rhoEQ7a8CRuYJkhE
eI6JQlwieChUAv03hBFQGEnmPOAHkE/XoLzmBPEPodUCrkUqvMbJUyQco2NikWjf
6Y6bzhGVQLpYSBx0iY2ubiWUDDVLbw+vdeToJesi2Xe0H85ItR6PeuIl7804lE97
IPpjH+rLN5aEVxg1w2G3bxMPx6mGXCdq1Mhem7N4n28qHSaQzp5zRB/9X+piIJiV
iNd9uY2XP27bGiPeTlY4KAPPEk1DNVqc/ttfm7F+jGjr7TiGGXPnrAfIHVyrCTN5
CfEOOtehI7HZEixjSa9Pgk6nF8DRAvQNVpaqTdRJxQM9/6Y8QPZkmHikrjkKEBUE
jVgv5fcY4HzyftF5zcziv/hdrhFp97tk4/7oI+7FBRsKjzxTXnT+zOBjfT13N1No
7lXiBL/kI85H0lLrM7P2qrgNMJVn5Fx/01hlihxWdHufNPJ4WskDAAj6lO4j7Drf
yU6K1Sblkukic4Ns7zQgrjpZDs5s4jNd6U7wDML/yuL5xnPt6s0y3uDn+b9OkICR
8bEkNe2BijzSm54tvOZoJalQdN5WSW+AyLESUT2vADapsaDsS9PyUU0oula7tCce
FIEOx5g9Y0CI79iy6zq3lOBGHIVnCN8/L7hEq65FCx9yoarG/n2a6i95/Izftj8G
W0qWrmPtnqqzYkp00RmudOiP2s3jOuYuRT5x4eQQktaoIu0T5+1/3ggnYT84VdST
Ru8+pwp5E3XlC8SmDhiYHBW+PgQhflIVXhxPzLTgnNvt3HPqoVpXoUlfOUpYlVw0
aWUvkLJIPM9APnBOrPmivk2xovtMY6+oGRIg7A1h15SQ1HZTL8LoVUpwf0+fwgSy
bagbrtDiKrGRA9S5L9MBW6o288oRvzMzzkFDlR98F3I=
`protect END_PROTECTED