-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
kb/fTAM9fofxKDlGCPI/UajpleARRn3mma+h55Un7s/ulGmblgD27kEIUfbbq9bp
jVsKZ2A0moe6S6KQr1eem++apBOJ9VckHumGapvnXVR/I46z4sIrP4ZzKOsFjBTI
X4MpV6MNMiD/E5fzROEyUrIT4qcK2V862kohyLSKQlw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5964)

`protect DATA_BLOCK
SO2RU8OjfL5v8wAmk/SMsOQcbvALbG/mop0r+jgyMLonlNAoXxpo7R4+xYJZdE6O
6DvqTj9/Q2iZXBRdbnd2R/O9gpgpvRDtwgoKE2tFGTaxSJjxo0Qloaf5mrTIp87n
0UNu53Z89Pwxti+7k4iSFVG1krJm/t53kzhYk0I62u/e5ssyoUTtiye5oIt/6HhG
EBQo3i26VaK/8YNvuSp8uHcS0CdiXzzqww9xyH0Y29OaS9js4ZhV7EJL1mLjithU
gn1De6TGPtsyo3R0+ZKK8vGBj/ROkg+jwwgm4dHzVh6GDfIKqRfzh/ZKWhHTcgJL
HFagBv/ylRz+tP77adamkPacAbXkBB7oZir3MZ5NcV4Xu6l3fyWWHjq6HSU1k3Z8
c+UAphqTRoTFPRZAhXlmxfqXCo45xGgWJ5zbaUYX8SxNgeZVtLDODpTIPLN1w2Q5
2cVnFvYVinOB8+J4ejgorIH6sjllXLGMi1wQLoFnDo0MTO3xMj79oY4nFrrTM3xx
eM8o2I2h0pw2QADASE0JoXfzC/r56MXxQ3LVD1gPEza8kMB1RgipFkDW4WUJpoA/
ciFdCAjwltHUNwv4Vw1z293Y6Qf7uYBhiCgU37sfaTWjyR6qNTqZt1TTnnesHzQu
vzahBIL17Uxaj1AeEQmT7iceXxD6+WfNnOHz2pm+YfKbqNyILwHIMvegpFVKc7rY
mpwpbcp/WK8k5olXihdtWbh2xnuQhgnfK+t7SRGynaM/sKc2VbYmUmtPXR6vsSA6
xJQQNG9aJTcIPY0jmMqYc31uKNlF4Lp1h/8QJKZ18owv3xsjHlM55slwYT24CVtj
yJc96KFpwLtIOluooKJbkmVt1w8woVx69qH9MZoSE7PLKlg4Gn3R+HjG2MBNIXLh
yECcX/bFCwec0p34oCTJR9RTEbA07g86j7wF/BK0FlFeQ4Y3AqRPDgfT33pA+wTQ
k0pu4p0ZBvU1NuKsOzBfFTbLjMkIWToeHxNtWVUshoLcChJXoX/GB5kCR3Q/av4g
p8XWsOw31yS7356DEt3ROsNOEiXoi1RSP4c4avbJyTcGFZHcYg/sP4I4gpb8LldV
ryC2jK+Kw4pIbc6L/Y2WRWq3yf9wuMpillAo9IInYaVgITmio8aSSH5AziIkKXAu
QB23HIvxWz1utlu/edRnAWySePyvGp81l6kZRQbuRq0StZ3dUBkbVKYQ9Kx5w2yt
KTL3AWsue9M1Lz7eZ9vBjPdMNClVTYqq7tQJuH6rPZR9NjdWejqAHMdXwPtBJx/d
Rf9gmSJewg8aox3WFUV36mFDdFBBDPmfElIla2PA0JEkVFkt9F5YydiMqULNmgVl
tbjnLcSZtDEsH7hlcQUxH9niA4aX64APZjmmUd+W5Oq6HXhpO7luLS9rNUJCtJam
evgPhqYCayvSxN5VA05SBKxOh57N/lSSW+GyKpFgNgld6kz+ajOvdULGWCVneMGR
3LU4T8rw4btRXo3DagQNVVTsQW7fYVSMkKksapc13ujSIfC56+dTEZJn30wYKeVe
mmogB3neqOyDT4AmYwZra0qIdjVkPbget1BZCQ/Dt1dGDAHqUkIamHcRKJcpkcg9
hpbuYwLB+hvAq1yOe67UMo/VfW2HRVS4unyAsxMx4J0MPCi16tHF6gkJ8ldtgTP8
5X94kBTIdpUPtKHZFtr6ga7K+aA5fB07XzLc9nROWr6gn3FWtr0yo6YGOYy3ETHB
vBvuSU+EZaSLg6ofeyMAP6r2UOfvYqoalPEdGAq4MXlW6C0MG/AkEdK4yRbnG2Tz
1N9WB9bbj00T3QBgyykeYLL7gPIOEyjtVT+yMeVaMgx/aJsTOTSDxah/XDLEJLGM
ct9zc6PY+DLb6o3y4UsVLuV0afgGVtKC2a6GP2Fzjui2IWZSGMKgReoF8kJq6ZqC
iaMKgiJZIlws2fQvROYjt+Uw72nLWr/3BYoaBfHmEz4sLsFID2jt8WwU8Zmt8OYb
28xFkyC6bXfGRvfEXH472GbkVrHc0iZGuO/5ZjaTZw53S4B6pvY2Kc5j/5hNWH/y
DKLpsoIy5rsxhYJ5FnYwriry4qcBhdLFXd1JFJa/99tqGavywIbCcifc7BW27rbc
kFaetOJd3eU7zXHmmFZW9DWzlMpT86L0FcSxQ/03XNkK4TZ9E5dDID3SJdru0FBE
iM00DbxsdO/NvyFl9k01gJadMizLi9CTVvWtqx2nriNpdEEVauOC8P0aTAijNinX
hC141vNWfd892xtT5r8EicZkjYY5VRkAGk51H/+04sbZjZVsEAmc1Vxpz225rtqV
Q+/3Ou5ws1kRufLJ6A8PKFVemNOWV8XlXn5Txzy76+ijfUWjaDZFeZOReKUyGzpk
2PwJJqCjvsInjlIQ0gopq3AJ9zgf64vQ4Ua0+wX6Jm02CAdXoV6AOT2srAhNGFXK
j3CK73buyMKmMlTsgI611OJ1XfFNcFKcgLSF4n4/X+txhwD53NJ1u54wfCYyDg0T
T11ATyp3h7v45xDOESGgJrJ6wpbydVphxjwakmItg+ccJ7+SIcyQzY+jtMXsTlDu
ZvhhJIN9ZKmOtDRKwfMT0Crb4/K7t9IV8jAcplKBQ4er/9EZ8TZx2dkGSpA8swRY
ag752vikbh/S2FhlDKF48R/4/txCwieuPAmT8CjK6a7ogHrst2PJdcQcuCxTWkDy
2lSy1ldXAkpF9PfdqpgrVYGOulaO9wr98qfMJ/2CcR4aTcdMKOj1v3rgS45ovED/
p1nLH9+ArYXXHuivbGW2s+QeazN0EuRbkISIU0yVFdYIDTqC87YcO6V1meiTphWV
qhdrLb+3FuYt6CiddAmSWBCU5gUsVXOI8hAynIjk8xCgU11juMcEp9SqnB+vFZ4u
NFJ95xMzgqSZqijC/9gM+AYAPy1x/meZajqFrbIMR7u490gWqjGUVCzRWH5e42Kl
IaEk981WqjEl5whrZhiE5XZ1wD034q1toyVC5/i/QhSGOaqZ9gLx363fiLOuejkc
mFCuuEicXM1sl2EWDK9nJheCzBbkBIjXogRFO/qsa1eg1yQEZEfvv4GSCuXP77q5
DXZBmA8nT0uXPIfTY1Y9bB0G7AA+6MtNqVxRK7h5oTwLp8TN3HCs5oWp3UxsbiPv
4wdjr6ZkuT77HBm7QzeO49akpeO2y9uMl4z/w8TZuHpvkoO37DlnPynLjWDE2iDB
9W5x14EM0Vv7GOLiDNrjBrLrHkmSVPNMgmjiO4KnKx+qx9YdfoGaAY/ee3itIK5/
yoHOLCK4pHSi0aztaoQFGZc8OI7MipQHDrqYiuAXFSJdblI/RRdhn8OjRvboLdY7
wuWSkXUjJQH5UG24N5W1RBHnqqrCN3KnG1DeEvhJ/7JjZc6scy16Euh/y0RwcegL
+G/GbZ5gXOK47VirZQLm5gP7WonjNAyM67ZMwUMuIa2pyL2x5sE0AhQBCbzJzt55
mI5leXC0FhDALvahmVfiQXswi+PEG8n/109tfEakEF1ngQvzVwcQ55QGtAdQiB8h
MF5GvEz2Xa3VFf1SgAIpQu4rpsx76t+XVA498Ip2tEBJWpn8BKIkoxV2uM7rcrtk
uZ2NEt3EkwEEp6nR8+hDof/gMafSU0tzzrJGWgSSW+tfmiX7FaBC5lX+Mh5Ds/cd
bC9fsN19yxSEl4eEr01BxmdUCtZH1Zrx/gM227iB2T93sUHAFTxMP5HyJWQdyikH
ZZRElmAS48zePxXGUEPirOQhGz+7AmACj26/gtWUmwiU2be57ytDKCZMBcNJ/QZt
qr5tL0oXJ9IfU2TpqaNHI6MShTJJCgyJmRuSlQKMQdelm0SpsbjDHUjwPt/eUNjm
RNuLEnLaYxCc7pmriuaXCXRLcrDqDdIx7/gFYecoiaSI/sPE8HugsbVZi8UsUmx3
6NlGhP691U7gEx9NfMV0V78glNXrqfzMU34hJFsXzu+pdbFJSGP/qEzAHxHTwajc
pp7ucZDWyvTCjtcvMC/CHX/KX9girCFAx0pP0Nwyer13MIRxopd1Me0Ti0PC4JyH
RPQVj4RZ3t9d+fkvbRUEZADIj1b/3VqRmgzSDI3q23iojk4i0dILfe50Pj6F21ja
Jpzk4CL7q2VIsR8Wg8+myE/30sDFnA6JhVpy29qFQlSO7bR1V54z9jexpu54Xs/b
xcklLMpZmEYFUp2XrD1jQJESWODgKjG2BG2NVOO9/MQI66uz0QtSCiLOaOF/FRgL
yx8aZvGrNKximMu+x3KysD3iksthXq+eoJIkmCXFyLjXr72htJBgbiMIErcBZWqb
vBxrlZziCeKGrN1wLTN2V+w6x63Ui7wCFbHWW29fgGd9BeavoXb/OLHxlJatB0Ga
eH/PqRex7KeHma1hstoYEUSNI8Q15QyI6o+gc4WCwUojnCKZSA56UyPzRPy2GcQV
em5Wbt/+Q053tnlea6xd61smnXyoS+OW1wU2PJPT+nESODe7W0+tkn0c2n/KwhPx
DXIez/rf1rjZtNqqkAUvgSc6NR/qcnzr0zJQyyoIDnZyuDPPv0b1ksQvPyVRNyZY
GxlXwWj+6Fx8Fcfjox3CS41sMy0zy7BN7eJ1ynN0RKOwSHr37BevdNWseEhGCR9m
jsrudKA5pDHGqG2nJhbK4TS49erFHLnRhgW40PRaUjzU7QvKAYnGjxNlFjTDNGtf
zhJ2g7jAE1Pvl9XdppFKWk6XwqMTswVlB9TY9EiLfP8bcFO1JwT3tXEWm7GXc4ZW
qtcHhHtLmcZOPXvVlfzhZ2Bo+0cnniDb6UMDuz0SRD6xid3RNHXNBICFK1+hZrdR
5uJgyaXhV7SWiXv3ioQsdMeyyXnmo4VfkF3R4b/HUDgNL3ByYu/SnR8Sre8xu5VS
+3V8HAuGXuOnR0rndKA0MzKv3zqYIrBNnRkC1HDZrSNy2oJ/UDNF/+upYPi5T9Fm
RR2g1s+7S0TAUh9ug4Z7eZkFqpMo4imjWWmp9gWFGGkl1lT0QSV2LLVYsYTwM8tE
Z+87/ec4Ff6fX46oKBz5ZPHvN8kbICl9GkQ7GUyDk7DiAogtr8q0sF/WO0ch4jIK
PMSs3nQ8EypbIyrejegcWYsGLmjuTRuj+9N7b4VSDJ03idRc4hnpOttX4tVOHgqH
I++Bb2lwXM5TBHgkoEgwf6NZQtNANmjyPwq/nNn1/slkH+yQmZdj06pdcQTVmVCk
7lmdFxGJrL/yqnocElLqKYgdEGNy8VhWCkwt7TVdQECSvl6FAd1G4FD0QJkAVQuW
2b0LHqlrU3929ejV+7fWimdBweOB/qhp3il/DyrAYr/91NNxXlJO/jntTZgKAY9O
xhlZMSYPAJuWKwAAfc2WaThAEh8G1ups1ghcpwIhCymW0BPey4jMDVFnL9pLKkl9
mhSaEo6EuzoIga28OLcHF34LBOnqp0bdvIfSXa9Nw5cXljORcGr4jsTdJ+KICJZR
HPXjeJiAJmRQ41PIcrtbneew+NZhXbqBrTQzZkTUAAB00e2tUTBDz23o2yp/Hkal
dCEi7slF5vLmPJFgzuPYu0ATYcSQuy9bE+QOiVtP1DGgFvuXbbLD1Y6QfzvvQCmQ
flZSC3SVnvActajPu22Khz4AzmgX9bwZ4CnLcYRplH0PNmipp3TwyYuYLBhoBxVl
Fn7WPI+fJtxGIfDJg+2GiYVvd5N7ldZn+trNN9+1kQJPz3fAD+mabVL3MMact11V
Mam88XvvQpG2cLaaOp6h16fSWVNRLSmtB5QvEmTl+8RPVR05kxF3KWqHlS2W0giM
043BshsOU/KsO8zAgbA7cKqj1TfXLjLqreDIieaqMNch9PxTXnhu/YJ4t4T/bw6d
ZPLoSjsEccx60w0EbKrmB4FjzalcUrmh+QVEkE5Yagz2fcGBYiYhoGFqQ9HK/3gJ
MueLZFJ+cwP9Ts07aHSD8btDveZ+574q8RZXMvJ7ROI1V7YWRXtZn0n/pE8ZrGPf
BwryT2ffBnAlImvrmGEVXFgsu+qRvXmi7UJs4NWpSXWBm+famciaecE6PDCoxqjr
Awd8ttI57/+Y/uVQvxOUkOaFgdg8HDMUOQXdjjzXW6R9ucx4kTByRQCpbaF13YmJ
lgZkoep+iendPlKOJ4QjKHVY8Bg9wJkmOMv4mgqGEHQ6X1FWihb70YXz3ekjaYzK
ZcDLBc18mcEiidgO0cNhWQ2Q76WGHGMG+8HK26pfcAofQNz7ON3SaQBEcyVaEkmH
zHShm39MYNFWwu6rl8llsbNcdp/IsWCLI280GWLMHtNZksiLr6MeXgZp2lR5M79O
G5jftSyHc0o8srZarYm8HpsXP9yVWUABaJlnjL77ZNvhzo7S6xOGNF2C8O1bb9s2
WHZWGrua0APA/Vdr5MOzU5HrN8Ru8FLmZeJrfWIXv9b6M8mbmdGSDosgd+YTVJH3
1adoOLOt5ulZrdebzWFsQQYVelq2iehLQGHuXSH+NmymTWKHUteydVMqBMvft5dp
LoJh96Pa+rWCUeYsDxc19iJ1c/CwboG/UHvQFQqvN3kwXngU7rAmpC9VbndsxIxy
gza2UxQ87Apao3tJ9jHgDV29E+Gu6UkCaHPR2twOV/UvmEqeoXONB7x0Tno0msgq
282e3xEX8VNSnboV7C7LDSaBp3LyEuuXK9MoneVRaaJCGGDnf5PjmGt/N9vojpN4
l3CIgzMZ9RV4Ra2phF4qXTT67c+s86bKrPuXRzZhJI4vuzqaC/mIOhkzssrdENXJ
7hpyVkUzDUVOFEKokPDnVDcgntsQlmVxJy7QQJqzYWMgrIJyqONncnwTSgYM4Ry5
D0NzyP9B2LbZ5niv+g2uubMwTyCmSF0lY+CoaXcZKvmY5/SRL15WgxArRIs2t7cH
xReAY+J0zpczxXzZzjJaIwhXsLic30W/8JvshIZxcDHcMx0iXu68AdjLIoo9WGYM
+6MHhMfkuK/8fslou2RCgj0jEHIHF56g6UNw8wU9oqPwvaGVhl0PKR6G7mxpj48a
BmDzYjFdSGtOjD2oStNKPgisZ1Q3urHVpXJcjY8Omp4HpAScmfbLmiIVd3rWDcBx
TOIgACdFXEpMspDb6uX7nTpEaqXG/VLDbwFK/ikXH0R70rxWnt4a5+H4VtH4i0ZR
UrVYEVubQpFoS/8gyAK8/TQ38jG282zB1f7Ufh4kCoR4R1CC+HHCLuixIGokkBp/
Y7FrfyC5hVFcL6yKa5oOGi05gxpKXfxmRNFwh6OfGSJN5ZrVnRoIWWhGxdsaDF+f
y1Xn2vBsM+PXf060bP7R8xkZ3NIG3GOJQPRxCVCNYTv7IsLSYGcljMBHMAhfguvB
RGdalb4Q3M/3f8iLdh+obm/J2ntKMdOigyCAAXtTd0LG1f5gsXKRagx5O0DQIa7m
LATGOWELGNqWoOhuRi3Y+upxwqBD2RCGHVoRa/QXM0jKxEGfJxt2Bi87DN+dTjLc
40/Mtz3dYDB+EzNrnbegpgJmxdumMVV6vGqeuWC7DemOUbMW2o4BE7Z2jRcuCYkZ
+SOpoWXx/Or4+53bCy7dzDCeh/LV2diV6Sdtju3f9+o+0egP4kr2ab89LCh+cV2w
gvcxrPapX2Fv96QIjKT3nC3ohdMog5BVQq3wDVWlsChgi3P1A5VAdVpUt/x8Z66b
64GSObAfM+y2GalnwEnEhVLO+drZDLdd1xCt279ffnSssytn0YhYxq4LeyyysXkr
qhGSh7dRmTR9Uxn0LKntYYODdXA132YreCS2uTA6CHNFhg0gk5Xp1L9R+89Ladez
xCzS5UT2pdx2WWYGEXuVwDyV4FTqDIUumbxiXJdJpydE5ZGlYxRvMLeKGvzkhAMa
9+PT/abAPSedleBxTLxStSxNTjWE35YRU3L9zq4JClaMPd57U4TXC5fpf3TEgM8Y
CQbKqs80/IBi6k2JMz37SXWHbr9BsY5/zGe9/s6WlKjHxTqzx89ctUu0Rjnwdm1T
GZcim2woa+hM4wrQf09HH10dxwSYwVY8w5ib9REjF4s=
`protect END_PROTECTED