-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uOwKoVMt1ANx0oAzzx4O/v5vnNHnEy1vwe71OYCZHaIXH9kH3GmW0pPxTFd6d7n4GkM+wIEdKcQL
sL+9LKLB8OOtb1bILgwK3ja039siyHUEtYKBPsSfKxT9KEWg7zyf6fehkB35phhjidN3LhxxpyJG
o6osO5E/yMT3sKli9mxpHD0aUvYkR6mSHWeKw+JtD7mbfaKbZ7SZHdip+O16CtUNDgMDvCuGItx0
gjekLr4twBiVUisgRQhImUaxudfgD8zJ3xTgHCOVCjiSePsFi0xtrmlIYM73l9pZZKvvC4u0mbvn
PtLjsgEVyPQWD+OPcHzEwjYgnxB1qlCBKXdBtQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5056)
`protect data_block
xbFOMXWY5kWpIT/UvWpT4mw+2q8XNZMAlU90rQMDuoZq1iZiw3jp9fsT0818PSvwuJ+aQWV7ugXS
3kZSpW/lzWbVlgYm2cZMSpDCk1LZIPtfLGqw/5LQBTshNm7k9VxUAtpukz8vbn6a8WlJbLx1TUxA
wUCxdojg45kSksLqXGKtwOgb23NOdwkrdNvnVxcm7LhuxE/qy1a1V0C0TIKmEzfeFoGcuqaLgTCo
2R7NpabOjK9ariefk4G+zsAj2lHgyCkgObc+VMLTHkf8P+EGXg2EZOCZ+Z7E0F44DWRSEDYdHJta
71sMok57UxABTqiTHoyrG9a1mKBAKTYvN3McOIbku99VyZGYm0hnMqx2JU4hvgqz5ypbNv7YlK7M
yGaksYzOAPsu2XqexRjUE/DQ0NGrEXbqSA/w/92yJLHd0w8ZxmqnqRC67T2U1qRu9hoxHVwt9re8
yxqW4vRqsF25WEm3j+tU3V2DL7eE8tCfVVrjPZrkfSXlbATsX4bsEJx8sxZy7B6GBz/4IAV9DzOr
TCeZfY03i25uz1nI7QNKOLOvSfWud/J5oobUDzn4LvIOyrcgYM1JA4lh/m0xmAyypkncHi9xU0+d
RRFbWGT5pNWXQ77uUKjnEG9pkcLWTqsXfRivWcjZBnrMHTHg0RDGn5Atq4kUv8xE8IS/A8xH1X3N
/hMY9yn5VnDVdMDBI4JpCkKY1pvYo8BMg83BI9VKIeOOX2dv1f9m6t6Q6Nh8/JTygw2vkoAGsltM
npTIXzWTky4X2GLlVCM8+DjWpRW/h5q5bMxMCJwFBHQztXhW4PvJHc/ozbgtird6C8IUSV6QiCkA
azylRMA4UkRB+aXFDRo+QiCeYcbpFepNf1LBZiagihmBTb5bWN+UC3SdtVhb/+WOPcLMKStUM5Ba
E81GNsZz+4d9OPhB5PjEzzR1kAD7Do8NvpCGcvsdm95tiCwdjrigmGb8wkeUOavj1sEWWUKxFH8S
aWDF3AQLzKtJAnmuthARmjOTcmxL1cVfn9X2Dgqyyb+Zcq4ONa/5daNtGeAAICPjxzG5zkcRb/MA
GHKOr+LJBO0Etf7YeUxE1plD7gVA8b8AIpyn2F567375cdSHJ3QODc5UmDDTRHHzagjiLECAN/Am
ed6T8XgF/kfxwoAaYr/mjKoWGVMruGHTDOczmWQ2Y/ue9VhMBfTFDwsJAJ2Eo/hYinOaC6lpNSpg
q4q7EyR89pN63QAkUibiwdhJb9F8KhjhjxzTMMlUReXHHK7Lxe4ZSa3R1zs0bFBBvmL5SiLgTLT5
C39hF9qKu3uJpeOpiiKFeGsC5HNpM4JOLRLTFqMXvgXYoKPNDIME2vPBGLf0upZbEjywdsL20rFY
AL3CgtUZ9NEu3ICUVEG32pHgCsbywumxrKMXmj6xpBxQVINlvxidWRfxGLXszv5fdODnqJmFklzg
5+2J59OPt8bGQoM/DNQynU9niL0Sfzb5RKXOUgMxc1K2oilr1bvyr4ePfSS+Be+XsHccX7vToL5p
YmKYg9IPM73bAPilnIBMlp+WWGqKRrm9XerZ3FdtHybTwXdy8Ky3PfB9MxElE77OuKEyaNwGptLz
s/L8Z06Rnm5rvJVvmK6h6Q8EtS0AD209QOGxzHA9z1JABtZa9aWhirn+yBpgxcPLqmrxL6iiM4Ff
e52DCw/ya9JddPX3jiLDkNB1Mw3RZ4OUMRE2XBIkO+5f97skHmAAtS/1smJypGGfEK5FBatq+g0h
O54KbzRrTAq677WAKvZQQN4E+UzrPRt1F6LHUh82pZa4HJXvtROIXI987AyGi0ghhQ+Wf0AB5FEy
PRso0NDr8yCFktBk0jfgGDoumlKR8DC+5c3+KPWqMeFUGc7cZymSJgV4XfeV2Cm7UIZ3ciuLxtaX
hqH5/bAxS7hrCgRUMyWBD+TACg/kNN9nNJwELsI2rlV7sz415L92eBE/6OELsePT+LasiolRtVIK
Ar9TTauhetl1Cr7alIpwzL2v+F7TZDYHYLvShxiJPS95JSAbGgldAbXml0XFa+M+a7gTE4Xwx1v4
p5d0oTrUxFN8P03zmB/lCvu8K8UNqIxBOMciomKJQ5sDkQRRPwwyY2Rak1kyP+RU3g661X2Rty5Q
mYRX9eDk/Iy6aOEmvZtBq9mCscpws61UTLDYdGfP7O+bz+9K1PbzcbSvNUJg0cVxdEAu01n7zeOk
iPXHH+BTF+wsfKjML4jrsv2iqDmzRbupdIaCaTE5f8PLtU9cNtLB8eWVIbmParzrgInxJfUcmiPV
eEZQd4/XVwzkv+1OCx/DYROYzycI9wR50D12dBI2m/aVWYinYnmxbA5w28jet6zl4Oqv3Yfu0pLO
M4ZTzELS/lEXbxzxJxcl8WhPUNJUcOJORpP4cj2MyLBmRjWHYlXZ77QDoTkRlHF7zkmsqlyAtPLp
fA6lqgrX0RR87f+ZfB7C5A5O0wLi3XgXPtLgH9Zc35Uc3eV/G1znzJSgD5t6yMmjWWDRwcIppAeG
ahILaBl1PjHEqfBB6iIgMufW7XHuQT4ojlvvMIep95V25aUl2y7CWnVNjBR2X1ryDqRoO77IHVgt
zt1aE5FPY0H2aKnAooFYjyxAvnMytjizuFyMI7GwhFCAg9ataiUUIPC5GJ9MV1cXXQRe1mWzlQs2
kc+Irkb7bNktRFl71XfB4nI5I/lPyYnMM8ULmt4bvMfox0kapz8zxnSec5CsZ/P4qnsceM7ehx+O
W307czsCNI/8Wqry/rBo/ZDDYkUxdziIYuPpaBseT4LH4JMCjqmblvlFApGSvxRfwaRSXrzI4svL
vN8eTzmgPnUY4pDydPSP5/YmuSZTl4xC7JUVc7K0V2522h+PrhVXcaEV9h0WCXzGNdgXXwN+xB6P
3s1cIgTSoiIbY6alQn0Z+KL4thloqAn7gFLDgepwo4zZVCxBBE8CSeRIQyGrcXxWStpUD0DEYTZ2
yszwVndnjgvfu6qQEMG0ko1H2+VnqdWgvui/8IuxvMX4yDmzaW+M33ZR5IbK5OyEfR+/J1qItA3R
EXouemIbe5hV22uqZc2BqriRP5Nr7/juwLpCAWcnQipnbi2CIquob5nwOz7R39BlmiCqGRW/kMkN
UISFAS+tP5xiEJKPGTbrcb7KE3r1EzCGmIUHKL5gWDoeHneAMLTPlfN8uVkcBudIgZ0sQe0iTeUZ
9giFA8QoJVLsx4MDueyWHkXybFzi1eL25VhlTIpIboh26aRkLyYQ5z909GqqYGdS9t6m7Ivrlof3
ucnlZfZqPMi3kz/dob+wPtRrO4mscOebGhg6P8PZoWTJPcsod919YmP7OQ8GSa0gPfRrb8XAv7tL
cbeuAdetLeWfRXA5gX1R53k/pnaAWz3N37RsDxNZ8bvUjZPfeKeS1XR2eAc1RNM45RQKR/78IIB+
0d6ZKnqzT/ggcwASEwfOMWVT0b1qYy1X6M5u4KzAhDiSqovTcy5+64XzgDq7T7uk/dPPxE/TdaaE
te9uB5BlsvePie083cY08+3YvhF4bA77kHHAw8885girr4+C6qy/2pYJBEMdBNiQMCGVQmoIBKuk
+NKlgHRvZB7DroYdy7iciIVBLGvVQbUgp7o0khA3NFS8w39vOFFbDY3I1NWp2gbx6T9TsyoNIiWY
vgokriT08UH//u4i9AmiRQpjAkowcUaX4saXqZmhGx+HMDqBpb6mzi5q4JtQY9vNZJSh12xjYw2P
HpXnczS+jBbH0d4r2m3Vm6+/VIto+8eTW0c4RBrLCrTeiKt+jjxWYKOMQ9xGf9RdY9NhgEa9yQ09
+xku4WY9VasdNhJ9JbN+wq4mW+QF7rqVwuTtzmMfrg7XaUXKGJ7HYIOCCHCC7d+sJq8DsWYmH1FC
ZkDBUXR+ftYb6mPFjeQEDaWGRXhwIzUfT50Xpo2nRtfVqrXnmMP2vCrMUnA3g7IWDIsvNe8x2pFB
ckFVUNptI8I4hhrWsFTBl3yZNCLwU8Wzpbyo/d/6B8PsIobhTLuTbaFK4UVIN984dIme4D0qR6TO
FN5W7SFOh8v/xOALNzMtuFghsEW0oBV6JGuZODdE3RFDNAztC8HW7XIMdN6qGgnSBoXkZD/XIimr
v2Ngek5jZm6bIoecYLJcIE17y+zThsWlbbel/RCikMI2lyTYoIXSqINAQagAsT1HDEe3Ko2fzLJZ
UvZZD5TnA9FaMQiANkGfqr6bnX3WG7D70+7q7yqLCJpf2gjuxztyUdnJBdbTpqn5ypXbOgJj/GK1
qc68zMh8v4Ne+VTH55xNlz68Zg2i7n7Tk3NGrFEVz+yyFwbM6KHq+iiIn0CCUhzhzrTwL6IJzhu1
ta7b77p1OeYHMCuu6fbcE/hEfoVTey1VO6W2CwlbMhMCqJV/FELIneaZ6G6JP3OlU6G9AmzO+nMx
hWudYrUBhHsUQGsuy3XAU4EdnmtAd0TwdfP1DuoFVAUFUfk1KghvelJaIOXJCQNQq4DlukEVz7Y5
v5xkDTnhkqkQpZEVuGjcpsY7zkzXc5kiTziuA00ANSnwBdmN3JjDeRzJJ5AcM8FIw5v6q8qnmjLw
puEQtFP7H0z2LWWu/rpqmboHHbZHj33YKvN4Ry7F67F4wKAeCnIGg/Ekf++7ZInecRycCqfwOGZK
918+w90d9FRSb1xQuiZTCfCN7c9SsjXgkGJiZ6fRP57E8+mKqCXkIfOnFVP3NkpfVMcUqA5a853a
o4gRiELfCZfBev2RFAAl7OCkzc1j2VHbvnF9ASPJvsynsWbpb9JBuX1btqJLVsvIKE65vUPpb4mr
iI4wd+5BLWXn98pKm8aJhn28Md07KXSyCCJ7w3w7QQbCBrUtnwUJxHmOrEO+wS95EQJ2KnBQxIjo
jmSSx2Q5iGZ5dRyPzzFL2Fr3uIy1V9quPipvEUo5KtKX97igQkXp3VkZvkMh2NhyOdlXzYh1ftVB
xca5+1PU+G8C0/M+n5jZqaEmWCG/lccOw3qaF77TYNPZzuXy+PbIhuK8ekV/cErQYBTSlm6WywrM
RFEJdM5K0mlySkdWVm8rdd9uef8t3TFXyJ418E6ylNFs/gXONfzL3jbj4P0jHRMXAyw8xKhmroKH
BBPix0Wk0epq1ruAKou2Gx0wzqtjqGaLdJO5KKkge/pkXKd4mYQVtNYA/6ddj7clQejqhLigaGBI
fUeeaPe7J1f97q247H+hHxSc91GxdJipPxAyKGlgTtTiw9RQcytgVDUCOz4c+hn8cZYuiEQLfB45
Dswc4BPD6d/4Ci9immqk57vXVYhabNZyfEWB6RDh9kDL5SJxGF+fCmWSpETYZLimcdPy7/vgAfIm
OKbQ28MByeDbbcE2IA04UdQhOK8XGp6hr8LGMAWuAXnLpeiIa+0ixFYn0pGsBNpBGftRyUO8f+Gd
84rLQYx/T3shrfIFGh3lsTDHNeOqsb1YY4EL/VQs3kFssppl5EafIonmATsFgkdWHQObT4lpF4Sj
uwZ2pSOAdegwFM2Qqwvl7pRmOGfiPTxThnQyk5yQ9zaRo1oiazCYw/MXotnGxN4wE1u7J/noIj3r
XUDlnm0uthfPfykIpkydAvPJPpCeUVsJ64/ss0/zCBsUKR8XUhtqxN9we5jOOZ62RibUCbKZWqOn
+f8B5o0EvQbOf8ttE4+3/Bo1h1LonlUvKIcMpsm6nIDpIBkhfqP5EwcHuKM9Au2hEozGokY8iNW+
smQcDLqRuaKJOPHhekbI3tmqhHgG5eRC19YMivJwVHGBlqZJ+8Ta88CksEaKdTmsMMkpe7w8SNyA
dhIev4cRfWtsRhiaHcMznVIIHmeMhKqhxZGT8baVIvHnf4wrgqTzrxU4rGZ+0+nNk9rlQ7ODfeFT
qZyK/3dQBto+zAefFkoxX9qsNTN3qKu8yonbd3Vb+V9gFCX9FvOUo2NSbBmoVo5rpWrVT+Z7QQLm
gQAAUvnSC/TkTGM98Z4xiAsLIKBza0B+tPmyiDCVcC20BOVcZYLaRaNpofmiN8hpv32V0vdcorFg
6igbPFR4c9o+AN+LNs4ZfulkxWnexJ0syvMTCNxcVu+0HD03ifB0JKMnlhrt9HZzNNeNkFGNPpek
X1CYOfWeyo5B6wrdXB4QO6kEvaWpPY3wjZm611Ve1ccm+v2LQNn52mcopvXHEuimokyRPI7rjANo
JUHyjnf70yhR7iwsbZjecadN1tyVQ16TTLwlXaTzL8R7gjdq/7vQSguGjLRS0Ev5jSmBv0b8+JEC
AXwebc7vMuv/0ow+sUDFsEMxvnIR9SUX53JUCUsA4sX2s83xq1pqVVithOya0BkBe4Y57sQhLy+M
byNlzFwbBd87Pbi3XISTaCOmaFmbCJIQcSmi4E7zp3NtB3uIvKttX7OdH6dyOStwJbSUq+HObdYd
sAGywF5rZmegAm7i07VYu1SXtnMCPD2Cv7WgQWfr1cyonoSEhlSYXwV2HaS6FtX8GIQ4YcJEz9up
uJaMaxuUO8ohHdNB4ZNP0u409Gea8iSIacODNNwjQkuB2c4hkGGe8v6UXSoy1Af9Gilw7IhT1LUy
pEFRITtQwIH5UN+w5pLt36k2vRawA8pxVZGellnFCzPMkhRjTW58d/IY4LDAkTE0Zgz4hCCZZZtl
yUDxyTAX6BOGllxZFyXuWjVNXP1q6+xp++E/ZW1hjTY0ZV06xqA3k/upv3BN0r1Mafn5U6m0FXGp
XxzR5xRooIkaoNbre0/a11J8DNq3clQ5G4dcD9nZaaBGGDIFOAfOUg==
`protect end_protected
