-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
4/wn1njKgw9FuVyebQxqzRIffrOjL9eZAKy2l6a0CUGSvu9Qh9nrc6Vbb/PpOjQs
ZUXOp/8DUfLyoNuhLdDI8k6D17iY05p/YoXONF6AtleD0YR+BmOu1RRqStSRBUVr
5T8c/lsfh3HLvOqL0TbzkqVf1R5w7w1RTg4K1wWgTrpZYVtdXWTK+A==
--pragma protect end_key_block
--pragma protect digest_block
r5XeQWenLTDYJn9MUPNWmYyurG4=
--pragma protect end_digest_block
--pragma protect data_block
FwYC997ZkOAVCbzHtY3LcajBsJrROxMvM+jm85ek0X4JYxKQp7OjYC0YzOFMIff7
6HM5j5xbPe9P+jpnN4cjfhEYB1+3ocUJOJJDf2tT8cv0+hzILSidc0hUKmxdzAcv
L5pZuEg+OmCLF8amDoFXGfuRfZ4h2c7cR9c5rV0blivayqz/LpD7TYx1W/o/6bDD
P2+1kEYdKUSxsMxpx5wEtvKR1Ff/dopoqVT26MhCaYpdgcvk9tAtSCY5sAZu1D3G
zQNBP68N6S/UILUOrLKSfGeqtME4LdUmfss27Lqpa/1J4fEOkWzJfXX2C3qJjcIn
9xY2CHdjl0/Ek+hVM34AIPyZZdT0lq5YL1+kZEPF+5wgyhYcRqwWRZXO0iE6BQtj
XWHgs+tJUbk54gwtzGSF542IpzdHPROBGpTOwsnjRDkYBULaE68N/uAZj+DyFPog
bLV1p+aluYH9qdRCOuVg4RsHs3TZ8oxZ1fjE3GiW31i+bQI7/IjxbaXfFNdRBXc6
UuDS2s+Pumh23C2wHDQVMJLRFoiWw4/uJvmclmdLilP3+6gqlu1KnbZCy1ueDAtV
1WUBxnxDDy2w81ahMI/da8zRaC2pn2w03rocMTtVhzHxvt28hpxgpdJKaTHY2zhP
IL23RGWqyw+rcttWVZ5jz91PftbBwScAN/3iGhK9LJ5ezEOhaWbMl6JlCFnF47pR
OdnrB0buNOY/y8b6IJL0oilTVt307LxLZSsViD3k2rYJMd9UNoQTXP9ESKksPDXL
jtSZsm8Mad5XpOYXhUT3YD3BfCXF9+MMsUSDgtLBeT/MDzQa/wLNQ/ae/jOD5GMZ
iH8am6drt0MPxZdmSJgAkAOlOYSTtuEnqnYOWLicR6X8M/UT50mYX3QO8oEi/7E1
d9jan7PI6WWKQYG2c1JnMhFSFynBM4EMHGu8uBLPWdECb930Z8nhDfKOlAMahnKl
9lwRwgcFDeduZPm159WgIX61aTjEO06llPIgiVNFhFbptLNFVYV+cclgvlrtH0Nz
VAUBbv4gHwYTHayIs7Qa9z0PgoVzNHla79RI0LeLljbDGAYViC4I7/OmWAKZPEZ5
nskzzE+wiIQcGnRNC4+Yd4gGmI8hLw1XonEBR5Kh9TjlN/I9htZ46tDvVDt628Q9
UMIapp2PO7POK3UIVpyyUrSjeChx8uFbOEqijfn56DyaS0cjlA7l6QDx/nUfXsdl
APKJfpHmZRGIfIeg/XK+fkJagiYKJImUoo5I64fhO1EsbL+53fgjJ14RYsZ/zhdW
buUQGgk79ces0Y3sbXZJboIKkuyfN9OLGS+oU/xp6+6eQr9blrzNb981RIELyKH7
MOtGY0T6Ww7IZStVlv4FsTHnm2w9ALOc8CnPGA07SqACUXRBlQkRApTG6qjpEmnk
t23wZAB25hW3Bwhx5Y9E1HZmq/yo09cFYs21FdQ9y4sHAdF1edh2q3u50WgFPyn5
CQYPPpSP3vzmmmamB4tkaF6qCNnZBvltgxBk+owQrSo4L29z2iGsK3K/IDOHCYC9
q7L6d3zgEQrm/XCpLSGHAFZZjsoFRogIipSoeYy7e/czDlVqx/sNFYM49W811Ffk
7hJNk6MTkVm+RyGZdqlKfHJMVocmxKyw298v7252Ak1On7XnuwGSNut8LsWDU2AG
yq0n7zeZP25xl0jPdmAa+c6OiH4w1RKsbGXSQrgH2WV6RLP9M9CWDUwtWUTz2u5n
guOQY/ze7QjjLuW3LZHQcfA7eCD0lcHDNJZfdtIEXvTu5A+n9i6A4iZs6L6Db1Bu
d0zXfxD1K0hxk+6QYN0yzs4zNQiWN86FfQJTmfL23mGEi42z+8xOquWKs+z9FHLn
hD0n48i/PxaWuVSc/alvyqXsUcOc14yYU4bdGHwv5jyjXunTBC98b0FRMMZzwP0J
WbJ3w+et5BBWzaz9SkD23DLipWPb/ONZCsWahHdSct60dgVfr3N5bfMnL+Kr4Tuq
xPIjbibCehCYcIFLSHe03J7DEBO/6/8yc3dOyAdXDvBrZ4Iy1QvYHZcWVkKFRKCl
wgMIZahH+OkwyjNTKnb5+7N5BvIxWhV6P6DQY95wSwv4x2Y/ETOY+F8ChgV2aQ54
cwR/gGMD9w1+065yhHhM2HymQbEbJ+XMhuefBOY7nCKWyTMVUIDhDILZvefSct8b
Q4MiMO9rYjHKDuwZlmIwiSYboo/v5aUcthjJChJ0wPQ6kxyZnnOplsn4uVD/zF+5
UHFDZlKZVqT5/MbTRuzIga+Uo765L2+yr5Fc7lDvndbh825yR/JsHMCaG8fJ1fM0
cviYMc3j5Lr+lqqygxoZkkGur5tLxEnu94UzWEvQ3mliYs+/uR6Cuv+2bwYWfc9V
r0o1a9BonB4uXtVCoHGUQ14kPTUW/fWrIzK8ECoK7ohmjDes/k43u/uFMxGJe70W
svLmfCV5kOBzal9Cu48bDawKQFL7p6V/S7CJXsRKzncWEJKX/yDb0NX+BKthwUOs
TNL/qO6gP4UleHlgTbN5s2PDn7sbklC/do15kecBBejW2cpdb95STMW0e+4wTvUp
o/6cbsiwoiiGNYDsItQl01pex9rlhk+anRGcdDlLExoMsrYeaQqTsklc06EqhRtu
m2bJuk4K8vUUda/nBr5qhwJC9iymYdulfO0qkK5Mn3s/iGDpVqZNKx/4K+GTej8v
/vuW898S8Y0uTrinVGfc8iFzmpJuFq2ym0MqwxQ7iqTABsZRxcezcBZL87TGKPjh
Mg2yVaRf/Gjdsix5RrF3aADj3uCc8ohT9C1/qsSf9IREv7ghr7Xq16gVps0R064h
fcaow2Uufd6C97R/kWdvv3vtZf3d4me01lPzZ0e7bHYHb6kx4AjcK3pKynah9+7l
8jTZyDVIZs7y8fo+T80WjMnBY5oBJ5sVzngC5POLi/UAwj+OdsbXWwoFaZF764Ps
2WgVDB2GRIRLyfxaO+GlKYbWlOqgLttNCj94gvsAvJN1azIJcAJDJwap7ZnhfXIe
q5WVz/C4Zw49H3nv18ZVD7jqOMciDj/eLNXUAV/Llxfl8YS96NQQvCtmnsNQLHuu
j5ltgw2wVB/m8t92JXAh2DCYJR+8G7XaSyduOZtA1pZ5qhoGdKwSmlses8JQ/vH7
atH/LtFuzW52xRx1+PCPFyOYVdQ+UG3RH60EDJkQ7YWpWke9lOB1IRDHZJEr1/Re
zUqgpyDTb2bVxbzZZtQjmCfbyuBLr1ch5kRo4IF1/Qc2pj+UvKC7tow83KiuEYhu
uaP0G9R9FnO23PKHhSfyxr0Sp+ax209Xv4Z5JJohrWMiP7smZusvV3r3Ha2L0nVT
uDuN0MnHy+CKDz/K60aTrlAYzrEyRdifk7SqzD6YdhOpeWt1g+j8nRZul3pLaAqd
3N6T53+gCTwY+Vg05U1iuo7j6jAeOOMbRxAwvd8fJVoTsSrokiaQjfnH8CCpRidR
P5s7lGNkOWSTYd4gOtZ8X0E5eayDlt5z/XAEx2+BtAro/3SnX91JdJzeXQ3SfZ6P
+8bPQbeeI/3ePHlzyGtb5fim5bdEedxs/nYTppdLfB7bA1JtO7iw9sCtYtL92TIj
+oQqGABjLGIWXlJbdb2yt4Rtnd/PMc3NpINNDWXGoU4j8TBRBe7DupdfT6aASbm3
yaHEcsqtCNk4Vpd0LTxEc+CtS/ZOgjXDnIziaQCtkXplcRfd78QDjmIakMAi6gjA
5FvL5uWH7yzfls51Wr2hyTyqxLfX96Ub28Aw/jVTjEau6cQ+9frSJXpWZMPakR0/
OK6O+LCHMW/R9kTK4JRqDFdrfGxNXB6dyv2PHszcwvPITftulthjBPmTQHfUw5uM
WofqaYbN7T8dHbLPaTbzLBiUHEji6SbZmHY6dVCIELmUYSdo2erh3FX+lPTdKh1J
OXvXesyFvnda2bmMs19D9ZE4u1MzFV8H8yF+Nb0H1Xf1Qpa0DMu71oj34oHuQD4c
Bz9/woCFKRwPoDDpW1lJUU6w+OZVZeNa7x2mRPcgXNR1SND0KfBwxSyahUNzG94a
4L1upTxkik9S8nWCMzzV86eAbaMJJrHb18gf0meNqplsOJwAM1mKK/jjA+nD52EJ
GeYLhImtrLEipnm0q0WxyRm9JZZyLkQywuuAU5VYTnBL8u/OxVJl9D2G9YEGUpX2
DullInq14G6t5KbKIexaMYF9pQMjiO7AKvgAP81RqNuMy1bqLD8EBp5HRQfGsJjW
8yhAuvU9GE5PdCsoBjyACmJyLfnrKGmAA7pCw12v/ETvChtGl3oc4ERrjWO6lq21
+dHfUu/vtpV8u9DWTJrSKCxYq6u/bS2A64BDdpAeyiTR8i4KM7LaBhs8EtDEJ60N
ZfSESJBJuFhvbrVWAhmuxWeRV7n8eeT5kpO2oGO92Kb4WZ6YN3DNfx1Wf8H8HTEf
O0Q4YSrSlb4DMf1ra1WOnCLeCzLlf0F4nZqmPHDloQDOo72dl7CGmp3SzaU5fDXm
Czob4eGIg3E2zmtj7WxABCKg172rh2I6wFWYWq0h0G19MYE4Q8G2K51u4IJwYLLB
GGxQl/VPHmFt9Y6wusFJCEHg6ZDS8oWXOdeYzADb4U/IOpE6uM8j6eqEaPXXrFkQ
UFFTsJYlX7wH6vCDL21OaV3s4o4OCi3S8gihuXGX4k/CziTaCI4bXnIwcaTNohk1
NUharG7KujzVzb1OO47hvp/gY8Tsbdbu7Xv+ZA4z2shPIZydrPGV/2yBISbROMtF
zX7idEcdnWfPjHEJlPvl4ogS2WGKN19X9oSbBNLabxHFP3e5rrDlUOJi8XhOWo38
yDdD8pMkHEunBFGn2xR0/D6fmBl3y2ahj0qwQIkcpUhmeB8y8kYzfuNVutYi0vsw
3CF+SqU/9tnKp7pxiJgiZMpV/MNyUn7B1yWCAc4fz0vtXk3in9JDK57FzUlySX4K
MqPDFMkZm/nDLFq8tpvKfzhX/7WetX8Ba1brhI14pJPqCnbb8O2cDKhw8zysrMK9
nRlJiAEp6lrhuj+OE+CCzb3whEVjB0ijizq/yFrGDVZ22WMbTexZwakhIyZMS3mq
bAbtRC0UiAl998tPYxEnR4nS9MgByaGWV7R7Pjko7Cing+i2uhVLIlWOWxfdc41i
mpzgjVxfIrGXp6+f1/NfU8Rs757IGktwAQAKvi8Q3rdRflTyco9AbiEBiy3oy0I5
00SlvRR7z52cHorrUv3RZwWWYsr4cyt2B22ylhArpGuTQcjSGFs2eU74q+M8P0OW
wfBS33PwsyqRjuJigTr8n+ykd6dtUT9YZqom/iWwlq7DDP2ZJDCp/EvH7LN9AFgr
rxRjNcZdD/ngapx0iUKzRDW+OQ37d3CQeKE/i2qO/HJsHewqS0cX/vOJnWnOkBj/
5X38Cux/oFSrdk/uYJM6tMkGdDGIGfBt8oeQHZNpwUpPGIe+1N+57Y524V4uS91/
ovV5PsgpRiy8qt7ypwULRGFVCsFySvcKud8ENA3+Chd4lWt+OouPFBR9SjB1Bhjr
wC/ufG9uN6UZNw7qmV6oSUGMBCnEViGSzxEksEW7RZHn6D/w18anrqGslxCLrjQ0
PyBYr7ias/RQQIf1t/LRJT3xhahrZY+mCH4uSGPOvChQ4+kaiVprBXC46Y2LYz0h
1Q8AZ7K30RH176x4Zi7W7pU4VxO3WIZlweq+VEZk3TOFr9ehA/fvB6xa2FquJjOd
wqmuUgXkitpx37iNHmEftIOvCxWm+qCutkR1lJVEaohW9FBDQqHT+D3MFm5YZPwG
hKyEoz5O+iXfCS6bz1ivfZOcqa6ALO3ySQtQSW62g+vlkE/0uI4daJeNp+HNkVk/
5ZOUOt/Mf3BGA7/rF3qSa/7yYb4IEQoBD4+7MCnCC2j7ToRKHh+qz8Y1SaaXuTa4
1KqVSsgR3jp8JPzyRUZMRfNw4Ju2Ee+kgyIjJ9sc9xmRft30c1WbZCj0anbZta7H
rnE1DaUsfFDBMfq8NHXS1c4z/VC4pdZ2uwxNWthB8qJi3ck50ozZppK5PngU4c1P
aVtLsr5bl911+rJW98RPjpyeo07SbVaRD2NgFEh7K+kiAZU6jp5gnD4SClj2fsoL
Ib52sbwmMMbE8+VXg6L54bZrJI38MIXz94Q7mduS2QrCbaPu16Mqjo15VUt7iUYu
Oa9M/Pivx45LoGljgIoyT64hQi80rkk2fk9MBHObhm7CMBejz//a+YuStHtgohYi
qCo+AuMsTHF0PLz9RVJfZYLUKtz+A1vXOGoha+SL0WzUEvZ5kfPx/Zzd69i6pqV9
g6M+GEdOfUFBuMKAu3pUHeHfSLqk6hIM3f0+orr/MFh11KQGigKZzNQlfp1ec6UF
PUyslCYJuHeCt0O75ew6aWABr2+dcS+ZM15TzVQmgZvw5QKg5mqo1reJcLLm7PoX
RPdhkJudw99tHOk8B6XWvuc1yRwW8TZwsSD9DwGku/l/dG7gNICOWAZsEmgyTp4X
yaKYxBW0aTDZkdjtL8wm5SxOunqLD5EEupyv0aMl+yn89pFlBifBmIcQkr6b4jcU
3rCiqkRfcOVd76OgpEKvUNGdSgWmqguSJWYDi7eiHRK0nVyAW+JOsTHNbydDTuH4
TY7lEDiYjPMEslzjNgyY7HOIGlC7iwm1i41d2pV7eqNK6PXcdlqPw5AeKSqKtN9U
icv8LvyxcFresakxOnGxUQRyKT3qPm45BJzryeO60nkA2pgv2oG8QUhRQWV8SQQv
zQLc5C7feo+AYGQRj4PzMovpHxFBEzLCzB9UKn0iUGp7rpEYqgGQs1vsD6yk4YO8
tQjUeIYhWPjo4+DERLOoAB9YBegVAp1wL+kb7xkmquClrJdu9tyX1etI1PTeGiW0
g7bfTZI0cFTXDmJwZYscH9Bh7lxE3VYwzcsZOsSae6sAIzKtDcBhbfRdBYPFf64H
6JGWU+nR2u00OUTpA+Svo1v6ZN8AzNl4p+VW7kVQIk06ORrRqglr2pk2Ir7WVHqj
W80EILyVZK4/zLXfv34r6stm0xitopB1Iv6WkKsU1Jyc4VE7UXa9+ePNCx2J9fap
lxp9FKs/jRfoa8rhejlE5l4HMF070QC0YSPmb8LmhrAwvCiozDT7cdD/917TTwVs
TKrFHtfN5hqwMF4voQWGLkGlBp1iQsNgtJXstcQmWUdO+TWyGMzNvBLdr2Ul7x2N
aWgjeXrQGe5K/hXlSpdn2d9imbWzWnfRZ5xIvXJPwDcJixOeUnWelTO+92esyj+o
KVz69sk0sTJ1UUjVWvndKVplne/E1sY/sr6M5eTKTFSnQrWwALl61G5+U9U6QDgM
4VydPxLxddx3/ItUBZDtowMlMygcXEBplMsQdSxziUdmofTaZXh7Cp/YUYFl4dbY
FmRNiXHaPVqmDJ7KJwAMHBa4qBrdu/EfqOv+Xp6Eqe2Fi+x1XJV+DFXM+Z+fU8X7
D07DzNkvFCqSw7RNseZL7DU4JWM4+O7VKt98yCIOSyBKTYsoCWk5QSUcLtihnclu
wd23an8/H9Vi/xXWctKurSjP3+qmsDVWVXS4sUkBFUGU/yahi9qoI3O/llPaPQTB
zJ4D+LI3YQB4qjpvsDP6XpzctpEfDfi16kxU9QZEFhwJkkhT1cEcQDesFrzk7rOp
L/WWTJL7y5V6fr8D6po0hqSZVnvdPjBK1u7oSgYQ3KKuk2gB43OmY/zWElx4TncN
zj+z6JSvXy2RZyNhY2WHKik0eWJKxlV4ZcCx7kY6Xu8xD3pry3tCY32qampIbiCR
7ie+Qafnx0YBevzn82BTpB3LlzEt9OO4taEKWezuWu3NFi3tEnRxWW54BcJVS28k
s538OyQ9penQ57qjISRtPp9n5HylsDArBetyIH1ro5To92lXuVFG47HQgBciKH3y
VWv820OwDW/ifyRXZLKmEQ4Zm81L2lRnc/lpBx41uLC6S+5416/K8t/wt1HQuP1A
ynseLgAX8ULP8fGJ7Uqpp+/Gg5HfrvtAvpSaNLpRU9Ub1py4gtouefw/v6pDkRGZ
kXgGqgps6VgwaB3x8u4LIGB+7+z3Qijd2bJXk9OuboQW8CESxAiZYUHvBJk1QAsI
t7eRut7bNlzUlMmrj+KzgNSQZiHVZXfUqLMoNUGuGZYaO/007RussCNbafTSmwHK
hA4KiX/X2whhyeKr8Me71mIGf26kk8xeGZGTSoNsw3EEEBjvAI1IcbYQJ4EfDqM7
p4OGQ8gjlLKEnB+/RJ9PGW98Gl4YI6HyYcgTDQIqGI+aeESmyJle3VXCNjvHOAMb
G3LzWmjgHRYI/fj+nNBs34mypL2CVhNVsSbYit6AAaPRkFk6ZxoiQtwXpNYlXB28
P5zERGs1/QveqtupU9cBqulP56rUTz6zhSN0XCmAvXDsxJcZuAM2TDPOIcJaazDp
6qWenbBJBaW4rs/SD49vZXhiaZqC21WU32WC3AKnSRjRqNYDZNOEMUr0xnoIvSJG
JKIolklXjDQg2XbDEHHpm/6bC+5nE28vtTbnE7PhjlFzr7v2zlIZ4Peq07DhrIiz
LHr77vSgTu9azAELjnrMDTJFQk3wfuTrHjRwcdXgO8mRHcMJZFPjlcMgBVL/i+A0
6GCr3jqPdKb3jpm2ubXMIuKqyTtUZETSyarGdnfLrZ0S6veaFtT+Z82LiSQeaXtd
7PIiYL8rd/Sb2zhszLdWIgssSiMrZGUExSnWNHHCGjL9fX58m/+7SuGk9Z7KIPdj
lUlOYrI3B23S7J0ZRJmhxZhQ7R/lD735Ls2mhyMvwUXPt7P3+JyvFP2w08333QnK
lTMREYmvASBvyK8ByflViLnkGYU5tHnnIcwZ2EBSMR22zmA1zYlQ2TJNX6wp5obN
jGkGW6uX8ilJfVUbLlnFBSCttxUOM4Z4sNOLvwupTrYZuVloHuw8OErsz3B+yJ0X
gI3DkhBQcVUwI++wludOYB3LZIC+vJaI0/0xTl+nRD5eDQjb/i48M8a4gsHECN6z
QpL7YyJ5IgqmVzLIffTr9V7N3WXu1Y0gYR2nG8c+B/p1dkApBdm9Vm0AwxizTEYK
evmvZUBW/3t0T9Ea3P6R2uPVo24pNLerc6+sky3r4qtAVYpOhjJi0iygnFONQ4pt
JuHPZIQZ1AxvwxhizJYrSeTPcdqSfo0/vh6/d8UOoY/jxQevBq+AtIy9Ul/5z+6W
ffRfamPz0n0/PJ0voo3QlreUrPSWiKp/aHwTew0jvEPu4vl24cf4ceREgFsCHeHb
CaJmMeMQU7hLKg9JGXIqBHQT+Nj/BdFLcgWpxHrJ8ezQyQy0HiRN8cYuDIw80CwU
fzP9JJOXVBBxx68hZ+bwiqBJvFO3XIcLp4jvXOz5+PZQ3gjFSLfMbZd150x+AaNz
R3U8es3ibsq/vdcj3EOYDwftQ/dj4T3iFfxPLq+BCJeYpMOMGk5orxZCmGZW1+lI
mFyYtzv4joJ8iAr51woxbvxctJtRNakf10/DQ7GEAroU/+qYHirVkgVqraYe71gC
kB5+n2qa/iVf8kR2kI4Iaxm09274CfmCb+4Hk6BKgBbatohOHg4IeZNl7nzxl0h9
ZX8o5Wi1peBvC0vYaJjjfqGuzGB0uaj3hP8cjKhFjeS4uGT3wCE4rVMLZ7EiCAQ5
d9vzxm9Kiw9TZqUH3XiqyqrlzvagiC3Zl4Zv//5MLlsaPjHz98oQiJMuW6iLrR9s
yqbMRUxnFWlsnqObTS4d5CSAn0XjKkL7S7DlvlmKn8TFREUbxdV3flabHUS8RGu2
upcR50tqzlkAWL9WWczaoJBbLZQqZfarUiOs7R9o4EsyNm8SfwUeYecOBhT5TM1w
3+lXucsupX1Ojz1TDhthyzeA7bjMJQra78+SZ1z9HOlsyqdti6ae4mqXXnJOSlBg
fcMDdsB7ajziDye2o80QM3m5o2ETmsltzrHIF/muJgm6vX9cw1njTk96OPkUDw0O
nnYl3D4888KYbIngTB7DR4WRlTICkSNVZrFO5uAV1MTBce3/3pjv5xbfoJXF8m2m
NsPdg/0/3XIRSrdvtxP0n3FyIkbtv7XKbia2LrJMotaETuKkcpjX1EZX0RiEKEs8
L5Q7ULELuQVVcgQkc9BdWl/43jhJvA++/UgiDTdORm897OqZf5tbaJXPu1ulGlvg
eocW77S0ASx/vSwogguB5QEacORDksIgF/N8ycSkZMJpH7JL0YjY+UEYWRGHZiCM
VXgZJqCQ7j8Mp9K+RZ+H4CSSmaQyRRL9uHxbqqqkUSEk/kvVu+rjE5LzPBVxqmWB
MMBgDVhy1psy/Ohw8/ise0S8FXS/uKFEcOeGbqlP2hrc8ilUelr6aRznc40DakFe
nxmTjBNz9/UfZW3RXx3Tq8fpeDLR6J5nvXAdqBPUJ+BZZUq764QsQARrjwbtZasB
s5dYnf68zpjQf+QuAIRYUUn+SUhmlGt53W4w1kuJrvLTW4zJMpGx5F2mVKtWaU30
J0PcWPvCL0X3gOG2iFZy19HwefRYF3P3DTjClXl7KSzoquh1nBx/UjC9oQGdRwaY
EHgzNWD2QG14pPXKW5oifasEQvrRNvVEZrJyqvhtbSC4YBWGkRF2L3asdia1Y+Xp
bgMAVHMwHlyK6JfJmtbT5pgr02HC/w9JBBW2RHwOa37u8NxX8+ltgALXY46S8hMP
nhY6U2NSG5gFqNaWqkSSOGng+05jIq2TBcn5rd4SN1c8OHFlcmywyulN4T/JDkxv
Y1GRK5gU88RofOwwETxtos59cQG9WwZYVmXw69gdZ6mxjOpF3tFgonH8s/aGwfZ5
aeeWaQMH1tdNKHM2l6ni7di/c6wUtRUuNoaNVQKExQIdoqvWOQ3I4Ctj0y5Wu2eT
J+RoCEFetCKRXlazNQLKbAUvR8F88kSY9MucvNxIOC/JhQyQUvXY+eJ/ZMF+WA07
bFd4GGViP9x76XTe/UHAvOGPgmktKKR7B5qdCPEJfsP+DmctJV/dFtXHgk2gecH/
ek9dmmd7HmVd35qLCnXNAVZZRcf5nnA3+3ggonHjF42TIyk4tgkucId6ywsJhXpS
InKYkPh8syuJXOwtBrFmzkrgfTjMdfROXtL5JZlSmdFxer29hKxz3NTZJZHUCIJ3
FBaegTITaJmoOme39RRzV6BARoWMsdHXWLkLOXymfmF9Mek46e2i1CcFIcTey0Qc
5w2Kei1M+EvHRYafy/Zo6OEXkHfGLyTShPGXz5PXYseNDDVgHWJtEIKSpi0ekXpV
wjrs+glpVjmkTE88UxISZBpxDGU7ILnXbJDrwv5838jR4bU5oe3r25XWvMjZt+s3
Ro1E+3WInLCV5e//PIHNmySU/g4LV5H205vzFFhHErs1Wli6bbh4kFKxgiNMcmnC
++T3GrSgw/URAoe1ttxIJ7rEC/0VWTSvX13O3+vz04evRpVdifZLk4Gjw9FiEYPi
lQy9FjonUHmrFszQbRoJJp1cbe/UdPVlIrCHfogK5mMBk1HaWtdhgDf+w3jPy0O1
BM+ntYn3BmTVGwydoc3sf9e5IAmofw465mQ7Huj5nEtq4hodZMgf66nV39KIecz9
mdCG9fiaSIOrDFWrkYtDBpIrbAbRzOcGSP3uHxoUkJx4GuYMaBGRy3MKTbqw7Kyl
Z1xmZOrerIYHimK3frum1b4plpub7BUhLzxlyAxTfmdGURo8q7XYt1GJGnuRcUiH
8CQTF3KjTl9nGhgwo5t0NhsOpZXyZR3TxE/k2rZbyW351rb92MVRAkOM/mjvyZsh
wpr7Dq0f51Ri10rKj6cEpVb6TtpfTsDeUGH+ImvWUe6VHGytAiZcFpVfNfZajGc/
jbAe8XMIgGY/GfzuztE+qwBPh7JLqGohpYEJABqWQTl3N0G64RbKlb1o5IRn8VGh
pdWD5Oi+Pq6sTTM8/gBY0xclN3bXSSp1SRAqe1wMnEdvu70B3j2qe56kFyAi66TZ
SiD+k1wfPLpp8bp71qFHo2UGR44G/4SgQOCVyuqkR0ooLzBcC2dbk5uRNJNvOLKV
jzwGEa+YOzGrf1PaANTyOVA19TIwskskCdkNsjECTboMvyNZEe1vV7xv8qLFth/u
A6DjTz0LpGKWgOBA2cBVldQUF5wb1UaD2+L+9HxjOT0IBcA88cKqeGHyPD1c/yTG
CGtVaH51RW/UcCMNfLRtoG2GX+xtAy70Dp3J/9UdmtER6iRpEOyqqAdqf4ckykar
e7d8m3s3Yvwteubo9xqGbIzpg1kN7KTqIkpBpfYQvnTXLgjwRgPV0zhnRPBdm1Kt
+rXGnkxclKTZ2qWJOpFwRvVqh+6sD+ZZDS1k73xwOi5MZcwPy4ij/dlnpch3W783
TzkuWSrEKefFSQRpM0AgBEwUke3VEFePYqZJs1gF26Zgy1DacjOic0A9/h18oGRC
B1p834jPeCs72EmyyVhx4fO3uVBGL876a0sBFcorIJ3IZ/pzXyPZzKBFJaEVYZml
N0W/uLMzE7SfTzK4r0q9cCNcj4eEEKs1Dpb1EjRHjLEirw6gqUDZOaqPM60ufuaP
Gd53hZe24toE1qzhryGBwv+l12quXfi7Ukem2XCuISjHY+EH5WLfAsUwMKD2FgeY
AzMargRl7EKVjg6Ik6vzKeF993l2mOtNAYQ3HtMYcCIhIETRFirlL/KNMOqUctIw
UnESokJDW9pZnl4C0t0er3G2xM6PRSP59m3cVHD0WrZMt9ja/qiRDJ+Bdh/BKTr/
cr8y5UsrMHTQC1hZNmdZ+fYn4tjIjtAVH7eVqXmmN4PQuCgZNjNhWNKao8+totnH
4d/aH7qqsSrKOQGTJvNkqST9U8tEpKC2ODZRB+9WH/U0O/UoBc0w13fcQsf9tb0V
Ro/kUtJf14uxO4GTwG7Zto4vkuqNiFzjn/1GsTtdFis7+p1/87zxMsfFFRgjWB0J
EmPcSqVRbe+zHwdy16X5SU2KKUs4O0LU9q4aYmcxCrEqIgX7Uj57Egv+gRY13ZQ+
M+QwkfDGD0/QbNMuKiWV3WaoPKyWoPcTe+NJ85FkDHlvc9k4bq5U/r5wLKhlYJLl
xozrikwPKukskSFhVWUiYZl92Es/8GZ0ryvXJT9+3iLHZp4friBImSIOgkUH7Fk0
tgjlMT//eXm1/JXd29fVyjjPtu0ufDWNGzbxhbD0aTP7ULsQ5i2yqCZxPVEAbjM4
6mJ/zz5Jky5/8nrHB0V11dmpcCVbGwXSYIRnhC0lNkg7eq5uGo8HCbULTq3Yut9I
V7le26p1BkP0INvde1bw654JUvdOHfeuq8NeWSe+pj0LBRNl8qywxGogPgVecbpk
iuxjBcXsEIDLolvJGneQmYlg/Nza2U2Ykvmlo91lL/7atbUrWSKCn3ZC+fKBMmNn
Tp+ANwIpH3ELLI6biYixCvbR0dBNsS8ixpy8aWPSHtDQA1O2tWQpfwA6GaKlUP0T
NfDDd/ZHP6NshQ7386EDcLrS9dq+3tQvWItYU0Y9S8eb5k1pKIlClZbdFWlJ0wI6
v4DmdMq6huKuXSq+X9eRsnSybCR6g+hNWmLVYyVK6TlqQhuWns7buCD0p0JxKY3Y
uPkQh8AKqeuEEhdhUE59cruQmqTLTgr+HHku5lQYZVvnqk4IIiwvy+sfiUCFgOvI
JThgCiXWGPLbvf2mPcdcO3W5NY0jXoX5/cokxPAXSwHzePoWOyJfLKAlFtWQBxCt
Z5APFMdIDnaPrcMwAid46TrLEAogF7dvzTE+JZuE/rS8uxtUCBmQINtIsuwZIp37
m+37nZrF6XV4ozdTEV/U9lThJRaHnyhmMr+hNaBVR9ua0NDxkOBEo45WMj9bcpJH
JYXf0AdJc9N0lLn13B3kl69J1wU1cNkPoMB2DSyowSw+KVkWjB65y50/mFEm00SV
R8K5zZVNIMhcBpdbWsp3vrz0OLVfQ1xnLLJN0VeFCGf4mw74F8kUDN4lfQ2KsGed
nwOey2gxlqYPt9oPJdBf263ALOw8BFFeIGgYlSIqbLRucDNIFC9CwoZzfMOMnzor
17ywGYI9MtZnFP0qJH4Qfijmd7+eqUgOy/ux8pCto04aXMfnRHbWaCv2M3lBHyUm
vFp7uiwb3wHht8xF0ZBDfJ+oIoNDChLexf+04WTfLRmVJ9VZO0Nb9FXJjk/e5SPD
2GP5UsQMpQyOXFXKliRgBUtbmL8sqAl+Vw0bj5l5fzBxIFMG+LMSpmwrobf/EDyL
8339X7SBYIqvEYGcnquRqjiHeSBog1dU7oYDIILmpWdoIvQcbr1Ul0dg3DfeP9Nh
pkZcJjm75BB6qnNtbjtqrIBm0smYTzJR2bAF50fGz3JZGWi/0483kVHiW5u1wjhV
jD5P4EiupMv3NzKZ1OZ9ZzdLTwVuwz+pzFRAY5Vkm2Z7zSTvOUREJHtay0yPZ67p
FfFyJYU+zIPr5jIgJ0ziElDXsiw68Skaq2aaLW37C2O7Pin8JtWslKr38hNt1tGH
cHSJE4KHmu1QovxUW0C2tPrFtLWTyGOLdxgqTeT+6NZx08gYxvi547vCJnfL+kZI
0f7JjhpOQ4XEm+Q5Suh+Fm7FKgrEYrDKqO6UiT1JaW1PHqiD7vANcvz+KF3px7gE
SfLlfVWELqdTfNQ5YcaNH2ktAap+d0MNx7hfyzSWOVFpF/HGY3XkJc8ojD2+wpD5
jiKc7WpaNJU6r/sYAVz0lxEFEPQ/vwfd7UqpmtY/ZIkNfFe1wRFMkNImchby+ZCO
vRRqYJihJwfpvTj3XO1DO8CW99ntfQTYZv9uO0aiUBF2a7N2vWyUdZUhOg4UJAqt
FYGcHVS4F7RfgjV3X8b6+KJfieYT1ApbkrP7FtKBvea0ORqoLwS/y5BtNAAQeO97
hgJgtFzrutpJFpsWXWaW9fsSiA/70yyDNID7fCRz2tvQ42tK6opvjziWIJhv6/nI
R5Q+OZUNlLEtmCTqYQ3R2omD8+5aFRbHSwa+heT5hqYDa+CdJSkBc49+HjzfX4AI
foN8BFhXimqRqCnHj6yvHfutYA6p2geYce/y/Owc6/XGXJA+B6qcQvf5gIPSQxrd
iJ7xA4A+BkOtAPPTU9DZGmwjQEOZ33lCmsy18NB4T4sOHP2H0zF2RWGy0gEk5hYv
E86cvP4pWk1cKJji3yPTPaorDXl3sGkJjHEctBzK2tlMNsl1vVKexsshgb4a0NIE
q/nmGT3h1xrPjVi2pWL9PVSv+lvXWGxhM6dnoIje+kaB2eoZ8h0CeZT6OdDMx3cp
+sVGmv1DZa++LJs2MvnjpWSBAMBgrj6wmuXVx6MpEY3UQJiA9+Ds3JBKK/Psh9tT
mgPY9TlPlOLgFO25be7LjEriTYm++pKSlHWAnmKbNG7AYfLHsBJclnko5HjlHlLg
5WB8yH3yvUJiRPKTfKQafyi9DOvnbZIWLIhOBJ7lGlaieGNG1QenpVBZEUAJ4g/M
2XXjh8NCUM3Mw14yRMbXHRlVJH0je57XaA5/fZX1LejrR3G6yjjQYO4DiK/S8bjC
qHWzs/5CHAXNV4nLsMrMVhSJ8pD8HocPhYXKwEw4VNTiAHtr3zQyAlfZaPShaFN2
k1fR4YLTMF1X4jBcjUge7Q08P4lZxOZN6OJmW8aF2TNScsDybgdxZkQInIQE7wi6
qqjqOdnGV+dhoC1EX6BbG0VAwwxp/FjvsLtGxq+3qgMYrEzVBGkhSdT+9//pnNg1
qXUP6FnMZMZbouWJZbaxTJraOeLcPxM+g82v3xf4rqtaMPT0wz2h8gBcnplbVsXm
VSxlloiS5HeD+67wOagOWVq0dvyZaXzfbh9jbl77Hqwv1t4KCzGPrBK7hkmYzHRx
Kl29U6WFK5e9t8nojqHnPWlJM0FJ2K4/283v0D1ysgN6l3khRa+pcakmiLR+7T5Z
GZSgfNYJrik1r/0AtRpMgparO8ziyQI+yBDRekqKTtM2TB1PGr0MQdv8LBdRuN25
jSU6ezph0/UQYsP3g+y7Sbyh94gzZ5vWOMWltRGtgw9VBS0s3qciR008U+7QR2K9
/o+HTGt3SnYilebnipHDx7eA8Ip2aUptHmYSU7dt3f4ua9PxPJyCWr1A96BEs6/m
FwUX4781P9FOZFvRENcwvOPCuDTksn1UAEzMG3pofSDmUYjgd3SloGb1DMTOKk17
U4L4kSnoflzHeC2H4hoQ2V9/3aB2HAPoH3tyh4tZs79abbWO+RtV2kx6lZr1fNV8
cKuulY+TJ1mDeOzxi22IEpCujN1wH9CuJ4E+enD3VaS/S4lXnLZ3jMO5dna4HS1r
aMEp5EyNLD6GT3cMPV0kipW4/IjmLfl1q+A3zD4eE6BQxs60ME3Yik4fei1EHZJl
DAwXAEoRvfqeHim4MUJcUmGbMYZZn4g4qcpMP/kMbn6k+lwKiM+cYBkxL0C8Mlem
6PQ4lI1XUN5ij9gCtDv2o653esq5ImFAeDMbPcR6ClEc2b0I9x7DzMGZs9XPgqSY
m5Wdwt6CQMJECE1hjDUcBLt7i7Gb2GDpRghbHNtM6W3wdEuSOPdHHPL97bW1eOkl
s5hI32PufN/R8hijYsWP1Cd9Jm3bBj1F9hFjXGOO5j07thKth7kBur/4sPmjqWZf
QSlnG0QI8JznGjDRdcSXtl/m5D0iKVSBD0BKXw4k5kEtI9DkDgq0aPm5//F1Lx7x
y/0O+bq5rvOCs98dnEMrGxIyP5sQ1d4725UsmnXhPXv2q5FU05F9OxGXX1A/+tWf
bBpCZjlbW1FD5XFRRJsCwhHwao7r3F4YRUYUfyB0PesrxMCtTCctRpZ9FyFCruyq
UcjDzCbspl5d1/4F0jNf8ovvOYqpVs7lWJ9464fPMhFbAwI0lwtm6aBaZObKmAwt
e5L7O4SVG2Tj7xGMePf0g49jNh28gohXHuIiXyxY438i+TuJMX4RLH7bmy0ZVe9i
a+M+jB5QAFsa6WtS1Bt6KTJ2OpxZ112gr8ohy6SunvDq/9zDIya04deehuJxJdD9
abAsIgx/fJMof7AW77cA7sQmi6xVgEGrkvCgsV/CSPCRqK1RnAL9ayaSIVMLkWjd
UWpv3ZJKHKEcYTDVAsvo39xqjYbn0//Cd8n7xWMkvKnjNcdIJ/zGUWR7BLYjFxAx
h2ws6dXW5CqOKRWj2w/2RkoIpYtpJCjWwTyCJ71yxvu/3pF5NvZhzJjBk7SCSfDX
nJ/jTGfMVZWqwa5Uic/L1MrzAzfZ0xxuIxNTymsX1x8CBURYdM1k4GBUBJbYM3bL
5Y+Fc1hXc5tVmLQi4P/d5bH8zQoDAoBRFPa0ApCFvsQBQNTfhHbYjnA3iC+ernnT
aUifOZb4ZO7Uh6TZsCEbBcmpaXycWRg9+vCkd5w3SJNgiogoY4ldW3kHsMYXOGVd
tIcSO705zBqL34asleGbppsMgGHJtyzY3Z9BSwqgQ5dG59EdIapzLm/dzePT9kid
f/wQ7LDPT8qPCwGJ+z+3r0stW4GLxyaexMFuJaCPc/Ac/kM/hy/vvtMW20WTum8O
NzR6V/zWBVdIvNMkmUc04modEp2VoWqCpHBxXqblm0N6ol3jmKm5qrAIBdeZ4xQ/
aqdxp6cqmy0nGDsC9mSmu2F21FOQFAtspW6bfD26y9AWdnOzmHP1552IrpmQRkIz
WfVxFrgg54ZgZ5eJeCO+aF0OHrMeMgZCv7a6Nw0FyLG9/nOx7kMg18KoZAHR5LyU
K171hxkUcNN2w0s5oxN2tFjrwrN/EHahLa7zrK2WOj2eYtzaTSZBSVG9bFQ3fJsc
6wjsJa7A8pPHLt1vKJkKypleJisbVhLXOZmPvp2wgee8Sy9/8Vb2kurplAzHJioi
AUCH7NeBYmQPbWVUFouElAWF3WUZhwEBqe98RApq8vp7cfiT802L1RXwtuxSVePE
B36Ejl4Rns9eI4W+T7qKrRwrVsj+ziYAp7MMA7qLk4Y5DETQshOwPcNOo5s1sE1u
16b233OiCRuXU43OXeYxed1A2Z0Kfs6s9WM/J+XyR/jonf6N3RUz5UcsXZZgPXeH
WYLEyEMMxIJ8iFu/BnDnT768Afjk5cnA4jmmGUHXJt59cavLXMzWzekf/3UN9Xd9
4XEVVDHyf1b9L9MP6/Zsu0qG1JSYCrOXmBTyyzdGmAQJH9knW54NoQwCala4aXLC
93fV3fEDcJg3Tw3EfK7wjyer14IFKgq1gYWHUIeenVRluODCq7nPNcso6b8OMY8h
Aq2T05MMV2RLfE7XhE8SW4M3m10s8uWGgVq4Rkt/Fwz0+/yAvvTeqLTWiG7HzCiu
vZejE6R9ZZ8cFVHn+oYD8WH8BtC1y3sp8KxzkdLSk64B5PyZRVS3uDkR1QNO3uG6
UKVccJREmOGuu38TBIiUOxQfFT3HDUwrGwBCVN9PLQdSTD8dqGMo5wXo/7S262Sg
dvGN6smWi/U6QtoHtJ1dQnZ7hhwlN5d83y+2hVRMXhzPZkRR+Q1VI66dth+FcGj/
ytPPIq2HoGugqWEc3yX5kCsbfvxEK+/CXU5eSTT/8yLhCNlARP6n4n+L511tLqmn
NtYU/0qzGCgsX7ePOBsWPxUTNvRJtq1nt93pl1g+TWRhx1FuXivrYspWA0b63+Qu
RRj5RDqNbiIrbUS5+TPej8HaFT5p2hL/XhPnQcVff61Mhrlidu0izkgYB89YkthJ
+wSHbf1cu0x6cuCrFga+sr7Pd7GkKPmQmXgPx+sGrK+3bPOqfOnB4mFygUejdLmQ
oAIUgn8g2G1kM2Lll2YIIirkhqECyFE4L8TbzYdXxT4g8tm3b+K2MRKSkNl6sp3+
75P1uXaQzz6Xp0Tf1JwP6YNkWoIyfVAi/nZc33hj8TUif+D1miiwOeEEu/LkUixp
Smpd2zNET2/s47cz0L2eZbaRbASi9wtjG9+ZRK9dMBr9ZQIeirrFZUaAN4rUnM2R
oJuaSZJDR6YfRVZaMo0UQzICmBQ1ccHvY8IdAd/7Db1CJLh3acg478jZXBXTN816
2cH43UdzHt4bt7swFru52RFnHMQbltvZgUo2FexZ3h+l2Mmy4vpYwGOQauoB0HxY
cKa2I60Kr6BlxIk+dEfpmceICqZ1Xaiw/tp3T+UUgpHZ6gUDXiglfZQasS9ps+9k
lgvbjc38QOv7uIaaqa0vuleeek3Mqd/mjZiesBG3m72SFWP/t6czrCyxRvQfrVSu
/hbn3OftpbTW9FJezhaUulzdbz7YwTbHD5JQephaLfKnXl71pNjeSFZlel3ZrWd9
2gZGkOKcuHI4t2wlsVMpvQohZmfdbvfhAkgpssGcxJDC//iJapuvfeAvXIfXHBBi
zlQORDfLbVK4lax+Fc/2jxhCNXprlTnMxdWPfqn/Umx/+UDhnrmuj7O/v2LtGnMb
O3ojrzTU7q5Z/2L6Ns2bJqa+uidTrJkS6mi5yemxe0yn4FEDcgTkF65Cgao9hR2+
Qadwznm6/LULF4j4g/l31FV0fC6M89gt++FpX+almPmfAa4FxO9s0oLTKsuQdAME
2q4u/DmBP+y3f9RRaOHBcVSrvU88sc94d4e9iybq92jYGQjAM/5O75X9HfZ/o2Yo
ScabQU88xh2jny3pVKjAmH0COrN/71CAzWCx2p81cMlVPhEwvzEWJbpzL+VHI93G
CocUifl6t57yEk+tQxQl6Ei3K/mVEiZUfD+fOe9+SJ95aySK7cEHxJCfpXkiPgQR
PuWfCMybIXEc4t0feZ7T9asdZ+pXgFz7vFUplgAihFGgNQwA1/JdcvYl2dPuzv5V
YOCzjbuXYHyCIJ8JB5DTeA3zrveyE9WZ4Bwqwy76wSdE+1/MLxvdL3ESXqv7oNcY
JWrZpZH9s+613AS/nRikJBv1M6kKTtYi+LScdIvSoYS9AX2WdKUp5hzUJjiX9lG4
9eokiq4FUKyf2da9zRjDyj54FioPJFLPreYNCIjgrfDyTwzQ5Pu3UQH6/negJJLV
aFn7/DwoI8sk/ERTTPNvBrWjUD66o76oyn3pHvb0njVVe3kt7cJ4fDupQi1DD9iF
SWSeWVrmSrh+K2VlRqhIKGasmFHP8XdeAF2wad2nqMC8LN2pOsd8S9XLpIEDcDI2
G2M8cBNajhhD0peQVyjkKjMB7LnZC9Y7DbnWSvDttvGnYL5/XKuMo3zHIGiFEq1E
46ZKTT8y5Q9QrY5w1hlNa14Cflo+tWJ+u59Czby+dpdCGvDGgWeAw3Pgc460VyZK
36f36PywI0rZJZ2aEQx3Brs6f08Ta0xTkiKCU0qXhis8+Px/hWqc9sDgpjrO8dN4
39FXj9thDjF7+pc4a97/IiLPwphqxZBlpaC9wcituVWnUJtJXLprTyjQZM9BvXG9
IoLQX8F2uYkEMk4y1C2TUiDmRJSKxZLjCEKZ7f4N2o4ORJQ+rDon4S/RYwU8JVvp
4JarT6MjIZN8mfa7bBDL7cADPsun5dl8GCZotk1zCU7rCAow0s+hNaSMKAQBn8Q8
s5pAdKhUkfa/RfIQzn4QaHW9oJOcm3OCz8ukSYdQUMUP6WZhXtzw6lyt2n5o5P5s
gAOGkSDPnfvn+va5k+vlwcm16YpKQ2ny2FB/PVj2pDXFWeLS0075vH5W7Dgdywkq
+TzOWec94IR5hnLrX8nOEfBt+NSAl7mnMR7X0BdzAqELGjLawPqjvApAEAbulJmn
evWh86rgs6QSvZDY7QZ9/P/nDqz4c24PciJkHjDKygicet7u3JYDvozUzJuYUtFx
giquOCtx8gKXu5kAIMdPP94xWKn8YmSctc/9Xhv/CnrGqp8RSr8ao/mm5CBERB4Z
8BuIJNW+hc/7kIloUReN/ISsP+Nugce62iO4n7PRuAkyVX1lR70SMYhR8pMvNnI4
7lP0PCWmAHq0LpyFQLN0OK7Jm/SiNm88cu8/hxW0ufVrfRTzsecbVqi5WOL9WvOl
yk48PxvPujRN3tvuBs+7T8Xz4gcJIPIUZZnfyFQZT0eRoEHjxnOGDTjG26xEoH/p
tzOUmm7VniAAwCvvQmHMhUzz4yvUhSaZpGp7hS87X0Yn4CEVDtzpRrlf1ZkLojOg
Ggh3Q6P6dgBNUAdlvxLLDvfa70q9wHao0mQ2yrVTIiOYlFS8mIQe2moaKPvgD+mN
PXATZ2qQY3OX4214sIsrCqwf62lW7Ug3rgyTL+v8wErJcK4cSUjKON8sAqeRPjIP
JIDGpL3zjjOwGNmgSznhmugiC6YfILx1Up8ZJPNikWRLrLIu2wPol3fRentJV3zX
OmXphPXr4AmGqZW3/Y8FVjAe2G812Edg6i/afNtV1zRQ0bHCzZ9gxMTf+IhqW9Jp
9qUtHBeHizl+nhntqd0DoAidvWXpuFeD4niJCRTcvKJD83sB4x9h0HmSgiQuwyDh
1jfXAVIq5Z5hy5ie0VkpGtAzWXnV25u4rncS04rNVF1xkbzV5VyX1DxTt+M7ySSW
m8em9K75XIfGV5gp5vGoCutKvNfDT91lWPxRnmk1QuthdIm8l0aVmJE5oZ1QsLMh
x35iO/zLneGYfweuzQS3D/uqjWRqqSBH/C5BSfiROCwiQhK4xwhDtk7J3i+DyeD+
vugLAsJuZAwUkou8Plg2gJtwPBRb0rajjjRbvYK6z89jlO7R2C849WaxtpaXt/fu
dZTBBNmIDxHJJp3/kXQtJbiNv4CybQqZUnd+2DO396c86ekLfgQL04ifLmicCGYk
G66XQDKOu1ykr2qUMc01G500ZI6SU3DAXbzxlntpqgfuOImGqxBEwwO/OXJyPyrA
8GxgH/afjpj4oEb7BZ3yOqCwC32iFzbPrPnEf+knZTdw6GDmt2Yq+urE2wXu6nIs
GteSmT7On9y24V90plsqGrPtT1+HiN9CMKAaUZRRl7kbV6RoO/vEqGnJLJUg2m4m
abQ2kCqQvucZXTDeRfa9CaQHBDfp7QXxOUSNArXw+CA1TNFOpJgBrgPrrY5kAUP+
JquZwlGu8z+cvW81DVBZucbjA7dqC6tqQc41R/emOFWRm3kJdNKDRzvbjUWTbHeI
Nac/B+l8ZL2s6FmukBdukW9bPWYHJXMN1DAgDqIhxTi6qpxDGtVWweAVLljJj55z
gjCPB7G4WLlHq/2Y2FyO5Dr4lnpEJ8FUdZXj32mK+WcEfl1Ds47VfJYx8148mEXK
XHPMc0xQb1+Mb2MDUDRllWOP3g0u5PZEVJRX51plPQ03vuNIzMRp7VSoRj+Jotit
K99pcvwViR1Jvl4JvIhz/B5Pvrn+Cwu8ffQMXWbIiMw8t0PzyKiQ5GdGSh43aVkZ
9xbgWox/7uvLVzSz/9L9vTujwaaqLnr6xJI3Wlqxr5uBWK9PHTKl2yLx2rUq98ld
NcJNPDQJ7Kb4+CP/HBviGV2kaMWiSCSAPLP3naH52beWKeB+/MpAsJ+3t/46QxVy
Zsg9osrk6Bmv/6+2KUs+NiaYuTPLlq35pHkgbBIImOe92i+b1CCqcjZLeqS3TAHr
8n4eGHCDUXHZQBBNPhxm/VJGoTOWcENY5RPVwarJm2vnh+OeZ1hPSDxeRfIhqi8A
SehkOnsBCUaLE+ktWYuzDAnwcSb8i7cLMUQb4BAjYNB/Z1PUpW2T2T7JeCqFAHIW
Om/UCGJ1mPk/ma39qL6Jku4ft2gr5xMMs3baCXg01Jy8SrmUTpushZz3BDJJ/pIb
ATF3PijZUNsIJ50N1j8thTDO+tboV3hRtjXuWZAna5gpzUqsw1tsIIQ/+Hyg4eTK
+ppbNVJGZvFQAZwN1NrJIcxL2haakvWcTYQcUkj6cOM2jGvS86NvYL5m1hpRPjdL
aaZ7/V/oOa/jMp+1ddFZe1AcOX+Dvv6qi5d7ExnqDgANAe707r3AeRT7MELIY6LP
0shrnhYUgspHOQnf7HKC7Sa1yfFnRKaWskgRUvaCa60Rwkf0LwE1PUWu2Mb/Ocki
1g8rYLuvwahVIqtQeMPh/4YT7HBsvIzCPz6ZFJ72nQYIJDa2sAZZAZYZGQluZmaJ
trZT6r0zCeJgZufQ1ii7a0Yd4hnYSv2E8BAcRSODCmR5VSI5xeqZZ9M2YejGGOVK
h9E57dYsfUu/p+WuTPl5i8ntiOVpQODPh785+ePCxkdaJXYfscLyHZMhYxdAwQGe
LtrYGvCcGJn5DfinEFlnWP54jZdXnavlMcTdXPedop0rS6Sd0bAh9kOLXbZVAGDa
xJXtPkI8vauS/flXJa1l6PXOSLCzv2aclz7Rc4LLX2gWuInghyKBUae82z9kp4or
IQyswJpKS1/PfOuBNnlr7RkBYHnbtVWc8y00I/nokHM=
--pragma protect end_data_block
--pragma protect digest_block
vGZT4ciZkVHn912VvViaiiZAWAY=
--pragma protect end_digest_block
--pragma protect end_protected
