-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
8iTWLVh8wHg8oHGHCRWMVEcLuPiI+/XPuS//MI+DOen31cWatFdGC2wPR8bzIh2Z
nsNwDtK3FSgrr8a5jDPUHog1ibE957UqzsouwrrnJc2UPTBem34oHGjYoS028r54
ycCo9/jtzoYbJILUULytce9j6UVFq4IablRDXDuBpxOug4BexB+/xw==
--pragma protect end_key_block
--pragma protect digest_block
oX9HvWaQOHjsnKPEiP1eaoLsBuE=
--pragma protect end_digest_block
--pragma protect data_block
MB8nQZxGZs8PUUHeVo4JlsjImyUCvKW5mUt9KiiBp6WVpNqjgi+ZTh6vxCKLhq8Z
DzB9rVcTbyPqwpTMc1m2bSIe7wRKWk8vd+8e/VlUcB+pvYB7/ULQn1nlQ7KOTJZX
7mdpFialPK9JCmeGP/FY8G8lqOv8eB4G6LV0ttt7aATu6oAZh9cGV0C2PR+EdJQz
vEiucd8vidalMEbpui6QYZz7yUeg/q5NNZzZfrNNj3sOd56mKoGbEza7KMF1qcFV
tbePrIuSdl9ibMTdyLI7PyfWI5paIJ18n54PLtseN7PHGNgPRDRXcHjBhXEVNXSW
HGE+/4ZgCajTQ7w0sn0XwhQtojNe7OA5W598VJsIsMga0LqRZWzZGFugu5+hRNJT
7fZnilQP8J654kRkxz/n8AOaNOV6WRwVG3vM29N1dko51g6mEdmZYtcKxcdUe5iK
UL0GiOD30O+yG+8/7LKpwCgf3UvIHxSG9prT1loyO1sz5iKTkEOzJDWZiC9URK8x
q+ufQB7oMsg2zcUxfjfxwPuDWb424+ZgSVW4hPtny33PqIlARdulXVSBOribl7wQ
PK3fYqyWMC53YaSOGOQP5BgMOOq5OuTPEFxC5tT9RNI79ut82XfSNgrD2MOzIscj
G6tQyoS1efSE2dyHe7l2ios8F/tTLveqrVQfCzHYC/czTR/+g81GU8tojYPw/em2
w3j30YJsfLVKZ4pA6gRyCJmX6HoJxJEKSxULdNVhnNYvko7gjoj1w6SrvF99Z5dd
VaUbYsEJTjt0GIM8JSD2a1T1t3j9OT6oGfL4G8mZeLR2b0tQWqodfgUmPlssIhni
jfy2CpVHmlK+7zpgTYy38TMJ0aEr4qqRVLCG5QU/GZ68EjVQQSglUS2eCaT6Dvxw
OyG+Db4gs7fwtqlt5YoNd0sVZSBQnue7Oz8kjfQLvrgOq/3zGp8Gx124oH410atx
mCDa0Wr7Ti1zUV8bHPPyDKDWe5IU4kJEW9taOM/ruKkMe2Jms3sPCt+rQ4GJqQwh
Wc+9aG7itgQnNkObMAmT/GuQZ9c4nsfkOv+M2o7ifTms03LNjzPX0yl5YNSgmqBX
STO0do5kNw9YD3D34SKftjzDXubJkrRIzMO4N91s+1Co0dPPKzcKKk7YX8il5C81
e/0QH+eI+Hwqw9iFhqYPAn+30DdqLsLSY08j1bH9/L1gE4nyz963UK3LYQ8ehUAF
bjQvM5cT/jU+Q58Wxjv4b4ySUh/XCDJtzsGQwHY5KBTUVc5Dzq4zbZa6xmTtn2qx
3KIsDJHZUsi7vIPbxkHA2dC24g2yJgwzyfTbHnQbT+vsB3MoR8hXJvoIJbsLiYd6
BWtjA8tziX9UfCon/AyQgI2d0uADwJFdgcvNINkoE8BoK+jOoSN/u+StaLwKcSBc
LtmH69jkOBMH/2MwU5wZnHyUal+NTjHsI2beis0HyqC+VyWM7+rlBmPoi+dJ5BfI
0bdy4VGkc9hiJk0wtRR+1yw5qEUT6Mt7MF2OEUA+zb7b10dgBk9uTMA9eRXdcKe8
r18DQM6idB5hliDB8DDgpJCmssgfIiBaCaluDS41F8YyfD/9cLPkW3o5gIRswUp4
bvjKdicVjvpzG7bviFBD2pjmc69aF67nwbVu2LPS6piB8miCO2DceBBrpx6NrgRY
hw95hyrtldD2K53bfXUJ8AP7ulsrFeepFnocsClvzJd5jbLNRF2blWNLCJ8oDU59
E7RGndhbkkMOIK4i6ztwzkXg9sgyj1KyWzB2pLt5qPhmvzm5KHkorHjdSgTlvS6W
FZ+5bqI88HqnkoSys3Lo0JOw4qYJV3q4bDWw6U+uxXSgYTEKr2f8nECmVKvYTnOL
2O5Ezx0dh7cAHCFCablyrnG2qzlAM7SIoVKSCWw3zrIkjJRvQg33keuRDEs/ETrv
oHdKwvlFvKGzxnkiGnSrhTfGvtaMXF/nRgJV0/BOGSSWdWmUHcQiQp4mCBfBNmzd
UmbqRWNMTBIkJC02JKe/+g0cJMD8WTJzmlbSlpvCh/+7n/pb+9kQ6GfzF01/qEGv
QARJ0EGc04Kg8n415Ct3VBNSK55mE7/0iGF/J93V1aVuSdg4gxXZ7Dpz4yCeVhRa
bW7q7WC4cl2NmulbPXHiE33TaGRkDP/FGeCuoBaK28dT5PjZeNtYf/PouaX7JIB3
JKzHVQAVLbdizBI1bXXrnu8Uo1FIoSD9aWIt5rJbh3iTfx6iZiPBLhtRTOpOKqmn
UX1ez8XOm1wr4zZVKKlTO78CkCmdR44n8jyrouHCtn/8Xvz5zvdeNrPxqjIAZpx/
YNtPNlvynRH7WvnELrWshkD/A3MVw8eyBh10Hw2vV1gGsEF1MEdGwQyprjPc7+De
PumVW9Vh88lYhK8f9uq2QFsGcK5qTsjZKbW55VyIIou0zBGH+VhxJqHdazeRqD3X
pD1Q2wsuLkpuHIHeq45mzAQLf8lfO//WoQsLpnDIhnl/EDN9gpM60Kfz4ORmqYxH
r8ctSXIX0WxLFx6K2Uv1GSuGA3UOsYJeDrtntG+fx9Jkz/7oEPBxeHcC2opNN+5i
OJIZpadJmVGbE+kCI2aKAwWjBbIi/8JsFT5ivCAr0CoBmpzbZX5SWDbtVRV2oJ3L
2YlFNRxEcPwF1OBkG65bE8aPU2qmLTcYoNtZebxTRzF25B8pXWXvpvEZtjAv16/E
e3ZVBVjCmcQi+wsmfWPFwkPiOLw9hnrdmLhgRMnCS+kWFPHO8aULbK1n86+JXDEk
icNPJs6cM5hfhI71A+TXNOvNMUT7Iw6dKElJQ2WYOFw4JHPjX0PRAuFMcJHe+qbf
IDJpEl4sdwsYoR8QIXY8T7PpMVi0Al98iel+AAhX8LY7WtsmmHMeVpU+QbaniHqH
r7YpenOeGEoLZ+Ce/9XvhbOQeBoTU7YGA16Lz/G25oqqRj44N6jjQnna/Ve3+Z0j
Wh+hDmH4D7RiQ58/5Lw2TWxetSyAL6/oI3H5/jrbQN/UZRJqUPS5hW28my8z+ChW
T678VacYnXL+rigDzYsL9aA9v8dUxBiYHr2TpowSqdvXnNtVgDFWiWW6tBcd3bZ6
cTkoxwSJ7rTuqgCwHXFny39SGb3soL9Mq7GaYiNdui9xX/2vgSlsY8kLJJJxerGo
RNTjEEdUeGORsMtJxilZJ8daivXG0qF12yBKJyC59DqhPw3waRg01+lXUCzP17d9
FGdCCeGGcgMmbeJSS+PhvSOXPRbhQ2vAYVGI1zDmfAlK3DOrcFWK/zt17p748CLT
//Ta3EcZ+0zV8KKafkRNLNRZNSdUlxSm6UqdSOGBBOXW8BkknDAeTi6m4c5M/pPv
gAi2mEj317VQ4B4hDQy1wIIYJ3dMqaxHfeMFSCW0Wj3Qsx+qmdmkAyHT+6GK7pGl
tw0uo6f3Ui+l09J2iYkGQqzktYaPj0aTpqbXvX0TGEUZPEDxlPecMGOGsJ3l/tDM
ZGdfJRCyHZqlph/DHY+cM/m1w77P2AdJwEVlrI6UiCHmqvfN/vTaWS3pHCNApIWa
5b2owCsewHpSTbmqAa7gSbFI9Q2blBEatYPixw+Hrc5aKmcbaD3yrhJydNHleKKD
XpkxJnmk5wa2q82se6LlhTBugWySnnoUu9gRYviQWBvMfZkOm312WFbqPdP/sK9u
ujm+CkDOkaf5WSSBFVN1gmzwoOs1KpxUWqpUdnyGlisO27e8/UdLAxCh42UXe7Ws
2DaK1HhdKhyaWINQbbsc/3AWLojZd0AY+r22lmldPLzqhFO+3bHPOVPe/fTT8nsa
+h2G72LsQfH2rDlD+GjYvuGbVhTO7HdcAJ2bBUvdnnawGoW7SSW/9vskxi057FfV
bzV5GzznjNQy1Ppf39K76lQe94j9qIBUXdAieEuQzYvMNx7vb1EDj4BkUYtZ7qfK
KXK2y3/nMR2FD6YBUDFxeF2/QYbnfFutJrlDu5531EBf411nVs2nSbWQ8f01FqRV
IWt18cNZ7tAFebn6TURkDhKrByUC0plyDy5bDF0HLfiO234JebnZtsLb3/A6s6uF
xM1B3EDAJcAerq3rMaE4Kj3xVsucCzILHZEYrpR6AekPjuCCrhLWy5+zv5cpQitL
o5h/p8mEf0LFHYG3RbsXNyuyDczfspVDI7v4g4O016+asv1S8v4Gk8OyLAPn7y8d
vscOqcqX5TXWsrF2t2AaUHobosRBsdSeCv2HbiAxeONQkS2tMoQ63FLYHc/skfaN
LBm0xCmlHSA/ZR0res2zCiwmx3gmTikcBmHY1nmqCXGCDD8ZtNK6+WadIIHZD8WT
bXPADkL/oJvHyRwJg4Ad+87GfrIndD0BE4hmbDYZLFOFu0nEA603moPtn//ACxn7
6WoAPHGU1dnzzLweSkjTIxUDNtmXrdx3Q1IBF3PTY8fJIcpVKqFKaxO2Wn+GQ56s
wT62AM1a9FX0SkX8advaAMZbb2ZYVcc1+7dc3TAXjiYd7BYRhwOxN8gjtiaISnbq
lcvc0wKGa6BlTfmwBguGzt2pOc1HsOX1nMoOp/rkOZuJl7RpoLIwrmvTi9tu3lTs
oxIudJjIHICt3s0VvSb8h8jITDfv78fm2/L1JJqeEnEfkIPhLs1jYREymxMr2sJw
SzN9T91Ce8z4/jPA8CkLXe9S7fgAJR2ZDbSk5VO89grqibajrGUePxfymEfLxpMw
NUnCrCu4Ry4jbTq1Mjm7KP8BtVBq4l35kh/bh6zTlhoBoGcHsRvj8GmyamPdu2gv
izAYw4/U40ZkoHJUPGTisTRKxrGVsI/OaA8+6wd1S5lbIO4VITyKGjvV3UFPg5m3
CdLTNAi2aIv8e0WbDVRJk/aNwMX525dPLYtNAoLxwMELcYTI7Rxs0Ui2bIIe+Pu2
Oo7odBv+u/uUrgYySloHhyOwsxHdx4HQYKO1x3Ep7gcIXLSiTJBiQkD21q/L2IZJ
Zlk51Comvwn0cEaYpZTtKzA5ZMMHPCNy01wLTQwtHRCDGNUR9PUE/cPllcPm1rJ+
SDDCQccgkdee+jpdxBKACAbB1I+Fvlu5U+FMCg+h0h0TMURGARebcI1Dui9vypyY
ht5KhNiuhqbhjir5OvKYLiXcGasBowHQGcLJWiu0w6CQv8gL3csD/4cchCFXxxlU
kASPTmC3fg/Cd6TAtZT6UZlMdYOveSVWkt3/nxjcU8bvPXFWU/9QozxS71W3EziU
gl/OcS1Hz+SIXabdiY+cu7vUFiVidn/8n/yTWEOTznIrYuTf3DPNoAzpCaqvNK6v
e/CAXlK0YllkGCU26R+tpAf046kavTdd9Hmrkadq1Lqqz6KM2GdPiV9vjt7J3qGJ
Vk/RkdRHEoSJ33Evop/lFFNE7Dv7E/TpRtt6/33jZT//Xj7yD+VTDn+gPl2IpG7a
TEE0+eSDXagIDijYiIk9tq8NSxAL2l8Q0DPXVO6kZULOC2kt1WEpacO53c4vD78s
tjnkzrf+TAJGb4U9aQQZZIRVgxNjgHFroGYOTX0NkHS4M2BHKY2d4LbcWY8RxW0Z
i+knq6Z1s8njpVLqABXR+Wt9k+V27WwLbr0q05ZU0NtfRwuZuIXdqlAIVxJscjAw
qG+YmT5C/7h8y7kAjWZQa65wLIgYSuHsrwyvFrsLxBPb5+xdVSwd5wFebSnnCdHS
pApr+ffL9qMKChiB9eMryX9b85hP65r3cmlmSbpcAvR4rXf4d+enQ8v1nadMOgkQ
CA5XW5RFKEQgChc1P3ObgEt1Q09HNv7vyU0WSG6BW3wDR0OAjtAKyYSOPc+mJ1wq
Az9MpgUoKc8nvlkW0z0OU+VGjmZj0mrop9U9rYFEL54tfOkZxgTabWTiilUfux+/
tLj9nxyiMlXildlEb7CvqCs/gX3YWzDOr11yzKepXFNiQwgmvcEeBBC2I0jxcQan
yL78/MU4R1Ats6jz+Syry+EMCrt0qB6HPq2818NgDBTXAD6p/EjwC0JxiTyOGBaX
8zLW8v0h8yY9aMsW6Q4t1sdRr36frZ9J+S5scd5EESulluRddLLzQtMLwJuXz9l5
K4kP9d7uHvep03E/Mkq/M56iWUKkkVkO8Fd1cKLpismhaURJ9R17s8I4qmtNw9LW
k0tQRqXIRtEfAmulPRsHubJZsXRh79PhpQnZXsPmALsQYM9ti1kFjodKtUYbJXhi
5XH0AaWrPLJhATILY5ioDlL+dRg3Z1AE+fJURJg3K5OKGIJH1YZiNpaNL0cNJ2kf
oStrlLmNIgNdfgXFqRD3bc9QejdNn8/NV/qjTPU8s7FNv7QbxX75xL0Kbq+69Hm0
sV7oabvgWJPwhfu+WQG+r2F+duA41QFzj49dbCV2MZ60nOLLH3d93Eh6ronmZ+4a
+FgcGqMVqrwW0KPTVSTf7KjCBy528P5SJbPWXpKe97dXiNzlajVlnpr+vIhLKO9c
rGcnZSE0iOHkFFTf3Cet3eT2rXG+z3qP3Pu82KLLnViQBZ59biCfu2IFcFwTtp3N
AlldAA0xK3K3ItJfMa3iiQxdjH1u2RSAotnQH1OEXAo0yzNW/vOCOH9B1J70AdcN
3/9DDWLmyfLhkDsWEcfhwIegkbQ3AJ9XIfk/FeexbyMMxg6WcNlzYnUwWxpNJrAs
l327UhlRmyqbWByw1VwXaKFUbt1rYSZUyO4pPJfPUy95eWZ85Gq4+Ouiyn0+zwCN
+4WV8Gzhwlos7GE1wn+9TLjAjQwRwNy1++2npYaBODHJBhYOqD1nekyKUXIm1oC5
BKbeE6PhMxfSMbVOEHroCrDRFBR7AsGRh1Fs03lzIdIaaeHuk5S1UjZ8zR5iBLZw
zr565FOTZVG7X2BM0e2zklb0rRd9UWzF6lLiPzPIux1amWHtHinqweu+lRtW3TdA
aneTiukGYKzSagtYh2cn6q9vhtQZSyX80oa4cnTJLeNVn6j6RyvmqAj4qMa4TQ1r
fA6H9WxxxwHHGGoE881vz4/K2t3MZRffzEmpJxgtiyZyUGIIAm3w2sVvflYdB75g
A3sGirHWeRjLyvYulTc95qr0J6njOJ42aicZ7zdxMYS1sHJKtBSA5+nh3YtedT6s
kfgxOKWOrKDroaZvid7zl3fC3Et0CzkfTnbrziJIL/ZQ2qwvOzFDYsoC62s48uJo
bJcWi04Tpm6fJaJffE/uLaGTBIKMau6vHxotMzl2b6ZlY6RbF/UmZOJBhjNDavBD
PFwGTvoPb0rthiSmJN8FK0eTFxARF3uTLH2YzEsTVu5UQGEO1+b+JQJ22E5zIFDc
n3J0AlzmFveHbLj/PbCi5KGvpL0EPBFSLQfCVx73iLbPSff5fyeyawLA+va7xI2O
kgWRUo9d1up/DBL2fnVCGeHQcwVCmlmyUYaCidpOw+S2VUrqy4sP43eEUatmUJvS
bRbtu90mGxDOPfNtF8v29Rpy4F81s7R9aLa/F2+ZhcuzsTvuk3vlCnwdYBHMIeXY
9bR1GlLcYlNN6pMi7tAyiedb9+AIpJk9fpadk3tlN1CiImPqzOp4XIZLy68Gavdd
r6iGaTHgocZIpAyo7r8N8l4+1cbzDDQMQNRu+JRKKVuSuTLZLwe4P8OxWH2Kg59a
KqmfBFFbRkKcA/RO0Y9YDsuMfLWCiquqk5hzT2p6Fu9nn55QoZD0IMf810BxxwXo
4EmfRRVWtXC0joF37/N33RAGLKkOr+BUEVKcu9gGcC1U29CI6YduIVBVWi/euhBp
olsRtHHc4KHrHgCGKmljnQHxwFp1YYJCc8ESB3fyJ3Fd9YATNYERDsgcr1BYhvKj
leDAhLvKWWr+zUph2iMmsWReGTi4THva3FNVj3ECZx8urSGdOh+BG8o/JtZJbyOJ
gkA6d+GGQuCSFlXFDOWU2gXSTpKftuF1WgBGjvKufbxJyitM6LontatdhoabsZCG
fB2vUoPqPCPDW5SX6upMuezjO6vSEt9WESn7fupEqisuPhnOvN/B/0W96QZI+2yD
XGiHZm/ePWTSuaqlFHI/7v/zO80nU45xHTnterdmneCHYnaQA+LB+XxqmACRG7Sy
MXJUkETTdwqH1+IGJy9lzfGXJ9s9vbv+84lVeS97YGRJHt2boyEPs0vAm7LtixMj
yyQXl481L4q+Cuq7L1/7A4qBcYjzvG27+9UKzrrKK2ljea/AuC2DVqXmXJBTSkBR
mfDA83A1J/F7nhxjoGkvW5s/Tf6xh1fVw6apGKm1wBJw1PoJMqjzbwBfDqu38Ov1
qLj+6EIRWonZDWejEX9IO65LZNoZyLG4hD9eHGodEwPadsqSUPL1ZPbJud7Iaa7/
Jp5NV/GyO0Um6jG5/7cVSeEajTnWXl58u9G2G9dh0VUyYrNrpvnI5Cy44CYi7UeH
upKjS78+A7xZgJ+azqR7LCoNOwAa+bbWzyTgzTj9cM/HOzc+Ma1f1eNXYbG3VW4Z
PndavM8NDt9UVB/pW8FIkRct8LVDJ10MuZdzXbzLuDZUrylzDmrmh9EPpjzGbZo7
teqZn+oV7osLMxb1S/Ave10eb7ukg7drD2nwMBwzxQH4v9J3hlxn6oUqLd/paMRq
A9FOnT02rSQ0OWNsUTWeigVWJ7nqnxm7mbgkj9D7gwcXPmBHtClGSi+m0nNupeTy
Mw87wLGNqw8GxWuT7vA2cc14KCK/aw7y8LUiGqSygWBEhDmbJv6FGh4CqbriUdRQ
NbYxheThrk6Pi79Oqm4vVDC2x1Z8ifvJpeOteixR0UyRb92GeAJE2we3VE2SlDXS
Hjh9UeDz7qesGoUixVBmLEuyT6AsHqsxGkajHYxiSC3NyvXJ8TvXQStYRk7NeV7N
ZRD8wkBCjtqRCXkVdQBoXufxCendMWokoAn0WS2+kzO9Xc2RqU6z4VrfMY6W7wOM
eBLMkXpuKxH4UeXrnASz8wIw7N7Cc9OMO44V7JJYi8n5SIPE0iV4kyWkf7iRfg4L
6rlLouW1D1St1ebX/c37lMGBYzYGzwi6jFMbvl7YQPmyYN7s0Fw0Jk4MxRiBTsiB
OxOlGu9gi5BsuBV8k4fp7/KboQplq2n6LickaykCfN+jTVFdnh7G50F5CC7NPa0C
iI4Ng3imRjS+xOEofbg8MpwP+VVa1osCfB+L9OAs4cgE/QtDuxeglcVU+YwAm+p1
JFXSvS199cPRz2TPtFbyojPyraEuINNNS7FOHpaCVlv2RL+1GC8sPtBPuInnri1F
DoiG8oCZtVodff0YGABtNHuzp4Q9Ehj5HQI1RGzIE/rACi1WbYvKlD0YEXionFyg
KGOdJLq3aGom0BEQeThxevXzPoIIaxOP4FtuJMYFQ2gWXuF0fdpHewRaJNscdvOB
Z2Vo7kwgDFqW4SfbvuPQq19kJWOfz/NJC/opUeqDdFTWHqh9WiHv0GBoATjXH0+h
cpQEgLd43lqS1e6NjAIJ+Bjz8gesUEztgbXOAljEa5ck5XyNgq1SGj/LI1D4/zpJ
cnKe2ZNRpOTtRcum3fys+QjXffrZKefdU+ivIguQpclKL9z//IqJMt5rDNmc/bF9
b6a0Uz7bJYd4HhF4T4GZGHV5ZrA8QuLf3MP6hS8L4F8xrazBNI3+OYCUmCuCHpwv
Lx0OD/++1OVSDM4erJdtYeK9r+mEbXgmr26FtW5CleGmEfZspbMqftF10NrMP7XY
JYhItdjDAngJ0EY84nn3Qz0Xy3VbgMpEHrc/UitPAIaZgdHtT1ge3grCmYW7cd+I
RGzyJ2Q2Yb2ke0I7hQ6eA55REZQpluaaGuqpZ9sNONXEnOk9aTIpDdR+SrUx2KTr
C3UMSZpOrimBFJ+O5qna3/cY+E0GSygqKYYs//XVMmZU0y7B7kGHUSV7I4MV0UU0
voPOH4TnXcSUyS7gf485WMfC6fQEVjVfHhVPkzi5WbkK8cMkhXJMIJC5BCqTYEoD
zhWTOx56aGVrQRwto/duEBJEqEyYXq6f8LiZP8Oto5cP0ToxoF8zUWScYcl2PJd1
UVdRE1x6Hs7iVN36IV46c2apgmy23B8i1TkiFopBjo/M3SXhyOiPzNAB9bjb/uj/
ioNjFeoegOcARu5HiAfRvgu10I1oTVOR6RGz39lyhDenZkZT2aKu00Ls8Q/C3akm
Tf2Ym/iZKtxUb0QDB387lOY9mG4K7fqmGqcGQr9NQeFi3mflMLbX65u34pYMf2Zl
ENaVafvADADdFsd759bUj1nKrd3KMbukqH2/Uo9OKWw8s7fNFOWLdRquNopyeERm
yvSuTRIcyDFl7SsHz9g52XoBrGCY0sgDxhXg3wug9i36kdzSfHvw4Zok9MRO5fEY
3Ha2e2yAm2HLn4enMJWM3JmDcMbOceF5yfFL5aya4eIEaGL9wP0UVFSmNHXhL473
QJ5/+DwNhQQKb6vOxZrPVOZxKzi/Eg/UwbyHUty/imeUtZRWBeAoL1irxkwvYwOR
VwFeseSjKWstsDT3TTne5cKTbBFzrC3+RhhdyAEXRgD1p6w5PfDgpV7mpP9fYxTP
cjZeh1R0vqV4iZtIdglttugor90ER/C/YnItI2MunS5PTDW7ZpEFNrrOb4T3R7TK
nFNNLe7PTz9ljGqTyj5przpN0DqXrhu6oL/Ycqi6UDTapI9x/RQnHd/g03g1KBhS
uphdK9wlh8KoHaXxTBtkYeEJ4QlzDJCgmZl7HjW4t3lU75LTxzyBjLosOeSMf4sE
pE8LlyCNdEd9cGYGJIEbewhLsI/Q0zBYwU3XyUR/f02cfEF06Zq/x09oFCe8/g/6
rQqKI0bC0wuGUPuDpj01dV8AKLg43SBAl/CIBhGuTEv91r/Ind8zu9Hzh3mqgdPk
NNfvmWHRDIXRppYLEeFcLPBaUD8q7HOSXbM2zypaqgFS5bR6pH3OXDF5ltd7tD5f
y6LH+ChUj5jWTxbCbbVOSikf+jPwUAkPeHoJddi9ASSGuBjTcrJv6G0hPy0AtTz3
ygPG7+RkTQh9OqJMvWGiy/rnYg4hdSoZuBBZtcXZPggjhJ+6qDWNroKXJJzogwGj
1OKsLsUr+3wdoPbe15191e0zlsp/taXDiuhzy0coLL3kpZFHXQASAF5mdllujq2c
YYrVdPAaTp5NKJiERYMSw+tdX2J0PvVr5V/wUKYsODWUprd2DBwS2irIuHWt1ahQ
m+n3Uqb9XgYbjxD5WNxaOHlyqE25HphzouNUiWXRIu4BY4z51eyIUEMBtIcFaVo0
PAfEgSmioq+hpDEBtUyGFWgz+AEV7TPBstXWmPMxy/xXs4PipA2Es7QPEqZOJM64
0K9Ij9DwBxlCEgB9Ix7XFfjTv6WioXeV7gswNzKbNjCuafDKromNU29bPLADEby4
c8ULQy/JJflA+fTY/xQBMjhu75GFCVYanDaih1wlSx/zHP2vME0rGry3F57c7iej
WzXuG9GCaRyhIvvhk0QwTG1Do+aiqvP0LPtwwLSqy16Rp3u1jkF2H7zIkuDebx1P
pGWgo/dMUE46+zRxJGrWvfiM9rx9U90eBpNFHAW0hQOoM08se/VtmrdM6Knpkby4
BXlsyMfCtlJIlJoPIAyR+/ZWMz5tOLBgbQjBL4AJ10wnNy5Gn7zwaCxiiULtit4K
VO9TnHb8vtrOO1OdSDUMiNJdzBeBkhxnQPEgY8LuDrzKU5FVORmwHaQLuXAfXLBK
JS7sjsKmrYfk3FCkE+L8AYV3GG6EcNf6irmH6nlHb9WK8QTEO/fjk/o/gppZFWXy
hIvZYOnt//odZnsxiWcBUywzF0Cr9vezEGjNTDlhSlfdOmbgELOJTGi0MiltGgJk
93HU8XFvda02KSU2uA6vzb2PMSIzA4KU95L3ix0XsyryxjJyv+I+uP4Z49ElhCXa
Eu0RxM5b0UfWYzYgBhtUDrv6GCKZmAt7FdSI+g4SihxLvzVpERyRMhi1plVnncH1
tzJtpjW1ZcWb8O6s93UgYvQsrHx/kTVymRR8Mgu9KJLKXCKRGm77BYPKU1givR/+
B0ebiMZfH8e+vr0hwGWU1VRHE6KE0rCJdhhUQQ+cBeSSWBLWXurcRi1k/695JDNb
HirxUTyc6tqE3NcsKV6Ew2RWMooly37a605uO96SpTqnHdbl3iSKZDv2C5XzV7of
v8z5x8lGoQHUr8LrwNxGq1o5wfdb0EeGTQCZeRDDxo8RJXcqDuEwwCk7+q7Od5fU
LJZrBu/HIERro/tV53SdbBySQPFjiuzZvJAXpovZ5Lo4OEQb/gu3d5uTrgj305Is
nsISghj3QtQ0dLp5XS+wwY7ACITXmTu1O8JmLamcGe52D20/jQIS0PbFGvt0C+Eg
5BEnR+5Ra0YV4Sw5LNnKDMZk1C2HDh+MxxNbECGf78nmvXPZ1GPkmxGnQM0Z9adp
U+rpnBJ4u3EnmVaxa7wErM9TDxwbdwKWjmvAoMPp6LTLl7y+WxarY/vTe0ViWEEe
9zio1aUFsV0EPb0nmhy+4Wj/TpK02MqVZmWCguc0nIM27NlzGFe1XLYLItSqtrW6
Tu2crlqXYpH842OdAIR1EUJvp4l6GmGFzRtoL3yt1ds36nglLC0p9ZGN2f/Ab17M
nhZfyqtJrAkW4HQHvaDd9c1d4UHncBBn45qJ7xHaNg9ciigKJe0ZN/2Ky+O2jtbK
1iAc+lFCM9Hf1YRUW4MJ/R10+USFKFvrH6FgGY3Qs/TdmYk9X1/Ibf1ckYMxD2uE
P4c6u3tGp7wbptiwJMYl1/o213rEuKvBxkkquSOCKWRlrI5pDP63nr3vs3dXM9Is
8oDtsmTrfR4D+qCERINse8K7aKTVet71UKvoOmtNxLuaTUw5ABpG02nA4nntnzye
3ID7HWV82or7rRliYpuj3kt8NmLGlS1JSx+A1IULMSfHJrc55BcqsJDGVpUdaybI
zshCQ54oCOFv1g46ukHFO6wNkv5TZgLvMuOUOQEk3F0vmIsNrEiWODhQZtxHUraU
ZNlSARW5dKsqA0Y6iYrZtwgch0NP+nDHKADhpz8rghDNkFaL2T5kdIz8a+RuNpOh
yXviKnyPPlJS2XaNGarHyVqR1Id+jqbY6WIdu38EeePWZrxXYR0RnKm5GVSghhkU
K7BbYzpCRVyqq8RadsPNQ5cMUAVK6yncCKHWDk9X5QbAPNe0rcFu5xuGE1d5CL1k
lm+LRFF9SCxqtsFa/Ey087aU8fKuZv1VXbu0vo0Fbh/7ntTtn3MJBb7fw1om4mkk
uBni7bHwBg1G+FMEAkpP1jBWIEboRiTTfLUjvE/CgcHIGeq6vXZoTcQjZMk+2flT
/ZhT7B0yUvBNgSH5T8fM7mIZf4/gEYD+wXChuhyXXFRdp1UXy+WRiTqKsRjS3dEg
zcx6cqFNQL787m8PloFgFaiUjiIt3EHBfG/N/qiqnyTdL5U18ksOPxKDB7wG/b4+
nhKOk8dwZwKKNsrrRdZHbqV9pmEmH6DEb9fm/hS36pm4BTw8nFT4VBvOQhBMzIrO
iJ1kcgvOpmdOywrTfd3BAQg8F8VboKjebyURM6av13f9cSrhW9WqT0lY5zUxSShZ
YkY1pNUH/VNH3waZdfXd4bS+4QzrdrBISX64/E0kouRlQMcQCkVkjah9MCQRjXm/
TAs8NICnRyOAa8mUTq+y1K5lmA2k0BjzXxe9xMy86Dt0tw4cz6UWm0apYQjZgwex
qaTOkSXk6SjmSJZ8RnlmRCOUCJQeB3Vef+cASOq23c9eOWH6aVwhwOcx8qbIphf1
DJQFKRDIlEZBH1UIQ98uphClZeJU9YMC1oSNHHIt36Pab3/V91Ya+Hgqyz1ySKc4
aNo5oELskkvEABZvDbPSTaQ+myBsSLlsVT47dRfvdtxNoBWz+hYMo4410OfDFKOs
KTGlOFPCK7Dd1PwXFMOchS75inP6Oz/+5fS9gD0uN1nMzX4jqDqr9vZ9Fg3Me7qR
aQzghX0b8lBl+rLM19KDM6FehuRg3Fi5THyOAjIa1e0YQHpKZFts+6BOshm46dxB
BxVYKlD3FTYWyK+ubZZCE5uIRQxLSy1yhSNuboL+zSAvG24xdHgINqDEWThEIYVR
1fOwHiNE7mrqv/FONz4vw1YhWBbDk95YrvbkSskUam5InlOrqHQaG2jV5tT2mhgQ
ySNS4omCQYI8Hl9uM8XHiW9xcPLl9ow8JU9IYqN9ogVmRrWSqjfFBmOME9axG9F6
rfpe2LKmKXiTiHkfhV+Dt+cu68DKo5oVFcJL4H9IGgk2RPa0oSW4i1rO5h1WhVdm
lUO6zeoKCQKRWxuVl7RD9N6ZjDvAZu8n4KRWwAK9iERw8+Fda/MYXNQFivBJrlUp
R8lU2/fPtSgna2BRETH1GpLaTBcrypTGWq+Hj2bUxqo1GHfXvknazNSVjbVVp1Jf
lEZeyKCYdSpXU3qSm/79ks23C7xRpvp5OyMxREpDmCkpSi44G/omOIrJtq0Zzcpx
EPf3RT8trVROM/p0BCYbS8ERAGZ0U3lTWwY96Gb3ngXeSDEAnf0X7I6PD/Aat6Dk
u8D7srPzgaVnKYLvuHY1nSwBcbNb+4HFRNI7S82ArgdYuXsOzLbvuFq49lpDMMTt
Q9AULywUSPniwt1HdxYrqdZa+fQkGSbylojBkxbCUvFlOUrWqj2L8T/EHKkzqfB5
UWr6rqSUswtzF1ZnxuUTbANYfdmbvVhaEZ+n1YBkrV4qd47YYXdrz3iB1N8wfum+
pUGX+gs1cm99Y6L/xB2GDlB6cHNCmkP+cKgJ6G+ZKmWWrMUfIIhg1YCoRLY/xJ8e
iHgatnz12HxRRXk1FKaXamsmiqEyzb1qlJPCGfITz3fQ4BF+76Wtso9kJkdfWs92
elD0X6GiogvntOeuGiFlyM7KYqqrDRMyZZQa8THVXAw9KMjbD/TtmziZgku8+ZM6
xwUgVxWBVuBzOj6Tgk43++VAZf7TTbONeGqZ3Nnd5APqDNZE9wyboykZYftMoWsB
Dl6EDvZcitf9ovq8Q5kU4hrVnqc509MN2K9t3Z4MKnJGfVnEja9lF5XQy0BQVPTP
w9YG/IPVOdBsXraFB+NzhW0Dq96RsU8LnGwfA6kMV5Y0wp8YxVeDvJVUTHVN772L
BO2q4EVtiNar6iZbfgAH+1K9Xp2B4B0dbpMNsz9X8+IZDafxzuxeAsia1xgX3w0Q
J8ADVtWhIYed+fLHsw7yxaD8b+jD1wFHXEktuK04QTC6kOJEkSzY7I/CxIKQZCqy
GVwX0ctZXRWLK8BmAUO095T9wfC0I+SGnSd91MRY85wACIJiLmfe4xC+g0HftnnA
Ik+sTfgUQOO3ZRsUTi10Tqe/XaRwa3WIiz8FoKOTrCAoeTCEiIiXM5cMCZTl0Q0k
mTwwH8jsisVNpdgWd6KEbQguYAt2hVLmJrcI0LFQJXhsMLvpSm+3lFdIYJmr0Ikt
/eFcr6NqYpeO1zIsifIeFVkKooriH2Y6pj1awsn0QTq2Jwu6oTpla08nnfz1QUBy
Og4OKMJ5Vv4/xHcr4v1RBeBNLVGBuYQgmmMg36clotMa8S2YZABPVmtD4S2/qOxf
XL2GrqDR5LvWR/+ag7B1Z+5x/9WrNjJd0wgW3VFc1zkHMmRS9srfncK8r2EmSqVb
ugCbnKsJVDs/EflZgnKazgN4DeEHCVo3ehPylsJNKdA1OKF4+JYiucF1+BZLyuAQ
PFh+VTZ26zOZ/3syphTtEGmhnQHr5rK7V7Kx/zlIqAcyjsS7ZAkyiWvSR7VzZUSI
6qi2abCXX2l5suM5muqleFc7Oq0C2RZCMTpqsE8IoQyK539lu5fe2yLERP+/BQWE
+QKcByWNjJ8ACBIbR8hw9NrHIz9cZTVW8TFsrs+GAem5kjvWQAqDOKoAPzNqhetA
fVKPNA4Fp6mAoA+qeQw5DG4ZrQ2HZHyeOBsE3AFJKfP6vSLlvJe/vslJAoFgbhce
CrRy+WYpnrn2xW4FChNE63icfy7UWRDrEokzDF7RiSBZqp3BX9dfs5aorZLctvVK
pOAt27CT4k3h6YszEttea2wvfDKhGniLkb1H0ErITks6HHcEN5o/zc4JBVfZFILZ
nw10mCb1/pamHOD9HKFbDZ4cmhyn5KzewR2n8FPIPBDn1Bg/Qm/LuHFFUmyBdfhY
0MUW410IcXMc0NHBI53w/PBq46KdrlrTyawJ8MkcIv43u3D+83d8lYS+s1aHBpKH
xILxxxpvZuGKVSQs76IbSaElVwsdb1mEHXAoE3EZ09kgTyx9PsfFMJtT1//+kKTK
D/wewCOhEBroEzSsvc/fWNAnrfqcvdxR829RovitveKWyo4JbQZYAcp7pEqc0sN+
W7qTaykU4sSR1E+xoJRLFQ0Ok+rFnQN04PmdtwmUjMCIhD4WdD7v/KdYTrc1psBQ
+xOUNcYuA0+kOYy95Cj6x18Ht3CaAd0pQSVsJJi5qQimgk2dfOBz06QlSdDmi7V6
aGadMUiueFsyPXhtfz24Pw1tPWgWg4ZCMV6+GT68nn9hCjZHmkpplRRW0rLC4x4h
KO2vN8k8owgSo3TAZ2WsbhIM9HbJK5VaRV4+DFa/hNLsNhyoJt24dR+TqlDcsyw+
5VbqIkAGvfxmJwMRg2RuDovNVjG1E5PFO3AHxof0B6b7q3OdGegoaU2+8CvupibT
mMgZaWsz3LZUxz1f5bJn4Syh6kvDEBv7kyvkLx3B0t5b3NbFDDzUGHGq2BfYAnRL
+v2CXa33z84YRLwYnFJu4/iOfQNIhisiIQ+nvqI8W7p7GL/IVW7zTyshAHADTjOs
Jqt9AZ5wmsrCOuLnNBBz4rzHrz+tTyCND8z+d0kTzBeOVS0bqZspBqFNJ9oPqJA1
d5t3+Zf2Y7Axowf8qwoYVTyTcsPIoziR9nwaPQq4Gk7p2vAAP7ZUCayo1+T1TppX
g+wNXBFWWdYl2/ALKOeRpYrzE1eul6lmzxkKBHFlFz+0VNeFbPOdk3237ZXZPPej
TVqzzFhr9F3ERHm5m8+bFSS/o7+BM8xmVujmALZhPRKd8yRUsdiHR7EGg863f1j0
WqiqG6UotRxOhOZw7WHNu3pADfy2tIOSlA8GwvMaw323kRRgp1gluqA2JMmKLgv5
2nELfuSQ9lubXybrgvKCCQiDht/K9K7q90U5CZcZ8/LRXe0fpZLozUZgH8rx2Cma
6MTmmCDcJHE5GvcQRy+EmOqbvCxRfGjeRQSGkn4jyrVqQECke+jLU3e6uuGcoQg8
AMyzgUehoXGYl7bCIpBFnhqZsHxT987xyuyCEg21pUDdZMcPaNxOfuqqfXTX3Mjy
BnX3D7/yKZ0QYrM+DJNekpcPzOG9PnsN6nZ58imnIQ2OvYPCz4goMrR9t8YB4DTP
Hq3+TaSvjvN4rW9qATlfJkQHPYj6jEaH8Y6kMiKG1YAk6CcbvHyFD63O4v5QHLE7
FebThbAN8XZUsVJ9LjGxv6e4u6k66UVzYURKe4SuEswVtciFXbEZY1aSPeV5ZCOp
9wccM5YW4xDZdCbjIOZQyurCHH6HFdiqmp8gIf3m+FlLMOUYoMrsykreilJeGAHv
xMakW9koPSUjzPwuyHjJmYorL3xRo8SeDnevhG1MLpwJ7hY1AnKmGEXW9c9yXQX6
UE30/jneKnh7gzLFKJaoB07c9kEOVWuCw8MDxSyUjkOLIDgIQehkAkLTgujVCga+
RjqLZ1h5hELHZqxiKvzl1GP3bpkgEcBwahoUgig2CGn80Gg5moKnk4GijNy33wzK
R6ATqsD+KJKXoYsOhEkJSSthcXxcCGgq1SAc0aGi5dVbWUYUm4+C+5hRI0upKfdz
JSJ0dVVWRGBjwFgWDWLQ4PRr02+a+VO3e9LNnkHXuZppnbheMzQTf9a4WryCd6CU
n1z6NeHesK7SWFEaZVKqdEklAUe4qygC77h2vE1qINZ8/ESAYkCcH2Jgit1VfvQw
NfaMzL3LcMWbvoUQMLRS/JsgPoghG0UJD50fDCcvy/1kT8awSWgG3Klp7r7+PXn0
tK1EbOmMohEg+G/9KxhKM/GY42xilRXz/VlEfYh0DNYposkjk3kGlsk/j9gSf0kH
mTGxRRwiLeQ/H+t7lrsUkxTeRDvZLwZy3hz/6SWUOK/FrGRUEd0qMdRTu/4PcO4s
MOkoFVDShS8JFfc6JG+eGFo5h7PLlbTib4yo/sf88qCwSGn5vvVJ5cvc+F5PQgHU
oPySkh/VmwEcuc9PyJx2Kv9qScwonAyA6ZsPBYMm0TvsWM/Jt+5WkFTShNzxqc5M
lSlL6KQBZJUWCkKtZ7UqmEjKlHT47IwrwtL4oKHccGG8tLIOhTYfOIB2cQIhoAeb
nJ45pvHFSBruedQUqPPsO6GqEY5JZ/8aaTFz3msXmVnc8vB0PCtyHkMwd/TLIHfW
ikPyRNjosh7UzOR3CsS0BMEPKqXXNba+PdY1i0flaUa4EpGsP0eguZY6aBXDLWA/
riyg7nnXCiJ6e9kP6LnHV5oVwRik1nbHHEsgpc3P3Pi668B0tuSb1gUZMfdPD1go
mGnkWNcdrP9EpDpiz3tW3viDIwGLMdQKiTi6pIHdzI9rAYpVB9T7uhyEvEAy3IPz
Ctkq62Ku30suG5Ff84YvDup0vQYP1zHIXXUPPFG6eUZ1ldK4hFISjOW1rNDW667f
MaTwlyLLwgtEbi36+1eeU/QNcqqgL+om0lKILCJId9XYDfnoGXryMmAfI+Z9GAKR
npWdDlkfNBay8uZzdGlHQB6Urj11HPl6o08yCGAipomJSCxZaiVwX5+t2mrWJaSX
3PIGT74EWZmTnLWZxJUwPFwRXNC0xgtA+lIJ8xebR5AWt3KV9oN9OzD0SGtRahZr
qnALSSU6vtN/oIQ8kH+hHJ7bS2Qhn1T6yBmNWNHhhjyjVU2yV5YFjsLwUMBidd5j
3qp4gj4g/KWu6ZF8+iOkCUoK+XxKC80kxhC2uwhzAvjqOQKjGCazCB+j2ZoXP/zN
3w8yjgGIk9c5muMchlt7MmPTwaU1Xz6Vb4M3Mk+0Yb4FE/wK62BluqtNmBg3339y
ybROKVXGCUrZuY0CCnbcJ0GOomR/YkWxwZv7NtgjI6xMte7OgrPu7UAnjyozsreS
tj4xHZSaBeDtFeOTanaZIuZcaM81uUogu6Xx8vwi21g3FNdFFEx2DEy6pfhaGNiq
Vr+87bmF9jrp+kAJ02FV/aTnvPGQ+abohcfVTsaPXK6R1zCzAGv6YfJL5Tvp0MXn
VjsB+fRQYH8Q0bpF5G4TntS56PG8zXlx2v1DDkAtMWWpRF/y1k/lIp26lkvvkIfE
P7wi1fcsCTjY4xqE9864Qti4RaDbVa2V3AAh0PC5IW6FeB+KNRnPyQd62qMqnaDU
tlSBjLXgLoss5BSGTeyed9jKyrpoCIkPtI6jOp6T4wlbKniE3uSjHRSQAGF+ZWoO
/joHnP703N1EeaZh7d13jtXvqVVx5Zg80cdNUokF7JcTcP3nMsaAw1icE3fLg/F8
K07NgpsLndEEUkIR3jvzstl6Vju/yBREcP7eoreYqa3xcSYQoN0rK1Lw35H/ld2V
8W5JxK4qwEDUsxEPso3i/E2V0Ej+1DjJm5SCA0ae2DfRYUIoyU8zhgPuYuVjF1XE
0ikmiQTL4Hj3/pENvdy4+TZR3/4NLncnsC08wPP7wOgPtNFYhEwXO5WB7O3KYfmi
5SsGF5mn7ys33gyx2DtM4ZUOpFgEvrSRN5YdqIbMlzmGPULbc4hdexaCKI4ezJd7
ujleONH8ZOCZisySi38D13olPKrW995c368ug2zg5SpY1+DlazatPAl4BhxG1mi6
UlNEaDGCnBGetFbfi0Ezniz/uj2N+P5t6uCyhz1ix+0Lm5gwO0ry0pZwWyenBSKp
V8xIV3ybwXglpS6w6c5sgvAcjkCIkzHLxHbsEw1rByVMU7o5xWoeLLjKIemM6bbt
W93SsvKDUsFOuogifGJL6+tXJoAIwBcWKcHqPg+SLP6v4N+7UNAPnuWWNXN18HlJ
8QxjM6qrZ+tJ0pr/3iQTZ19G75Dg0dALvoH6QgdKJbbOCi8QSMFw8zsV6vhIsee5
leEfV4CIFwYtMJeUSHmEKnRTS1Ipr7wW0UXNHLOPVVYMKLrx+ekPCRGG2M2B229z
gcsA4SVyz+uQZfre9+2BNMX5B1hLHRAiMlzTmEIIKZg3WF5D8kJuuin5GmKLTFGL
L/p+BpdfQ99YBahQ8E1+i7pEc21+kLd8EVM0D4XE78bdr20PSDzWqX6QJWUwftzg
Yu7iwob3pKW0i0wqQJInZZiCGhB7Dswfg6GS+XwWYxpI7lwk9pojirzDki8Ju9oP
DrMWVVqXBYYP/hJmViH1tGTcHy3Dbmnd9lV/ne40OZ6SCEHUR5D32zL7wCXrho6B
BjRLQclE2ubd+tTr8gCS80CZ8Nt+xEM1zbPEsK5swL7i9wHZJVBjt1VgdAaolHj1
gvtjQiy1yGCtn+i+VeffiPs9vKR1uSZg7YICcRUl6yfyjGlOoA1K/R9TTkDlB9j2
vLeNqWqE2nxzy1L/3R9Rh5SbIDlYqyKGSte/5VXemuEaY6Sk6NMXdlBm9yZOOq6F
XYbE6w8jt4AcdCWt2jPtRjOH88/9wJ0i80wmrWJ4CAGfhdVRSpm9lphXYcNB/flr
dkIL5yxhNtQbtmpHC/1MjoLE92HL1n5cjxwc2Gkt0BbUstUlcbQEK7CnhGXV8juH
YjbGWhKdKPkY4FenfDQ6uQs5JFPhPv+ICQ6pQB3tEJrutH+J2NxXl0myk2e/yL7Q
wWpVQugR9T20PLVGYEn9aHvCtnXoYrJFta2xvHgq9Ra2cwh88/rPRjwwHbLg/jeb
Oh2jGBoLmmgMUl8BwSf6XNte/oIW2bIiSe1MeeavKo5NcGK9qdTbyEIwDx46UOB/
4oHfP7ZkTQRM0VKJsDjdFBH/yKXqoW9Aj8aBffEjI2nIxXNS0tKga6lO1C86Mwfa
c7+VTSLQE7qIfh7m8/+jVrgsLxwnXYYvWkqabIxeykqeZSGBaAqJhMorcEv5/DHO
wLQKiS6kw6jkjhhxWewPeSEp5vhHLHWaxKYXqxzYRQ10ORDX9ymtmLrhpCnrV+I0
rlzPaGzPXO14fdgkE7gmRQbjCMbjN3R4dbV1AVYhKvSu9MKRtLkTRMpV5rK1RYCn
Elx2mjkNF1uvae1Z43LNSF6vMoP2vuj6OR9XwJCA/30lhrYAwr//RZ52cC+3nO/g
deuibWb7GBcs8vaz2geqG2k39jCaz0r+XbSUxIg7ntXumq2lq3O6JnMiEj2ueqAT
xB0cCfwAlL+GBW4zgyyEp2kevQH5Emhyldc5UwkBsm6AXC2R9xfH8R8/M5cavDs+
LvfEsZz+/9S9a4y5b9DrBKBnn6tnzkR12FGcpaHbclEK7myexTpENvDoOD7qUD52
fxr7xzxNA6bXIZfs9DQ7weV18TqEBy4TRyvE4QvIWkF4FwPwO5REEqESoh273+Ou
3ZQzw58OHsGP0yDK9dCw0r1FeU0GuEUkmDwXyd0sR94J910TZDau6LNliHsU39C3
dQIrcVJ+jxB8tiUmAysdUR01ZfTOrsJ6FYnvPVIwhKoqOavMXFEexGJhZOwr/YMx
IhPGoGiYNFL4xgzwBmbdtDHgNd7jCJEWfkpn4f0pjfaEOPV+K5BH1GYGYsE9fl4X
C1/O0ul2mHck7ZqGk/11zvSHd/ywT1wbz/zMKKrUpqhT6iFDAVXd/K52KRHOExJF
8RYxqe/4Mvlc6kdMssaSG6RKLsIjy8U36xyfIK9v7oep5mEoI807hSniT5cHbJws
JybrQXhuMcwHDhR7kxBcpHiv+zQgtombeKGqyrEY/mnMKFhi6MT7wrhu48Gu0lxh
efVrYoXdGnm6RMpcsp/fNFkuzlh2FYzIRb8+908ZaHtlVdYnzBBAVIv5ouVr8aPu
ucNtPLx/nYuXEWHKpNgtiMG3vUyzBE+iJWmRXDyvntZd7bWcQlidmKgu4V2fRG3j
pzfL0Rv4ET8/D277JjTZGpHXXBNQOEjph8cMGQdUeEBoNL3twCqMgA2MH78m0C5u
ndqyk92uNLtkLNwgw+AUNem+afTlKXvRAm/KKo+18grzi/gt5zJJzndTgoFZ00I7
akum2shZ6mDPOXDykorWCcRd/zZVv1YtZQscnI+Qa0DP5xekNVMv8umVsTwKmrl+
llIHM6G4CFAQatkQs5Cbis2fxaPd7VMwSqPVVBTi3xL4if8ZSmEnA5g812QlvFzo
x+k6yKEKbZBuAFmwRD1cD1+KYUZxjGw5yXRdFTnY9GRmK3FkduLjGX6N63t2vXHn
0K/aor/vzqFZZhm5KedyvCtGDkCmhHhrgNDr1TlN5j2lgBdSjSnMFZyNzlNLalkj
Luw2GZ4v8NItPTMb12+rW7tbgx+U0vgPcoEF3d9yOpYGD9Y3v3FgvQkSypB8yPbM
0cDq42yLt2QlRhS8I+JcXJzFkoiZPSdaYLtIl2Vqe/1eC0GCwzqeHudBftE58e7d
cANaIlnH5HFc1MWh7odZ6RTplzwKGsh7PD+qV//aOgfLSEvEHY8E/dsDBegWURC0
VnTkahI5JM2NDzPAUdHDybYTGcMKwd7CclYXKfGIjffF+4dzqJE+A++tOznPeHjL
8WG3vbS7xIy588WnAhi2Dr2kTR1hoL685vElbGxcJYi8zYEnDoY/vP8ktTc3o79Y
x9xcr59JHFTvmQQN/ww9/x8iTCgM7ss6IcHAfvm2pZpiCGJWD7a6nORDimr8fCBr
SngJ33r+0r5Zq/07S3sqjZNcQGK4Hd218cQbqvMPhilrnSPJkOZxLgQL3T1GVDra
K7ZsB5lNjYRlEuBwpyzpN4x92GCEu8Wl2D3V10xueYAE+5bVelhxdbKxinkf0XHK
SowE8xLFIXvdv4/NLtcsueX2/YYex+4t25g5wDiW7bMZQPeNhqiexiLa22i/wOVD
uLvnkEe/hMp0qj+/O+ZiPsUjm3CMVrjfJijsDE/mUgom8lLIdr5sJ2+rYD1k64M8
4VIZjkxRqK92UgUMylz4Zz6PFCTkNwaSemqJnlhkWbn3t+1mNre03Emvj+A0UKqG
UiH3K0F0oAiXcyQAP2NSSlUbVQnL2jAC73KJciuaJXQctO1QiKwfUJWCs3v96bl+
DLZ5jyDc5EcCCjbBunTy1gx6Cbd9llEM2KfkhPXOpXsbJ8csdGXm9n7rfUiRUsoY
zzupirqyV+tUGEk+fDnfZ7gjfFvYmp5e5fgZx2H/B7fae+241YhYcHXDlIwzmjL8
Izmu8yMBbS5yMHEUdFffLW2KF9tbFlkZXaYunVYF+Hbxo29ttEkRFhdTDMxocJhI
zW6y1IrxSfFXPrikjEhYK162AHJWnu238rwSEXeJdHTDuRQEWb+PctsXhSpRCKFd
yxfW10kovvqvEMFeU4zqATsDOT4yxKorG5hcxblHUk37nGGSFmTRmxbAEtSLCe5w
kpQC6WUPhTbMLw7R588p8cB3CPEn6qif87CDn3p+sT6gsZqwbseMX8FVKEJl2SIS
dYdwgOlluwqFs/dLwVt6xx77JRTy0HVCbGNjHsOrfG35rMP8A2vARSmL8+9Xkql7
Jo/UY6FJV9WqDRphn34v50M1rDYZvN/Vgnk68hgCXhE4kHi6SjzPVhVzycZOu9xM
YbRFjl13Ipgb1WNJSf9R3eWGvUofOGwMAkcWHdKaLPXRgojInukuE/ljg3pdrr9E
Gzdy6kSkPWWarXUjhQMK0cTV07A+DIvzzi9ntm1J5RdT8TwlGNEZ4uZo6Eo24CUZ
enXG+RIGHFMPJ3zRMzNcgevIuuGvTmaKS0UZ3BAEAZg3puBmgsE/QQ22zH4FuqR/
nKJgBZcadYZL3qXH3W+3IzbOr84617hDHkvKNwJnEM5AAzVZKSGrxlW/0o59YdVx
vosJm4OO4oYEQius3BVHhK/iUlm1L4CO9fUckmLgusfh2wOLkSsA9FFjJi8N+/le
7rUPJMI06yoIOfEgifP0QMJ+p/8o1Qy6D8ief9mcyOeIYkJ59WI6OFi8jSGAjOGw
ClxuUJb24dEyaWWV4J9I68XErDbel9uq3ol9AIw+DydIBvmO8lN8+rmAhKuc2OVk
4ZGh+Ls9btHrlHtDU9e73JLmDjHu50uyQEKWgzXUxsgwmmtSg9xxIsvHeRZ0olrg
j7rHG3N60pc9jL5dIdPYv/LX9wfhdkRKqw2DOk0HF/SmotcJ5nMu2JRRAvkW0mwh
tZKfC36aHEKdw+tIRGDqDUnakb4iO20zjxooFXbO+T0qMKLRfDjzgHMxjqQXLgNC
VCjXUj6ot9r8v34EsILxsIFO4idVFGLh2S90nV62xY5sU7BbRhIYa5LXX+fozEwz
ZV91nMNF86FQ6UVEvNyH0rCVDBgDdKzmXBADbzi587dWxMtGV4CzhbtqvJdXQvZ0
+QgSFSrc/zWH4nNii+NPQmV9xwaUCxdoUtiDJgRnVugdsJVJ2/fYt94fXdzsREk7
9seNjLEsAN7UBQ80v428Cal/HIL0ySNmagK5ZSMVN4QqacyEgdvUb6No2+XJsOLS
U9a1V/LKKTd21VvYEO3cvccqhSRWrTL1lPeP/PyzwfvxfNfuXfFGIjCI7mz1k7Mv
dshzuYC1HIW0yKeCSC7gzMJTjtgh9wvmY3S3Ab/Dam1a8gSNll7PURGaVdoBwDSQ
JLcZ46RAa30sO65wtITK300hruyqbqWvGx4vimfypFXHqW4PfYZHBAUSIB9V32oQ
QmVK71Czn1IpG0KQJDOfS5FtE4u3IofHmR8KO//Q1UDz/Bwd+uVuJ0jhFc0Nlwon
d+A3VeNXBgu8Vlgk85k9/Ms6a7B1rD2iLKJ8ICS4AmdLcP41k2SKnp/AcxgVsxp6
gMjQGIVeAF4d+k0xIa16jdVSTem4IjDbWJUxKTXIqHG4Y6EXsUpC+2d57pabw08J
Jl0qFr2EYtLVqSUqLUvbg8PWTOTpqecP5ZZ5FCj7jH7UbWQG5nxMd1azMs5CwAQz
cZkxW1DWN++TX5k1PA/YgxEetH9YPkvsl+VP6wlQG5kmZdBMPLLXFjz4WW5z88TF
d+14lJbiW4cZQaq2pwWKEonKn9nGlKOt/BpT1Fv6ZzmYbOr13TazvSK1FyOmJWWP
Ylkpv336QdxlbKKfJ+BoK9R1ku4NHZX6csYCTbjIXjoyZTbOdWNaJSordxv0XUQi
3V0L7HZtUPVcpEZAs2okGIZiO87nBULqtlklOa6gJPwBpjbO8d4bVeTaSkT7Ga5u
tMGp/sv4JEjrA7VPjMQCrS4tnc/NXKeJXio0PyNySgWRL8+sE2jyHaUO+E9EQFBM
DukXn1osigL4W/Py52R6Fu5bKXUL5gtboxNN019o21r5qQhox4sPutcq7DC0DQ2V
X489TVUu9dB008Kw5nTHQ2u9hxf2Fx5MHPNZQgMyUiB1FD9JVN3GucOR0olwifZS
H+Man9dMoBZMN0F6oQH+vQNUB5oUYodVYmB4tXF3OGsj8T3CSnLr3OWoJ77uPEHT
Fh0npkf4bMNa9lEGzoVGQ8Qd1LFJM7RKVuJ65Znv4ywWJwjLvBAPGsueLCG8HeXv
10ST/SDfay2HLGRRQE2Cd1/vl+FekMcJk5dxEBDrRzvSlzXumwYnWyayRu+uFnED
Z75rWkXrBVwOAdlGjqIAVwMMPrKiX153THnpFwgKokM4kPhaZzQSKGd7srstTSgx
yKHOT4nd/Q0xJnXofWTt8QIzswHjy+Ta4AK+VwxNOqSxXgEdmnTH35yWs99YblRS
QY7JNPbb0WwXCaNZl8gNawLv0IksOdgm3xj2ssxo/ussp7ME8nxYjOd+5bDA5NOb
Oc78ncSIaebGw/m8Oyyi44o4ExfvdxxMDllgTo05E10I8EWXLsdTUCWouSRKgAzh
WigOWP/d/aBu5fw7+TMYr+IIgHHhSHs+46BQlF6QBVZtfDYQiTdH8S51yDEThuRA
UiU2zJS1RFpsjWzqhdqJyGEopHYxwu9c/+iB6pTO9aL+HNiMtSyF9/BF4V+rMw2c
DCFviEEnSIu3rPVcfZ1H41RkMW5iuU9SJY3lmrHjF16JUYM02LAc8ZVSy0zBwp47
eNFAtRhUAASNcKTboWtWoK6YaPn/pHRu9BB8fakfQ4IpdqtlFN5XvxP3C9glJJMg
dVR/pl+Yc2UHftnrf0+Z6Ca6GFxFLQIUbTNC9C4jBW3o44KKTIpnRon1kIVwJ9xX
VPV4Bo1gtq0/IG9JZUtez4r0yzLWUPV7qmfbP0IWFfjeb2ICRx77pxx5TefABTcV
NTbGbD/snc5MrEGblayagRF1HfDl9IyEtN6Agr2Tff52/afUb3XeULIRiUlFd19a
00QAAdyzWzvKi7ifaGI5jJJzsqRvPbimaGc/776+fd3wKU8wkg8bvSVluyWoGHlb
fJOJs/fm1UtLnmeRZJLUncuH4jIu/v5YvT8J2y19zIyqSqClnocNFqewtMhWj0oX
xsTud9ev/y9BciKxc/ExLCiev+bgGZ8YNkJSPhpvqyaQpnCGPgI4XmkAvP5L+hGU
wM2j1RPxETT0cHtN3S1uoCncc0q0L1L8QWybDW27PPfmPzeV1TbGKlow/1cdApT7
SuuDvkmTaboYivAtBsryKQExr8zzzyRKpkUDvLPxpSMyoAkMJ6tortqYqmYdgS6b
rL6IUJoyvKD9JML5nLd5w0tWxKLP1oF5VyMlCQPfWy5vzFFdzhtZx6RR85SsGe/c
qY6ZRp8Tg5q5JMqhhr1T4exbuNTgieRoRIrJqsZctnc/lqM/UDxxrsrGaUbKnGWW
U94BEvp7dwR/Cvqs1q6iqyQiPQHNlpJrT63prVwibsVOfP9bxU8SSFEemH7EADkN
hXW5s7plIcmHvoxbFX/ykrR/vb+h5xNEgKcgypSSxCKT+iChzHcXYentPv91ENB6
yy7m+jD/LjqzH3LNFmS0H+pvauzOb5iBSdjP7dgvE++wexhR/5WiNjxbiHvFJx3J
Lztvw73TYHXqXRZkerqxrZQRtAB749FyJpXXW+oUNQMSHBYkUewAR18naL9PSBN5
f8+v90/gg51V5tG7nwZ8+DbGbSpxIIXAqPOiKjVKC+/GhZLP39hbcLfz7dnKMO+F
BFuT+7UyLYd1yLm7ZKfaRVOYNhgUODSN4/JJ26uetg5VsdXwX8cOLTlP2lFpbVRu
vSxdebUmyFPkHVyxGoa53yrSaTjNOSVfIUgldBsHMBt405PXbLrdnk7SwPPM3TI2
R4k/AprtHY5DMUpaHjpVAlydm55sY/j7/0Z366kdumpjV+XA0SH1xQqNBdFctz+V
7QtwgStqA3PnVUAI3D3s2qRS8ujQvYNvPyNI1Y1d02V9wbqJWwlKQnrbdbVyLAyQ
DXp1PfTWadf3GtYFN64f2a7QyXCvUAKlGxVkRiOT56PJ2W2n27f1u5wT7YlcPa+n
+0KzzswspMzz1c1enycX8l6QtNc4knxMZPzDBuon0wd4NYBQXdQm3190Tol0GA1N
zm96vyRRpDo1qX/laWhFoxIx33ihQY9nb3zdPDTT8TsUviwEeuaB0gvxSVqiuZ0f
jt4A3/7DKlfxHMA2KTOXj0Ie/fRt+30QvPpXir0vXywHCPDLUluZ0xqnP5yC0zSr
PCwGsYQTXFoMJmeCWc250XQ5SFhE2W0WyC5iVG/+Iw7H6Fm/4yXBvTGNVzriq0lq
+RrW8wxaaUFCuXvzWd1lI0I0G9O/xLXNsM96jf/XxEeQK1fskqpGHrqIKPqFdpm6
P2duUiIsiRh6zDps4pTZwo0UWBxEJLH2zSEMyKkDJHqGbrnGxzpFEDMTXqinbaOH
RR73OcHBlIXKc9LOpX9vOxIaaPupibrN5mKtip8ZWhjmmXISyuGPkr5OrSU8OeNE
Ukh4aoCeu8tDROBggJyuM62H7mCo4AyxCOdVMzQbMU1ksQjaLyDYEmv3QE3lnmL/
P1wyFN+P7gC8b9S4c9SiDsEW1C3kIUwpTUqmw+neVpdc+O/6GmBfSdcEOinohPo+
1fX6Rsg9Ks6e3S86qH3ERd2aiWsge5qhq2BlQt9zUqC5/btaatCm1Nfc8iIq9/px
3ov3aEzd7/tBSi5qd5S+gSK5NpjlWR830r6khvJXlELN14Q1EHq/s+PLkICdsI+W
eqbpHtyV8+Cc823eVk63MCUVIVbAlzra5SLFvTrRi2NxFc+lTDg0SHOzsTIDeY3g
lccibWbejc0hVx+P3n14UyjQjPOlNm4VdTuFRqNnn4jIwkYyaXyHDr58VMxKDAoW
Z/DzaJw7RuJuxapHCyoQwEyyJk+4Gl34Nu8zWEO+woPYd5Huml9blWbB4ZxpcbUn
Q2SBHX+dVvfEgrLZ1qDvcmdP062ktf5sE2Z2utHRgCiIjLFZQzQmxam1spW7msoA
tkS5bGv8c5IT51HUn48BndUOOy9A49MxKmyWhkmuPhom0r47mY21ZFommZHFOsWq
U5wF/bipZ81yKZZMWDcYQ0+NvdE8pE8Tm5RtSe8G3cRQ8IEuUs2Regc9oD1ZKYLV
r8YqS9DzIXGP6nvRRu/ZNNxWfAWEBerzx4G/bysRf0D3dQmDvpO95r3aePQFkvrz
+Pbjo9aL/IJfV6a0xkxg7NxCJltZAtj+6gGNtESjnY7i3cQcc3ptR+RkBHIpSDmZ
Ub3RvKV73awNJf/fFNNEK38fnSlgtvTAltCFDdPB8DwZ9ty9heGzYKgLCFzoTKZv
+yQsaTPpLtpAgKF3c2huS+ahqh69KjDUAJT8NMUkofDm7XBVoey821ViURqddqNx
qUuABuA6FYX9HfmMoCxVX8XNN6xQdVhJT/wETjRc2SfG6mb3Iv1jz8CzSZhqj5Qm
1okKVv3uD4wcflHNTwr3lnYNPfMooHWevcDFwYu2X/R1Amkt4LQZv7qhxO8rB/xx
+UdHdLvy9vZI+C34Rl84VxWvLjnBPCrswcj3J7CkAxUvXEyAP8p/+CWO5C9j7BqR
BiYgm+RRvbynbK8cN9H+oroag4cFB0LCJ+1Rb3iZ8OulcDtq1xl8oBrngsUQvBgF
D9wAREVCNXtLtmJTE1DTGoqJtQzG40/dOJza2j3eFN46+ffBhkMYbxERihYCNRKq
Ko+dIgtbyH+AhXTY4B/LkfQtIXgBAimfBYVRSktxjqTLcZ7UWjdaSM8/CoqV/6hR
t4DJ6Cw8SiwjhudBiSUSqq3xoRSCI6LI08ONemdgDD1x+NkfLvZvyN8K0SZxVhoX
uO+h4mzmNLuGACg3sK/aTfAKDw6B9ms938ZvTBF5XVseJDmH2ckSvED3csI3NLcP
Br6aqOwR4F1KfQiqQnQXmMfuXvvNGEKR6VqB0T+CR2JloKOCPdSQ1Er4hZElg7Ht
EjBT8PcJt+sIJa9eif+od7Lwuiu6xy1sIVBYQIstpP7vjvOphYFzl2eNpWvychhA
mxupAEUl2K2D8zWQwlEYYgSrVHxB5VmwqtTcdnahBD1t8B7aaKVsMrWqpaxGt67g
+ahAOH0Ay4r4ra9dFwY1GpuD9EgvHlQIQdXZSyuFdgFC3IYx56jBTRxiGEiS6SJA
Vm0oF7vLzG/sWFNddm4FkwBYfI7nN1qFDgMiOjRphFA52ujZdekMNMp47gfGRzuj
VlQViZmF4dto+FauojIKAYfOJba7x2AWfjYaf7c2O8zuEhIjK1LFPQgwEndLoYxj
jNdfYE54+fU4jsL3lflnv73YoXyzKfhB62JEPJXMzYEAGDwHI4aAIhKd4uIxVpQ8
/PrYSe2U7ISfb8dVSCuwgbyZzxHpdfrrUBJSfi8QCItioULB9vSXRAoIa5vJ4DYT
438/6AFj7EBWFqZGroA3oCakociaUn+LMKlWWxtQcKhuHpIaa8nYCAdFFrGjCBTN
2/D3O6CdYIRXygTV/ULAqu4ulQj14jLX4SF/y3IntM+EsRW60dtNt0Iy1NVZi3zA
zwe6iO8+tIRPZdH2Qd7m7mOom8HwPXUF1kqf8glCF0Jq5BXUjoou/nydS2h69FxH
NeXnYBQdxEbnDjzhLUOMzy9Tptaw3YPMKpn01M0liMqKxf/869anTZFfcgSmmaDu
qiagdFHuiYuxV/oWoWjlwk2gzMMw4hFCib0AczFo6tpEEmmpWNqk7SjhQr+PftAu
m5AvcbMv8sfzCLJlwvOEZ+15EvA5fLWwqLdSFbHF7b+OtdoXb+EOMP2t4p2BDQUK
GBKeiwnd4OKp40/P7qlm6648k3by8QNxIp2ei2y9Nm1kUbajJUGE7UXte3U+iYeg
NXxBjFMZab/TfBN870jh0fy73CA2wOVX9BZ3cboJxUyxZwx74O4YJDFUiWw7Bm7L
xGICT7HQLmRPoE09JZ6VueNPy4PpSflulP17DhA6uK2mcf/pSNlBHj1TpJzbXCjr
oRmYhIk5y/RrKhr/RNwc4qOnoONsfpmpXjCJDf3CwRc0o7mgxPJPB3KpgI9vGCq8
JHaA7D7STmiJYlFZUir9rWs0X4judc1/ywShEmljuL8Ymkouzyaw5xkbP8mjamrp
HrxA30+Ro52RBHJhu7IGh+LldmAC4/9mLUB9J8kugvdyjW1Fbl8NGuwbPsYLTVNR
CTmea2tt6DNRHUclXwxApx4+sU471NG+RjeTp4oD9Jau7COEWGCcsCQ2qfjKJJLl
De0dn4YaJZQ9bYapYAo/0T90DbCTS/Syof7zTdvUlf1KhFXDruXmhyao3UQ0Tt1j
AOSl5rccOZ/cwJfQKdYcw750uK8vMX10OXyxj+n23798qKtEJWDudlMniHlmebc/
9h5KxdjfMmbjHMEzH8FDLa1iiAzxyRtJxcyRjJukiw0PWxQ/iaDmgXeap4FZp9g2
2h83vR/hzGRpIGTlqLcehubWfDEAAvwgvzULTMo5pGH0M0jvJhucEdgiS7jxjNKB
WTGhcud9jD13iq+7SCz7Iu6kKdmBEV09oI0W73jS6YBPFT1gztVoqSMlIM6BW/EF
1YJfwe4gKzqAeLTuK+yggD3Cl42VKd+fCF/BbHDDYJzy68/xyHFdrINFCXvR5O/n
oO2bXVGNW+lFLvd5yEgJJJfHkU5KJa/hSUg0x2dtNHOWhl5jFVU4WLgfdSNTHCaF
LHNqToStnABok7oVZHrPXA2se0VlEjwIAzP5FlZl4sJk4p0rRx5jTd/dtQewqH0j
iLMKLNvQk2ZUNS6+yd8BszzFar9SDxI0sCPCVm2I+bBXBwkrQg44g6V4+xrUpp2X
6jsYTEXGLlhZ2n8kTMt/Iteq5hu4cROTZOhqBpZV/nbwdPWbcuvRRhPz54uv7P+k
TklftN3ZLiXvRIQQDY4HR0p4U6NydErh5dir1+YIVAxZzdKA2RFuPgqUYYlX/3+n
ju+OokzXL9X4/79SXY8QTiEJVAAZjWyBmuUDEvjnTI83FO+nJCVCi7+/3MoHmG6j
aOivSO3RLFbCYvxNDq+pOnHkPOSzZbmKgoNsMMkN5atdJzFUoj/UgAK27JxY+k4I
i2GRkuuvs86wAVASGEZTOABRXX2yM62Fh8eH5N1D3YYleD4K0PptivAmMgRkb+AK
n5tsWO20v9zHmt/5a4QuiXyheBpPPZ4htZHss4xm7XyRX+cS2qLKTQnpJAB4v/mX
zbYKpS/IoKKmTqWFJd7oH8eV2SQuXmNoLdv/yxul782WQcAZdvXDxE55MZeZ0+Gs
yYUBjppp5nUQq4cPeRXRIMNjNOxSN6GUuDdjGM8MibcK450hcD4AmLP8ah0wCVcE
gXiylw0LGKTXTSQ+GBywBCeK6Yx6GSs8xUUIxdW1chO36BHwVS4RRihYoPIVMcXY
bQeezcIFGSVMus7vbin29QLPO6EaP6fg0ZH6luOKYGenODgg8QbplrBMYH4WkIto
Wkd66X/W0A1E41/k2g+oK5tzEys8tJv5POa2vpvGNu/jiYhZ4C0lw5zrnEctdxYU
4Biom4TzXtOnZbquSrTn3kI75BzK4rJyoORGRfxgTps1ac7Qep4Ff7i5i8Tiph25
vjnVigt0qPQY8gvhr+2UZVOsgKglx/9E2P1BIGAGTNNMDSPkUmzfIB4O8VgAV0dR
BrSc1TAwemWg9gWYwvQcWKjJYJFqa4Yhwls5N8Yq7QRpqWu5g4vOy+zk6OqUUJZG
Pk5UtkcOnZQdEiwrfiBBtEAxcZ/Ez7z/CWUJgmDSbz/OhqcktqlPxCAQvXNvtzc4
lyIsH1sOlzwgzECwv8IB6iPzMMlDpdk9WMpqCFnHvuSCOCxosFyHhsCvqYfX/Z98
JU9fetmmd0O92Q4RM5AWoEO4RA1iSf9dYNvOW8VfGvq3Mxy3Uo7/w3xnKqHPZeVJ
SvWoDWXEcjrE3ACMcB5yzzT2/VcvdFDc/1EoDWPCOaaplTnEt9hQex9nseXhh+ja
qJpnHV7BCRd/L5rUc+mKfHzpE85q3Pxlmihy/1rlpfdK2V/c2oHEIi/Xjk1CuU18
Ewl3UEDrhgs6MK87Kd2Xe0hM5J6A2KpPIgrcz+a5d0fCTf/vxHpdB3bs9tr6tSkG
yFtzX0dF9TuHQrMjwrw+qnFXGUB+LtlLhDACeaHrfDm1AjF9g29U6c9wGzvP1OVS
P9ZmW+gdmmTAygAmXXhuXj/GV6mlxzqDo6C808IhUTndhSvCFgrCrf4ehlGWDvPT
95noYp0Y3PJiWQD8O7dhgIxzXAmDIG9ottQOi8jjFdTn2gJAAakTJWRMWfR8kAHR
d0j5Y8nlmqdH16CCy7i07brBT3gvOVYd0S2y+AqJ9cl9VXiOjTcj55TTDDX0pHs+
aWHaJhaqjz47p3t47KalN/rEhNHH6zttfQWQ9OREovTnbBt6wK8poOZYl9pZm3Br
PDMWWmLPgTPpXbZuCOPdOUbrbBKNXC/yk8OZ+hlpGEY6FgPoirW/PV2TWWXjTi+B
xQCaCRVW8ZN2LIkijnbd+Vmb5CEhOL3M0G4JfuStJ2qtXEFtnl1C3tyH7Gc2PG3q
PlsFjkXTEI56zS8gGRv7pjaqh5tnismefLNl4ev3cmGlFqxBbHi/9nAtdibK/0K7
h0ZcUS99X4mfy0Kt8qr081eJffYXo1vGn5n4ysJvmbm5a+q0AQUiRl+IS+gipTa8
5DidfN6eW46+uhDCpnVpRIEj466fgmdc/2PDIUydsQzmuqj3KFqNPGVBj8/k1oRL
2A3WDARh3AjPVwwbsD4lPJjun4e9Pj82FpZcrQloi1E3goxW8SoBMJRBaAfUiRqQ
G4m5gbLmtFJHRobtoaCXywzt/375920xwH6aisDt7xYSNfS42CL95NFyiyZowLQZ
YEGYpCrId+ancQe+oirP9scgB5CzBCRPHlJhFXwYawO+Tk7ExPdYLPyorrwj1dhG
bPv35fPrc7tjcy5HiSa8bPzhPEuWJ65HHq8DOw5WKef3FWRHF6z2JXKbjmr7MLFh
Pw7lKhjLsdob5aUkGpAvxI11IFwmodIWFV+Vf9njSiTLxF26iYtwUitBUTtXBlcT
HESqCUM9Ryzsq84pf0RVFYZ9Nn5O0EjYQPW8BbxWB4jKy04YdvFc3kqNjVjX+NDS
3cr5mnsmN342XL226y0T9h8So+r+0AnGNJaGby6Du5S5AygiwNOt2mewa1sBm+GT
T7J0XJmadOufMECNd0feZ3WnWFFdLITdKJkr9UquMddY2pMchduf5+7MrdvMRK9Y
0v0lnP/vE1asE+cSuM62tgygoGplduFkO82DIoMv7ZkmatROOlyYZpwTaMhkjN3O
4JWNfrORTwjkYfA9stT/pg/U3cL9BTnax6K2ML+8IX84yOpKxIuvfPrBjBWt44Li
OAdjv9xGvd0XrV294c6GpY3kaUjfegSlEhawbKMlvTzEiEXLYrOk5B2eiNYBvn0e
mqfq9yRZETD3CjwQcdY9ZDkUFwNHhx+iPD15akShVq1BCQomSXCDQ0mnogP43E7O
c6bpmb6jwHOyjNECj1ZySsp9IEygQK4KACiYxSmxNoCqWacsEbcaxUetmRpvQNmz
vE0K9Warj81ZysFoSYs3vSduVA0QsqpYkh19cQlx60ai6DCLDc9z+ANu9wWBQYTu
ir6eSn7alRwfjbagHFtI/LqhgwHEoKidIYIAQEDdHdqkdZ6o14bJ9F5XQcR3Odqv
3sreoJE54GHzBm6Se0IC7CMXOl4HNBq9lg+5P7cnwQAdlG1DvFQwSsYjAGxelSg4
81kOSlnf4LALP4F5WT8Ngj1Osw8ML/kU5DDywpH+GoqV28Jr5pDy6/4N6quj0a+w
UW69KWea6Dcz0582a/CnSMMEUZ5AfUTZw4qP3IeRdu2OyvWqwFIF7LhU0iUZEH0r
fA31OJsG09NCMbLsN5qPToh4UX4OuRxiqPiQ86WwoGi9Zzey1Myvkd+gQ3FmDHkN
/AUYylSXX44nn8i59F2UrPrKwrRrguUbzXKX48DeY4UFk0eznpgFCJ5JR5oudapV
vscrEbn04rkGSQvHsgbm1H5LguYu61GHP3RFBZAJs+rdrlQPljiCnATaOa/Ub0Ci
zdYGmb7AVygskDLxTOGIuWZ1GQvXrKuqEjoLDLPBEl+etPE1i2zGakTBkqwG2S2o
JbmfdUZfFgOl6VlPaOmorm5MO7oiybh5eNp8u7eN2ZXWn/7SU5obKeXOctaJXSnX
e+Zs8tPUFyoLhPJU0kq4WsNzq5GuIOPzETJOs5WI+jOjSq4HpxyV7WHCUYTN9p0T
1k6qCUkoPPW04rkKo95vQ5OSMcMUNfh6hsvB5jOZo5gWIFZOiuoACrNCuXY/pWza
FErBrPDOhweWe/dlCXJ2B9bTKdxD7y7nXBNEEg5HiFb2LYFO6hvTSM4lZr1b6HMt
mIB2wJ9NJnMZZE3hP0KaEvhfi99nNIUn+x9tyMiWLFNfYOTH14U3KL7+nCMsSe/M
nCoiDR2+s9Skh4XS3ewnkd6S0HrSLjfyrDpV5bU69xVDR4MHcaCKSG8k2eaDJpEP
pgdBGrnI4oMWuBAv+3BGXXZ8UuMlRfyekdsQfuuYS28tdo6mnT8b426opaY4CZFX
EdILhdN+6asFoDGgBRfynqucACqlMYfkruMD52GEZuuq1DMPfy/WL2k582XXVSi2
uHAfbeuYc2wFQRoH65miUtgu7eWlCfv8Ij3twruGNa2InbNSynpGzQOwNoRLdWS+
pvjqVRfubc0kPaQel1g1Y3suoCQrsvx62FXpMaFvzzrQA5dqRHh32GkNxo7AwU3e
G1xM7k6b9fGCAFofHP1CYgYTzLw1JEpaqTM3Il17cGDT4pxLlI2K8+siWKRYM/Xh
vE+MGnVCdOExpAfjTbVFsCzyWqoHskY3gnfcbxjFCMEXLxY+0kaPRT4Upkk/NGHx
zok6tcRVSONzEmFhYXYuYf+QTveXk+x+42nCbo+c5o3X4gtnNNSD6LfHD9dYz+LY
aB5fbnW7XErrJjlKp27EPIGRZtA4aslx7E6psqS1yNJBJSArkcUiw6566yAKwel1
GeMqiCPnYTXtRXbBTB3Nh5hz0Htj6TqTd7LZD/gP/z7rv71gxl/wCQKKarlveafK
ib15ediuWgmzdHA7XbEpRvSaD+uLhImguyiFb7+ZK8Cwxu1wwo8sFSEjD6IKTsSA
ipXjowQE2soA+sFN7zjEwTc7kCf2bKL5agfYDlzpBUvO0hTrv8SkaoVLx2pAUAN0
3Wd3WI0bQdgMWHAJrV794cgWLRJ6c9F3NMxRhJFKFg31d36MbD23Dv3tosNXrCGR
ynZ3Sl0JTVIK9K3KH+uTaFSt4ugUGktFTQysUQv8gi8Vt9GVWHI17Bg4IvtccmgJ
HoX8ZLhMNZ5mlAFxhLoixDDqKNBc1DwkjO8tgLTQLaRHMCtikrUPYkXEMyaZvvIG
BL3IMvE+y59gee7/PF2xnaoku2au+VRaleiTZTLwftRjsq3tZ/tZeRB/A6MsHJTF
ABQ7gH24Tjchg+3/vFA82hhJEF0FrDiIITS3mN3Bo/smVxb2saTthv/pEo193YqN
I6chXDh9XIl9S7PXWqe7ecQceQ3UgRzDXUu7P0uoh/4TS49aTZ7eguh0JfJYRVLy
0qgI+MfgYpDfN1/eBJjLbMIJpeUuiaTNZX00NYNlKzQjWnhx+j2b3CyI1DOrN3Tt
S1laBRWbV7osp1icf5iIYYv0MKmgQfAzFXXymFr9iKxrRHhsEb6kk9NeuRGt7gI9
Zr/mfFj54dgJNEDRoKcnu1VFtWpG88biEzx0fN0gfwLuGQxOG/mGcu1xfD73Krxw
vG94Ctqrunp1CgnhmeZr2js0CwUYX2WOcFsts25oNfp4FJDL5JcsF+TpDqRtZWi/
fMGw+qeSTkKqVIYdSJefbEShMNavG4oLNbACbkFYoS2l3XFAJeTYtmbi6cjSu6Sm
3YlPvPbfeSjre5QzkwHG/1IyzbsFzQce13+kSTcEw3Djlx0aSSjDZvMtjRWShGK6
+U8Tvoj75Y7mj8rowoZh1hLHGfPDTxYhLA+ud2R3sR5oQ7BxhcEVJ32Mo/TbLinj
CwSsovw9RKvNwWXFIwhJFKwp+5ROzL3lh+hM9kXC9QxycbIWD/I3ot9tupXE6P29
kdEfuJgAQE8U+jx93B/Vhzpea/XbznCZDAX0jSG1EHbYDN8NbtJ9IcZbD78tIp99
fu0qZT8/U9rd2MKaNJu9RvNL2vaPRX3cU0y0xOQaCLOOIjrkU3BdM0+HmwmJLp32
zC6TN+pwDiUxZNm7zbZ5FqzQasRNtjDT/rcgscRT30QXb76oUDk/iHG7rUZ1x/4D
pu7yOooGNYvujHzafe4g6h3oG1lJqaS2xF0tc/KeFNrIZQio0yN/aVAXVDPFKOVX
uXWpGO/voUr5PsuejgvmJtsjU2DqRtDgDmIcGzkZnWtslYFF1xrtZhiLJzMZzsl5
q8uWaL/e351v/oKF7BBHdq3vq5olE85OUNKeis3218N1ZN0c2vn+0tI01M50rLyV
JRfAPFJqR6gqIpB4nVsd01ymGe23UJ0b89j0u4bVHkBTu5VzV0RMYGDV88M4kENU
o9zV3TNJrrkskvLsVVJSG8ZDQhM8MzXQzG3VtbJ1fgWkFfp+JfRU0fd0RA8noiIY
1NzYvim8ejO2tFfZBhEToJX7cxLGu4QeyXbwfOMVCyf7pmKRpkcSX5+z6V7Ip+2G
08bQcwzNMUoza+npdf5sO+hfzXKg0wb0r8kwpmKr+XEKFI7GFVvSsl8gbV1/0fiG
PNWjWE+j+tyzGaPMlMioCR3kWonVK85XuUg4bHzZsD+nFbtbGtExCZSkyDZs57uH
1k1PiVsj9n5LM1MAoL0rd9kdidNUrs/rdDtsN2oQwTAcHmVApfJqx9Xs/MGXOvBV
w7HIqDn8LrsWZYfQkPsxiDInwfpYMIMmCIMNt+rVkQDtF4gNexO4oTmSlgS7Sn9V
e8xiFcLkSOBxcRdWfeJ2UpH4pYC8dd6xpU+k0AM592uurwsrJZPLp8JuVpbN0wKf
/Sud8lZmY5qMntTrnnqyMa6E3R8BazLb7xHg3+K0mKkm138Pkf5x3a/R/yj7Ymct
apYqGRbFJZXHA/UTcUraHdxH9TSC/7u2uR3pAJG4fzg640Em2h+qatsi0u2YWP1Q
2IKHwA9pMqSsjaACCYd1Q0XxtQK4WXq08mrZ2KHFLXfMqN4sfxek+6mKJKXKDG7l
jSUkfws5swPhji59XUTCI6/VmTxwSMPp4nvhdjbjlTkMCywHqNtywQ+DvePm6KfP
zmGq7b7rQE2qySKNbElamDdTbQylSA9XOkwP+NsxsjEHQDOgsOPMNu0T1t9SRWKQ
obEJxymek+/vDm5mxcx30q11mJvMvUdNKAjezmXWFfOFQml1yy9yVBXgZAnmgWIm
02D6XNpeVniKhEIGEac89GFn/IlS5Re1aXUUxgZYCjSYfBiGmGX8mWt5MNnCFfbd
IDsZzmJKb++GMaFqYdVMXPu6pn1sK4hu3Nu2SYdvbBjOIKdEGlUJjrsaYMyP13U1
O6YLFz7qYaMYjP7pWO9cRDh/IoSphrOAJ9H1KxIvI3ZZ1wVcQkbWAseyzQBHpgxy
yzvv2n8GZsiLzPzGCNdJtoBdqbq6gFfWoEdpC0vPSqAhynbUs1jxyXu5+J8USmhe
BeiTxbVLoW0vXrWr7Q5dd6GYUB/tjK38Tp0J5vIhgu2zZjX11sK5xe3OMMgOsfpq
epXhAkbG3bi/xGuP44+r3mV6WSYTyskXLPlCUuDUUwa9CTEm5c8Q6zmAI9Cah8hx
8pHdNbMKzLyLA9DUwhNy459EME3Duo4aTddPhs06I+Rix9XvA/qXnO3xFXXe3Otz
6oVSNEHJ76DwJAUoMJwGBJQZxcmqE/JMCk3JwPoBmQ0mdv7BZiVUwFXXSZUAN+Rl
jqe3lvx/uFfc0tZdADqOiMqV9dLCupkK1tdrtRjsYlUX/UQlx8U7mj3iOR+xEpFq
39q61UsGa+QSAF8MFm0lxNP4vNznGAHOXYS81jBUvXSWDzLnhuX6BUMR3U78LXlL
p62AZfMJtEjVgKHSPEFiBTnbalEsCATa+L3jbSOomiuviTOZh/qkEJ/yipKUcX84
djOqjn7c8/4k4EVDvhv2dqibb478W7Og8x+gFXonH7XuQ373Lg/9lAt3OzGMB2iN
553sUdZhvTnUsnEPMkkEj9igvblsNB5aJCMnQHKAH2nrphg1Ob0tWmQHiAXeRsUh
sMcphgnjb/7HJLgEHSRehUTAVsMtzxaHiSx8VW5awyTdePxK/Ip7UJPDc3y4zNtx
GwoMeVTXVL7T1WnbIxCXxCkExeKwAHTn0MFdtusNyYBPnrCj1ow+MsGkQmaYP7tT
Bp4nhyaZg8WWTSuv9BVHGvU4V9Qg46Ry6NgFQC1InAhWYfAOselpMeqJJSUIo0jg
cD/jH4DmV9dRjSmv3m8d+mkKq+vq8VhgtET19LPqUVGgtAGvB3NHW0QGegRlAeEV
JTAHTWymM7Xf65CFgnhN3Z7BM0oJc/kiR/ox2S6B4ffAMJWxOV8HtQ8MGezA9Pq/
cCRtDGXNismsBZ6TsIofnc08DC+E+dFxC5qaDER6itQfZ0GzHbakKZOMOYxyaVA1
VMnakK52r05tgEmTQFTDaAQ++HZPtLY/1CR5Ve6TCALcGMQoek1hVhda2i118c9O
wF6VD8F24O5GTFBXss0QM8u6g6e/+eRzdcdNre9F5ZwplwSkDzE/HoD+D/bwIWBZ
JpDUeVcNR/E0wpvf1bvtOzfxMkJ7ZcuyvyS8PUZtuI9n0yva9MRAT91bpD+PSr5W
DZ+rp1AVHD6KmlqgS04dHDun4SCmJA5mcSFmQV+BIPV/TI7U+apuHAUQpB/gvEbt
mpyOZuMwrP5w9swU7n23E5oAtLLrgcBOcUhZ4WT2MwWiG7bCgopBSq91zQnrG193
1mEe43t3JWD4Iiz2FD54ooDaDTjlD3QqF3GQzJC9LA143uSOn/Kcc7uBQpk5/k2d
Dl6Ga+cJtzwEa0R70+KNyHERgDyBfAVjMkmmFX789xbD17NkuDbjB4Php1cv6IXf
qSgRyX+Gtu73HNZka5SQe3ilh8GDGCL++gbbXqxwANtbsP5tXPwHFkm9H7kZBVNG
CJUFgMAlhumddKtBckj85JfnL2Uo0XtekUu/D3xDIx3eMEOAdFskxamEwc/Px5QV
Ifs514Kw1jh4Gq4QucFB078arK/NPncnh7I8i0+zqLWx/OctZq9jQLc4EqwQ0VtV
+A1X8WTAz6dgmxD/8tJAlbM2ba2oEtw+Cb8es42BV2uBEgCUNQZ+bAslT4YiqvRm
uVtMrS/Lrz2DiK5E/Hm4MIocXFupAl2J0eodfwXlrtwPB4qIrsj1g2K85vgAq3GP
gC5r2iUjGqB1f6GqDkqv6dXdbAh9WOydO2Scn4Sj6aX9Dq7TDIgdknnQKoRlDebm
klu79kJgavyVfanWkZAAxg1zjTVVCv2201P7oqC+8nbBvJQBqHyTuvkiuhftiG/d
1oeh98BbN/BCdp57HcCV/cSlEzysM7AtprPj1DwaeoZduDsQVOPn6CgdZzzf16s6
Cgr9LqG6ps+H6kRSQ6bFNk+WDpu9xcwwCjQx/nc3gl5vIsEZsvOKGzsT6Qy9qZME
ASr9q7Nqc7ZM2tfoCq9oflaay8v5JKYcZCF4fB6324ouVpZm7NifezU33EdyeVfv
60a68xElcF4OFL5arbwXmncI+6e6jev188Y+VdFBAec3GMq35ciKAQCOzg0UTYXF
ROATAvI7XmKHRJA7jzwYSp2Qdp2AKSAP167GJR/vH4nWlTrR77usez21gSRZgOTG
RlH+WKnIpNU2UAEoxLAgF0jfg6MTc4XwejLOgqLteXjp2+Cv0N1XvjOmR3ubZ/Bu
0R8NssaHpso4DY+Xtifef7BOlOjajafGS1gNkZmMp95Gv6jWRy9cYhwXk5lyiTDC
JOOoyk5XD46zGKtKwTZRoS3MPS48qCm8ieZTebz11JS+CcPuJsTVKPIhQ5UUdO3I
FetcHBK059Ul3ePwO4AwWO/mgyfkciP3qUo7YGBbdsOIwi1On3+JtmOwgTe1qUSn
JX+xQZMxDZS/dWzz4xwHTwnMWST3fWivjrRNMZoJnVIx70whpG/7AbiIt4EFskFB
fpn+IJvJNGW3F0NkELdzdS/l2/GMwz4JkAycZhaDHwXAtGw80GJ5w0aUYmhoX+ic
+TSEoVnwG5a+WfUG0unXIe4XxsZP0mWN0GpTlknnki+6SETXZTfsXUcZBpweUKmW
DmpvhM2BV65oUcqFpbgBUxJbAazkaENrN0mDxxanNwD7KVckPuBgDp2a4xd2XJQM
qY7hql3UvNM32X9ALo/V1VetUYTxBvJuYCli8MDmPSroWCgLN2NMw+OmylxSpF+8
ISuyzGAFvE3DM+OvCqtoIcf1FUORRAfTbiQyC8NhbGMrMsBNbLoilUGZ/SPgBmkT
r8ELgo4bHRMpnDAjQ6OP//et6IhKK18A3wPzgg7WZjYPvNlzTbRKKsdgLIeAX1e3
s0VgC0GWu/tzK4f4N+DWdVoLK6JzQLsj712s4fes7EDZVvxshxB+sCY0Mi2FAhW7
TuMlxg25Zcs6bkjmTEslk/52HWro+ZobCIB98Gq5a2l1ikXX/e7kcX8sVvyAdRhA
jvhcd6Vv5Y8omNvDZzIlOxjRRtxG1FDJw1ffi20I/ICygagkRUE8cbJnt9HJfCa6
PxcXsaEiO41SGE3qJzS5d79ssgixFueOWMQPyd4qA3RZDT9H1MWeXeGpxzMKlLWH
lLcmrWjoQEot1pQ03sPNi++/44d6CIjG9UvBJMEreqKHQfmwfNq1otmXrPqSx953
rcUMTsF3Uaw7xsD1OxW4iicQ6hZJCD6mxJpyqTzJcNgaeA+dAE3sHTu5UoullZey
9gtL+MZQP6AA2WWHpqbJ81lAEeSIFyR2tTTOVfv2eM6WYZNoIUSfeKodQsDszLLY
GTALngZEdTM8ofoVVI4Yi6AIciLDj51koYPoXnbWUBczraqf/s2LXPrE5WCnixFF
nj0dCynjVAkVAPs5IkwzuanjrZKlcnOWMcGXmdK4+2mXVkqb4z8m61rgbsDdGl9m
+RmsS4ErMod5xzmYGpgspBlwicMUVNxgc/fgYNHxKT8O46+AR+MvtYjFhfD4pg5R
KUFc50zUcwB+l0C+qOf0awDPnZkyykWeZcrUjapF0MYZV10eEsPiHYELBA+2bmbE
t4gk/pIONR5AZ2/xYCLKK4zsZifsa/dwEIzE15IcDTz8bC3pa/tMemcw75DCJk44
1nXtl7sFZZeDnuZxOQfl/a5VegoOWSzlwxRPfzpu8nJU2379vnkExxQvLtkHsC8E
TQo27ybHQAavxKjrNSGs5xfkIknYa0TjvCyuqR8pUDWOEHlxLuc7vwW6FCU3q7DK
T1whdVhCdxpwtUXejFFqYhxCA5L1SzlAtq21hDA6GjodojAfp18/tZzed2trqHw2
I1tPLFB6jHLaJEsQOvFHNxHJsGj4wULlFC8moYAVzC31iuQQ36pX1zrVBxTpMa4y
V3LNHlCZFb+okmeUuZjMRRjctzTAGgRniyi84l9yMmOe+HO/8uAL1vKUWHMzgaHD
5gOaHfF8mpOsH67RC8/J9uq0DUtP51OwLaXE4Him/XOenJerQoQLBW8R/yMQaSjA
2nGsDry6IfjKt+6eouD9TcA88kHlJmgOK1oHAyXJeBhPyp5rY/BZOOA3OILOmtdo
y/YA92xr2glf/k/YKalOwcZ5JH91XSXgy9WhhIE+Kg0obiT+P4viQvAwQj8fGqAJ
EOOlgsPfPkXOCOpYyTPxUgADGV6skzYP5lCMM11RMPpwe9Txr4Z98vTrB6DjCJJh
Rqi5UksnfpC/W6RxDMnYV4WGbYzefi17q0rPA0NZKCHxKUFELwkWzPbO0k7F57v8
Fu1haDHsxuHJLT3dk3f23ceLB65jBsnimUuUx9djqeYar4TBU7Ftu/7cvVhZfmTL
bEIgeEavPqfbWfgTS8909TJ9gMhllowxCmFcTfqn7RidsNhKTXbzke8z8GjYathJ
HC26PxoJ0lO3r/v7LW0Uw4nTfk0QJGiTbQTTj5pcTeStulrQoUntStdixbIFl7qz
po34Jh/eBh9EML2g6JQbaB13zIZUjPQjIEoDNcjFyalFHD15AD2mptvpDzH1qreo
tfTvlfILi8qs+3OZ65QGGI0tstNIZnUHlKi99G228/vk49CDWl0LJs950dkZ7Iu8
OGjB6bOPkm1YeVKeY8tSibi9FLnGUxAQNGHxBTYOybsjJLEUmnBAN/SVLGU26maL
p/PBXhjxzrhE145jb63+FuSRDpgtjiCwJGv+fRKJrQ4/xlRQyJygcp1mMCL5WFSf
y4KfewivszixrffeDWh0l0dC80Lphcdw+X272sHuJVQNvuAHW+4pWaVRQ1mBtLuX
7UDNcT50hwVC/NM1UFJaxRBW9jv4a4nl0YCFGiw5vD3jgOqp1XEytigpdmuNSXaC
SkXa2oeREmxIjskWdJVHYP3rn2Wz7O8Qlf1NZoytKV8fYBOaijhJ8epnU4x5aNDU
XEKkXd18xMNvdjl7ff+qKX6lyPIedrD6h6gBVHYdzyH6ZyQ0nAwvP9PMOKUyzroK
mXlhmJhedbkBs2KLG9u/207BpSAIy7KUsN3ZFqfoUlXFRZs0jBRGMCIE5kQgWK8m
hFIemhUmJjhopUXq5yHJEUtuPPxgIO2IORdoGlFcGKlg6pQCr3yqcG0thoS6++wj
eZY3wApkUkcoYaaSzWPwXI3nYHYNxQoIXstJRVzlKASYtRC4XHaprz8y1FPbM59h
nAc2dAT++03t7Z9hLe5V8Jy8U5gr0V7jKtHUu/eUiqlF9vEOw9s7dQs0nFKfmN1K
xSWJlpuoluKw6BWEP9oPlsapvlpFrWYn9s6HnKloKvQtwGH6ZAOVRKfWjdhPaxra
kruafk1iF+NMntm5DL+VXObsrr4IM6cWVq/7Ak/vnQPomTSJGPImMPYRJrx3VQ/p
imbMQBtYY+S+oGjE+LsEHE/+aNH9h4tUh3jvhzkWaDb3WVPlg2mra+DvMVfy4OfB
y7iJw4+0GFLdVJgpEDo9UNCmm6JJ9RtJfXZn/8Xy46cZ+WXwyJjfH6iJk0kaG1Y3
660VX49J9NmUJfGnwJy5TMwjYOupz90MBRiDPOS2IflukBSvBgLc/VAA/XyyuJ2v
BYCSxKVpTWy0oH7rTgLC6wQU5lysJhHjmZVIqhd4oLMPGQxoQi27sxHwKYURxR6j
E1mLElHJLj/QGIz2HN8F/4N+fQ++Hwwmj+pDyexz/Xt9IiQ878HcBIBehvVUYXks
/SkEfPN09HTiQka+pF7FozEd2TrjJrJmQAF/fNdTyNfHQ6iLjiqDPUzN83tpKuz+
b6lNDFHwtrCIlwuj4jaa0wynxFz1pzZ+YM3Ci1vHvqisd/6viP0kl97uKHWW9SKd
YFprU6Av/z1zTU+7HtIiyZpzGfld6NzBnDKpxiEcHlceih77KCag8xTfPDd/v7gd
V9N2Pd+apm5mfH15HOBRydjVbREh6xw3GF5aKsaCXslYBIF3fypmwq7cw+Ub/q4Z
TJFjNM2rIoSVBMUeK4AkjPD/0eCPnc8JKLMn90vmOxQyavKQMPKTPfTxcMasTvtE
DfGvhaITnEBo0mOvT+hXFswxwMdiIGI19B0/9s67ooRUydcbIH58dwHo4vtgsHqp
YMInHeHrw+xlhqFJuINSeI08IMnMp0+ew9SUUh5+UMqC1zNfVZqBr4rCMOJz+9RE
wuxWArnt86UzWY4VlLohxcUvOzcSQAq0Un5FFAPGLo5kL6kzv9N2eB72gJN4jZEE
kiPZ7LbgFx81igopKRqAqnL/ssQqtnr/MeJngIDVAiJr7DSmJMsK7gwiE9hk+oU8
2T2kV/zVOvMN7L48t00nuIaYeyJCd/cd0UZ8A0e47seUstKbb7Xo5I+eQ9uPZAd+
KvM3ufYwuDvyyqcfEiJkHO+jOX/9+XpPg0JqI5kzqSoeNQMgQhENSxfLWMbItS5V
jLpy4biPUpC3cWCE2P3tjmBVOWWo2pDsc4VnxfCAOKbal02OwxNJeeRCAirFRiMD
ADhI69lWk+OnPnUVsEQR7pswom2d5gBFvL4ppIbgK1Oz9h1MHyRkvbMS38jv5equ
VIZvRgZ3wHT/QNoWNZ85NVr+YQpVDBPa6J474Wocpd1ND+VXxZNkk2TRnFPGz+yE
o5O/NzjEDJ10ErirPxtp86YzSSExNecDD/HdZ5xJeBKgBHbbIo66PBrnyMexJg8p
B+QHFHAyN8L/KAgay8bvgea8qRfTH78fRd6oTgqMCH7v78DOiR5AHZLMAPhBr0Tf
b2OvaDJ2njPHG5V9zoa7+eMMXlCFtcdz5RXXYf/M/jKVG9255FtP9n+CvzwfSkLV
ph7lZWtuT5DW+/wsDxyFvo04OKSlqV0zpfQMrWO2poCLogV/x25/vSq1pkEisWJF
SgRM0VCsuZzFYZpFFGkg/oOOWJVOX3PZB1WNkc7GVA1l0y4NaZ+eDTaH+cobe/28
iS42XPv8eveR+L6cCdGyUHtmU76YuBNODFM+WPtWp3yGWhEQ379DSKDONdsapS3a
A7g+mwkfcOdzDfhfSteeE2oRc49wj3jEvZboJ105ezb86cgDLsGy7+9kj+PRQYCq
sRoZFNLS3BbDn3ANH1u2sMOmbE7BZhkmOgrWgV3yJ1kPTglYExVtPxrAiur2T7MH
YwKQH+prn27SEVvMB++aDHYXr18W0t3GI6EH5LGV4KhuEqzdIdIb37NOvktsNhIJ
Hxc7iUso6Dv4RGlB0MbTmFhae6ONwyc8DGjYQbka5EU3RJTtkYngpU3MVUsOO6qx
PA5NtbY+RXTZq2qqo2Z9h8BYKp0e+hxbxYvmxiKm5IQdsX1Sf1VVj+MD+HZZiHvu
tcWKW6Jrs7ET725DQBIqs7WF8Q+11FzcMLaUgMJDuflSz19KhPUqjEzXI9S4K0sd
QeeJ1DyLbfbUH8+un5A/n9w3lQn6VnoPCY5gYDNjxjlW1IZUoxd34tTk8405C9x2
1sGhaOcIhSTBIDGTNbhqc15me6G/1z1ddlEmsnNTECIZ8VMEwWhgIQx4aUfIrLcY
GGRnPLuZWbUb0klDc3UJaKBp5DOFGzDQqhguqHTxFBOMWJ/fmAsdeERUzsmsOCJA
hjRI3QMB44xmiuICP1fjuz6FfuJNSqxSkeDVIsOf0iGzW6li5fCtfXyrq/4zpUmo
IaDRKG2ZgRbCivZdFvNLwkjwYUBAJwD/GdPaRZzYOltIWUx0jKBiMDHTRwvI/ciZ
Vg8QUD3ZimIf1w+X60OjrSoCjaQIo3427eJUwdGlKEhrdd2XsmqHPq4dDX3HgfpV
jkAJBHi5OpAjCCE1uGKU0yabq2fier+dAS1Kv8Q9y9JatUo3oRDEvXHYqBraxCVK
502PD9Jvnm/WY0CTf3DUU1iZesOsim2biAnDDk/EhkiMAkUEelk80G4PwDeG8UFJ
1/Em7NZ9Ivn/wxHchWG6Pi2/16MPjjEZM9I6ZD4gW8GLlS+uHb15NHfrZ5KOenPg
7Q+dyHrr7vHRpoDRbydAIvCbTPBjjEAIh/sDJyJFKFiRHX70vXZCNO7+mu3YAPYA
RUb8Jnjm/F957Rp53Hbav6pXiC5qFXtcSLTQbXksMFiBsB0/u6jkrHa4zc1AJ9fK
oa8LGNeyKIhjUFvP1E6Bf6KsSIxEHgfgteF6FinMzzubV6DwavRyL9ZzBCQWkZ/R
/51cp7ejcw59+6YEymdXQQA1e4LGT3tB61kXVgKYkfBcoUA5rStayvAMoI9eygCj
B7v3DjHHH6vJ0fKesM3cr8Q6oXWheR4JYxilC8XSGEDrcN9SDcw3mPsJRI7JVI+x
u+nl7ub29nsiYYuGs8RBc7wjW+Do82q2QTcP9gpTEf5ooOre9erqpF61fcQ22gFf
LsIDyBNM3ZGFMSqovcd+LkDSlZ7DpBOMQEFlAe4aX++YuUseOa6azxJ4Ki8OFXq6
Nx9bO9MdzwGGM8Rx//Vb9TLO/rt6r+0ydSrjeu0jrCMh9CyFtF+Q8mk80DBG2NWG
l53wITZpNQ2bjxDItgtPt0S8aYFlseYkKN5fbr9BMXxoNUhBLvbMdAUYk2oq2Pyj
w/NiHaMTSzncTCRXK9upzanxPOQ/oOFt7l+G25C2Lt96lXQ4hiR1/6B9rlUI9CGM
jF0Zz1aE/72iVGmvCEddSTpnN314xfAuiC+fWsEKWMHSdVAPb2yoIeqrScalcQS6
LdrP/Uq052Rbovi2E8J8MJpVvJeocsznmUah7zsv5p3t85aW8XrqWGgXILWxM4mL
ZI/XqpMtV69FjRo8v2oPVEGQfJ505Hg6pVUjNru3vK8mu2n9oh+LOzYRQx7/tpqz
7V6aGSypxAe7Yub4bEoAX83degPfgcHCka3K4hfFsG32mXwnXTYaABn/NuLYSsYR
T6rgnQmnHUnozLsxrLwuQEyKvJv3m3E7I2eA6MbuR/ZbtrT/sHgH4iv1odMXq6LL
W54KD6WfTJuljTFuZTGAhmaGr8u5tWcbGHiA/J3DSOhhltvC4RkIue0Ltkmam9mW
XM4oTNIkcpFtKh3ZR+t+JLGNFevfIqdwDP3a59yROsjdZryAtneHBAsNlZz7dULr
jQ9jysn2a/SJTvImXSzEJXBcQdWJXyd2d/SWAj7D0H2vqPSYfkSPaCr07ZdEkvii
KUGCuELjggfaOyL77hwz4HVbpS/6sjkInUsqnMvP/FNfvGdkHj9h9EfTY2qoCbL8
v9n05k6q2nJP4ZNsG67TzZWB+nidauxcPl3rFUk8Pv59R1gjKgNOwDY5E8vYe6Uy
bNOqcXWUoBoDd3c2KnMVOKymY8+u7Slgts0ng4PeedPNurV5Xti5V6FK+qxgXXUy
Vt9mDmp0UXqX4u/29/+5/xDSbFlzb2aNyUE3cZd1RWsM9e6/MHaBErEEoi+rqPfv
JEmKH8CK/5f+NBapG2jP+/q+IA57DFVKUUWO8XCmD9II+F47CPqBg2ml7JMcyTku
ml8EIXlapiW3RT6FYjdq1rNZmboVuglQBRSeiyII4taGE1EAJkTGcXFHbMhh12sF
uV3AUFcbjH9/9RLbfZegWWTUQvvK6MparH4rKyA+Ls/OCDdFEN7gmyTu0GIo6P2Z
D0tKwyoPFEG15orLdAzwsRAJDRUaBHlcksDWXtwduerMngaiaVNdLAnblAKPG1z7
kT8KMoy1v3TFbU0AXprjs0a8Wz4/1VfXSi9Nd5YLzBJDGaR3Ch2ywCeLuYYS2ejK
k73EmJe0x+Tw/53X0bynVbYk2hYTUOMnv9gNWquIVr3OGxTA6865Y2CN9ubHW1tZ
F2RhRoQOcOTHcr0pmGTxt/26Dqmic4IyyYPggEMqylA5CnrqJVJgJDMKMwXsAmkq
XasLhLrEU5AlTB6mSZLenYCQ+WkLiNWYX465NVVeV/+XmTs8pLzZ0u7fe91309Uz
IJ1fybHAVy5OWYxLDpTvPsndrYG87QaDSDElrJxMGl2yMk1ozejBSTvKh173pUb6
zEMxnymC6CzERg4CoLt1LYLqntghws6lWQOtJrcWALE/T66n1y1o4C9f/SAnA7RO
6T9njO4rkbBQhXFp7J9d3QdMqH/ilWyRvruv10ko4DmDMqGYT8POvKI6xo3LdaL+
MjIa5cCrROdUjFVxLd4wqVPl72JbckLronVzsf6VDOUctu5EzDBEB1gwYUYy9PvV
aJdBi+/7SqHB6CXp6pMvHiTaJ71Ps8ZS1iWOh0U3eykV2s4p/pjkAoM2FwnX1EZH
/tbCfk4UCjHfKMCIQKZuJly/8eifvFEmtocdxAbYcRGjkwWs0yCgXwitmhs3GKNJ
MBZjXeZCW8fG4h5fthV9BDrO45Z9WnIM8TPVc10LO/4Ht8Agxn1x8PIQ5nvmtJ2F
KPlxHaM1NVyPyCE234o8q5cV2RuO5vqUKh7AwUWLyxex90CVc43RfojuthKLzFPg
ccoYNNdP6zpcYjsHFjbGK3qCbk3Smd3rDbIIXpcaDgfXgF31hYG6HFadVKAIfiAI
TxaGxCjJRK3fXzBck4VHrIN/aG76KAxxDw7a12ftugut683+I+0OTsoH4oZwUo4I
bHw8sSug2t2fkk2murSL76vE3Kp/PcKMujVwTbxh6EDVfML+ovH+mw32x7xyEzym
EB1h1RK6lAkTgSRLR7kL/00M9aIh7cxcTDP+YoSk7DhOSarZ59IvNIMb/tg0yPk/
qHHbg/VuuAb23aHOlXPuDsIBuqc7WwnzIbS4+1WRUIh6zqDayL8sWStK+6teLFHF
KfLr+QlLUvuy6XBaP2NC4sDw1THrHEetvjOsxWa6srS6OGucnxIWltxf7Nh+0RO3
k8K0coGUU+5s4jTxCzayJaeYHQccATXm4N5MVs8NEq1dZl53h9ap5mGk5hxZoy0Z
pV4plBhjsu9/DhL9Ga8FTfX27fxpO77IU2eXk7F8/Lygtclk9U6iIeqjIkv+EMvo
jp0/QlRgNWrZoHIFnnCTC4pNKjeAAs8FRKy3DCg60wZPxDs7Y8ZXRd8kNvXKyxNn
2fiGQHfivDeTXOvzREZW714PtlWxN67jl+4+yIPfVXH2lMXDcCdLWYXUsKOH0mu1
7laY9/pEBjIOnTXZaGOieowdxWeLYyl5VOzSVDTgd0SMCKCs0ePRL6S0V3gCxHrh
Sk2uAQD4p3MCqDJvENaaVd7wI3/wgfKvFswSIbtV+8gRkVmLSQHniUtHprPw39Fp
dKXl+Q/J8Zj8zS5IJLn+U8GOGUlQHA1Rv3I8k/Ils6YQmoLhR5YED7Jdoh/lExUr
8+aJ/J+y0rT35klfe/1/7PELu3/i+QA0XJeIrnCwZ2/V9A3QKMafE9oX0HnpXrJ8
FXxtz+VP5OxdU1FOi519Ipu+OOibp0JiznYj8Y3vkcPuNdJz57YfESIMD2buk+lo
A+hdyIwBFPG4tYYdCG7H/TvPHkw9zi0g1EK3E2LIBFMB9FX5cuby5qSqtL9x8oii
2PuHA9RaWt3hW26+lxhAkpQdSpMh0oZuPMX3UD3VVeuf4912OkdqQ/9Or1GBlAD4
ZlCupKVvNXJOl8aOtJKGo+zskhNP6cQ3uxLLYKN2m456uGpfpYJHOi4KtM2wnp2V
dVT7EctodhdMi8qebVptxfLCMVJNzg1IzsmgEpI2LlykH2TCqURrTElJB04smk5A
sOQaNeohyhyCKvwEu8sha2ukwvERRzuFwuYEyWkWLGD15NAH+wUEt49ymRxIMLya
+jUjCnxPAzaFZpQ6LlshPna+mDl+l/dDn11AqDnaUBmunRZ+2Vld21h7smSAXleF
ZAKo+ocTVHiEA491DPNOsTJq03MAthinwBLtqDa7mstGlqZY+sVXBoT9leV4zz1v
ozDLYING/ce4+nPCLXWYWj4duVxuMgKlKYyafuy0/RtZlunLaTiuqyq4v5LscApZ
egfz/5w4DYl+s47PP3qxdHF1On33SyLl8Uen5LHfTzS/4jWbPU6rLt5ACBTlURhK
zp1ofMY6dbbh/8AlYsDB3IxdOmWE+RM/RJFUYGcO6Tdhb13CG7ZfOqILA7n6tcmZ
oYQezIb0pVs8Y/K/I9nVKXSDfAyHR21b4MQsxDiKj6UhDUngXwzh0Hp3sHHIa6hK
jYzwT+dQd97yZlTcShFrsS1fvxSap2XHVrJF2+7/+R+759T5QhTvp6i+1tdqHydP
YHU+DHw/1rXy3J8Z47Ctx77W03i4sr6yAlJ07L1yqVRf3CnqFEKViWp1RiIlkQwv
nZVe0QB4jbMu9uFFtysp/uWm3/jQPU+a6t6yO85iynOD0RDhXnkzYPMk4F0jirKg
p+qhDiNnCH41/fJ8zHrxC/sOybdNivHiuE0GllM3gVF6/2lG22A7jYS3IPcrfoX3
GBpoclbV3fkWYBOeNY6cgNAadTHu/G+kSucy2WKrgCoSZbU5/rpOh+EEZIjL/qjC
o5Esm0BtwfOYiigQOpnJldiXyTKhHmMhcR5z2Lu61HoJ96Q0Q8/sr/epHc86qr2N
97pq1Jdd4BBg2FNM/+LHZ/s4WoTHEPbxCsXLBochyShzCkVECUw6YaRC68pZ4SDa
JJ/oWwnwK7ykmbXP0TVCL1pfuf8nXJUn9b744fBk4R1q7ZjAZXl3rh2KuWItkCLV
5WeQ3tBLisrd04M9t2rllpti0midn6ZhOypJfE90p3jH1Ax1gDq+C2QN5KCliHuc
jan3RTnesbuJyeK39djfGHfPtZPIZs7dA3YDVnbxzIZDuid/A/4IS4bg7+cl+c2i
hr+h4KTeFHgi3vic/WzPE4S77ysODmAc+9tBZfPCzkf9PhUWS78ekU4wZ4jSZqDw
3935MEY8PIliE1YrEoWsO9RAjhY7hzvaNT40qKFxq/GPdOuUKIasSqhSE0ieY1dU
A/mgFNP5UvhlLYnWHNYefr/tARSTGIgJik3D3Ug8/mixFgQDmvO0sRy6GkDzrE9j
KL4Td515Xvs/gTLEx1R6m843HT027zRdAVR37Ya5SvPxyXRPGVZjlMq9/o+lEozq
xsGAWSsS4iuF9SJGmHvQv7TYwjjjv3CWCgimz0Vnwbu+JthAxt3GFrZzMYJzNZjV
k4mOJEM3FnWeUcnmLUwgOdGc29l9JqpF1UYl2bRFPN717ROU1t3bN6Qpiw/uZmKn
vK/Evp2whTUqJAHqn64dyFSdqXGLLg6MAveoGn+OJeMCx+HpywJFHJiLyAI0suUh
AdOVJdA3kBjo4srmhP1dwCRkRwuY7QFXq6iitqlD4ssxnI2b4amFqFfXMpjQjRZT
VE4rdukrt/RkxZCpNIsCaAsAI1x9bUCZ/QR1DHTHg0NZZ1E+aeTvrXCEEPjz/TO3
V1IaFhAYb5ntI/C0ZKJP3k/vTx9fSOE0hztzfelHKRQiAQugOSRbDRs75AGx12jh
WEiqMYqPi6Wank/71UCukINpQs0ZSxHYQXrxDaRcGxZlk6OX1XK53lpE9WVrwwYL
rjZli+FniZExI8mBi/L7Jom6p7H2FO8e7ENfknkVPzp2MYPkbeHww45+KMZ/fZ+Y
AnjSZ5iVn3PRDURx1OH94bNIlpx/xqJFvmPGqYQOEibgeYDCyeNSGjY1g6UWNiGz
GF1KM+1F1LPmN8qr3kmsgtXtxVYwl8+iJd6dE0vJJ/5l9Tbv9JNVGGqvDjFq3wY/
q8DRfW4LX49yrsp1eW0PdrY0/pXbYq618R+NYPHnrR9FiYe6YW/OzqycwpgCxNv1
Ky3XeCxdNzI1yx0PYgpmsReM/xNyvehIxaY01ZTtLHXSpbIXlEkVW5RiAqWAACS/
uQ906p9B0qi4LS/7QXlnCE/SYhfB/dxNv2zUYsGnkLvoWu6zcmU/8M/NglRK6o12
2JsPiWxqkUQUGIrT68/fhsz/GwAHWAICQg4YRzspnSjP462xPE2eCknsvwfmq/aS
/xK+g7RYQbCI1dVaLDFtKMrjIfPpih2NQFa+MIZr0z8BvyTT1D8VS/hgEoWAUnCP
jFRp05oqYDSXNYmb+HYvuVbefhLHU2bBc8E4zMbj05RGmYuvFFPHwPFdquWqMrbX
8WByloz4XcVYptfg+p/oJ/3cPIHqlRhjTg77IcuWuSw7HzfamiWyGqB/N6Clg5w0
1GXBf6ImVUL0V+XpGLbPMrIQGxpzDrO8UgZu+x6ADDAmACTio5R0c6HSVkI9UIwP
aZscMaCcA2to7H+kZ/X0zHmizdaSmU3agwN24ia9wj5iU8niywmQ5DZqaQRKztTM
a6qmvkwszhLrHWAU3iChVtnxInmcZsdCgI3LJGsfrM8g/hL1AnXUbz/J3TQIr+jf
qRv1W/WfIUoeuNMbrq2jzKOT1G0o+4jDV1iZEmjqapunEwPddO0zSX1kWLRnEoIn
8/sZPwG3eJXj+zMlJGlrMtducxdqi/qxmmtvJRLNhmspRaW+G7vKaiYoo6X+xp/w
2Ke1pSw06PFTfDKftAoHWpKYNJmYQJnM/k2z97tWtyuDFxi787KBaP2ctLTf+0wp
kRDVqbaOKloufytb/GobT8yDfvI3i8Zc5FUf2KHfx4uT9dejZY4yg+1ViYPRtvrF
XtDikaEjGVU3CJi/D/rQ9hnExWnpztPWpW+MJTdw5xjiMnkFI1IsoH65L2ENbzXu
FxggcEiw5hWPXyvVsRCkwDDIEn8mT24/0opQpYCXdrvfoPWnVyYmg82Y/iYJ01Jr
x0GBg39JRL4Xq2ggVEsLft9+s3V66nSiD8HWdHy42k155uYBcwFdAuG0W9Nb6KTj
1+Y7SoKTnvZPwyPU2XqLoYYFsYSEScAmi8jtdHxqdR7iOvgtTwOM8SSdiUY31Tnx
1lDRikzZZUTKI0JD4mU1yWk4wNBVbjH0zD7KQUYI56/ME5v0rBuUHFNcgmC8LFmU
jpk0UsAtZQutCuMLTuSDa6rreevuFnZYtyTMWWKRMiu8gg9n9zHxGn0PfLxluLQ7
JDmOKj+QIodqqYz7mm6BriKWZw+AlzHE/VxgYTb0gvS2v4257htYeFgO7MPLbr/S
g7nLKF2X+wBgZQ0/QvzWSNatgnCxsNw/ZDpeU5T/jJiflYjgYU56VKbmQPVwY550
pf41jjVXSCeGXdR8ELMaIz0YmaXt9LLR1sIpACiUNI9Q+8NlgugQ4s7LEIPoCVNW
FrJwL6w5TvJxvSyIXfkpQ9Eg7WbwTEjX3emPEitjJao9HokdA66CL2NpST5O2KRN
9gmymlWofVeIdyBJ+eBKOkhS7SdAU4IDIZfzSauus2DWFKFOwuxOOYEcxx0bh+9d
ZlCwVimPiiP3jwSxkyvpvzEQI3toOjIBTXr+JiewXD6VjAimXXqbS+/zO+4bB6Bc
S3m/qTt4dNsDmakLsxqzN0c+TQx5mrhnv4xf8ITGH3zBc3bpo5fqiHtH4E0FTzt8
mcpGqMkZUUjAD0UWdvs44zzYlphDqYJiQ78cCke3Jxr458P+1+JSMFC6r3gQ2Qqh
l6SP709h51DNF1gVV3/icVEGTaPNIj0N/WP9If/Ngpn7Qy6fKo3eAmslbByKVav5
ccaXklblECANYjP6hyiVco4m/Uu1SZ4vlNAcgSbMvGR66x5zE4SPEj4XRqNubIYx
tgTGbeqiL/EBCPmrNfQe5ugnF6FFRL8XWtDS1FBqUsfiybTFqKngSvRf9XZk5tj4
Iejz8hhV1fOZ6sTb72D2vGxjhnaHTwNXfXBA9CT9AlxU7bRHd8qadHRpRLRWmtTp
9mAylej9S2zCll5ufz6tmG136yIsqNTVCcQmYHzg4Qod8mAgWG6s//gX3X9ZyprU
gQ9ECaUGWvTxl4g4UswxmWdikbOA3J+TN6d0KtdFRhkSEn4Y6U0O2EuOZBIoV/y0
5TYSzslz7giHwW1EwkNVkbEHiqasFv1XJpS+qUcQXPK1o+ewgP7EYFrGtlWmctDp
nAbQfC+rs7ZiFqreNKV/KNs7QZQmpVDpPJK9oMaQn1a2F1cRZfYVawqRy/8xf1Bq
zkugeBsLayjS/mQJHu0aYr3FcNHMK8dVktCsw/tdE9C1XJlisoarVpYOTBxZX5Zv
6BIbLCZMTgdszQZbuCM/wRF2VF27AaeTUfi1hdHRXU/3Hh4MNY1FKh0XFVqHsxz+
1od0ubxWPQEHyjpG+yl5pErI+hbNI84hhKQduL97yJGKkKP5sZoavF7HLmpbQqsJ
2C+R65DOzdKPjNsVqa82oB+vo6+ABxphUb8tCv5fFxJbycnhgnN5GJgXLwy397Au
B9acy30gNH0NrcYPxoyxeWBjTv8R5c4DKkHqoAsOZVSvR9M8YaK3K7O2HEVnmd6b
4NfMe3I99M8z6mofugosicMr1XZL76VtQti4dwtFPBnim3DsmZufd6IhywM1CBel
rwUPJswC3UdK5eEIykrC1Nhw8SCDe+rxBxqMTkNL1b36j0T/FzA4C1qhSOTSXM+z
4hjP7TJpw+Jp0q8XMAOKYlk8ZUMrszOJ4yL0IXW6tRbdhukeGEQ3AGCS1MfYFzwr
d8n9AWEyHnfBETRwDTFVpJiKperaVFkzADpJvLXmf3csNvfsoBMXg+9XnlrTL2GY
YyenmWTubZd1u5L3AYadlJ+2dEkT2jHg9fGe8H2a4BId8CutVz1Cxhff5qET+Tq2
0BMcS/ZWjN0Khpc7lSIEMiL8kAGNMs+/smxx7ReUgBXPGuCiI9Zt8MFS7t3k6DKi
pD0KcpHwO+opZWxtBfFCH3KQsVEmzhxS4IbKWOKT9JRKA9Y6FGDJQ6swoVMJMD0m
hfSIIAlKhtBNzV+kWYPzLJ6eNP2Q6gaTSS6ASmAzN7xHg22JpcdPLbXVxKGmymPi
1e6LANrLDBounADVOeEd0708a79JBIhmtMv9jO1etFDtdSI9sP7shP6Xfwc910HY
ipXy2+3iKWA7L+m8lOknmrYE/qv2UebqrvKHLkM+MSkVTKO5dI41ibabSq0u/3Mr
wU/Xz2s2H6KAzRo1E31ftNFkaKM34KOxKHWkX7+nzwJ5jjtcZte6+qMNFkLlPPAF
nqfnU4+tTMYYz1EfS717amB1/lK7SO3yRsHw0ofiZn+helIJo60waQP6xuXHC5Al
lPhaTR6/lULLlZZffOCEMiBBNTEyp2qXj7WsusxwS6cz1V24k5/6J4axXzWlwNGi
5Xe7dgRFFH/JAKj04MAn2cNF5DlJw50JrbXEmMzcHasL87budCd0KE4Qppl78e1a
na1CuJPXLFzAcOafbM8biPj0Ixl4geyb3eCbjzL3U7Q4vEs7D7GzrIaUMset2c30
JvZvL6V/y+DMOGVLi5u5hfx65NN0/OyCz1eXLHxiE1WpSHbtW0sDyHhdyejK4XhT
YwVfLqCB6gFahX06pQUF5dhLsX0X3rQN1Qbl9tLt0mO9Vxqi1SV6ca6f090wQJZZ
/cgc1k/XmRWPdHncHnvidvPyFfU8Kvq5GNEn3tenLBwuwevdelXK/Ap8hUUSFka7
h9yWbix3WVdjGdYBjZWURAeikz3kPTGvs8a2/kYFzmn+YZ9WS7hV9f7mnFcVyf5L
dPu6XpE2Dm/NM9BirrpTBIR4CBv0UjWgdGxSrnPUjqEzCL8DYc0cYKulBoShcb9X
IxlgdmGpOoQnjI4qEeOjNBtVyn/7rX8l7XxFcO9kmOYDNicRnYCTXOR3KYB0O1lR
5+DfoqPDt9GKk2F7q+us/V15ZnFBoRbl/jmdZB1wgaG8ZzCENkjF4w3ot1mECSY1
GYZZZEW5EMfSVAjwNA7PoMCXX06qXiHnNSNfxuRuJoChYGe/Xyrh/K91DSpZu5D+
K/NubnnAs5aDeSVx7n5yv5PbgXL4PluFK4BmFYD0axyCEsT9HUF+hO4v06IwSwQX
QymJQx8R9jxbBuHzYmjRgMbzRrX8XB9TudKZYu/xrNCeO04I4nBV0C+evu/ktIdH
IaGqjpPoecYSldT0TfX/OL4pW236x3SKrfEtF6I5qKrTPOuhFDODkbqLgsF8ot3A
tYD3EM4ZOZaKxNDi5iI40CJgAb8cuQjq7hvP0AI5gETNpgT5eecPLBUdM8Qje9BC
bhnIUraqdp/tF5PrDyRrOxB03MgcNHgUmpjOPynI5uuN64E36I5AVXS0pU2VfyPP
KMuzMUhdKxuom8f2nlpYWZrsa5PP9jgGnCa9TD1rK9q3prRj0enp+oWtZwhK/Iw4
F8uE/nt8m+LR9OJ1K3bxqD1oD7CjxYbYZRQj9dzsdZNQCx0o4I5ESb0Ivd/69DGe
Ch7lkvLVN0oXI15/CL+0xSFzObHihKrf5dvL0t70Oc4PmsQi+YOlPAluSIRpLPnR
2EYkRjB+xKTm5lmV/WevpHn/Zfee/8uQcxo/jr3qHlq8BJXJMeoODczyYASOhbgQ
35svR4NSMRo/XzOZOnLU/SZs4qk47je7c3/nT//51yLL5+jZCtJDFCwDaPlzhwl1
uQI1V5yAUjUkZxOAkMge72MpNtGWkIjzpQwRylYOUxdWqOYeOxt1JzPfoXiFYr6Y
rBP0R0TMtcZQPcnteJ2qxOrYM2zVA4LrRZ7NFx8dK8WnZ0/nrrNSsPJQs2x3ixMt
HSDp6M46/0l2qix3kjSeyipqQdW10A00q5MB5PrYQwJuofgxwA8JxsNU9CKxD8Mj
+YhUmfgz6OAfA23b5f0v+OfVu3TYKJjSF1EGUKnAbxibosaky3w0SKGvGqMRWZo7
RbO/ltp9ah7g9gbyWjHr4ExPjS7Pn3udBoeBKZA65FuqAm/eT5E13y/rhqncQqpQ
vZwK+aYPD5Wl1trgx7SJiswTCv46XERRX2suoKoZEPXktYUlY8dLTV2ZnHMT7sqJ
PTcEi4KZeKgVsOWXNPgXvZ+6iPBYlSGSRGKYae4/0wgcD+nrnfWGC+F0crZ5yEub
MKdKE0YbrGaGwwU6EjwY4MRiWzpHBldTApknjb9oo8k9R5xxgTQIgO2u9zwKbdDF
rRrwhJZvEVNDSKsUZ3kwcV4l5AtxhdP61cS0b8B2NFAzlUUnhgMDsr78rneeuc1q
e/ge7eJH/jt1qsCiqC4tF4f5TPUNEYR8t+33a4sv8U/1yg3a8J8NdBVcvZFmnSZu
xlEqaru5eVaEG9cmbNUdq967T8Ntc3J2sBRVKR9iOmGkY1g0FhBKZ3lBXSWV50kI
XB1u3PX0cvl8gU2Ygjub9ZKO6u/OnMghUIqg9h6kwJToJrv1XDrtja0l1aMPaO9J
/0OSDMKniG5efJBJCoJxFj3bF8MpbB1tl9wYCqERn5unupgO7pfgXEUeJ4qO53jx
HEsXxcadqF3jRY9IxA3Eel2CAMgdv/vfLsYg7KX61aylITZ4lj2WeXX6HdEE4YMK
Rjq1I5rtzVovaR6A5I9nu7PNRRDSfJY3OeDm71mXHoUaqCx7kwJj0AwfOUdo5Awe
iYEBHeridcnyAbhnSLI1kZ0qVrt7FwXvGhM3CBMgW0Cb7wZevzaJeJEjYy4pxLvr
F/V87Z3r/dFJq5yyecCPKosQLLtEIXfNK+DcBfA0J2nrsAoLHSx/TDj3upRfaVVs
UU+1FynwuZwv7LQpcD16hVAoHq/5BeeRDW0Xq1W1O2gRjY/Zw5xM/kyhSIKEIqCW
d12H4iSL3dedyFg73oijrC6tsrFvQzk5oqqrJ+jdVBOsiLEFhYY4TDH7N/6e6zBL
ce5Oez64oaXNlB3NHgPIfSOikFT6hC1ugJ/GeGkI11yqLeb+C5Bjpwt6KzpqSuJj
w+r/xSFhye6ila62PPljwyelsSHUHgpEKnQKi9UZtum5t118zG5rkdyfxekCCV/0
va2atYYE/KQoCzZwJgRkGXT/9b4rqKfp28GQKLfkjNFor7lEWKkpJxnp3rX0fMac
ysrm5KeVzmllB1LXqKHbLTxqWJwAOQJMvFx92iNN76TIvCw1r7vid9rMx9hAfN7i
DIB7FNQ1bAgTUiSfbJzx/VLszVJ7p6+zgZFMzWvRjhCxQNiBhaTInFUkJ9iAi/0H
x/zeN9kyr/kCX1l/Er27VDuatfGKiYnJjOxQEnGuRVHyuWNws6rPrkONR9Kd19bW
hMAhWaWR9i/JvgPknoI6onURK6qDqpUyNZlEhYGuQ0joVYhwza0mxbS/6jNZwJMh
K/GdvgQbd7IwRbbW3FWGA0uhX2B21SZsbEAY/TBB4/yA9vg8lALOnCHQtwRhm3Yf
pjZNuLOt++cqmcTJo3HrTOtkrYP52T44pzSJOVIZb3eBxprotPTYm/RilUL/7V96
UgIXEb9jSwi5UoRMJwV+ZkS2EsIJFv73PFOgX8zOZDaTWm/zfJJWS8BHlUPVTgTX
Tdf/dA9Q80LRIu6LnXFJzaiwtCWM/SE7a9euJJco7YuFfsVn9YMkVv/QTl4yxuod
kQVZDf9nsIWAxzB9vaHAIDLzZB/Wk134u6DYtDjKS5S7wNPwCA0fO5qwcODc626w
VbEv2H8wOl4dEUWPvN9Rt1BTWL6OKAr/vvJ6tyhcLErV8sj3m5bE6X/40HV5Z5m4
ceZI77vrpqShB3HBOj9i6cDn3QGPR1YHkhBxz7ZxAFSqM1JX8/o4S2kq2WyvvKww
OJm2crLxfICyTj/wubRdCFd/2adL6XIGCdkh8a0ALxGUxrqNpzup7vb8XHxgp7Fn
vsVJV/NAHwGSW8Xpz3pTLHOPJqXniNejCxKolYh4AAodfQ5iqdEmy/zzuzTmvgep
Efq/rdElvbChhHqhCekA9A+Bljv6Jg+SY+3sZaGvBRxJPVa80sBbDey7ixqiD2E8
2NRyltEI9fod3lvXF23NTiP6qAzVj7mniMQibNgSJvAS7ZND99oUqhxHbQGJZdnI
k11AyytdUW4rAAjMcqtw3nAxe35QHI4um76u1SrxNO7+qH+7vs0hR00Pw+Q2sUYH
4Mk0REkOLkUStk/71BLOAauGhg1lx7IB9p0JESjueXWm0RcPZdxEeSsl0voNvdM6
j6QL9LLgDhZX87WuchH+dkDvJsvL/Wh9M1XGpKr0BXSSPdRk0houKF/JXaLbGX1T
Xs8gnJQJ6pcbWbX0F6antnJcD99S5OEMuxx2T+2Pq9pc4MhXg5Ra1qbklKR5pur1
XMt4HPN9uuY8e1G8Z4FwpvlKGhY1E9evrRHVXi+Kuuga8v82GLemjtHJy/lC+rs+
6aBZcF5QnfzDooX66uv2zpql8PwYdxeDyy0wpFcr6DC2X1SNWBjObcy/6pV+KDJ6
WscUMyGnk64vFUOXM6dTFOfDFTLFwIr6y0wH2xVQoiyCp1/ZxQBpMT3gX1iWlzLZ
2bSHaGo1Bhfz/4QrTRKiqLt2BSj8AzQwzAp+yoXQvGdYvTY25DcjM52xQXlP9IbG
Cxd7+ovr1IV0Ga/pS1tvJ1QM6BvvEm/SS4OwO851JJvU73dXIvNrS6H6EUyMONAL
iMqXzDzRV198r0DuPkuThEj/u0AqPxf0txIdiWxFJXNgZ3iu5cFzcMJbDLPK66PJ
RDU2kHgQCexRCCzfvpvNkoY7xD/sBN9NRusdmbc65+aUXsAP1UulzquptEIdswuY
ZULclemW8B7Ll56s8zjAJKchyDcd6fK7uVLOa5u/E0BjEAHjmxNrKV0QVLV3zVnR
tuDCb+n2cXfLI94HfDBZHcDlOkjfKFdkxVhS/lypn10CYqcAOMsNXagbo2OnpkJK
OEwQj4LjDNp5MobvAuZK7dD/civp3wK5mQCN5m+dLik9O7ZRZ+XtYgc4vgV+wfCB
RHvcwSd26iJqYRAYLDM6RmGUvmqbGRUBR228Mxqv8q91W9r2/Mx8XCMmU9M4atbS
gzSpkeOish5FxjMhdtW+WuheqJk9Bj+MaXwkCB03tFYrls38OSe1aZ0dMsMwfOjl
lV1hW5CwkgpiKOv3NpmEE13nqxGMndUz1i0kr1EuseaW1GSUKa1cMqIoVBEn5tr1
8LTxxfbXEfmMHCloQbnvPaJRo0l4oetXq/Zz3F4tbrULAe0yEKSE4mDyvkLI8Ab8
NUrNpX8DA/VkyxJqfoV37Qyn7a2/+UY8YAeVo9L4i8NiQwwcyXDiVpXP9BVauT6i
bZ9rGNYvchVRh62BvZ9cAOr4w6gkscbqERxWoGYXp8v2rznSPlimXyLhO3hERgVV
OSB/IqXKGVrMtY49f05znW7qfK0MK9Z++EJ3pHqi08T5tBW1X1haDG8VC8rrPX2v
JlfefqT/qNGDSSLxPVHwHHIw1DZ6pVhV1C20WkOcvP9bV0Bo9R9VxeshmQplel2O
M4K6+4/+4U3S4F0I6qIBGz0z0WZ6BhhQVukVmxj1YZpAJ/8plpQpAlP8iudR2UHv
XlUlA021FHHZJW7LGb44GMRzabBQPF3dMabB5dVl3F//sQvsYbZtBWMP2hAmziUY
YhB/BkskEx2SgMlenU5LvIlNwvAr5QsLazWNBNXTEFEeKQB7cqOfIfi6i0WE0BQg
Qq+x/zrvH51iau4Ev7CJ+FGX9nUIKJbkg0wqVBoSb1FKCw+yqnhXieBeuAhwFghy
VHgpOvG1eeO4w3uA79a7+oSKutQMDpyPV6iExo4I6wS6qlOrrn3HOZ4cq0bW/B0/
dbb8ID9+0auPTdvIYuI6Y8zS5jCvUkCTYk2YVaAxr1cCFz8fcZKQMUZr8EOILdPD
aslbSAtqma0csEE4eJKwfj7T4pa8lVkdA7L6ruAMXnDQJ7/bisMLoOv7XOI1NAE9
i9p6BnxR2c5lazVt42pAyYFzPJ5/PBjqbgBSkR5AI3yRptPIJBmES8Qxab068qeW
8CHh1oNQDj5roLBuoBR+UafivBBZSI/MXfRIgbSuCBqj2kRUrw8Vr9psXyHKTlkg
nU1wQQyZcjcBlfLca1ZVXnA5KJHeTho+GQH49LikkJN8DXhcy28YhhdFLzlh+J3V
nQa00qLf7/HoNXQP5rbI4DynJoH8kznOBLo3Np7bdfnk/oQkeJTcWOHgXRonmEFY
J9S/MfGF47qOTLylSk3vvyMpJ8MLBZ3u2b9Edt4frRAR0BciFvAssfchD2Go5bif
ogBeehnWU+LAJQUYz+erSUS8uvtjxPsgB5ZUUourYRv9df2HY45lIuqFryYupwi2
QOWKKRjxcy+5a//NCrkWyk9wDmvp+pKDq0lqKs0AUl40goRt5wYSZJOof3gbSgxa
tHxbDfV15neHSjU00p1pYzP10/WkyH+EmonG5t0oyIWE54CxBsKsAnLUrH05db/9
7/WGIKCuspV9jG07Fjjf69vxMk5k8y7g+YtzOSSarr0AdEPsq1CBtF/QaSlrV99Q
nRdEZxbigsnajEBAiXllOxlGtnwUz47XvmFA7O+JsEcih4ItsBmXKSKXuuHZF2mY
7jSrJVr/LgfuQiLYuRJv41VCLeThD6EBLjjtnh/K1jAB4TnYb7M0afaMRdSK2QzU
gtB2yUIhVEX2628Qn2ydJmUJ2UbEwZ46SMIc4/U1ftwa4T6tArLTUErgFtqABx1K
me+Lx90DyEueCJ+0YIQIauwz6C2/4E4fF0Xqt5slQuNOiiNColOI9tK8cZ7tpP4S
1/KnNLsl5dvweiYZJa5HceX4T432ZW+kuSWzMkNWmLJOE235kw4qefMeowDwwMHo
pdc5cpLlM7puMzUrMfzBsj4gvTm8KeMa/nfuJMTXRHOjMwcqDwPTd9L79918YF1A
Tq4QQ6zSlDbKKbk1BZgI2m9Gg9K6k94x+aaMPWVgTwtbCoKB3TgPSybNj8o06wXU
G2EoH4qJP4wMbKScxm5S8ahGPgpMF5j4oyX3lLigAHEIkH0mFjrjziRqv8LM5/Vb
OAGUt9SxDwsLwsA0qOgNXEvrV4dwRtEo2A/DnMSwFn8rAOwZY/JiBq3VU5LwYwUf
N3+y2splhhdAdY9hoc9yxPRohixnC4bSvgPsiF8KIgkBLw48lL+cUTZbxrRyHRLc
c1gZLcpCKvjRD0lLld8sPX7boha78gxhKKvxIbHxzXG8o4qwoAw4KjD3+OT8qJjE
KmSXg+A8bI0afCLxwpXdMryv5xhfyUSiGVsoKvraISjkKfY/CkNtXlv6ejNZmngP
V0KiwtAhV2AISUvQJVHbytfEQGlOwQkL/2WTivSGqO9GhBrPI9UCKuxpv5Ql+SaI
YtGxZSiLfmYhdGwhuYqPHk4cEzZGuODYxk7SUSq/9gN248EnGn3RrHchGobaRmgL
nZgh6C1MYqc/5GyMvbIvAtw+fLobF0YZ/3zayX9w52qKYv44dltRySRlVgXbjP8N
gz5VDOHPlaX0+LOs6Vc95FlS0ggtWVb0iMN5nFFm2o8Mi1FXSI1FAqA7grdMoUrt
tyPEgr587jQGqvv1GFvPiebvJy2yt4vKogb7umEYhPiEBUuKzqZ7aQHzEWB5nbE2
0rJZEhdxXpk4n1aL4avGiI94U+tJJ+L5uz5ciVe1fB1t6tIJdvmrp96+hD7rjn90
PJ7xPiIX4GGZdCI6TS4sEvu+cLE4HnYBiN1p9t9agM5Q+mKsFazGuJk1QP2u+/BX
/LcsKkuWWuykTC8X687GQoCThrq+SnaYcAa+Eo2vq4oPdeLAbaN/FisGyaPEw2pH
inUEb8c/vZ8SdGVOF4I+6ABzz6T8Ufb9p8OGmtXmYU8h6cs2ZNDzvEqqQqANoYF2
GzIGjZkcVoTXZBBignBQPj8MN6bo9dZh/3ZucVS1hwmxv2tcw2hfp4ObZmVEhDWX
XgbUMANz+DEv6r7RwZeTa7MWVdNf7CpOWhZol+FAUirbIVt4RZ2zz3RtLVqA5h5t
N/VOYtJBFOcX34R15PFjZ1ZsAIGXCoif3wtDnrVVeLahFoVZQiSgpIC5mVmcGrG2
KOXG8ADoGOzNYqvgaF52PmnY7TlEsI7hy3rRYpJUH/3hMhiNFIclrVl5UgiObPA2
APqRVuoKTiZdl6PwQkwMyMIHB2YoZjJQJ7sHcwoGzumYNyOL7pCJiJSMnOw7z98Q
yxCI3Niy+E5ZFV6RtbXaJjYnSzcQaEkTiPy8GzpPF/SVyuAqyWF4VTEkjudDTXoy
uuPnw9D6pwPmsong15M2WrBlvc/Sk0p9PoftKDzBWOhhxCl6D4+pKhxMv6viCDGv
xCyJ6kTFrKU+zJGGiysmP0r2SzqtAvP0Zk7yN3fQToC9ANWW7Voo16P2XXZiHAWy
SSPLNAww6jMislwdqFPLl+g9wYuSeOBkUyrIgLAanWk3ZqvaFNZmjcVKK4WweX7h
UW1Xt9NIxRbKmcmhC224to6vyq7i3Gl7E6sCKeg62p9p6B+hIfVhfhk5pZ4U+Hd2
3uylWdZqvnEuzxVk//kijRWBobd4JteVAE0Y5R8Lt2sV+UfFVp7Hv9IOxIgmOhbm
tincQXwd1gROE3AxCJKCUS3oWvlM8JIqA6WSTQMQ5n2u3Xnfm/icafgWh0CGcxYF
smJIV4LSU0Ly29xa0rDhs80xVE+5WxuzQniEwUTb8N6FB4wYQIt3/x5TBq4WySXf
w/ok3qTUoRBOxpER0btQ1iX4ELgmc2t/rEiSsly57kbFkuBOrQrd8Kkm3lWzh6nE
Y4nLpEpyKVlo15iUEgcmVEINQyk+pnKeOnSa3Ai/RuV5kx/1yQIHsZgY9A21Yynk
lMzh8jq2J8jX9D4sqrd1O0Pgfojgz2pbKIwgEQCI43yYqK6zP/6ytRQ0oNZBzA+6
s+MLxBUsvRfZWIy4HiF7NvhSK/WTFvu4MPA0zJUlSsSzm+xjL2TNyUE0Bou12oGn
fOEG6pL8hjdgAaECxYVSOrDVLCne9teh2oQzf8mkTbM0UeWxj8xhYcKi1uEDzgRo
boIEDe/sPG7kJcFVr/JuEnfvbTSx2RM73jWDy+acHK/j+f6PDW0I4kseGLKSJe9I
ibaGbZjlnxqCj7+t5WRBvZlDTvQ12aQQ8wPXCvXAPpKrgAnutTIBTGB7dI6Bankl
ZnLmi0epTdnAwshts04Hi+uDzjwJ9y0jc6i33lsjNteEThwd85scp1bt0ZirsTG4
xNXOd6EnPGucRFbOdu5yXasJbEUbpPMYcnhvGQlBsIEBKoJz3Cn9JvKdUB/owNKy
cucfTbqZXgXFuFnId9zopxHxqPzirN7lQCEbRTHaYW1F+pdmBUQEWVSJYGYcbJ8u
Dljz0JiY7MC4cihia8MqrW4IpYnhfp2AfmtK0v95YW/ORXbyy6diPkyFuYiDtDIi
zOPjfpLTMYvT2PSKh9vNoq9hgUGtZVxMVMtiDmGJSeMY1UFEE+xv27H12KlSyyJN
c5R7i8DYuNBv34E7uMmYh87cvxDQ4IdlN+htr91oaPqHkigobe9sLY2+OBngDeGI
qSppri7VIVejc/FT70CkSB/SFnSoSg/ZKQZb2GNRgOEHep5PdhpdoKM3QmlXMGLB
GG9ORJhb7Ode7hhQqCqy6qdPJv4sq+6DZVk2f6pU0ovfiWd6sKoXEeNDjvbirNxZ
uwf4PIqTlrsTsiHiB7dHVdrmg2CR7gO8XUCZgWZ3jik2cOCvz5H5Ho0p4QnGy5NX
Sk9E/Dtnxx8/Ze4Jd4ALDiccM35i6fTKeAc6zwYM9mmCzQ2Qn0CuvOlUW+OteAnj
GkLFUveRLzB/EiqCEWQRLukV0o9RCG23XvV5LeJFj7JDzyip5URmkligMwkkuK1b
OOSjd1DKSWqDqivOuKcR40J5+D0Na/F1XawSkda5Qh6hpiGdTa/+BIO7Nbo9Ai6N
H1TMd8ggn5Ktx3i7sAoCgJ7F3RQH8Sa9AtVQ3z+KCB0J0HW6vx5lOp/WW4Xx7L4J
f2rhpXM+eG8NWZffnByZq79h9uaKxDiEmWeUr7haMU0++3ARgUDJodCgf9ZT7IVs
ElK3fm/XGJowiFlabJxF0wLCmJHVlDKWfkifiZXKJB2o1IVH+YwkRONu9L9wS9DA
8NNFz2UNz2o2H1KkTX/w9nv6t3HtZP064vwZtptGAe3V3VsuFsBoREg9fWJOMGmQ
VT/iPdDbwOAxfxnVqhLVi/y61/Sq/kHyv04IME9CzF0sBtxL05wjTKi2Nw8W17bg
9JqjOL/vVlN34x4fnXyaC6sPldyrBTZBuCFuRQCh/N4xQni6Na1HDOHocJ8k2Mfg
sth0Pk37Yjw5p5lJSlkOKfpTGlU+34iYnnaWagnylL4KYk2ryXMzElU7Gp12TSvA
1FIo7wiubM8HU6fZNeQ8gdBpkIHNwYJGrtjPV+bEdkrKiatltEXRoJBR/2PTw6JI
Ze6HMJ+nKy8liW6czGGlmK/VH5se/KnAX5xzHI1PlvJl/6USJyyVf750u4AglRbP
2UCn50T+Co6/1LCGEj7gxnB41thb1wTOyu0A2EvxOxbt4w41vqzYPlC4Bcj04jdL
AypB89A1VvCNg6l/BHaYdVVO/tfCzAgtcR5ZJcgqgewYe8NxebhI6qWigkOMQahe
woIZwtCsyJrn3L+s6snZJg8351R2tIydZIWfwKNbup/IWRNk68ZT0NxfQWv27li5
1ttsz7CYHqaX56k7Lb5qP8s5BVkR0BXcawLS9HAl+NdurH0QsL7/0Wa22cmIpoLb
XjKXEwwh2b9JZnSOWQ1NnEP7egMdqtaGWuEXfHmybXIak1TbTW3e5tTCqkP6Arz3
+u3DxhjZQNPyGQBWUnGTi6ped9CpRnVBBjSp0QFmgrW8nbwKzYFJmiAIpkTxnUb0
CU295W6IT14+yVfcwtrW4dveNjtBg9vCQbFvUIWbg7/hoqlkJLB03lcveTBYuz7Q
wXXuAAoNUFhSS9YCSEQdVpEu3EQ/OOF3rcQ7QCOxrr5MCM6dW6bHlXBcMwWEVx5Y
n2gFTqdnl/qpafGKNcETV4FT6Ts/wGqMOARtvs6FShvlc6DggL5OwbqO9jw6jUFM
0SON/3VY0O3gSCZPVuHvYFHRlZoY/Kkwv4iu94I3yzkKnuTBDXd2UU5fNVq6j+A/
6cnnRazZOSwtKKugSEhwwwrhvUmAXisPZ0stGipqS127LqYqpTdkRczYglmt/0WI
Fz6xzhSPNjxMMZcIgNbgM029TwZVMV1lRaCv+UBTEQMguS4WFaUy6zVp0QNStww/
7y4GXFSNxeZwh8IknD48eayjV717voq8B+BMsAxCb61hEcJvig5akXQ9O2G9QMFq
vdwJbZuA7Qy2N0izIQxxyO56ziboUBsl96L8wAjZsjQJZYCNQq3CpBcWgOXljZE9
mjmVOpsaXWMeEN+SnsRxNQGtqocZrbwspIN2iWWepw01HtIzaPoSieyK2fwhopN3
qI+likbMOqGqW3qIxvN0aiRrN1TWlhqdwaWcWk0mqVxXLL7yOeZAm74vWQcp7rY5
2o49l3GVoB+pI5jqys2YA9Xb8HA6lKgUhLO7Q3Nknci8324zr+aUTxvpXozCaS/N
OuRezJg9okAp67DbZCcrclE2RmuRoLwJLJ627zgCexGNp2CB9kYkcf/EMPNllOyA
vUvjNlO1s3va0UIcainsldrdzHHU8pk0dkF7WpjT7fQ0RB3Dp8HnkHG/nhNzVrW5
cjmWPfHh4RkUY5JBrrxbVFHtrkQRzR7+J/HaJ4bMqKIl2hC38LZiwK/E0pSf4Ykb
heTNIW6GIAZKoB6FkjZV83d+E8WnsDt8rFUwtT+TuyFJJsQzD6ID0SqNFOKHAI6f
EBwd+KveyAXjAFOxO30mb+IqmaE//YGYrtr98ka3Kk1OJPcA/0z9fCKO1tNwSZLY
CeJO0NkYyrYnQD2Ke/BW0/CcG0RkGA9Uw0xRtusun+j3O/vGNC+0nUfnSn2VgHLt
r3IA+4Oy1RPsN/nzjVx8TL6WTZDwjUZ+s+SnZWxbyqjBBhlCKmKFQN3S9HqNtkQe
aOmEP/AVu8gUrnzbd3YYZCooJj41LHFxf7hvu1rBS7v7vW+/U+kK2mazKzBbVtwE
GkVoJZyiC1Qgp+T0KTo7klHR1N9Lb0djjYiiNloK3dvnMFk1bEcAAZJWI9bZnAWt
w29LUyRM5X1kBHevM23RLJdnx2ZCJSrTbnQD6oxz/3xoumYVcQ9fC4k8I31gG3AT
eRlpWa5HpCR0skHWo/xCjKfB8/Utwv2FDWwdZvIy0MPR/kMl13JnTDBCOq9fdX2A
1zJEcEYAFo9XKSaaQPO4aKVZ/fQ31V1oY1meyfY+IhNFWghVg12djGU5R2NewzrY
GxJfyD5/vvCRU6cVe2P+GHgEIvpWTFqJ8hVGaI5+jOkXDxi0p5Dr5bK93gkyv3yf
JT1Ads74SAtVve+zdiuUAahqsQolvWNjjo881B2O8IIMj9Py5GKFBKiWrhWiIip/
zBpepEpTLAf5z2ePy3gFj8I1djbxiMXWYrLTqFTBnaFzRK3lOu+k4T5YDVzZ/12e
OTX0Y27vIpsDaVgqyj+HvzM/qPe2JkddftezmbR2Nh4rEj7BbvnwuHUa37kZcDlL
9SKGaswF2x2pm0DSrwuooRZp1Tm4i57+CPAXuBWm6W0ljnUY0T2W44s40jvPXk74
Jng0P9QHtzC5lsA7/Ygc/a09OTfA9bEN5WfFsio1XwISprJw+SuJpoc0v3Ist7fz
7LtgSKYlo4GQWf4CGWDciswskWBJr4AVe7JjmY0w6LnhhmQhMmmaNujGrwN8/0vb
qCRTgwR86oJRQfYKDmpR8AmUleRY1fdk2SJyG0bvBdTAozsenAS0WL00JNSnZYdN
XtVrZZw7DOhj3F42g+BYwlR2m0SW/YEpbu10ON2Rx4x9nmCzGzw++sQZ0uh3xahM
YXJpEcgEy2bd7IipIOyA74jKrBHUx8ryRZ3TeHZKnyMel+1wiltdDzsJJE8anzk/
3R2eEQONVBotguOGRG5OJC/4agZuaTbGg8dKFCn0KyhQtgu32QivvFFSzw5pNgGn
gfBzZTFLXO7XBKjmVnW3Xh8/aKIGw7s0xNr2QaFjUc1qCo8mT+I4OXwnNe1imQSy
YLQxUTzk2xjeC1a/xlNJPgp5FpHmsafwswvKOEp2iOI2U8/+jo2mG3et5wd9OUuw
nJTX1El/S4Zvt2NHD485K+jr8Ii3DbKkwc15Vyvk+Hpmby6yYznTfr1Ydciblxc0
BUsaJxSVemPdCKI2jVPV1N75fdT/a9lST//w6zYzoSRbIVZIB/cltp+g44KUiCP2
SepQrzKY63uwm2CsuCwGY4P8rAFMM+9r4KdCZUl4vEs8op7C0RhGok7pDpJ99Igp
NS1buW12mGAzsEQIKrGh+UUZCBwxlKMrHsU+h0e4H/ND2b2OSn6MrE2enW2AGIKV
amVXVqBKF6Gua1W3r36PgC3r9xZ7Cx2r2e2njVXNVYC55ybG2rZF1/BHZu3XApGS
ocMSSc8wLqArneqWpo18WiOgh/r18z94svy2HXbqN1BH4GB2Y6z3WeIOYOJ41Val
3qcT8V3VIDNf8oOXt/KqXAnPVHCt1l1+2DvximXhgmI5XwBPgzrfLgHuFyTaj5tR
Wn2ZreUutq/0RE+7ufDuXauzHOvhd5aVSmKhtzlUvFJCTcWzWECVsKh4oCuZYCUm
JaQTMyQYo/jYTQM7IBTpm2MwqsedKOF+hy6g5EO25tsEL/AZuJK00g17llp8Cb7r
XMLRVtXsFLTvlKsjIv7zXXxg5TFH5fCrIXcDL4A9yvLq0tmUM7sP5bnBNg54HN4q
o3nJp200imQvpisQ/B5jIPo4AK+z/k/taxEtRm5N3/iRDM2DKBRzbhW3KTNS0/Z7
PVjxcXv61xxP/grgHKoOyH+BgfUEokbVUAptseYbZkNPWX97UDj6hXz2NTbRR7KH
uusoo8k8wXl19Iwfb9BBr4Hs/g9CvJB87NN/S8IcxbsuGrHwOTSHxYBuyeCX5cF1
YT9SSRuEdnqlm4sFf6mKlL1yzu4RixlcgaEMYp77e1mQ1BH7b0mBqY8T18LfMPT7
7pdbCB73aoWtNYKO3CgGBImDG+mHsgk4wkQCE3pNUxGgQv6HHpqaSWFOGgImMOjZ
AcG4I9P/GL3gki5odgRpfgtNDrIA1bqFzBiJPwtcXQXVgr+KRSK2Ya5U45T0xbyP
IomP598UbuU8OZj/iaBJbAKq3Gb8T1A8iVgQsncSumIOZ9g6RFt+pXI7wr4IudQy
mWdTVCrxTpuglFJZjwYFxYO0A0dBMaMg89CsyzXK5LAbXF5qlBbH8Nf5z533zMzd
xm2diWjcRAHp8KRdpb4l4wAAaY0ZNJ1roE58jB1WxK9Go+/1ekffd2BpLlCiJtT/
4WBnsuV6XVhEUIyv/A6R0hQSn5Fpxgs9LieUVWgJHXjb/n7xaDiYFEYF4B1/9PcS
IOsx4/4+GxeuCgvjiwIrMzPpjJVplAi1hPdwAx/guWZrsYL7fzNXJkKyp9/jYG11
9sNKzt+Z6EE7JxWAbsI1e0c7zpRvscaJMvKoSvwd1sA5Tj2ljPzIJYjcT+WrBek4
AtM/RllhY01iMYEUPzSEn4Xt1Ar6ta1aObhd8lxZZcVlLCF2g584N2D+X1gElr7U
t5HJi1ytRHs78FhsEV9ULOqrVUp71IOPLZ2lGTiIzuZY35l6ZKmemViZzLzH7Eer
bTXx92En0WRZaSKHWabaP5fKO50lCKqEp2aTi7rgEDcb+VKFe/McNNXO7GnnhWpm
FnBrx4nN3L+JWWh8v5ZKME+DiuLxonJPpzGqgNhjIdgBd6MakJoh8B2ILRwJ4zG0
p40ATfIHKn7/8ENkpe3LQovMQTJqHswduB5t5f1Zle8B/YTzN+rqJ3sDaWiMDE0/
WG5hJRk7Se/s5Md0xKgUhT9kxdjSdOhz8YUl32tzC4vZq6xQGk4rg8IC2UAcjyFQ
YyLTwFJb4fwXwbcpBCDUm4D/beEUS2tlrL2xwJ8bP31+k11LnQ4gzR5ogz/eWKl0
hsE0hz0efPaaXKENH9cVkET601I9cl95gJJhRqYkSkDFake3Hc5kvwDocUoxPTCj
KgKZtD4gFITpTu3Rumt/ffZ7tz89uRgfplE0OemrNbg46VsQUJY4YLcgGgCK/6GT
QiL8m3BYUVseaUHRsaikCBs+CsdZ0EnDQECAwbWYbt7HNnJsY+jZbTqH2KqlUOfz
AGbS8rfhA1TXWUPpE+NyvwKfgw9+KBoct8BdtfXENSOv/RPuYLvQOjsPleDUAh/F
rVe2Du1nU8PsHJ6j41D/AE+uAeiHF4lzsuTiUTXOO/mGqiV/WK0xyh3MTLRHlTaQ
C5XSrBObQJZinZuVDFEr2CtEvDKh7EHuqC7iGdOnhV+dw+ruAE8bI5uaSmP4oBCm
Mo98BLHFh6Ck239C6gP2rTZtqoB/+kpH9dueGl1XGL1sssM1W8i18uFFw229gcZE
2yNMvpm2N/eNN4KNWKCyjvphlq7fHC0APTLIdE1RciWa+MagyzE1acUGt0/lZde5
gfeHB3wqT216aICKLcr/TmoQu9fv/G1Nujx9obK4yg9V6ZaACxUN+wCGh0Eq7FQm
Rmc4dFiDjANqPS1JIA+7ZqV0bKXu5TxCJ4x3ICbRslZbXu+tS60SBSMYLQzG2610
kR/wlxWYQNBcUNDt40efD0TYdK0xzSSBkEIA4ZWvhgjjdbRDXEDTGpKoPZ4t8xq+
qEbuP6FFvo7YmMSQL4OxC5HbS4mUxVxst+KV+cQWebn/TKXnAg5oe0PQpGCKh5Gi
1FBaU86aj8jlx2e2qGHiRG9ZX5ATULBA0x1kq1h+iE8/T6GKotcQGGtv6V7kOXow
3UqGd9iOaiwGDRkQSPLkSseOSKfNrOyaIjZtTseqYwbhP0EhQ1RwQfNa63Ia6jJh
eBNPg9fv5IoDp4bzUwXOwD4pV1CuMvLlUUcLEs/Erau9vNJrSeyChQ4W+1l9XQkY
+iGVjdnaLA45Wng5P3veKUGbwzXrvQik4yqngbr7OZijskM41KorVxBPmkRuUxg6
thyoM1LC/qEaq0DD5/hjzaQPD2guQ1BvJ1w2847kC2E/uCnPYBVzlkiouQwslMpF
sKUyUw3PYr95VQlSS29OgDysL+kz1i0yqfvLvgtrH4KUWMqbiwEQcgoR7TL2jV47
OzAWijhjMbhlQTk11K+jmfaJGXlMfPE78vHuz4lMKnLIuKAeVewmMzHQDBqQs518
45V9QQzzhoH2YVyzFNYpHJIDsywKMqS52LO+GozbQaTUsrE4BE2OxOPz75WxNwC5
Fgfa0Bv1j1+fXtIdU7Cnv1SwDev38u0mfc6eP6I0FIf5IWQRCF65QI+pqP3gxflt
fBQOkjgxD8ErwiwovaATfb84vTJwwyjot0kAxVCVbZTNyLObR/Yyv+w7ac3F16KT
py9esJsOC9Qmh2vEqcbhEzm6PWJDFlU0rhb6xDpiZs43Y8TfVHzgCeQU2tW+gLq9
QBIABf1eyVaML79gCJZsSU+diI89sz/fKjSEwLS+17Rb+dLNJBG7A8Q6WR+cJu2l
sMmQnQIofUR1Ns6BJF6huTi2gV++214ElONhxPcxu3C9FP2uWo7v1dSiFHXdm9vD
0STRr13LYeGWYkEF7qPpFWCblgZ3nQeJJV9SX94MXDbPo37qgXX3JuNsZ9OGIyq0
oRm8ln7Ts3L6xzPKwt+huWbb0Om9h2kzg33t9hu2y3+Ruqir77ybdN8Kc5Ppucjz
kaWk19eZdLNeEwhN5ZhSVb+vjHoN/+OGdyKK1RsS4lNslU4zaCPAF5lUMHfmyDXE
ru6DCVLSvBUk3FI08wOARanEE5Q3ilNmRHPgeKT8vHEX5s8sYalChPiv6drnTblP
Q49VxsAhnAnyrTDW1DApRpPJKnZfrQy7npP8T3BSwFUj01VX+yMkCPn09/0AT3+X
9nBsXNZULmYm4+nO8T9d7JASZP4h6lqEBoPchvWw830b5WB7sgcAjcls0o0nhYxh
Flw3sM1OM3za5eskAm2bphkUyo37t6szuHb0zK0SdPl6JZgapH25FmQSoZGhiEis
9CeLE8sN5/Rolfhqcvn3+IU2szGDPlGix48GwHXqM7BnYtykgvruLNtJBBSg8NGW
Hrhp10EbPSJIAAkbViIQR277d28vB9F6f/mDQ4tHJYUQw1/PvifCxKf7n6KEuHSp
ni3tGSpBKhobMp6lUaWMBAoDiykq3rdtOfivE3tTJ12PAX8IoGjIPRi+KMONfonp
8fjSDxbuvby2s2ZhjhP6ftP3tRfWrC6tmGnsj2BvMZQY3jWeayas0LmmBlc60c+s
5UYB4Tdjw7Kp/6di6eAlGImKZIWx7rCGu5WSHkaZe5qNE//lMJUtnnr/miSFtIfb
Z3Sn2AV2Ggc2TJ+Poxgpi39u8h58KiF1dF0Dt8iGNh+q0xDMiP/9UJvL+lOdANrE
JZKn/ckArprGnKE6++gJQ7btNSobeR/TuCdNuxbw/RtNY1QacXJlbsUaYZ5Wb3GZ
/Mt0lYfdzrKWUkcAsi84THClDl5oVgEAmPk8MuZznffX0j+mgymafO6OVMyN0Lgk
gQAdahWBOzJV5ZD8263ysNVpYNyNQab4Qz33W1x1s1m3SVtzK1NQ9ehCyrt2yiG3
GdIlDW4PKjb9aYJBG68APyLEXG0flPSRwNR56iYZU2TJK04GLM/iH2oZch6OgExQ
ppTp3y+XIWk1voLGBq5lIXuyAaziA4hesoBKiiUZObo0rpSxsP4LXm8TFGJ7w4mI
wqTgJZ2NkfNlXpSvIh2Aorelw9ehUNRHXUX4TOGZ/64eqHpnSxab/7zkxlPHo/wr
l72bEv9yT4Z/Q4KTyzqoPY7lms9T6RBouaaogrM9BQ/elz/fbm/1c+08U+dcx4cj
V03gxmhL8m+BuOsUcJ8iWeK2+hnnScYQuda5ADI8+wNv6fNpebpvCINu5hODxvG4
kln+h4sSpI/rEFs1Vsw4Tyx/bTi6k5LDvtfoPENYvaJ9CU5t4AacZUyNZyMlRIib
wWG+xZwcasELLXn8v9Z4Wk4otLlshU3u1EXXH1OC6OgcuGJypcFe3ka+ZzRbzvDF
pAUQ5Vz9GncvafL/Y9eCflAQ2Not6vhnJikPGbcGsmS1yso1dIw9wWIV/djXT9Xe
cBsHNMxwhoFFh+8QLmnM3ORXHNpSSrrb++slTzLFV2FSUu8slaVkerWpOUIBcQC1
MkEzByg7ux/Lnq/S0XYEYT3tGIMPjjXvmXfLBH5kcu5SIqHTU4hE7Tbjwli/2K+s
eWnhyN4z1XZh1XUhoHb/VqR+ZC0KNuxgzyYsLtDUYbKfyAeqWDqMkQICys1azV0Q
XoUUxIWHMAaTymlXt7UfhQ72+5vATof1SJDBzk81CsAxfdDtFRa7B39jXo5fR3M9
lxMPekk+LVl6W7rh5hv6M2P48HaX97NB05B7yTDPzhejsQvQV5l1JkzY+EVKEROz
B5uc88NPZMv3BzWAjaul45/FIpP9Y5t8OyrkCDsjiyhK/NV0O4bp30Z755t38WbQ
q3i9sKKArDTdpma7o4JNTnO+BmTahErY5bXLANR+mmMNo7tVY9keeCnRGIfoEIAZ
ouLg3HxsHnDko299hii7JAZqOrgw6HWwFktJmOwDZ6IL8WMpOuc7iev5uaZPhltQ
aOfsOc+df3ZsTzgpR+y8G+dxbKZ3eenRX9wMUsqvLl0lICf0wODFYdId2yFkj1DJ
LcmjIV0ewME/SWhZcNsIOVX6JL8Cmwo2V0lsrNIe/Idi5NlG1oVlK59/ENO3T04G
RNY+4DsUqj+/J3pJ6xBem4NUcnL4Ra9Cm2SOerFs1+teAXn0myvwa2NcgFuKYqYn
oupJUKou9LHh7A2wVlBMjVNdyFfJ3UpHeymzeg+Z+xAGecAl5XXXiWqo0mqTzWos
xuMeZrznywytz1DakpuLg22MnPdEJd0jY2IVyUSQzGzEt3pcYQ7TAVQIEMeirQj9
LR/T1ndk14wM7HUaEjfumLPUlcMMa2upN2jY/G3q91N6tQLDy2/FLYmDS1zfVmFq
RNAzkk7rMgW43tVeFPkkflpRKuEUHBayGwoAeLej5DzamtkTBk8P/BP2pheWbtRb
OofIEZ7L5QC8WWyguH/ILlb3vPY/iLs18skJqlx3s0N1+9ueYd4ncZYbFrp1iThj
V6o7rTZoTgdOufJlhtSXdUSByfZzDnuna70f0JbW2/cBje0koksPf2PPW8gwpOpc
xN8v1pfJWFkl/Lbe2lJmoQtT9nJu3wtQ/H/vok6uHm4iVEPP//YtWwM5zPnK7DpR
zChyINPH/h6oSsSuQDei/9dYZi8LhfmFC5eSNQ/rxxc0YzLzQ1tuY6j1fNB2z/te
B5g8PSw5urZYCsSRTjbYT1DPKVeOxXNNvN3w3SDYu22gxdjjQQBySfNRBe/jEDVa
L4trZG5fKJz/HLw7qHAIdbJCLYvjuhIqGCpukZ3lVSt9P8pGa+695Ku49YkTe1ZH
/cMRHjBXHTfQv5JsM/XNLSh1gHezOpNzC6eWUobdqEvrakG+bdQiOWrSTUdFFL1/
S4LW1WdUOzJdyWkOv2RA3YooxnSP337PD8gjdyzOWIrNgl+PI4O2XUjswHPf9Q1u
mtpeSOpCEmy5K2qsEKquWhiEog9i/J8zkzCd25ipuMYpzORgwRFhTthdA1pzrbGd
CbXU2aOvuAgtUrFkwnIeyjpDa5ehqVFpeQuctd6GQsP+IMZpD5uIf3UCd/1Nk1F6
FTTmXDJbCAZtVTD8LvfJXRtQt1aCm+jhbIMG+yHfkdZvrx/iPQrFTiXOz6VMPt5A
Izr8ThsE5lTDD1E0gv4iAp1mCkK4UbxfLVxbSjCv+gjUjvmDXIJGiqnRQTfy4Lu1
R9HnyIOqEMrqMok+OLSqWVtcJ7uxGDtxUwzblEAaiJv+CYLmBc0ARaAwtsbdIh/r
64B0g5Mkw5h1Om+fMziLYV0mhC+YHQj7ArVjsgZkZnmOUn07ZP1y5GJa7V+rzolp
eD4NKoETzDNzW01VY+jrJBKCFRRExHvMQchD3jhz5IPPoE1PCpSyplj3tJ0Ba/HK
BKtX1XiBHGOHQUV1yQ58+yTFeaE8KDAktO7DYcjCmEWHUPK+nQ1Q1MFGGvbjDWOO
JY6QcbbI08VsM9WpLfEl9H087hZCL0BE1QMuXK5t+vdzI/8Rk1MlfAs8zpL967On
MW8OSkEGYBlR+JXQdXVwpWknT2vi6nM0Vx4zRfSvQDrGX9D7MGPxrjocmx9F8tAL
oCOS/hGfVPuddLCiBhG6VChq0H2ZNKisgbIh2Am110OcrD/b4tOFixivcFAjL7L2
6aBYSz3wP0Bz/auMoso9LSMFam732vTJWoHxID5KqQ+gGQITBaluGHYbH8g5MfLK
5PxofJ2SkVArZnW+lPl+t+OWHTLYcw3JEPfS5aZFGsK1ZwaaV6Hen5DHBgMbm+2+
ZZiMZUqtf4xitwLvxMz+5wbKnCvWfWVEe9G1X4I9U3ufz7tym452tCrbtffWiLVb
9GZDQ41HE7nn+VQdDPN+Sf7PGVETWbnr9XiLnqGyDUv/BeHq43xGK2GhyB/JSLLN
X/+DVOWUhSr6eoNnwb9yi2tprjpX6aOYz+sKuC824uw7+Bzt+135P/BqUt3K6fHS
cL33H1iR0XS7z2XnalzUwmmAD23dPYEKwBiXLYqs7WNapqn4DSJ8tllW8DjkUZKz
samy/iyYSxE4xlToLo5E4Xx0nXyTJO+jypE4YsY1wkWCED9VuuMgOcy5dArbQMJO
kLUcWXH4Bv9xsp/4e4RmaeALkJL0oM+E9D3zDIOx3ljFyCzj/uKuye94P96Jzez6
TYZ2o/HhLzgpF8j0nrFO68aXNR1o09Xfsbu32J2a7OuSZlmYF3/2JIwIb5fT/Asa
YyTHDkGvUHRd3V6b1MylsHB0lHh5J986sQxk0/fy20IWyf0MK2jX8EXRx2d6uOd2
YWqW2L5wjOhoQ/18fMRXtAkyyCNCK78Odt8J5DhGc37P5dLkkfwSS0stVxV/Fr62
qu18dQC+XONkSnx6rbPGHZ14kt1X3Qx0q7V56h9oGggC4VNOBi1uN/PeFMMoIp7D
SnQm/2vnXbEYHnVNE6QB8F3iRLlzdtJK+KeHxtunOX9QQpFacCPDKi1iS1R9uHrS
Pzr7s1WOl4miFvbvE32M4cFBY6uOyRI/GHYPSRevxwLFKdld5JTnbTSdU9RsQb1M
RCkWnFtvLBYz+cNqM8K9bJLUnvwlheXWjwBBDSi2urYCHAzPvOJi20xHWHQllOww
RJOYBFdrn/AInONAmTMJip22X8ePWOFd0ylw1pf19x5+jp5VvVvmSKYWxZ6EeH4L
cLmxNJ8JvG2qa2/TChvdDcaJ42LDvDHul2Mw/s4NuxAzkTv9BRJmLLgij5FQbqeP
8u6qO568UQN6WEF2EJrGvBlkfY7POjutZyqjql3HovXwRzTH2XOqhGsn4mQ0HNVP
PdXCWGwVeeckeSKRgT6I9s2Lph+yE4tgh/63n2POGMaD7TtrO5u2WjbbbT1dlkVS
CohRR5X7W+xGaTOG8iKGmtzRtBTktCZn4arPGSqEHz4a2GTvsvpc3cD30t3lfn77
osh+YQwnY9qg5F89miEy4sO8/0qG+wRaRd24foGfK96Rx1iR711Yy/k+rdZOHwTr
jTS3vBzbLGbsoUBpr44QxomNU9Ow7X4ytikMpQv4qvnm6jOZs1AN8Az0Z5XvlFb2
HBu0wGuOKdk7nunlOfPGaQHQz6Y9FoTPSMHDw8Ah1WLMCtB5sa9exc+i/qOcEowL
73CvNeiJuSPvYsBhGPS2bQFOC+F8CPGT8uI3/k2yo8VWoKxlMzYS7XnT2hugvfdC
becQkeuioldFD+sk1Zg7SI1K++ZnjGnfNYjK9963XdfHaI1LgiylLfEnxP2Qgb5i
SN7mg7H13bK97fZr5Z650iIA+caja/a7mdPWQIOlUPY1rFw6JLfCSsFOMoAxR3hl
OpkvoHiBi4XQDqVmIwn6RBvBV7LonLw9Ee6cpbHxpGptt3FCPR/ua7f5sApusUQQ
BK61RaTkq0fzYQhA6wN1T87dorIEZqbAQ4NUq0OAHURkGYVFGjywVK0qB67I5IIQ
3PvVjgvH3//4hb7JWZLwEJOQuu8eCAMu5XFZiufngk0lU1TeOVzEJBQEClB6jZbA
AmvRd6/IGp8pfTzTBvG8Hh9au40z+nPXzPBk8sLvk6ZvZwVKbbp10fYHC7X1mBlK
/55wvzGAh48CWk6oE9W1OSppDlqt/SlM9L9JC7rE6nzbkkZ/AAJcm4IJ2OyBXPBr
0MMOiu0RdpHzxu9K3T/8JMMBrWtyMhcmcxa1oqjgJIn8blczZVYvVvPevZ0YKO/E
g7sL0gLWEmVO5764py7XE7F8Ni7mj+Tp7d7fbgicRPxxUguJTu2bK8J7npgVZlYm
l8FVOghJR5G9YudjWIRh3ixCQZsqzhTbv+5x5nasj6pAbvc6S4/eSg2/+TjmB2XQ
WXTDNB7oqsHtlBEDw3mlT8hwIjn4vzGZVZBkLcHYKo2lvyxZOSwe0rGo/LcTP84z
1VzRy9Q2M4i+w9BvphDAgyWJMCUy8hZfuWXUmpcXrH8hwy0mSONqSBFwtbfhaDKN
A078vrOdq8FI9GsAMLleS/m2/GzlkC8lnXME3A/1fFHxeRdqZVL0NV5BpzyHSh37
f7fAE3vJXEB9PbJEIchnPaenAJTuoe0L+j1C9b4IWCczIbQszyghDVePNXpYGzmQ
Dz+xw4q1OKPWaJXp9bFSbnQ3uQWz8ljV38n9IEs1Y4INN2F8Hwe9wkAJ9yR8fTdh
f97ekdxTj5TrRF8H1B8Ti/giUCXGdIul01DgJuBE/9e6t4XRzmGt3W5JGk4nsILL
ykYe2RFfB9CGvUYnWq1zcsTYHA2R5/LYuboqsFleVz/nqbPlaKFfnNVDLDvA3e+m
0eH9BK0Kh3NpmuaNK3SmqpzP9Ae+kXU2eHJ9sKBGE452/iPrb89MhrMO3gjMj+6p
p0HGwqymDkl/FsHihZcFoyFIdbgfTC+CdbCDfbdFNSFc6lRls4/gmEqzNfmtMwUH
m2CFw5V8BoaYSndJVTX6p5rcffA6A4TRv7A3LahTNY4v1Zw2dDhOdYk1GCHlM2Up
C8DmMFskZBDo63A/Tr5kBAymM/szWabeLpPgQ2bUaYCzblRnVo9Btt6XbbC1pSPF
Dfa0AdyARcUAM3OYaYDZ8jsP4QHFtJJoGk+tTw39S4C+bjkpHcqIWb0Ad5ppGTMZ
p+Z+acC4hTnIRGvt6CbxrD5/rVqCXbszIdCjcVKDvofGifkiKv3vyteQlGS8k6MM
jm2H4RSweo+BgjXrRpH7QrzLqvEqc/QjENDlL3BbxPYTb115UPwZpm4i6UrRRGuW
ek9jXL7hxgAs2q7tw+OmyMOuoWydIvzlWElqtuSgrdcU6JNoCRXKhHKIisazCs9K
ytXumXxOdJ7mPyj9qyS93ViN42Ixv/V82B/hZFWxS51miV6fzKG9Avpui200LlXg
QnWeU9RfKppSyr3dDtOPM+t8WZUMyffCfHaIYOjseJ008C9ai74gYEwL+q4cx0AJ
bjkFB/cdP9qgUG4SofNpUXBRjwjpHUnLgOthvjHT5yoJOjcvH5iitlr6uNMLDTi+
x+gmucT8myz58dL/43M9jkoldhjuo7RvbXBwSxZyGn8AmgtAjAqJigWbxRIbgvva
wXbDXB0mFXhdc2OqtGlKjMpm1ySVs3yf9X1PpeKIHdKRhqAJHt6TE3NGgUfFvveK
BxtLE5BYFBhIGiwLlSRo+CtTCAC01bU3ZSlqAacz8HCcqNhByCCy60Z8ngzTBAqs
2IEAo0YeJhr0F91/gvG3ADmMguf+DNpduncO0jjuwVkuifXGNcH5oo/FGVe6jtbk
2rVuSdaZE+Kph3utoxT4TpZnD7jd66hfmtsgzDmSqiArEHD/nADygrU/1lbqEKZg
d5cHFr0U26qag51SD7PwxqIzrW3/s8syc2TON1Lu9b3Xrl8oTHFOA/kgU6i+EwDZ
pMhqzqZ0Yjt6mFnF8MTSNyvNMzc5wA8aAJ/kNAlswS+Pn8ltM3KrNAesyLcmhAhH
2jg9lNuAfW/asyzyfZn7FQ9f2lQtegx8CO9TM2oRl5TwE6wLBnV7LTb01slgP0xc
yL3TbWID/UuPTmhPiiwWzK66YUeGPbJN7rPGAFIjYfCUqlJq3LGFbf4hhn1dL2Py
92DrvS+PcvGyzU06CB1/DECYpULQiZQ10EN1O98ID0IPTwgobjNNbMWKp8waTu2g
J4s8MzNSPUALxHKDmAaDtk87QZOf/pJbp1sea+px3TyJdiW5SL6IATalRjVNswYv
o2AxiMVEGuEiTQTJouyEtF2sbyuS2t8tAQiz5G5GzdFfJBiEai3h2HRfddpZweNx
0fqLTk9fHk8YAggj0XJdDcLj/M9wmckPEba7L6nUegzQa0hLE62J8+mb5WJ0UlpY
uPetJdAH80C4PTaqDu/QPQob/kobnd2FmbmIHp6M5dCUXu2RuuOKx4uIxdg5MW3v
igw5gEd6P33sZ3HK7bjIez1qj8EEm20liz/D4gsm4tikeWqefts0VA46ghq6NSRr
WaAiZ0p3EvpLMRwH+JH+KEGruH24gCcAodc7rvGx997/gpdRdwwHRWJ6uov/f/uF
/Yi8YFN3IqJZAqKXXWvdUy2w56/i7wAyeygE3mjcmQDMszxaWuTZcMlUDVF/QeZg
p3z24mkG9aGlhS6M4KBaYsX5Ss55X0szXzi7Gb4AY2+jKcuXJDT2lSYqoJP11Nmh
GVrcK++rn2Qv/G09koPW1F0+o6kOONGnBjCYuj2nBldgQKPahh56W18VyUF6sPgk
zPR+DpQyQCPtrPhWCdi2ai/5B/KD678aaEo3KNxSNawvtVZbtxclhA144buUyEaQ
hlIdsULWG/HMuCkiD9CRcP737Rqfh611tOtxsF7VdRxr5vBhlTXtYqKk4PnUm/h0
QwA4MGUiAwDcpT2TwX4IN6nc34Xot0btFH1oJyH8ruC/0z8dRgXRqkiJQ/A8RLQG
1ZDEd7Je5pxaN+uL0h6RD2aMW3dAXvFIouGZ0mm0pEqzJHFsL0Bk9uf4u0UdXEEh
2AiiYek+3HvngGXwtp7QHrhkY++NeJ/C0+PcPcMdQ6zLr04gL4xtPvUwgHzcfBL7
CcLVQrb0vYvl1GRYDYjK3w5RvRMj1GLQxdt/WcW6qIR0Koi4ZbsyqGRHs1gCbnGR
webeUKU3Eaj/XkGwSdCO+Q7tqY2A++4BjZhbONKAjCGwzQp4YEZ1mnUAQp86BT4S
yUSkev1tkcdU1mp38yz9GWjRpgDl28TTSoplZRHSb5HpZJkXHUei5nHemobrEDel
1cgQgFqp5yAJthB1IGzrYaD4FlEqTyB40AnjdjOKQ+7r4HXFSJfjYywHlbCO90oG
pn0gTkavMY9dv6BFNX5ICIO+XwfW8odZolrZl/arXPRxXNnqsBJz0d6Omwi9GkHg
ZC+sAw47xWnBPWjocU0UmlUwQR3b/sDstxlNztRAZ0jOaITulJRVeErrULT5rook
ti5bGW5Pc07QqNeXZD+JXfFXR3kIyFCesx59QXVRdsKlqh9h+Tprr4qHmN56dwvp
BlVF3WeVV5auD1vAulCJDeE7nPRMuPU5vU1jBe5dalIGxa3tM4EwpziuRRiDt7Hf
w6ahplZMdnwY9F7zWUMBtFb/06n/5svMtzl9BvTFH05BIA6As8Xd5N5FZsnVksrg
V95Xi2P+z7bBMVg7PA5J8masyLx9rPxugc/M0Wk6yzzgomYz2EH57vvIw2xVCwyh
g1Anc8eSxsnhpLL22Ml/uafxN/B9ml/iQVoQg8Q2xe6zlJfuljuGx9oKA97IlZ7D
C/jnyG1ayD05l8szuTKK740CMGIhdoTjCjzlt/TQbVT1P9DVGDSQo+Ap1pjBRlfZ
EDD0Jg4+FWGOoV0urcGOnEJ6bN5/mo+4Hder8V7hsgrZAZ2zcKAFX3aqMr0HVhln
YCNb+NtOpvaF43w+hM6dFaE9dku2N6gbX8U0ZZyHQL++11rKaTr8sxnLYU3cwq8D
y9y3l3EBul2M0bH2KGcw+bKcITCdQAg/l0Jf0+6RUBMFuNd5LYRF6zTT3UYiGnuQ
SORtsvcadB/xBfLR2tYB7lDAex98NNTJf3bfmivq/E5JBAfX0sdF1BdogNQCOBZd
XTFYx6PllbLqjHeUvtbpY7CtuYCFoglq4ZxG++KSI1u5rnr4jrdbbfoe0Ger3nW1
+M8Dj13VNMoTTjZCMGgjRp++3PUala8hoRJVEFz0xWLLsA8k5Wayvk4yMj3e3ULX
slxYvjyGQpN71sKvYOw+8aQJ28DXtXa9ISy56eQvS5qSmVUpvJbWizz+PBN+JDdo
//9Pb7nEgWOtoS5ShurcAl9UALlSO6qHkaAESnTVzM7pOA9ZJOr/I7DTT380Bp0l
5xsh9mLERYhU2xCxb58wjdMcrHxyUlRD9HkQUvwl0BbbCOG4NpmrEhVgZkW1GqAw
iNXvOHWihjtUGA0jkyWNyTQEwKbEbiRI4sWQgjpfmsITnoqXJsarQcKcsikvxjw8
YyNRQAuI7AomuzraaaoO0wlQlYxU23E5NzpCcIxA+LOfngJkPN+nYxpJjE1TdDWK
uYBUl/Rm2JHhbVn9JIdIDECkfhns/1SKxGMiX7sWq+UvMXPGBMfukVn+WbZnlMY9
xG1cpCb1GzCX7UXenQOVsZx8oZue2SWothUxqAw+g20KuNDvhiyN/NZQG73Yya9Y
SSYlLiSKsbjWJ+zzgsATUZ4xBGK3llQ6GWNwEMjgA7D0/kF123feH0rqu2GU7xHn
8rM0Ulxqmt4PEv+z57IBUukNU5p4mARpy/4mSLCdlS4zKI4wT6sJJwbvLlW/O/cw
KxhDz5G0Y7UMBd1l+xZSZtjcQG87T1mRNVhqJAP6J7AyWy7l+7dMx+4fXyVTOw4v
7Y8Nty2dchq8p0NDliOIkFDMVq95PDZl9uPWlxFSYXlf7T4vD45wQPwVcaB5P1de
nH7CagT2NSJxdWwMCuLGmzlIXOgILXE9+EHyA6JuYiFGJiH+MhX3grheeTX5LNNT
M6YS63f2P7R772FUHpIGxSsR4kq3+VsW5ykxDISgM6UO+Gn2StuRE9YhZ6i1sA+a
W70aH0WeAPgS8FxEqjEIj5EJ8FK6yV/aA23eSL88yrhQlMgJPgeozeCyzaprQQXh
RySwiCN3D3adUXD0UxRUv/A+w3eTkjWrIpaspwVDRwuY855P90fRSrV9aSZNPysT
U8kmLLGj8eFEN2+HMUlG7tbBM+ImeWScz54FhCjmrTuTen1bK0TvS+rfyMBWC4C4
ky44+0YprTQH3RYpdpgJjY3WrDuEFWzmSIYTMl6P1Z1xXI7QxlD7gFAuGjB6Mv1s
eypi8Dof3PiCpDXXZyCSSiq/MYQeqRVnIP2xhC/dIA9nMiLyxJb03OoVrAUTWClZ
KqQvFM6a8IjFreDx2m+239N+2uEEeIt2nOOiU4X1uoI3S5oBYCn3kWNc6k0NKOyv
7WCx7JKTyswE+OamfYC1Fg9V9bbfAFnp6RCx7tWwliBY4S9UoFCfSkcBlYVaf5FO
yC331aKgVC8ZufHLxcA3J6iySUf4+gy38p1iq77M3dnjX66XIkXMfx3UKAiP3BpW
CmobrdJvayduYYiw491AOnlx3BvvT83p8YQUFUflV5innFktYXvUIom1/IMfWIDn
xW1d/jGXwlB+KzabYacYnzIgrocOF3CsmDLf4ynx6TsGwud/Vd3WO593igjPoQ9/
URAMOt7WKTTWDBG45Qj8YqRMenA9oPy3mYHtP6RhnCO+4UlOMyl6zL1698AKclNn
TNKtCD+zxrT1MVxWdyKf9xdraZ0LeBTmunGy0Z3U/kosrdJJZdo/1+2KkBrzCfK6
fD2G3cztQr1A1OgN2fk6XSzIAnhYU+gnrfbWR64pqEo8TNGeI6HAie0bjFvXVqJF
gxsmlHgu/7MstNHWEo738CxsmM/vKmswJRHksCRTbrp4cs3Jym6jkW8D0ZD9jkOE
a/uMCd2XElNmJrP0OfrP+cjGKHrvvfZYQFnmj8rSYf89fLdKTyOu2b9GsQTRDEla
qzufM9YJMQw7cjHv/E21ecoG8BJcbJGN99UarYDUdIUWRFr46S6c67mn3CN+Xp5w
SbPuu3Gi9qahyOUTJ9yUdwN1/YZpSH15fTl4/QDo3obZdNvg8lxy0D+OJY9zUWnv
wkrl1U4QR77NVQWwucDUMVqL5Thz7Ey7UWkToiTbFLnxzuF4Sk+V/gnRs0FZ9KO1
R2R8lUrElzO9qV9FsN1CAP9WX8crpaeipfbLxSjVd0HTR5jQ6DYtlAWRdSHB/jjK
mHZ01SZTjxl4n/cNE13mTE0FMdnHMheSkTv2Ezu3QLtU689FrZpN+v53sMXq6SZu
fkWXUSQB9gkZqYNIkFEwu5MQ7idi9G2QcHqPK3cLdjzlcfR5ewqdXEBxuQovxVRM
pxAW2F8tOatGlfyx5az28E1Ntnpnp5/qmhwK5nRgfQJhFo3OstLLDM7E2nAVRJb8
nsvmdUAstRviwpd396gHr5MaRfO3ZzybeNIYmYCE+6DM7izUyVEyellFo8fn093e
JL0+TL6CcZY91Ay/QjMF7YRKwKvWvDPiXCFsD0b0jHEoDKQnQgCWdRODGFQLbJld
nOBHUifgFyuWBo+X7lMgFAU97xk7ZhuVe8SXzlexNnCgn6aTqz543Gkaw3jNPY6u
+taiZt1GAORejinuLGnfiIiNQJ85qTZhSpZ/Hf4dYEUU3Mtjg6O2qoNsqyjUp1WY
iK5bBRifvVFx60CwTlbB4tQ8W1EBfyAfR+U7LojxssuUq0pyg5Op8VJz3PArbbgZ
wAODFIlRj4dgNKGwtIweQqpgPhuXPBug+eNBhMG6kyIoFyYP/jj/mw1hCb02ntVj
HvRuhTeUJWpoN3ymdMNCtxvEveQPxUEEN4Q9OPkpJ/WXzOy+yv6Mq6coM0Fm8SUO
6SJK5rZqAzZXxW9XTmS27cUN8M7i55L9vfc/yy6Nli1JYcysoL2pMgoGurNvNCWL
mTMuzDyXEo6Vri7yYXy3psL+ApSoEC3198KfTW9tpdezMvjycoMAOx7dkrgvjX/C
ewFKxQfMUPqwq1RTia3BOEbTTyh5ztcgbM6FHQ6nu7FmY29RortA8hybN2ne9INP
byzPh0hwBBfHp2glBvuv3pUHsG6V/3mex07vyxuRycj0e8uwrsbI+Mbi71l3smIZ
2JyK/vyE+2+Tw+kv3J7x292Dvo4NrMYF0UU6/LJeNMIOmsWHNIHFrz60akFnxNtC
3mgZA8P+Gmg46t15C8UxfBMhZnWlb9BNhcFch6aoxXXjf+BigDZkvzRV+cK1lXo2
5thys23HRfu5JrFgGFsqehQFClCO5fI8p245txsoKEt71EIIvLknZU++CXLPPXEk
jW20zfz9i7pwcqvpVKu6eA0scu29oIcPE11+Ik7J/S64TtkRcMERCZ3/sO+gimUw
uD3O6cMZ1Vn6gLJMHG0Z970CKfNMyLCTOsJjqwoyHKt62jAjX2YpRHRqba5/Hgde
3f7b7hvVvD8Tt4oqgqs+XwIP7dOm1jeaSijg0iLST5nReUnPjgB1YF+721uVRQui
pLFyFYc2FyeflD12N0Kif7DORbB/F1b561g3G+GptCstkUesY00Bh1pO6fli/nde
nOFleshdDGaQYS8PQGKB046RULSTNZHMvBKYPDN5PgjMtBlvXVDH1X5qOEnV3/X7
Gt0AdQLlzfuubf4Y03nZfm/YFDoqymKNtWUnUBdld9T/vl1vuZ1QViuEqeJloce2
xsNX2rG2Kw5b4QrcyW2h7MEn1w03WhRjVS1XkQEjlU50X3WV/UiDFgmNZmQwB2By
wEz1hMSCzdnEfP6497oZ77079IDTLcOxy1Jt4LqJolSntZM6CmnpyjAZh0SWnjAK
B94r1j+hf+K8X5lOacJLY+LCLBcLffZSW93iL3yy8MwpNdXaeAGKMH6/PM6InpJN
d5ZE1ebEpq6EArIZyLnczjQH5nVaTWOp+j95UnclaIb9MLZOos6LMkhdBYcarVIA
QIfZSYO3JaLW24cLQ2iWoVXYwboDE2D7PsuHxXZuThgtJIg/06w1xzNyyZixfYMj
ALnM6lezFEhs6ahDJysX5gW9C1BHWARooFV6ihH+3WKNwhHTSeJ8W7wkzqKbITPS
IXrk+XrvTegXKUnXsdSM6NtUi89CFESsgVnaHAn+H0XQ8lxSXqgQkvJ9QpGP0B4P
2Rj8kuuypF7t9BsATOG/T8YL0T8AfBHWThTOwzKmPCKoaad3qVE7BnMgbUOLHAOA
DzUZuNRSsLG6cMfS7FjE68FWIT/rBkCQtIdhh8rQSQXkrZewPCQI0shvuXBLnbpt
Ov/E0+zJgGGfwjSwpK6XXLhhmJvsjHvucbtKmXsujX8nNo2b6GtS+u79ChGmNzlB
8JUeCobAJAnRhqePVXCGgCqeZY7rRau30DhYLlPhHYeHjrI9BKdGuW0zz+JYcBW/
XvX2iXiPbV7cJdUilhcS1gFDpZQTI5VouV7/bihbsU/KNxAooGxUogTrhhYfRcb6
62nYpL+XDEKEIauoitnCL1+oJufR+uDQVGcKwfFWp+MAtc38E0bW+SQJZrwaIb/0
x7JzkyXkJ8fPDVPI2VISLeOcMUsPPWPEmL9+z3WoqTeFIVySd9Hpu2VRv5/oKwme
1MXwUwVN9vWq79FF8Yy4m5wmowBTzy8HhNTN1DAWIeQd/2GQ24K0D7pSoWs2SNM/
PMtnyXpduSDllDiFTHbQLWqlBRxszaHo/BI/KOhpRxdUmuiZSyzyIdcevEh7+hP1
Z0rOGQNGCScUuNpL/IXGQ0FgcZnLuiKxkbWjC8ObrjOkn/A5mRwIr2t03NeTl6KY
9hXeZc4raeGtu7NEbI4wrrhBACvhyxG066AqqQFxMY9o13/dcUSuRKYrv+CWO7b2
TEnqmkj13hj/lgp/IXFZGrQlYfWdyFyvTEBdWNMoPtOYts2C4xcrqda6tjsqv95o
0u+wMgQv7CX74B4gXKFjOynyomzei5I5EnFpOjDwr+yXJIK+WBVlih8lDavWk4C8
kqCh5Kh6l5/a5nrT/y0/FQsj6KBvqZ6qxxyZj0qZ1V5bBDUIYG27cL9T/N29olh1
RxnmOeTUzcOs8BUAiB/21ku+UUYgl962Yx9ywgMSoTi6uD50PrJD8HVCpWur+gpZ
Z2KYYoPP34+ajYNJrAMNp+Rq9UxtubTZylFnlS1get+4tnQ1sarCQtCHYvhvj+Vo
Zt4hFvxT5SOB6HPaeKVZNkmmdOLuPONP0r79pdR7c3q2p69GIJviQTOqilaSerc4
sRIMuYLEsVHFonAyQOmXgsyMSkc9lLoWu63PHDPTCZoyFe0d5wnnqBfIPQu9jbmq
TWEzn4hsIxRegrBUb8Ho057TcbExd+aY9qtbLxxVCqPZKFndrhEjKGnku2DVV2OH
9J0V08xInzXfsq7GjetchCayTCCYM/e6cWzq/hrn6suC51xGfpi1xy2wzUkHkUAa
HVo4Gk4jXhHjAeB8z+4EvLRr28chnueHyK/0E6qJepyXBnC35IiNB5c7Ag9ZELcl
fH9ICu4ym3Bf/P/3/U+AWZ/eF8UOg8kNjVh1NtAKMfVSEawQvkx/ZRSNm1JncTeG
j7455q7LRYg1PkEnqdzST4IyNiGS33WWD/I9Je7zRxrWghp5ymNy964QpCKPEa6j
FKDNUUKeu7nbyY9q5nRE65zyI/u5bMuFbP5htJEmRbO9uPYGURPvXi7FvYxuKBR7
PrwZ/NTGAHeT9dCsnCrSA/7DXWY1blV4kEmoyaQtpaAEFhMohu1wSTpb0O/j98vz
2/b1ELo98jQIHNfS9kpMLoih8FmFxN0LerlXwn0R4+HZnrIoastZZTEOgx/oICHA
Z9uq4jdbu6dpQuhipAJ/d3I1fMFXeX7utG6Lijb4l9BxZGgRHhzHcamP44BI4Rw8
/WnHcAEmzU9r/YUPOWbOPMHcshlzrheTccaHAcDbvRxNsQdVhFgq7pvpTMTjdLPD
dcIT6xIcBfTbesL/IxJjjaJKtP4WiHcGCYQAfy+1Fjz55KUpupDxDB5dBA4JrOcM
XG/nhuc3xngy6/8AVg9InCbFDJ51pZ6N0KgRqt0Q5npH4qp5uNwvfsCrev/6ibF7
9MfotMtIqR8jUdXLVdKRg0WuYbXFkznoYRrGPsde1XMO+coqAV2Udjk0phm6Uc7z
KxNFBm9AAs5yFE3FZkDd+x8LN/3/yfUQOsSYXXwJ60IBUIBy2XaDlNFjulXqPh5q
vdx+TQTvNUvfoE918TNxMnC9UmI3iMKqznlkG4Fh/PHG4z8sLEYKfMfFlMXlGM0r
TZSr41D1n3AFKo0v9kPgPJjere/UKsPJdNbWZvVPo/ckJDd1j9CV+oEqgm+Rmt5l
FyjwY63YIhhqZnPBXONYlXxCeOZArLYf9Vk3AR81H8ueDIEAbGtEiRelHNte/J7i
ypQDw7Rrg2LVeJxaKjba/O/oy214IXFThVbm+OASsGuIVIz9fCpoBzbnPAvKX33P
QX3/7Ohz9wwFbJEKdfauUFwhyc+J0EW/FZ62ZVm12NTL2oHRjEqsjBVFaM+JSZ12
lyfWhH3Ga6sB/87Hm38/hMYGs4by7fKTocdvu69FN0BwR/ErMqbwF8Y4cmOtMleg
P1drcSF5VDKQ/N1WTpJfriV97P+aBIPpAfNZijxszRx8tbsXR5/pgSml5ahgu5MP
xg9Gt88bwGrTmtbEeuDcyKZjURvRgk3+A4wKw8AIINUSUuxNmvYz0NLwGFizWv9c
bkz6kMkO6cIQqAX/b24djDPgG8thyMFuoPR/vFVlBy0UCYZn5ouKfU2+5aaXoJJR
cmQ4gFyh/qzYmmIRTGq2Bx/u52UaCFzBVGges/5qBjNGW5x3Vt392s57N2iVC55g
TnSgbNw+Z6f66KoL6/sqZisWS3/BICsVhUSkSiiyIHBu271U0eKzPScQ0PU0EbOx
74l/eLqIa3+kNgL61S2ZGP8Qp9oZZQyvxf4EKF+nSUcqKYeKqiRWBEKfI2ZroyEb
LQVEwvA0DIAETvTgBH5ARnPeLjX0KBtVjX8mbW2BrZNm7/YBi5uupA/nm4PKynhX
LyGL1ek9af/YaqOrAKEMZ4WD1Ob0/5qDtscS/HF8qMUZEWda81AEpiWPRSKVkyaU
mOnTI/iblXk2erKOyShI0kbA6JZDDDzDvgjPAJAyu4SY+8dWQPv7SFgH/fOyVFHs
LBzpN1MtTVaxI67R0pqp2rkBEEmsvzHHZhWBF5d4hffliPKa8RvllzISEmgkW1a9
LNCYe5ZMnZyqu3OrnjDkRXushjL9MxJsyAaG2KoOjeh2E0AS0KyK2A4mNWPtAC2L
KMYQo/NrvLAYi2W81afcP3oDvXPxFFnatafSLwa7mWez5zwkin2WiXViLMSWTK/0
wJsIlm8ZY8jCH7lkXQEsszDDDcZqa3Q/rMgQCxgtxXNXGUV8cV4BEw6fv08sD7aN
aDb4HpHA/Glx3QKjohs8Rd4X5imMvLZJkQS2zL0jNT1w/Ldw1TG00UsVbbcr1Mjo
vTWI53Chu9T9te7au5pC3qV3lVA2OuanwH0v1FnwBgL2OV/VTWd5xpRCJNnauksV
PhaI6XDQKP8Bv3oo6n27PG5A4qi7lrIGXvP9WXvMzacLaduFmyilLJbHS5KIftkx
7Bx3HqSIanRbI/7jj93CQ1KyJhM/Bet03ErURN7q/EN9jL03+AIPj8AT3A/AR45r
rs6pCf5HZuzS66eVPwPx5/iipeCSTW0gNE256uecKMWU6GSd9UEeHIv6vRQdLexl
ilafBvJtUtNhrJX3L4NW9IaFB+JSXYQbBioqF4OHYe8Nc5e5W3INLA8fDWwGxpJO
+x21FYC7ub74BdgYMunLMQCjFyxlh9/j4xIliG4tUz5mRm3K18yQXU/hfmAf9yqF
BSV6YGS2apHbVFFNplL6wqB1bEIXDbhxHieVt55wK6licjIVFLuyoYvNOOruBySk
YwlND6Mr3h6EkWDlAZbWueoMYT0iYPfyh14KjYTys58ht9krNNf4Oa7r9bZD3TO6
V6AgZtXGfQAgaQ/M3AZM+wMDFkAJmcbM2zOurUOttbp2B0kfYzaHZAZAVPgqmHjs
iXo5u/bVm7EebgypzhDJq5StpqoSQB+ryGL3roR7gcCtM+5RQ3SUF/mDZ+pFwy9A
dTzBEhuTFlQWReIdXzAPNn6dPrvL+TldE02c8w66VtHg8LafgVWIchyLTMT/xRd4
C4MMEx6AeZIK1wlog4583wdW2jG1D9ycqTHJSCFndACQa5gK0CpV6fQsIlyifi+8
snAkyZAw7iAC/ZaGd8liXBxnKMr6i/qf2MwuH7K65jcK+qQaeBen3B4opy96yeKa
GtHWZHR5Z+KkVrCKC3Or+sx1dn8ekPXvjG2JypZRz7RzWYY8jpXWNkBbpkEuyYYN
Z6niPX1Sa50Hb6JfytKhG48ksoZsh8a1+Kwg9nRg9taMs4sv5QCm9Uj52g5qm0GS
Yfmn+F4KEpwVaX93mSs6HI7RpPakIJgJnrOjLQJU0BUy/zvFDR8+x91IMVHXVBLS
w6eckPG8bOA82w1CE92kBdxIEH0DGC2kAI+YzpYzGJb24rJ5SvYs9c62In/ljJAe
uczEFSwDSaeqO5/rYGyxpcCXHI8IU4wO2DTEEsHVaLEN6dTD073spLpNREfmLe3f
lDOBOFCCmVDxpC3D7yDvhJtLWxSI9IJQmK5Qh+lOxjrKFQetZbuwOSI6LQq8mpOe
S+Ao/YaAuFu5nUGXmy9YXrRBBRgT4aiHaw1GRfQXqGjSXyuBuuaqblXdMMRwcRok
BIWJmc26ILYQTe+3HAYZZrx5Um3j0Ywy99327xNWoxqJ1iqZtm5XhZSVXjqGPvDI
+ahdQUSbxA9fKKlbIRPnrxcjCjlyr73I1it9WhgSd44Sw/N2rlV0/g6qJmTcJult
Iv+fBeH3p3G0zBPilhKawIj+faQDYQ4dZ4IjP7j/gC6UFXun1TJg1MPFOoleATkg
R3UU8sz0O/KeXjgtGjRL0npooqME0GJogJ7O0SIgBlDWAIeGghkl48XAq2qDSU1O
Ph7JPmOK2HSQ/cQcaPta6vUkPHSf3YurZYllBxvMeauLAjNpsYhdz7bBj3bGEh/z
Kqtkw0StinXv3HVv7OtTYcx6y0h2YPi6nvinvZCG6Dd1VyRdwLrNjks82Qo0zoQ9
4xHkS7oT5HPxXLmJUZLw6ye6jhossuyRWl+yr3pYaHozWw81Xrrs67eFrlL/j/En
dA9jSpPt7dn4eJrDgZiyuvjCvIR2cRS4VTwtSCZwQOwj/TjZw+VdKuffbgkvb2iK
mGWSwD9jMVnC+jBglLuBVgaVkYt/YsFkklhzV7ug2DrFvw81oWcUbEOsQ06WzSGW
nHswb11BZFw1zm9bFXwj7kWI+a7NtatRLcksGQ/SPHY4Z1V/3nK0jlfOPte1Ggfg
aVEII1obCdunQPl6xdPNBiFZI3bc6r4bUPJYSNcAF3bFhdppWECNlsGCwx4BAgvu
Ri2tGNUlhEoNwBQxbANTi4DoIUIu+Qat2/3XGfT/HIjDm6EH6df209pb/0dzwf08
dfsMF+D8my8D2iCVVztelI2UQOyjceYY5zs9zX4OHj0+82IvS0ILuiP8HsG6wKVA
/fBsj8Vs9OIQJfDd95qqCmmx0GkZTHKil5mqwucAhjSXZlEqK0M52vw1W9RxuI+p
TgPn+chGrlwn1yF/kTSlmVzBhfz5C/mvMkGzA+vkV61G/QdY7OHBfSU/3q4l+wmD
zGAeLwp5ViChlvBuP0nZ2RPm8HMjwKPiRUrdSdmnRRNy2O9/cx25T/2iOCK/ENQ4
Q4KPEAC6FfFuCImYLuQEe7sHoOplmE/sXBKlXB8OdgmMOwnC/XLOEeBi0Kb6cTsI
91sM+oRubi71wbTYamqT/v9HjH5wAY/xjEQnnIaGHvI0RTcLdZZMamiDwCGEDJUa
78BiliS8iz1WNwrpulZYMuoOBvOCmMqCn7xPehTs3AMR2FgN1S7L2MDPVWqS92qT
VxtbtkTH6qWg9uYFgBDX4q6/YWVxU+IxlN3oHw6+FFgRxDGf6d2u/y1oPLi1Zq7c
bO9RvOkQ0mH/VAMEPjRqCm5HZJqKK6M0cPUnscv7QhT77/pqueR4joTZTyo7V0NO
H5cbu550qzlwzsYmqyzwIHqmNjwFGlFjg8YLnJ3MhRDUPMD3wdzmbEqab0FK6C4D
dlkwgOdBqnqhSEMcgE8ZCpIHviZLlQfwLsJfZ1/GZ7cjWTO7GhD2VmS/vc33ztHM
so12dsHZPYPDfZD0CRpgqAyF/W0d1ZK4K8FHFLjCK6hdZxzT/Os5g4eaTHmba2jV
JbE/T+Tc7Y8CVxYSrbv3ctaN6Ne8gZ6MRbrpCePM1Rd89PnWVq4aRkbDtZvW7Y4K
sRgwcuavBN9DbWugic39igksPteochnchTq+f7XjvHjijH0WkRnjvjrvXj9sqGJQ
zDGm2d2ye5vzekGr/U+iBjdVd1c8TVGP3EvxGYEeTfO1tedsEOVaLq8zvbwOzryE
ITGdslLq32Dg1rVjsu3OZJUjBY3NyOnfnCwnPKuQ3E8uVuLfVwJv4CXC5gMY/nm9
F8BFVCzMsD3EZgR1fPrJdOq355YVzHThZn09MMI9wj78l20h52Xp3vpBkv71es7n
HzWdf5eOCe7iOmC59C6k7JldOIpA+ZWOw7pZuByt7ssxm8N/iNwLgJkrYmkrrnP3
Vw7UvWIrhLDMwju5p2yGUtsbKwzLJjTd5mLNDU0FUyki6u3/4oZ9qpWiMUTQyFqo
9ghAfxjLp6T2IzoQ37LsIJiCYE08YPgVCY3C7c3VZoRPT8EwSxLfD15szmeEZ0xg
QfcOPK4ZgIwRq8zd1djqomiDDaP3WcMktSN1/vChm/eCLgQSKhKzX8O5lrEzoYCi
TBJngl8+rL5Y6I9hhBgj/9L5kfMbYS4R3BqwHBz5cgP+AEV0+lZ1fEaHO56c5uaR
vPDne5TGYkKpGm8SOp/b2C944LFnx9Yi1H65XqYLpYDA5WrnsZA8QDWQZaVwl/oT
jpvUL9WVpTGrk0146VNDrWCNKjlNqvGrtOWv4UDlaG6BQDNdALqJP3qLUYuZTWvR
yBJGTKJTrO4fYrtyp+Bg5SVeloxamW3R5tyXhpYY8C2L81SdRKE0lOo+VkqRlawy
0EzYJnzj/OKday5ovCj0iZy3f3Ru4+ta3OTZIFyEc4Nqocx7vdVQXq8slVGbugCU
E+7A3WJOD/TnRUrQXltLeDyo1xe6h6ZfXRJ9uJNEv4zLf91I8vDgYa5y1yCZ5UUT
FIeLqsVH36ly8/6rRtxG5iurN/ezK4xS6bTS9c3dh3idPyp7Fzoz5I9zFnR0KYeQ
7/zdj+/uQDAunu+d8LsuVBZB0fm3Ixu+6zlwRLxXEWzYxWGnWRSK+zt5LQKMeG90
jyCB3WlN7NPUnhG7LiMPq5AASV5XSe9pCKSjRUsSUlqbTGQ97+kYyImU5EKNZTqh
sAzKEliR0L6mKZopyIU/FwTEGxg6u78h8deuL+2RiwkHg1iT70w72tFc+fx3Dr2q
T6cOXAhRDvwPCegHS+oTpW38ZkNx6n/58hy6b7CpDBmixxVLGKE1ifaf/8Yh/9UI
bKBn3TVKxXoQCJiiIYPjFKe1MfYUtY0f6N8pDyEBFvkWGUtXP5f4kV7j7plDtFw6
Jw63wZTMwdJc+4/veFP5MylxDpkzY3TvA/BEafj4X9Wycub3EIGr3n6L4hjCYSQF
FWK9t43499LlZ75CKusvHRBHAxi8/bVhNkNtPXfMjMd3F8v7Lk206vW8LSCbUcdS
+WzUAjBTjfPyO/tL1d+o53Cm3cwD4Ew46kZvsyzbICKF7nc+W+HntmiNBnJuy8O8
Y0iyO4U/HBNMZJag4op5km5DfUcs/391NhwwPW7RPYfJ7o/eRX/tMTjlmxHo3WmJ
yOJ5lwWjkMqMYMvouzvEvKH+sueCLd70BXk12XxcRnkzFMThbLq/hsjNtiHindbg
k7CYgXrzaDeZYb2ydwlyKf44ENJcxtO8vT9Xe/5lLBzKDjWI0joTzc7bOXxID7yk
q3Uic7UMJJj8sUHSQYUvoOjYhSF6muNTR6k1O8CcYqh+ErmXtprff4DhBzCg/mwr
qXtPIgpc0NFW2ItWAw9vyWHRTwd0/JxjkcsHR7GQWaH5n00jEJl6rJkuJRAXXCx2
NlJA8k5NEfCSHQ9it/xn8wtEjJ6utVJFV9J84LQ1ULzf5GMjgI3tfxm7tc1v8lUt
0NvyAiTbTh9zc/7RdT/HO42kKlsyzkaBP65CgyFwhRymjO8WB2a0g6QRmb5RaJWC
7ae/sTycLIrqNGyqQQv5sjQGBxDIoU12I8YMeSzMSLK73ObtTVyUQt0VlMC0UdkI
55qLa6ZmJJEvZtmjPTB6AH55q6P4uRWufbsogkfv11arb7kNZO11qBjhexR6MOLw
pg8sUmMmtbD42tizDJNCKdFjm1/7K2y/t93kVH6n8cELZtRiYmjfyHc0/Z5fye/o
4815SFSserg7lKG3mnumGogIDWTMCuygsptO4+xcxjTjN2jLhYVjBr12kqEfMjU8
GdiXXD79amphDe6P2PB7uqDfZNlBZ3M4A9G2zdooK3naYJs+Edh2L4r+TPPoHFci
05b85XnTViTXctDKIey4bbs8MuVmLWL+8x4ZzjlE+Oyk8N3xVRZ8MuySlU5ElVUh
AK4GkdkjAb/7DFdnc69tn7L/QYRaXUx4DgK7gA45uvW1oFGimlBfTgRZ3rPHrk1y
W2TWd8IR6GEnwS/kNxoDQPCSagXL8Y6QhMvFr8zUaxdDFbUO8OmAQWqZUM09Fvio
+T/PxJcdwMgHkYywlDImcc8Vde36DqZ/6buFQK0CH6rycP5G+BZTBPkCuuyPaUvI
jSg3IwJng3tDI4q8sFg+Kr8PYK7g3ADW+eaIxUVkfNgLESx6OmuUB77rrtfzEOWH
xWEHsADLJS2aMyy8r9GNQlkwmGOZngYTpkzYVblz50ILHwvt7YFe4PSQjZeBEHs0
uzu3rNgizm9k+dhwGnDtg3Rsy3x94+KaBL7v/lfspWyc8YwMcBMCS4gnqkJ52fmn
1EkKs9wuZOXAdwvJYkrjIolT0skLA1R2ia6SnH5ey8LAQb+Se5DQUthhZHlfm010
A6nXD3bfnv4e4CpIkZ7DBQhEbksrh8Jhp+94fGTJ82K6CjmgUmxLwTypE3nM+KrO
bzJ5Su49aJlP+OkbsdqeIzasfZaoIJU+SGPC9fnUasN6EdZg9c+bXcyCRL0/jXCA
oY+2ezOMNoVKpgP4f7DfiKzVq7xoBsJaVx6rYxZOb0bTlKTyUhT8BbyiNya9TIjz
vanPsd0aybQcMFfk6ORMT8FYVe0gviivPS0GSidF0+Duj3wvo4WBqIcuu+hUmyPk
Qldu7euyTYURZ9KRd/P3GydpGAAgqfj0zYhWsyWnB+G9C0BorVGakXA6jhiPVZUS
ET4nNL66Al4dJZ2fTPbyYtZdWXvr3CWKR1S7H1TdofGsDvX216JRFJt2CkgyL3/R
RbBr1phKDMirYWn2QwB6uEmaryR6g0I2dPyJEhxGTLYm5ggQRfxid3IVVLF40uW0
Amazz/CTxUU3OIezpLEyVMyjOeoCnCi5SCC9VNwZPsj8AZN3ZkJRXiPZ8KTiPQqt
56GHrVMNf8G6KcMkpvXGz7HS/ltl+URMHV7Rjpcb9ZwGPMYcWLS9FYMsep/ICJXy
4iPt95N5TcNTCNG73vEoOdXik6BQKtqCjbUrnBCyQhh56ks70S/kcHq2aVYTzFuW
IhK7lNqfWCqxOzGBiHn6dRmz4qLIRJgNBGDCXilv0E4H2VcRyUSz2Kii9K7ll601
28qWHxtWrcqp+65k7aPQWUMcVySValFG75sRDX0pvYH98CA2DAUFCE9kkerM//AY
nugzJ8ugB2g6IlRT12jc/1WA7Sa5xO31Px1cfCLj7oTHVt5lojBtOeoNBiYUzzEA
t80pTpa7CWeEgqJ2EWdaldIffWdWnuApEk389yfooEgIfOqSUPjQ4SCqPGmXQBSM
wl8L8cONIV/l5jaoC0QcRUDWNEjz5c3Keli4u0m2e2H5H2eg2ZwOihGZlM6VQRMO
LdZhlPDJUpihCU2Kyd/0aEbdhs4D70t+5vcHGUVAHUJ1BRKizPS+1AJoJjgDDRc7
0XTKefr9j/h4evciKHL5NwDsqwge/U5mHIm72ZbXVp5LSut37g4kqoJ5AQaRBHiE
KfvjTLJIQDFgCyNUV9oarZQEe/umlfT63nSumkIf8SzRPbxEGeReX/IQtDT+5b+q
gyGOIlweLWMNYY7OfF4G5spl0l5ky6hCT4NkFpal8/oPUTVjag+JGqgjpkSmPeLT
VQNwufj+JaTjXfUKxE0gAkiu4mZQcB/Bz0BZD+VgJzVs0G0kDSb6MibG9W1opcPr
kOcordk/IKQ84mXwtRPD+aRdsqTVoQFHk0EthQY6nKWqJ31sojC2b9Gw2dp7L94e
0JdzMhE/FQPQyfA74DKrXvRtOorZjO9S5euOmf9Y1f6uDza+DcZBwnlU4wTnCwdP
fWlpBmN5MzqNJcJcsLfEamRo6d8Hs4SkUGlBdtLpSd2pA4YQr7QPJfltvQodz5L6
F9w5hsYrYMFseFbOABCW1XiFCRpK5bnpHvvyhJo12bGqJViUF71G+uTYrz84QnPK
+hC8O6k/U/t9/yOUGD6nsWgTaw9A0PpOqe7X53DGK1PcsZDEBqIv2ByVO2AAuBi6
B2oTP9Kp9y8m343qvEIjZ90emeSO2thmMuBSpuQzy01KPbq4tUxZ9Au9C7t4Lgeu
YV97pwTI2MWpzYucD2HwOFHLv624wV2RM8Rai1EYrxzXQddxOpLTyZ4S2pTV1uTq
sOorWgJBQq2oWXHssT9I1+hsmt+7GRf6+e8s8Lu8hNgCHH81Vkn/CjrpCGx9VUt8
YYSYUgsWC0w/3SYjKNTaWUb0HioatrFfEuIaKjf9BVzh6SgGHLPk/DUJitd3WdCi
nH8n12nvB5/DPbgItN0DDrNZpGnqi0h5I5n9z0y/Z9CEYKdF9eRjx8NogDJ2SH/5
zLO5JMM5jaz27iQePY2PZ06g1p6a166dg3P6VgvGcQh7zA0wn4AW7JCxPr9TUlyu
GOyC6LOYJ4UORUqpzc/cx2hTsFwBZT/BNuckcnJzBlaxIkDNCbzKfwqykqumXNbS
tH+34/9aLUcD69qNMHVhe6s3CWvUpapbYF5P9ZFQ9ufzvjofnGx4Q9/WA59VS/7+
Df0QLFY3jpkVLqhLvrXMBm54qldeQTlWR7+lTdbAgaOohjZnkPZgONGF6x49nfaz
aadvzkJb/T3QUQolBN4I47Z4zr4Kj/xhwDYL5KIFCNqjire2xOxg8t0Rhgg+ES4r
o3XE46HYrw8XRy2hJkCGCvaOUpDerbI5Dww8Qx+uNvvHXL/CLk9eBxtkV2WnlxiL
2/aOJYGRHP4w/bMsJNXkWvUvD2f967Nk7AibPlhef8pSoBrxGpthfr+TJzgswLL1
4e0Qcaml9HrymDXPNf39GGET4PsMLWqHvlNDGpi+FpNto6bG6W76nbuFrI/1Mmuf
b0VBvPRJ/MQu95ZuclC8Fiv2nC68lPw6AnIjJngGuD/ElBS72mB82rq/Hbev1d3o
P+DXBwzGhGr1XBX2z5U6ZtHvXZoExDqhq637xxOYdzTmYuY+odAywUfBufTbHnDj
gRpm0EReuqwG07qDIKHr5mv0UZQZJW8wI2AKHeaXE2stfExi1eqysE1ad3qKE176
baoZjpz1dg0Nu7Qus2tDgDpvm0EsxXrW686N2avxlZh5HcXVIZCtCdahNuzJ4WmM
6TDDqf/r5FGIEnmeKRQ+MoHKhUYWHkFBr4syHODZA75QxDkLIIxBQaX9EoJlArtm
QDji3ZsJqQtQhvA6xoJ7jBQ74USoj7EMcBHJTMeCwA0+hppD9NA/3Ae3p+6HyFMe
bYPpltQATFw+sZ6DSzFesSK75Y4+GiEetyRXzN9BC0e6B2bjFj2fIemtDJ9jTRsh
2rTrwIA0uwfn9keelSrrZCXmdxyn6SFjUaSiSBwYxkip3XcgfY3d7ceAW6sXTjK+
cXHAnmNiCDZXQ0XM1KKqOH4UJ16Y0Y+LI30iwjkjQDtm9UG3Ye6cSx3abvYO+Spd
Us//zH9jWEG0DBmQLeQtuqjUF4r/fJ5VVgXMimVNs990Aq0/VgHJ3Y/7S5r47BA0
HboAvA+g3rF0iACcWYxAWhXmZmzTJ35OdK9rHOxtGBxcEwsjsW7xJcif3kddXJYz
H/QLd1sE4xfkigGOYehDno5lDnj/HVBNSAFO8IM4PczX8fLPDuubaqoOsbi9GGrR
KK+WytJjS+7NK9eqSpQ/vH948fzE8mHvfyQbgxC4x4W5al7CLKStb/Ip5syN8yck
vAXI1DIKQQFgSCjrUR+o/Xv9qyoqqfBryw3iwG4TCsha9eNlrLsWOI4D5gYWovbc
B53qT8OyjlOiLx4BgZGsKo16f1UQdTMTLgiXcOUnFKgaSGcJqda/Ncv8bVqbBKTe
WfzpTqonp42YIYkjYN0mFcZ/Nv0QMtBGT1eDJjJXQTvbmk4pKabSeSLX2aB+CRRI
HGumUkMzpeqKiHxlKVT4iHzyp0O5owh6BvEq8kpaqMUongONwyXWktPRfDw0/SXD
9u/B1a61XUr9wYrchWc/pdCc1GFa0LgevIZGnPchP9uSsjdH9OEuHCtkVV7gJj5C
rXzbJE9gygDrAwjPim6oqBmRbSIUv/hSnrcv1DIeWA2n+zSwEbNtlO3mz/di1xwz
U/Fi6FOYi2lZesGpeqlBNyIk0liNIjhPaoiqOMA2W1yNWmSCNl8b75MwNh1GZdvJ
pUalgPDtC3ANpYXXMyku4jCAE648nCkD79V1g4n/1kDK+fLWLEnth/cC0cie9JTF
NoTCKxdSR+qgX9U8oPhi80F085ftUeDkcGb1gatnVRPQGzOYt6+GdaS2rBQVRff0
yrGDSa8c62rx1ev0AXOtjV38WnDm9STfYtR5FyNrb5eTalE4FHVZ01mBcjd090be
xYq3rqU6iJWVMqqjzxTT6WufLNAmFj9qnV0g0yWuh1rrGm5uh/lAxloR82+Y5NhV
amSS09/KVjcxy2bOZYNZfxvu5aJ7gF/e6QABfpIBCMGijzx9DvMMI6dpKfo3ySD6
vpw2WCKfvSVU7r0It7GWI1BAnswltmuUtGxpqJLbQ5Q9sgzYDHwUmlu9vUyAupls
mlFjPCcmexWon4guEDXTImcGC0be9FWqvyKGcDfgeWFU3QXmpmQ5LiiInyPQZ7An
NRMo5Dxsi+QHgRQDIHMlRtED9AP3wjNBsd8eD7UOVZ0hJxNb37fxaZULtNyIWEX+
s7kpCcl8rJP6x8yC5tSfglFyn+WlONS/MLIV9ucaIzfuafddrQjykkj4vRstKdk2
2UQ6SH1LNr8lt8L/XJ2rboxlJJgGfDX5Yuwba462mKXv1w6qh2Jm+jMXTGGEeSTp
qmvq/1iwKTGPhItWC972PQQ7yZIYBFsRjBMWU3Nc52YE9nqDM9S3nIJSPk2lXkYz
xW1WapN8D1xNBPG2whlPh8etmq3BG5JjiRVgZ63YbqcVMQDf0AH7HYSTZy1WocJ4
E1dNrF4XntVfnFPGz1QXQ3cZmAZSebyS8WO5dN3UnBSOyYa5K48DHGjoEExksic8
AlqXVSq8Clgr8a1/Q5LqkSUesYOox37RmWLNbgGVB+IBsyK1RXtnSDztsooH4XKD
C955/Uou/v3Btbpgz7m5ovY+rMsrHIU7KOFLVJL6ZP7t56Z1nLeW02CWMT3uPgDI
GFKGHaShCZ7EgZAJM5MLIw49PlFMxuSlzzU2lOcOfwLIp7b75KnjdT1qBU6Ni8Tm
VsMF6HHcyuK/niMt6bVCNpGIQE+eNOzvSH+Y9AEPYGhU5i4cSvAuYIeFu7sXwW4Q
F0NvUs0GcUvYOPmRlidDQc+X1EgD4gDyQquw0ymeqSM4BvoiUFKX7kylLweg9ME5
utbYXJ0eKTWZVRcbIDhiTeRun2FpP5LDrMsn+tQpf3oipI2a4xQ7QqtjOgfzUCUS
knwYiE4k+wdo7hWiW7EzR57SeCv7eDPFHXYkdghe5N5bwiN1L6AhBsL7PVohFQ3Y
MBDIYfmT/hITb9M71QX6eVW1mqoEdp3MwSz8crWcIi5pD7X9jtmJOOtqNSzrUOl8
xRm748RNBLbhhX9qWd9GexuYsuBjPJXzowE2doUik3YzNKmwS2dtSl3hIMcFr0is
mxUH+3+ZJYvOVlB2nCLpGny5NdE5DrTxf6J/tiizR7F4+6+No1RQWRU36aKLkerl
L5WoAC8h83tzncpO+/yVM2gqi8yostuaFe+z3KqyrUr2XZPVhrHHn6mGcC18Qnfj
DglZn2QZM5XrKlAFPu5cMWAVOxGR5QeRTq59zqQpd/rrAEf8Sdy+O7XlUX/6l4si
OMW+P943cElfk0HMffUCg0EupkZha042Bg5xjOhI4wJRnUDYV/mdrIuefx6FA0hq
nw6bOfEbovWDFuJvZOd7GdMnUN9Vm1ZlXAmZGbLz5CGlpMq7jY2adp9XxseBYR5X
aWktCsS9QYTPhGZo5OPOuK1bm8R7os/+aAQ0VRXhVcykLOI1dXwP0SUZ1i6FoQx3
NSQQdVuAd/j+bEaCyv1+FeQAH7M+7vGp/8ZOC5sHvs8NEcRVa+RDU+shj5UyGIsu
lmEgb//mwlUvBnNXoI4OynvZ7eZAMLhzfZntMH6t2e6ifumLJBS61z+/9CeH85UT
sO8q7fT1ylFWGff5L6E65elDGmSiQtnc0N2tTEMp3zLXO9oqu3FRL32EUAJY7aGe
ZsDF7ruQaPim6UPKAGYHB/ynqlKqR0QfpeQv6/963k3FEta+akK/R8kSQg5dwheS
iwOTpgQveEZXtOt6RZNIEmKj545/2MgPCVrGtNIv/7aQB491eTiBJoc4PbuolM48
FscMmRGWGLKeMx7DSbcr40jatwfqR/5hWJAtJsrJSyEJ3bRo+iruzXOOk6XUK2jz
Mzy8JW03P4sZRd++peFNKbM+vTkbgf/qBCjje6gXKbcEfiHeM/18GzLOTBLooQ1W
qbnP3nm0yUTrIfKuteLdwwr3z4ZhCLwPl1gwyB9K+JRXl2reTFLWOTvYUnTM/jIk
20uKFKSp24/MASdx9fruyMqmUF+MyzDImpq2N+aBRbabkCZDwuPSJKxsPTIkpLI6
vmLOodyKiAv+zmArgaSKESpAUOa5QOn3z2d2a47LyLGMsDMdtb5v9qGGCg+TTOwj
RZT66hLhlG0PoZqyfZizrTeZ499m25h1Z4u2nXjb1vkm8yCjZiYWSY9DCjGGnas1
IGg37Efmtgvm5trj19OKuv9t9+SxFj8MaDJinEmdSuJukXHqoFzNNPsbS949a9oi
jcZIwDTIF25LLi+4BmN/UgLd0wQ0rqfzX8rYs+UHTHDlpyn5+N0872EB6Gb1jebp
KjgEmsxcKY/z/ttGcXvi2KFI1NOu4FzJb6Eh3LKEU/0qpR4aUxnMWv/29R1gnpyY
rLj5uNO358Mg2XiUw+uTyVcNktsY4mA4puRYcKU7YZBDV7/D8BB5MaikZXAbAgQw
x5FbApjx5mJg5YphehgdHOsz7pw9Hrte7i7ARVitq2yPQrbwa3gcLVEFblaQbwoX
NFgt4Cl0YjdS/NNotAfXbtTPykrDVidG7+325ypy1ooK6neDCJ2CoPb0Ca/8Uym7
cK21yCQMPisZKk8lZvoIIsYDZO1MC3BSX2chbfujOB5DGK5nWIz77NhXyx0PDIPp
6mc1uM2gMeZOIsM3Bf4WiuwU3P7Mq0ZbPXpyuiGLbhUWmgVoerT8IRGTBxGX7Z2Q
OP7LqeN0Q/013PNcwWPttPd1lkNhwFx+isRleHoAU7uDaXwMGPuWRC1dFgb4mzoM
aStahsH4DKAmLhrwLYYoGxnnql3D+JhboT59zm4wFJHfh+bQ1bMA+9ZzdTYBovii
rTnJsv5nPY1dc7zZ8ZkM5N4r2C1W6jPo/rzvJd74zXN0+IMftZzyKd0kQJGf3KAE
CFErG+MNUb8pN0R0mE1hP3nV6vwDA9fBNcztqnz97oABdpVAIrT4Yk1j8b4BxFqv
YOC2fQDPDmaTnxe1Cj/MHHAJhT/6j2j/C96WujGZSiyjLaevCZl6S/du9zfcB06o
IUpuqpWHCWyLOjg1Okdy/iFtFsJstbRIoNvoz4kD3wpOXDtr2wGStQnCwFSkqB0g
H20rnZXQVhNdDXXe/sEEvPud58ymyRHH6XxjON7lGKEryogHm5/EI1zOVkaw3NWv
oxrCY4fDAkCCzGmP3JpWmjhdpei2eCvMAQBmzFEbFHp0Ge2wk73OhTKXf6sCkCKB
Bc/EWKQ0xOJ5Oz4/WpiWyOfGfC+zvVXlbzC2Qw7tciPJd7JBp4u81trRttV8k1AT
msikQ7FF96bG4WCvzdZXK13Ox1vMiAF/GJaufAlWz0dK7bl9dhE6uNm7PyP70n0u
F9ofXVQeNABldJ+H5AED/DUkaInRIpQtJ1vWkXPKKAM2z6s0GksFQTd+kLKAbAc4
dFGGoJeDQlQGwXyHE/mA1RL+XPJXT9wzuDb2KTLDFZinySq9Q+yWWtFu2zeMRkbA
U+14nlghAoeL5IAhSojfaKcyi4u19Dhw4xB8RwHpTvaR2Ily0kuzVKHllJlfRm/M
xReoyqMK4ZH9Gq6U/u94Do/BwAMIS+FkZUcrFXw4K5tIhxtw0BsKVjvqAE0Cmo74
Ty8pR4QsVXsr3nPpGtaV+RgAhppgyUrSWnG/kStnOwKF7qpa8OxnuSc/WtIMyzcP
Jj2EwLcyIuIIlMMb8y2sDYEhUalzEJjxay0ZxN3BkZlPdOiIKrut8v+zBZeBRXEB
hJQuyhDaYuS/FKzwOa15rH2Qan4+JOa4guzEF0hCc7pbJnsZm7Qfd46BkgJXGr40
trFYg469ckiJTmn/qSKw8H8dNhtQ/JXwcPkFYkz1QvRas6GhEnW7n9mKlJNKY7Y+
ig/s9n1Qo0759OCJOjxM4c0HgyIlmJqVmO+c1avwsTMnd1fjlrZwOSyYyvTXHZgw
EFojbsiw1rr8QAUBxSWotcVCPAoB6q42ro9FPRFd5FfGtX5NoTxCJc3gxqa4McU1
jw9q7SidBmbztZBg+1SwC+hnKAeQcNNYvPMwaULpfFEU5D2J8XWl2YYiboKly8UL
dkvJdwbg3akNljv//fC0RukiOIl4CqXwxx+rGp7DGUtHXsZcp5Bdim3HOwKwnnAm
zDI+Nu4gJp6hAMRHAv3ksVh8vix7EFCtHXtkVxjNTHVN8Cjozo2V248bbkAM7akI
cWzLJis4LwL+e9Y+TibLU+9O6qjREJXy1kPgS1kjAZj2fZ/IODHSKasVePSNc8SB
qPj0bPqXljyMPNbNZt/vTcITrM30ri49gauGFGE74cgrmMdE8R80kOYBaV8dPC8X
5vx2cAxePdXlaZlFr6tVkFqDJb44PwG7QblJj2/qVaArjdmabOuiPLOFf75EI4P2
TvEG39u/lReBjXLL6FTxyeMw6Chsf+jSGPSGOXS6QOI5tHBpxLV6ET+5XftsgZCn
WTvzZBE1IdI6/ZC9z1zPn7o7w0iBp3Xivr8z5BQpOPXPt3BuPuupZ3zAIVKEfLyc
GTUn9ibCKvMuScnsTr381DK+FHgaOIU4A9EYNQHmz4xShj2j974gBBsLrYxmsz5G
cqiaRrYe2jaU6CEFF7LVerPseuJ7AMR84UlY7TlwJy0MAnAf6m+ZwGbgp5ZGeynT
IComcqPihZk26u25iB+ojYtCaTasceK7TzSLTqpxa7bbEFUoKN8HfHr61hqkDe1h
sW9BtnyqvOEDXLDx62cVFJ63VwIwHtR9r3ADEr3HG0FoiCJc7anQYnfCkHRkvmlV
jHXK9aQKYP9/9h4CxA2SgO/2ixHmb6Lklcvlrj+2iqR4ZEnsR6c4ApluHttgMzuZ
ALd4/swHphA4iAOYWhAnKNpViVRV8oxc4aB4X01EI0uTaXQDEZcddtZDRZ3miJbK
+Pw61tBuY9Q3QNGLqtnZjCZBfgUgCW5IorbwdFzuoafttK9qnzyarCZ8AwMKUhjN
1C83JSSma1tXuRSIIBvsXkzF7TjqE7a7L3UFuCKqR98mHi7K/7o3iDfUo0Msl/bK
kdxOHeB0Har4IzfN7/qxBsKzvKz4X20DcN+CzBRUWQeeXflNMWPG3r8lAGRMdZvt
nGGNKuH9QgXZ8omPlk3CuLIoPkBjILn96TfONq6CmtFFet6cPWzacjIoVppBY/A6
pIyqtkliW4kvU3e54Tr6K1SUSRSnRX/kLYqz9qQ78TTZk1/2v95DIQgLYSHSn+Ir
CLKCmRKd356DwVpivkOUcUTMRGLltBcpy+a62VCWl/2cd56Bz46zMM+5HEK/iMUu
YZ5JN4WvKL2gvvqcUakfuNnKZnZFcRUrTaINuMm9kWMmbJs71maCSa2uQj851Dbu
i1QbBY2tI3t2fZlLrj9CBFpoDVAZ19tE3IZufehUyFXcpugmFLqkf3Drujqqhr+U
FOxpeVbJlsBtEPEMlshIbq7mw0u6JW0ASK45lZfFGopxqgX16ckUf+pA31v2p/gx
8ZAPJ1StDnfXLg3kVxFDmVNMbfSYkUwvdgEVJDrr62Zppg5Oj0+692LzNPO5ZRfJ
9RdgRfGP4CktwmDChrIlTmq3CezCueIhk2N+/cYuIST6JHV4QFHTr9ozDrd5H+Eo
dR2lf7cHrhfkD9czQ+Izy+WKsNAWWv7U1Ki9fPjA05Qsk0cz/1ys9QzFqTv4zA8b
RYCNjBCSQUkIxjcWy0pqcw9q35dmUshVzabQx+7erUkb5JjCtFD0czTXcTFs5zMs
3l0LFj4oPoqYhmcs1+hdPj8clpsgUFVaWKi4n5DCDH63Cm+W3PlVS1BIyIYdurqJ
nQMAEQTPFAKeCK1RjqxpbuS15gnfHP8WUD1Dj58E0iTsF8yiga6QAIBN3qwJPB2N
2uVK9sqUu/yUpqVilPE8C5Lua6d2cbZ68eweALDzTJMz3FujixFz+aKNcEJraGGb
k7t5aOP9Gt+mOrSxQcIFPDxdn29Ll4lxNHiDrC3CGhcA0fc/n3lswIfmfzofen+L
UXfjdlMHmjvdlQ66rjBi0w5FOe3zKn4Akxx8WESjOxzyDVmIJowq2ajnKG0K6ojm
rfeHdT7ICQn/sWD1sdHhtg8LdDQlMc2QlaHs/pfr5SNedpEz7mPbSeX5P4inMt31
7yvVwLvhxtq4rAldvAZoQ8VruT50e/I2SRyKfbKzZvOaV/05p4GUN8jOkeNYGdw6
tGY8eusd0DTPmdGJ+/yPo8cCv9jgMR75d+ilI6DAM112X8BIcaZLibEyEuUVQ4Sb
Sz7Mn3gtpdTfy6swIqZdudYq2ViQNfJf4VhdcB+t+gsF77SD3u1Nu16ZU3v1iaNF
5HRbU0tm04hdcGRfC7nfkEBFQ+lfhdRXq4gjYLATrd6FPoSVtzXSdjKtNcZUT4Ab
bA1doQy9IcoU7EM/hC/y6E8FiodiUkNixj0cSvu3cOcCVQwnGa+Lo9eVZtJiDdZG
64tCVoOaHeYVGr4ZD2HK8BeRVp5YY1DGYUBXZRDcKYx+hSxk2h/YF0GjFBBajl1e
0+9uHfLRVRg8WmUxWMoAs5Ef4L1rUq2Ix0ZpBGkb5FIunX8PYUBU5O9a1km6jkqA
HZr2pcETRUa+nh6xzNJ4pxlJSx+M2EEQuprW9oP0y9EFSE/OdIz9t2N8adZxJpY+
QYNI2dgDY/LWJrE17gOQYPSeKoSF1xExqu64WMaphXcqkpANKFb08fPobO+6Q4VH
+KnnBtDDR1aeOlhWgkTYXUTbwJcA6ceI9iXDLcyoxCqVBJAOiwhFX0St7HyGcbtp
hVodO0P7jHDnbxwWpniDNz9zIMAgp6yn5NF4GBEr2i3l+3ne5MNS9VX1P8Lg3gNI
noRg9v8uOwCn3hSvH96cis2q5v4n2mv2gWelMP+Gy6j5xVqOk3BeceAfO1o8JM1j
izRWiSxBL8tcsMOliM14xGCPQSIJ2lI3INBaEdCIQL1diziiCuWao8jEZixBtUR0
QQHVOF/CwDpqp9ENA55+dwqZh/1aLFLN0a2KwOi0ZFUdJWhc3K+hzcM+G4pWbeYY
BmJGZkQrN2gN8stMyo71iDR5NJ+WiCdnTvKjGKGjn513efgJcGJmsSYHVGN5JJU2
ABPuFopFOuURyqOHXUXEbEn8liGrsPRgiQKJRUM76pwXraYQ0WMY4w0qZOPbwgyo
sGlKSOSDEmsK0OWZDhlrT2hVfU1sr7rCZ+zG1BwQm12OM/RFYfqQUvHxqgDvlYda
o9Q9uIT3UJMgqwLHdxz8o+wP6laZTbVYAZS0jaeVyS9grbSCjvSKaN53ofVw+43g
iBS64tDg5Z0iYzTI9MpYu+MnN/jH7iNXSGCdNlafColTm4hUVxQ4eaCD+6dHraRj
LKIIwAi/RUm9wdWuAm/ApXQguKwGV1qHufHvr56Ph2dHHU57mxvQmMTDWwKP9Jif
gw5Gqo6UZh/cEiIc4mNxRLmuzBcnD1kFpBjGatxpx/a1cmqHZa3gYltM9y+9g9Ro
GTkxatqgn0xh36vYXZfNqu93KizpHW+4q0c+TU5qpcL/sABZxSGQeoPhq/KxoP9Y
tUi0gegvtrHkSp+bKQoRPO3dx4aVLVXiVeKcizRDieF6ZxePtvXnAxiDQ+mQDBFt
umSDUJYlkxbR8awPweCV/MVqq6OwXJIrmUS44fTPWR2G3mZMFUQ9ZImAuzGWFGrD
aj9vpqSg0M2pPeA+wJHhLPumOZudSn/6cZIrsOqP+2kmb4mKpz2GNV1qhdydbsY6
Lov9AS7fZDJp6bOO3v9WaMFOVW8M/4tjxQ5ywQnWmfXu3Ay5Ktrm7K5c8WvgSC84
iqtzzsxmRdkGYW1LpLHhD+ikNQI1wAccGRYuvU7Gqm3JKRpFIRnm9QvvQPzejixd
vXVNUAa3CxJOAK4JDstx/fKclYW6vvDvXiGFmud55+KT8aIMvlkGNRAU/G5kHH+h
935BoMfktTW1GZDzpUNo+gpmrtvSj3LvpIRUoJ2dVivMG1KyjZFU2osDDiUo2qTj
e65bVEb0xeem7JrV0ceyhM1fHykR3sPb+RAFX/kvunvuAseUTnS/A4hkqwfjYXZq
3jnOAacvB4yymENPQvVWQjX2pEXx4ej04WKcEHzx77Ei5E+g0AfbMlWteKI7yUAW
xGbVOy6Snija2rHsp1lrKggclKFwBDkoOYRBrNQEan0Vg/BsYwFJOD1ZrF9pIY5H
XaPi3byMxWq/pQIAPboDqar6FRUMtzEhWMIPDOtd8+ct+z6dbWcieXLDxMBG6UZm
jU7enzyYVJ3EIPi83VZ7CBoi4koZpaS240lziwoQiaakwBXINLalZGS8MJSrE7ow
3p3tg0uJU/jyGP0LvrPtVKJHB7nEafX61uLJmxSuGXx5zVDCmcXXPJDKuNjuREUV
zBkjAuXB9cHR7K0xdEwhA+casnBtNEndh3wovB/2zRUTk0nHzRgH10rJaun7mnBK
1XE6JLWQZK7RsTtu+cH1sjD+Ac75P/YwtrtF68dMIuLOZaAzsOoaUQcjJiEVhr2D
7HAyPW2IXJaXvXlafMcfh++ylq8H8haPCENBMOJR3Aaf+fajEyzNogC8gc/eWI2s
yLzRD4VaIoOVKxbgDcvEr/5tC7uja/DInJEK4SV7tyVSzR33CCNz/1GPtYC0gc3y
TRFHDutScmJfazQdNwNu0Ml99Gn725HJdxLuxNhWp4kkmIy9BNVZ4zp1Ac+awVxJ
+2+ia3Cmarc/5YVE8y6zyT0Xij+XwVTrhxdzT0J9kfKi2qP5yGxMrqHDbktrWM8h
4iL6G34nY9I+X4lvdTg1eCx1EvqkXpn9VNyaJqLfgt9gPTDVuCmtSultmvT3zZ0R
4IpR1RGP1jVy0IeoHtVrrq4+kSj3u+EhMoSz3LWrfwgq0Wvs/4R6G9BY3/Y8HwPD
5MImJr78U70ZCpb6SrsQlQY3+RyXc2CrVNwOOWp0aZzDsTw1p2pTh+69ABbZVAyQ
dL4VYCV1I+HvvIkacPAtOOAfq5ZZQ9BZVcaoxjSQ1Ld4MnjWW94qsFp5goycyqA7
exqhiEwbNLNLpgRI8l5FQ4DX1c3B1diFIaS2r4Gmw/Ekutm0mp+eASwpMkzVU1DW
AMYwDMiJ/KfSVspK+KHPpbL1VHnM2AVyjnzxOeo9QU15P9hB9nVjv6MdyQyaII6t
JGGUXiwDac5qOOecYwoXgBFzfkTEdcY1Da+LuFXaEQdwVUkQN6O3YYfaATyZB752
vSlJjT3Jm6CbhMFYIAhGdG8U5A5wNLaBIql00Jzevvs9T91jjgtRXnlqbz/Vw2KJ
c7w1soWF3+749Fxl1GvNUjFVwXJYaxLXhAOa96+Gi6uNNR6f3tAgEObsfApW7W40
OeXzPemdcQ/04h8rZ74Ud05+zX6c/IuCJInr6uyWCBbud+lBt4fIFjOdi3yGXrth
BPSupqG9AKPECtlQYDS58VyW3xqPT9Oy8majDXGyJLoPsqeWluBmttyzAyBOxCVr
dh6aBO8HmAgH4Qq5/gvZRPpJL3KALOqeBn9GVlOQTxNixHJx94sxkcaFO4WBiB6X
US5abG2/91nq8BrhAFHGrtVNxW5lEyqAr4AmfDCRC2pBKOqLg46nab2koI5WbWKn
jutnM3Cs5MhGZa654koW2f8nmF6obIe7Zwu1/6MDNDmTBa+ljZBgXG4eXvDCIpcd
feKMX0rielNBUAmQbDzJGdKDKtiKSDJj4UmknTN65r+6y0FqXYQ5vZwaUL2+n3gv
QO6zQOQiGw2U1q1cqZmPaiqfLnBVGif/UDGHKH6PokBaTZP2VgH52rVvr75aZru1
1XqrvVDh/4MCYv+cZB1Eed/pOGCEenOE0KrY7HbysTexObhIAg2h3kswDETCe73V
6FB2PcNITmx++QZ1fDD3uH9Sex61V0NlLP/Xyz6ILLELuyyQwORH0ttXj2uCFluk
9IIfTd8y896fDy+lxwcS4P6SRgsHcW8iPSG0bnUHDae54zmk0YoBA69ExPScW9+p
wt8LIRiW1sGb2ayTROXMbS0pdxpDWTSwe0V7X+HX3MHxGZ2lNn90SqNVtjFxXDi1
ngYyg5+hRA5kn+cG59cig0qhKTfNnSx0TqCO/YsBR+RS854tgWX8hMAiEFokSI38
pWSPvUdUntp/x9Ky+nII/Gogn3y0Yq1RNyMPHpmvd8wjJF7jcKEPZvObO2HyuoE/
0+AS/KQ7VijrcMRHppLMVJlo1AapxtClk1NT66VrV77a1rvU6WD/zyaNcBmLmlKJ
1d/ZQQNBwttKOLQPDQWACMEmbUD7WO8/CiiTbjxVAG9VrUcfdwtccorI6UM1+Tji
C8AnQihCkaz3d0n/y1LOLqhVoSeI4fDiFF6hEVTCEi+WsCM5XrZgn8rXV3r96IdJ
T9PHA+vYXSqnVrSvUXvM35FDdM4romkqeOom/uU6EdS3GD+c5y+oPrgj+sIDsMv8
YxinVRj37AD0p/lYbNJSsRWzLozxDvSIlSgOZMJGv2uhs6O7iODFJsH0UzNQ7dWB
w4gjWg8SOM02vha+YbUljTYkrxFcQhKLgZCddh5u/LqItpUK+zbAyWJT2SjK0nCP
eXMo5kG9mf1IpT9pbc4xTM171tFacrahhIMGyMhDgZIGOjS8U/wtIRHK8jrtUnPG
kLAaQBb7oICxHxOuBG7WRrjpqvuRyDX/kjlyW3rnel/rfyZ6qphbDC2aHJ6TPZmH
jsJbiWFcf/kvslhy33bT0Pv2ek7WqTAOF1kRZOjzdAeDpCQ6sA0Rvj8cGV3tkkLs
cSfK2nXanntiBpiJw/VWVaIvJsS54ee+IoBY10YqRWeSvYabo4h4tvxa/Uh3+8Ix
DgiL1aTcWxo36N+Zpj9sUVmdfWx0ieU0XjogTmxgVIkgXFOPUjBkK/UJNHvxlOzm
9LF30X2MfNTcWF5xzsEur3t5r40pcpccmKXlmQ9zZwv1VP3DSzYOYXsRZ6ovzm0C
rT2K5sSYCLSD+4AWfqsbSIWinBEXmIIXLkkYl77a0fgNP45UMtP/q9ZM+rGr4Eaa
rHRlF2gbjQrfkz7SWxKRySQihdQPLpyWP5NOq726r0TL0fi+BUOO6yOFAC+GaIrz
hxXjeGoh52bPkeW63T6LdayuM8Hau6/TiBU/5nSAO8fWw2QUkw5ZWDHZL9RZV6Oz
56jjclnJwVpCrk6Fm33NH4RD1QlAwjOAjFPbNbi+/IcnFAmlEOiGt0cjAu8ux1us
zZflL6nIi7v+r1HxAJ0MnOnOVFcB+meE0FsfgrbyGzEMkDSZE5MrraLQ7E/Itanv
F2rJANJWyGJyycZOgFA3UW+vQQ6vq19YS+dVgWlJgd2JQbj07ohCCsw3ZMMsN4zT
5U1DZFn0leeBjdbvzckoxITt80vJBgQgx6ZW1AvqgJ1Q/Cq+keMtAVa7Bxw7mT8Y
favMSD8q5C6vrBgxu8dWlZ1tM1OeQQExXdOO1nNV4bqav19TWbO1/TJUIrFwupCV
z8/eB8ChKyaniv2XruzVnYQ01KLwja5uU+WBLPNcz08fh10en0CuJ6yMZm6ct1G1

--pragma protect end_data_block
--pragma protect digest_block
OoB/xz4X//ABHHN74cXgeB76hts=
--pragma protect end_digest_block
--pragma protect end_protected
