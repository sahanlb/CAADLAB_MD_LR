-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
mIokNtZ2t2Lum2HVqswipTghQBDKYvCu6XlsT1MboWv1jK2dQzE60Q1NLtWQ1Sb3
Fkv8Slj8AB0IjIQLBQ/aOqWEFX9Bx0sCGgzUdo0opGiOjtyqgmTBxFQ+bRP8xw34
QG25RCpBw3S9Y9s6SD5JWnEzGQI2GpOA37keE8J7OTY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 20095)

`protect DATA_BLOCK
VLTQVa0Rvu1clPSWxbsnnVcf8d1WpcbqZ1sjrTMDzQpirf2wvhSIq/GLPdyxGLsi
IHAr6aNWYsQfzhJMIJCJpwD7Q+IsZlZMkNDCtOnaK/cc4IbngHQeb+5TLQHZ7D2v
237UBln8bUGEErrYrLVDESlM9IBlvCq4I1YxBCmNIYbki312AT1nWP/LdFkt3p+4
Db9R7G1QijhDFAQ+cq3lJxVEgbWoEcqH6M3C4jbj0LT6lczaVqTwfm74q1L2Sbcp
KBGWw7GuHKoyS4gGwIjQMdSF83R3YLzysJsjZFTPZRepjaheQx7Oo0YRnz6zi05i
G2aNUv3E1L3dwUPDpWvc4aSDtSte4+BfBuIIicaMF62J8IcXv+G++UvyX5D3HuMy
3jkWCz05jXunHUxj5IWs8C2D7fjZrkrna7QjVPE2d/J5xhlSc0tLSJWrNg1sSzqR
OykG9ED7A62/Lm34zWGlZ4bYtIyPDyP2SecfnRo9/+DXCdA1SVp9MX5tP8MaxKCe
873RsmvskFwuUR/f80GHD+XtzAsTpJsGqnYGy3mHi9HzHk4jGZA5A0QmV9BZXY4e
S1h8uH2PevoClxK4yIsoUdCWOqWseAnCeeKdkK5VOC9EZmcua5QTv4Un/VvNC/n8
tplYBzrjk6X/tz9ZoeXzVcHehncxuu8d98W7Ns/gHZJywrV3RO1Zypgo9bkiSeLj
H0yIBPc1Rcnumj2XP0wdvWDma4aHnQ6ih54qxjg2kQQeLRmwp8ztu7uG3QjzPH5/
9+SswGp3xUUcbjW/y+VYvqyzW6IdFM4FYm7Zqo5Qo0zb8D2lJnT2Vi+kjJidK5td
f6SFPinKEe7OAe7wm364XDITyrsOZRTvsYcTRUN4ORkLHh7NuGrqMZtMkAhXkh9Z
A5P3V1SJnNAVrL7BXnJKf1JlHBkSitrH2jX7icUCV6J/MkOizzSJQOXf+csfaugJ
1yjuuFLAv93ZkZhG5FBnOC1RQbHF68LXsnm5MTiSN94uHwOKfQuGtQjt/PTE+Qrq
dK4UMb87J11SOo0dazQ2R+QLMAN7Fh7rsIRFMdIO428GDOG5CmhKWTiqW9YZerCS
M7wCSx7KbfCPM+RqKOp3I9Z/C4x9XqQFX52b8lkRz7M7DhN0wQ7woUVsxezqekQH
j44ziR6wrhem/zx61Qj8OysS+5afvLM5dkEi+ot/c/ZuqJraQLu1y11FolWGT24g
69QYt5yGTRaEkiosROmfPPyrpnE3xWZX8SzJvCPv8V2mMPHsNG33tlkHzxUAfDwX
ubFZ3dEuUFt9lKGaOLb2ETWlJvadAUxGmCsvqztpFGPr1q7+PnECQA8z9SNTeOT8
15as+fXimqti7+xc0eI2SzVFBjIxZblWR9rorSQ5MLAkGXXVrAJIlxzvoYiJvsTI
m8m5BroiS81xYakp8CmTzHgp/17GU385auajDUo7bDwDQki5rDfry8kQivTlnfeX
2gsmB7ZN0924wePsqKkjffXv+/oLJS/SFbww0cLqxmsxlrcoS4DmHY79PrrsxCd3
yKrd3geapl8SgN32YvdzFvNNcHljZBvDffeBz5ER4YyppsnY2UDQEps7vc9kpiCU
k6fL9LhFHi/KT1qZNM9RIYL5QsfuAJFLM1lG9X2U0FdHhNe+mIPre81FdZ7qiPVO
XeywD4XF5XHW0WO2TLs+ylQzoArooqn7MdNYx4x35C0PemcattbbQZvqvKS1rPC4
qqPH86pgbDkK/len+KYE+zC2mTFkel6Vsv5aQoZRMOtNtHB6JHDG/ezXsdPlWYSs
0/lMgZIlhmN60VNOznes3WLwrSpau43khDXektt2jgwH2SMcFG0EF0RB8M7ElSgN
t9IzmYXXOTH65VYBQ++iBK7rmWCOlCThsE5j+wrqkbt8HE8QiWNqUG3KutyDQYoc
jFbGRzD+2wRw6qcOGEExcXr0DImk780FG1yazAgw5Q+lmqW+fxSySx9Gfk8m25ig
hlDh2HvEEgiHt1CN3lZi981g9WnZh0j7oRms7hVc77BaxAFUSFj+yELBn78RuAcy
OgxRGTzSIfDo7qEFwYiUJhc2VvtfYC2NHg8bhYqqhbuL+U7yHDn18/IbNROROgnW
gtY2O0kmeJQKAyvrgQvQC7jevxKkDwk2tcI0lASbKR/U9Ojpym1JDBeCmpy6IAId
IbsVVY4H6MwyqZDbKD/7nszjuRETR66vEZSP/8jUm3dcGNm8XLLs1+yoUy9wijfK
Hae75mi8hAvwk4RXKAOuKviv30WO0IzIhs2W5sY8/w6Kg8RyF60sYfhbECmXdNno
Jo2XISKJzGbxJXhqYcjavl4bPQKRPeerclkAp5bwernK7PC5M769Zmzs3jpYg73I
eatsl376KjgkHrWoilHC2hP7epgp9R5LO/2wBXIxkNdgter6tsWew+QdAzEIYGd6
uadP0uGluAAe09yosSAf8oQv7T+kJgDlYNn31j8iwgPr0yAT8o/PQBCX0LOAL1nd
RlLt3F76rNvXMzKD8dV5dk5pVBGiMCKnN9QV/EXAM00XdIPmZVTv55nSI9p8HXuv
ynM07g4B29UBQ9r8F2uBoZTH7U0+9ksU0yYCxIJ6anx6C6+WtiU07a160TfzcyEo
cAnLjI+Tin8T/gv4SZwzSa1ztuUFbSlJFbKQnbqGfhdS4k+VJNiGNkWpaXCuRJMN
EnXO7okjE6CGlNKb5b2lB5yU3/M9LkHqKx9d/KSitIBKSGItIsa/2gocFKfQr7D4
pK7YgAcJeHhza3AJst4mapreIRBoMVq+4+bwB1CkafEsjU8bLZdVfe5qCTFSO6VQ
qDDxXVnvUweVXwMMoUQNjrgG5UsOec/K7HU0gX0gYv/+HGiF8bZQBzGa906PN6e2
jaf+0J08QFlk5M9tRwiNBGqBW9ga3zUd+nkgLMdjD4jwV/N73KiLQApec9NI0NSh
JzKQ2GCq3A+5HBueRzTev9k+rg5pFYA/Jc5+gzc/lttorrdycPVsPhBJsCbf+8ot
ejObe0khdXAoQ0uf5xeqo4QcfHdgc/w2xQAg0J7FlkXHZj5kChTikQoQCX32H6qg
MC7lKNP0D5/p+tbQcB8bTHt300dBCFrlqrzGBy846kKtIBTMn0ExW/cNA+G2Oo1g
SfqYRW53dMTzM1BRc2mtIafGbM1IWa8l4tKF8tYBwLzfMW0s6itTRyIimc8quuSn
uwvtuhjBtSEEluO7+1HfO37/kOWulFvjrfkMcWGpq1VQLYZ8LXERvFIuLW3BDN5B
apAtCuSz2YVRVhrjvwDaGpnA/UPIIvPFrM08gDgMHYj2Rog2UkXsMZSx1RBHYZK6
W9rvdgIrQaY78ko8ofFA3pk23UgReCE8lrg/iw9+8ZdSFuiN36jdI+aceZyXbKtK
1Ez4UhJMpTG64s26SWEMN4XKzAHp1EsmXH1aB/aOlmvt6J25WDwI3a6oBLpmxO+S
zmBRYNseu4b9rWXE5B3lRpYgq59ryvST3iPW0I6CRQ0EspXtW9ZK54avRrkZ9wl2
5VFgcw0NhLgWI1/nNkdyq0fPWtjfkEIS+N2bCEIuSP90UBdGqCKjGvuRmnaH4B/X
F6e09kbQJLYScn6sFZdcIADOW2XqOuMW0M+aGnJ5O7npXLEhuRK5C67dN5MTWK01
9HVjVe0KDE86GSZJM4cLb7FLcQO2ytxHihE89zsJzCcdam0zsAPREdXYw33K7Wyn
NXpVIJKez7gKGmjSMoj2/7hE1zntgandKiVQTXUcOqkhym7/kUqpU3tmbwYNxrd+
apdQD5YT45pUR36wgcIH8lDu6z3U+Ollq4btEiEICUbVJMp/EYn60o2VQljeqP07
4hOcCNy/bt1qwvlHA1KDChOG+Ox3CRdTFo/NADvOPTB4ad713XLmbgZg5kLS7sqV
Mr60Kurv1qb+UXiEeGsXQpHI6Xhd1K3fixcdk9OS1XjGzNjd3VPctuR9g5p5h/kE
AQBvoIR7HPt6eQn7xECiyArN2AfTrSyuqFz1spwT4lW/1OgmSo2wp32ekcIHgaEt
360QkClM77TLICK223YypLjKv2M1YWVRdn6AkzjPcS98KVv6oogBgcF/dA5KQYwz
cgqTJ9rMqGfALHVuP7R9O/FLc0wZWy6GnaCG/jPit26xZxLKvME9Vs3i4iZarqu+
C3XG3xy0a9en0t46YyIaD9WyRhMHlep9HW+CJJBMxBHqAHAaYaS66u2CAx+sxsLa
lGEmdcBX8UP0dAWVG7epc2lvpTUw8oNWDnUqf1eGMtpTmxaH3D5mqdpo3056b6il
ocn/qo/VciEBqlf2vMBVn98FVo3kal5DXdpkFyjj7ahxnpXDYW6ug2PIESda6rGm
C7yqLuv/Ay3u3JFHBoWOIhPA1e8XPNnub6slXMSsybBgkY/XNlku6MlabEvqvRRH
wr3hbXu+52v4ihxyWNin3QbKABMeDmB4Vep4Y4qaG/bSLfOhvEpmH7DG5s2NRGxL
VoAl9KbNCKG+n2IaMgw084L3Rp9h495IdZ6Xi5jEBch3y9WXqhxZrQFXABZp2klp
bKCANTajRcU3pDo7TJVvbp1KfhONCxPU7mbYYOlt56O0hqHMY3ahBpqgVyPrsPN8
bM8pJ4YGq1w899A0mJ0amq7DnYvlbOl15uucvkq/hCdeXJuniwYupwRZDq1z+wOQ
h6lwCA4/VL6e/4BFEKbhRIdlfhBWcDcdP5NLjyNnpOntRRo521q1JZkibJQdCazD
wrR3QMRjQkaID6PTxuu88XFOlxbNidAwz+TU8ci6/RSEeTFeE2hsqt7u2TWvekPE
J4QhzQvHoo1K7MG5KAVIaPGNwXTcQnkG9supeqQleGyQhk7zv4IbvRu3X8YlY8M2
O3cSeloF+Y4NyhxFCXTxexlnPwgYSHoyN+zYt+bJcCnS298vV3RRe0f1qH+X+B90
Au3y8OeWW3SMd6oOJnTSFKtJdl0dYbpxcP8Ox7YKQ6ydrvuvuN3z+eajPimjJmB0
IzEpzuZk5fjuoy2A227V3YKVX/04I0LP6IqucmkWhYegQhVuwxC1u/jEp7bcloI0
Wq+nZyjuyVyLIn1N6hkYLdv5DcAAYlSQFQup5R5s2z9xzPKQwQGEmGGK8H4hRmCb
q3GbgZeWtAiGmxo4gjbDhDRZhcBClk8ExGlaObqw98hR4GlS8EUeaKSLxwnrN+4g
NjOJ5KMtM2TKMOFB6BhPdxBkOIl3O0Uz5q6JsdpA/zT1LcWX/zNPUg4YsSgEva1g
s2LAL2bx6YClEUN6gqwVF7aEo17HaVThPapapkGEw1HB5TxV/IIT9Hqk505EhLCD
3iJkrEQfBPH2j4mzpeVk3IxNkygb57ks5KNH9DHA4gS1ttcxg/nVI9u/rcdfTf/x
OhmRm3W42I+on3bcfjPrOzC5rZVY50vBK9uyO17utPoMwAuoX3bUsfWkvO5Dmjh6
VUqkl3S1kuXLcOt3z4Gzcq770tqGI0X00KFGUcId+hlpaBjHJcFSMZTZ8AB5VnXi
Zg0Jeg04d2VljgqabEbPKM3LcS9/5ZH6m9UNpprK4NMRMnVzsda6z9zh56nA2i23
YGptq8KlRJkAEflzj/veWWvX5tf70c0Pjg8jUS/8gmFbfRAB+NLhNwL5GcA1uWuo
QvaYr5zIKei0qApVajQn6nZxzCOrKwpXoMQh18Q21F2V/GYP3FVpPTWwctEWBKfE
Xo0T5kbZJyB2AKrQpRkM/7Oq3viwp8RGO/CV4uFrD8ldg00co+rWj9ZMP+HqZDYP
gvxl1NNSh1xaVPN0lIAhw2sOgRWudTuN2C04pR14uyOO7kaanZ4dHar1LQBlTubO
cWT4mqqnU0oK0Kscr9i59hY5jRP+Y1m5cw5jTkpRTxfcYnvSyNwd8Up7B2XKIxOE
+cBcu2iRYbxCjr0sm1lZmFdP/kM8XJKF3NMHUaeZL9Z6yAhuk1+NY4o/Bk7Ll/Ed
EBkyzW8lnVtlccQ2CEeH319NEY6xdfeY9A0CfmG9YObEcXDdDV37g0uCbs5TL6w3
v4505TF7SOUBAaekztteg+vRXIQ+hRhZX/sgbAEHR3d6JWJADFEmMc+5bS0s05AV
BHerYwqTo5T9qQLaMCv6I/t+Rs2wKzGArwD0RWE+C8rogMsCaTi2BlWMt+joRYrx
TjLPhNXymattPFs5avW+pc6CLYpFXt8E67ONptj54O5tHgXicUTcUcik8jq698zV
VA8igxgxOcfXiIvroQlOl31Xg0wHMMFjqSu+Sv1nPyre00vw/t0MPev08yDBVAlY
66TlDCApbIjI7gS5y9VSTcM8RFsCco+C3v8rAyNcxm01jiIuDYmxvb8ofqe7oeZ/
Db1kpgl/6hf/1VCA3GLz6WV67Uq12oORql7BlmEmlKFwprVTdcRy144yxM/b+B2n
qE4T3UOmQDb/zMo3gUbrL37fu9RgSa+AWLhf1NF96pm5jkSZhGiAL3t+nRXK5o/f
lRDGppXsF1jsseZAa//JbiEOrved9Wa57XZsMOCqWWVTioMdxqCoNzLCLhbRDu8Z
IPE6acsEfyR06LsTT+sBw0itnYf44xhPkl+AYq9CQPlg8V2dTu7kFLO61a1o7ZJb
Rgnd6fYU2UPGqESVCb1Jikjq98KwdjP2ALbFNUD+NKXxo9BpSp9vLKTDy9pOJCf5
/D+wofzM6na0/eWnTXHNh/Lfaev4lCY0DPZjMtaijlcdy8Pf77Le0V39D0TY7Jjz
jr/Z7jSGZhtTK163rhM/36cOWKy6MJnxTAqLbni6AuNMnukHmGHjy08PLMgY3LeR
Za+XpXBdMbqIPi6kOGhkugtlrfe74DmgQHLk1uORquS/sUOBay4J/0oRla2EP4QP
R78bHKCx8/Rh2Wc3CU9GYI2VhwiyFJ9eh4TChmDwuXiY+c6bFjj+4RDm3hpeuZn+
or5YXnDUrSn7/rc1Rfa4kd0o6+Matg3lVs7xR3Co2mR4KBfmlWnYgv4B8wGohyUN
N/v9rryemy6nTZNmzYI3k40ClR0gpiw7s4wROw3H3rZZdk1okh9aKwWzexGBDx/0
p8xfuVCiwdNKAamFavx6ZBuDV/xWOm7foK+4gwysWliQaRKOh6I6jsFLp9Z8/kbu
cdrEeBG05qTZxxnIgZmjlDwpldQlyuMCUrx7J3co9SpFKq1QMhLBrp0Lhl00Tnx0
4Ab6QjrdPf0+ngjz8xfKC+uFIEaYg43u2cs3Dhwmkoe/pgAGol9+NOuZWKe6kpYU
MxhcWd6ofvb7PtSusG8ofHRb/LIp0m40uaXxZXc9EJTOo/owFMnvf0dmQcamKmTJ
NOsxkeYenDUEUq7xwiDKG8cd7cAl5enWeZVez855RslWOQN/WfG/4Wg+6hp6joTr
OWYO3AMhxbYQjriFzUjo94cjBGUzCQiw8i8oM4dvOoUvViyKWcsqqnSbJ7+FlPaa
FgIIYJ66Y0pLZWc52Z0a1z9ssA2L3c5FBfOFtgait6ez0HOp7tip6dBe5V2HfVNT
VhKmQkQtL6vNb6eKJdQqn74UsdyCsKeXpogur96Vm/Dv7ceGuM01sqWHvnEavJAi
KkG90atl/VLrIXgjhrgE4k1D8nrbY96ZbIDAQ8w7gImz1oPt6CP4+bV1ge57jZGC
uiopUi2nT+ST0vVXQZAqLnTrcbtY6p5H/w3zbMLvAiitvb0aBcItmLdIjMHLkelK
071SOfCjLP6F4Bjdjn2sqpajcuMwrIZgLcLJeoEzKA+GCnqsbPZaNKq4fYw7WdlA
/9c29DW0Fyc6bm50bzezUSKofiWVvsBREmJDfeOHsPdGha+PV5UBISlIgMYLF660
lSkSzgtCko9XiWgjjtfpZ310Cvhao7m/2/bJsHREbUD6qthnJ1xZ4+xSspLYovZ6
UnNDrZOzd7ADhUxTYxJOQqjhcMQ+4EH5WEKzB0gqhTclxkPhaSNjW+Z/RQY8pdvQ
1ei32mJ0w2htkCFx4Ugj3EGxugf9W0YgsyH1bg9qOV9LEDoEPCeOwKNlg+VuIXyp
oXIRFuQb9pBgegWGIAfuARL6e8oX1aJET2dtHyTw4Hx/FIx1SLZAci6lCx+Rf643
5WGa1HJpsRgxMC6x/fn0HPGYy7EfoPGVDzihJg6rr7CWJkWusBNZKXaOIPS/lKLU
f1ao74ipVF0qh6M+OWzVWS+yGs5ooPMimyQ4JAxqMorRVrpUUphCwvBNGcYER+EI
XbX384/9PDD65v0jyoxFgOdxGHDm8/DyeGtrlmfl9IkZdvo1AutY3NOf1SdDu9Zc
o2VUKqZwLlrhmTgwo6PV6gr1QKRE/g9DfobwDlM+/yunr9nD+HJKek7B6UJRpgGD
KyoVSoxpTr3vnhqNLVyh5vhCRkgbyQOKjfkKQacOc1ipip0jZol9Dmo72jT5v2Xp
1lOP+ejygLnLf4HTKEfOR+6gg1VgecbRh9zBWjxiC9gXxbJUGS5vAnZ22ZWjxsqT
zuHK/VcrzJMFGu3c6ewlMjla/5mB1iDzXNrgTqVNrC6PCNn5Nra6D7DGelWvb+dp
LyXCxrOvBiMsEslan1kTZNztn4R9u5n9HWDzF0Db9gtkyo48ncQclfUfgq/eAqPK
REaVrOSBdue20IDwA4OuMPkKZWp4/pDpNJRJMTl+4tnP/zjn1rZWh8+aDsoyDHlW
/g5EFrxz4lD5kbn1ZLdFN2Dag9mC376fvEbUpTPJdU/eDDM6gKZxg2kPN402tHk6
klhbRyqX9LjW/6JTv1sCpOrPWSxd0pBvlYRBomR5jNf59b0Ie2GjnGK/MKAUewIS
59pjOnMqbxRRd1VWDwUczE/PtLfdb+WOa4K5Z6cmjt25oDQe8NsnyZ8/+q86ou4r
f+E5ZhZmxs5BqP0AHHhln7GLoZIL2lUIb4offgOxyHoez/4CO8T4+vbYD+gNzfRo
NNOIlUjN5uBn6t24j4M/2vcmjByvLiElkK9dtuZMq0q3u8WyUO6tNL/iH3l2zSJh
VpC4omIAMYJarskLJuEQgc4aZBnVnRaFoUnrj6aKtWHLndywnE2ACmYpQvs2im9d
BmXPVyVTGsAKaVX+DWbLna6spiyeFH0tzKkn4D+nL71ExD91+c2OqDAj9lNreayq
BTZQUgG5Ns1Cu0kY/R+fcRE3wV133sKu9RifuLNWwlSxQEQIhG7x8Z+vAT87t1ym
UjeNc5Ng6BzdzbpQAiB750ew4Vt9gSny8V1UXaYuWKgYQZ9vV48xoRSW4RYVqjNC
qc8wv42Efl5JEhTBQJ09sOkKYcUogMleYAuLp0upxLO0ZDxpcBKwOxKRFqfoVgCg
oX+e2ve9dnMuDe1X3UTImtFVsoHdv9xdJFJUCLEXNZ6VzBH8OoT4GfUB6RHKJ6fU
mUCCCPNKSeQMRAzNG21Fo0EAStwXMvzfTknZqYc1L8XcQeLo2dpgWUKIZj8g4fsH
nkKzjiQzr45lts3mX8Nh6UKUgteFlr9d5F3naMtHQg62OkHXxlNgc7Aj49kTfcul
GQT+wxLUfZkqMx0IzaIwrG79gZPeszN1P+ZqYcsnq7fZuuEF7dl4xDl2v9WCQnr8
WFEskOn6W4SsPENmn1PoYKwrCSy+yTVG4LXF4+gvo1iCUX5QaP4icKaRX2L6FJEo
wa6QA1hkIt3QqiPeBaTmNfw5l0lPY0HHTEM7KLPa0Ur8r8QPhNIR8b2rsWqn8epc
xHfQ35cNwER/bqBzbIWfiQQVFiioa71xuX9UgkA8bw3JTwXA5RDlUAxUVNdBL2yf
d0qY4cLlONSuUD50ClRBbMbICRirZwUKMqkNcWEXizOs83Evpmfx8v22cyytZfXq
kUaSBQIaiRhiQlmkziY+PzWb307246uru/cPgxbS4c0Z3LyXKYC7ldH2GW9lzaJw
GsNC315MJGCq1uRUOPOgxYQMHOeafFaCD9igt19sTOA1BHEguAruuoQoeV+QV4oN
oRsMo7+EiGs+U3x/UwK/toMKComLDh3E6jVabH0DOJVQQtsoDndYoa3ku5zpD9+G
Dte+h3rXRn/JrraRf1IP4MGNgRX5hxB1/QFo/4rwDZ363ggQkkX8zOUVcIv2ZuOC
aXBgMVKZB4mB6ivqFoOUQquOcgXbwf2EdNIfHucoj8lQOTgpBdnDVHHjiV1llbik
3IPxGwQvXu/FlEyX++qTI3aFM+6fqum7I0ewOhONODnNoSwQWIEnQXOxzLZmSo6T
JzJiM2tX+75Ch0Yd4lQE4XS7kcEw4JihWOCTue2SfsoI8mA0rHYjlMVjErG45hWZ
prVM4D5CO4931yOjyUEsPteb9mOUQg2e+Z50g/lY+BpDKgB7MKXFIjc8IcbI1RqM
6cR0GYRwoWkBnF8FMoptPCSFUWhYddb/J7907PzMeVeYRfmq43EtSi7Y/B1fhp8M
aKqkXJl4ETtuienTOn10blzbRSFI1FhSEx+kqE1opdcxuRym9kWBaNWSS7my9DsR
XFdkZY3/oxGBAhNOMt7EDBt0paOeRtUOlyrhbN3NaZ4RLlvV//dbElUvmimHi+zw
GSBBfgB1xw/DaAE6XdUAz4XQcc+nuAsZH+fiGhxHRnzUi7o2UzFlkDOErbxAzUvn
eBH8mW9t6IVe1DHC7+fztQaNtaFRm000cdmnF4yXFOE66V5nJ1ZT8Wfgg5aUDvO1
LfmEEiPENXI8zPzRtWnGU7fQXueiHyly6T97k3YJRjFiXpsBjrBZDShDDvm19Ir7
pCRTgz2HMITSENymz5mmZ1saHk+XLNAGfYNjVXSExkUqXnFddCD488caceINrwtd
it2g5d81M2fOsCquksOKIXpfqLIfssTMU+KD73eSXNTB7S4h6M8axICq8b1WT3+8
Of253rL/Godsv36TLrSozW7TpdvC5Hgjuzhos4xfMz4wYdezvo6U7MOLQIsdemi7
5y0gnQ7Xsr48XO/6bGy46RU2JKrpedxaypMYo4GIQE29hNv6MzkpEnUeidpyrt0u
DHWzbbQJ2Uah5pGAzbClPuAlDgNrPdv9xv2+O4lBZFuDwZm7LEjP+fb58p599cjq
KHMH9VVwmEBJiWlVqo2KFQJh2OP7nlpDX5BrMokb3EcTdGNicnyTm7DkHHJH7Wqr
q3xRo2zN7PMLybn2mrfU1mFc4y+qPVlwcZhW+RDACddJqfXnOK4u+0NUEsD0zK23
WuU9jTPIObjFhbgZ0JVkzhjn9QjSeCai7eo1YIAXHySu8tTrFO3y0+YLGarjK3ms
hvGln2/tA78YeoWOCehtwbvsOOIv7Cl3OFaZmrwGXUevke2qM/OZCSysSovQGzcr
nIDzkJm8ksPZ3x0EBkwxrN4JI3SM2ijRid5lUdMTs8gMn+ox9dbVZhjBbS2swvBG
3sJjiIh98Ty9qMlDzzRsvKxK0qG9zeU9sYHz2y/nyalZxwZWwWvwMQPLV4VYo/Io
hXMj2Bvs5qBfZpVhRocWL3OMfBfP05xFB3RXPtPNuE8nJ/MBsYKyiLcq8173Fg1B
UZLJM2DNI+R9TMKOVXpRSs+CUKRDRFCb70UqW6hL9GqbZplU0pvRD+rirFlkIbl1
9I5bTZ9RInUprnciwPYOYqXUX/rEZqTjyLUftiytZvxUisepmlC3QRUCqRcW0OsR
7wkiQJPuRpq8EWpFihYdxofTeypiyXrYCCwAcbPIQUNCgj1+V45pV5Fp26Zr0iAW
8qrr1qv78sXBTnazbtGHhRJkXqx73mRtzh5deQC0JsbybDG94mPk7O9MqDaLKBhm
SqP0MaVh1yAu2FYOCStI2ptfrllqYP+cN5q0wHMN7JA75eno2JDkLYKVXNIKNb27
Mcsq9bkfoEVdzQl0nrzaNCz0TJCNX4ObOc8uiQ1Go/UdYho1ABcBr5rEfjC9BMRO
9NrdoN8X1ldausR8hdZ66kb+LMguaHBTBab0JVi7GZL7HKi5EBTo+kR0h1YGfdwo
nPWsSIdb2C44qsQOyYD5q+dVBSrBOBUm4CtTQvr+xIwNJejKyscrq3rX1UX1nq26
S+jd1LxnIoJ0O0DLzf2ju60u0dAonoITdf5dmoub+/+VsufPPoLoXkTPT4Cyebrn
3Sf6mpWzrftncTlCcG5QCMWaLAJycRyS7/pwJNTMlwxPk/rdIzCIImgcWApoDsoV
qMp+cyhU24c+VZr2MUIhfAOUyfWxfkYGkTfpnm8eArksSQwQ/CtoYsjrem+sk2Y8
sNud24f1NP9D013eqga5h/SBu/dDpjDY01vE0QMJ1NAxGOls/mJ4q5ANIJeCqDsS
o7uCHTfPykmri9ZV6+4qVh/2qwRGAtoXw4qicnFLgdppMZ0uk7+YkLE1XolQnKgh
QbEPq9VDYKRIil+ukbeSklDrWN7t/XsPoRaE+nfpnSQH/m1h/O5c1QTHbdGa5kdP
opLyaNs+frEhx7+y6L0TtvUNEG8zlfeveuhVJawf0Qhp7BO6EWZWp2fWxm3IBqch
X35LYdoYH+kjMyh4dWWso2nnOZssZw/39MLl8nsEdHBsafOFCBKjwkPuvUbpjfJQ
/T8Ogismnf3IG1FZlpmTMtywgxzWqto1goWZtPJG5rh4jAS5PIWOckfhUvifUvor
q5srhTVMISJOOwQVgmRt9lAqBC9ag265iF7DEej/qnFQMSM/Fu/gXgYuj2p0kZ8y
a97JQ7XRp9kCNW6T41Gde01UG1dHQmxl869XBj2H28usvjVeZLomsV4qfOGtv9qM
u+/lmCXmOd6DVZlGqe5alNWigOpSyAWJXknOOqiHT1GnJKOOlOVvSuxNNVWogyKz
oava1s5JNUaFRjO9Rmt7iAksrX5kdEV3FHWkL7qJM+8/ZCLeaYIRlS+i7IcJsHDs
3tSa3nfOkr7+uCaikIbJOInQk/mbxq0cXufkEXmLanGpE+3Qtso7tIFhx+/4Sz7m
icY/xTavrAXsYmpOe3kwn1siUfMKKnR+gahZbaGsRFzXnYO12CSY77Ot3edD+hRq
ljUNoaYljxQ9RKyzaQoAQ3L000PX3xucNHdceTTUdJOu3N/3YY1+C5N6ewTiAsLu
gclMKoqZTgxWTyIR9KMkQi4+tSRTTADWcvp9zfT0N/FgwrIWDPzPxjMfYGDH/eqw
0Z4TU2qcsEMosXaFv2eSNxA+2bZDosSTrXONb11oOm+XO/UAzsOZxy0PrOlw4dH8
we9SYiZDaadmcgglBEBE+Px8VnKN/jtbd0cKpu0Y9b5bhom9H51i958hzX0bEeL7
fzJRlOnk0DnI3tk4Sct2juT8UPDwiH/8nkEfCthyG17GCZ0k1p0kJ3De3oSVjwJo
+f8hgtG3jDjno0sO04HV2hftkj366S5U+j/T0aYJergrkpTPjxL3B5vkiYatzUdG
l1iYgxM6dNHMkM1P60nu7fr3wKv6f3J/MhPfGIWWqY1rQjnzfTApsq8mCsmL5Kzu
tw+k+Iu+kmuAD8YTTsL9u9pAL87KjL3gglLcJak/DBrh9DP2Y8hzkkAMEBvQiYbX
mwu67qZoitOVDn8v3J+eyJzO3Fe90zO+KWA+1AznTkpvlT74FNSMqE1A8hYpsua6
ZoYJ0bbqV39XLPgaAiKoWa/qW+uEEBGm2JlPqXomgjB/FLr4l74ASIkxSKp8wwqz
oP0/4wGj8nvHnHyi5+6eaTfQG4pCOMSx2ybS5W7nd26cPrmbhrz9SKSP7uwH6uNG
oRmtZ1k26GiUQTym14+x9zk1MaHJkQ6QvLjLDpgxxvXdRSJWrOzW2cCDxV5DFFuo
Y+MxHQRKwxR3yK5MhCePwjtU/1N6mdMXrIY8Av/I4kB1lkcSng14zPWEJj81hWiS
VOHWrQ/SLJEENvuTqYggZ7j4I0HqmG1rIkGA5YxW3ge1XOSQ5kPXDtMzlMRdm+qI
7MqV5ix7RyCZDurgxT+Peq8XdCDKw6OsxUkMiwY7p1+bd1bzTqC15uksylpcp+Lb
1Eo/2TC+M1NVxFxs0OhV1ksMl5F5DqJaxd3kWeYG3HQM/tDgG8sKlAUTsTD4dPup
RPloepvLEXaei32PkTmmm0vS4qub8ux9EzG2yIsIJ/8SYCYHcSr4UlY8D1M6dapz
ARIbMork8pnpzuRR3KsZ536S8AKZBexXQQydIIxxTyu3URAtsiVLpr2tpzZm5bWb
D5QNgq/U3bVm27ch+xbV0pGMJFSsehEgfrtJeEIKeKmZdIleXqYzzp0Br3/i0Y1j
HxjwyGM4z+NYaD+O1vaUO47i5FH7Zfp6FkbGPwJ7P46oj6jOhfZ5zLVJzmRxwX3Y
dpihakmgJfcZqBs05M4ft8G8o2b956amaFOARVpB4/5zSHGaNOcEVeZuKcbee/+O
bcFJT+ANnv1uwPgjIrRepzNGW2SE5sE57L1uR2OUFhz9yJhPE+TcUAjVi50YzXOf
sPjRSoEYUFkHyaLY8bBY6hKKbqPW6y3k7ey5sNaVzqFwe9snaicQTh7gTkmxEJEm
lAHzQv8JlIhkUr4CBU1isuR07/r1HRQa+kw/91wYPaQXivbcuYonFu770IR4CMaH
wYOHUYFSGiEvDVuaOOwpDlSzqXfJIrXaypX0Qyjn1VeIbxo5sEhLV1t0pyV9mKOd
q9ygP7x78z3UblziFLug4xQ8w87Q51e1k4a+pm2rbgWYd/eZSy+j6L2f8LyXxY6X
PqVqSLyFa2sjHibUeah4EqW27zzXnd4PhHwqG9PyErRF5nRQWOYXaIvsDSS725Ou
rQ9gq9NdHR9OrL5tsWCayLqQM/ivhvf9YaRhllrGOf+gMxJ9FX7blTWgtIHkHmxk
kXTLFFhRuCM9wTmL60zA/3BpiLU+yPWywAu33H2ZfgZ5OFLbGryWbUxHBFSvDkrv
ZsFEcR6AOpaN4npNXOixZtzqAccgyzckBgkvWhi0OX+IpX/bZW0QOh6s21OUHx+W
xydJtuwsRnIikGn9RUxKmlAbBiUc3u2NoRdoWlQAtzD14CPlzxChz4gnJLD/poZ5
UDdJyw0WMr2aAToiDhc0CpUcrSzAB4U/hPavH9Xw5bPIPUu02Lnj8tz7Z4XeSddR
2BFzVU2rhQq3LsXl8LL8TdF1FHgI6tL4H1xIid4GAHFt6+yeop4wneXnRF/P19xo
k/1bji8kmFPCkWeMBmC7sd87pG7eFUUfAmFW050HL709QhIi5+zs9PKGEOIamjIB
/UgDBrpbozksbwpj2ixRpXK/UJnHXFuJPw++HacPJ6K5BEyxtFR/qlsMcgbQLDXB
3hWZlVlipbHMzzLphIaZn913Ina9Au/09gcvGtYnDUYmkgfNiBd9BoDSulVwHWew
qws34J13QqDuMIEHIQjvNOXp6CCDn0fYFvMPxg7BkNifCbp2PRPgpaHDLlc9VsxV
5xEst/wFK4X+VHWNzP9aGL3OZ4zIZm6gDjleX/2ZMgg3bUafAfe4mgrLR02Z7ktV
hwA8WEoRnRfn3VIhmUWevxGkeKosy8XgI5bo38o4E0MZMjAO6OhIzNE116/cMsYb
PO4KfQakW0Zj/+DpWNSKVfw+m/PtjMu7vjqBCRBINCC9dKz/wUvRyvOBPVk5XIQS
Iq2vYeOy8eLxe0Q2EMcKu+2L5GYpOgKFPK/OWCYpmv4sSMJB5iZPj3Ug5rnWmvV7
cPQR95E/PGkiTSQbNzGQn7K0jxXX2kVOMC0V1zX3941nHvIdX1e48Gz2oKA27sW8
KhDMjMZB8/euVLHvXk7IL8lkC1uaKhOMdi0xjNkiG8TjMycBUglZbbsEEg6xy5Lq
esEBzw5BjarJAQ4DVYobN68qiGiwcCmy9n1yljvVGyS+X+bd5kWLCjLUI19BM4oj
DtgjDPZIDOUDMXHTLYJIohyzE9+eulpW8jiNGhpnhoL93Xl0UAemNPmAI5fpWCui
ceiI6Ta8MKl9dBCWL4Pz4ZwSdJINjPZWbkF95z3ilKrnmkukzd5iqB5OXsJRbL7k
CsYSMmn2oM1HPFrNHbV1wUC3SN0gzsXzLbV9lWzi0sFOrHzq54rHyTzqF5ax98JZ
WK0A6Jt6KCXGxa7WiYURzzz0M1DXBrm9fgpZghBs0DmEl4l7G+D9INuokRrP5PPg
i7TdQaxHL38nF/FTKUTWJnZGvxBUu5fGjvrT27Y6b1QLvuNPXvTFYxFibuF/Zg2a
z13ae8ZC8hqxeGuA+wgXjNFpgwGdpjriFMUim7CsdjGgBmCcefnaMF4UkO/EcuYy
UkllItv+VpWBYdlR3ztU21uycsnv0VJXMRvdMrzEiqaHN2oEJljNzLepcA4yEKXM
7ayssbAhAQ5K2/G/d/uEzmL7tVRWheVf8sMc6XWjKYb/fyXUZe9B2YBkeKWW25nf
ino6SELsSkoWEJCLV0uHlKhCzK06UjEUBSBnvkKxJGzTH0+cQil7mJ0ecNRKDD9S
L4ex5qtXWcJXouVPxA5fKRavgCxIVjHe9pKdz5INS2UIghGNs5MCSaXLsEFGBw5O
ylrKqjzMTlgAQb4RGYEsVKZ4OWiAe58jksuccBX4D7PnT5Fu1DGY+bmtxqyhs6+S
GqR2LgU/1uqHYEufgZY1IjgY5G0qgDyDlq/AXx0fxznl/rdG6Ndhqg+P0AsovrIi
pvwFXzOMdNFveLI4ey43bsWkYOMEgDcilhV3uhBr+HyfcJ4mWl7xQEcZOd27ywrT
vPi72NVmSmLfkpdikZT3Z2DuOibLoXM9DmCKP71+SHeN+sBghxpde3VcnixoFstO
LLNbAwAzFHL/zmAomxnfahFVJeNHaPRA3c1LGc1W/pJrVMwUlAwNEO6mV0S/xj8d
IYX9i9rcuwhYqqlK+g4vbciwMpB97rG6jbPpZvAz9XUp5UIF9mmpYqKefQuz6ntf
sFRKrf2EYyJ641x/9nZz85LzpE8Z6EY06eXq0Ml6vLjgucYiYGgYxa2tuUuI3InF
CdpEXDXqfhndotUSTYtmU7NGQgr7xG9ojV/wjPYeBMeZwrJ1loFPq9EGmZCapm2R
8o/PTHbeJf4mqJqr+sDy3Y9GoyOwdTApPKTtbzfwD+3WrhjJh1gAwzP9KI7bF+Zt
WU4Famdbq6ReNPLsobip8bOIMhSgyEfZZ2CT7eumQ4N1EjzyNVqDGH/mv7M7QSRr
NF4OivZCz6ryfpNfrjQtul1JMCKfz/WqS4iI3JzDPuP6mXR9+HsTLJlYq+O6g2IA
3J4SyGVDYRExTE4+eThGC4/G9B2+1HejJv3wInm+9cUm93Ev5xGa42rgj/a90HQI
CjBWmHt3IfWvbI+uCd9qTCJzRusPdzdpNr46oFPV/POV3FYQcZ5rL51pOMhXi4iE
Umix0c1G37INJjQKdsYyE6XmQbTG0n3HCtgeCXWGrR/16vCjkeL5Wb/z3T6DzX+0
NJ7J9C1AviNNONM0oABkbwUypZqvMJ9c1H6DXw1QgSruY9CDBOt3ujyv0ARFkeRw
bNeK3l+2KuSi9Q132nilKeuk/4n7vlBhBaYsiywu9u4r+21I8T6lsqHjAYaaNzRS
feJauvvUjS53G1QTE9HccrmO8JnXyZj/80A2Z0PYl8/Q8A1ldMz48mjfl+KdUss0
zTMaVbM5wHjZWL52HXliKaOtTA2e8dA5CPsGhij8BeqJF4FDXV6iEWh1cFjBm4Lu
coecpbVIerd7xFdWs8qj/lcHSlVsvwatK0Cwg7OY9PPv2vvOiVCFRXENLxgvxVpb
q+ly9mcn7lu7pjO3Fw5JS6fVL4jaTzUb0xMzodZU8W1wgliLw9YaTzuUP92Y+1Zw
Pc0jHcUaAzTpJKzlA5VBuV3KfTgWMN4IbCU8qVox08uA47vh1Mi+TBpVFQ9PP/yu
RTXOZx1aAM9vuhTmNHgBwpoX+BghA620+oZ2dIGvIAesyG/esV4pGlHEDDmfOc5Q
uBHqrDM/SuL267SGnnP6BQ/0oeeRjrRdif7Dvpl7CmV1MgnDJYPc6jr1HsOEPE7O
TA8EB3hTbe9fgOgZJ1qN8pFQowLyiXBuV+OYKacy2ccWnzHp+n36wDkHES4KV8UA
MaABl/H0V3+qzRAYbRgj1+xLXOZ1+qcB84QDt4o7ptRjgjP8Zo/EH+WhvDhkgPfY
Gqqa+HSBP7PkbHjMM4RfBOjh1wgzIfakHJu8oZ38IQVeLuoT/WGYUagTE21/eJRl
/zijZFIXOIUE3UF8hOkZd+iRRzXi1Pbpt1D86gM4ihLHauDUnPK31/vxzMkhI3BN
k1qMX1/wq97FpJSSXFrAc2PLJ+pQgVvROXdgGOtdibAge7NOdOOa+uvlcxWSewY1
nFhhW7H6tag547/nJ0yWVoFaWQyInh1suwgoKaq+2/kQzmNJMGIonVZ66k4SHan3
/14aKOgA7ZFXKfTS3YVEeMzAu1a+6hsaJm7oBaLlnBl/HnBUbs+tPvF4txPINCKE
Su+lG9NCRhiqnYpuhOQ6Umo4P44LsRtyXkkb8XIzgNQNJ9Wdqa4X6BYB5wVf1lad
crFRU8SoXBuXfUXZUYzYfcqpV709F0XHAkyf03ezkQnWPcn1BPOyPWmbbn5TjGU5
uF1ch9ZzOI3p9STCQBfNY9wRorTj5Z3bwVOdjTeP7bUifEG0q2wkzVbaHjninMti
H1j1xc6UMOpk07ILVJ+3o1zAa2oZdN2c3+8VZoBtIccJ47w9jlPbpqY8V31AatZn
ckf5cjPFiW/SnQzCNRClyVw1M7RwR6vhfIDoJDOMyCiI0krMgD3nNVvyeKk67PXY
E84C/JXEoKoJUnG+tc6mFQ7kWwS6hjyKtI3qfTatM8HggTssKIUK/uhMBYh3HcjI
ONBk5PgCz/y9+A3BjgfCoAhwChGl+/3qTkU2gui86KI5Bwb8vM5rOM/gwiPlHyvx
jIdKuuRM78V8Zd7HMMZBtKcn7hQuKKs+XtPe23+GOjDw6USe25fDzYMbfBswRigp
vt8Z63Gms6d/xYMOamVG1PGqPEtaHXk20yywGFl1Ry3AqcuABRNTJM6GRcSwxOGu
hql3JHFMnJvdXU5Kh0WpvJRRMOmMCDWx8VJRtO5oCLjRFvmzUMmP4UgbVuyavfgS
q4I9Z5jGLowaNROKM42O1lDaV0srjJoKs2ru9/1LBZlTkSj4bZ/4b8y8hiO3cImn
sEzjnBQfC2Tbq/gOzu5u5J1A1fPnMmwWd9+mxOuuqhCdFV0uVX4oebZNETNNr1nn
jf6wpbYYmrOHaARxfrzJU9f69FWGTQPfG/OgNEcTrWbt2VBAbI2b2yc44eidw+fC
J+J/IG+C6N1JZrVAzMqph7JA4Xppk1DlXLCR+6KSLtWkcaSkbufSOGXPR1U7Nw7Z
gKYQsmAsz/7K+BlblmXX+grrxYkn1cxtgJQ8WI3upGJcyufOFioM6y6IZ5vVxKCh
Zw6TIXOQxM356N7ohgj2QuR/daesdoYnDIkgms5l1Q0SRGSg5xY6tOpDVllJPdx4
P8ftg3SvmkSD6ZJT7Jx2nrUSp1r8grxD9Srz7ZoZBk/vdtHmoqrCmjtyM+zsyFbu
IDsZahs6wUpLyNT4WYchpeoLQ4c1NS5vtXUUSWu6n7TElnPAatQ1OsPRumV3RfOo
9y/jo/wpRBB4uOzLHdKCzTvT4RjM2OOqP7vyQdM4Sopg3jj9iUVXE0PUMqVznKL5
dMN4/lUuscz4mimyESF6X8QMbyXFv5GxoajNYUBAZYjo8OvALMhGYrvFjUddM5bk
OKIr96E9u6hUxmXK9/WoceeSbBHR75aUYaFyRi4vRdHlnw+Ttlq2xsUcBuJi4o6r
6oL5XqliKHwJdyq9+n9cHyl2N9nW4chK7znSxNtfuEtWLPQpDt4tyA4qs7h3mVb2
1vtK4Yw8h/enLd/586qmia1h3IHq8tx14mKZCDKjyyZUSDHOIsZYvVq5H/W5yhGZ
qgWZI+OAPzucn3GDaP/Yek9lfe/0N0AkTGrnYyu9H54A2t2k7RWL1/yEQ2iYMw62
7KJkFq28EPMuyK+8xMJV5JH8Ziwing6V8KQq/Iy8mfKPoX6VUgywx1KkMdvJbl+l
PMLBUql7t5snlOSx2aSaL4I6U9wPPxbnmBqlrZDmewrk8eM2whT7W2JUZfk2JRj6
y86PrOccMljA0sOQZ17l6f42ZT6KaFvmfnE9qVR3ARGORAtRlqUO24q44yhZ7oK7
OFHDSxR0lHP3cBDFpe4AveO/AFM+R0U1g5H+AGcvZ381qCY6BI+nTYe2qF7kZ4hS
v+xUYnvWW7LZdGiZc+GtWwbTytYI9k7CbHsqI+Zu0/23J8ru4j7fGVmAnhub7LWO
KtDtbJABiLliN6Gey3huFftto7rwtSJQSUZ34h37UE7wGDbKhCJKRmzmuiAgz9cu
e7CAziTQXj91Zoe1dwou1g1YwA0p7oZ5UKQd0eB1M7kbRU3vN6Kv+QaHhAGK3cIh
X7lWitn3CE1yf3/5GuS1ay6SVM+xtPu73Y7mN7scWSttkpk0HemAeoiK2ZjdV5/k
IHchbpszjgGwZGxeUqW6c9rGleCzrBud3lZuiJemAa02MVGIVV+Fr78bHC3d3CsN
VQ9CSyhHcPR7i10pu8O77yszZfC5nCUhsn430pJJIvpqBpmMfm/ZSMBO7b+51g9c
+NSTtZkSX6/GHTR9RS+TSJbKO1iBMvitdYJbeXVz3WcspjGV7aWMzujNQTwXVwkD
o3jHMMR0LRRZmic0DDsP3rCmjuaMvS/x0Ea1gxUGKsN52/7QC/vQwt6m89j0zw6s
G3Mn7hpN0ghSPqK/rrJuybacwlLIX9gZMeaWcYKZOfkMjR1/I/lcctOrYK6n7wif
1S82RDyuoOTZ03kMEaH7Y5/Y5fWSyZUZaD5FDltpNa0CljDVx8sfp1fgWDd5YviH
5ATcNnJ7ou7eC12WQ+c1HEJ7aFfpZ2ZDrBbmnW2+SScYPg+Yjm256bN2uDGW7eOW
t7USi+cLzGtoQ72N4lK2AyCx0nOTsTR8tMOmMeKSjsgNWFW6uh7Hlj0ngtwJwzIG
XwbXGKQe3tSEfViJqH8sWG4xhlV1YghARbrm1nWjjtVQ2WclPGzHVTd1cTftUYjz
PxlQzS1sioRSgBWTjCmxz2w+8Jfy6HizR89Nx5jvMweKFAYVXbIPQk9DBA8mA4/O
OjAU5/5rqcU2/+Bkf6YA/ptmrn62e8WypD6Wk4/dnm71VUhMFfOhvP96CdY3a+le
l1+agYWdDFzIM+TrF/3L0X3GMAa6WT+eITJaQ0Sl+S4mghHLkXeV80FylVtRoBaM
uNl750h/y8k5YwqtAKtTvqaV/XEubHzPWopmPCso+OVSpfuKb2DUIMFUUfV+nD9S
J0+JMt0Ao9UJaNs1X8JhYj0kJhgQggBoi3h5P5IT5P1PjVKcNIs5ero4tMSiweiv
/OIdLXJshUVfzx6cB6bMa1WpKnn6A/K5NxHYnLjqL1f26DYUijTy5NsbJ3t+iQJU
OGSjU3/LDSV5syrNot8QhzBnV/jC0UJbgzLU7Ve5kmoJJYouWPEQLrb37fxZH4Kc
tzVEFdaecBjzK6WvT9YiP3yyPq1WPwLSTglMGdD7fv5L+6tgR/gUZkmdbYwW7bxV
6k6y5JwbHoI84YYivPxx/LYnudIEhyweBz080GHvwN4ELkakN5F3aDJVuZVvNY9B
ENtXXnl5eUXMxdol5Y2p4K6BywSgTIcb77XkeeMuMxRNrmrKEOMQNRRYRbE37aEa
GKolB5OZPUBpN8jRxA1hEll88UhHn2AGmuLo+8A6jWwty/YQbP90cj7TlyzXHWjq
bL7p4la6kvVReDi51VIGX7PioJUnVDqM00RbbuLcBl6b8PNnqCJDXYOM9XPOY4ZB
B/k230Xe5cfAHcpYM3GMSYlzhScBterJNN5W6STqRy56jIuyx5LN/EDrT1yoG2we
UIsJMoH7a5ecMGzbnZf4CJ6Mwgxn/Lh2C63jufaQqGpz+uPjnPcxANM9R50udDvb
UjCkn51LI4p9pC2EvBfJ3oPhDLH00j243xEGeofN9oaUjsyJHim1+4udaxcfCR16
RDrl/Np+KMdPznrEKUfNyp65EifPS+gTND+55Tbvd8YA6RFnzAWBpHFDkCb3gc6N
70yMLLy+5MUu3ladvmrhbgcbzE3yaiMfAtOelvA0deqL3saKzweam2cu2EWEJo8c
vRcITuDGmU2TNcW+RnAn0U5jmFoxvngRRqIFBbkGHY7q/S0sLFAOGLRv+pvmylri
AbFXIosV4Ndgcu0DHG1xtF84QSVX/Yjk6HMVwveyQ7SiPXYQNvIWoX+8ag6Sx4f6
RNN8633K+eljbSzx/zPcRv+ZHGDjkOjmSOC8Gf3/ys5a0w85f5Od/5r9NtmcraaB
Ie0e7/9mll20YsTMLvflsRks9BxFc8J1bpYJPq2oedpmbOZXc00UZIGL1mEDiB5E
UtmL6gpnQ6ofsYzNCgEUDI5E4hUGq/jWzqP5H85NF4FuTOYe8AP+tSkqvYqEFj9w
jHlRZTjIxQDkDW9aStm1eYKnaydODdeSw+wRf9Y/yei6XB46UKBM/ltoy8eRUjBX
U2bQ9tQcs0bL7JrZgBYAjTQk857+hDWtDVvG0Yurk8O0YFZevwsceOnekUctvNx2
wlZAGEThqHYHlvVLax3Zz3tc6GQpg2gvSMStHeguNShTXU8+6VcVzE/0hFHm/dbj
k5f4HT7UOQYRb4lI0x3+bGk9XD25HUvqkZ9udvigZd+rr1b97kSyZQEXLXTlVlNR
LHY+g/29/kJs9PnKXwu67+F5NZSPYxoMSSyLW8CLQoO693fZxYi8190aTmvl4qTq
aRgHxe9DfKwjcUvXzLZSOe57wrx2hUW5N6EQp6UnpOrf6nln9vCQ/UxcXyzQdPM8
M56ehEdNNrgT/rs5afHX8Wh4B8w1DlwEp3R5hPci7oZKUNVqSSW32EzwhsPxQbJO
nXAJ3KTvS0X7NuUTJ7OmDU3yH1XKu5nOV0LmziaZyz88RkGI2vpeKseeJZ4sS8fm
pwuqhxS6GFW6XhOd0xXuu4ql26lGO1Lj5djXcCiA56PVE0iUCwSra+OZl/gDPa6N
LrB81q2q8gTJTzRtUAw60RID6VJU3AYCK7WWyWPl7HYEKgmoxLnqCddQ1g8P7ahV
kFRtrUzjKdZ1SqeOxIEFsEYWoocr++tSO/C+A2b9ojo4zUOnP5b9XLw7ofTCMKG+
UYKoawjKUQRwzbi3mTa5SGifID1NRHIIGG8S5Fgk6eZ0W0kVqpVM5ecn34SzC5N3
Sp2+EgkTUolJjDA/To1vN4ctlgUc/VL3G+wJfSQMdsjkrOHjndhLpGCzA8pNJmP7
2LHxWVauSMr5F9HKmcuS5dreeQbUFkCvMSDTqHI5fpPKcDqZWVQBD0l/2Dqksc29
7vH03504wKnG+Fs864O+J9VhL/4W5BQE7hRJ1d3H9aQT5OSTOCPGPbDnnXjJIIXm
vBouADyBvT4oGw9v74wz21iEZ53PqBsIIuFAPQHxP9z/BDUsGdIpwWRSUCP27MfC
zklKHEplroAsIiVS7G0FOJ3FFQpBnK3gKpvCerDNhsR5dpBGMbzsH/1cxHZkXR4L
QIhVQOkyY+w82HdsgiUniC6fJZ/4LsSIrIKrGQASqRdkuQmDsPfr4dtt8HqmPlbJ
jD1UnCU1kjm2ekTy22WvH8wq0mfgAXjaXj5qpJjNgbdZM1O2UQRoadA3AX7kyXtf
F3RRTu9/ZJnFsA3pkgTwZX6tr2i7ZBnHmgyapUYUEW5wxj6pjvTpEpGdbZavHBTg
rtKmU3chS1DDQ1ZDwapYSGWuqQz5QHT9chOBStMdPOII+ehpXJ7mGk86h2yG3EE0
RuihB4KyO94dGGxHOZK4S1Cc3JXKOLaxsaWCp/bUandCUxqeVHCbpglLFo52BkEL
OyCEwx7K65PUTKAaI4Ra6kUKQeOvZiiM5orK7JKyfxAaDmbwCUaPJcEMS4tiojL7
DyOuXf7RRJt6nYP2nMenXJm8aYUpNOJ9+qqvWZxi2XGerbDMpBBHSzIJxAPTiiFx
WxYkGqINWjxMuminy3GyD4BATLwQrM66JUxpmYOwNAFmdAvrrKzKyoWxaw23Nwag
Cuj4Mvj5EtcbjIDwV8Z+UDhHDKRE/eU282wveT87GRLT9KvNzLxrd4tJykYmg4Nn
+g3ZWir3RLUas2PY8WRTw6qlSz3mwkKP80xFYs3UAsl2WqgUt+atCqW2KMGri+d8
LcgRN8rFXwgBwr69FZUFjqymH4ziO/mC7o7an4fskzSIo6FEKS+K1vCjbbwaTtE3
qTv/s8pZ614/nvanCaNsRrT0pTPxUAoxl1pjemXHteF+Yj95maCL13IFf1ImtNKB
moQqNgROmH/d8P27PALhubQpK5p832zwdoo8l0TQOH742/YfNT7CXnRRmSyBPt29
kzQ7lAatuKwR74wNFZ9l5cnERGgZgq4DqInkpZ4v9wYfpDceVvL+aMNlTspqmJuw
1BSddTq7yr3F3hgzEaC+nktSVy3FhwJ9DJLMFmks28+chjSgmDY239xCQ4yDlxwc
LmTogFX1LfkhV68eho+4v6RVs/Pt2ZQaXzyGg9eGPlPXsbc8SpdId6TDAtEuKr2O
W1KneXEUkQVDn5pCfaN3+OZJW9QclRrmXLHewbzOsPvI6WWybEhnVd22tx178hPj
CXFej1swabHyyVnCE57EjB/1QB7xohfaJbrv4A2wN/ew84rJGBuPfGK7M35Q7eYo
q+i9B0BctePGyir7HPL5VfaoYxrq52bcU5/6qjsd8GH7sswD6yWRtCn8rYlYIbjs
Lo7TbJnt/Fbr2PeOJbFg/PN9wOo4CufkPzdPRcj3oLEVZcE5B8arf0UudMQrSWKH
qVYupHlrSWtBAHbySm5lObU3NcNvuP6pVFw6922OMioUychTsvyM1nux+frAR/Mg
yp0yA0dFtbuK1wJCJe27xp9ULwakbpSaJpYMWjmfglFtraWCt8MAc+l57Pl2sQ7N
PKfhF4q9JwX1lD5koQQAALSZaqwmZv7UfP3suXNeCXPWnZXZKs4COAfPOJWVqApw
PLqLtngFZgQ7pRhuxnrO9ih7QZN0ACSYh9WZhP5awwoNA+MzZOr8lT3zW9+6Sfn9
YwNtd0kmO9DkyiJM+pTjQv+vT0vv5ZnA88XSTLFVmHGDfuOrr4XtwFs8JY0GCzxv
mSTXZ0gtbOH20yCY18rJOv+zoF6kY5CE7TwK94OJFz3y8Gd24Vgm67KBh96PwwT/
g9tf/QccDBuwWJH+e5pzsg4uAbCXfEc6hS1Qb25kZyZzuYmO1p+N7DvsS3EEeVkP
AbNZLjot8hqooV7QABCUOLcchltBRKbNtVeTpI+YBv1u4YCg4l4t6sqOqDZDeZjE
U1i9WOkZK+6rf8/eID+D9jfxA+GL99rGzYW5zLcMDWMWsJwPEV07Jrs/D7g7lvd9
GNEzD/P248xQ1yioub/KzpbM7aq7Ys2CZxU1yKPYuUVzh3fW/JZ6t5UjfEUmEnD2
s52TY/EpMdTBewPF8wzNbrN0JYnYN2eiJPhlx1JTOiiv0sJubqxDq/aScNtAdG0Z
RCeMfyq5T3uUELKuTnh2FKsyk7fj21daJxohlfe+McaQruEMoj6AhWzJO/Lyhqqv
Qk7UYe7DKbGubH2abhMCywiWURg49Xlex7phcuGOsJiIb6GDCsx/WNU5W31cDpIr
RV/7ORsPal7f4L1asrG8+RrhGmQ8BZSQdj5FKE34aUTlFfE8q1O82J3Y/LRaP+ue
RPHFTQVMOO42FaxeRHmr7aNXX6IMQAIzfW+fFvhGoOxdy7U3AAsn2MGMmnRJYtjy
i4xblVYYz7af0C6X8+JMSpfAAh8vE8zh+nYNQfu0PpKKQgyfrqIdJk6qs5iyoq1R
uxFNSmNbCNv2CXuPsHYw/NJ6qCo462hdaoye+7zdrxFzfd+IJ0q95QaETVr5IRN3
ZUwUOj0pcDtMq0Y53/Q4Ksl7tUcQxJD0tWohOu0izDulu5esQgR5ybt21rCT/C/r
6nubKlJlrAAjKz9m+i7UMbyq8vpXTLpDo9sJPTV8bwJpCPY+r5oTLxpFmhHZsUmy
tKn2pIoCAM8mgluV6Jal4bzhrmpBzvada0kfT3buf42gwqsOm9h9ENDb6kp3AYOb
qGEm9QlTlE5tJBKebq8q6Sb/L9NnsYUar097tdSoptVWLPvSatY3SeP7AjyLjV8g
jLKQUVqD+XRuRGhBM7OX4lTLeNVErw+79yf5CKqpSZt28Lch35BciUjXKROGpT/3
8GDPMJPgZEBqyl0BsxNe6xDQNV+ByncXSz/mUzD6SwiJElKAZ6wFtoRP2A5QbBGs
/H7gbvuflGzn7GiHggE23xFwy7Cw7GLQmO9zHTitI/1rZCiYVdlaDXsx3N+fw1dH
5bsBpiEX6p8QBwF/CmYUMc8l9z/axUJDOUVTh3imolpQ9C/Om87fjpMODKMRRB1F
42+rDT2REZIzn0F9TEtYkhbFoIkJRbGEAZpyDYlDbTlRYgGG0w5kFytcH23Jaq+I
CGoDj3FdGKG7ZiChHMgSIRh2hsDTPwGfexnAQEHS+HlwRr6xkH9f2JEMP/gLOGIw
hlrmR2X2Lg+bA2X+dHPrx+AF2CZeG8bvJqfJqeCpGOR/5oY6jbiiTf8ssaHQ29hA
WjA2fneRJSRZ14FlaDrW7KieXGFzL8nZbw8HzU50a7g7119pZpvyqSYWd+4NkV3E
CZOQNkgh9pQSR8sbuSfKOyCBGDtJuhRgvHIzHM38nzIX+nSewzn8BfRXdjf9Vbl0
lvMFI9VKCFvzUAykSOjK3WAWYrdLFGHFG7iUP4XVk3SqA4XminPTXJ1YXV3VvxEs
MzzxKHTZ+vZg1KVGOROzjki8tGt2qRJTDoF1dQmokXhECDe5GBpuBUOrDPPyFoc/
uN0I0X740e8C+N2EIjRwBa5+kuyT2hlMVoK3+kCwBJIKChA7re9RRxm6l1doM+Aj
`protect END_PROTECTED