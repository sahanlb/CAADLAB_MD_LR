-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PH3PqlAlNrPMXKiZy0vsgSGNVMz8hEq+bzacWzG2suDwJQTV0J59DT+jp16eqcPPQjq6aLjiOPOh
ncxRT74YJO6tCLaZhOJhgh5gvJ57PaQZSGEA4V2qKBbMoINX4QQVQ+//2R+BnbPk8Mt1dIxVTxuc
O6I3AQIT11LmazWUEucPOK8dIkW5kESyahrc3oM0tPryybZNB0bY2T1HLr2EPMcm4mU4u31ogXcp
sPLb634MOZnIZQgJXz7qwCkxU23Aq0EmUuWJTR5Qig2VTIMxVywBDaQ6jnMJE78YoRNgnaN1HCIj
85ySWakDXNjtkX4a77nPJOEQPPctLXxN3BkMSQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9280)
`protect data_block
dT/F51VFyLJeZ/mqogzCB7HQ0qQXAhaKm/Xsyn84hzRQ9LynDdOItpm/XUVxGD7DVIwtbYWOmE+W
rb9Ofayc7+R0XRVQxAOENszglwA+/8glv8L+iDvPn1zyMZyCbt2jG0DHrKg9ctgEp1A/gVh4II1o
jgpbzSl5vbmulkQ+qF5BKcubida37bSjhXNpFyjWyJB5KqtFuhcvR4x273cX8q8qiu8uNeYk6X0y
xeajDpyPRHTKGZmBaZO5Zan8s5aHKfUkS0evhitrkcHCsGc0zxK3suVxcXYYocpGkWgiAIwWgMxn
z9tJcCTzc3QNZdC9ZsHt7j8DCiTPmi61nNRvAmxvoqvlVy95GC+FnqSiQT1fPOijWQRP5BxJ4VW9
+WXa9RL32/TW91XrisIIplAbNakhUer0f5GrdD17pdDrBzvBQW47ci6JPuGdex0y9cFOZuiwSNcO
6c7KbqpvCISLYm+ASRoLybTphg0/XPT1qQG9YqYKNJgZNKK0I8prT8902bySK5TUywN8UUNoiH5v
U5INTJ0d6P3z5inmGdPASlmQ8YZIzL7unkMI3fmK2hl4948EG/OjLf0jZvtfmg6SNEG/C/HlQIVm
bNgZ70VIW2PnSuBmnsxGI7+Wbg8LYG2rbixqreURA0QD2fvmtCQL5lXkFfp0KD3yW9b1jn5R3w2s
pmN2x6G4eTQD0F26HdkGQyDjKJqSk5CGXBTV2qaNEiKHmz65UyRTesKNC5J4rlRt2jiNtUfBgAlK
v+TQRfweOpWJLwSWMeViKAWvSP9++kEgyhS9TPw0j5RjemCM/t7q0gXhU0cB74NfnCmX11BxbM4r
q6LQe4ngV1GWr/bZKr0k1mcM7B5pEc9/N6txUlbBWmj80bmfAR5GoXD4dl9wlfPjNuHYcqCmQkyx
vW7HVu5IS86IxpNRx/wrgN/GWZENjUK9qb4Z69C4nQjqsrz1txgpYz2b5UZYRJAKHT2pehAqENyH
bQvxz8O7sb8l0bPVN/ZXR7pCnR4EpLx8NmS69dvfKZPXOybUJbsqyCKAELrn0uHuc+uU8pENUWxI
1W5FWkpmFXswqcyQOfo6aD3eY2o20KvDrS+nN8R04gXiCiJ20iKP2+LXFnvJsU5IlP5VCrXRQx8L
/zdvCHsqyXEYwk0hG8payGAg7BN7nXgMf24Nwp0llr/cj4UuDcu3hZ5QJLBy+gQfoT9PrpdQL+Wv
casIi6c7dzOEJVo0REicRAM01cBF1QGD6EoK1wSCdIxLJX+eQguE8zMGyYMOv/0imsw8qIamJD+r
1Ro3CbbTqZtqKtV8vOCFcr/87LTGDKdaFgs5kRfMlltXpiJXnIEuSmK980BuoBR+9u/FPLrWjINi
LaUnSDw/naZyYTDp3t16slhsNitimZul3V06e67llXH8xx4TcT6VJzuvYUxzTNLlds5ysa5w7y+k
I4/SACccuWnuaTjQa4zQ5qVXgRK+FGCjiAN1uWOO7j+ODsSUx0rTjkt13fx/OVTsnEOJp2R3qWxa
ognCvMU1gMoS5o4dvgQNBPeT01n0Vki1wnOuHngLsgk+mKr8u3k0Rp2zYsKW2tthItG6M1IqVydH
gj6EE9A+Q6+cG0Z0Xt6uxGqRyYHNo6jwvkfmO9O8vW789GhjlAcOfebHS5jCrgCil4GwVsWesmkO
U8DqAxM9xo4/EYMxmE3Ry/u7l4fsXh+IksT01UbkRO05ZdzMTK/0ivpo72i5/AZanReghKzwnTQ1
Wp+WmhXwigX9qUzU/xmV9PPDWSCnawZSIhib2viPB8rlARf+8ESr7LjbdvZ+GXZiaTQIBoW8f5wq
t1GBzwcRUpzrt/45acce0gEGWZ5B4YvEmkGXO1d201A6yTapAlJ7TCOkkAPXVG5XwZ1Sc5YWesdv
pkrJQ9JqomHrAuhLBxckkN7JlzdBN97OBEb6J0gA1m3B9lk1ZNt9EZMpNDQKL21I3EraY8is4tNr
IBXae5lRfm0DvMAkB69vfHkZLtCdykMJBaNXdmMAD4YYrazLfls2Qgi8uhmYTq1P4dv5VFv9NkJk
7X6UqwXRukSPVgpP24iqbuXK7GTWbyOOVQyEt446e4t5tvkoshg4fdfywv7U3yUyxTrY/H5RNWQS
ybSRMUIpK3X9ztHUTYGlo6J6CdRcybq4MwiC9NA1uKo5/TMtaJTulK1b5BCrsb4sGZGJJaf8+7w9
1sHkDA1BeMSBOmB+ejUpor96tyzbV+f+pv0/XRpdigOmwJUfuHndxuqdmBT3Bhnz0t9Kq0X9CAe8
o4SW0sVjHrlGMvCw5tEFtygYs57q9se7wzKOdgSvk8gKc8f9yfykTzMnCyDYvDFUps0jd5nWzsPV
05vWdSUP5sW+iCFLL5alAEI2orzvR8uX5H2pID48LjYtQvYX9Pqsr6ItDJry4aLOFJJmumlAVmrX
IaTIydddw7Tc2ycXR6yL2FJooYyeAPVJgNT4a/BILGCCPAOCEwTHwBfK4VMnIRie5E3lk22YJ3+R
i7gdpitu2Cu3QKPbjdUFSqkgRFe89VopByvaQ+FokeEUfeFiVUWKTNve7SWEvEpVN4onik0xHE5u
gpsPinDh0EoHDJOSEKIwGAzYSC1M0YfdH+vEubvS7sYZw4URZKyCiYLwi1Rf4S/09ydFp+lF54i1
zJMtO/BG5l5C0xgoWdcIJdryFsdxJc58Eyh6qWa0Yav+Dl3Jnspb4AEylzlxSc2bqd7mqiL1yLxH
k6xW2Xdr8ka9TuXvIuaMYuI0SzYn9RWH2c7rjHsrTw1IUQvYV4WGxs8xuWRvpS0yYWD7k3JRFD+5
0lX4Up1hnEQIqD+HXKK/GPYSrv7XqxoC4xpPjYcU2anxOskLQAA67MKt42/CWhEga9itfRTKF2PX
NWw/AmF95YjwnTuiL8MWZQ+l7NfrYdqwTgQN7DcvsnBWDcFXH86GaQ9ZmjHl5PAApLk+ymYV19Aq
k0MADz3roIrD8MBfkPK/HvlM00y4LyD+0W26AfsrGP8tDkxJI977WvH76XZeTVXM5vt4ocgYmwKA
/cKz6LRYePUy6nLkvWyoeKupFSddutUWToWOT1ERuDYAQPZd7K9XXMCqcKPCDpZNLfe9EkpTMmr5
QOiSBCbVnZSnC2wmV+AZp+Egi6wWWSZFQ+/WLpOMj1uos07GMKJnBDqPyKO6eKVtJEIApaH+TZx4
udwxFhJpUxEvIhJIVosPU6+Z17sdjjlwu207Yk+8n2JwHD2dDrrCAtUGOH5UiMLHGXb9e7u6TiA2
T8V3b/8Gaf6ynOmgaesQ+RAw2Xnos8phg8IO+arcDG3SQ6TA3opSSVMQw7vDKuNDJzAT3zvZETbK
kP7T5ZtxTm9jg2A3Og1Q3UGmNCtaWXOZ6rMnqmevSfjK809ykILv+WwCRPP6esiMm0J2eckfEOq3
7NvzZYt48yCz4KjatfZWws57XpBD0RHYPQU8L9dYL9wCqFM0Inz7+eTtr6ThmAdKOo1sNL7GL6SE
bho14eTbb2xCdacDH94IlTivuCF5nXiLZpC6rI+mVUOkiDNLDOFv/vRZuGzsz1TyoXZtJypEIcuy
8M21PKujDUgvQkQylWXLMLhC3K25uUVsmLL3H3s2u15ffguwy2Rj+QlzoNqaPtWuT8CAQEvbO2C1
fKpJRZfJgtqdCSBN9SMJiGp/9jn2HjjojEnvP5Dl3BNUmXkaiGY15VP5iF/mkBQ2eUMwQQsFoZNM
O61EkRICAaTtkmAz3LjsYrQNt9PZvAlwoMtswxZrvZsQ/nIVl4I2lPwDE0iHhqZm9sl8K4Kl71/S
ICcmoceWGE2sYLmPs8vSl9OW4+Io/V+pMG8ZJ/oSoztOxurt885TBmyfsStk966rvF8xvejNM0Q3
ZSQLiINwVKCIQ5LiQAgRqyF7aHyU6WVZ7LiOJZ3fhuUoxWIWKMy4fZIHnv5ykCU4RMI4uyqbXsP4
3BdBG6Yll5AnTkxw65ITnFt3q+YMhjxWBHzCETkJz7Sk4cv0VNv7c6KXawmoDJslE9I40XvwzLN4
SNPjuIByTYLekNEr/GDHsYYRYFU5BxVkzkjhu4jYMiLtngug8qvAKBUDcHSs0YgHGBXkvclYMbP1
ZdghXo+IjPYzW50e79EgJJEAuqIyC2BZEjxN4F8mNk+gBjzkG6345tIGzkCxBT7zH8/PGjEAZIQw
o+ynDc6aJ5MDlVVieCOPYtUImGvBridE1/mxFt91yKUMLvsM1+8Y+gkGsewlJiHToLm4awsadayv
K2gYm2Gou51OgiAPvaU83YLN65es1gIwvTTvm8UhuUDbgxiD64ng3z5NAC9BwnZAlJ6KLxYa834K
4/xxx9tDjx/c/VVooCxxPcjsNbQbY+bgrs8Fb45TJCG66QFoQoFmud7Rrn1JKmb+7qamr8/77af4
f/Ayz6f01YMqUDE3UDKU6//tXXjfIworxjGDi3U8qoch16RxYKiqTdn+WR/4SBa8VrYsWmvnLaDI
QKk5P8SPBgs5iCki+o6xvOhs8g5uR6uQ3DUwYyYM1H5tkbfhK0ScFJzEj691GXexEJ0rVhbcfUZ2
kUUVdOAhJk3tdZP+4PfwWvYQTiaDPRe8RJIpFxzsY8DINCkKrvw54ctqFeBbpknLxFiZtgqNkm00
5ELN0RLNg7tFKiNeIPXfI7C+Y1gWcfS6Vb5peYN0hFvSfLe0jEFPwMk1aVVv0yrRYQOEaVQpQraP
Sx36398NsEJjSyfmT7lnMsZir7zSXZbmE1aLnBc3NSo6rYbkEUsnL3LuNFYcmAuQ03O09wHOmtcM
czBHeW/qQfjA1dyQjnNGybkTGh0eh2M/DH7JARqH5mPCqIkaVab6YHH5YTJe5koBx7nAF+hdtrbX
JkxCW77/8AQKH99YwfEEIYckxtizUpIbqFHyV2FisrBentqy3rOFb0GjDwn7B/MpnkenisGO1h00
QJqwuQdldMAfbFC5/mjPBQDRNviI1JgqW5MKu/XY1rNJcNXXenVyEZSPc4kQngHNXsS7J/SYDEl5
BWRAdud7lTNDWzZN84ElmOZEqrT1TFQhEcWX8GIWPSlB9uSziRBcdZRPA737xFkAcbWtpMDInmXH
ZHez+Telua4jOr4tLD0UKGkj0frsPXA1Z2bDhaxEnEYPZs1OZQ6HiI7Fmdl5Th9nuTuXlwQQPEuM
Oo1wS5JcHrhebDGh5SzpoL5H0c8KrupnWUUoMjf5WSIjwZ+f5pMP59i4UbDMVG0huTkgMLAOCsIc
M3aTWO++8Cbes+6apTSxn4p3i2fJ69balNKYft91iiQqlQoo93rlR6GvgpHxlMBtzKyk28YWuIT0
tVZP3tdeFUcClFfEuY+cqZD3Jx0Xa8pGgwC58Pls94jn+lqQmSQiSYevauGX+hQvLd1NFeM9cv/P
I5qHtmJ/eZH3kW0aNTrg+Y5hZ2VW0XoU+cPonCavvYJ2BgoHcxgDYKYFLT55EoPj7qGHKXVnwYVS
QmDqS+zh3uxYPGmfasBvM61FxZT/j6ngqfgtwkJWk031xa4g5yKMTfXCs/KWblPGsV35uq+zQRsz
ODw7WtMsxCFGoV/Hsg7aD2J4dY6FwdW4F2qkpmKepwEvxfNGal1A1CRfplrCiZZQ7IrPnyik7N7Z
ZTV1UqKoGQ27Aso1XkRmx6piWe3VkBEOAfQb7ujtxIr0oDYh98EbM4fQ3zcLq76NqD4Y7ayg4e8b
LSCpxvHC9onNc+O6mVFl59YQZN3BMGmDj2p0i9FSvDKqnNwXsAvXEsp85cOMHGvypqzRhO1JZEmh
WnhAn3yvL5zjRgxRDufC6SWSMmtbrxXcNOCub7Ot1FPF6mIO3e8AZZBLOeEVGLtbZyCBBwzGY8Qt
sZVj92xSIOAx1tfz3fCxS5020z1/MaktfyXOxoWBiNk5Pr7x8GRfAQBH7tJo9q7mKlEjdSPR3Ich
0Yf4P2b/a+GFltXgTSc5+av36UBL9FMJYpky2UHFhB+92iiYRuXfleMO0lZ1yH1L3NoNwG4m5H9Z
U7LLgYv5W0HF4bOQdGcQ277ETGdftrp1Fy6i9HrZxKOUE1NYd+FzETKPqVw73yq/vQQu8O0xABhC
CVUaekGlX5DpjpXNh2awbRT64zyvuspf9ciAkOXbRoJMkfCVhMO4k1xtgcj2Guu/2o3aCrNDQhqO
FgxDVURJEBllFTHznYe8kD6SC/v903hhm2nPBXo3kb4l1y1cMhjSkvSwOUEL2xSMdgOcZbfdNOSx
Wv4HWlxmAM2OI3kMPJ3TEhxp7NDfp4pTkSxEfRQIQfm01uTr+S1rR5ODbR2+KZs7jJPHrCLkibxZ
OEkyJK6zGPcqzevxEErV+/fxPtA/gqKmBQsY9E8loEgTaBX6Vdef9xEzuYHGUBIBdMWS/GFdIDOc
WtOvfFVoj5SZA94bhpBTfpKemAzUHtKJju6LTCKE1SJjLPKmcsKvOHGL4/Ein4pQXJhjmq2y6GQy
DAqyIT9lxcvke1UZaY4uFHIlZ7xOo0mYe9PeRsHXHg0AO72LDvpyPmBCZxC9yKvofxscduOurxBV
k744EZAZvPZLDXxfotNWTVeD2JlzpEsMwrqQ58tuLx7HRsY2WiEZwJeqty39WXuYFKeb64tjbjS8
fS1QGlKL/7mxq8/jdhgM0DfaGuXPFWC++NL4xFYstBWRHwLLdWdszLoqvOzldhdqTQ1kTAiAHdBF
7zk7QwXYrztY2kQ2y7PzedyFGZJoii8CLQJoVTTTTNZDQgxmE+17IuR3Y59dNcot3Ys6i3q3A1VQ
XP8OQAX10/iJIl/7t7ZCmY+Cq79PZTpm2UhDS7E8PKmkcOm+bMStR/yEl0OnbFWbnkjk+A8Suf73
c4gBjzZn2eOqZW04Siuwn4ZxQ4u29OsMubmq87j91oIixYJipQv5cJl/m0rPi/FhFsm4a08wPQ8W
ycoJ7PyoeQKjkD6qvHnzvnPeajFyQiRybAcnZ3noLzzGptr6XtFchNJvhokNqPh4JJxBoo/imvMF
x4fJds/+MKCBzxd/VvzOyrhPRHdSWc2DmqiYyOfcyJJhQBwLB7Zmj571cUGpAcIcecK6A/U0xwX5
2bN3E93aW9cUrYOh5j9bI5XSKdTnnI82q7qW8OSIQ5Qqs++hwm45ce1ADgmz3CR1UWOqBoHCY5yJ
PsO/+2lFl5vAzGQCe8ASbF+8Q/XdBO9aXmLSszg/C+2rgfr+6h8nEnoCOWLczKJsg6ROCTwIdlYb
JPJf0ok+8wg2p8ly+2sJeSvS6DkdL5Wnt/FPFNiuYDC4gCWRQ/WwAQssouzCZbPQJjTiMAQYVKlQ
Mqh0ddpTXJ/HFmkWw4q0rWq22K/OqteWKQixXVXovDYrmJ6Ap6vDBded+C7DUXJ4EJKt41K4CQIO
QGOLaoqVNFmSEbx5lUtZSTrvLkQquT9vXUdlZoteARwp/jraShuAW+XxQl6Sqg5Di6X8q18gqmPI
Mgmp+A3TxViQ42BQtcbqKP5eAhphg3wW+mt7x7r2t/TPQ9InppHXDScdLkUzaXNP3VwPLcUo5PeJ
zRlyOPVKV6Xu4mCkT/hE344taCUr9TlkkF2gk805l+M/tdG80ur0/AMK98b+GAikDFCIvRb8nkBr
TaOgYUAzpOHPM/LU8xL3mep8Z1z9ERoUgjOwGeRfO+JMF+DiZYLcoZ2DQKuFZNX5LhjCNZ53dM/u
wYv8Fe1xPW7kY3d6E8mRogjMXR1EBErrNxsWgEkcaLgmCICrFGALBSkRDocOl5pmfIuxGJsdSM8r
przryvzNJp6+1sOZtnmNVAwLl57t35kZ4e/fiZ6fPAF5GgrUrrvWE6vTzTTwUIpSkTdU0H1HAzPi
FqiaVcHA06QRR2cPBhCcD2clc2a4op/HLtRcb4c5hyMABmqGC8jhwfiN+FBxytS9CgXW3LwIljda
kPu+L3+Q6KCIbreTFHZNrUBAAm6xd+9iwcPgN8Kk0oOQfW0hoi4clV+82cDdM9cDD+/LOGISdjZ4
VhqrZZm3kis1m6gvgfwu7YZ5Jk3LFpOxBJT7hHRDscA3ps8LmD9KGpuS9t6jfNo1YKBQ06A6nlDb
4gS/ajaaJO20dATMg3ngiDjyCZOdc+4/cbGDrW0EGxQ1yIjEtVbIXacS5oyh3TSJuQFTS0a5stdp
qqJo7fiMw27CgYnkROq1JVIfRso20S5Kkl1OCbOmOjvw73b5l0EuYg9KGqEPyV3+ivEzKAOgstNb
6My/EPVqJSTt0xuYge+UdwqWFHLTwOmnyTwR1zJDJBE1aTnSemDXdDIDZNBpfFgOkHYd/g2iTjp1
sFl/XVSP5+UOQBa60ulnNizwbo+9pIyKTe+IM459dwKh4QVyKrgczI+EjDNxXv2S24HmVycNeYKF
NgEEctf9I9HeHizD2/huZZH+Hhjrl59NUz+idYjai/0KlrAC+Pw1yaBJb30zB6XUsKPF+DQihZMB
/n+Nr+HCRLKUDevtNjg9dMJsWfbEZYPXQt/uCj0JGE5KfVUQF6hVvslzM2s4gvQB3Lsm+ozxfkBW
n2MPCgqpettQom6raXgmLVjhHMQzzC6hFVWS9oWK0pvQOKGhsBAXX9hu5O1GFZ3Fb74RAaKLfdYt
5fc8GJmCYyrL7X4GLOJLzvrb86qbAZoAbVAtD6jQ06Osxyoe0pBFNUNdM++VCJVuJP/giBU5Kww6
Pj/8oM2I8iyTuRj8lEd7Y/7oVxLjYRlF53C38QyJXRmcU2GU3NQizzGyZGzm38ZV6E/pGw6heGWx
Evld+XoXTd84RVk7sdshhEv7pl4BHtCuJbJN/rGmfigxLYS454JOsugIL665JXxqgLuiGBit7v/5
AAszU8/TMpPvzC2KJEeQLyHzX9x3O6rB34gOOLWXL+THxnTEZ+bCOCWbN3X/cQr/t8a+omNlUl3w
cI3kA2d/7D5iSfgUJZypNdyNqtBdMCRaqwhwa9qg+tE6N8pIl5gRvMIlB9Dgmyvha7cWg98jFhlT
M1SLtAu6i5kovPVFkXCkRYD4dLkj7b0buuL+xvkWwQAXZjAMGdb3jg57a/+wNS+vz3j4iSpcwJYQ
Y0RHZL+jjnr0wmKKH21vqthEd9y23pBfCApGaorfdkNVQPY806uXIuXw5Q7BSm7MMmeKVd02QdtO
X6srq31EChb+6YFv+gWto0WzCh3aPO3U7qHlsGUL89kXxeABHlyaQ0Bwebis6+w1XEANxpc/oeIU
cokk/b+xBXwyNnlo6MOPan8671aUFSfRBje72oqhLo1Bun0aC409D0SDdXLMdChZjTY34kR3ITbY
dXarNcQwCmUWzP5KTeGu+fAt5XARG+c0DYaArXcsSBocX6QAsGYP0aNIo4fKDe71bt3xM2FS9Rpg
SNugOMGq7Q8mu7rK9cIoJL8EDugkgGmGMZGoCVK+LgW3tivQyfaGn22ekaTdLMJ1JKU+U9uWFORA
HG1HCtsJsVA7KR0fTeWNcfy7K0BuKRdivBaCCEDs7eQIxc1pj8M0ALJ3FasmVLV6Yx+3qpCzPya7
UJO9NzjwD0HXYUctn7ZbZOYQEnhvEZQw355pnrOfhMocmY60gVH68XJR8E3DicxI9MMAESrfh48e
pj9zeTmZOKTMMyJH/dxQqpn2xMvEgGUIg823t7vcgJ1YZJa0d8bdzVEMvBrwU0fwRpnabKVp1Vsk
8lAqWNhw6bTSG+Wq0DDIEOKM2VfZ+DUkhstfT4EIYXFH9LdVugg8dx1VPtHteF5IQi6bk5Hqo0XD
x/oX1Qn5AUowjkwCRTv4R0AZVDaLNLB0ykK6T1cpElctRxhgOBpjHTFf8nuYBUSskW+F7N5dJVv2
srW+2L8oTqABUSxDN+AcsIOG8LjQ4ofQzKkiXkZw9aVPbm/AJkm03yV4//u4VbBkj3cX1Gz55agb
AlnlLeeokHpLf1fpeT5FqFeOVSnGlO6GFVXPNwRDgjBaivHMeMFeURMrKtmih6hbqKTs2Pv5wvwa
WFs6F2643Q01GWANJWr6LeEnX6bVBhMDTgLOQfMuyjvwEu8A3rwSyPPPk14mu9PGV1wL34ALCpm8
9v1yFRSm88LyZp9/gvOSFZEhHUc6wLgW3jBcQUm1bHltQbBnqMq1ZXH/WzOxDF/mG0CIcZFmifQ2
fJ+ZmI+qNqpV7FxE0OI4nj6F6pujt0C5puiC3FFjqRzATPB5rS29Ji6iYqE5sOp5spJBDcXo1MJg
ZGuPshauxgWQoy+BCvwaRdfBPfqSAV0IsKW3hGWxxo8T8pE/MOOfObnzYxFJFDBI2/CHpnX0FtoY
jCazaw9+F7RPUnQGHQW9Qprkt91CqNoAl9UBzbsccCgKmQJIn+ZnATdkijmd07f6buIhP1zeE+gn
FZa+Vq/fszI1ffH8W1iEz2/Em4zqODmdOweufdVAMtt99yhGv6vReLpwZtCARmIzZDLwO28CxQst
bWmjGdNV397ZBU2IkvvBMdaLK2fUYxHJmYDDy0IGs8jer4OT5UmD93zGbt//GgP5Zzz+rRpHhQeF
OePXudd0l9+hNIr1TfAUNEB+PhSvXPMxt3A8lKSPS05vSPuPeLgwpoi8kjoEUKWny8lmbzIeDqk4
sBdCWwReUZxFXpRxo55tb3uZX94xZn5bZv46qveWbM0LpP+6GMQYXiEaqc6GgIZIQNi8x62j4O7q
O3FX6pj8YVZO0nG1+cqK2dHoJJDfmEfyyqXF6rxHDAvR0cE7mHtso1L1gLfWtrCje77erP9bNNVi
gOXVMzxal/jOpaNFgVUIBjqsuF+xxQPAmUnk7U0/wiZ61T99soi5meEKisMq9DlcT6Lyp8HgvXM+
MHMaIQegjudIxIkews0gi+M9o9tL9/j0LFHailFTA6VBURgWZZdWuwLpAnrRtxwKzoEhgRm1LHqL
4XnLOYzTokrhlVoRpqxxnSyUC+tuOpATTDItQxzWWqH0zs8sOgkvOLFFHeG1X2TIVi3qYuoVQ8sc
tV8A4NRJOCIbUjo21Iia17RQXuYS2+Y6/sVc1TWFIv1DVTLOPcm/pnFzv/joGPoh716XgAOkVLTc
rc/GhmYClpdLzMbfljbdAyBD9wgtVUsShhys4cil63FkoUFZ6TTU6qKClcWcfko3lLMYH9jPu0eq
AfagsxlEjUwigJOgTRNWqWvdWaMmq6OMS2I7zHquahiVfdJpBllV4ZDOqTVF8NNEz7AIbgEUgot1
VyEvwUQ9DBDbkAzv5qVhZjw4NM1SpEwuxGlw7Xff6pwOZYDgkqUg6okov4qojsTIqrPPy7qUHvcL
cX3FdE7zuyQBaIpGN25K6gXgyYbTmGiVgVuaFH4Hb3ZIYtqYHCnD6f2dev/XwNA21mZ7mqgt3AOz
K/7ZtV5Ir2BtLvszbLXHjSnEnUaPclHiV4gheS7kG5mg477eIlsXYopyRcOlPc3i0k0KDySI9/5c
ydaAx97lPAxbsHNnHb+hqfDDjONNUwBHPecbxketYkZpXKgVU+kUse13vEUgNVkn9f0jA25Zor/b
bzvQoEnPOX+LSQmIpNljFOKmwJngNqquH59qaNk3X5iKPNinXeWUG9uFSGy4U5TIEGD3gJnkcdI2
mu1AHaEYagN6vsUnVxGC3O4Y6/8VdtTmybIb2hsJ4qAHFrDZD0XYjOveH/Ygg9dZcnrrO0LHFKhx
PjlBgph60Spg+LBp8VwYvsoJ/HAwzD+o0/rz6L654QF7PTR4s4nBMKptqptQMT+hzWs3CuLKFyBH
xcOoHrHXSQSbLRZyW65lBESO8MI5hGJoFvgsuEsHc9upCcniynOB0a22Kz0ysaFo5N3jHDMBVpvS
SnMbNhnUScXQ93f76H6L3B6hQJRUavqHM3i5uf3ppec5UYr8/8E7MAhopflS1s4LWhldATd55WxX
OfZGkl7P56FXYS8hsmUZ8pBpqMOfH5ICLYT+duC+99vwFmOWH0dRguQkAsAX3Ds41WQGleASXyel
9hwSXX0sOEJ7YyS0AYgsF/xxQcwgwc0BNVoobmChmfHeKdZLuqH+YwHcu0r14F9G3R7t9ZZ8e3X4
oj4SbiJX132jyxRX+QoZeO0HJjXSknHuBCyFcCuNStL9xfnXR+GiqD6oJXS/TS8C8rTxOizW9RVm
93eYinwp2QzaUlvGkvspbusI+ZjFnuNh2ojQCVk+rEjxomryFGtR0/aP/+PGCAHiTbYjOx9yYgTE
gN6tmxbZJkNCoG91LZRNXxmFsO1UcTCYNYIFvRhwAO0pD9SGlH7Y87d3beMV4VyKo9FlKR8k62qz
d26DGLb1OGtEO+KMUNDi1Wx7X6teH/DAkehEeO3xl5QG4qRJ9CRMP8rAPFzAbU+OnEWcI4u8EpZl
0Cp1ZMiS7d6Hf+zKoIqoF/teSPIl/MpNndFPybXJDmauq6ZOh2W3EkP8bxd8Bg==
`protect end_protected
