-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BITHeMA/PnLXJI37UXRH+IqLSykAtbgirG7LmlXG4f+EidwW6LP1vdB5fGRaYXC+
taTBhF4PD33y2twjZ+yRvJAE8xUY+elsB9i95dlERsINiGJMv82JWfTYByJHOHUD
U6kOOf70n4gkjsruVxUCjdHZ17U4CKN8PALDF/FAnI7V0OkUOLxNvQ==
--pragma protect end_key_block
--pragma protect digest_block
ySJG3LF8/GsxXzV4nhdcb9coG5Y=
--pragma protect end_digest_block
--pragma protect data_block
uAY7gVH8RgZpRAduyR51sk3XexzicYC/+CEoxU8MD8CY1rFvsgGxEDF+yUF8764F
W35c0Dvuby8J+4V3PUwGefb7Qt68wQg9I2LbhDcxRb47u279ao1uAvlFR14MbzoF
cSozB3y5erTpzunTjGBEslWUeJfKzCKuRFX4dqP0ltlVi4+YU2+BNPb+85IYtZnt
99jXC+s2efKuZabLags4MTTuVuPl71kgT+GLQrgMvX5lIjru1ejzoPGD0KLiqqp7
ibiPJUBkNVfzI1LixzdpDp3tevcuehuf1BhHScNEzYFII5qA59vamQNEdSkCuIok
SUoBAVFVgaqAe3mLZaD4Y4FC7IMlxTheazS80Ut9z31CpYRWV6T2jk4P8GUPi3J8
h9AC+8IYl5phFXuyK7Ir61U/xvfo0KhPWbCpZS7T4FonfhDkZV2eH0d763xaXewZ
4zQLBorI910/Jfsc6/RoN6hzqtc7YAKj1XqxcB3WGtnI/4E2yXMCb8Ic8TuT7tCM
yTu493u7lQ05oKFYmUzMOSvRJzGgzSq0A5mpQL+sCBh+JydSz4gzDO53rscK4ZvS
geF9t6+ArouFxtMiOXKNDh1OwE6s1nW1aCQspwDO90mk0KdWZ8tb5h8LKpJ96Gkk
e4ixO2v2azM+RPWzZW5wc8TG5NHOc/qkzPMXhMRNE1c1XD2Lpdq0g5lzqIyomfp2
5PVlA4FovoQhkhq9nZZIqBQyKzo4CwNrIlJxi8/mw/B/4S+kN4Y4KVw/Qn8T4xpj
kHyzfBsAPE37LHvwCcZWIaAqXATNCh+5ogcXBWGyNZktdXvlAQ2PXbxyohNCf2vC
jNjQ4uzvkgphk7Z0p+r22IGETjAGIWDgPQJdK8Y/NtxJATeUZJ1AZ5bKzEWRevwx
DXCxLOeSytreebWStu/MVLG4e6ten/vn6JjzrV+gt3yp2l+Gkvb5f/Yj2T6wD2vv
196eyE9NcxTCx51/LqTo3Ps7x+BzFY5uSs0VwDLm6C1q456TljXHQ2BX2CzhlU/V
5DYI2WEQAK4Xqzmu/ZfrljITKyGf5GTk4mvsCxWY7suFBe/c9ZxwNPyDD+LXXqbW
HdE67VC4jOLBv9F+Dfk+kviYQJdfe+Rxe86zcWS+WyaFvuM/EvQCauxspyCMzgMM
7kn/z427cCBf/9oPG49IvBMxxqBNXzLyqDU3B78NmKOnUiaeY2que5K/u0tv6btY
sp14StkgSewB0IsHPc3Df2jwZ3z758mCqA7FFHliYHjGjRb9FEkVcADUiaL7ehL9
ZFAl5M0bLMqBT+46LKJeUlDuZkosp7RwVNxx1JcUh1rPpg7gPUKRAwSNKoOr8+zX
pw02gCeAeb9Zz8v8a/yQf36HBC9H5w0opVGOP8SrhB6YOnYCn2QwvHj6wg7Esl/x
rscK+iGlHwqogv6ljo3bLJCD3XQLMhgOn2hT6ami22mkqm8V3u+Sxj420SdpYZBY
vqYllVnF67NqTpk5KdevwH9nirM2vfw+/8ZTiobPDc0yTmTaFdKCdKPkiBAt5o7H
mM5g34VpNHiA50duIoDna0BsB0UwJalEXAL+n7tPNnHzwWrXxaFTFXc3qFjtygTH
Sjc52NeJ57y6OfTsFv1VRCOb7RcNSWUvQZDOUPF1LiaVOxxcvCCM1a8fepOwiiW2
CguFYZPB1IE/O/8TZIoXgTRZl0Us1FLD903SswfOnQLTfQoFjbmGVhpIxCdmzH37
ZGjNv7kBrHCEz6nBnJRStL3wvzp/abFfwfILkwoyKrWxa3hE5qlyY27GZA4hjDlV
oElHwW/uK2Jz4ChW517EHLhUZHV/VHDpAVQhUinCDs6NnfM7cLUUCyLeCtPux7vw
uBtbmJdslhbY+HWdQz1XyMEr8KHhb+vnaMDUTbzHdV4I/SaCAOJ2kF6W/G1Kexnk
jOtY7V3txywl0ZPLRb19Q7D5L020xl7YlddEgWDB9cbNhYzArTZxkwZ4wwmTfcVa
h/G2Q7Wn3vvofpHzdFsOs0AjbsSYSJ1mF/XaF0g9wu7jhghRTim89hbYn9DpM2lM
YYSqaXZjB/A/ETdYPn09F1Xpfhlf6xE3AIaFOIMrtdsSs7gRPWflcF359XgvT4iI
MMj+rYV9uA1ih6E3LDYPMmoGlgPxl5Yx6XwAXDd65izNZpehaqtc3I0DTfeg4DJ1
9mMdBmGswtIueaI5ZgO+bYLthzRIuvGJ9Tofnwbsvxzrc9cM+JTKcLnV8oZZQGzw
RwBpy5SXk8uijtdAhwKtcXP7NP91OsNP649I4kc6yfvMsvr6jGRxDaLXGFadkBXL
k35x5g6XlsXiu/PZZF6IWYKSBCj6gTvJ84sTtw6Tyk/f13XjYQ5qYLZBpW9SEEaO
wjMe9V5fnrz4kzm6NWot8BGX010oZ2f/lGa2JIghBRoXY6hT2nj5Bv33QampaCdp
GFdLTgpixwvFF1pY7Hiiy0BUXmQZOmE7H6ROaglAfGERYonHJAsKXHjEt0g94R/1
MUCo9urM+zR0wJ6gXort7fyJgNprx2+v0Cm99xzu6s+jCHX+endJD4BclQ/9S0qH
2mTi8T/Y+ZfbL5eGp5iOaAn8u13BRzEzK2qMDoCQUwIb42BdZ4EGQf9nSrLdQW8E
HXJMD0VEC4Bx7stSRO2cbSNeIaJXmnE7lCRsdttdKknw7tTLC9s6HI05ZMNOsyxL
ysmwaxE2vKSelUvayxN2Euso/8HlVGC3KYSbqZZpGNKAbdmc8ZpficP0UD/Er0an
P1PMEU72OtDVdF8hJwHAdu1heaHSSSqcLoNIqrHIRvAGwFixCPFSYNaNiUPtkId0
5f/6P9BHigsxlkCGT6Xug47YL/Om5ukLn1gzAp+sirUbkVkP0Sa5y3o+Sh8i2hns
pqF9dXYauwShmuwa4eK8IUcbiWLDYZiqbtvi0iPn0t3X1AECfM+Jq7rNMqXlZmBs
0Wz+uqVp3hDO5iehDAkRc/PAscgJAVdTvK23s/ABHx88FY+HRumNjLNZ7EGWkq1Q
j1qrETHlLVTJae8+3vrMToecroTqrvBXXQH/GWvd0Gt2mDq5a4hyZsV6jnsJYwAB
Pf2Ovl2Rl1w+CjcNuyXgxEMo95wcOIWiKWg1hvSrkzOI/hGU7nUEEIu+vmjRQlP/
gZk94QIDOWHH2fx0IlC151jo1lO7quN0m49C4iVamvdjiZYjrffU8TmDUXi+A19i
krNFBtpk32uMMJRcDGZmFvwV9QKm4dr+cqSQ3q6A1kbQWZLCe2ls3jFjc4+3TNtL
ryhKgEqwLys+Y8Ng8hCdOnHAFjNZiAhi3Bx3OyO8EojzF13ZvnOBGknziISGh7TX
6T1lqinutf0usPvtFM6WcLCQk/ds5XVm6bU7rK/vcy6fWdB1+lIASZwy7crNuMgL
+0Rl1LWNYYVoToBSrEx3SlKdn5aeZO56Ke0h95B10Htc1Eie34pNIN3fh/rbcetD
d2pyQUmk/evvfzLrnXMR2Dwma7ZEUSqA5uxOqS7LLJQTq5v53h41BwJOYjKv3EUe
LRPnwx9+ot7e4DUWM9Zaedq7IqUMUrSRfqHstvoqBcvrNyE8+ukIUB7OZEb/EK8W
+Yl020AnIXq3B8nYyjLD4zJuuM2ZUFaSIBglvFNFTiO6fE9wTjGQaicHwuiVcVAl
5uCFy/L8g/QMnv0dVY7tXtGGbjLRqL/s8c396gxZZ2VHdlfF8GyIfEr35rh/n2gJ
fMRiq68/r150/0Tf7n49ku5Mi5jBUJuh8tSjE4SVab+W93X0sjPTexHuqRSrzMvd
6yqvxI4rhiaCIC6jMxDSwYk9vUiSQXHRjRKwRD/IkkQ4V0PXvzn4UX2sygKbCFtQ
4PTXjzZ6VUsYWymAEJpbReHYetudmJUeqNzzIfZ59FkJjgBSpPtORloARXnBN9mh
r9K3FkZ3j3P7jT6sY+9bD4M8crhg9mNO5NWK3OzKCQu1gl7rV6YNDwLn7d1wX8+Y
1zVrVWBIz55afIUcPqIoT8B4I15GyRmXqg8Rq8dSiule6bOYBafpl/RrzqNaFx5B
XSyhWllL8h1Ts/C+eWPGQ1nhHvr86Eb38JXFnG5/V78K4Mur+nulUTIItA6B7986
xwOu4xESLBom1uR6YHdYscwQ7PDLsrzN7fnVvig9owvrvFmkYawbgbHry52De6ja
jFV9r1Ir1SYkTdfDecxTRhzOTbuhRZ9ol8IH3KHQgOChcE0sDZdZlrSdih4Vzj50
tfkpZyAzWJK8aavvD52rp8ngNXv8edpm7oXceWNFiZdWALI00tu0eWOwGKxJrgIe
ZLQvNMwGfT7DDrVeUTQN81u/1W8S27H5sur5cPHB1Cv9E2pwZ8qWq6H/771pbFTB
9lP/xh9SuKdPJQN4Z4mZZVHHDF/UV9Zgbbj87Bnpiafea8ZK315yYYt36CIb7SJq
VX6MLnUhYwIHyvnFIUUmou3Pmv9iljHYsmaaZcbFNxQrofTECwJp5R7VyYXeWNNc
fPaENqdT7FA3L1eBqR0C+0Unl70CWbXBbb6RzFFySV4wekSFC6Nsopf4FZMQrxcI
+j1cqW1lDVN8EFlCn5rmcAiMdc5oy6P/3ei4m++7tw4xdk40fvAvsFY6hLBZJFxX
7ZLbtpEJVyynw5KpMqOpNs2ZwcOGAL2/LvcMDI8uuSuUzC8z2hkRK2XvGyU+f1iN
GuDZvpfGvFbvrJWOn3jm/z6lhOEpf+iQRG1TbHJ0DL/xmPxfqVOcGLfYix+ET88l
2/YkytBbvmwhiP8TJAlShI51vx3vkJJDQ8qfnV62lT7xewMOn2gs4X+N5W1tjYaG
wjtd483u/w8sphHF09Z3nLPa53iJIN3sludrKbFCOeNYzFRXcrrFR9SZNHYwQTb3
UfyXR1n41bWVE2XpNf1HEDguEmCxe6JJm04b/uo5I0fm3luE/2HA+I2GgyuqsPRH
o3wzQlbsPWTwAL9QHZCvgwAgkjJxW2hdeqISaJ47MSTH3XistXPJB4uYvF/0RYmK
6ut+DFVknriS6m+g/UAypIrTH6sBQSQkTLRvChVOKPdBaeHJqMGZkyUQAUtwguAt
kh0PaONopusZ1hpPmhM0u05vt5BaMO1UQw46SG4yIYZtardMOyS1nitnt8vo1nHO
2PYuP2tMa7Cp7wKlMytzupY3texuQ5sYWxyzMMpcF7gA9qsYAjDYK3v1MgQN6QEw
1kQDYjvwPmP6FTRQftCZ0egPLJLVKtVqVM1Nmhe9eRtQxKshnMvb9nfBIZxtHwm+
9WIdEbQ2fkMsi2yCJTJlJct/Tqm7UwC4UV5HEBnnCljWyaM40jmGaV+vXyV0Kfw5
s75jRYrRpbexqQTBede1g8hVgO8hBbYjPjLoSsMDUU332hCfyFFM6vO/E7CoqdK+
mvJIIF8PiBQCXJIzgYv+zJWN6uD5yH2kuBOdJdx7FD/6r+2uNL68MU0Ev6ypv4ya
ss3mCikH/7WpAmV3RTw2xGhDuT3FUFB5Ku3Or5qx85w5hffTgJ6M1CbBmOOsugFU
DvJ9wMdYQHRCVeCUq6hDezOf76fc4fC1vSkQS4bOnKMlAABU+53pVUkz3B0clIYh
in6o5XYJcrlst3R64oEEyGTvKP9Zt7ZgvItZTCIC+kgvdoTjn3yK8rzB+Y69N+OO
2svFfE/Q9QIlpVkHK4VLvUfs0cPDyJ/gN+JPLqQ8pAOAueSj9+fZwyrZQXc2Ucis
e34aVel8O5afILBNvI70IJwFKJJXhGjDggylyw19Zx6DFJ8ehVMyT94UyluOwUHF
w5CzMQHZcdUfLQD0+WKw5GACJJwdjK3MdG3ZJhZUd/MBXvpLbkt9ak/DACBBcgzs
8HKSi0hQjwG0MwSXsf3ttbGZJqk4C4wTrcQudGM1bV4kMJ7/45bzBn2p1G4u/kEC
kTTq4eG59cDc4ZJE8VwQG8a1nOG92+FLRsSmoKZ86lWdDEDBh1oDhRVu4vpl9frG
B9uTv5/4CW9+5rO93GoDOYxyoGuzKdFNakd/Dyb0BfIL9xVE9lTXVbwoZvAYn1eH
zF4ezkMg+VzWKwA/2YsK28bNGjDNRYGFsSoRGWPR+Sdh5lm05k7swDWnG5qAfaLZ
gLAj6mZUx82R3Tr+qPhhTHAjwFxjkb/njbKuTgcfnDtJOXdidk6eGb2QFsOXo235
q3sdBTan5gKYN8dXpv2QLxNVBWWeGOyY//dG0IR8N9nA05dSy9OkKwbaMiRI34dO
6yCA40cE+PuhqNg/aDmGlqK/ZtMV6IG17mNyzCtTavZewmrcRRJcYCUoiOwmIc1r
BpHQVTglzt8LFdOfqaLc4RkSetIbZVjpDoNyFChf93D4zV1Ox9kiDWrl4CIwEMRc
qjLCkZHPGOA5LMc2b7K6TxCnIEosQqWqP/0T6AH/fyjzHLsSMFTNjSXMUY5KCd1E
gog8orNhF6JAzs6V4ocOPJItlcPQwSp3B92TzvGJiTvZLRtI0ceV4qv6YJupnWfk
sXjNMugO1GfhEQfKCmXrhFXcVqQQP6GXD6LN7oYj7O/tYheuNfWcLK1jE+cyEYQ5
51TmBKbNgYLZ3o+R8PkCz4QTV/tLpFxT2hP2o9SVKyV7l33of74se6aRTe5B//0p
zeL1YvRLLM8VWjzyPJzD21wwrl9gZlURuxEOAfsEb+oe7GhElV6rEO7rNnf4iK1D
9/iRWMwSSGvKIQlwjyQ0PW/1UCyUggFW80UxhBcFDrU7qjTW5ybdydjPn2nesdrt
4GSd5SOoHiQS+tV3TA1VwR4w9lKrH7N3cZB0wWdDxqypp7dkvfYEO4/uXLTZ7N3C
b0P13xTtJx2J1touK2J+1anoaF68hQ/Q+2i5rvdJLsRZznGaVRxruQM8CPils73Z
RMtvpRpoQU/EaAZbr0in9cv0xBNheGRm1WC5AthaGiEm3uopriJXTZzRNfaxeqpP
NjzqITEF3CNwttwOPDX5lTCAONpsSF3iur9jxNoSLgejz9XBt8O7QIlwBKd89V6u
lZqg0+sb/pZU6EXwq06JHhq1tT1UFnQVvxV/qtCNmodEc+8b2VjvUU4jcW7dsHqB
+qaWW/+VNSQZPVUE7NSdYYlGmvRKNbXFNQc+9bfRg83/SNGH1QzBC03E/wRoNzmT
YCx330sXW5yZfqMEVQ0syp85y773/iCal4hOloHtiaL+Br6n/h3BiQftoGsyj9Tr
la6Hq/uREFi6Gt9wKQVA9JMvAw6PXIUIisAcSVd0Wx6jdmkWKGX8aDSMW1/llq7G
8x3nitk3/eV29BF1URt9eS1KzHTrnOPJiQAbiHRiQWjijpZ9vCIZ0ZYGL+duCUzh
82cONpTn5BbjcK6f3CMEg/GGY0l5FJR3UQk891deZ5BdH7dYc8WsqMKd8luEaxuq
sLcW1Xfcu57a8994z1l6HTgiHkXiobi0wqmG6wjHsNxSug6/x0S7f8qGREXtYTBj
Akd3NZWIBbK+XsoXUgbuSIGnVlxiDGdZkSWFWU6x+mm5oyXTOrNlBMbFLrH/rI1I
NQaB2bYRoIdNhSr0NYF53mwqpSVUX4JMS18jUux/ch9C26ANsABGpa/IgV0CD9dr
/IMU36ofbsVYS6GAmpBzknuNgD7Rfc57yApXO0A+Ht8oAJavO/8+4xpCM9k+1wAM
Yit1tgCkLWy7iu4zGDsv+enTVc+cvcySNclXquj3QW0seYMxP/4TpSJLxIZKmGuU
VJ3gOKUuJ8Ggr5JMklAhRoXfTLbGJmJ1mojaSCpYY655ZKA8bI2iF+5l17Q4Z5HH
K37Qfg7bnV7mmVWSe1JsxzYNXDP4XnrQmS4SK+921xDmDUlnMIe214Qu/JINBx0L
C8dBOecTOwyYeGkcrfqaMeihy1OIzhVbnUNfozSvZYG8OQ0k7TnstkVcGDv538WJ
iG35IqVfadzqajW9G+ud0Ej86wnIrUZJRB7FJe2oNYboghZiYU6wW1Gw3TcrPtD7
ZpRzKlbaen0M4PvXg04iF/Z0kE2vfGTw/BheEPwJp83gTz6CLg0keUnWwbVzrhv/
RQayr2OP3eNg1oSjtrPjgT6A6jmpq1ll37TxZNpE4xzWUoLcR/tPmMIMV8wY20pf
xjvbWI03osmnxO9AEItAJRO9jRLWqnFGVM+UaaTKEOHDGXwY03KOAEmoXMdNA+RV
MCEbrqLxQ3mKpnvd7LFQ95/a0DBhiaeQkErAluBTjf6zIQRv1OcHm8kC8TtX36GK
kzAgvNxNknYTGW9fytzj9ptkQDeoQcbJr5wDN3LD6Ts8WjyKYyDwrbAguK+PHHBt
zS5gmcAyEy/sivn1ZequSOvTD2c86oEpIovdHlshbojMNjtbfQxzRkIGcr9OKX/9
ZRF99F/UMqZTAA9o3HzEf44YtojDkQ95LJmF4GRaui5JvJlok8iyaaWYwT0jZQCY
2901DlhMfQi7vfyzqC+0e5cs2EiGmJZpMoMJ4/c06IdIlsGsbrKuvQ2WvosknE0G
wnJ1vUpJzAZC3YalSoHabmfJ5d6k2uXZLwN0ZZJ8dQmDJJgCyBAzWwVRVgnvfFTe
DudaA3Q0XGa2iEAKTcNtkBJv38DaGGLOrQuLs9iWdzEQU/QVzW5Qmnfdx7V31jVe
CNQ1rU/w2851qvg4nt7mndHn24fa/Wf9dRE+Po4m5sfi0kaaFj8CcXuWgFnA32eP
sIpL/Ppzj4cTN0kpqE4rC4NZgAAWrCOtbrGvfz+W2kSm/OrkIjtG7e7L/lURcngK
i68VDrihtOy5Nwo0Bl9npzQm2TYuybTUCuTLB3rIRLbbqy0FKQvhPlfRSuXSd7hz
3qUSgWlfnZhSmfwKavX631vl/4nj/0J3U4wz4AGNmriWda0dyMLiA8VRqDYe8tXz
NQOotPF0/lr13SVhQ26ub3F4AIe/C/86tPIkxOChAPVYO6KJHxmoVV4gsqnPITFP
umNnNm4VMq1LIJTepYmVduhdddc4dRvcw/ikS5gQjPDdeGcSDHJHS10/FvA445GU
Z2DnkF9roq63cF8RECPuMdr989xz8CTlLrhEI3x6YZ/U5+Re6yf7xeVnHtq7U8LH
lH4hmCTRxA9qURPHbj0cwwNfQAa+uB1QYfUG8BPgr9tJdAepiMgvahhMCVUP+Iio
o5Qc5nn4dPhgdFRKAD2TeVYKo0g2MD79Ag66SFi75TBAAGG9SS3yH26FHYepEy4Q
cxmx9woM43S9yj9g/ZVL3AJqo4TuuNobceUM3LMP8qQH9f51IEnLtlJZ8KqireDY
Viggi1Iea5J0r1Tee0T/bYBptvpUe9zK+eEcyi2T33WX6V8n9p3rSOYW0LDWSvQd
OTKsZvMwASUnhN1syGEb00R+NSLRmOM1EgdtHvDV/a6BrKYb5QnmyGXEK55jJPuO
4IY/W5kHh6qM1XCNY/HjONshU2suIt/ymCjEcZm7rubg2PSG7wA/nMm7QTI13v9A
87gqSHtHAzCfzWuauV37UXcHxHBtXKjoa2NF+oai8qfqz0B0e/avX/N975p2Q6Po
tMIrVK0fNrVpHBxvTlSDRUPzMfLyzXYf5G3JsCM/C+7QrKGqR+MVe5z7Y7P8a8Sz
xxa4B+Ls0NVYhoNz1kbjVsMCE4jFHlg3Sw64m0wLR2PN6Z9XdQY0OL4J8Hf/0rIe
gzXkJowJCj0TwCab3EBP0JavoLLu15oqWTV0blqYmpcXEJMNXufrVWYiGhylvCpM
Nh6IdsPukLDJ2MqRTDUtrdH/chzg0aHXubG3jF1NVlK+Nyr98kNMNbMZoTKMRxq7
Fk5L/28WJXWLZI+t5QTA5HpLoyRwdYY9S7M4WXfoe/jBJkcbsT9WVTNwCuqVxHVL
gLxP749xy3m2LX0kXVZEk/tjMFzPQ8eq2ttxOxOVJPBQIzSu8x3a7PDCZpjHEf6v
piGdTak2Wufsm6xcqCj6YvjpRGxHxtwfaJ9Ypd4TQL0pAIWNsfAyDDUat1Ru1k0O
4dGwOwRMJ6fhxbDbFPX7qlh0sa7aYi5n3feOICm7h3LOMy+kbUTRFwxyzpXcNhjM
r07HHVJdktsDPqlSKOqTll9rGTrZM8VCZNlXHFw/uVbNrzlTJmCu6NA9HZgBD3VH
Qg3BXK/iz3P8ePKu/ygxb4oArTxSr1b+Tty/+NwP50/wcgrFO9MK/ljxgyL32aoc
SZ/nwaHz6DNx2pGxqhqhE9GWE5Gi2Hkta5vGP1dXoztbtePnjqyorB+Lz3KIlcBy
jfytvosJsn3EPDdEs8ohZ+SUI47XSgi2aev/IyTy6gcNGUwWcAgmAusTbMA6m/KM
3gYtnCQUfVeZoVV4dZAqL8t1cbq8rVSjEgF2BUiTHp3JH2+Bqvs3KpM2BdVWx9NV
BtQRQ6jzOyPNotgDfzS92aJvGBZFPHpc8qmtjxoZKKT+6EjRVv+mERd9//usT9si
A5lPrDF+Nd7gS97iczCD/pE8OGDCJDDHHDSivkTfGPzpxctRvXMdMrZScSElxKPs
M9AfXwVd5ynG8gYjzUiER0QWAyCnNyIXc67/HFqc/yzmHgWNip8fcYXcqyddFrgE
s4ja3N2R2gvJUzNxXlEUqRh51SxUqWPYsj1zO3ZfX7EyXVxT9Bpg7eg2p3C1EcQz
OjrqVgttbdjNYjWnEDcZofL8sU9LsImzZDXb/4uQw/ZRddCLjIFI/5O8mAQMYNQF
S0convDzGzdk2MXT3goUPlW3l7mvkQ4iLxyrY56m/Fx89WJYwB95XFa4KJyLbM3b
ImjiQdokWtWQs4huE9Wvw7FHq0/UfDYk3uvnIYxTn4GruAoY0bHyLjruC8jEhRUY
hXioKyBJTsP5gcyFeCquSq5fNzomirAn2yOGv6oi4WFjDz+chxZ+IEkXZnYh4FUr
5Rrv9hXLcRi8WexOvsGVr6kzVfRYICObxHkNVe+p7qT4jJ1oDolFs3pdQJ2H2uun
hpOBDZhSvDpWEopZUoJCe4G63oPZZv1mODzUGyazsNstztCgqJdL3yhk65i9pMMr
uQQbdL77LrmlDiND4TR2klMR4O3wSUnWiIWSOUp2/3kj7cCu3PdRqseLn/uQnoQP
LpLEYG1/cb3EvxKzqMwsZWgRDRK9abwWT1UO5nE99G/39h0QdXwapOIxQ7kn+bGX
teSKo3EBAIShIdk84mpiFKvSKrkVHo8CwYC3xBEOf6inJ26TraLJ92lO0al+ZE/z
hscM7gsy5Z3gl3xd8meGPllf5DNs57G3IoN8+BYopbt+rPDUIDD3aJcoCDKa3FyO
B49GlDo8aKJt4rwtiThq8De49RiG2WOY5VDbBwW1tTTdTzM+zjJUv72F0wAaOL3A
MzWvHQd5qa/tFShptO2KhLzwpBl295/uflZ6Br7CxTQfS8bp5pJrHef7fNF7QnB7
y6yHiqDwVeOvxK0HVh8/Gwzj5sfa7NVBM1WtCrLBYQpVQ2hyGLQ3UV6ZOW1rfzWI
vyD/g9WS+xqWqMlr2j6sdcBvSb9fm7reZtpyhux3BXYYRFJUHJoozwEBmkR/9aip
w/y+dBf0gG7ezs6SKl1Pp9H+Rqylb5P++ntCv1wRJlVwOyax3h9DEkV8ZmkQYpTC
S24MioX4RMsEvHGinXKXW5OfxKm1Ts5jMctt5CoMn00Z2aBVdbCLS6KzLgpN0vvi
mqLb9WH+yeP1jJx+woMArGsFETfSmvKyZqYU8tu8EUAKDQbRds0D8tPC3gQqh7to
YyFXSNTTqIM+gtk8AONrytlTlvqTzTwpQBhDAfjrSPgU6GrRxTvE9/0uVSLtR6MR
8GMT0Kd7hOBqxtaroRSnO/o+nBmcO2oUPSvyAvIQXa4DL/nEYkTqIIg9nzL0xRSR
v5yDcioI5QxEmY3+LCfq6+HYtGf5eKPGoKBxJ+6Q+UvmX/1NhvSzoMpKJ8qxregG
CMSY1oO3QDGTZSeDp0McDFpheMcT4avFAyWspUFzyW5v4B3z4nLTZWCRngcrv2Lx
fMvRo7rxjGl1fwV58GZ31zLHBUXmc64QRcGa13G8i+0CDK7//u3l+OhVjn45i3oP
UjjhI9rqCpBLe16dEpjWJiwTbJ/3Gmy/kzrnzsVp8Nveo1T6yvU2BTWJefH4cm/S
CE963SsG+lL5TH2liSWvggKPdsLeH9tyxzl2KA0VrU/tCuoKeSLdNshyrFQU0gZp

--pragma protect end_data_block
--pragma protect digest_block
5Kk+7zbZRxkpihvj0NqI95I5ftk=
--pragma protect end_digest_block
--pragma protect end_protected
