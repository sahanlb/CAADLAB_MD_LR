-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
AbXIDb4OKNwnh/qiRai9hvQW3kRBn8bh9483rwt2BOAYsOYpMo8qiJomK+h7y5f2
mOPUo4OIzqMW3THhNJVoezpJ7xFEkFj3Ci1xeyTWV5Az01l1mROtNSwQszZKq/ZY
wT1oBad7p0YZ20JLF91NcSVqpa+Y1QCG4fwEwqBL/7tklltIbQH+9g==
--pragma protect end_key_block
--pragma protect digest_block
r3THakCLPEiwTZahRczQEp0c3AE=
--pragma protect end_digest_block
--pragma protect data_block
GSFtHP6Euy975mb7AWJS7iY7ZMvCzOBND+rZImehWmBuohvuAcOq5mR0J4oAPToo
tCVsMyAi2CVPZPk54/+bWc+wY7MQlas4SFyEQGFRR/y9agRpBm4g6dKWqxwzAS54
uM/bVgnyYiUVOMgi4yYEbnHv4tQX1ht8c8conptFnEgnhsqLpvINlXlPnQXF9KrW
mFh4n0Pv6FdaF17DyKTvHO9++Lvs8Go9bSC9UMHj8lsibj1D1lXcxYnZOLMcTmrr
X21SGZD6we/5AJXibevqVHI6g0OlW8OjjnmT/BX/2b3rfOu+ju/4N9bLqa5YNKya
SqDZ0n7iQU7BFJkaTA3w9SWCfe56zl6I2suzQc7u6ZOc0JKY6kUAWgZKlv+g/J+I
0v130Ay1bUCYFHkG9uuwVGLd1m+ApK5D5T4zo0N8y83EKJNIO7QQRuhthVIzjJ9E
bebz7/JoB+R8cXI6kglQ152gW+AavEtDJHL6weSFflvHo/UmEFMHXJEdrwef5cLP
fVJMiSVWq72rJo/aZH3wTRtSrhHArB0JayxUX/4FiHQeLnSSAg6fairAhTBw7NSo
zeW/WMNYslzqtf+tT87QMlEFy25vaIFDtjSezUHw3+Qroyc1Zs9I5pLH+fNUH8Wg
Qv8FTv4kOfZWalhMJl0dacM4qYbThMsyqIOqovFgf/97NykGd1Smgu8mQ729r2zG
3yI9NKecxawdql5nYfbOpvgqcniFgFdtzCZXGfOGbH+rWEaAGJH37TJCN/Aj4Qwg
VKy9L9D0EhpcQVXnRtLHDzh0osWs0V00k9zlTuFA6yRxnSFq2LghLODAYlBbgrur
HNmlGXtLKrVBrQD6LckdxTWLqPZR0rjpIu09VWPcIZaXt3sjWJQbk6EDsu/mnsvv
Lj8aET14lgDB5z1DUk/z/xdUBKEqqcz+vAYWqJCBtzz1wFv6uWDWXGufViXOdPH5
Wn60jlymFkmYwcGFk2M7oH9M4urFtPklj4ISBoZzyMfwF9JK+dmpZ8gnb5VV2GJi
PTYBrHkfaPOl3zQlLYPvcDgpU3j0bHoKtNhGuudnsJYsNNR0kUm/JIT394DK8cl5
jBW4fGbyBX3EHUhcpqWwjH1qWWD90/w1/7G5UVTPe9VRmfwFSMzAmxkc5T2FIur7
1VB7URqtGrHQJMTWkTPM5qF3SU7nnUwc1QhtcHU8g2szapd9bH+94Yx7kgXqm6cY
s/k2cCWktSLyYdHB9PCqGbdvRuKqMQD+ihlaR0UPDgya5qRSUfYrvGkhxWvW+4Zb
QgHvGdUBhGZf4ZjqXUxQyH1bkw3f0NxapyaycQZiQNd9G3bnfwsqhJy9qgkVQ0le
e+SwzUj9E5/0Ps9ZCMgtSGVFrbXXO73sCWRCllVAKFEiVvNQcSANLqKlH5uDTX4l
7yzsW0+B+PVOnsg499MYf33a2sdICzNQJMiWsqGPPavOhYLGVgJs38NpvoNgsfsn
NiaqyzKBq/O34f/zHTBmqCEWEhkbE3ezmj/VznopgCoamwuWjBJlvSBpnlNup9X7
cmMDCi+eDLx0O854Izi/27uQ7Gtu8+DsFmqTg6r+qQRzDnftza5zKkIvXbM7AA06
3TPa2qbbFF1dDYkeuqbzGeGBf3WAAzf8ZDozE0JFk7EXcSPbcrhoD3O4H8up5r0f
2aKmxV2YWup/zeJ41C8/AyCJYbca2lNg7dkp4H1G/sv+gGgvddy96JHxinujmfYf
eckkiXVerjTOvgKNk5edHDIXk9PD7twvfW+I9x8ep/K1jKWdKu3cAPlVd+661N4k
ldFP7E3DqMgCws57eMxysXSEHL83lWaiysXz5IZgXzdHd0okHGtgDyfiC1VJE0Ta
fEzsnq7nuU3NV17jsDomsmka/qV5UOSCPk+F7+gSPZHd1OS3NjnUyMYI69ecrxIM
Z1b3xBSeEXqRNSWEKHPPpvOgbOKCh1VFgQePSBUaRfKI/H98a7E/q2aYCICc8/Ov
c3m0excqoYSEZlmWlN3fX+M0iwkLPUxWEWA1aYfFPahvTGcrfWmj/bzSyfuCAg5G
JVCbTva6Oxli/m/OBia0e4Svk2lI9swwgRAZ01S4nb8sjMYUUYZXJkOeYDgeCEWm
DQ2DjzpKImbBADQxiOTZtjta9VWFRVtyKvIJSTouuC6vEpXsokLqSFs7rxo5j1EU
iaIQAPKR7uhwnfQjEUqhlgnGPsPQVLlBCGb8FPbLemul9KrQgYRbIZg1g/9KT/pk
sYuxnrKGFP4PCiqTZFCNJS1gI4SdDzv3TWaQYc/mfuAKj4bR/cbyHxyykzTaE0+f
vd53hu8auYhk/f5B2qtp/OrwthVnximaZfqhL+I1bjoCrf4nOGdfUEF+n8x9k8+r
Xkb+Coao2Gg2VJgRN8leLv93a+VKBthY33kpUypME/qYONcIMuWTHSExSTLShWNk
KLvOG0VPs8Vzj/qZpQCIfbcRGOnUM3i+K6ciqxPbhtf8sP8K8gGR+FJy9BVyxeqS
ojXld5aSA3mSSfLOyLhFNLgrIeeSApZxTKoXeP8G7EULsx23BaFHbrD3jllMZDcb
xlBGif+xFIEd9A/4SGFwBbXvzH5gKVBaI1yXUuKIStRks4gZ1LReDtkaaMPzAzBV
bt0QY4nUXz5Qnhl9GayPOZ9IxFhHJNDO+FN8/6zD4iUogpYVT/894DkrWPP3f2Fg
6/Zv0nxq7Q08Oyx8YsV2SeEq8QgSva8Qgic3Aqi/mk/4B685M4EnoumrNX5swgYW
XkS4caAUdVDT2uOGK5PZkeiQMEa4+ymEDUbIWcSSY9uNm3idJa91Et8xK3oX8vhA
sc2/1PQY7amsxt4NCAiMdlreDzBY9shVn+bcKiaW7HiX+iDxyt8pKyxe/D88FilA
gILJ1tVJTGgj1p59/y41Wm94l83rR0+E2/FmAxuCCe+qki2SGLCs/PJrTH3RZygf
NUcHqTHoq4Tojrhn/ADwQYHP9zuvLeEYB9FR9/N+Ta0ZDzRZagFf7EqEDMqqITdP
OPkFQTEOG2Acb+Ae73k0vDhPiQ/MPY0PlKnfS7I68Cql0voFzMEWTwB1i5s3Z8Gr
F5al1ihUqCwmnL0QDelYhX0EtiRThSmp+3eksHPzySKw204lh+H+i0wOi/fjEeHb
0l//0rKOID+G/be0V3OMthIxwTDYNMl7JZVZB8JlPg+4msyHCKZDijzNWJCNyA2e
rhrk+CRM9TjE4xkRa/t6/4ycFukaqJGBdGJ0i4YavqO+zFmLXIBCbyrJCYqajsQ9
V/AdFtuYr2MgNj3KaNuj24arhLZaUM0wpJiA7yeiIq3o9C9uxmxcTx9S+fVQMwna
96+NSQY7kTkiKzCfDXtUQzDDJe9MEmyKiJFDr42khpZ4bZ7Y0tH37McAtnIvsbYr
1w5On529iwwdMhAWPNj3BI/cAzH7sk/zqJbpLnqHQ+hOeVzYlMxsjCR9f2653OZV
fv5nVtI5Oqb6pMdrXfuzYDv6BPLMxt1H/Fqt9k0GfTrOl2LlxKEwQ8L0Enc1w0JS
yqXh5QDj5Fns/uaUH2GJZWmNWl7aGLlv2iQe6kVaotK3gUmEM4Fp6KQplZxGV8oO
ZbjMKI+DAloeeRdS9r63ZKqST/bTb4ycAjsRO6NsONNsRHZuFENm3K3SIlxpCjfq
9gbTEprwXJq4W7QQiSCpN2UD5F3n60TwGFGyHZm+U+qgM28g1kBLofBXuii1p2xl
xkN7rHSBMZVFNqHpDz6PKlbLV0ixMlV3uDZdnW4v6PZvgFUnRX4QReFddklg8Anh
m3LvTYVGilNVjJDdPOiPJfYpV9ejem1FVgu26S2/3POFtAWpKU3DsMx4b31OSA5v
Zul/+8u8eVzIHIUZLli6cWOlae+gMQKo+Mn4qnPw/g8mFwYlOk9hAal5sMRwz0wi
JRz13YyjjS17NnadLqdtGSr+SMz3nb2wZCQhbPmmVQcH1sIOM/sz/qEo3pgSNw3Y
/2N9Snl9zP75TpPww12hKylVMPwnMNonfqy5EvAc6c0uaT5V9pJDze/tyjSBNSP+
xzKk1LzaIVxtZVU+8nCXQlkIA2zmt5LdQSGVHhhIHzCDWN5hYiZ8CbFie5zBKmvT
jrFjk1BXSdR0lCxIShXZVmgY26+xLyZFklUqO/iDhvPaK7S6sccIUwgmxNquKcoQ
SITHERiqfTStNRRbmGB/L4VLszJuZTioxe9ecrXHQ8pMBTUHu4KdzhlNR0/jlfNk
tQi975vUzzzbt7boRY1OI2IBE7Z0C0RwhM13rJh31AFVpB4Gg2YrrGQvOijBzPkx
J9PixRZnMp5lj8ph1hPbWgqcF5ryWxcdDsPVgLV6HSPN+cI+elgH7WZEzDg6ETvz
KlFf6hEFQlboEwjtqTHriBcxdmzcE/FMY9VuuSagNSd9eCDhxuJBW45DjTdk97Jc
q2cAjwcCC7zha3iKU5z6XFbjBp3wFZFO7G15V6GQd4imJxdNpycroVPo/oVuRppY
OC4G2eRaJpeJQe3BDLSyn3/E0JDiqxRsBHPoTJI97Wjmcnu5f5EMAlMzzLVMZdIK
IQpi8O735Yk4IQr1WVAqM1rMDQE+y8mdJEcH+VFOXoY2NCXNn+h/GPXVZVpub16e
9twajCfpQJccbfod27DBhvR/Tbrs2o4Oa56AckGNGGvwdvPS8xNRUkeU9qDxau7u
1fsLr6qSzPkU98SWBXuAVJpAVXgB3PGwn1yszPoQ97J4tTrmV4dNX91tGM3Z0cOk
nTCVxRA/kj5FWQHBhh/jwTatUjY3ck6C4QjuQFgk51MMoiljV+F/4daQ88uRejAE
4SYM0Tlkq33MGmtGkeKltp7YDImgtiWYiBe25mzml/A/s4vKh7lJ3FngZG0o+fOF
3XW7oATJRLWw6g8xkQH/HSsqWREev3tKZrM0Fb+B1F9zu+aQEahVqtPAkik8ldCy
VTmcJh00QQ8nVi2r5yff7QsX4pI7UYmRmSddVqMT1uzN8A83pRGnOikctKUIdU2I
+5BwwsR0VgHlqT0vb2Arx+1HPEgiBTqkJIcOHVxb/LwK9RxmJrR0waFgpTzNkMn/
U7yUmKULXaYkFuNqYSoOG3FEnIxanpLdQJ/yFQiRbmH0erMgDT7Xf2ll+MsX0bGc
d6N10Smn6c1UCWA8KBqEfIuyRmP+ts1NS097VjxJHejPutzBtlDIXRgHg932YhpC
OelZsDePQmMhNE/RSvFdqZ2gzMy1ZGASPeVpSlAHCKslb5BMUrk3001AJ0yJw5SL
04yV2ED+liJQ/gb/Qi+QFqlzCiutLqVbG2hVb68fne9+T346mb9vIDb7yXszja5f
UOFta09WZLdqlP7KqCOQmpF+qfeZ9oq0GhutGODSEzcPBo1t/Zk/b34HB8TcfYXB
d/DEnirHwgEDl6j3lkaDHNf4bRk7o9dvgBS1g1hqDTlPHoMfLkOCKHl5Vo8tBqUR
JGfMweziX/y7UE2DvZNf2MHlUIBjLM0S5JL22uJVcsTMz/jDYGuayUGi/SCQndqp
Z3NDM40Ze13uU1v03P0QEXb4cDT7l3kK3YnCObsYCLp5zaOBdVqChw9wjN9vM4fP
Edvqo5YWnXfaPKtmxNevgVIs3wWerJiR05RWjMGrQfnMKEhQPcwQP4qfU8znUA3S
/Tww4mobctr0rRq6N8xDePaQmTSbnVaJ9kztyqoRwRVxHD4XAta+6GgixeBmDTbz
GTEVMLebDp3u5rxhJjGmTDnHTIOiff3uUKHCSeksrtbo8EmML6vtf1iZwwZsq2bE
UH71VhAMzu2d6d7UK9ABRQVClzb0NhmtWNbNXAw0BfDA1QBPeVa/6H/jUgRLan+w
LRGBGFa8GRFF6lH5k88VNlUeMyGMQ908H/J6yP9l9bGM/foWoB8pQ1+T+aE+4o/i
Hi8bR51hE7JPINEkf5bYMf3TMnlP4rP9jW7K8z8aXUxthVBxntEC25MgBef1RTjN
RW+o8cMeDFtxoe/TU986YDh1MwySh9vK5XpK6TZGGDbmHB/9Ba6uNTA2RBUEkpUl
/UYoDjrkbLJm8inCTUjvOGluIfrIXxEsrvDsgtMr62xxtWDoiqTV6lQtq1p41Bx7
J5F6hVEGgAVz/0MuJFK+zPArLCulR2+Pc839P5CS86EuOpD1iUq2SCMfykQK2jVx
THdgIRVFKZn6o3+hRHxJ6VjRZIQYTiDCZN69OcOPL5o+uQQWHPKXR9QKT7AMemqy
dg4tCWLAOzOtZimkB4tf+54+3HfIDTFNxoTJgpqJ7Rc+bCSaKVxH5x/+gWouLAJ6
7kBlJfIY6Rkohq7Gm3fOUZXzZ7XPN4hlnFHz6yMsw8iLO9uCERiGuIV0Vx3R44Uo
28biKPiUacDPllAWfCtDDWrKlRtxA++D2gLzGhejUYJmyeqnY2JfzGfXOZMC3tun
w6NKczHTHdvk1UUP8LH7fpKJeAsmZQbp/LtHWqwe0ppnaHB5CuzGeo0A1mhg0oOv
ugW63sxoxdlz/90iMXJl3ooNntFO3QC202ckl6Zj0iMemtfED8nT8EO7aig6nWEI
NnEaSwYcpMWrUBGXwIUI+QBi3eA+KY2XiTcn2fx1sz+GS7WrUlO81uCQC0IDypoq
YI5+M/hGQFK0Qrv49FUvEoUznd6FgOlZWigKrHs0jFxWsT5X8Kq3qW/fcAH34AVr
Nag4dyecFAqIA3M1t0u1BEqeBvnC+oQdK25Y+pGXaJsZ2QYf3TlqHEk3+a5tPg7o
pyuVqQCJ5p24O4gY5f82fjhU6JBronOgA7Pwk4uVUqUhJrOPXmgbVfytGDP9skvJ
/n3SmGkm6mJblv+LqwRBQyaBcjHGCmlDY1CIeV1QeLFkiwXerZQyLaOgJVcm90Md
yTthv7mfQBnXxC8Mrb1FUu6MCH/S6lV629dfr+/V9yqMi16rX2Mj4T7l4mvJVUz4
RnzTGuwtmkfwMORDfMr8VgAq5pFQuSTMvZhcI36+g9GHTE6pvbTnKEqR4gSoA37f
7Os60zEH3+0Gu+G/NWVTC6JiwbyUBQ5hoPKoYima/UJO1wtEGjLHPS9Qvn1HaQIx
ug+fujO9jd7nmwBfpDperKSQkZz85cl6YiW0JDqrcHFbPCR83UtB4rzRNuNSPUBs
7/Ujetm23jTPgkX6usvLwn1tXNWkEjZZKfZqk4fq38SjHR9h9ak4b4nplqloesq+
iHBisJCfrVcC27EYcvZidZThcCQ7wNhqHGbNqL9t6hnsVJu2/g5gOqlO3NwQu3qI
acG0VZjJHh2VnICK9DnIJQk4D0y/7Ii+nW80FKEfdHYcpGh52058CBxmQXmQKaV0
0ZX1nUP4YCjwZk6IyVPP31fkcwp2tgK5i4kW3DROpHX95jqINQ1GX9eHtjZzQZGL
AOzPeGZ3JR8PgN8MRzxLRf2XLyOKGw43yTOp8TO9hDc87UJQWgWMn6DYPlfJrag5
PZ9HLWVCXv1MSPhhOeGalUMEjGC+9rt+Kaifi1DcsRsSg5w6x+F8SYkCuX/xSybG
hVku3neCbUadjChZmZdBf8/Zqp7DhZ9XtZjNzdX2eei1iI8JHmCMmH7KlPzxfmg3
jppxKRN+XjcZCaR4UEdS5Niv9h4tLHjRIZJebGuANByacFTWO3uUBuTTRs9NLKzC
tw5qpa//fbf1taCgWnX2N3pkAoMi50tdBYgFoY47pMTOr1HfEhTsxht02g8Who8F
I/Ao8842Kb6iH0U65IUh8C5dp+audc5PY9QBdNMvfPE+O+PDfCijAJ7JI3o6t6h7
t9390UQTna91ZqASrBYlE2gpqTdtpYlf3J3CXSb/MfIgCbzncAi2REyZ/ySN0fOT
ol7Q+P1GJhoC20U9rUOQIP1fTwYlnIixfgot44eUIRMEb/qjwTjn9/c18BchzRaf
+VL0bjUqswnlpxzhMBR0toyLkFL1Hi6Evi/MIo9TZ4J4yZMgMSoFoTL9UANYgrp7
WMYOJqhimsuN0CxdXq7hVR2NFE2j5w8OQ8aRf8E5TUq12RbjmT1Flu76UEOcRW32
RkDFthFd1Fj2HGm0YP+Xx+R1m993LDNVdmeI8CEOW2SY8lg7ePEaypM+rEXRiW7v
a0BLeKnHzda8eHdNkSr1sS+yPU1YFLXiIEPjFOMQ7iZ3RkNdskdiIJ9B2JT8ZQpD
5x6nzd+U0QbFXv+0rdKUczuBkbA8XcdXbzsb/wnCMLDYA7dzLycJuoVwHqMhi/A7
zFuTpNtHOaeuk6+qHoCjRx7vzEwSlzNJ8aprH6mObriI3kYYj704zrprBpM2tEUR
FEbHc5iTei8WuI5vd9o8przUU00673HqKi+KP/qYbQ4mQapySWEhZlkpEzxW+g5T
K9r4CNUZo/R1AxJvJhd98ePr986o03JA0lJOoea/cHycQueu4qbEQCkj8FNrpSYQ
C6wNT7AnSUhoSShwBW1tcBgkskTGof+xal3xygIkjKYDSEeasWKjAl1BE1/BKqmH
WxvKY44ZEa/vljGM/KFB/d9kMcLMVG4AYwag3aPT/v1D1lNjtjSaG9wI8ldxX6lh
MtvOSHKzdAhqxcruhLVJwi4rOrHm4+44BJ+fy1gkyEB7LSL6IU7cIoWceoRgu7Z3
E4brw/0UZQycXhRg9EYI/WfIpVY01xnGD9d/dJx0PSZ36IWa/MMrvQUnbdQcrVhq
hnz0huVXCHFg/r+EssC9lN0n1N6PjeDQUZxnYMtCy0OBmjaT2u6jfAW6cVg30jjP
HTW1AibGM0WuNzrZBJWQEyHoiitOGYwvMz8ZsMVc/acAzQTAOjfx1/AesDfWV7C0
DePO0XGQBzAbScdyiC5/o8eMEfaETpMhwB5n0qvROzY2ruKLbmR+inaYSRIGKiD7
VMnh/O/nEnsBNkP+E7mF2GUPoUeaaNttqSLniLqoL8ezZFiI9ZhvhtrvPN+QOmhs
yU8Ima1yjWrGJ5gb+nOM2EzBTtFsefw0C67x6kjLsbotZJ1DInXa/ltB7AoHbq+n
baEKjAHziMgYBVh+P69kjajiOmGVPvXtyvdJ9LfwkrnXNdtcnqbyrcB3W3gOth/d
2AGEoSHDO63jzpcRiVe6PtaFVqeSZXTCo+Ud7U4NbTCBJd3BoDe8bi6lcAZ978mi
GoY5n6gn5lTmgtkGjAIOikJKig4VmEVzWmFC6D3yU6AqjH5UMSGHJsLQNN9+arW4
VQV1b8FlHvedJGpMTRH+7NzzP2SXuffjtUwTQKplSkLOq2tkqAUbzCxcDWJbY/ur
5quKHbfHyOZfbvuHO3hbOZzgTC0+YM7w7KtebcCBESZITsP+VmNDRcIQ8dFwXllM
l39p0jin44vtPLd2KCus6pT6nIwZ8pEL3/mKsaWzzB1Tt2TWg5kz93VUCvvwM6oQ
tl8bIIi29hToYIhkaYPQ1MyIyNidUv15tE5olgrv3isBN+GWqgkPsdp2pAU8UIm2
Qsh1b7YV5VylwA+6DuqOYA==
--pragma protect end_data_block
--pragma protect digest_block
ZdabI3jkach7x9Gl2TdU+d+AtOA=
--pragma protect end_digest_block
--pragma protect end_protected
