localparam [0:34428][128:0] P_INFO_NEW = {
  1'd1,  5'd1, 27'h0000031f, 5'd4, 27'h00000174, 5'd0, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c8, 5'd0, 27'h000000de, 5'd12, 27'h000002a9, 32'h00000400,
  1'd1,  5'd4, 27'h00000121, 5'd3, 27'h000001e9, 5'd24, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000378, 5'd11, 27'h000003f2, 5'd1, 27'h00000374, 32'h00000400,
  1'd1,  5'd4, 27'h0000023c, 5'd11, 27'h0000035c, 5'd11, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b6, 5'd14, 27'h00000328, 5'd22, 27'h0000025d, 32'h00000400,
  1'd1,  5'd3, 27'h000000c5, 5'd23, 27'h00000381, 5'd1, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001d2, 5'd23, 27'h000000b8, 5'd10, 27'h00000247, 32'h00000400,
  1'd1,  5'd0, 27'h000001b5, 5'd25, 27'h0000014f, 5'd24, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001df, 5'd0, 27'h0000007b, 5'd3, 27'h000003cd, 32'h00000400,
  1'd1,  5'd10, 27'h000003a7, 5'd0, 27'h000001e6, 5'd13, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000004d, 5'd0, 27'h000003e7, 5'd24, 27'h000003ec, 32'h00000400,
  1'd1,  5'd15, 27'h00000129, 5'd11, 27'h00000142, 5'd2, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000368, 5'd15, 27'h000000c4, 5'd14, 27'h00000071, 32'h00000400,
  1'd1,  5'd11, 27'h000003e9, 5'd11, 27'h000000ad, 5'd22, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001ba, 5'd24, 27'h00000075, 5'd0, 27'h0000005d, 32'h00000400,
  1'd1,  5'd14, 27'h0000017b, 5'd21, 27'h000003cd, 5'd15, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001cc, 5'd24, 27'h000001fb, 5'd23, 27'h000003bb, 32'h00000400,
  1'd1,  5'd24, 27'h00000359, 5'd4, 27'h000000b5, 5'd1, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e0, 5'd2, 27'h00000149, 5'd14, 27'h0000014b, 32'h00000400,
  1'd1,  5'd25, 27'h000002fa, 5'd4, 27'h00000071, 5'd23, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ee, 5'd12, 27'h0000037c, 5'd1, 27'h0000014b, 32'h00000400,
  1'd1,  5'd22, 27'h00000236, 5'd14, 27'h0000039d, 5'd13, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b2, 5'd10, 27'h000003e8, 5'd23, 27'h000003ad, 32'h00000400,
  1'd1,  5'd25, 27'h000001ae, 5'd24, 27'h000003dd, 5'd0, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000133, 5'd23, 27'h000001b0, 5'd12, 27'h00000231, 32'h00000400,
  1'd1,  5'd23, 27'h00000301, 5'd25, 27'h000002b4, 5'd21, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000093, 5'd4, 27'h000001d8, 5'd9, 27'h00000001, 32'h00000400,
  1'd1,  5'd0, 27'h00000199, 5'd0, 27'h000000c7, 5'd19, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a4, 5'd2, 27'h000001e2, 5'd30, 27'h0000038e, 32'h00000400,
  1'd1,  5'd3, 27'h00000376, 5'd13, 27'h000003d7, 5'd7, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000037, 5'd12, 27'h0000020d, 5'd16, 27'h00000132, 32'h00000400,
  1'd1,  5'd1, 27'h000002b8, 5'd12, 27'h000000d0, 5'd28, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f1, 5'd24, 27'h0000025e, 5'd5, 27'h00000290, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd23, 27'h00000377, 5'd16, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026f, 5'd20, 27'h000002fc, 5'd29, 27'h00000226, 32'h00000400,
  1'd1,  5'd12, 27'h0000027c, 5'd2, 27'h00000390, 5'd8, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000294, 5'd2, 27'h000001e3, 5'd15, 27'h00000368, 32'h00000400,
  1'd1,  5'd10, 27'h00000362, 5'd3, 27'h0000009f, 5'd27, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000276, 5'd10, 27'h00000229, 5'd10, 27'h00000110, 32'h00000400,
  1'd1,  5'd13, 27'h0000036e, 5'd11, 27'h0000014d, 5'd18, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000fa, 5'd14, 27'h000002ab, 5'd30, 27'h00000100, 32'h00000400,
  1'd1,  5'd14, 27'h0000019d, 5'd22, 27'h00000118, 5'd5, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000212, 5'd25, 27'h000002ea, 5'd16, 27'h0000025d, 32'h00000400,
  1'd1,  5'd11, 27'h0000031d, 5'd20, 27'h00000392, 5'd27, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000106, 5'd1, 27'h0000024d, 5'd6, 27'h00000077, 32'h00000400,
  1'd1,  5'd21, 27'h00000014, 5'd0, 27'h000001ae, 5'd16, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000132, 5'd4, 27'h0000019e, 5'd30, 27'h000000bf, 32'h00000400,
  1'd1,  5'd24, 27'h00000054, 5'd12, 27'h000001b9, 5'd8, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000008c, 5'd11, 27'h00000022, 5'd17, 27'h000000b4, 32'h00000400,
  1'd1,  5'd22, 27'h00000074, 5'd13, 27'h00000390, 5'd29, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d3, 5'd24, 27'h00000354, 5'd9, 27'h00000018, 32'h00000400,
  1'd1,  5'd21, 27'h00000259, 5'd22, 27'h00000311, 5'd18, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000f7, 5'd21, 27'h00000149, 5'd29, 27'h0000038e, 32'h00000400,
  1'd1,  5'd4, 27'h0000025a, 5'd6, 27'h000003de, 5'd4, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000171, 5'd6, 27'h0000039f, 5'd11, 27'h00000071, 32'h00000400,
  1'd1,  5'd3, 27'h000002f3, 5'd6, 27'h000003c2, 5'd23, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fe, 5'd18, 27'h00000209, 5'd4, 27'h00000112, 32'h00000400,
  1'd1,  5'd3, 27'h00000192, 5'd20, 27'h00000089, 5'd11, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c4, 5'd18, 27'h000003e0, 5'd23, 27'h0000000c, 32'h00000400,
  1'd1,  5'd2, 27'h0000027e, 5'd28, 27'h00000108, 5'd2, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000283, 5'd30, 27'h000003df, 5'd13, 27'h000001a2, 32'h00000400,
  1'd1,  5'd3, 27'h000000d3, 5'd30, 27'h0000029b, 5'd25, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000271, 5'd5, 27'h000000f0, 5'd2, 27'h00000174, 32'h00000400,
  1'd1,  5'd14, 27'h000003fe, 5'd6, 27'h00000100, 5'd11, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000255, 5'd8, 27'h000001ca, 5'd23, 27'h00000087, 32'h00000400,
  1'd1,  5'd11, 27'h0000020e, 5'd18, 27'h00000379, 5'd3, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000be, 5'd20, 27'h000000b1, 5'd12, 27'h00000029, 32'h00000400,
  1'd1,  5'd13, 27'h0000009e, 5'd17, 27'h0000020d, 5'd23, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000376, 5'd26, 27'h0000005c, 5'd0, 27'h00000080, 32'h00000400,
  1'd1,  5'd14, 27'h0000023e, 5'd29, 27'h000003e5, 5'd10, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000035a, 5'd26, 27'h0000002e, 5'd21, 27'h00000166, 32'h00000400,
  1'd1,  5'd22, 27'h00000323, 5'd7, 27'h0000022c, 5'd2, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000024e, 5'd9, 27'h00000104, 5'd14, 27'h00000019, 32'h00000400,
  1'd1,  5'd20, 27'h0000031b, 5'd9, 27'h000002e9, 5'd22, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000024b, 5'd20, 27'h00000097, 5'd0, 27'h000002f1, 32'h00000400,
  1'd1,  5'd23, 27'h0000007c, 5'd16, 27'h000003c7, 5'd13, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ef, 5'd18, 27'h000003bb, 5'd25, 27'h0000017a, 32'h00000400,
  1'd1,  5'd25, 27'h000001e1, 5'd30, 27'h000001d9, 5'd2, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000339, 5'd30, 27'h0000010f, 5'd14, 27'h0000018c, 32'h00000400,
  1'd1,  5'd20, 27'h0000031b, 5'd27, 27'h00000121, 5'd21, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c5, 5'd5, 27'h00000263, 5'd7, 27'h0000004f, 32'h00000400,
  1'd1,  5'd2, 27'h00000148, 5'd8, 27'h000003b4, 5'd16, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000012f, 5'd5, 27'h0000038d, 5'd28, 27'h000000e1, 32'h00000400,
  1'd1,  5'd0, 27'h000001b1, 5'd17, 27'h0000030e, 5'd8, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000038e, 5'd18, 27'h00000261, 5'd16, 27'h00000244, 32'h00000400,
  1'd1,  5'd3, 27'h00000388, 5'd19, 27'h0000022d, 5'd27, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fe, 5'd27, 27'h000000c6, 5'd6, 27'h0000023e, 32'h00000400,
  1'd1,  5'd4, 27'h000000e8, 5'd27, 27'h00000362, 5'd15, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000304, 5'd28, 27'h000001bd, 5'd28, 27'h0000004d, 32'h00000400,
  1'd1,  5'd11, 27'h000000d7, 5'd8, 27'h00000342, 5'd9, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000142, 5'd9, 27'h00000234, 5'd19, 27'h0000002e, 32'h00000400,
  1'd1,  5'd13, 27'h000003a9, 5'd7, 27'h000003eb, 5'd29, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000089, 5'd18, 27'h0000009d, 5'd9, 27'h00000132, 32'h00000400,
  1'd1,  5'd13, 27'h000002d8, 5'd16, 27'h0000034b, 5'd15, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000054, 5'd18, 27'h00000156, 5'd26, 27'h0000036a, 32'h00000400,
  1'd1,  5'd14, 27'h0000028f, 5'd26, 27'h00000182, 5'd8, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000089, 5'd26, 27'h00000020, 5'd19, 27'h000002c6, 32'h00000400,
  1'd1,  5'd12, 27'h000001d7, 5'd28, 27'h000003fe, 5'd29, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e3, 5'd8, 27'h000003d2, 5'd5, 27'h0000021c, 32'h00000400,
  1'd1,  5'd22, 27'h000002bb, 5'd9, 27'h00000337, 5'd19, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031e, 5'd8, 27'h00000237, 5'd30, 27'h0000019d, 32'h00000400,
  1'd1,  5'd22, 27'h0000007f, 5'd18, 27'h00000380, 5'd9, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002a8, 5'd16, 27'h000000cc, 5'd19, 27'h000002bd, 32'h00000400,
  1'd1,  5'd23, 27'h00000148, 5'd17, 27'h0000025c, 5'd28, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000005b, 5'd28, 27'h00000230, 5'd8, 27'h00000181, 32'h00000400,
  1'd1,  5'd23, 27'h00000183, 5'd27, 27'h000001b2, 5'd16, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000382, 5'd26, 27'h00000259, 5'd26, 27'h000001ca, 32'h00000400,
  1'd1,  5'd6, 27'h000001e5, 5'd0, 27'h00000149, 5'd8, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002de, 5'd2, 27'h00000083, 5'd19, 27'h000000c2, 32'h00000400,
  1'd1,  5'd6, 27'h000001ff, 5'd0, 27'h00000232, 5'd26, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000019, 5'd12, 27'h0000015e, 5'd2, 27'h0000036a, 32'h00000400,
  1'd1,  5'd6, 27'h00000090, 5'd11, 27'h00000289, 5'd10, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a2, 5'd12, 27'h000000d2, 5'd23, 27'h000002b5, 32'h00000400,
  1'd1,  5'd7, 27'h00000070, 5'd24, 27'h000000f2, 5'd2, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000004e, 5'd22, 27'h000000b1, 5'd11, 27'h00000200, 32'h00000400,
  1'd1,  5'd5, 27'h000002e6, 5'd21, 27'h000002e7, 5'd24, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000267, 5'd0, 27'h000000da, 5'd5, 27'h000002b9, 32'h00000400,
  1'd1,  5'd18, 27'h00000266, 5'd1, 27'h00000149, 5'd18, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000169, 5'd3, 27'h000001de, 5'd26, 27'h0000027d, 32'h00000400,
  1'd1,  5'd16, 27'h00000204, 5'd12, 27'h000003ec, 5'd0, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002e2, 5'd10, 27'h0000033e, 5'd15, 27'h00000088, 32'h00000400,
  1'd1,  5'd15, 27'h0000020a, 5'd11, 27'h000003c8, 5'd23, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003a2, 5'd20, 27'h000003f5, 5'd1, 27'h00000328, 32'h00000400,
  1'd1,  5'd16, 27'h000000b9, 5'd22, 27'h00000203, 5'd11, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000026f, 5'd25, 27'h000000e1, 5'd24, 27'h0000011b, 32'h00000400,
  1'd1,  5'd29, 27'h000002ea, 5'd4, 27'h000003b0, 5'd0, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000257, 5'd0, 27'h00000191, 5'd14, 27'h000001ea, 32'h00000400,
  1'd1,  5'd30, 27'h000000e2, 5'd1, 27'h000002d8, 5'd21, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ae, 5'd11, 27'h000001c3, 5'd2, 27'h00000010, 32'h00000400,
  1'd1,  5'd30, 27'h000003e6, 5'd11, 27'h000000f7, 5'd10, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000019, 5'd13, 27'h00000211, 5'd22, 27'h000002b8, 32'h00000400,
  1'd1,  5'd27, 27'h000001bd, 5'd22, 27'h0000038a, 5'd3, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001e8, 5'd20, 27'h000002c6, 5'd10, 27'h00000398, 32'h00000400,
  1'd1,  5'd28, 27'h000000c1, 5'd22, 27'h0000023b, 5'd24, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000113, 5'd4, 27'h000001c9, 5'd3, 27'h000002a9, 32'h00000400,
  1'd1,  5'd7, 27'h0000002c, 5'd3, 27'h00000006, 5'd15, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000349, 5'd3, 27'h0000011b, 5'd21, 27'h00000097, 32'h00000400,
  1'd1,  5'd5, 27'h0000036d, 5'd13, 27'h000000ee, 5'd7, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000353, 5'd11, 27'h0000028b, 5'd18, 27'h00000025, 32'h00000400,
  1'd1,  5'd9, 27'h00000040, 5'd13, 27'h000000c8, 5'd27, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000227, 5'd21, 27'h00000020, 5'd5, 27'h000000f6, 32'h00000400,
  1'd1,  5'd7, 27'h00000185, 5'd25, 27'h000001af, 5'd17, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000386, 5'd23, 27'h00000327, 5'd28, 27'h000001c2, 32'h00000400,
  1'd1,  5'd16, 27'h00000255, 5'd4, 27'h00000037, 5'd1, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f8, 5'd2, 27'h000000e3, 5'd14, 27'h000001f4, 32'h00000400,
  1'd1,  5'd19, 27'h00000282, 5'd1, 27'h00000134, 5'd23, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000375, 5'd14, 27'h000003f0, 5'd9, 27'h00000009, 32'h00000400,
  1'd1,  5'd17, 27'h00000228, 5'd11, 27'h00000282, 5'd18, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f9, 5'd12, 27'h000001ab, 5'd26, 27'h00000240, 32'h00000400,
  1'd1,  5'd16, 27'h0000025d, 5'd24, 27'h000003cc, 5'd9, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000016, 5'd24, 27'h00000057, 5'd16, 27'h00000369, 32'h00000400,
  1'd1,  5'd20, 27'h00000186, 5'd23, 27'h000002e8, 5'd30, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000349, 5'd0, 27'h0000024a, 5'd5, 27'h0000036b, 32'h00000400,
  1'd1,  5'd29, 27'h00000009, 5'd3, 27'h000002a4, 5'd19, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001d, 5'd4, 27'h00000332, 5'd29, 27'h0000018c, 32'h00000400,
  1'd1,  5'd25, 27'h00000382, 5'd13, 27'h00000389, 5'd6, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001ee, 5'd13, 27'h000001c3, 5'd15, 27'h0000035a, 32'h00000400,
  1'd1,  5'd26, 27'h000000b4, 5'd15, 27'h00000043, 5'd26, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c0, 5'd21, 27'h0000001e, 5'd7, 27'h00000250, 32'h00000400,
  1'd1,  5'd28, 27'h000001cf, 5'd25, 27'h0000016c, 5'd20, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003c7, 5'd22, 27'h0000016d, 5'd28, 27'h00000078, 32'h00000400,
  1'd1,  5'd9, 27'h000000a5, 5'd8, 27'h0000028f, 5'd0, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000326, 5'd6, 27'h000003bb, 5'd10, 27'h000001ca, 32'h00000400,
  1'd1,  5'd9, 27'h00000346, 5'd6, 27'h00000222, 5'd22, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003f8, 5'd16, 27'h000002ba, 5'd4, 27'h00000341, 32'h00000400,
  1'd1,  5'd10, 27'h0000010a, 5'd17, 27'h00000031, 5'd14, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000273, 5'd19, 27'h00000286, 5'd20, 27'h000002fe, 32'h00000400,
  1'd1,  5'd6, 27'h00000316, 5'd28, 27'h00000238, 5'd2, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000185, 5'd30, 27'h00000163, 5'd11, 27'h0000028c, 32'h00000400,
  1'd1,  5'd9, 27'h000002b3, 5'd28, 27'h00000141, 5'd24, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000214, 5'd5, 27'h0000019f, 5'd2, 27'h000000a8, 32'h00000400,
  1'd1,  5'd16, 27'h000003d3, 5'd8, 27'h0000010c, 5'd11, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000397, 5'd7, 27'h000000a6, 5'd20, 27'h00000349, 32'h00000400,
  1'd1,  5'd18, 27'h0000036b, 5'd16, 27'h00000372, 5'd4, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000036b, 5'd19, 27'h00000239, 5'd14, 27'h00000334, 32'h00000400,
  1'd1,  5'd19, 27'h000003d9, 5'd19, 27'h000002cc, 5'd22, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000160, 5'd25, 27'h0000037f, 5'd2, 27'h00000202, 32'h00000400,
  1'd1,  5'd19, 27'h000003e1, 5'd30, 27'h00000338, 5'd10, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e3, 5'd28, 27'h000003e5, 5'd22, 27'h00000176, 32'h00000400,
  1'd1,  5'd29, 27'h000001bd, 5'd6, 27'h0000007a, 5'd2, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003fe, 5'd8, 27'h000003ff, 5'd10, 27'h00000292, 32'h00000400,
  1'd1,  5'd28, 27'h00000158, 5'd7, 27'h000000c4, 5'd25, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000263, 5'd19, 27'h0000013d, 5'd2, 27'h0000013a, 32'h00000400,
  1'd1,  5'd26, 27'h0000007d, 5'd16, 27'h0000024f, 5'd13, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000191, 5'd17, 27'h00000263, 5'd25, 27'h00000213, 32'h00000400,
  1'd1,  5'd30, 27'h00000113, 5'd27, 27'h0000005c, 5'd5, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000134, 5'd28, 27'h00000033, 5'd11, 27'h0000003a, 32'h00000400,
  1'd1,  5'd26, 27'h000003e0, 5'd27, 27'h0000000f, 5'd25, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000219, 5'd7, 27'h0000026f, 5'd7, 27'h0000024b, 32'h00000400,
  1'd1,  5'd9, 27'h000001a9, 5'd8, 27'h0000015f, 5'd16, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ff, 5'd6, 27'h00000074, 5'd26, 27'h000002b0, 32'h00000400,
  1'd1,  5'd8, 27'h0000027e, 5'd17, 27'h0000020a, 5'd6, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012f, 5'd18, 27'h00000112, 5'd16, 27'h00000261, 32'h00000400,
  1'd1,  5'd6, 27'h0000000e, 5'd19, 27'h000003fe, 5'd26, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003bb, 5'd30, 27'h000000e6, 5'd8, 27'h000001d3, 32'h00000400,
  1'd1,  5'd7, 27'h00000091, 5'd27, 27'h000000a6, 5'd16, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003f6, 5'd26, 27'h00000133, 5'd28, 27'h000001e4, 32'h00000400,
  1'd1,  5'd18, 27'h00000239, 5'd7, 27'h000003c7, 5'd6, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000237, 5'd6, 27'h00000341, 5'd16, 27'h00000026, 32'h00000400,
  1'd1,  5'd20, 27'h000000d0, 5'd9, 27'h000000a5, 5'd27, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000007d, 5'd17, 27'h00000056, 5'd5, 27'h000003be, 32'h00000400,
  1'd1,  5'd17, 27'h00000296, 5'd17, 27'h0000019d, 5'd16, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000031f, 5'd15, 27'h0000024d, 5'd30, 27'h000001f7, 32'h00000400,
  1'd1,  5'd16, 27'h0000001f, 5'd30, 27'h000000ba, 5'd6, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000397, 5'd27, 27'h00000387, 5'd18, 27'h000003b8, 32'h00000400,
  1'd1,  5'd20, 27'h000001ec, 5'd28, 27'h00000388, 5'd30, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000347, 5'd7, 27'h00000183, 5'd8, 27'h000002e3, 32'h00000400,
  1'd1,  5'd26, 27'h000000be, 5'd8, 27'h00000023, 5'd18, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003bd, 5'd5, 27'h0000012b, 5'd30, 27'h000002db, 32'h00000400,
  1'd1,  5'd30, 27'h000000de, 5'd20, 27'h000001f8, 5'd6, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e9, 5'd16, 27'h000001f4, 5'd18, 27'h00000109, 32'h00000400,
  1'd1,  5'd29, 27'h00000318, 5'd18, 27'h000002e4, 5'd27, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a3, 5'd27, 27'h0000006c, 5'd7, 27'h000002ba, 32'h00000400,
  1'd1,  5'd30, 27'h000001cf, 5'd28, 27'h000000e1, 5'd15, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000385, 5'd26, 27'h0000039e, 5'd30, 27'h000003e5, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h0000031c, 5'd1, 27'h000003f8, 5'd2, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000029d, 5'd2, 27'h000002c2, 5'd13, 27'h00000089, 32'h00000400,
  1'd1,  5'd1, 27'h000001aa, 5'd1, 27'h0000006d, 5'd21, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000f3, 5'd13, 27'h0000006e, 5'd1, 27'h0000029b, 32'h00000400,
  1'd1,  5'd3, 27'h0000022a, 5'd14, 27'h00000011, 5'd13, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000254, 5'd14, 27'h0000000a, 5'd23, 27'h00000377, 32'h00000400,
  1'd1,  5'd5, 27'h00000008, 5'd22, 27'h0000015a, 5'd3, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002da, 5'd23, 27'h000003dd, 5'd11, 27'h000000d9, 32'h00000400,
  1'd1,  5'd3, 27'h00000092, 5'd21, 27'h0000010d, 5'd24, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000298, 5'd0, 27'h0000007c, 5'd2, 27'h0000001d, 32'h00000400,
  1'd1,  5'd14, 27'h000001db, 5'd2, 27'h0000020a, 5'd10, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b4, 5'd0, 27'h00000351, 5'd24, 27'h0000038d, 32'h00000400,
  1'd1,  5'd11, 27'h00000262, 5'd11, 27'h00000108, 5'd1, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001ba, 5'd14, 27'h000001cb, 5'd13, 27'h0000028b, 32'h00000400,
  1'd1,  5'd14, 27'h0000011f, 5'd12, 27'h000003be, 5'd24, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f4, 5'd23, 27'h0000035d, 5'd3, 27'h000001d3, 32'h00000400,
  1'd1,  5'd11, 27'h0000037f, 5'd24, 27'h000000d7, 5'd12, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000355, 5'd22, 27'h00000355, 5'd25, 27'h0000028d, 32'h00000400,
  1'd1,  5'd22, 27'h0000015e, 5'd3, 27'h00000273, 5'd2, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ba, 5'd3, 27'h000001d9, 5'd13, 27'h0000006d, 32'h00000400,
  1'd1,  5'd23, 27'h00000009, 5'd3, 27'h00000051, 5'd21, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000299, 5'd11, 27'h00000203, 5'd1, 27'h00000062, 32'h00000400,
  1'd1,  5'd23, 27'h000002dc, 5'd13, 27'h0000020c, 5'd12, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000375, 5'd14, 27'h00000109, 5'd21, 27'h000000c2, 32'h00000400,
  1'd1,  5'd21, 27'h00000166, 5'd22, 27'h00000092, 5'd4, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b3, 5'd22, 27'h00000036, 5'd13, 27'h000002c5, 32'h00000400,
  1'd1,  5'd23, 27'h000000f9, 5'd20, 27'h00000374, 5'd25, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000039a, 5'd4, 27'h00000262, 5'd9, 27'h0000014e, 32'h00000400,
  1'd1,  5'd1, 27'h00000248, 5'd0, 27'h000002ab, 5'd17, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b0, 5'd2, 27'h0000005c, 5'd26, 27'h000000e8, 32'h00000400,
  1'd1,  5'd1, 27'h000002b8, 5'd10, 27'h00000209, 5'd7, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000053, 5'd11, 27'h000003d2, 5'd17, 27'h0000030b, 32'h00000400,
  1'd1,  5'd2, 27'h0000007b, 5'd14, 27'h000002a4, 5'd26, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a8, 5'd21, 27'h000000bf, 5'd6, 27'h000001b9, 32'h00000400,
  1'd1,  5'd2, 27'h00000303, 5'd23, 27'h000003c5, 5'd20, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002f0, 5'd23, 27'h00000035, 5'd25, 27'h0000039f, 32'h00000400,
  1'd1,  5'd10, 27'h00000391, 5'd4, 27'h00000231, 5'd5, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000113, 5'd0, 27'h00000361, 5'd17, 27'h000001a4, 32'h00000400,
  1'd1,  5'd14, 27'h0000035f, 5'd4, 27'h0000001a, 5'd30, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fe, 5'd10, 27'h000002b8, 5'd6, 27'h00000325, 32'h00000400,
  1'd1,  5'd10, 27'h000003f6, 5'd14, 27'h000000aa, 5'd18, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000161, 5'd12, 27'h00000212, 5'd28, 27'h00000174, 32'h00000400,
  1'd1,  5'd12, 27'h000001e2, 5'd23, 27'h0000004e, 5'd10, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000022f, 5'd25, 27'h000002ad, 5'd20, 27'h00000085, 32'h00000400,
  1'd1,  5'd12, 27'h000000e7, 5'd21, 27'h000003b7, 5'd27, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000cb, 5'd4, 27'h00000254, 5'd9, 27'h00000066, 32'h00000400,
  1'd1,  5'd23, 27'h00000210, 5'd3, 27'h00000032, 5'd19, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a8, 5'd0, 27'h0000012f, 5'd29, 27'h000002f8, 32'h00000400,
  1'd1,  5'd23, 27'h00000033, 5'd14, 27'h00000400, 5'd6, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000006e, 5'd13, 27'h00000004, 5'd18, 27'h000001fa, 32'h00000400,
  1'd1,  5'd21, 27'h000002f2, 5'd13, 27'h00000346, 5'd29, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000372, 5'd24, 27'h00000331, 5'd5, 27'h00000280, 32'h00000400,
  1'd1,  5'd23, 27'h0000015e, 5'd23, 27'h0000004f, 5'd15, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000f9, 5'd20, 27'h000002d4, 5'd29, 27'h00000136, 32'h00000400,
  1'd1,  5'd3, 27'h0000024b, 5'd8, 27'h000002d5, 5'd2, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001cb, 5'd10, 27'h0000013b, 5'd11, 27'h00000253, 32'h00000400,
  1'd1,  5'd3, 27'h00000023, 5'd9, 27'h00000284, 5'd22, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000106, 5'd15, 27'h00000267, 5'd0, 27'h000003c7, 32'h00000400,
  1'd1,  5'd5, 27'h00000048, 5'd16, 27'h000003fc, 5'd10, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000025c, 5'd20, 27'h00000157, 5'd22, 27'h000000b7, 32'h00000400,
  1'd1,  5'd4, 27'h0000036f, 5'd28, 27'h0000032c, 5'd0, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000012f, 5'd26, 27'h00000164, 5'd14, 27'h000001fa, 32'h00000400,
  1'd1,  5'd4, 27'h000001e5, 5'd27, 27'h00000037, 5'd22, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e4, 5'd9, 27'h00000045, 5'd5, 27'h00000027, 32'h00000400,
  1'd1,  5'd11, 27'h000002ac, 5'd5, 27'h000001a5, 5'd12, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000141, 5'd6, 27'h000000f6, 5'd21, 27'h00000272, 32'h00000400,
  1'd1,  5'd13, 27'h0000014b, 5'd16, 27'h0000037e, 5'd2, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002e8, 5'd19, 27'h000000ea, 5'd11, 27'h0000019e, 32'h00000400,
  1'd1,  5'd10, 27'h0000032d, 5'd15, 27'h000003c6, 5'd25, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000083, 5'd27, 27'h000000f8, 5'd3, 27'h000003c8, 32'h00000400,
  1'd1,  5'd10, 27'h000001b0, 5'd25, 27'h00000370, 5'd11, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000147, 5'd26, 27'h000003d7, 5'd25, 27'h00000353, 32'h00000400,
  1'd1,  5'd25, 27'h00000120, 5'd7, 27'h00000311, 5'd2, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000397, 5'd9, 27'h00000226, 5'd12, 27'h00000314, 32'h00000400,
  1'd1,  5'd22, 27'h00000307, 5'd5, 27'h0000035c, 5'd24, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000029f, 5'd16, 27'h000002b8, 5'd1, 27'h000000f6, 32'h00000400,
  1'd1,  5'd22, 27'h00000225, 5'd20, 27'h00000189, 5'd12, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000335, 5'd19, 27'h00000019, 5'd20, 27'h000003e2, 32'h00000400,
  1'd1,  5'd25, 27'h0000006f, 5'd28, 27'h000002bf, 5'd4, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000322, 5'd30, 27'h000001cd, 5'd12, 27'h00000006, 32'h00000400,
  1'd1,  5'd25, 27'h000001a3, 5'd30, 27'h000002a2, 5'd25, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a6, 5'd7, 27'h00000121, 5'd5, 27'h00000326, 32'h00000400,
  1'd1,  5'd4, 27'h00000173, 5'd6, 27'h00000237, 5'd18, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000347, 5'd7, 27'h0000025f, 5'd26, 27'h00000110, 32'h00000400,
  1'd1,  5'd1, 27'h000001cd, 5'd17, 27'h0000014d, 5'd7, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a7, 5'd19, 27'h0000036a, 5'd18, 27'h000002b9, 32'h00000400,
  1'd1,  5'd2, 27'h000000fe, 5'd20, 27'h000000f7, 5'd28, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000014b, 5'd26, 27'h00000024, 5'd9, 27'h0000039e, 32'h00000400,
  1'd1,  5'd4, 27'h000000db, 5'd29, 27'h000001ac, 5'd18, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003e7, 5'd30, 27'h00000379, 5'd28, 27'h000000af, 32'h00000400,
  1'd1,  5'd15, 27'h00000060, 5'd7, 27'h00000103, 5'd5, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f3, 5'd8, 27'h00000013, 5'd19, 27'h00000228, 32'h00000400,
  1'd1,  5'd13, 27'h000003a9, 5'd8, 27'h00000166, 5'd29, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000062, 5'd16, 27'h00000354, 5'd9, 27'h000003c6, 32'h00000400,
  1'd1,  5'd10, 27'h000001f4, 5'd19, 27'h000000b1, 5'd20, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000284, 5'd19, 27'h00000304, 5'd28, 27'h00000004, 32'h00000400,
  1'd1,  5'd11, 27'h00000225, 5'd26, 27'h0000001a, 5'd5, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000160, 5'd29, 27'h00000012, 5'd18, 27'h00000031, 32'h00000400,
  1'd1,  5'd12, 27'h0000008e, 5'd28, 27'h0000014a, 5'd28, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001e3, 5'd10, 27'h000000b9, 5'd7, 27'h00000228, 32'h00000400,
  1'd1,  5'd22, 27'h0000019d, 5'd8, 27'h00000078, 5'd19, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003be, 5'd5, 27'h00000227, 5'd26, 27'h0000038f, 32'h00000400,
  1'd1,  5'd23, 27'h000001b5, 5'd19, 27'h0000033e, 5'd9, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f5, 5'd16, 27'h000000d7, 5'd17, 27'h000001f7, 32'h00000400,
  1'd1,  5'd25, 27'h00000128, 5'd20, 27'h000001b8, 5'd26, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000342, 5'd30, 27'h0000031f, 5'd9, 27'h0000001e, 32'h00000400,
  1'd1,  5'd23, 27'h000003eb, 5'd29, 27'h000001e4, 5'd18, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000377, 5'd29, 27'h00000103, 5'd29, 27'h0000032f, 32'h00000400,
  1'd1,  5'd7, 27'h000000a2, 5'd2, 27'h000003a2, 5'd6, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000005, 5'd3, 27'h00000202, 5'd16, 27'h00000188, 32'h00000400,
  1'd1,  5'd6, 27'h000001e4, 5'd2, 27'h000002b9, 5'd27, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000cc, 5'd10, 27'h00000185, 5'd0, 27'h00000135, 32'h00000400,
  1'd1,  5'd5, 27'h00000285, 5'd10, 27'h000001dc, 5'd15, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000259, 5'd14, 27'h00000367, 5'd20, 27'h00000399, 32'h00000400,
  1'd1,  5'd7, 27'h00000252, 5'd22, 27'h0000038c, 5'd3, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000049, 5'd21, 27'h00000362, 5'd11, 27'h00000018, 32'h00000400,
  1'd1,  5'd7, 27'h0000007b, 5'd21, 27'h0000026f, 5'd24, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001d7, 5'd4, 27'h0000030c, 5'd9, 27'h000002fe, 32'h00000400,
  1'd1,  5'd19, 27'h0000017e, 5'd2, 27'h000003ed, 5'd20, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d7, 5'd0, 27'h00000338, 5'd29, 27'h0000026a, 32'h00000400,
  1'd1,  5'd18, 27'h000003b6, 5'd13, 27'h000001e2, 5'd0, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000003c, 5'd11, 27'h0000014d, 5'd10, 27'h00000365, 32'h00000400,
  1'd1,  5'd16, 27'h0000002b, 5'd10, 27'h00000247, 5'd22, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000039, 5'd24, 27'h0000026b, 5'd0, 27'h0000021d, 32'h00000400,
  1'd1,  5'd20, 27'h00000116, 5'd24, 27'h00000213, 5'd11, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f2, 5'd23, 27'h00000231, 5'd22, 27'h000001dd, 32'h00000400,
  1'd1,  5'd29, 27'h0000014d, 5'd4, 27'h0000018d, 5'd2, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002bb, 5'd0, 27'h000000bc, 5'd13, 27'h000002f4, 32'h00000400,
  1'd1,  5'd27, 27'h00000247, 5'd3, 27'h000001f7, 5'd22, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000348, 5'd15, 27'h000001a2, 5'd3, 27'h0000021e, 32'h00000400,
  1'd1,  5'd26, 27'h000000cf, 5'd12, 27'h00000189, 5'd14, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c8, 5'd10, 27'h00000371, 5'd23, 27'h00000217, 32'h00000400,
  1'd1,  5'd27, 27'h0000025c, 5'd21, 27'h00000104, 5'd1, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000165, 5'd23, 27'h000001ae, 5'd11, 27'h00000133, 32'h00000400,
  1'd1,  5'd28, 27'h00000383, 5'd24, 27'h00000382, 5'd21, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000296, 5'd4, 27'h0000020a, 5'd3, 27'h00000254, 32'h00000400,
  1'd1,  5'd9, 27'h000000c2, 5'd0, 27'h00000231, 5'd14, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000252, 5'd5, 27'h0000000a, 5'd25, 27'h000000be, 32'h00000400,
  1'd1,  5'd5, 27'h000002b0, 5'd13, 27'h00000291, 5'd9, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002fb, 5'd14, 27'h00000197, 5'd17, 27'h0000027b, 32'h00000400,
  1'd1,  5'd9, 27'h00000210, 5'd11, 27'h00000016, 5'd27, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000006f, 5'd21, 27'h00000141, 5'd7, 27'h00000372, 32'h00000400,
  1'd1,  5'd8, 27'h000000d2, 5'd21, 27'h000000d8, 5'd18, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012b, 5'd21, 27'h000002b5, 5'd30, 27'h000003d7, 32'h00000400,
  1'd1,  5'd18, 27'h0000036c, 5'd2, 27'h000002e4, 5'd1, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001a, 5'd2, 27'h00000045, 5'd10, 27'h00000222, 32'h00000400,
  1'd1,  5'd20, 27'h0000015e, 5'd4, 27'h00000160, 5'd24, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000227, 5'd15, 27'h000000c5, 5'd10, 27'h0000010b, 32'h00000400,
  1'd1,  5'd17, 27'h000001ab, 5'd10, 27'h000001a2, 5'd17, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011d, 5'd13, 27'h000000c0, 5'd29, 27'h0000002d, 32'h00000400,
  1'd1,  5'd18, 27'h0000023d, 5'd23, 27'h00000150, 5'd7, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003f8, 5'd22, 27'h00000328, 5'd16, 27'h00000332, 32'h00000400,
  1'd1,  5'd18, 27'h000003b6, 5'd21, 27'h0000008f, 5'd28, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ac, 5'd4, 27'h0000038e, 5'd7, 27'h0000006a, 32'h00000400,
  1'd1,  5'd28, 27'h000003b2, 5'd3, 27'h00000217, 5'd16, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d5, 5'd3, 27'h00000394, 5'd28, 27'h00000214, 32'h00000400,
  1'd1,  5'd30, 27'h00000074, 5'd12, 27'h00000172, 5'd10, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000274, 5'd11, 27'h0000034a, 5'd19, 27'h000000ff, 32'h00000400,
  1'd1,  5'd26, 27'h0000022d, 5'd12, 27'h000000dc, 5'd30, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a4, 5'd24, 27'h000003a4, 5'd7, 27'h00000099, 32'h00000400,
  1'd1,  5'd28, 27'h00000288, 5'd21, 27'h00000107, 5'd16, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002cc, 5'd24, 27'h000000f4, 5'd29, 27'h00000345, 32'h00000400,
  1'd1,  5'd6, 27'h00000224, 5'd10, 27'h000000ff, 5'd0, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002c3, 5'd6, 27'h000000c9, 5'd13, 27'h00000343, 32'h00000400,
  1'd1,  5'd6, 27'h000000fc, 5'd5, 27'h00000293, 5'd21, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001fc, 5'd18, 27'h00000400, 5'd2, 27'h000003e6, 32'h00000400,
  1'd1,  5'd6, 27'h00000350, 5'd17, 27'h00000198, 5'd11, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000101, 5'd15, 27'h0000027b, 5'd25, 27'h00000080, 32'h00000400,
  1'd1,  5'd7, 27'h00000345, 5'd28, 27'h0000032a, 5'd4, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000161, 5'd28, 27'h000000b7, 5'd12, 27'h0000017b, 32'h00000400,
  1'd1,  5'd5, 27'h0000019c, 5'd27, 27'h00000176, 5'd22, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000107, 5'd5, 27'h000001bd, 5'd0, 27'h000000ed, 32'h00000400,
  1'd1,  5'd18, 27'h000002ba, 5'd8, 27'h0000002c, 5'd14, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000220, 5'd7, 27'h00000339, 5'd22, 27'h0000000b, 32'h00000400,
  1'd1,  5'd19, 27'h000002f9, 5'd16, 27'h00000019, 5'd2, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000019b, 5'd16, 27'h00000189, 5'd15, 27'h0000000b, 32'h00000400,
  1'd1,  5'd19, 27'h00000197, 5'd16, 27'h00000095, 5'd23, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000262, 5'd28, 27'h00000341, 5'd3, 27'h0000016c, 32'h00000400,
  1'd1,  5'd18, 27'h000000b8, 5'd29, 27'h00000108, 5'd10, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003b3, 5'd27, 27'h00000356, 5'd21, 27'h0000032d, 32'h00000400,
  1'd1,  5'd28, 27'h00000288, 5'd8, 27'h00000065, 5'd3, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000375, 5'd8, 27'h000003ce, 5'd15, 27'h000001c5, 32'h00000400,
  1'd1,  5'd26, 27'h000001de, 5'd5, 27'h000002ac, 5'd23, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000022, 5'd16, 27'h000000eb, 5'd3, 27'h00000080, 32'h00000400,
  1'd1,  5'd26, 27'h00000219, 5'd18, 27'h000001f0, 5'd14, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000001b, 5'd17, 27'h00000100, 5'd21, 27'h000002dd, 32'h00000400,
  1'd1,  5'd28, 27'h000001f3, 5'd27, 27'h00000060, 5'd0, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b4, 5'd27, 27'h000003f6, 5'd11, 27'h00000044, 32'h00000400,
  1'd1,  5'd29, 27'h0000000e, 5'd26, 27'h000000d5, 5'd25, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001b5, 5'd9, 27'h00000125, 5'd7, 27'h000002f5, 32'h00000400,
  1'd1,  5'd7, 27'h000001fe, 5'd7, 27'h00000327, 5'd20, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001cb, 5'd7, 27'h0000030f, 5'd29, 27'h0000020e, 32'h00000400,
  1'd1,  5'd8, 27'h0000002c, 5'd17, 27'h000003d0, 5'd10, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a3, 5'd17, 27'h000002b7, 5'd20, 27'h00000225, 32'h00000400,
  1'd1,  5'd8, 27'h00000222, 5'd18, 27'h000003b0, 5'd30, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000026, 5'd27, 27'h00000194, 5'd6, 27'h0000005a, 32'h00000400,
  1'd1,  5'd8, 27'h0000037b, 5'd30, 27'h000001cd, 5'd18, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a3, 5'd30, 27'h000000c0, 5'd27, 27'h00000319, 32'h00000400,
  1'd1,  5'd15, 27'h000002ba, 5'd5, 27'h0000021f, 5'd8, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000023e, 5'd9, 27'h00000132, 5'd17, 27'h00000103, 32'h00000400,
  1'd1,  5'd19, 27'h00000306, 5'd5, 27'h000003f0, 5'd29, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d5, 5'd18, 27'h0000015e, 5'd5, 27'h000000ac, 32'h00000400,
  1'd1,  5'd17, 27'h000001a4, 5'd17, 27'h00000308, 5'd18, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000036f, 5'd19, 27'h00000195, 5'd27, 27'h0000004f, 32'h00000400,
  1'd1,  5'd19, 27'h00000248, 5'd27, 27'h00000222, 5'd6, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003fa, 5'd28, 27'h000002d3, 5'd19, 27'h00000148, 32'h00000400,
  1'd1,  5'd19, 27'h000003c1, 5'd26, 27'h00000312, 5'd29, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001d6, 5'd10, 27'h00000060, 5'd5, 27'h00000174, 32'h00000400,
  1'd1,  5'd29, 27'h000002bc, 5'd10, 27'h000000d3, 5'd17, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000041, 5'd5, 27'h000000fd, 5'd26, 27'h0000021c, 32'h00000400,
  1'd1,  5'd26, 27'h00000145, 5'd17, 27'h00000124, 5'd6, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000087, 5'd19, 27'h000001a1, 5'd18, 27'h0000035f, 32'h00000400,
  1'd1,  5'd29, 27'h000002d6, 5'd18, 27'h00000019, 5'd28, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000016b, 5'd29, 27'h000003b7, 5'd9, 27'h000000bd, 32'h00000400,
  1'd1,  5'd29, 27'h00000257, 5'd27, 27'h000000cd, 5'd17, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003e5, 5'd26, 27'h00000341, 5'd30, 27'h0000002a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000013b, 5'd1, 27'h00000270, 5'd4, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001dd, 5'd2, 27'h0000014e, 5'd10, 27'h0000024c, 32'h00000400,
  1'd1,  5'd0, 27'h000000be, 5'd3, 27'h000003ed, 5'd21, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a4, 5'd13, 27'h00000369, 5'd1, 27'h000001f8, 32'h00000400,
  1'd1,  5'd4, 27'h00000243, 5'd13, 27'h0000018f, 5'd11, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000056, 5'd15, 27'h0000015c, 5'd24, 27'h00000219, 32'h00000400,
  1'd1,  5'd1, 27'h0000012c, 5'd24, 27'h00000276, 5'd0, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000039, 5'd23, 27'h00000380, 5'd14, 27'h0000001d, 32'h00000400,
  1'd1,  5'd0, 27'h000003f0, 5'd22, 27'h0000038d, 5'd24, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d6, 5'd4, 27'h00000230, 5'd5, 27'h00000042, 32'h00000400,
  1'd1,  5'd10, 27'h000002bf, 5'd4, 27'h000001e9, 5'd12, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000007d, 5'd0, 27'h00000195, 5'd23, 27'h00000208, 32'h00000400,
  1'd1,  5'd11, 27'h000001f5, 5'd12, 27'h000000a4, 5'd0, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000288, 5'd13, 27'h00000171, 5'd11, 27'h00000067, 32'h00000400,
  1'd1,  5'd11, 27'h000001a3, 5'd12, 27'h00000146, 5'd20, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000353, 5'd21, 27'h00000239, 5'd1, 27'h00000315, 32'h00000400,
  1'd1,  5'd10, 27'h000003e2, 5'd22, 27'h000000f4, 5'd11, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002ad, 5'd21, 27'h00000290, 5'd24, 27'h0000036c, 32'h00000400,
  1'd1,  5'd23, 27'h0000039c, 5'd0, 27'h0000037c, 5'd0, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000019d, 5'd2, 27'h00000194, 5'd13, 27'h00000026, 32'h00000400,
  1'd1,  5'd23, 27'h000000dc, 5'd2, 27'h00000144, 5'd21, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022f, 5'd12, 27'h00000336, 5'd0, 27'h000000c5, 32'h00000400,
  1'd1,  5'd22, 27'h0000026e, 5'd14, 27'h00000144, 5'd12, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000187, 5'd14, 27'h0000006b, 5'd24, 27'h000000f8, 32'h00000400,
  1'd1,  5'd24, 27'h0000033a, 5'd24, 27'h00000020, 5'd2, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002fe, 5'd24, 27'h00000199, 5'd11, 27'h00000218, 32'h00000400,
  1'd1,  5'd22, 27'h0000026f, 5'd23, 27'h000000a9, 5'd21, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000336, 5'd1, 27'h00000334, 5'd6, 27'h00000228, 32'h00000400,
  1'd1,  5'd1, 27'h000000c4, 5'd4, 27'h000001fa, 5'd18, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000084, 5'd5, 27'h00000005, 5'd26, 27'h0000027f, 32'h00000400,
  1'd1,  5'd0, 27'h000000d3, 5'd14, 27'h000003ab, 5'd7, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017a, 5'd15, 27'h000000ad, 5'd18, 27'h00000117, 32'h00000400,
  1'd1,  5'd2, 27'h0000036c, 5'd10, 27'h00000292, 5'd30, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ac, 5'd24, 27'h00000023, 5'd5, 27'h00000147, 32'h00000400,
  1'd1,  5'd0, 27'h000001a4, 5'd23, 27'h000003b1, 5'd16, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000f6, 5'd22, 27'h00000232, 5'd30, 27'h000003e4, 32'h00000400,
  1'd1,  5'd13, 27'h00000048, 5'd0, 27'h00000113, 5'd5, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003a5, 5'd4, 27'h00000236, 5'd15, 27'h00000283, 32'h00000400,
  1'd1,  5'd12, 27'h0000025e, 5'd3, 27'h000002a7, 5'd27, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002b4, 5'd11, 27'h00000120, 5'd9, 27'h0000016c, 32'h00000400,
  1'd1,  5'd13, 27'h000000d8, 5'd13, 27'h000000ee, 5'd16, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000344, 5'd12, 27'h000002e4, 5'd28, 27'h000002d9, 32'h00000400,
  1'd1,  5'd15, 27'h0000019b, 5'd22, 27'h00000109, 5'd7, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001e3, 5'd21, 27'h00000260, 5'd15, 27'h000003f9, 32'h00000400,
  1'd1,  5'd14, 27'h000001be, 5'd25, 27'h000002f1, 5'd30, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000217, 5'd1, 27'h00000361, 5'd8, 27'h0000024d, 32'h00000400,
  1'd1,  5'd23, 27'h000002f1, 5'd1, 27'h0000012a, 5'd20, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000271, 5'd1, 27'h0000024e, 5'd29, 27'h00000013, 32'h00000400,
  1'd1,  5'd25, 27'h00000103, 5'd14, 27'h00000267, 5'd9, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ae, 5'd13, 27'h000003bf, 5'd19, 27'h000001d7, 32'h00000400,
  1'd1,  5'd25, 27'h0000016a, 5'd13, 27'h000003d2, 5'd27, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d5, 5'd22, 27'h000000cf, 5'd8, 27'h000002f8, 32'h00000400,
  1'd1,  5'd23, 27'h000001d6, 5'd21, 27'h00000248, 5'd19, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003cd, 5'd23, 27'h00000304, 5'd29, 27'h0000010e, 32'h00000400,
  1'd1,  5'd4, 27'h00000204, 5'd8, 27'h0000038a, 5'd0, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a4, 5'd7, 27'h0000013f, 5'd10, 27'h000001b6, 32'h00000400,
  1'd1,  5'd2, 27'h0000017a, 5'd5, 27'h000002e9, 5'd21, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000b7, 5'd17, 27'h0000034e, 5'd1, 27'h000002b9, 32'h00000400,
  1'd1,  5'd4, 27'h000000c2, 5'd19, 27'h000001da, 5'd14, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000012, 5'd16, 27'h0000014d, 5'd21, 27'h00000093, 32'h00000400,
  1'd1,  5'd1, 27'h000003a6, 5'd29, 27'h00000202, 5'd2, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000373, 5'd26, 27'h0000033a, 5'd15, 27'h000000aa, 32'h00000400,
  1'd1,  5'd4, 27'h00000335, 5'd27, 27'h0000021f, 5'd22, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003fa, 5'd5, 27'h000000e8, 5'd3, 27'h000000ed, 32'h00000400,
  1'd1,  5'd10, 27'h00000291, 5'd10, 27'h0000008a, 5'd10, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001cf, 5'd9, 27'h000003e6, 5'd25, 27'h00000064, 32'h00000400,
  1'd1,  5'd13, 27'h00000073, 5'd17, 27'h0000039a, 5'd4, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f8, 5'd20, 27'h0000017f, 5'd13, 27'h000000ea, 32'h00000400,
  1'd1,  5'd14, 27'h00000269, 5'd19, 27'h000001a1, 5'd24, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000df, 5'd27, 27'h000001a1, 5'd1, 27'h00000117, 32'h00000400,
  1'd1,  5'd14, 27'h000000bc, 5'd26, 27'h000001b9, 5'd11, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000dc, 5'd29, 27'h000000c4, 5'd21, 27'h00000372, 32'h00000400,
  1'd1,  5'd23, 27'h000002fa, 5'd7, 27'h00000189, 5'd1, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002f1, 5'd6, 27'h00000199, 5'd12, 27'h00000045, 32'h00000400,
  1'd1,  5'd21, 27'h0000011b, 5'd9, 27'h00000043, 5'd21, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000092, 5'd16, 27'h0000025f, 5'd2, 27'h0000035a, 32'h00000400,
  1'd1,  5'd23, 27'h0000028d, 5'd16, 27'h00000293, 5'd13, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000048, 5'd15, 27'h000002f6, 5'd20, 27'h00000383, 32'h00000400,
  1'd1,  5'd24, 27'h0000005b, 5'd26, 27'h00000205, 5'd3, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000251, 5'd25, 27'h00000358, 5'd15, 27'h000001f9, 32'h00000400,
  1'd1,  5'd24, 27'h00000267, 5'd28, 27'h0000009b, 5'd22, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000175, 5'd6, 27'h00000195, 5'd9, 27'h00000281, 32'h00000400,
  1'd1,  5'd2, 27'h00000123, 5'd9, 27'h0000029d, 5'd19, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000022b, 5'd7, 27'h00000097, 5'd29, 27'h000003c5, 32'h00000400,
  1'd1,  5'd2, 27'h000002ec, 5'd17, 27'h0000016b, 5'd7, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000007e, 5'd16, 27'h0000034f, 5'd18, 27'h000002fc, 32'h00000400,
  1'd1,  5'd0, 27'h000000a3, 5'd16, 27'h0000007d, 5'd30, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000277, 5'd27, 27'h000003c5, 5'd7, 27'h00000173, 32'h00000400,
  1'd1,  5'd4, 27'h0000025e, 5'd26, 27'h000002b3, 5'd18, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000031e, 5'd30, 27'h000000de, 5'd27, 27'h00000229, 32'h00000400,
  1'd1,  5'd10, 27'h000001c2, 5'd6, 27'h00000058, 5'd7, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c7, 5'd6, 27'h000001e5, 5'd18, 27'h000003ab, 32'h00000400,
  1'd1,  5'd13, 27'h000000d4, 5'd9, 27'h00000325, 5'd26, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d4, 5'd16, 27'h00000085, 5'd9, 27'h0000001f, 32'h00000400,
  1'd1,  5'd13, 27'h000000e5, 5'd16, 27'h00000111, 5'd18, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000036, 5'd19, 27'h000000ba, 5'd26, 27'h000000bf, 32'h00000400,
  1'd1,  5'd15, 27'h000000ed, 5'd29, 27'h0000026c, 5'd7, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000162, 5'd30, 27'h00000176, 5'd17, 27'h00000031, 32'h00000400,
  1'd1,  5'd10, 27'h00000272, 5'd30, 27'h00000270, 5'd28, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001c9, 5'd7, 27'h0000002e, 5'd10, 27'h0000005a, 32'h00000400,
  1'd1,  5'd21, 27'h00000168, 5'd9, 27'h00000139, 5'd17, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002fc, 5'd7, 27'h0000018c, 5'd29, 27'h000003c3, 32'h00000400,
  1'd1,  5'd23, 27'h00000393, 5'd17, 27'h000000ec, 5'd9, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b3, 5'd18, 27'h00000279, 5'd19, 27'h00000141, 32'h00000400,
  1'd1,  5'd21, 27'h00000147, 5'd16, 27'h00000331, 5'd26, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000073, 5'd26, 27'h000001ea, 5'd6, 27'h00000312, 32'h00000400,
  1'd1,  5'd21, 27'h0000035b, 5'd25, 27'h000003ff, 5'd18, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000030c, 5'd30, 27'h000002a3, 5'd28, 27'h00000205, 32'h00000400,
  1'd1,  5'd7, 27'h000002f5, 5'd5, 27'h0000002c, 5'd6, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ed, 5'd0, 27'h00000218, 5'd20, 27'h00000003, 32'h00000400,
  1'd1,  5'd5, 27'h000002ab, 5'd3, 27'h0000016f, 5'd28, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000016e, 5'd10, 27'h0000028f, 5'd0, 27'h000003d9, 32'h00000400,
  1'd1,  5'd5, 27'h00000217, 5'd11, 27'h0000032e, 5'd12, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000131, 5'd14, 27'h000000f8, 5'd22, 27'h00000231, 32'h00000400,
  1'd1,  5'd9, 27'h000001ce, 5'd21, 27'h000000c5, 5'd0, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000277, 5'd22, 27'h00000035, 5'd11, 27'h00000068, 32'h00000400,
  1'd1,  5'd5, 27'h00000316, 5'd25, 27'h00000233, 5'd23, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000156, 5'd2, 27'h00000009, 5'd6, 27'h0000014c, 32'h00000400,
  1'd1,  5'd17, 27'h0000001c, 5'd4, 27'h0000002c, 5'd18, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ac, 5'd2, 27'h00000171, 5'd30, 27'h000003d6, 32'h00000400,
  1'd1,  5'd17, 27'h000002df, 5'd13, 27'h000000b8, 5'd4, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003db, 5'd10, 27'h0000032e, 5'd13, 27'h0000036f, 32'h00000400,
  1'd1,  5'd15, 27'h00000236, 5'd14, 27'h0000008f, 5'd24, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000382, 5'd22, 27'h0000008d, 5'd1, 27'h000002b8, 32'h00000400,
  1'd1,  5'd15, 27'h00000392, 5'd23, 27'h00000021, 5'd13, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000016, 5'd25, 27'h00000207, 5'd23, 27'h000001a7, 32'h00000400,
  1'd1,  5'd27, 27'h0000036c, 5'd3, 27'h00000325, 5'd0, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002dc, 5'd0, 27'h0000032f, 5'd14, 27'h000001b1, 32'h00000400,
  1'd1,  5'd28, 27'h000002b2, 5'd3, 27'h00000127, 5'd25, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000004, 5'd13, 27'h00000089, 5'd1, 27'h0000008d, 32'h00000400,
  1'd1,  5'd28, 27'h00000137, 5'd12, 27'h00000158, 5'd11, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b5, 5'd13, 27'h000000e2, 5'd24, 27'h000002d4, 32'h00000400,
  1'd1,  5'd30, 27'h0000027a, 5'd22, 27'h000001e2, 5'd1, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000031c, 5'd23, 27'h000003d7, 5'd14, 27'h00000126, 32'h00000400,
  1'd1,  5'd26, 27'h00000150, 5'd24, 27'h000003ca, 5'd25, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e7, 5'd3, 27'h000003a4, 5'd1, 27'h000002fd, 32'h00000400,
  1'd1,  5'd10, 27'h000000aa, 5'd3, 27'h000003d0, 5'd12, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003e8, 5'd4, 27'h00000210, 5'd23, 27'h000001e0, 32'h00000400,
  1'd1,  5'd6, 27'h00000265, 5'd11, 27'h000001f1, 5'd9, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000341, 5'd14, 27'h00000344, 5'd19, 27'h00000058, 32'h00000400,
  1'd1,  5'd7, 27'h00000041, 5'd15, 27'h000000d2, 5'd29, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000305, 5'd21, 27'h000000d0, 5'd6, 27'h000000f2, 32'h00000400,
  1'd1,  5'd7, 27'h000002bc, 5'd25, 27'h000001b5, 5'd18, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000386, 5'd23, 27'h0000033a, 5'd26, 27'h000003af, 32'h00000400,
  1'd1,  5'd19, 27'h000000c9, 5'd1, 27'h000002dd, 5'd2, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000162, 5'd1, 27'h00000011, 5'd15, 27'h000001e6, 32'h00000400,
  1'd1,  5'd18, 27'h000003eb, 5'd0, 27'h000003a4, 5'd24, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000130, 5'd12, 27'h00000141, 5'd10, 27'h00000058, 32'h00000400,
  1'd1,  5'd16, 27'h0000025b, 5'd14, 27'h00000302, 5'd17, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025d, 5'd12, 27'h0000027a, 5'd26, 27'h000003ba, 32'h00000400,
  1'd1,  5'd15, 27'h00000376, 5'd22, 27'h00000063, 5'd6, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d5, 5'd24, 27'h0000038f, 5'd17, 27'h0000017c, 32'h00000400,
  1'd1,  5'd17, 27'h00000145, 5'd22, 27'h00000191, 5'd27, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000248, 5'd3, 27'h00000233, 5'd10, 27'h0000002c, 32'h00000400,
  1'd1,  5'd26, 27'h000001e1, 5'd2, 27'h0000038b, 5'd19, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000210, 5'd5, 27'h0000007a, 5'd28, 27'h00000042, 32'h00000400,
  1'd1,  5'd26, 27'h000001e4, 5'd11, 27'h000001d3, 5'd6, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000396, 5'd15, 27'h000001a1, 5'd17, 27'h00000310, 32'h00000400,
  1'd1,  5'd28, 27'h00000260, 5'd12, 27'h00000337, 5'd28, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000a1, 5'd21, 27'h00000338, 5'd8, 27'h000002a8, 32'h00000400,
  1'd1,  5'd26, 27'h0000002a, 5'd21, 27'h000000cf, 5'd15, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000035, 5'd23, 27'h000000cc, 5'd27, 27'h000000bd, 32'h00000400,
  1'd1,  5'd9, 27'h00000010, 5'd7, 27'h000000af, 5'd2, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000004e, 5'd6, 27'h000001b3, 5'd14, 27'h0000019e, 32'h00000400,
  1'd1,  5'd9, 27'h00000013, 5'd9, 27'h00000203, 5'd20, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002f7, 5'd20, 27'h000000c1, 5'd1, 27'h00000280, 32'h00000400,
  1'd1,  5'd5, 27'h0000035c, 5'd15, 27'h00000204, 5'd15, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005b, 5'd19, 27'h00000165, 5'd21, 27'h00000343, 32'h00000400,
  1'd1,  5'd6, 27'h00000234, 5'd26, 27'h00000295, 5'd4, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b6, 5'd26, 27'h00000346, 5'd14, 27'h0000015d, 32'h00000400,
  1'd1,  5'd10, 27'h00000039, 5'd29, 27'h00000132, 5'd24, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000060, 5'd6, 27'h00000384, 5'd1, 27'h00000398, 32'h00000400,
  1'd1,  5'd15, 27'h00000385, 5'd6, 27'h00000283, 5'd15, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000363, 5'd8, 27'h00000296, 5'd22, 27'h00000042, 32'h00000400,
  1'd1,  5'd17, 27'h000000fb, 5'd20, 27'h00000095, 5'd1, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000099, 5'd19, 27'h0000024e, 5'd12, 27'h0000038b, 32'h00000400,
  1'd1,  5'd18, 27'h00000005, 5'd18, 27'h000000da, 5'd21, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002cd, 5'd28, 27'h000002fb, 5'd3, 27'h0000016f, 32'h00000400,
  1'd1,  5'd16, 27'h0000032d, 5'd30, 27'h000003f5, 5'd14, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000125, 5'd27, 27'h00000020, 5'd24, 27'h0000020f, 32'h00000400,
  1'd1,  5'd30, 27'h00000023, 5'd8, 27'h00000233, 5'd3, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000003a, 5'd7, 27'h000001e1, 5'd10, 27'h000001fc, 32'h00000400,
  1'd1,  5'd30, 27'h00000099, 5'd6, 27'h00000072, 5'd25, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e4, 5'd16, 27'h00000018, 5'd4, 27'h0000019e, 32'h00000400,
  1'd1,  5'd28, 27'h00000339, 5'd17, 27'h0000039d, 5'd12, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000143, 5'd17, 27'h000000c1, 5'd23, 27'h00000144, 32'h00000400,
  1'd1,  5'd26, 27'h0000035d, 5'd30, 27'h000002f3, 5'd2, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000022, 5'd27, 27'h00000340, 5'd12, 27'h000002d5, 32'h00000400,
  1'd1,  5'd27, 27'h0000024d, 5'd29, 27'h0000000d, 5'd22, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000331, 5'd7, 27'h000003da, 5'd8, 27'h00000160, 32'h00000400,
  1'd1,  5'd5, 27'h000001e7, 5'd7, 27'h000003f3, 5'd18, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000161, 5'd6, 27'h000003a5, 5'd27, 27'h00000382, 32'h00000400,
  1'd1,  5'd7, 27'h0000029c, 5'd20, 27'h000001f0, 5'd10, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000172, 5'd17, 27'h000002e0, 5'd16, 27'h00000211, 32'h00000400,
  1'd1,  5'd5, 27'h000002e2, 5'd17, 27'h0000003e, 5'd27, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000028d, 5'd26, 27'h0000000b, 5'd8, 27'h00000141, 32'h00000400,
  1'd1,  5'd8, 27'h000001c6, 5'd27, 27'h0000018b, 5'd19, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000018, 5'd30, 27'h0000017e, 5'd27, 27'h00000210, 32'h00000400,
  1'd1,  5'd20, 27'h000000ff, 5'd8, 27'h0000017e, 5'd5, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001da, 5'd5, 27'h000001f1, 5'd16, 27'h00000052, 32'h00000400,
  1'd1,  5'd16, 27'h00000247, 5'd6, 27'h00000204, 5'd29, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000072, 5'd17, 27'h00000081, 5'd9, 27'h00000025, 32'h00000400,
  1'd1,  5'd16, 27'h00000171, 5'd17, 27'h00000172, 5'd17, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003f8, 5'd19, 27'h00000038, 5'd28, 27'h000002c8, 32'h00000400,
  1'd1,  5'd20, 27'h00000024, 5'd30, 27'h000003de, 5'd7, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c6, 5'd29, 27'h00000028, 5'd19, 27'h00000051, 32'h00000400,
  1'd1,  5'd17, 27'h00000298, 5'd27, 27'h00000280, 5'd29, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003d0, 5'd9, 27'h00000069, 5'd9, 27'h000002a0, 32'h00000400,
  1'd1,  5'd29, 27'h00000296, 5'd7, 27'h000000d6, 5'd20, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ed, 5'd7, 27'h000003ab, 5'd30, 27'h00000275, 32'h00000400,
  1'd1,  5'd30, 27'h00000017, 5'd19, 27'h0000035d, 5'd7, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000036d, 5'd18, 27'h0000010f, 5'd15, 27'h0000027b, 32'h00000400,
  1'd1,  5'd30, 27'h00000092, 5'd17, 27'h00000093, 5'd26, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000021d, 5'd30, 27'h00000322, 5'd8, 27'h000002b5, 32'h00000400,
  1'd1,  5'd30, 27'h000002f6, 5'd29, 27'h000000ad, 5'd17, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000011b, 5'd27, 27'h000001ab, 5'd29, 27'h000003cd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h0000009b, 5'd0, 27'h0000037b, 5'd4, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000156, 5'd2, 27'h0000008e, 5'd14, 27'h000002a3, 32'h00000400,
  1'd1,  5'd0, 27'h000001f4, 5'd3, 27'h000001c3, 5'd21, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f8, 5'd12, 27'h00000036, 5'd5, 27'h0000003e, 32'h00000400,
  1'd1,  5'd4, 27'h000000dd, 5'd10, 27'h000001a4, 5'd15, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001fe, 5'd13, 27'h000001a1, 5'd22, 27'h0000003d, 32'h00000400,
  1'd1,  5'd1, 27'h0000017a, 5'd20, 27'h0000033b, 5'd4, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b6, 5'd20, 27'h00000340, 5'd15, 27'h00000081, 32'h00000400,
  1'd1,  5'd2, 27'h0000020f, 5'd24, 27'h00000353, 5'd22, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000025c, 5'd0, 27'h0000008f, 5'd0, 27'h00000220, 32'h00000400,
  1'd1,  5'd12, 27'h00000123, 5'd0, 27'h0000022b, 5'd14, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000225, 5'd0, 27'h00000324, 5'd22, 27'h00000398, 32'h00000400,
  1'd1,  5'd12, 27'h00000105, 5'd10, 27'h00000324, 5'd3, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000035a, 5'd10, 27'h0000038b, 5'd15, 27'h000000f3, 32'h00000400,
  1'd1,  5'd12, 27'h00000278, 5'd12, 27'h00000160, 5'd25, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001fd, 5'd21, 27'h00000283, 5'd2, 27'h000000c2, 32'h00000400,
  1'd1,  5'd11, 27'h000002f1, 5'd22, 27'h00000284, 5'd10, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000334, 5'd25, 27'h0000021c, 5'd21, 27'h000001c6, 32'h00000400,
  1'd1,  5'd21, 27'h0000007d, 5'd4, 27'h00000146, 5'd3, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002b2, 5'd2, 27'h00000320, 5'd11, 27'h0000005a, 32'h00000400,
  1'd1,  5'd20, 27'h00000341, 5'd3, 27'h00000128, 5'd23, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000364, 5'd14, 27'h000002b0, 5'd3, 27'h0000035a, 32'h00000400,
  1'd1,  5'd25, 27'h000000e0, 5'd15, 27'h000001f0, 5'd13, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000116, 5'd15, 27'h0000016d, 5'd25, 27'h000002ac, 32'h00000400,
  1'd1,  5'd21, 27'h0000025a, 5'd24, 27'h0000002c, 5'd0, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003cd, 5'd24, 27'h0000024f, 5'd10, 27'h0000030e, 32'h00000400,
  1'd1,  5'd21, 27'h000001f1, 5'd25, 27'h0000033f, 5'd22, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d8, 5'd1, 27'h00000322, 5'd5, 27'h000003b3, 32'h00000400,
  1'd1,  5'd3, 27'h0000004e, 5'd1, 27'h000002e6, 5'd19, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000069, 5'd2, 27'h000003d4, 5'd28, 27'h000001a5, 32'h00000400,
  1'd1,  5'd1, 27'h000001a8, 5'd11, 27'h0000002d, 5'd8, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001b6, 5'd11, 27'h00000006, 5'd19, 27'h0000023f, 32'h00000400,
  1'd1,  5'd3, 27'h000000d4, 5'd11, 27'h000000d6, 5'd29, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000273, 5'd20, 27'h000002c1, 5'd6, 27'h0000000d, 32'h00000400,
  1'd1,  5'd4, 27'h000002ab, 5'd21, 27'h00000322, 5'd17, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000037c, 5'd22, 27'h00000012, 5'd30, 27'h00000322, 32'h00000400,
  1'd1,  5'd15, 27'h00000059, 5'd4, 27'h000000dc, 5'd6, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000db, 5'd0, 27'h0000033e, 5'd16, 27'h000002bc, 32'h00000400,
  1'd1,  5'd14, 27'h000002b6, 5'd4, 27'h000000d2, 5'd28, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000fc, 5'd14, 27'h00000132, 5'd9, 27'h000003c1, 32'h00000400,
  1'd1,  5'd10, 27'h00000305, 5'd15, 27'h000001b4, 5'd19, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000272, 5'd14, 27'h000000ee, 5'd28, 27'h000001e2, 32'h00000400,
  1'd1,  5'd14, 27'h0000006b, 5'd22, 27'h0000005a, 5'd6, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000121, 5'd24, 27'h000000ef, 5'd20, 27'h00000080, 32'h00000400,
  1'd1,  5'd13, 27'h00000132, 5'd24, 27'h000003e8, 5'd29, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000144, 5'd2, 27'h0000030c, 5'd8, 27'h000000ab, 32'h00000400,
  1'd1,  5'd22, 27'h000001a4, 5'd3, 27'h00000381, 5'd17, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003de, 5'd4, 27'h000002c6, 5'd29, 27'h000000dc, 32'h00000400,
  1'd1,  5'd23, 27'h000000e9, 5'd14, 27'h00000236, 5'd8, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a3, 5'd14, 27'h0000022e, 5'd20, 27'h0000014e, 32'h00000400,
  1'd1,  5'd21, 27'h00000374, 5'd14, 27'h00000208, 5'd27, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000199, 5'd21, 27'h00000203, 5'd9, 27'h00000210, 32'h00000400,
  1'd1,  5'd21, 27'h0000001a, 5'd21, 27'h00000099, 5'd18, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000332, 5'd23, 27'h00000014, 5'd27, 27'h000003db, 32'h00000400,
  1'd1,  5'd1, 27'h000001da, 5'd5, 27'h00000288, 5'd4, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c5, 5'd9, 27'h00000242, 5'd14, 27'h0000027d, 32'h00000400,
  1'd1,  5'd0, 27'h000000e9, 5'd8, 27'h0000008f, 5'd25, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001aa, 5'd15, 27'h000003ba, 5'd4, 27'h00000113, 32'h00000400,
  1'd1,  5'd2, 27'h000001b9, 5'd18, 27'h000002bb, 5'd12, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000392, 5'd18, 27'h0000011c, 5'd23, 27'h000002ed, 32'h00000400,
  1'd1,  5'd4, 27'h00000019, 5'd28, 27'h000003fa, 5'd0, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002ed, 5'd28, 27'h00000368, 5'd13, 27'h000003bb, 32'h00000400,
  1'd1,  5'd2, 27'h000001f9, 5'd27, 27'h00000302, 5'd25, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000004e, 5'd5, 27'h00000190, 5'd2, 27'h000002c2, 32'h00000400,
  1'd1,  5'd12, 27'h000003d0, 5'd10, 27'h00000079, 5'd14, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002b5, 5'd6, 27'h0000008b, 5'd22, 27'h0000025b, 32'h00000400,
  1'd1,  5'd11, 27'h000000f2, 5'd18, 27'h00000180, 5'd2, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000002b, 5'd17, 27'h0000039e, 5'd11, 27'h00000065, 32'h00000400,
  1'd1,  5'd12, 27'h00000015, 5'd16, 27'h0000016b, 5'd23, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000209, 5'd29, 27'h00000190, 5'd3, 27'h00000392, 32'h00000400,
  1'd1,  5'd13, 27'h00000374, 5'd28, 27'h00000017, 5'd14, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000036f, 5'd30, 27'h00000048, 5'd23, 27'h00000272, 32'h00000400,
  1'd1,  5'd25, 27'h00000249, 5'd6, 27'h00000269, 5'd1, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000033c, 5'd9, 27'h000003fa, 5'd14, 27'h0000002d, 32'h00000400,
  1'd1,  5'd21, 27'h0000002f, 5'd6, 27'h000001e3, 5'd25, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000018a, 5'd20, 27'h0000012b, 5'd3, 27'h00000303, 32'h00000400,
  1'd1,  5'd25, 27'h0000003d, 5'd17, 27'h00000115, 5'd11, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000120, 5'd19, 27'h0000036a, 5'd24, 27'h0000024c, 32'h00000400,
  1'd1,  5'd20, 27'h000002bf, 5'd28, 27'h00000172, 5'd0, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001c0, 5'd28, 27'h0000001a, 5'd14, 27'h000002fb, 32'h00000400,
  1'd1,  5'd24, 27'h000000c9, 5'd28, 27'h0000020f, 5'd24, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000001a, 5'd6, 27'h00000190, 5'd9, 27'h00000393, 32'h00000400,
  1'd1,  5'd2, 27'h000000bc, 5'd10, 27'h00000154, 5'd17, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001cb, 5'd6, 27'h00000088, 5'd29, 27'h0000015a, 32'h00000400,
  1'd1,  5'd0, 27'h00000398, 5'd16, 27'h000000a4, 5'd10, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002c9, 5'd19, 27'h00000069, 5'd19, 27'h00000128, 32'h00000400,
  1'd1,  5'd4, 27'h000003e3, 5'd20, 27'h00000253, 5'd28, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000264, 5'd26, 27'h000001d8, 5'd7, 27'h00000046, 32'h00000400,
  1'd1,  5'd3, 27'h0000003b, 5'd28, 27'h00000166, 5'd18, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001da, 5'd28, 27'h00000191, 5'd27, 27'h00000268, 32'h00000400,
  1'd1,  5'd12, 27'h000000df, 5'd6, 27'h000003c5, 5'd5, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000224, 5'd8, 27'h00000001, 5'd20, 27'h00000059, 32'h00000400,
  1'd1,  5'd13, 27'h00000322, 5'd10, 27'h0000009c, 5'd28, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000289, 5'd15, 27'h00000349, 5'd6, 27'h0000010f, 32'h00000400,
  1'd1,  5'd14, 27'h000001b6, 5'd15, 27'h0000037a, 5'd17, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000aa, 5'd17, 27'h0000020c, 5'd29, 27'h00000258, 32'h00000400,
  1'd1,  5'd12, 27'h00000374, 5'd26, 27'h00000263, 5'd6, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000077, 5'd27, 27'h0000038e, 5'd17, 27'h000002af, 32'h00000400,
  1'd1,  5'd14, 27'h00000179, 5'd28, 27'h00000380, 5'd29, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000ac, 5'd9, 27'h000003fc, 5'd10, 27'h00000151, 32'h00000400,
  1'd1,  5'd24, 27'h000003f1, 5'd6, 27'h00000261, 5'd18, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000182, 5'd9, 27'h00000159, 5'd28, 27'h00000017, 32'h00000400,
  1'd1,  5'd22, 27'h000000d7, 5'd16, 27'h000001c7, 5'd9, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000066, 5'd16, 27'h0000007b, 5'd19, 27'h00000216, 32'h00000400,
  1'd1,  5'd23, 27'h000003a4, 5'd16, 27'h00000348, 5'd26, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000000b, 5'd28, 27'h00000054, 5'd7, 27'h0000031b, 32'h00000400,
  1'd1,  5'd24, 27'h00000123, 5'd26, 27'h000003b0, 5'd18, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ae, 5'd27, 27'h000003e8, 5'd28, 27'h000003f8, 32'h00000400,
  1'd1,  5'd8, 27'h00000335, 5'd2, 27'h000000db, 5'd9, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000251, 5'd0, 27'h000003b5, 5'd19, 27'h0000039e, 32'h00000400,
  1'd1,  5'd10, 27'h00000132, 5'd2, 27'h000000f4, 5'd30, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000156, 5'd10, 27'h000002ff, 5'd3, 27'h00000365, 32'h00000400,
  1'd1,  5'd8, 27'h000002a4, 5'd14, 27'h000002c0, 5'd10, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ac, 5'd13, 27'h000002e3, 5'd24, 27'h0000022e, 32'h00000400,
  1'd1,  5'd9, 27'h000000ba, 5'd25, 27'h000000ba, 5'd0, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023b, 5'd24, 27'h000003d9, 5'd10, 27'h000002ac, 32'h00000400,
  1'd1,  5'd10, 27'h000000f3, 5'd21, 27'h00000338, 5'd23, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a3, 5'd1, 27'h00000097, 5'd8, 27'h0000023e, 32'h00000400,
  1'd1,  5'd19, 27'h00000255, 5'd1, 27'h000002b4, 5'd18, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000024f, 5'd0, 27'h000003fb, 5'd27, 27'h00000385, 32'h00000400,
  1'd1,  5'd20, 27'h0000017d, 5'd15, 27'h000001a7, 5'd4, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c2, 5'd13, 27'h000001c5, 5'd11, 27'h00000137, 32'h00000400,
  1'd1,  5'd16, 27'h000001d4, 5'd10, 27'h00000236, 5'd21, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001da, 5'd25, 27'h000001a1, 5'd3, 27'h00000243, 32'h00000400,
  1'd1,  5'd17, 27'h000001e0, 5'd20, 27'h000002ef, 5'd15, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f4, 5'd24, 27'h00000106, 5'd22, 27'h0000035e, 32'h00000400,
  1'd1,  5'd25, 27'h00000373, 5'd0, 27'h00000331, 5'd4, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f5, 5'd0, 27'h000003e2, 5'd10, 27'h000003af, 32'h00000400,
  1'd1,  5'd26, 27'h00000240, 5'd2, 27'h0000001b, 5'd23, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000035e, 5'd12, 27'h00000320, 5'd2, 27'h0000033f, 32'h00000400,
  1'd1,  5'd26, 27'h000001fc, 5'd13, 27'h000002f8, 5'd12, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001bd, 5'd15, 27'h00000120, 5'd25, 27'h00000108, 32'h00000400,
  1'd1,  5'd29, 27'h00000210, 5'd25, 27'h0000010a, 5'd0, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000265, 5'd24, 27'h000002c4, 5'd11, 27'h000001cb, 32'h00000400,
  1'd1,  5'd26, 27'h000000ed, 5'd24, 27'h00000093, 5'd20, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000162, 5'd3, 27'h00000216, 5'd0, 27'h000000cd, 32'h00000400,
  1'd1,  5'd5, 27'h0000027d, 5'd2, 27'h00000038, 5'd11, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000025d, 5'd3, 27'h000000a2, 5'd25, 27'h000000da, 32'h00000400,
  1'd1,  5'd7, 27'h000003a0, 5'd15, 27'h000000d0, 5'd9, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000132, 5'd11, 27'h000001cc, 5'd18, 27'h000000ac, 32'h00000400,
  1'd1,  5'd9, 27'h000000d0, 5'd13, 27'h00000164, 5'd29, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f4, 5'd25, 27'h0000031e, 5'd5, 27'h00000325, 32'h00000400,
  1'd1,  5'd9, 27'h0000009e, 5'd21, 27'h000002f6, 5'd19, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000384, 5'd23, 27'h000001de, 5'd29, 27'h000000b2, 32'h00000400,
  1'd1,  5'd20, 27'h0000013c, 5'd2, 27'h00000103, 5'd3, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000026a, 5'd0, 27'h000001a7, 5'd10, 27'h00000345, 32'h00000400,
  1'd1,  5'd18, 27'h00000079, 5'd5, 27'h00000099, 5'd25, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ee, 5'd14, 27'h0000014e, 5'd5, 27'h00000241, 32'h00000400,
  1'd1,  5'd17, 27'h00000399, 5'd14, 27'h00000023, 5'd17, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000b2, 5'd12, 27'h000000ab, 5'd28, 27'h00000082, 32'h00000400,
  1'd1,  5'd19, 27'h00000179, 5'd25, 27'h000001ec, 5'd8, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000080, 5'd21, 27'h0000037f, 5'd19, 27'h0000007b, 32'h00000400,
  1'd1,  5'd17, 27'h000002b5, 5'd21, 27'h000000df, 5'd26, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000258, 5'd3, 27'h000000ab, 5'd8, 27'h000003e5, 32'h00000400,
  1'd1,  5'd30, 27'h00000024, 5'd5, 27'h0000000a, 5'd19, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d0, 5'd0, 27'h000000d9, 5'd25, 27'h000003c4, 32'h00000400,
  1'd1,  5'd30, 27'h000001f7, 5'd14, 27'h00000072, 5'd9, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a2, 5'd12, 27'h00000380, 5'd18, 27'h000001a6, 32'h00000400,
  1'd1,  5'd28, 27'h000000f3, 5'd15, 27'h00000174, 5'd29, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ed, 5'd22, 27'h0000025f, 5'd5, 27'h0000027a, 32'h00000400,
  1'd1,  5'd29, 27'h0000000b, 5'd23, 27'h00000238, 5'd19, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000258, 5'd20, 27'h0000030e, 5'd26, 27'h000000ed, 32'h00000400,
  1'd1,  5'd8, 27'h000002ab, 5'd5, 27'h0000010a, 5'd3, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000332, 5'd5, 27'h000003f8, 5'd13, 27'h000001d1, 32'h00000400,
  1'd1,  5'd8, 27'h00000272, 5'd8, 27'h00000138, 5'd25, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000d9, 5'd17, 27'h00000008, 5'd1, 27'h0000026f, 32'h00000400,
  1'd1,  5'd6, 27'h000000a8, 5'd16, 27'h0000037d, 5'd14, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000015c, 5'd17, 27'h000001a2, 5'd25, 27'h00000188, 32'h00000400,
  1'd1,  5'd9, 27'h000000ef, 5'd29, 27'h00000034, 5'd4, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000371, 5'd29, 27'h000002f2, 5'd13, 27'h000002e6, 32'h00000400,
  1'd1,  5'd6, 27'h0000030e, 5'd25, 27'h000003dc, 5'd25, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032e, 5'd8, 27'h00000197, 5'd1, 27'h00000234, 32'h00000400,
  1'd1,  5'd16, 27'h00000185, 5'd7, 27'h000002ad, 5'd13, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000109, 5'd6, 27'h0000027b, 5'd20, 27'h000002e4, 32'h00000400,
  1'd1,  5'd19, 27'h0000016e, 5'd16, 27'h000001b6, 5'd3, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000222, 5'd16, 27'h00000283, 5'd14, 27'h0000018e, 32'h00000400,
  1'd1,  5'd19, 27'h00000018, 5'd18, 27'h00000033, 5'd22, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003c3, 5'd28, 27'h000002b7, 5'd2, 27'h0000003a, 32'h00000400,
  1'd1,  5'd16, 27'h00000251, 5'd27, 27'h00000277, 5'd14, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000326, 5'd26, 27'h000003cf, 5'd22, 27'h0000022c, 32'h00000400,
  1'd1,  5'd30, 27'h0000016a, 5'd5, 27'h0000015f, 5'd1, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003d0, 5'd10, 27'h000000df, 5'd13, 27'h00000198, 32'h00000400,
  1'd1,  5'd26, 27'h00000385, 5'd9, 27'h000001a1, 5'd21, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000015c, 5'd16, 27'h000003c5, 5'd3, 27'h000000bc, 32'h00000400,
  1'd1,  5'd30, 27'h00000118, 5'd17, 27'h0000016e, 5'd10, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000010e, 5'd19, 27'h0000032a, 5'd25, 27'h0000002c, 32'h00000400,
  1'd1,  5'd27, 27'h000001df, 5'd30, 27'h0000021e, 5'd4, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000331, 5'd28, 27'h0000033e, 5'd14, 27'h000002dd, 32'h00000400,
  1'd1,  5'd27, 27'h00000110, 5'd30, 27'h00000331, 5'd23, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003db, 5'd7, 27'h00000206, 5'd6, 27'h00000063, 32'h00000400,
  1'd1,  5'd7, 27'h0000024e, 5'd6, 27'h000003a9, 5'd19, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000031f, 5'd5, 27'h0000037a, 5'd29, 27'h000002c2, 32'h00000400,
  1'd1,  5'd7, 27'h0000009e, 5'd18, 27'h00000173, 5'd10, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000364, 5'd17, 27'h0000014a, 5'd19, 27'h00000132, 32'h00000400,
  1'd1,  5'd6, 27'h0000004a, 5'd17, 27'h00000297, 5'd26, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000150, 5'd28, 27'h00000234, 5'd5, 27'h0000030f, 32'h00000400,
  1'd1,  5'd6, 27'h000001e1, 5'd27, 27'h000001af, 5'd20, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001db, 5'd30, 27'h000002e9, 5'd26, 27'h000000b3, 32'h00000400,
  1'd1,  5'd17, 27'h0000014e, 5'd7, 27'h000002cd, 5'd6, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000194, 5'd7, 27'h0000027e, 5'd18, 27'h00000309, 32'h00000400,
  1'd1,  5'd19, 27'h000003a4, 5'd7, 27'h000001db, 5'd30, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002fb, 5'd19, 27'h00000209, 5'd9, 27'h0000014e, 32'h00000400,
  1'd1,  5'd16, 27'h0000026d, 5'd16, 27'h00000271, 5'd19, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000035, 5'd17, 27'h00000309, 5'd25, 27'h00000357, 32'h00000400,
  1'd1,  5'd17, 27'h00000233, 5'd29, 27'h000001ee, 5'd7, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000097, 5'd30, 27'h0000025f, 5'd20, 27'h0000008b, 32'h00000400,
  1'd1,  5'd18, 27'h0000035b, 5'd29, 27'h000003d2, 5'd30, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000087, 5'd5, 27'h00000145, 5'd5, 27'h0000016e, 32'h00000400,
  1'd1,  5'd28, 27'h0000007a, 5'd8, 27'h000000a0, 5'd20, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000025d, 5'd6, 27'h00000294, 5'd26, 27'h0000004b, 32'h00000400,
  1'd1,  5'd27, 27'h00000146, 5'd18, 27'h00000055, 5'd6, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000374, 5'd16, 27'h0000005b, 5'd18, 27'h000001b7, 32'h00000400,
  1'd1,  5'd26, 27'h00000173, 5'd17, 27'h000002e0, 5'd27, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002b6, 5'd27, 27'h00000003, 5'd8, 27'h0000019d, 32'h00000400,
  1'd1,  5'd30, 27'h000001a8, 5'd26, 27'h00000141, 5'd17, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000f7, 5'd28, 27'h00000343, 5'd27, 27'h00000206, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000000df, 5'd3, 27'h00000068, 5'd2, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003e8, 5'd3, 27'h000002b8, 5'd15, 27'h000000da, 32'h00000400,
  1'd1,  5'd1, 27'h00000290, 5'd0, 27'h0000016f, 5'd24, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b7, 5'd11, 27'h00000395, 5'd5, 27'h00000013, 32'h00000400,
  1'd1,  5'd0, 27'h000001fe, 5'd13, 27'h000003e7, 5'd12, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000393, 5'd13, 27'h000003e7, 5'd24, 27'h000003d9, 32'h00000400,
  1'd1,  5'd5, 27'h00000096, 5'd21, 27'h00000047, 5'd4, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000342, 5'd20, 27'h00000320, 5'd14, 27'h000000d6, 32'h00000400,
  1'd1,  5'd1, 27'h000000df, 5'd23, 27'h00000352, 5'd24, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000167, 5'd0, 27'h00000125, 5'd3, 27'h000002c0, 32'h00000400,
  1'd1,  5'd10, 27'h000002b3, 5'd0, 27'h000001d5, 5'd15, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f2, 5'd1, 27'h000001fb, 5'd23, 27'h00000018, 32'h00000400,
  1'd1,  5'd11, 27'h000000c4, 5'd12, 27'h0000024d, 5'd1, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000111, 5'd10, 27'h0000036f, 5'd14, 27'h0000009a, 32'h00000400,
  1'd1,  5'd11, 27'h00000095, 5'd13, 27'h0000016c, 5'd25, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b2, 5'd23, 27'h0000014f, 5'd4, 27'h000000f0, 32'h00000400,
  1'd1,  5'd12, 27'h000003b1, 5'd24, 27'h000002df, 5'd13, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000089, 5'd20, 27'h0000033a, 5'd24, 27'h000003bc, 32'h00000400,
  1'd1,  5'd23, 27'h0000033a, 5'd3, 27'h0000006a, 5'd3, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000360, 5'd1, 27'h00000070, 5'd13, 27'h000003df, 32'h00000400,
  1'd1,  5'd22, 27'h00000018, 5'd0, 27'h000001b0, 5'd21, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000269, 5'd13, 27'h000000a4, 5'd1, 27'h000000dc, 32'h00000400,
  1'd1,  5'd23, 27'h00000234, 5'd10, 27'h000003f2, 5'd12, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000127, 5'd14, 27'h00000011, 5'd23, 27'h0000008e, 32'h00000400,
  1'd1,  5'd21, 27'h00000083, 5'd23, 27'h00000286, 5'd3, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002be, 5'd25, 27'h000000ae, 5'd11, 27'h00000351, 32'h00000400,
  1'd1,  5'd22, 27'h0000028c, 5'd23, 27'h000001d2, 5'd22, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000033, 5'd2, 27'h0000017c, 5'd6, 27'h00000169, 32'h00000400,
  1'd1,  5'd2, 27'h00000133, 5'd0, 27'h000002d7, 5'd15, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000d7, 5'd1, 27'h000001ae, 5'd26, 27'h000001f0, 32'h00000400,
  1'd1,  5'd0, 27'h00000058, 5'd12, 27'h000001de, 5'd9, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d6, 5'd10, 27'h000001b9, 5'd19, 27'h00000336, 32'h00000400,
  1'd1,  5'd3, 27'h00000369, 5'd15, 27'h00000025, 5'd30, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001cd, 5'd24, 27'h000002a7, 5'd8, 27'h000003e8, 32'h00000400,
  1'd1,  5'd1, 27'h00000379, 5'd22, 27'h000000ae, 5'd18, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b4, 5'd21, 27'h00000259, 5'd27, 27'h00000159, 32'h00000400,
  1'd1,  5'd15, 27'h0000001b, 5'd3, 27'h000000a2, 5'd10, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000028f, 5'd0, 27'h000002e5, 5'd16, 27'h0000037a, 32'h00000400,
  1'd1,  5'd11, 27'h000000b0, 5'd4, 27'h000000df, 5'd26, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000077, 5'd12, 27'h00000388, 5'd7, 27'h000003ae, 32'h00000400,
  1'd1,  5'd14, 27'h000002fd, 5'd12, 27'h0000005b, 5'd15, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f9, 5'd15, 27'h000001f5, 5'd30, 27'h000003ba, 32'h00000400,
  1'd1,  5'd11, 27'h000001e4, 5'd23, 27'h000003e6, 5'd9, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003cf, 5'd21, 27'h000001d7, 5'd19, 27'h0000030c, 32'h00000400,
  1'd1,  5'd14, 27'h000001b1, 5'd24, 27'h00000293, 5'd26, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000002c, 5'd3, 27'h000000c7, 5'd9, 27'h00000388, 32'h00000400,
  1'd1,  5'd23, 27'h000001bb, 5'd4, 27'h000003c0, 5'd18, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000308, 5'd4, 27'h000002c8, 5'd28, 27'h000001eb, 32'h00000400,
  1'd1,  5'd24, 27'h000003a1, 5'd13, 27'h0000026a, 5'd7, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002fc, 5'd14, 27'h000002a3, 5'd16, 27'h000001a1, 32'h00000400,
  1'd1,  5'd25, 27'h000000fd, 5'd14, 27'h00000029, 5'd26, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000068, 5'd21, 27'h000002d0, 5'd8, 27'h000003d8, 32'h00000400,
  1'd1,  5'd24, 27'h0000020d, 5'd22, 27'h000003a6, 5'd17, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000153, 5'd24, 27'h00000053, 5'd27, 27'h0000034e, 32'h00000400,
  1'd1,  5'd3, 27'h000003be, 5'd7, 27'h00000181, 5'd4, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000041, 5'd5, 27'h000002e9, 5'd15, 27'h0000017b, 32'h00000400,
  1'd1,  5'd0, 27'h000003e7, 5'd8, 27'h00000130, 5'd21, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000af, 5'd18, 27'h000001e7, 5'd1, 27'h000000df, 32'h00000400,
  1'd1,  5'd1, 27'h000003cb, 5'd19, 27'h000002f3, 5'd13, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000020f, 5'd17, 27'h0000000b, 5'd21, 27'h00000245, 32'h00000400,
  1'd1,  5'd3, 27'h00000375, 5'd30, 27'h00000279, 5'd4, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000f9, 5'd29, 27'h00000075, 5'd12, 27'h0000013e, 32'h00000400,
  1'd1,  5'd0, 27'h000003bb, 5'd27, 27'h000001a2, 5'd24, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000028e, 5'd6, 27'h000000e1, 5'd4, 27'h00000090, 32'h00000400,
  1'd1,  5'd13, 27'h00000116, 5'd9, 27'h00000101, 5'd14, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000fd, 5'd5, 27'h00000377, 5'd24, 27'h00000232, 32'h00000400,
  1'd1,  5'd14, 27'h0000015c, 5'd19, 27'h0000002c, 5'd0, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c4, 5'd20, 27'h00000076, 5'd13, 27'h00000175, 32'h00000400,
  1'd1,  5'd11, 27'h000000eb, 5'd16, 27'h000002e2, 5'd22, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000296, 5'd28, 27'h00000365, 5'd4, 27'h000003ca, 32'h00000400,
  1'd1,  5'd12, 27'h0000016b, 5'd26, 27'h000002f3, 5'd12, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000172, 5'd29, 27'h0000031d, 5'd20, 27'h000003ba, 32'h00000400,
  1'd1,  5'd20, 27'h000003f5, 5'd9, 27'h000002cb, 5'd2, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000176, 5'd9, 27'h00000390, 5'd10, 27'h00000313, 32'h00000400,
  1'd1,  5'd22, 27'h000003a8, 5'd5, 27'h000001a3, 5'd24, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000355, 5'd15, 27'h0000038e, 5'd1, 27'h000000ad, 32'h00000400,
  1'd1,  5'd25, 27'h000000cc, 5'd17, 27'h000000fd, 5'd14, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000388, 5'd16, 27'h000001e9, 5'd20, 27'h000003b7, 32'h00000400,
  1'd1,  5'd23, 27'h00000156, 5'd28, 27'h0000006b, 5'd1, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002a8, 5'd26, 27'h00000200, 5'd10, 27'h00000246, 32'h00000400,
  1'd1,  5'd24, 27'h000000fc, 5'd27, 27'h00000102, 5'd23, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000342, 5'd6, 27'h000002f0, 5'd9, 27'h000002c2, 32'h00000400,
  1'd1,  5'd3, 27'h000002c2, 5'd9, 27'h0000026d, 5'd18, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000361, 5'd9, 27'h0000006c, 5'd25, 27'h0000039d, 32'h00000400,
  1'd1,  5'd3, 27'h00000214, 5'd17, 27'h0000000d, 5'd7, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000069, 5'd17, 27'h0000022a, 5'd19, 27'h0000036c, 32'h00000400,
  1'd1,  5'd3, 27'h00000234, 5'd18, 27'h000003c5, 5'd30, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000377, 5'd27, 27'h000000aa, 5'd6, 27'h000001ab, 32'h00000400,
  1'd1,  5'd3, 27'h00000316, 5'd28, 27'h000000b1, 5'd17, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d2, 5'd30, 27'h00000252, 5'd29, 27'h00000393, 32'h00000400,
  1'd1,  5'd14, 27'h00000243, 5'd8, 27'h00000296, 5'd8, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000351, 5'd8, 27'h00000253, 5'd19, 27'h0000034f, 32'h00000400,
  1'd1,  5'd11, 27'h00000253, 5'd7, 27'h000003fd, 5'd29, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f9, 5'd18, 27'h00000187, 5'd6, 27'h000003b7, 32'h00000400,
  1'd1,  5'd14, 27'h00000202, 5'd17, 27'h000001db, 5'd19, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000201, 5'd17, 27'h0000031a, 5'd25, 27'h00000369, 32'h00000400,
  1'd1,  5'd12, 27'h0000029e, 5'd26, 27'h00000083, 5'd9, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000259, 5'd30, 27'h00000009, 5'd19, 27'h0000030e, 32'h00000400,
  1'd1,  5'd11, 27'h000000d8, 5'd27, 27'h0000023d, 5'd30, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000342, 5'd6, 27'h00000189, 5'd8, 27'h0000020b, 32'h00000400,
  1'd1,  5'd22, 27'h00000326, 5'd7, 27'h00000248, 5'd16, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003d6, 5'd8, 27'h00000362, 5'd26, 27'h00000018, 32'h00000400,
  1'd1,  5'd23, 27'h00000268, 5'd19, 27'h000001db, 5'd8, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001e0, 5'd19, 27'h0000006d, 5'd20, 27'h000001e9, 32'h00000400,
  1'd1,  5'd21, 27'h00000139, 5'd16, 27'h00000319, 5'd30, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ad, 5'd30, 27'h000003f1, 5'd9, 27'h00000318, 32'h00000400,
  1'd1,  5'd22, 27'h000003fd, 5'd29, 27'h00000297, 5'd18, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000022b, 5'd28, 27'h0000038d, 5'd26, 27'h0000038f, 32'h00000400,
  1'd1,  5'd7, 27'h000000c5, 5'd1, 27'h000003eb, 5'd6, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000008, 5'd4, 27'h00000035, 5'd19, 27'h00000154, 32'h00000400,
  1'd1,  5'd8, 27'h000001b4, 5'd4, 27'h00000189, 5'd29, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a6, 5'd14, 27'h0000013e, 5'd4, 27'h0000016c, 32'h00000400,
  1'd1,  5'd8, 27'h00000021, 5'd13, 27'h000003b7, 5'd10, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000130, 5'd12, 27'h0000018c, 5'd22, 27'h00000295, 32'h00000400,
  1'd1,  5'd7, 27'h000001ed, 5'd24, 27'h00000243, 5'd3, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000007d, 5'd20, 27'h000002cb, 5'd11, 27'h00000249, 32'h00000400,
  1'd1,  5'd10, 27'h00000074, 5'd25, 27'h00000118, 5'd20, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000005f, 5'd1, 27'h000003d4, 5'd6, 27'h00000134, 32'h00000400,
  1'd1,  5'd19, 27'h0000013d, 5'd0, 27'h00000230, 5'd18, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002a4, 5'd3, 27'h000001fd, 5'd30, 27'h000002e1, 32'h00000400,
  1'd1,  5'd15, 27'h0000022d, 5'd11, 27'h00000009, 5'd2, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000130, 5'd13, 27'h000001e5, 5'd13, 27'h00000249, 32'h00000400,
  1'd1,  5'd17, 27'h0000016a, 5'd11, 27'h00000397, 5'd22, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000325, 5'd22, 27'h000000b7, 5'd1, 27'h0000012d, 32'h00000400,
  1'd1,  5'd16, 27'h0000037b, 5'd20, 27'h00000363, 5'd11, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000247, 5'd21, 27'h00000336, 5'd21, 27'h00000240, 32'h00000400,
  1'd1,  5'd26, 27'h000002d0, 5'd4, 27'h00000200, 5'd3, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000246, 5'd1, 27'h000003e3, 5'd12, 27'h000000ee, 32'h00000400,
  1'd1,  5'd26, 27'h00000337, 5'd2, 27'h00000280, 5'd23, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e6, 5'd12, 27'h000000e7, 5'd2, 27'h000001dc, 32'h00000400,
  1'd1,  5'd29, 27'h0000004b, 5'd11, 27'h00000285, 5'd14, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003c8, 5'd14, 27'h000000d9, 5'd21, 27'h000003f9, 32'h00000400,
  1'd1,  5'd29, 27'h000001c1, 5'd22, 27'h000000bb, 5'd2, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036c, 5'd24, 27'h000002f5, 5'd11, 27'h000001b7, 32'h00000400,
  1'd1,  5'd27, 27'h000001e0, 5'd23, 27'h00000356, 5'd22, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003b8, 5'd5, 27'h00000041, 5'd3, 27'h0000025a, 32'h00000400,
  1'd1,  5'd9, 27'h000001f6, 5'd0, 27'h00000351, 5'd14, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000009e, 5'd5, 27'h0000007a, 5'd22, 27'h000000f6, 32'h00000400,
  1'd1,  5'd7, 27'h0000011c, 5'd15, 27'h00000094, 5'd7, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000064, 5'd13, 27'h0000033a, 5'd17, 27'h000002e0, 32'h00000400,
  1'd1,  5'd9, 27'h0000025f, 5'd13, 27'h00000336, 5'd25, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020f, 5'd24, 27'h00000357, 5'd9, 27'h00000197, 32'h00000400,
  1'd1,  5'd10, 27'h00000078, 5'd25, 27'h0000016b, 5'd20, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b0, 5'd23, 27'h000001f2, 5'd29, 27'h000000af, 32'h00000400,
  1'd1,  5'd16, 27'h00000057, 5'd3, 27'h000002b4, 5'd3, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000018b, 5'd2, 27'h0000021d, 5'd12, 27'h000000b0, 32'h00000400,
  1'd1,  5'd19, 27'h000000b1, 5'd2, 27'h000000ed, 5'd21, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000238, 5'd14, 27'h000003ca, 5'd9, 27'h0000013d, 32'h00000400,
  1'd1,  5'd18, 27'h000001a8, 5'd12, 27'h00000160, 5'd16, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000236, 5'd14, 27'h000001c2, 5'd29, 27'h00000328, 32'h00000400,
  1'd1,  5'd19, 27'h00000127, 5'd25, 27'h00000180, 5'd6, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000030f, 5'd20, 27'h000002c2, 5'd19, 27'h000003ab, 32'h00000400,
  1'd1,  5'd15, 27'h000003cd, 5'd23, 27'h00000380, 5'd26, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000272, 5'd4, 27'h00000174, 5'd8, 27'h0000003f, 32'h00000400,
  1'd1,  5'd27, 27'h000002d7, 5'd0, 27'h0000037f, 5'd20, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000367, 5'd1, 27'h00000118, 5'd27, 27'h00000102, 32'h00000400,
  1'd1,  5'd27, 27'h000002e3, 5'd14, 27'h0000005e, 5'd5, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c9, 5'd10, 27'h00000355, 5'd19, 27'h000001d3, 32'h00000400,
  1'd1,  5'd27, 27'h000000ef, 5'd14, 27'h0000002e, 5'd26, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000e6, 5'd21, 27'h00000287, 5'd5, 27'h00000203, 32'h00000400,
  1'd1,  5'd26, 27'h000001d9, 5'd22, 27'h0000011f, 5'd19, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000009a, 5'd21, 27'h000000fc, 5'd28, 27'h000001c5, 32'h00000400,
  1'd1,  5'd7, 27'h0000020b, 5'd6, 27'h0000002b, 5'd4, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023e, 5'd6, 27'h00000147, 5'd14, 27'h000003dd, 32'h00000400,
  1'd1,  5'd7, 27'h0000032f, 5'd9, 27'h0000006a, 5'd23, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000182, 5'd17, 27'h0000029f, 5'd0, 27'h00000094, 32'h00000400,
  1'd1,  5'd5, 27'h000001b5, 5'd20, 27'h00000061, 5'd11, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000038f, 5'd20, 27'h0000020b, 5'd23, 27'h0000033d, 32'h00000400,
  1'd1,  5'd9, 27'h00000198, 5'd30, 27'h00000080, 5'd1, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000304, 5'd30, 27'h00000341, 5'd13, 27'h0000000b, 32'h00000400,
  1'd1,  5'd9, 27'h000000c8, 5'd26, 27'h0000018a, 5'd25, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000019f, 5'd6, 27'h00000287, 5'd3, 27'h0000002d, 32'h00000400,
  1'd1,  5'd17, 27'h000001d5, 5'd8, 27'h000003fc, 5'd14, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a0, 5'd6, 27'h00000332, 5'd23, 27'h0000025e, 32'h00000400,
  1'd1,  5'd17, 27'h0000038d, 5'd17, 27'h000002dd, 5'd2, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002f4, 5'd18, 27'h0000005b, 5'd14, 27'h00000211, 32'h00000400,
  1'd1,  5'd16, 27'h00000112, 5'd16, 27'h000001ba, 5'd24, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000020f, 5'd27, 27'h000003ec, 5'd1, 27'h000003c4, 32'h00000400,
  1'd1,  5'd17, 27'h000001ed, 5'd27, 27'h000002b0, 5'd12, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000246, 5'd30, 27'h00000338, 5'd25, 27'h00000264, 32'h00000400,
  1'd1,  5'd26, 27'h000002d6, 5'd9, 27'h00000374, 5'd0, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000268, 5'd9, 27'h000000c0, 5'd14, 27'h000003f7, 32'h00000400,
  1'd1,  5'd29, 27'h00000028, 5'd7, 27'h00000198, 5'd21, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000013d, 5'd17, 27'h0000005c, 5'd3, 27'h00000042, 32'h00000400,
  1'd1,  5'd29, 27'h00000201, 5'd16, 27'h0000036a, 5'd12, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000028, 5'd20, 27'h00000250, 5'd24, 27'h00000273, 32'h00000400,
  1'd1,  5'd26, 27'h0000032e, 5'd28, 27'h0000038b, 5'd2, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000033c, 5'd26, 27'h000003c9, 5'd10, 27'h00000214, 32'h00000400,
  1'd1,  5'd27, 27'h0000032a, 5'd26, 27'h0000023f, 5'd22, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c7, 5'd8, 27'h00000083, 5'd9, 27'h000003d9, 32'h00000400,
  1'd1,  5'd9, 27'h00000005, 5'd6, 27'h00000064, 5'd16, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000211, 5'd8, 27'h000000f5, 5'd27, 27'h00000057, 32'h00000400,
  1'd1,  5'd8, 27'h00000164, 5'd17, 27'h00000225, 5'd9, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000154, 5'd16, 27'h000003c7, 5'd17, 27'h0000010b, 32'h00000400,
  1'd1,  5'd8, 27'h0000014f, 5'd16, 27'h0000011c, 5'd30, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013a, 5'd27, 27'h000003be, 5'd5, 27'h0000025f, 32'h00000400,
  1'd1,  5'd7, 27'h00000269, 5'd29, 27'h00000110, 5'd19, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000026d, 5'd28, 27'h00000233, 5'd26, 27'h00000089, 32'h00000400,
  1'd1,  5'd20, 27'h00000085, 5'd7, 27'h00000160, 5'd9, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000207, 5'd6, 27'h000003f8, 5'd18, 27'h000003f1, 32'h00000400,
  1'd1,  5'd15, 27'h0000035f, 5'd7, 27'h000000ca, 5'd26, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000083, 5'd16, 27'h00000279, 5'd6, 27'h00000096, 32'h00000400,
  1'd1,  5'd16, 27'h000002fc, 5'd18, 27'h00000377, 5'd18, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002fe, 5'd16, 27'h000003cc, 5'd26, 27'h000002e6, 32'h00000400,
  1'd1,  5'd18, 27'h00000014, 5'd26, 27'h0000017a, 5'd5, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000032, 5'd30, 27'h00000343, 5'd17, 27'h00000047, 32'h00000400,
  1'd1,  5'd20, 27'h00000274, 5'd27, 27'h00000337, 5'd30, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002e7, 5'd6, 27'h0000033f, 5'd6, 27'h00000037, 32'h00000400,
  1'd1,  5'd29, 27'h0000032b, 5'd9, 27'h0000010d, 5'd15, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000022e, 5'd9, 27'h0000036d, 5'd26, 27'h0000022b, 32'h00000400,
  1'd1,  5'd28, 27'h000000c5, 5'd16, 27'h00000203, 5'd8, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000028c, 5'd19, 27'h000003ed, 5'd18, 27'h00000246, 32'h00000400,
  1'd1,  5'd26, 27'h000001d5, 5'd17, 27'h000003a4, 5'd29, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003cd, 5'd27, 27'h000003d1, 5'd9, 27'h00000099, 32'h00000400,
  1'd1,  5'd28, 27'h0000015a, 5'd26, 27'h00000319, 5'd20, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000292, 5'd26, 27'h0000038d, 5'd28, 27'h000000b3, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000005c, 5'd4, 27'h0000006f, 5'd3, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023a, 5'd1, 27'h000001e4, 5'd13, 27'h0000005f, 32'h00000400,
  1'd1,  5'd1, 27'h000000c1, 5'd3, 27'h00000001, 5'd20, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d1, 5'd13, 27'h0000024e, 5'd3, 27'h00000099, 32'h00000400,
  1'd1,  5'd4, 27'h000001ee, 5'd13, 27'h000001f0, 5'd13, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000088, 5'd10, 27'h00000283, 5'd21, 27'h000003d9, 32'h00000400,
  1'd1,  5'd0, 27'h00000292, 5'd23, 27'h000000f0, 5'd4, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000013f, 5'd23, 27'h00000222, 5'd14, 27'h0000020f, 32'h00000400,
  1'd1,  5'd1, 27'h00000054, 5'd23, 27'h000003bd, 5'd20, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000206, 5'd4, 27'h00000339, 5'd3, 27'h000001fa, 32'h00000400,
  1'd1,  5'd15, 27'h000001d2, 5'd1, 27'h0000001c, 5'd10, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000337, 5'd3, 27'h0000033e, 5'd24, 27'h00000310, 32'h00000400,
  1'd1,  5'd14, 27'h000003d2, 5'd14, 27'h00000147, 5'd3, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000000a, 5'd10, 27'h000002d3, 5'd13, 27'h0000027a, 32'h00000400,
  1'd1,  5'd13, 27'h000003a7, 5'd14, 27'h00000067, 5'd25, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ff, 5'd25, 27'h0000005e, 5'd5, 27'h00000073, 32'h00000400,
  1'd1,  5'd12, 27'h000001b8, 5'd22, 27'h00000074, 5'd13, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020d, 5'd21, 27'h0000038b, 5'd24, 27'h000000e9, 32'h00000400,
  1'd1,  5'd25, 27'h000000bc, 5'd1, 27'h000001d0, 5'd2, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000366, 5'd4, 27'h00000101, 5'd11, 27'h000001ee, 32'h00000400,
  1'd1,  5'd23, 27'h000002c6, 5'd2, 27'h00000381, 5'd25, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000006d, 5'd11, 27'h000000a1, 5'd3, 27'h000002c1, 32'h00000400,
  1'd1,  5'd21, 27'h00000042, 5'd13, 27'h00000235, 5'd11, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000046, 5'd10, 27'h0000036a, 5'd22, 27'h00000195, 32'h00000400,
  1'd1,  5'd22, 27'h000003e3, 5'd23, 27'h000003fa, 5'd3, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003cb, 5'd20, 27'h00000325, 5'd15, 27'h0000001f, 32'h00000400,
  1'd1,  5'd24, 27'h0000006c, 5'd25, 27'h0000009f, 5'd24, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000370, 5'd3, 27'h0000021b, 5'd7, 27'h00000259, 32'h00000400,
  1'd1,  5'd1, 27'h00000067, 5'd0, 27'h0000025e, 5'd18, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000150, 5'd1, 27'h00000075, 5'd25, 27'h0000039a, 32'h00000400,
  1'd1,  5'd3, 27'h00000160, 5'd14, 27'h000002c0, 5'd6, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000000a, 5'd15, 27'h000001d8, 5'd19, 27'h0000011a, 32'h00000400,
  1'd1,  5'd2, 27'h000003b3, 5'd12, 27'h00000324, 5'd29, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ce, 5'd23, 27'h000003ab, 5'd6, 27'h00000253, 32'h00000400,
  1'd1,  5'd0, 27'h0000039c, 5'd22, 27'h000001c2, 5'd17, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000379, 5'd20, 27'h0000037a, 5'd29, 27'h00000169, 32'h00000400,
  1'd1,  5'd10, 27'h000002f2, 5'd1, 27'h0000009c, 5'd6, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a6, 5'd2, 27'h00000252, 5'd18, 27'h000000e9, 32'h00000400,
  1'd1,  5'd13, 27'h000002b7, 5'd3, 27'h00000006, 5'd30, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011c, 5'd10, 27'h000002dd, 5'd7, 27'h0000033d, 32'h00000400,
  1'd1,  5'd13, 27'h000001cf, 5'd15, 27'h00000183, 5'd17, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000311, 5'd10, 27'h0000017b, 5'd29, 27'h0000016a, 32'h00000400,
  1'd1,  5'd12, 27'h000002c4, 5'd22, 27'h00000355, 5'd7, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c8, 5'd21, 27'h000002b0, 5'd18, 27'h000002d4, 32'h00000400,
  1'd1,  5'd15, 27'h000001a8, 5'd23, 27'h0000036f, 5'd26, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002f3, 5'd5, 27'h00000001, 5'd9, 27'h00000399, 32'h00000400,
  1'd1,  5'd21, 27'h0000005f, 5'd0, 27'h00000116, 5'd16, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003dd, 5'd1, 27'h0000024f, 5'd27, 27'h00000196, 32'h00000400,
  1'd1,  5'd24, 27'h000000bd, 5'd13, 27'h00000072, 5'd5, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002cd, 5'd14, 27'h000001df, 5'd20, 27'h0000014f, 32'h00000400,
  1'd1,  5'd23, 27'h000001e7, 5'd12, 27'h00000149, 5'd29, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ff, 5'd21, 27'h0000022f, 5'd8, 27'h00000260, 32'h00000400,
  1'd1,  5'd21, 27'h000001b5, 5'd24, 27'h0000007f, 5'd18, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000142, 5'd25, 27'h00000221, 5'd28, 27'h00000193, 32'h00000400,
  1'd1,  5'd4, 27'h00000354, 5'd8, 27'h00000280, 5'd0, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000087, 5'd5, 27'h000003b5, 5'd12, 27'h000000dc, 32'h00000400,
  1'd1,  5'd1, 27'h00000323, 5'd10, 27'h00000077, 5'd23, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000080, 5'd20, 27'h00000274, 5'd3, 27'h00000234, 32'h00000400,
  1'd1,  5'd2, 27'h00000262, 5'd18, 27'h0000007b, 5'd13, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000016e, 5'd18, 27'h000003a4, 5'd22, 27'h00000258, 32'h00000400,
  1'd1,  5'd4, 27'h00000373, 5'd30, 27'h0000031a, 5'd0, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023a, 5'd30, 27'h0000001c, 5'd11, 27'h00000143, 32'h00000400,
  1'd1,  5'd4, 27'h0000026e, 5'd30, 27'h0000036f, 5'd23, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000075, 5'd5, 27'h00000121, 5'd2, 27'h00000293, 32'h00000400,
  1'd1,  5'd12, 27'h00000287, 5'd6, 27'h000000fb, 5'd12, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001f4, 5'd7, 27'h000001e0, 5'd21, 27'h00000095, 32'h00000400,
  1'd1,  5'd11, 27'h0000001d, 5'd17, 27'h0000036e, 5'd3, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ba, 5'd15, 27'h000003cf, 5'd12, 27'h000001ce, 32'h00000400,
  1'd1,  5'd10, 27'h00000195, 5'd17, 27'h0000015e, 5'd22, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000ee, 5'd30, 27'h0000036a, 5'd3, 27'h0000026c, 32'h00000400,
  1'd1,  5'd11, 27'h000000c6, 5'd26, 27'h000000d2, 5'd13, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000335, 5'd28, 27'h0000031a, 5'd22, 27'h00000181, 32'h00000400,
  1'd1,  5'd24, 27'h00000014, 5'd7, 27'h000000a3, 5'd4, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000276, 5'd6, 27'h00000122, 5'd11, 27'h0000024b, 32'h00000400,
  1'd1,  5'd25, 27'h0000001a, 5'd5, 27'h0000012c, 5'd22, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b0, 5'd20, 27'h00000183, 5'd2, 27'h000002f3, 32'h00000400,
  1'd1,  5'd21, 27'h000003e8, 5'd16, 27'h00000219, 5'd12, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000302, 5'd17, 27'h0000017e, 5'd23, 27'h0000006d, 32'h00000400,
  1'd1,  5'd25, 27'h000001a6, 5'd28, 27'h0000015f, 5'd2, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b2, 5'd28, 27'h00000289, 5'd12, 27'h00000247, 32'h00000400,
  1'd1,  5'd23, 27'h00000103, 5'd27, 27'h0000028f, 5'd24, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ad, 5'd7, 27'h000003e3, 5'd6, 27'h000003d7, 32'h00000400,
  1'd1,  5'd1, 27'h0000017e, 5'd7, 27'h00000120, 5'd17, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000022, 5'd9, 27'h000003f1, 5'd29, 27'h00000099, 32'h00000400,
  1'd1,  5'd3, 27'h000000f2, 5'd19, 27'h000001e5, 5'd5, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000102, 5'd17, 27'h000001d8, 5'd18, 27'h0000037f, 32'h00000400,
  1'd1,  5'd3, 27'h00000379, 5'd15, 27'h000002cf, 5'd28, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003be, 5'd28, 27'h0000020a, 5'd7, 27'h00000259, 32'h00000400,
  1'd1,  5'd2, 27'h0000029e, 5'd29, 27'h00000264, 5'd19, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ce, 5'd27, 27'h0000016d, 5'd25, 27'h000003df, 32'h00000400,
  1'd1,  5'd13, 27'h000000be, 5'd6, 27'h000003c6, 5'd6, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000371, 5'd9, 27'h00000244, 5'd19, 27'h000000ff, 32'h00000400,
  1'd1,  5'd10, 27'h0000031e, 5'd9, 27'h000003b0, 5'd26, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000239, 5'd18, 27'h000002d7, 5'd9, 27'h000000d4, 32'h00000400,
  1'd1,  5'd11, 27'h00000193, 5'd19, 27'h00000387, 5'd18, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e0, 5'd18, 27'h00000022, 5'd27, 27'h0000002e, 32'h00000400,
  1'd1,  5'd11, 27'h00000105, 5'd27, 27'h00000313, 5'd8, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001db, 5'd26, 27'h00000265, 5'd19, 27'h00000386, 32'h00000400,
  1'd1,  5'd10, 27'h000001cd, 5'd26, 27'h00000105, 5'd30, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000029, 5'd7, 27'h00000358, 5'd8, 27'h000002a5, 32'h00000400,
  1'd1,  5'd25, 27'h00000051, 5'd6, 27'h0000015a, 5'd16, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000252, 5'd6, 27'h000001ef, 5'd26, 27'h00000167, 32'h00000400,
  1'd1,  5'd23, 27'h00000278, 5'd16, 27'h00000103, 5'd9, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000048, 5'd18, 27'h000002cd, 5'd17, 27'h0000006a, 32'h00000400,
  1'd1,  5'd24, 27'h000003fa, 5'd17, 27'h0000031f, 5'd27, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034d, 5'd30, 27'h000003a8, 5'd10, 27'h0000012e, 32'h00000400,
  1'd1,  5'd23, 27'h00000149, 5'd29, 27'h0000016f, 5'd17, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000006b, 5'd26, 27'h0000006a, 5'd27, 27'h000000ed, 32'h00000400,
  1'd1,  5'd8, 27'h000002e5, 5'd0, 27'h00000383, 5'd7, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000129, 5'd4, 27'h0000010c, 5'd18, 27'h00000080, 32'h00000400,
  1'd1,  5'd7, 27'h000002ef, 5'd2, 27'h00000183, 5'd26, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000dc, 5'd13, 27'h000001b4, 5'd1, 27'h000003a1, 32'h00000400,
  1'd1,  5'd7, 27'h00000000, 5'd11, 27'h0000005d, 5'd14, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000154, 5'd12, 27'h00000313, 5'd21, 27'h00000118, 32'h00000400,
  1'd1,  5'd9, 27'h00000099, 5'd21, 27'h000003be, 5'd0, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000368, 5'd24, 27'h000002fa, 5'd12, 27'h0000039f, 32'h00000400,
  1'd1,  5'd8, 27'h000003d9, 5'd22, 27'h00000009, 5'd23, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000011a, 5'd2, 27'h000000b0, 5'd9, 27'h000001b3, 32'h00000400,
  1'd1,  5'd20, 27'h000001b8, 5'd2, 27'h00000305, 5'd15, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000008d, 5'd0, 27'h00000137, 5'd26, 27'h000003e9, 32'h00000400,
  1'd1,  5'd19, 27'h000001a2, 5'd14, 27'h000003cf, 5'd3, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000008d, 5'd10, 27'h0000017f, 5'd10, 27'h000001f1, 32'h00000400,
  1'd1,  5'd20, 27'h000001a8, 5'd11, 27'h0000028a, 5'd20, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001fe, 5'd22, 27'h00000003, 5'd3, 27'h00000060, 32'h00000400,
  1'd1,  5'd19, 27'h000003b1, 5'd23, 27'h0000009e, 5'd10, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000009a, 5'd20, 27'h0000030d, 5'd20, 27'h000002c7, 32'h00000400,
  1'd1,  5'd25, 27'h0000037d, 5'd3, 27'h00000250, 5'd2, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000dd, 5'd2, 27'h000001e1, 5'd12, 27'h0000039f, 32'h00000400,
  1'd1,  5'd27, 27'h000000f3, 5'd4, 27'h00000266, 5'd21, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000026e, 5'd15, 27'h00000105, 5'd4, 27'h0000033b, 32'h00000400,
  1'd1,  5'd30, 27'h000002bc, 5'd11, 27'h0000036f, 5'd12, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000024c, 5'd12, 27'h000002b9, 5'd21, 27'h000000c5, 32'h00000400,
  1'd1,  5'd30, 27'h00000363, 5'd22, 27'h000001e4, 5'd3, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000207, 5'd22, 27'h000000a3, 5'd14, 27'h0000038b, 32'h00000400,
  1'd1,  5'd29, 27'h00000095, 5'd20, 27'h00000333, 5'd22, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001f8, 5'd0, 27'h000003d3, 5'd0, 27'h00000158, 32'h00000400,
  1'd1,  5'd9, 27'h00000312, 5'd3, 27'h00000282, 5'd11, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000377, 5'd1, 27'h00000110, 5'd20, 27'h00000380, 32'h00000400,
  1'd1,  5'd8, 27'h00000022, 5'd11, 27'h00000259, 5'd5, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000215, 5'd11, 27'h000002ae, 5'd16, 27'h000000d3, 32'h00000400,
  1'd1,  5'd8, 27'h00000378, 5'd13, 27'h0000032d, 5'd26, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000030f, 5'd22, 27'h000001bb, 5'd6, 27'h00000296, 32'h00000400,
  1'd1,  5'd9, 27'h00000073, 5'd23, 27'h00000222, 5'd19, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ee, 5'd25, 27'h000000ea, 5'd27, 27'h00000180, 32'h00000400,
  1'd1,  5'd20, 27'h00000256, 5'd2, 27'h00000044, 5'd2, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ac, 5'd4, 27'h000003bb, 5'd12, 27'h0000001c, 32'h00000400,
  1'd1,  5'd19, 27'h000000f9, 5'd4, 27'h000000c8, 5'd24, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000e2, 5'd14, 27'h000002d7, 5'd5, 27'h000003b7, 32'h00000400,
  1'd1,  5'd18, 27'h0000002c, 5'd12, 27'h0000003a, 5'd15, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d6, 5'd12, 27'h000003b5, 5'd27, 27'h000003a2, 32'h00000400,
  1'd1,  5'd19, 27'h000002be, 5'd25, 27'h00000052, 5'd8, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000366, 5'd22, 27'h000002e2, 5'd19, 27'h000002db, 32'h00000400,
  1'd1,  5'd19, 27'h00000394, 5'd25, 27'h00000289, 5'd28, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000389, 5'd2, 27'h000003b2, 5'd5, 27'h0000034d, 32'h00000400,
  1'd1,  5'd29, 27'h00000138, 5'd2, 27'h000002a4, 5'd16, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000030d, 5'd1, 27'h000000bd, 5'd27, 27'h00000272, 32'h00000400,
  1'd1,  5'd27, 27'h00000357, 5'd11, 27'h00000052, 5'd6, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003da, 5'd12, 27'h000000cd, 5'd19, 27'h00000048, 32'h00000400,
  1'd1,  5'd27, 27'h00000209, 5'd10, 27'h000001a3, 5'd26, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000133, 5'd25, 27'h0000029a, 5'd9, 27'h0000003e, 32'h00000400,
  1'd1,  5'd28, 27'h000000bd, 5'd23, 27'h0000038d, 5'd17, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000336, 5'd22, 27'h0000022b, 5'd30, 27'h000002e1, 32'h00000400,
  1'd1,  5'd10, 27'h000000c2, 5'd7, 27'h000003f5, 5'd3, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003af, 5'd10, 27'h0000001e, 5'd11, 27'h00000244, 32'h00000400,
  1'd1,  5'd6, 27'h000002de, 5'd10, 27'h000000db, 5'd23, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e7, 5'd15, 27'h0000028d, 5'd0, 27'h00000011, 32'h00000400,
  1'd1,  5'd5, 27'h00000339, 5'd16, 27'h000003ff, 5'd15, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000d6, 5'd16, 27'h000001f4, 5'd21, 27'h00000151, 32'h00000400,
  1'd1,  5'd9, 27'h00000085, 5'd27, 27'h00000331, 5'd2, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000003, 5'd30, 27'h0000023c, 5'd12, 27'h00000172, 32'h00000400,
  1'd1,  5'd9, 27'h0000028a, 5'd27, 27'h00000148, 5'd20, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000012f, 5'd6, 27'h00000362, 5'd4, 27'h000003bf, 32'h00000400,
  1'd1,  5'd20, 27'h000001a5, 5'd9, 27'h00000163, 5'd13, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003f4, 5'd8, 27'h000003df, 5'd23, 27'h000001b0, 32'h00000400,
  1'd1,  5'd16, 27'h000002a1, 5'd17, 27'h000003b1, 5'd3, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000253, 5'd15, 27'h0000030f, 5'd14, 27'h00000243, 32'h00000400,
  1'd1,  5'd19, 27'h00000148, 5'd20, 27'h00000012, 5'd22, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ea, 5'd28, 27'h00000385, 5'd0, 27'h000002b5, 32'h00000400,
  1'd1,  5'd16, 27'h00000194, 5'd29, 27'h0000030a, 5'd11, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003a6, 5'd27, 27'h000002f3, 5'd23, 27'h0000030d, 32'h00000400,
  1'd1,  5'd30, 27'h00000273, 5'd9, 27'h0000035a, 5'd1, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000173, 5'd9, 27'h00000273, 5'd13, 27'h0000018c, 32'h00000400,
  1'd1,  5'd28, 27'h0000038c, 5'd6, 27'h00000125, 5'd23, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ea, 5'd19, 27'h000000fa, 5'd3, 27'h00000362, 32'h00000400,
  1'd1,  5'd27, 27'h00000349, 5'd18, 27'h0000038b, 5'd12, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001e0, 5'd19, 27'h00000286, 5'd22, 27'h00000086, 32'h00000400,
  1'd1,  5'd29, 27'h00000386, 5'd28, 27'h0000001c, 5'd0, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000078, 5'd30, 27'h000002bc, 5'd12, 27'h0000032d, 32'h00000400,
  1'd1,  5'd25, 27'h000003b9, 5'd27, 27'h000003a7, 5'd24, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000c2, 5'd8, 27'h00000161, 5'd6, 27'h000003dd, 32'h00000400,
  1'd1,  5'd10, 27'h000000c2, 5'd6, 27'h00000322, 5'd16, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000231, 5'd9, 27'h000002fd, 5'd30, 27'h000002dd, 32'h00000400,
  1'd1,  5'd6, 27'h000000fc, 5'd17, 27'h0000025c, 5'd9, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003dd, 5'd19, 27'h00000078, 5'd20, 27'h00000136, 32'h00000400,
  1'd1,  5'd7, 27'h00000131, 5'd19, 27'h000000e2, 5'd26, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000178, 5'd28, 27'h000000fa, 5'd10, 27'h00000089, 32'h00000400,
  1'd1,  5'd7, 27'h00000296, 5'd28, 27'h0000016c, 5'd19, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000112, 5'd28, 27'h000000cd, 5'd27, 27'h000002c4, 32'h00000400,
  1'd1,  5'd17, 27'h000002e7, 5'd9, 27'h00000337, 5'd8, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000104, 5'd8, 27'h00000282, 5'd18, 27'h00000259, 32'h00000400,
  1'd1,  5'd19, 27'h00000063, 5'd10, 27'h0000005c, 5'd26, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000019f, 5'd18, 27'h000002f9, 5'd5, 27'h0000025c, 32'h00000400,
  1'd1,  5'd19, 27'h000000c6, 5'd15, 27'h000003b6, 5'd16, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ef, 5'd16, 27'h00000015, 5'd29, 27'h0000026a, 32'h00000400,
  1'd1,  5'd20, 27'h00000181, 5'd28, 27'h000003a9, 5'd7, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a9, 5'd29, 27'h00000398, 5'd19, 27'h000001b7, 32'h00000400,
  1'd1,  5'd16, 27'h00000191, 5'd28, 27'h000001b2, 5'd28, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000037e, 5'd9, 27'h000002d7, 5'd8, 27'h000001cf, 32'h00000400,
  1'd1,  5'd28, 27'h00000371, 5'd7, 27'h0000024f, 5'd19, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006a, 5'd7, 27'h00000086, 5'd28, 27'h000001da, 32'h00000400,
  1'd1,  5'd29, 27'h000000e7, 5'd18, 27'h00000003, 5'd8, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000c4, 5'd20, 27'h0000010c, 5'd15, 27'h000003c8, 32'h00000400,
  1'd1,  5'd30, 27'h0000020f, 5'd19, 27'h000003c8, 5'd27, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d6, 5'd30, 27'h00000342, 5'd6, 27'h00000197, 32'h00000400,
  1'd1,  5'd29, 27'h00000012, 5'd27, 27'h00000198, 5'd18, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000036e, 5'd26, 27'h000000fd, 5'd29, 27'h00000250, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000205, 5'd4, 27'h00000073, 5'd1, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000207, 5'd2, 27'h000001f8, 5'd11, 27'h00000013, 32'h00000400,
  1'd1,  5'd4, 27'h000000de, 5'd2, 27'h0000012e, 5'd24, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000394, 5'd15, 27'h00000032, 5'd1, 27'h00000115, 32'h00000400,
  1'd1,  5'd1, 27'h000002e6, 5'd14, 27'h0000034d, 5'd13, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000363, 5'd11, 27'h0000006b, 5'd23, 27'h000002db, 32'h00000400,
  1'd1,  5'd2, 27'h000000bd, 5'd23, 27'h000003cd, 5'd1, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a4, 5'd21, 27'h000002c4, 5'd11, 27'h000003ea, 32'h00000400,
  1'd1,  5'd0, 27'h000003a4, 5'd22, 27'h00000271, 5'd21, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002c9, 5'd4, 27'h0000038b, 5'd1, 27'h000003db, 32'h00000400,
  1'd1,  5'd14, 27'h000003da, 5'd0, 27'h0000036e, 5'd12, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003ab, 5'd0, 27'h00000375, 5'd23, 27'h0000021b, 32'h00000400,
  1'd1,  5'd10, 27'h00000225, 5'd13, 27'h000001a1, 5'd5, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000179, 5'd12, 27'h0000038f, 5'd14, 27'h000002f1, 32'h00000400,
  1'd1,  5'd11, 27'h00000063, 5'd12, 27'h000002aa, 5'd21, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000355, 5'd21, 27'h000000bc, 5'd1, 27'h00000048, 32'h00000400,
  1'd1,  5'd10, 27'h00000208, 5'd21, 27'h0000014f, 5'd15, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ec, 5'd21, 27'h000000c9, 5'd22, 27'h00000149, 32'h00000400,
  1'd1,  5'd23, 27'h00000302, 5'd2, 27'h000002a8, 5'd4, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000002f, 5'd4, 27'h00000200, 5'd15, 27'h0000013d, 32'h00000400,
  1'd1,  5'd21, 27'h000001f3, 5'd5, 27'h00000044, 5'd21, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000011c, 5'd10, 27'h00000287, 5'd4, 27'h00000315, 32'h00000400,
  1'd1,  5'd21, 27'h000001ec, 5'd10, 27'h000001e9, 5'd11, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000355, 5'd10, 27'h00000273, 5'd23, 27'h0000009e, 32'h00000400,
  1'd1,  5'd25, 27'h00000099, 5'd25, 27'h000001c0, 5'd4, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000327, 5'd25, 27'h000001d6, 5'd14, 27'h00000311, 32'h00000400,
  1'd1,  5'd23, 27'h000001b4, 5'd23, 27'h000000b2, 5'd22, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000012e, 5'd0, 27'h000000ce, 5'd10, 27'h0000003d, 32'h00000400,
  1'd1,  5'd4, 27'h00000136, 5'd1, 27'h00000395, 5'd18, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000331, 5'd2, 27'h000000a0, 5'd26, 27'h00000273, 32'h00000400,
  1'd1,  5'd0, 27'h0000010e, 5'd15, 27'h00000135, 5'd9, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b7, 5'd11, 27'h000000bd, 5'd16, 27'h000000f7, 32'h00000400,
  1'd1,  5'd1, 27'h000003bb, 5'd11, 27'h000002ca, 5'd26, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003e8, 5'd24, 27'h0000033f, 5'd6, 27'h00000046, 32'h00000400,
  1'd1,  5'd3, 27'h0000028e, 5'd24, 27'h0000010b, 5'd16, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000153, 5'd24, 27'h000002c3, 5'd27, 27'h00000310, 32'h00000400,
  1'd1,  5'd10, 27'h00000358, 5'd0, 27'h0000024c, 5'd9, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018a, 5'd0, 27'h0000005b, 5'd16, 27'h00000042, 32'h00000400,
  1'd1,  5'd11, 27'h00000140, 5'd3, 27'h000003f2, 5'd30, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003a7, 5'd10, 27'h00000248, 5'd10, 27'h0000007b, 32'h00000400,
  1'd1,  5'd11, 27'h00000342, 5'd10, 27'h00000307, 5'd20, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a6, 5'd12, 27'h00000053, 5'd26, 27'h00000061, 32'h00000400,
  1'd1,  5'd10, 27'h000001a3, 5'd25, 27'h000000d3, 5'd8, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000028a, 5'd24, 27'h00000098, 5'd16, 27'h00000154, 32'h00000400,
  1'd1,  5'd13, 27'h000001a5, 5'd23, 27'h000002af, 5'd27, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001d9, 5'd0, 27'h00000105, 5'd5, 27'h0000019c, 32'h00000400,
  1'd1,  5'd21, 27'h0000023b, 5'd5, 27'h00000062, 5'd16, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001f0, 5'd1, 27'h000002f6, 5'd29, 27'h000002f0, 32'h00000400,
  1'd1,  5'd24, 27'h0000029c, 5'd14, 27'h00000008, 5'd7, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000003c, 5'd10, 27'h00000374, 5'd17, 27'h00000069, 32'h00000400,
  1'd1,  5'd22, 27'h00000206, 5'd11, 27'h00000141, 5'd29, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000007b, 5'd25, 27'h000000cc, 5'd6, 27'h000003bc, 32'h00000400,
  1'd1,  5'd24, 27'h000001c4, 5'd23, 27'h00000098, 5'd18, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000074, 5'd24, 27'h00000235, 5'd28, 27'h00000328, 32'h00000400,
  1'd1,  5'd3, 27'h000001c2, 5'd6, 27'h000003ea, 5'd1, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002b2, 5'd8, 27'h00000005, 5'd13, 27'h000000c2, 32'h00000400,
  1'd1,  5'd2, 27'h0000015f, 5'd8, 27'h0000012b, 5'd25, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f6, 5'd17, 27'h000000e7, 5'd4, 27'h000000f7, 32'h00000400,
  1'd1,  5'd0, 27'h000001ed, 5'd18, 27'h00000367, 5'd15, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001de, 5'd19, 27'h00000304, 5'd24, 27'h000002fa, 32'h00000400,
  1'd1,  5'd4, 27'h00000126, 5'd30, 27'h000000ba, 5'd1, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000264, 5'd30, 27'h000003e1, 5'd11, 27'h00000151, 32'h00000400,
  1'd1,  5'd2, 27'h0000021e, 5'd28, 27'h0000007e, 5'd23, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c7, 5'd9, 27'h00000240, 5'd2, 27'h000003af, 32'h00000400,
  1'd1,  5'd14, 27'h0000005d, 5'd8, 27'h000003d7, 5'd13, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000269, 5'd7, 27'h000000d7, 5'd24, 27'h000003a7, 32'h00000400,
  1'd1,  5'd10, 27'h000003b0, 5'd16, 27'h00000324, 5'd0, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000003d, 5'd15, 27'h000002eb, 5'd15, 27'h00000184, 32'h00000400,
  1'd1,  5'd15, 27'h00000165, 5'd17, 27'h000002d3, 5'd21, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f5, 5'd29, 27'h00000182, 5'd5, 27'h00000099, 32'h00000400,
  1'd1,  5'd15, 27'h000001b0, 5'd29, 27'h00000188, 5'd13, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000325, 5'd26, 27'h00000231, 5'd22, 27'h00000263, 32'h00000400,
  1'd1,  5'd20, 27'h000002ac, 5'd6, 27'h0000014b, 5'd4, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000232, 5'd9, 27'h00000366, 5'd14, 27'h0000035b, 32'h00000400,
  1'd1,  5'd25, 27'h00000215, 5'd8, 27'h00000295, 5'd21, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000006d, 5'd16, 27'h000001df, 5'd1, 27'h0000001e, 32'h00000400,
  1'd1,  5'd24, 27'h00000031, 5'd17, 27'h0000035f, 5'd12, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000125, 5'd16, 27'h000002d7, 5'd21, 27'h000001bd, 32'h00000400,
  1'd1,  5'd23, 27'h00000229, 5'd26, 27'h000002f4, 5'd3, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003f5, 5'd29, 27'h000002f0, 5'd12, 27'h0000025a, 32'h00000400,
  1'd1,  5'd24, 27'h0000013b, 5'd28, 27'h00000109, 5'd22, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000105, 5'd9, 27'h000001c0, 5'd9, 27'h000002aa, 32'h00000400,
  1'd1,  5'd2, 27'h000003b6, 5'd5, 27'h0000017c, 5'd20, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000186, 5'd9, 27'h000003dd, 5'd26, 27'h0000003f, 32'h00000400,
  1'd1,  5'd2, 27'h000000b6, 5'd18, 27'h00000147, 5'd5, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000019c, 5'd19, 27'h0000029c, 5'd15, 27'h00000351, 32'h00000400,
  1'd1,  5'd2, 27'h0000015c, 5'd18, 27'h00000317, 5'd26, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001f8, 5'd27, 27'h00000280, 5'd7, 27'h00000155, 32'h00000400,
  1'd1,  5'd1, 27'h00000354, 5'd30, 27'h000001e4, 5'd17, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000008c, 5'd28, 27'h000002f1, 5'd29, 27'h000001c9, 32'h00000400,
  1'd1,  5'd12, 27'h000003f2, 5'd5, 27'h000000bd, 5'd8, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000342, 5'd9, 27'h00000209, 5'd17, 27'h0000023f, 32'h00000400,
  1'd1,  5'd14, 27'h00000364, 5'd8, 27'h000002f2, 5'd28, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e6, 5'd15, 27'h00000393, 5'd7, 27'h00000110, 32'h00000400,
  1'd1,  5'd14, 27'h00000044, 5'd16, 27'h00000296, 5'd16, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000011d, 5'd19, 27'h000000d7, 5'd30, 27'h00000226, 32'h00000400,
  1'd1,  5'd10, 27'h0000031c, 5'd28, 27'h00000374, 5'd9, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000391, 5'd27, 27'h000001ad, 5'd17, 27'h000003c2, 32'h00000400,
  1'd1,  5'd14, 27'h00000115, 5'd26, 27'h0000004d, 5'd26, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000031f, 5'd8, 27'h00000143, 5'd9, 27'h00000335, 32'h00000400,
  1'd1,  5'd24, 27'h000001c4, 5'd5, 27'h000001ed, 5'd17, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001d5, 5'd6, 27'h0000032b, 5'd29, 27'h0000004a, 32'h00000400,
  1'd1,  5'd23, 27'h00000308, 5'd20, 27'h00000272, 5'd7, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000f0, 5'd19, 27'h00000185, 5'd18, 27'h00000383, 32'h00000400,
  1'd1,  5'd23, 27'h00000320, 5'd18, 27'h00000107, 5'd26, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000282, 5'd27, 27'h0000034d, 5'd9, 27'h0000033d, 32'h00000400,
  1'd1,  5'd20, 27'h000002c0, 5'd27, 27'h000003bb, 5'd18, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b8, 5'd30, 27'h00000178, 5'd29, 27'h000002b4, 32'h00000400,
  1'd1,  5'd7, 27'h0000018f, 5'd4, 27'h000000d2, 5'd6, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d4, 5'd3, 27'h000003df, 5'd15, 27'h0000033e, 32'h00000400,
  1'd1,  5'd6, 27'h00000214, 5'd0, 27'h00000300, 5'd30, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ff, 5'd14, 27'h00000234, 5'd5, 27'h00000009, 32'h00000400,
  1'd1,  5'd6, 27'h00000277, 5'd14, 27'h00000139, 5'd10, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d4, 5'd14, 27'h000001e8, 5'd24, 27'h0000027a, 32'h00000400,
  1'd1,  5'd8, 27'h000000b1, 5'd23, 27'h000003bc, 5'd0, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e2, 5'd22, 27'h00000199, 5'd13, 27'h000000a1, 32'h00000400,
  1'd1,  5'd5, 27'h000002a4, 5'd25, 27'h000002b1, 5'd22, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000035, 5'd0, 27'h00000087, 5'd7, 27'h00000226, 32'h00000400,
  1'd1,  5'd17, 27'h000002c2, 5'd3, 27'h000000bb, 5'd20, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000030f, 5'd0, 27'h0000030b, 5'd27, 27'h00000233, 32'h00000400,
  1'd1,  5'd16, 27'h0000033d, 5'd10, 27'h00000370, 5'd0, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000001a, 5'd13, 27'h000001b8, 5'd13, 27'h000003b0, 32'h00000400,
  1'd1,  5'd16, 27'h0000034b, 5'd14, 27'h000001d1, 5'd23, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a0, 5'd25, 27'h0000029f, 5'd0, 27'h00000330, 32'h00000400,
  1'd1,  5'd16, 27'h00000077, 5'd25, 27'h00000138, 5'd11, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000211, 5'd20, 27'h0000038c, 5'd21, 27'h000002c6, 32'h00000400,
  1'd1,  5'd26, 27'h00000358, 5'd3, 27'h000002b1, 5'd3, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000056, 5'd4, 27'h0000039c, 5'd12, 27'h000002ec, 32'h00000400,
  1'd1,  5'd30, 27'h00000298, 5'd1, 27'h000001fc, 5'd21, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003a6, 5'd12, 27'h0000001e, 5'd4, 27'h00000176, 32'h00000400,
  1'd1,  5'd27, 27'h00000194, 5'd13, 27'h00000127, 5'd11, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000080, 5'd15, 27'h0000018b, 5'd24, 27'h00000333, 32'h00000400,
  1'd1,  5'd26, 27'h000002db, 5'd24, 27'h000003ed, 5'd3, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000367, 5'd20, 27'h00000327, 5'd14, 27'h000003c9, 32'h00000400,
  1'd1,  5'd30, 27'h000001b5, 5'd21, 27'h000000c0, 5'd25, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000028c, 5'd1, 27'h000003fe, 5'd3, 27'h000001fe, 32'h00000400,
  1'd1,  5'd8, 27'h0000034a, 5'd4, 27'h000001d6, 5'd15, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f7, 5'd4, 27'h00000236, 5'd21, 27'h00000074, 32'h00000400,
  1'd1,  5'd5, 27'h0000029e, 5'd10, 27'h000003ff, 5'd7, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000367, 5'd13, 27'h000002b6, 5'd15, 27'h000003b1, 32'h00000400,
  1'd1,  5'd9, 27'h000001a5, 5'd13, 27'h000002f0, 5'd28, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000038b, 5'd23, 27'h000000b1, 5'd5, 27'h000003c9, 32'h00000400,
  1'd1,  5'd8, 27'h00000071, 5'd24, 27'h00000285, 5'd19, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000247, 5'd23, 27'h0000024a, 5'd28, 27'h0000001c, 32'h00000400,
  1'd1,  5'd16, 27'h0000000b, 5'd4, 27'h000000b7, 5'd1, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000038d, 5'd1, 27'h0000015b, 5'd12, 27'h000003bd, 32'h00000400,
  1'd1,  5'd17, 27'h00000181, 5'd4, 27'h000000de, 5'd25, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001a0, 5'd14, 27'h000000ea, 5'd5, 27'h00000108, 32'h00000400,
  1'd1,  5'd19, 27'h00000217, 5'd13, 27'h00000258, 5'd19, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002d7, 5'd11, 27'h0000006e, 5'd29, 27'h0000020d, 32'h00000400,
  1'd1,  5'd15, 27'h000002fb, 5'd20, 27'h0000038d, 5'd8, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000171, 5'd24, 27'h000002d7, 5'd16, 27'h000000db, 32'h00000400,
  1'd1,  5'd17, 27'h0000025a, 5'd24, 27'h0000009f, 5'd26, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003e4, 5'd3, 27'h000003b9, 5'd8, 27'h000003c0, 32'h00000400,
  1'd1,  5'd28, 27'h0000027b, 5'd3, 27'h00000025, 5'd20, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001e2, 5'd3, 27'h000003ea, 5'd27, 27'h000003fe, 32'h00000400,
  1'd1,  5'd25, 27'h00000369, 5'd11, 27'h000003e5, 5'd5, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002e2, 5'd12, 27'h0000015f, 5'd16, 27'h00000340, 32'h00000400,
  1'd1,  5'd29, 27'h0000028b, 5'd10, 27'h000001bd, 5'd28, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000eb, 5'd23, 27'h0000027b, 5'd5, 27'h0000032f, 32'h00000400,
  1'd1,  5'd30, 27'h0000014c, 5'd20, 27'h00000369, 5'd20, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000f8, 5'd23, 27'h000003a3, 5'd28, 27'h0000004d, 32'h00000400,
  1'd1,  5'd5, 27'h00000178, 5'd10, 27'h00000014, 5'd2, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009e, 5'd6, 27'h0000025a, 5'd10, 27'h000002e9, 32'h00000400,
  1'd1,  5'd7, 27'h00000069, 5'd8, 27'h00000379, 5'd22, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003be, 5'd15, 27'h0000033c, 5'd0, 27'h00000264, 32'h00000400,
  1'd1,  5'd5, 27'h000000e5, 5'd19, 27'h000002e7, 5'd15, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000038b, 5'd16, 27'h0000032a, 5'd24, 27'h000003fa, 32'h00000400,
  1'd1,  5'd7, 27'h000002ea, 5'd28, 27'h00000231, 5'd4, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000166, 5'd27, 27'h0000000d, 5'd12, 27'h00000057, 32'h00000400,
  1'd1,  5'd8, 27'h000001d0, 5'd27, 27'h000002c4, 5'd21, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f6, 5'd7, 27'h000002a1, 5'd1, 27'h000001b2, 32'h00000400,
  1'd1,  5'd16, 27'h000003ab, 5'd5, 27'h0000022f, 5'd14, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000176, 5'd10, 27'h00000003, 5'd22, 27'h000001e5, 32'h00000400,
  1'd1,  5'd19, 27'h00000390, 5'd15, 27'h00000358, 5'd2, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000367, 5'd15, 27'h00000275, 5'd12, 27'h0000024a, 32'h00000400,
  1'd1,  5'd17, 27'h000001af, 5'd17, 27'h000000ba, 5'd21, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000185, 5'd28, 27'h000002f5, 5'd1, 27'h00000256, 32'h00000400,
  1'd1,  5'd18, 27'h0000013e, 5'd30, 27'h0000038d, 5'd12, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003bb, 5'd29, 27'h000000e9, 5'd24, 27'h0000012b, 32'h00000400,
  1'd1,  5'd30, 27'h000000ac, 5'd8, 27'h0000031b, 5'd4, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000095, 5'd8, 27'h000001c9, 5'd11, 27'h000001d6, 32'h00000400,
  1'd1,  5'd27, 27'h000003fc, 5'd6, 27'h000003f3, 5'd21, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000030a, 5'd17, 27'h0000001e, 5'd0, 27'h000002e0, 32'h00000400,
  1'd1,  5'd25, 27'h000003f9, 5'd18, 27'h00000122, 5'd15, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002bb, 5'd16, 27'h000003bf, 5'd24, 27'h0000024c, 32'h00000400,
  1'd1,  5'd25, 27'h000003b0, 5'd27, 27'h00000041, 5'd4, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000bb, 5'd27, 27'h000001db, 5'd12, 27'h0000002a, 32'h00000400,
  1'd1,  5'd26, 27'h00000087, 5'd26, 27'h000003c2, 5'd23, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000121, 5'd8, 27'h00000211, 5'd5, 27'h00000276, 32'h00000400,
  1'd1,  5'd7, 27'h00000068, 5'd10, 27'h0000014f, 5'd18, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000309, 5'd9, 27'h00000147, 5'd27, 27'h00000351, 32'h00000400,
  1'd1,  5'd5, 27'h00000171, 5'd17, 27'h00000039, 5'd5, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000026d, 5'd16, 27'h00000261, 5'd15, 27'h000003d1, 32'h00000400,
  1'd1,  5'd8, 27'h00000147, 5'd18, 27'h00000143, 5'd28, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002f8, 5'd27, 27'h0000031e, 5'd6, 27'h000003d3, 32'h00000400,
  1'd1,  5'd6, 27'h000001a3, 5'd29, 27'h00000240, 5'd20, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000303, 5'd26, 27'h000002d5, 5'd30, 27'h000001b5, 32'h00000400,
  1'd1,  5'd19, 27'h0000037c, 5'd6, 27'h0000017c, 5'd8, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000225, 5'd5, 27'h000002d6, 5'd17, 27'h00000397, 32'h00000400,
  1'd1,  5'd18, 27'h000003ca, 5'd9, 27'h0000023b, 5'd27, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a5, 5'd16, 27'h00000209, 5'd8, 27'h000000eb, 32'h00000400,
  1'd1,  5'd19, 27'h00000160, 5'd19, 27'h00000038, 5'd19, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000174, 5'd17, 27'h000001fb, 5'd29, 27'h00000024, 32'h00000400,
  1'd1,  5'd17, 27'h0000031f, 5'd30, 27'h0000027f, 5'd6, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000108, 5'd28, 27'h00000396, 5'd17, 27'h000000f9, 32'h00000400,
  1'd1,  5'd19, 27'h000001dd, 5'd29, 27'h000002a4, 5'd26, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000035a, 5'd5, 27'h00000102, 5'd7, 27'h00000089, 32'h00000400,
  1'd1,  5'd26, 27'h0000035a, 5'd9, 27'h000002e5, 5'd17, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001e7, 5'd7, 27'h000002b1, 5'd30, 27'h000001b9, 32'h00000400,
  1'd1,  5'd30, 27'h000003e7, 5'd17, 27'h00000232, 5'd8, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000366, 5'd19, 27'h0000010b, 5'd18, 27'h000002b1, 32'h00000400,
  1'd1,  5'd27, 27'h000001e1, 5'd16, 27'h00000102, 5'd26, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000311, 5'd25, 27'h000003c4, 5'd10, 27'h00000014, 32'h00000400,
  1'd1,  5'd30, 27'h000003d1, 5'd28, 27'h000003fc, 5'd18, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000fa, 5'd28, 27'h00000271, 5'd27, 27'h0000017e, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000088, 5'd4, 27'h000000bb, 5'd1, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000224, 5'd3, 27'h000000e2, 5'd14, 27'h00000320, 32'h00000400,
  1'd1,  5'd3, 27'h000002c7, 5'd3, 27'h00000026, 5'd24, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000f3, 5'd14, 27'h000002dc, 5'd0, 27'h000003a0, 32'h00000400,
  1'd1,  5'd0, 27'h000002a7, 5'd12, 27'h000003cf, 5'd14, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000244, 5'd14, 27'h000001d3, 5'd21, 27'h000001f0, 32'h00000400,
  1'd1,  5'd4, 27'h00000097, 5'd21, 27'h0000030b, 5'd4, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000111, 5'd20, 27'h000002ff, 5'd10, 27'h00000378, 32'h00000400,
  1'd1,  5'd5, 27'h00000049, 5'd21, 27'h00000344, 5'd25, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029d, 5'd0, 27'h000001b4, 5'd4, 27'h0000000e, 32'h00000400,
  1'd1,  5'd12, 27'h0000013a, 5'd0, 27'h00000308, 5'd12, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000c1, 5'd2, 27'h000001c8, 5'd22, 27'h000003b8, 32'h00000400,
  1'd1,  5'd15, 27'h0000008f, 5'd14, 27'h0000016a, 5'd3, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009d, 5'd10, 27'h000002bb, 5'd12, 27'h0000026d, 32'h00000400,
  1'd1,  5'd13, 27'h000003b3, 5'd14, 27'h00000073, 5'd20, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000331, 5'd21, 27'h000002e5, 5'd3, 27'h000000ec, 32'h00000400,
  1'd1,  5'd12, 27'h0000018f, 5'd22, 27'h000001b0, 5'd13, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e9, 5'd24, 27'h000000fb, 5'd21, 27'h0000001e, 32'h00000400,
  1'd1,  5'd21, 27'h000002da, 5'd1, 27'h00000196, 5'd2, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000143, 5'd0, 27'h000003b3, 5'd11, 27'h0000020a, 32'h00000400,
  1'd1,  5'd25, 27'h00000173, 5'd2, 27'h00000382, 5'd22, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000036e, 5'd12, 27'h00000349, 5'd0, 27'h00000161, 32'h00000400,
  1'd1,  5'd21, 27'h0000028c, 5'd12, 27'h000000b8, 5'd15, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000022f, 5'd12, 27'h00000329, 5'd24, 27'h000002e4, 32'h00000400,
  1'd1,  5'd22, 27'h00000155, 5'd25, 27'h0000002b, 5'd3, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003c5, 5'd22, 27'h000003eb, 5'd13, 27'h000002f2, 32'h00000400,
  1'd1,  5'd22, 27'h000000e8, 5'd23, 27'h00000297, 5'd25, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001be, 5'd2, 27'h000001f0, 5'd9, 27'h0000036b, 32'h00000400,
  1'd1,  5'd5, 27'h00000047, 5'd4, 27'h00000400, 5'd17, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000327, 5'd3, 27'h00000310, 5'd30, 27'h00000069, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd11, 27'h000003e9, 5'd5, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d6, 5'd10, 27'h000002d9, 5'd19, 27'h000003f1, 32'h00000400,
  1'd1,  5'd4, 27'h00000374, 5'd14, 27'h00000280, 5'd26, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001e8, 5'd21, 27'h00000395, 5'd9, 27'h000003be, 32'h00000400,
  1'd1,  5'd3, 27'h00000172, 5'd20, 27'h000002c3, 5'd16, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c7, 5'd22, 27'h000000f5, 5'd27, 27'h000001aa, 32'h00000400,
  1'd1,  5'd13, 27'h0000035d, 5'd4, 27'h00000005, 5'd5, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001b3, 5'd1, 27'h0000008c, 5'd16, 27'h00000102, 32'h00000400,
  1'd1,  5'd12, 27'h00000293, 5'd3, 27'h000001a5, 5'd27, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a3, 5'd13, 27'h000003ab, 5'd6, 27'h000002ba, 32'h00000400,
  1'd1,  5'd14, 27'h00000062, 5'd13, 27'h000001da, 5'd19, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000024b, 5'd10, 27'h00000193, 5'd30, 27'h00000306, 32'h00000400,
  1'd1,  5'd11, 27'h00000177, 5'd22, 27'h00000031, 5'd6, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000197, 5'd23, 27'h00000027, 5'd18, 27'h000002b4, 32'h00000400,
  1'd1,  5'd10, 27'h00000185, 5'd21, 27'h00000164, 5'd27, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ae, 5'd2, 27'h000002b9, 5'd9, 27'h0000017c, 32'h00000400,
  1'd1,  5'd20, 27'h000002d2, 5'd0, 27'h000002dd, 5'd17, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000027e, 5'd1, 27'h0000011e, 5'd28, 27'h00000233, 32'h00000400,
  1'd1,  5'd21, 27'h00000061, 5'd11, 27'h0000016e, 5'd5, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001b8, 5'd14, 27'h000001e3, 5'd20, 27'h00000037, 32'h00000400,
  1'd1,  5'd24, 27'h0000038f, 5'd12, 27'h0000021f, 5'd26, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000271, 5'd23, 27'h0000033f, 5'd7, 27'h000003ec, 32'h00000400,
  1'd1,  5'd23, 27'h0000009c, 5'd25, 27'h000002bd, 5'd20, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000198, 5'd22, 27'h00000089, 5'd28, 27'h000002a4, 32'h00000400,
  1'd1,  5'd1, 27'h0000032f, 5'd9, 27'h000001d8, 5'd1, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000032, 5'd7, 27'h000001d3, 5'd14, 27'h000000ec, 32'h00000400,
  1'd1,  5'd4, 27'h00000032, 5'd10, 27'h00000102, 5'd24, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000028e, 5'd20, 27'h0000015d, 5'd2, 27'h0000012b, 32'h00000400,
  1'd1,  5'd1, 27'h000001ff, 5'd20, 27'h000001e2, 5'd13, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000030d, 5'd19, 27'h00000252, 5'd24, 27'h00000036, 32'h00000400,
  1'd1,  5'd3, 27'h0000005a, 5'd29, 27'h0000010f, 5'd0, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000359, 5'd29, 27'h000003d8, 5'd15, 27'h00000057, 32'h00000400,
  1'd1,  5'd0, 27'h00000187, 5'd27, 27'h000002ec, 5'd20, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000006b, 5'd6, 27'h000003f8, 5'd4, 27'h0000035e, 32'h00000400,
  1'd1,  5'd14, 27'h00000238, 5'd6, 27'h000002f2, 5'd13, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002dc, 5'd6, 27'h00000368, 5'd24, 27'h00000352, 32'h00000400,
  1'd1,  5'd14, 27'h00000154, 5'd18, 27'h0000018b, 5'd4, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ce, 5'd15, 27'h000003a7, 5'd10, 27'h00000334, 32'h00000400,
  1'd1,  5'd14, 27'h00000053, 5'd19, 27'h00000107, 5'd22, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000361, 5'd30, 27'h000003a1, 5'd3, 27'h000003fd, 32'h00000400,
  1'd1,  5'd11, 27'h00000052, 5'd29, 27'h0000019d, 5'd13, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000332, 5'd26, 27'h00000205, 5'd25, 27'h00000038, 32'h00000400,
  1'd1,  5'd24, 27'h00000310, 5'd6, 27'h00000122, 5'd4, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002fb, 5'd7, 27'h0000038c, 5'd11, 27'h00000307, 32'h00000400,
  1'd1,  5'd22, 27'h000002c7, 5'd9, 27'h000003da, 5'd23, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000035f, 5'd17, 27'h00000310, 5'd1, 27'h000001fe, 32'h00000400,
  1'd1,  5'd20, 27'h000003fd, 5'd20, 27'h00000120, 5'd13, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000278, 5'd19, 27'h00000262, 5'd25, 27'h0000020e, 32'h00000400,
  1'd1,  5'd21, 27'h0000022d, 5'd30, 27'h00000050, 5'd2, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000053, 5'd29, 27'h000003ee, 5'd12, 27'h0000022a, 32'h00000400,
  1'd1,  5'd24, 27'h00000247, 5'd27, 27'h000000dd, 5'd24, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000037, 5'd7, 27'h0000036e, 5'd10, 27'h00000119, 32'h00000400,
  1'd1,  5'd5, 27'h00000059, 5'd8, 27'h00000221, 5'd15, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002e3, 5'd8, 27'h00000174, 5'd30, 27'h000002eb, 32'h00000400,
  1'd1,  5'd4, 27'h000002a1, 5'd19, 27'h0000036e, 5'd7, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000096, 5'd19, 27'h0000002a, 5'd16, 27'h000000b1, 32'h00000400,
  1'd1,  5'd4, 27'h00000036, 5'd19, 27'h00000178, 5'd30, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000281, 5'd28, 27'h00000242, 5'd7, 27'h00000042, 32'h00000400,
  1'd1,  5'd1, 27'h00000024, 5'd30, 27'h0000015b, 5'd17, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000013a, 5'd30, 27'h00000123, 5'd28, 27'h00000124, 32'h00000400,
  1'd1,  5'd12, 27'h000001dd, 5'd8, 27'h00000325, 5'd8, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000395, 5'd7, 27'h00000280, 5'd18, 27'h000000c1, 32'h00000400,
  1'd1,  5'd10, 27'h00000389, 5'd6, 27'h000002b2, 5'd25, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ce, 5'd16, 27'h00000004, 5'd5, 27'h000000f5, 32'h00000400,
  1'd1,  5'd10, 27'h0000030c, 5'd16, 27'h00000016, 5'd19, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000015b, 5'd17, 27'h0000001d, 5'd30, 27'h00000132, 32'h00000400,
  1'd1,  5'd13, 27'h00000095, 5'd29, 27'h00000396, 5'd5, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ee, 5'd26, 27'h00000085, 5'd20, 27'h00000242, 32'h00000400,
  1'd1,  5'd13, 27'h000002a3, 5'd29, 27'h000001d6, 5'd26, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000120, 5'd6, 27'h0000011c, 5'd10, 27'h0000007f, 32'h00000400,
  1'd1,  5'd23, 27'h000000b1, 5'd8, 27'h000001a2, 5'd19, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b2, 5'd5, 27'h000003aa, 5'd29, 27'h00000301, 32'h00000400,
  1'd1,  5'd25, 27'h000000b1, 5'd17, 27'h000002a0, 5'd7, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000209, 5'd19, 27'h0000009a, 5'd17, 27'h000002b7, 32'h00000400,
  1'd1,  5'd25, 27'h000001ce, 5'd20, 27'h000000c9, 5'd27, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000013a, 5'd29, 27'h00000219, 5'd8, 27'h00000128, 32'h00000400,
  1'd1,  5'd23, 27'h00000148, 5'd30, 27'h000000a8, 5'd20, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000008b, 5'd28, 27'h0000006f, 5'd28, 27'h000000e6, 32'h00000400,
  1'd1,  5'd5, 27'h00000373, 5'd1, 27'h000000b3, 5'd7, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000026f, 5'd3, 27'h00000014, 5'd19, 27'h0000013d, 32'h00000400,
  1'd1,  5'd9, 27'h000002c3, 5'd2, 27'h0000013f, 5'd27, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000014a, 5'd11, 27'h000001b1, 5'd1, 27'h0000003d, 32'h00000400,
  1'd1,  5'd7, 27'h0000015f, 5'd11, 27'h000000ba, 5'd10, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000b1, 5'd12, 27'h00000054, 5'd24, 27'h000003d5, 32'h00000400,
  1'd1,  5'd6, 27'h0000027b, 5'd21, 27'h000003bb, 5'd5, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000077, 5'd23, 27'h000000ff, 5'd13, 27'h0000011e, 32'h00000400,
  1'd1,  5'd7, 27'h000003ff, 5'd24, 27'h00000184, 5'd24, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000353, 5'd1, 27'h00000196, 5'd5, 27'h00000232, 32'h00000400,
  1'd1,  5'd15, 27'h00000372, 5'd2, 27'h0000014b, 5'd18, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002aa, 5'd0, 27'h000003eb, 5'd27, 27'h00000280, 32'h00000400,
  1'd1,  5'd19, 27'h000000b9, 5'd12, 27'h000003bb, 5'd4, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001bf, 5'd13, 27'h00000069, 5'd14, 27'h00000055, 32'h00000400,
  1'd1,  5'd18, 27'h0000026d, 5'd11, 27'h000002b9, 5'd21, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001bc, 5'd24, 27'h000001e7, 5'd4, 27'h000001d0, 32'h00000400,
  1'd1,  5'd16, 27'h00000134, 5'd25, 27'h000001b1, 5'd13, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000bf, 5'd25, 27'h00000234, 5'd22, 27'h0000005c, 32'h00000400,
  1'd1,  5'd26, 27'h000000f8, 5'd2, 27'h0000030d, 5'd1, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000fc, 5'd4, 27'h000000c2, 5'd15, 27'h000000fb, 32'h00000400,
  1'd1,  5'd26, 27'h000002d7, 5'd3, 27'h00000157, 5'd24, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000074, 5'd12, 27'h00000073, 5'd2, 27'h0000035b, 32'h00000400,
  1'd1,  5'd27, 27'h0000032f, 5'd14, 27'h000003f3, 5'd11, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000103, 5'd13, 27'h0000034b, 5'd25, 27'h00000128, 32'h00000400,
  1'd1,  5'd30, 27'h00000339, 5'd24, 27'h000001e2, 5'd1, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000a9, 5'd22, 27'h00000045, 5'd12, 27'h00000370, 32'h00000400,
  1'd1,  5'd30, 27'h0000030a, 5'd21, 27'h000000af, 5'd21, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a6, 5'd1, 27'h000001d9, 5'd2, 27'h000001a0, 32'h00000400,
  1'd1,  5'd10, 27'h0000002b, 5'd0, 27'h00000196, 5'd13, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000025f, 5'd4, 27'h000001ac, 5'd23, 27'h0000002b, 32'h00000400,
  1'd1,  5'd5, 27'h0000010f, 5'd14, 27'h000000ca, 5'd6, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000013e, 5'd10, 27'h000001b9, 5'd18, 27'h00000396, 32'h00000400,
  1'd1,  5'd7, 27'h0000038a, 5'd11, 27'h000003cf, 5'd30, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d0, 5'd23, 27'h00000390, 5'd6, 27'h000002cf, 32'h00000400,
  1'd1,  5'd5, 27'h00000312, 5'd21, 27'h00000352, 5'd18, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000339, 5'd22, 27'h000003e8, 5'd26, 27'h000000ca, 32'h00000400,
  1'd1,  5'd18, 27'h0000012f, 5'd2, 27'h000003ae, 5'd4, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a8, 5'd4, 27'h000002fb, 5'd12, 27'h0000033d, 32'h00000400,
  1'd1,  5'd17, 27'h0000003f, 5'd0, 27'h00000269, 5'd24, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000080, 5'd15, 27'h000001b3, 5'd8, 27'h00000177, 32'h00000400,
  1'd1,  5'd15, 27'h0000023b, 5'd11, 27'h0000031c, 5'd18, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000212, 5'd15, 27'h000001f5, 5'd29, 27'h00000044, 32'h00000400,
  1'd1,  5'd16, 27'h0000013d, 5'd25, 27'h000001d1, 5'd7, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000038b, 5'd22, 27'h00000284, 5'd18, 27'h00000256, 32'h00000400,
  1'd1,  5'd18, 27'h000000be, 5'd23, 27'h00000057, 5'd26, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003ad, 5'd4, 27'h000002e9, 5'd6, 27'h000002d2, 32'h00000400,
  1'd1,  5'd30, 27'h00000093, 5'd2, 27'h000000e7, 5'd17, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001fa, 5'd2, 27'h00000070, 5'd28, 27'h00000317, 32'h00000400,
  1'd1,  5'd29, 27'h00000090, 5'd11, 27'h000001b0, 5'd6, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000083, 5'd13, 27'h000003c8, 5'd19, 27'h00000265, 32'h00000400,
  1'd1,  5'd27, 27'h0000039e, 5'd15, 27'h000000cb, 5'd27, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000351, 5'd21, 27'h00000318, 5'd7, 27'h00000073, 32'h00000400,
  1'd1,  5'd27, 27'h000001db, 5'd21, 27'h000001a8, 5'd19, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000025a, 5'd22, 27'h00000349, 5'd27, 27'h00000177, 32'h00000400,
  1'd1,  5'd6, 27'h00000203, 5'd5, 27'h000002fb, 5'd4, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000010e, 5'd6, 27'h000002b3, 5'd13, 27'h000002b6, 32'h00000400,
  1'd1,  5'd6, 27'h00000359, 5'd7, 27'h00000358, 5'd24, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000008e, 5'd19, 27'h00000240, 5'd0, 27'h0000010f, 32'h00000400,
  1'd1,  5'd6, 27'h000001e4, 5'd16, 27'h00000346, 5'd13, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018a, 5'd18, 27'h000003d0, 5'd25, 27'h00000284, 32'h00000400,
  1'd1,  5'd6, 27'h0000006e, 5'd29, 27'h00000273, 5'd4, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000016d, 5'd27, 27'h0000009e, 5'd13, 27'h00000378, 32'h00000400,
  1'd1,  5'd5, 27'h000000e4, 5'd29, 27'h0000015b, 5'd23, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b8, 5'd8, 27'h00000281, 5'd3, 27'h0000016f, 32'h00000400,
  1'd1,  5'd18, 27'h00000016, 5'd7, 27'h000000a3, 5'd11, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ba, 5'd9, 27'h000000ac, 5'd25, 27'h00000027, 32'h00000400,
  1'd1,  5'd17, 27'h000000ce, 5'd20, 27'h00000110, 5'd2, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000004b, 5'd17, 27'h00000014, 5'd10, 27'h000001e5, 32'h00000400,
  1'd1,  5'd18, 27'h000002e3, 5'd16, 27'h00000296, 5'd22, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e7, 5'd26, 27'h00000057, 5'd1, 27'h000003a1, 32'h00000400,
  1'd1,  5'd20, 27'h00000288, 5'd29, 27'h000002a8, 5'd12, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034e, 5'd28, 27'h000002cf, 5'd21, 27'h000001b1, 32'h00000400,
  1'd1,  5'd28, 27'h000001c2, 5'd7, 27'h00000301, 5'd2, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000255, 5'd9, 27'h00000105, 5'd14, 27'h00000352, 32'h00000400,
  1'd1,  5'd28, 27'h000000bb, 5'd8, 27'h0000007f, 5'd22, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000236, 5'd15, 27'h000003ff, 5'd0, 27'h000000b8, 32'h00000400,
  1'd1,  5'd30, 27'h0000018e, 5'd16, 27'h00000009, 5'd14, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000086, 5'd15, 27'h000002e8, 5'd25, 27'h00000045, 32'h00000400,
  1'd1,  5'd30, 27'h00000325, 5'd29, 27'h0000017a, 5'd3, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b2, 5'd29, 27'h00000292, 5'd10, 27'h000001cc, 32'h00000400,
  1'd1,  5'd26, 27'h000001df, 5'd26, 27'h00000095, 5'd23, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000285, 5'd5, 27'h00000113, 5'd9, 27'h00000156, 32'h00000400,
  1'd1,  5'd6, 27'h0000029a, 5'd9, 27'h000002ee, 5'd18, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000071, 5'd6, 27'h0000007d, 5'd26, 27'h000001ad, 32'h00000400,
  1'd1,  5'd6, 27'h000000bf, 5'd15, 27'h0000036c, 5'd7, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003aa, 5'd16, 27'h000001a6, 5'd20, 27'h00000003, 32'h00000400,
  1'd1,  5'd6, 27'h0000033c, 5'd18, 27'h0000004f, 5'd30, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a4, 5'd28, 27'h0000000f, 5'd8, 27'h000003bc, 32'h00000400,
  1'd1,  5'd6, 27'h00000390, 5'd29, 27'h00000310, 5'd19, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000020f, 5'd27, 27'h00000008, 5'd30, 27'h00000026, 32'h00000400,
  1'd1,  5'd18, 27'h0000001b, 5'd6, 27'h00000252, 5'd10, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000308, 5'd7, 27'h000001f8, 5'd15, 27'h000003de, 32'h00000400,
  1'd1,  5'd16, 27'h000001b3, 5'd6, 27'h000000b9, 5'd29, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000210, 5'd18, 27'h00000131, 5'd5, 27'h0000020e, 32'h00000400,
  1'd1,  5'd17, 27'h00000070, 5'd16, 27'h00000353, 5'd18, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002bd, 5'd15, 27'h0000024b, 5'd27, 27'h000002c8, 32'h00000400,
  1'd1,  5'd20, 27'h00000122, 5'd26, 27'h0000009a, 5'd9, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003f0, 5'd27, 27'h00000300, 5'd18, 27'h0000038b, 32'h00000400,
  1'd1,  5'd18, 27'h000002b2, 5'd28, 27'h000001c1, 5'd27, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000002e, 5'd5, 27'h00000142, 5'd6, 27'h00000196, 32'h00000400,
  1'd1,  5'd27, 27'h00000219, 5'd8, 27'h00000117, 5'd17, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000002f, 5'd9, 27'h0000026c, 5'd26, 27'h000001c1, 32'h00000400,
  1'd1,  5'd30, 27'h0000029b, 5'd17, 27'h0000014c, 5'd7, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000181, 5'd18, 27'h00000390, 5'd17, 27'h0000038b, 32'h00000400,
  1'd1,  5'd25, 27'h000003d6, 5'd19, 27'h0000000c, 5'd30, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000137, 5'd29, 27'h000001b4, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd30, 27'h000000f0, 5'd30, 27'h00000378, 5'd15, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b9, 5'd29, 27'h00000010, 5'd26, 27'h00000400, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000002f3, 5'd4, 27'h0000020a, 5'd3, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000031f, 5'd3, 27'h000002b8, 5'd12, 27'h000001aa, 32'h00000400,
  1'd1,  5'd4, 27'h00000121, 5'd4, 27'h000000bb, 5'd20, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001eb, 5'd10, 27'h0000018a, 5'd1, 27'h000002c5, 32'h00000400,
  1'd1,  5'd4, 27'h000001cc, 5'd15, 27'h0000005a, 5'd10, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000022b, 5'd11, 27'h0000006f, 5'd22, 27'h00000309, 32'h00000400,
  1'd1,  5'd2, 27'h000002c0, 5'd23, 27'h00000176, 5'd0, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000023d, 5'd24, 27'h0000022b, 5'd10, 27'h00000272, 32'h00000400,
  1'd1,  5'd1, 27'h000000bc, 5'd22, 27'h00000059, 5'd21, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c1, 5'd2, 27'h00000339, 5'd3, 27'h000000d7, 32'h00000400,
  1'd1,  5'd10, 27'h000003ec, 5'd3, 27'h0000028b, 5'd14, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000e8, 5'd1, 27'h00000338, 5'd25, 27'h00000163, 32'h00000400,
  1'd1,  5'd13, 27'h000000e3, 5'd14, 27'h0000039f, 5'd4, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003fd, 5'd12, 27'h000003c6, 5'd10, 27'h00000290, 32'h00000400,
  1'd1,  5'd14, 27'h000003dc, 5'd11, 27'h000002a8, 5'd24, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000083, 5'd22, 27'h00000066, 5'd3, 27'h00000272, 32'h00000400,
  1'd1,  5'd10, 27'h00000169, 5'd21, 27'h000002f4, 5'd12, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003af, 5'd25, 27'h00000183, 5'd21, 27'h0000011d, 32'h00000400,
  1'd1,  5'd22, 27'h000000ee, 5'd3, 27'h00000120, 5'd4, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a6, 5'd3, 27'h00000272, 5'd12, 27'h000003f7, 32'h00000400,
  1'd1,  5'd22, 27'h0000007f, 5'd0, 27'h00000305, 5'd21, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000098, 5'd13, 27'h000000dc, 5'd4, 27'h00000274, 32'h00000400,
  1'd1,  5'd24, 27'h0000023a, 5'd13, 27'h000002e5, 5'd15, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000028c, 5'd15, 27'h000000fe, 5'd21, 27'h000001c0, 32'h00000400,
  1'd1,  5'd25, 27'h00000002, 5'd22, 27'h000002e0, 5'd1, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000015a, 5'd22, 27'h000003bd, 5'd13, 27'h0000025b, 32'h00000400,
  1'd1,  5'd22, 27'h000003db, 5'd22, 27'h00000279, 5'd24, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000091, 5'd2, 27'h00000062, 5'd6, 27'h0000027d, 32'h00000400,
  1'd1,  5'd0, 27'h00000166, 5'd0, 27'h00000337, 5'd15, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000030d, 5'd5, 27'h0000003e, 5'd29, 27'h00000213, 32'h00000400,
  1'd1,  5'd4, 27'h00000026, 5'd10, 27'h000003a3, 5'd6, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f3, 5'd12, 27'h00000258, 5'd17, 27'h000002dc, 32'h00000400,
  1'd1,  5'd1, 27'h00000023, 5'd15, 27'h000001e6, 5'd30, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000002b, 5'd23, 27'h000003ea, 5'd6, 27'h000002a1, 32'h00000400,
  1'd1,  5'd1, 27'h00000306, 5'd21, 27'h00000080, 5'd19, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001cf, 5'd23, 27'h000001e2, 5'd29, 27'h000001d0, 32'h00000400,
  1'd1,  5'd11, 27'h000003ad, 5'd3, 27'h0000038b, 5'd6, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000013e, 5'd3, 27'h00000144, 5'd18, 27'h0000037e, 32'h00000400,
  1'd1,  5'd15, 27'h00000148, 5'd0, 27'h000002ed, 5'd26, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002f7, 5'd14, 27'h00000132, 5'd7, 27'h00000064, 32'h00000400,
  1'd1,  5'd13, 27'h000001d4, 5'd13, 27'h0000002f, 5'd19, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017c, 5'd12, 27'h00000226, 5'd30, 27'h000002f3, 32'h00000400,
  1'd1,  5'd11, 27'h000002d5, 5'd24, 27'h0000021c, 5'd5, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000325, 5'd23, 27'h00000078, 5'd18, 27'h000002d0, 32'h00000400,
  1'd1,  5'd14, 27'h000000ad, 5'd23, 27'h000001b3, 5'd27, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001fd, 5'd4, 27'h0000038d, 5'd9, 27'h0000016b, 32'h00000400,
  1'd1,  5'd24, 27'h00000177, 5'd0, 27'h00000218, 5'd17, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000039, 5'd1, 27'h000000d2, 5'd25, 27'h000003fc, 32'h00000400,
  1'd1,  5'd21, 27'h000000c9, 5'd13, 27'h00000164, 5'd6, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000263, 5'd13, 27'h000001d8, 5'd16, 27'h00000163, 32'h00000400,
  1'd1,  5'd21, 27'h00000102, 5'd11, 27'h0000022a, 5'd29, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000031e, 5'd20, 27'h0000035d, 5'd5, 27'h00000257, 32'h00000400,
  1'd1,  5'd22, 27'h000003d7, 5'd25, 27'h0000033a, 5'd20, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003df, 5'd21, 27'h00000190, 5'd26, 27'h00000005, 32'h00000400,
  1'd1,  5'd2, 27'h00000368, 5'd6, 27'h0000016f, 5'd0, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000053, 5'd9, 27'h00000343, 5'd11, 27'h000002b5, 32'h00000400,
  1'd1,  5'd1, 27'h00000366, 5'd6, 27'h000003d5, 5'd22, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b3, 5'd15, 27'h0000038d, 5'd2, 27'h000002d6, 32'h00000400,
  1'd1,  5'd3, 27'h0000039d, 5'd18, 27'h00000306, 5'd12, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003de, 5'd19, 27'h00000219, 5'd23, 27'h00000397, 32'h00000400,
  1'd1,  5'd4, 27'h0000001f, 5'd28, 27'h0000022a, 5'd4, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a3, 5'd27, 27'h00000121, 5'd11, 27'h0000037f, 32'h00000400,
  1'd1,  5'd3, 27'h0000012c, 5'd29, 27'h00000229, 5'd23, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000007d, 5'd8, 27'h000000e1, 5'd3, 27'h00000387, 32'h00000400,
  1'd1,  5'd11, 27'h0000039b, 5'd9, 27'h000003d4, 5'd14, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000015f, 5'd6, 27'h000002b8, 5'd22, 27'h00000106, 32'h00000400,
  1'd1,  5'd11, 27'h00000297, 5'd19, 27'h0000015a, 5'd2, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ff, 5'd16, 27'h0000000b, 5'd14, 27'h00000120, 32'h00000400,
  1'd1,  5'd11, 27'h00000197, 5'd16, 27'h000001e4, 5'd21, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001cb, 5'd28, 27'h00000092, 5'd3, 27'h000002c9, 32'h00000400,
  1'd1,  5'd13, 27'h0000014d, 5'd30, 27'h0000035d, 5'd15, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002a9, 5'd28, 27'h0000027e, 5'd24, 27'h000002e0, 32'h00000400,
  1'd1,  5'd25, 27'h0000024b, 5'd7, 27'h000001d9, 5'd0, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002e1, 5'd9, 27'h0000034e, 5'd12, 27'h000002df, 32'h00000400,
  1'd1,  5'd20, 27'h000002ff, 5'd9, 27'h00000185, 5'd24, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b9, 5'd19, 27'h000000d6, 5'd1, 27'h00000059, 32'h00000400,
  1'd1,  5'd24, 27'h00000013, 5'd16, 27'h00000106, 5'd13, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b3, 5'd20, 27'h000000d1, 5'd24, 27'h00000100, 32'h00000400,
  1'd1,  5'd20, 27'h0000033c, 5'd28, 27'h0000029a, 5'd2, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000225, 5'd30, 27'h00000001, 5'd11, 27'h000001f3, 32'h00000400,
  1'd1,  5'd23, 27'h000003e9, 5'd29, 27'h00000325, 5'd25, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002f, 5'd7, 27'h000000f9, 5'd6, 27'h000000e2, 32'h00000400,
  1'd1,  5'd1, 27'h00000290, 5'd5, 27'h000000de, 5'd15, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000071, 5'd7, 27'h00000074, 5'd26, 27'h00000209, 32'h00000400,
  1'd1,  5'd0, 27'h00000173, 5'd17, 27'h000002ec, 5'd9, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000033a, 5'd15, 27'h00000359, 5'd16, 27'h0000037e, 32'h00000400,
  1'd1,  5'd3, 27'h0000009a, 5'd20, 27'h00000209, 5'd29, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000385, 5'd26, 27'h0000032c, 5'd6, 27'h00000286, 32'h00000400,
  1'd1,  5'd2, 27'h000001fb, 5'd29, 27'h000002cd, 5'd17, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001aa, 5'd26, 27'h00000235, 5'd29, 27'h000002c0, 32'h00000400,
  1'd1,  5'd13, 27'h0000033a, 5'd9, 27'h000002d2, 5'd8, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b7, 5'd5, 27'h0000021a, 5'd18, 27'h000000eb, 32'h00000400,
  1'd1,  5'd13, 27'h000002af, 5'd10, 27'h00000087, 5'd27, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a1, 5'd18, 27'h000001f0, 5'd7, 27'h000002a3, 32'h00000400,
  1'd1,  5'd11, 27'h0000034f, 5'd16, 27'h00000217, 5'd18, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000019c, 5'd17, 27'h000000e9, 5'd30, 27'h00000121, 32'h00000400,
  1'd1,  5'd15, 27'h00000097, 5'd27, 27'h000002d7, 5'd8, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023f, 5'd26, 27'h00000145, 5'd19, 27'h00000274, 32'h00000400,
  1'd1,  5'd12, 27'h000002e6, 5'd28, 27'h0000035e, 5'd30, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f7, 5'd10, 27'h0000014e, 5'd7, 27'h000002ee, 32'h00000400,
  1'd1,  5'd22, 27'h000001a5, 5'd8, 27'h0000007d, 5'd18, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000012c, 5'd7, 27'h00000095, 5'd28, 27'h00000037, 32'h00000400,
  1'd1,  5'd24, 27'h00000046, 5'd17, 27'h000003a3, 5'd8, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001e7, 5'd16, 27'h00000347, 5'd16, 27'h000000fc, 32'h00000400,
  1'd1,  5'd24, 27'h00000155, 5'd15, 27'h0000036e, 5'd29, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bd, 5'd28, 27'h000001b9, 5'd5, 27'h00000288, 32'h00000400,
  1'd1,  5'd23, 27'h000000ef, 5'd27, 27'h000000da, 5'd17, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000182, 5'd25, 27'h000003bd, 5'd28, 27'h00000161, 32'h00000400,
  1'd1,  5'd5, 27'h0000031e, 5'd1, 27'h00000255, 5'd8, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000030c, 5'd3, 27'h0000034b, 5'd18, 27'h000001a6, 32'h00000400,
  1'd1,  5'd8, 27'h00000198, 5'd1, 27'h00000207, 5'd27, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001de, 5'd13, 27'h0000039a, 5'd4, 27'h0000013d, 32'h00000400,
  1'd1,  5'd5, 27'h00000322, 5'd10, 27'h00000385, 5'd12, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001cf, 5'd13, 27'h0000023b, 5'd20, 27'h000003d1, 32'h00000400,
  1'd1,  5'd10, 27'h0000003e, 5'd21, 27'h000002c5, 5'd3, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000198, 5'd21, 27'h000003c9, 5'd13, 27'h00000320, 32'h00000400,
  1'd1,  5'd8, 27'h00000374, 5'd25, 27'h00000281, 5'd21, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002bc, 5'd5, 27'h00000024, 5'd10, 27'h0000002b, 32'h00000400,
  1'd1,  5'd17, 27'h0000037b, 5'd3, 27'h00000029, 5'd16, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000232, 5'd0, 27'h00000074, 5'd26, 27'h000000d5, 32'h00000400,
  1'd1,  5'd17, 27'h000001e6, 5'd14, 27'h000000c1, 5'd1, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b9, 5'd14, 27'h00000172, 5'd11, 27'h000001bd, 32'h00000400,
  1'd1,  5'd16, 27'h000001ef, 5'd12, 27'h00000197, 5'd24, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000112, 5'd24, 27'h00000301, 5'd0, 27'h00000058, 32'h00000400,
  1'd1,  5'd19, 27'h00000092, 5'd20, 27'h00000379, 5'd11, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000028c, 5'd21, 27'h00000277, 5'd22, 27'h00000243, 32'h00000400,
  1'd1,  5'd28, 27'h00000019, 5'd4, 27'h00000292, 5'd2, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002cf, 5'd0, 27'h000002b6, 5'd11, 27'h00000214, 32'h00000400,
  1'd1,  5'd30, 27'h00000272, 5'd2, 27'h00000296, 5'd23, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000027d, 5'd10, 27'h00000188, 5'd3, 27'h000000c2, 32'h00000400,
  1'd1,  5'd29, 27'h000001c7, 5'd13, 27'h00000206, 5'd14, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ec, 5'd12, 27'h000000d7, 5'd25, 27'h0000019e, 32'h00000400,
  1'd1,  5'd27, 27'h000000c3, 5'd22, 27'h0000004a, 5'd0, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002db, 5'd22, 27'h000000cf, 5'd10, 27'h000002c5, 32'h00000400,
  1'd1,  5'd27, 27'h000003dd, 5'd23, 27'h000003e2, 5'd23, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000006b, 5'd0, 27'h00000327, 5'd3, 27'h000000f7, 32'h00000400,
  1'd1,  5'd7, 27'h00000044, 5'd0, 27'h00000104, 5'd13, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001d5, 5'd3, 27'h000002e5, 5'd24, 27'h0000014b, 32'h00000400,
  1'd1,  5'd5, 27'h00000388, 5'd11, 27'h0000000c, 5'd10, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a3, 5'd11, 27'h00000144, 5'd16, 27'h000003db, 32'h00000400,
  1'd1,  5'd6, 27'h000000c6, 5'd11, 27'h00000287, 5'd28, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000224, 5'd22, 27'h000000f1, 5'd5, 27'h000003ce, 32'h00000400,
  1'd1,  5'd8, 27'h000001f8, 5'd20, 27'h000002bd, 5'd16, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d3, 5'd24, 27'h00000001, 5'd26, 27'h00000338, 32'h00000400,
  1'd1,  5'd15, 27'h00000365, 5'd3, 27'h00000380, 5'd2, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000299, 5'd0, 27'h000000dc, 5'd10, 27'h0000035e, 32'h00000400,
  1'd1,  5'd17, 27'h000003d0, 5'd1, 27'h000001fc, 5'd24, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000096, 5'd12, 27'h000000d4, 5'd8, 27'h0000013d, 32'h00000400,
  1'd1,  5'd18, 27'h00000387, 5'd11, 27'h000002c7, 5'd17, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000042, 5'd10, 27'h000003b3, 5'd30, 27'h000001b6, 32'h00000400,
  1'd1,  5'd19, 27'h00000312, 5'd22, 27'h000002e4, 5'd7, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000205, 5'd23, 27'h00000091, 5'd18, 27'h00000111, 32'h00000400,
  1'd1,  5'd19, 27'h000000bc, 5'd23, 27'h0000029b, 5'd28, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000099, 5'd1, 27'h000001ed, 5'd6, 27'h0000023a, 32'h00000400,
  1'd1,  5'd29, 27'h000001c6, 5'd2, 27'h0000032c, 5'd17, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000030e, 5'd0, 27'h00000391, 5'd27, 27'h000000b5, 32'h00000400,
  1'd1,  5'd30, 27'h00000384, 5'd13, 27'h0000017a, 5'd8, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f7, 5'd14, 27'h0000032b, 5'd20, 27'h000000fe, 32'h00000400,
  1'd1,  5'd26, 27'h0000004e, 5'd14, 27'h0000030f, 5'd27, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c7, 5'd25, 27'h00000021, 5'd6, 27'h0000035f, 32'h00000400,
  1'd1,  5'd30, 27'h00000019, 5'd21, 27'h00000173, 5'd20, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000241, 5'd20, 27'h00000393, 5'd30, 27'h00000239, 32'h00000400,
  1'd1,  5'd8, 27'h00000358, 5'd6, 27'h00000016, 5'd1, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000297, 5'd5, 27'h00000139, 5'd11, 27'h000002ba, 32'h00000400,
  1'd1,  5'd9, 27'h000002db, 5'd7, 27'h00000113, 5'd21, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000216, 5'd19, 27'h00000175, 5'd5, 27'h00000008, 32'h00000400,
  1'd1,  5'd6, 27'h000002e4, 5'd17, 27'h0000008b, 5'd15, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000024f, 5'd18, 27'h00000317, 5'd21, 27'h0000037b, 32'h00000400,
  1'd1,  5'd5, 27'h000000eb, 5'd29, 27'h00000189, 5'd1, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000003d, 5'd26, 27'h0000019a, 5'd12, 27'h000002b9, 32'h00000400,
  1'd1,  5'd9, 27'h00000022, 5'd28, 27'h0000009a, 5'd23, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000307, 5'd8, 27'h0000010e, 5'd4, 27'h00000300, 32'h00000400,
  1'd1,  5'd16, 27'h000000ab, 5'd9, 27'h000002db, 5'd12, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000157, 5'd7, 27'h00000269, 5'd24, 27'h000000df, 32'h00000400,
  1'd1,  5'd20, 27'h000000ab, 5'd17, 27'h00000259, 5'd3, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003fd, 5'd18, 27'h00000275, 5'd10, 27'h0000022e, 32'h00000400,
  1'd1,  5'd18, 27'h00000259, 5'd18, 27'h00000059, 5'd23, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000299, 5'd26, 27'h000000cf, 5'd1, 27'h0000015a, 32'h00000400,
  1'd1,  5'd17, 27'h00000140, 5'd30, 27'h0000023a, 5'd14, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003de, 5'd28, 27'h000003e1, 5'd25, 27'h000000a4, 32'h00000400,
  1'd1,  5'd29, 27'h0000027e, 5'd7, 27'h0000021e, 5'd2, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c8, 5'd9, 27'h0000036d, 5'd12, 27'h00000359, 32'h00000400,
  1'd1,  5'd30, 27'h00000261, 5'd9, 27'h0000009e, 5'd22, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002b3, 5'd16, 27'h000001bb, 5'd3, 27'h0000038f, 32'h00000400,
  1'd1,  5'd27, 27'h00000306, 5'd20, 27'h00000177, 5'd11, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ce, 5'd16, 27'h000001da, 5'd22, 27'h00000218, 32'h00000400,
  1'd1,  5'd27, 27'h000003d6, 5'd29, 27'h000003b3, 5'd3, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000021c, 5'd25, 27'h000003d2, 5'd11, 27'h000000c5, 32'h00000400,
  1'd1,  5'd27, 27'h000001a8, 5'd26, 27'h0000036d, 5'd22, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000032, 5'd5, 27'h000001f8, 5'd7, 27'h00000062, 32'h00000400,
  1'd1,  5'd9, 27'h000001a6, 5'd6, 27'h0000005d, 5'd20, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000192, 5'd10, 27'h000000da, 5'd29, 27'h000003ea, 32'h00000400,
  1'd1,  5'd5, 27'h0000036a, 5'd17, 27'h000003e2, 5'd7, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000004, 5'd15, 27'h00000365, 5'd19, 27'h000001dc, 32'h00000400,
  1'd1,  5'd6, 27'h00000040, 5'd20, 27'h000000f9, 5'd30, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000037e, 5'd30, 27'h000003da, 5'd8, 27'h00000312, 32'h00000400,
  1'd1,  5'd7, 27'h000002fe, 5'd26, 27'h00000060, 5'd20, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000237, 5'd30, 27'h00000066, 5'd28, 27'h0000011c, 32'h00000400,
  1'd1,  5'd17, 27'h000001e9, 5'd9, 27'h000000fc, 5'd8, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000a5, 5'd8, 27'h00000207, 5'd17, 27'h000001fb, 32'h00000400,
  1'd1,  5'd16, 27'h00000192, 5'd10, 27'h00000066, 5'd29, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000168, 5'd16, 27'h000001f2, 5'd8, 27'h000003a3, 32'h00000400,
  1'd1,  5'd15, 27'h0000023b, 5'd19, 27'h00000113, 5'd16, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a8, 5'd17, 27'h000003c8, 5'd30, 27'h00000317, 32'h00000400,
  1'd1,  5'd19, 27'h00000075, 5'd27, 27'h000000f1, 5'd7, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000021f, 5'd29, 27'h0000011f, 5'd18, 27'h000000f2, 32'h00000400,
  1'd1,  5'd16, 27'h000003e7, 5'd28, 27'h000003ce, 5'd26, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000273, 5'd5, 27'h00000377, 5'd10, 27'h00000133, 32'h00000400,
  1'd1,  5'd28, 27'h0000027b, 5'd7, 27'h000001ea, 5'd18, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f0, 5'd6, 27'h000002a0, 5'd30, 27'h000002cf, 32'h00000400,
  1'd1,  5'd25, 27'h000003c3, 5'd15, 27'h000003e6, 5'd5, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000201, 5'd18, 27'h0000026c, 5'd20, 27'h00000012, 32'h00000400,
  1'd1,  5'd27, 27'h0000031e, 5'd16, 27'h0000002e, 5'd30, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f6, 5'd26, 27'h0000026e, 5'd10, 27'h0000000a, 32'h00000400,
  1'd1,  5'd26, 27'h000001bf, 5'd29, 27'h000002b3, 5'd16, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003be, 5'd30, 27'h00000193, 5'd30, 27'h000000c4, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000257, 5'd2, 27'h0000013c, 5'd3, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000339, 5'd3, 27'h00000366, 5'd13, 27'h00000066, 32'h00000400,
  1'd1,  5'd0, 27'h0000035d, 5'd5, 27'h00000047, 5'd24, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000031a, 5'd11, 27'h00000160, 5'd0, 27'h00000072, 32'h00000400,
  1'd1,  5'd3, 27'h00000262, 5'd15, 27'h0000010d, 5'd12, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000343, 5'd13, 27'h0000017d, 5'd24, 27'h00000070, 32'h00000400,
  1'd1,  5'd0, 27'h0000006e, 5'd25, 27'h00000204, 5'd1, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002a, 5'd25, 27'h00000280, 5'd13, 27'h000003f7, 32'h00000400,
  1'd1,  5'd4, 27'h0000026d, 5'd24, 27'h00000354, 5'd23, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ab, 5'd2, 27'h00000066, 5'd2, 27'h00000155, 32'h00000400,
  1'd1,  5'd15, 27'h00000154, 5'd0, 27'h00000143, 5'd12, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003b, 5'd2, 27'h00000303, 5'd22, 27'h000000e8, 32'h00000400,
  1'd1,  5'd11, 27'h0000025f, 5'd12, 27'h000000bc, 5'd2, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000158, 5'd12, 27'h00000343, 5'd12, 27'h000003e7, 32'h00000400,
  1'd1,  5'd12, 27'h000002f8, 5'd15, 27'h0000013e, 5'd23, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000037c, 5'd23, 27'h000003f9, 5'd3, 27'h00000046, 32'h00000400,
  1'd1,  5'd12, 27'h00000183, 5'd21, 27'h00000211, 5'd12, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a8, 5'd22, 27'h0000039d, 5'd25, 27'h0000007d, 32'h00000400,
  1'd1,  5'd22, 27'h000002ea, 5'd2, 27'h0000009b, 5'd4, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002c8, 5'd4, 27'h00000035, 5'd13, 27'h0000002a, 32'h00000400,
  1'd1,  5'd22, 27'h0000018f, 5'd3, 27'h00000287, 5'd23, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000006f, 5'd10, 27'h00000374, 5'd4, 27'h000002ec, 32'h00000400,
  1'd1,  5'd23, 27'h00000269, 5'd12, 27'h000003b2, 5'd14, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000a1, 5'd14, 27'h000003a6, 5'd21, 27'h00000037, 32'h00000400,
  1'd1,  5'd25, 27'h00000128, 5'd24, 27'h00000291, 5'd2, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d5, 5'd22, 27'h0000030c, 5'd12, 27'h00000032, 32'h00000400,
  1'd1,  5'd22, 27'h00000377, 5'd21, 27'h000003a3, 5'd21, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000063, 5'd1, 27'h00000200, 5'd7, 27'h00000004, 32'h00000400,
  1'd1,  5'd4, 27'h0000002c, 5'd1, 27'h000003cc, 5'd17, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b0, 5'd3, 27'h00000346, 5'd26, 27'h000000fb, 32'h00000400,
  1'd1,  5'd0, 27'h0000035a, 5'd14, 27'h00000395, 5'd6, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d9, 5'd10, 27'h0000025a, 5'd18, 27'h000001ad, 32'h00000400,
  1'd1,  5'd5, 27'h00000057, 5'd15, 27'h00000082, 5'd29, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000044, 5'd23, 27'h00000180, 5'd6, 27'h000001d8, 32'h00000400,
  1'd1,  5'd2, 27'h0000019c, 5'd25, 27'h000002a5, 5'd16, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001c3, 5'd25, 27'h00000323, 5'd30, 27'h000001dd, 32'h00000400,
  1'd1,  5'd12, 27'h0000032e, 5'd4, 27'h00000162, 5'd9, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a3, 5'd0, 27'h00000392, 5'd19, 27'h000001da, 32'h00000400,
  1'd1,  5'd12, 27'h000001f4, 5'd0, 27'h000002f1, 5'd28, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000fc, 5'd15, 27'h000000ef, 5'd7, 27'h00000303, 32'h00000400,
  1'd1,  5'd11, 27'h00000207, 5'd15, 27'h00000144, 5'd20, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000129, 5'd14, 27'h00000400, 5'd29, 27'h00000215, 32'h00000400,
  1'd1,  5'd15, 27'h000001b2, 5'd24, 27'h000000ff, 5'd5, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000120, 5'd22, 27'h000002ca, 5'd20, 27'h0000006d, 32'h00000400,
  1'd1,  5'd10, 27'h00000381, 5'd23, 27'h00000393, 5'd28, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000115, 5'd3, 27'h0000002c, 5'd5, 27'h0000019b, 32'h00000400,
  1'd1,  5'd23, 27'h00000068, 5'd3, 27'h0000002f, 5'd19, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000238, 5'd4, 27'h000001ec, 5'd29, 27'h0000016a, 32'h00000400,
  1'd1,  5'd22, 27'h00000283, 5'd12, 27'h000003d1, 5'd9, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a0, 5'd14, 27'h00000277, 5'd17, 27'h00000115, 32'h00000400,
  1'd1,  5'd23, 27'h0000013a, 5'd13, 27'h00000179, 5'd29, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d7, 5'd22, 27'h00000253, 5'd7, 27'h00000339, 32'h00000400,
  1'd1,  5'd21, 27'h00000019, 5'd23, 27'h000001f0, 5'd16, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000294, 5'd25, 27'h0000010b, 5'd27, 27'h0000028a, 32'h00000400,
  1'd1,  5'd1, 27'h0000032f, 5'd6, 27'h00000014, 5'd3, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002a4, 5'd7, 27'h0000000b, 5'd14, 27'h000003f0, 32'h00000400,
  1'd1,  5'd0, 27'h00000034, 5'd6, 27'h0000020f, 5'd24, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000085, 5'd18, 27'h000000f4, 5'd0, 27'h00000031, 32'h00000400,
  1'd1,  5'd4, 27'h000000b6, 5'd16, 27'h000000d1, 5'd13, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000034d, 5'd17, 27'h000003af, 5'd25, 27'h000002c5, 32'h00000400,
  1'd1,  5'd1, 27'h000001e5, 5'd27, 27'h000001a5, 5'd3, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000041, 5'd28, 27'h00000236, 5'd12, 27'h00000282, 32'h00000400,
  1'd1,  5'd1, 27'h000002d4, 5'd27, 27'h00000189, 5'd24, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000021b, 5'd5, 27'h000002fa, 5'd4, 27'h000001ba, 32'h00000400,
  1'd1,  5'd10, 27'h000003c5, 5'd6, 27'h000002c7, 5'd13, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e4, 5'd8, 27'h00000155, 5'd24, 27'h00000018, 32'h00000400,
  1'd1,  5'd15, 27'h0000004b, 5'd16, 27'h00000062, 5'd2, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ae, 5'd18, 27'h0000020f, 5'd15, 27'h00000194, 32'h00000400,
  1'd1,  5'd13, 27'h000002d8, 5'd19, 27'h00000026, 5'd21, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000200, 5'd29, 27'h000003e0, 5'd1, 27'h000003fb, 32'h00000400,
  1'd1,  5'd11, 27'h000000e0, 5'd27, 27'h000000f8, 5'd12, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000014c, 5'd25, 27'h00000377, 5'd21, 27'h00000127, 32'h00000400,
  1'd1,  5'd21, 27'h000000cf, 5'd7, 27'h00000241, 5'd1, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000015c, 5'd5, 27'h00000215, 5'd15, 27'h000001f2, 32'h00000400,
  1'd1,  5'd23, 27'h0000016e, 5'd9, 27'h00000391, 5'd24, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000396, 5'd18, 27'h000002d1, 5'd0, 27'h00000301, 32'h00000400,
  1'd1,  5'd20, 27'h000003f1, 5'd19, 27'h00000190, 5'd13, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000276, 5'd16, 27'h000003ee, 5'd24, 27'h0000034f, 32'h00000400,
  1'd1,  5'd21, 27'h00000367, 5'd29, 27'h00000030, 5'd0, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022a, 5'd30, 27'h0000005a, 5'd13, 27'h0000008b, 32'h00000400,
  1'd1,  5'd21, 27'h000000f3, 5'd26, 27'h000003db, 5'd23, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c1, 5'd8, 27'h000000f1, 5'd6, 27'h0000034a, 32'h00000400,
  1'd1,  5'd3, 27'h0000034c, 5'd9, 27'h00000146, 5'd15, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000164, 5'd6, 27'h000002b9, 5'd28, 27'h0000006e, 32'h00000400,
  1'd1,  5'd4, 27'h000003b9, 5'd18, 27'h000002d7, 5'd9, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b0, 5'd15, 27'h0000023d, 5'd20, 27'h00000105, 32'h00000400,
  1'd1,  5'd3, 27'h000000fa, 5'd20, 27'h00000211, 5'd30, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000003f, 5'd28, 27'h0000021e, 5'd5, 27'h00000115, 32'h00000400,
  1'd1,  5'd1, 27'h0000020f, 5'd29, 27'h000000b1, 5'd18, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002b0, 5'd30, 27'h000002f1, 5'd27, 27'h0000025c, 32'h00000400,
  1'd1,  5'd10, 27'h0000030f, 5'd7, 27'h00000176, 5'd8, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000391, 5'd8, 27'h0000021d, 5'd16, 27'h00000228, 32'h00000400,
  1'd1,  5'd10, 27'h000003bf, 5'd7, 27'h000003e0, 5'd27, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000223, 5'd20, 27'h00000237, 5'd5, 27'h00000164, 32'h00000400,
  1'd1,  5'd12, 27'h0000039d, 5'd15, 27'h00000284, 5'd19, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000132, 5'd17, 27'h00000151, 5'd26, 27'h000001f6, 32'h00000400,
  1'd1,  5'd12, 27'h00000291, 5'd30, 27'h000000f4, 5'd9, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000018a, 5'd27, 27'h00000131, 5'd20, 27'h0000026b, 32'h00000400,
  1'd1,  5'd12, 27'h00000296, 5'd30, 27'h00000073, 5'd30, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000022e, 5'd8, 27'h00000290, 5'd5, 27'h00000183, 32'h00000400,
  1'd1,  5'd25, 27'h00000153, 5'd5, 27'h00000229, 5'd17, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000012a, 5'd9, 27'h00000139, 5'd28, 27'h000002eb, 32'h00000400,
  1'd1,  5'd24, 27'h0000037e, 5'd17, 27'h00000097, 5'd9, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000027f, 5'd17, 27'h0000017b, 5'd18, 27'h00000078, 32'h00000400,
  1'd1,  5'd23, 27'h000000b4, 5'd17, 27'h000003c4, 5'd26, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000019e, 5'd28, 27'h00000282, 5'd5, 27'h000001b6, 32'h00000400,
  1'd1,  5'd25, 27'h00000004, 5'd29, 27'h00000204, 5'd20, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000005, 5'd27, 27'h0000036b, 5'd28, 27'h00000019, 32'h00000400,
  1'd1,  5'd6, 27'h000000ce, 5'd2, 27'h00000196, 5'd6, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000019c, 5'd2, 27'h0000021c, 5'd16, 27'h0000015a, 32'h00000400,
  1'd1,  5'd5, 27'h00000264, 5'd2, 27'h000001e8, 5'd27, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000059, 5'd11, 27'h00000223, 5'd4, 27'h00000001, 32'h00000400,
  1'd1,  5'd7, 27'h0000024d, 5'd13, 27'h00000207, 5'd13, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000c3, 5'd13, 27'h0000006a, 5'd25, 27'h0000009a, 32'h00000400,
  1'd1,  5'd9, 27'h000001a7, 5'd23, 27'h000002a8, 5'd4, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000032c, 5'd24, 27'h0000007d, 5'd12, 27'h0000024d, 32'h00000400,
  1'd1,  5'd7, 27'h00000331, 5'd22, 27'h0000000b, 5'd24, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002f, 5'd0, 27'h000003eb, 5'd10, 27'h0000013c, 32'h00000400,
  1'd1,  5'd17, 27'h0000027b, 5'd2, 27'h0000012b, 5'd17, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d7, 5'd0, 27'h000001ad, 5'd28, 27'h0000007b, 32'h00000400,
  1'd1,  5'd15, 27'h000002c9, 5'd12, 27'h00000224, 5'd0, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000360, 5'd14, 27'h0000003a, 5'd12, 27'h000003ef, 32'h00000400,
  1'd1,  5'd18, 27'h0000035e, 5'd12, 27'h000003c4, 5'd21, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000242, 5'd25, 27'h000001de, 5'd5, 27'h00000007, 32'h00000400,
  1'd1,  5'd17, 27'h000000ad, 5'd23, 27'h00000069, 5'd13, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000020b, 5'd23, 27'h0000029d, 5'd22, 27'h0000004e, 32'h00000400,
  1'd1,  5'd26, 27'h000003df, 5'd2, 27'h0000001f, 5'd1, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000de, 5'd1, 27'h0000001d, 5'd10, 27'h000003a3, 32'h00000400,
  1'd1,  5'd27, 27'h00000093, 5'd1, 27'h000000aa, 5'd23, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000dc, 5'd14, 27'h000002bd, 5'd0, 27'h00000252, 32'h00000400,
  1'd1,  5'd27, 27'h000002a6, 5'd14, 27'h000003e7, 5'd14, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000038d, 5'd14, 27'h00000268, 5'd22, 27'h0000028f, 32'h00000400,
  1'd1,  5'd29, 27'h000003cc, 5'd23, 27'h000002c0, 5'd3, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001e5, 5'd22, 27'h0000007c, 5'd12, 27'h000001be, 32'h00000400,
  1'd1,  5'd30, 27'h000003b8, 5'd22, 27'h000000bb, 5'd24, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000359, 5'd0, 27'h00000374, 5'd3, 27'h000001c4, 32'h00000400,
  1'd1,  5'd6, 27'h000000bf, 5'd0, 27'h000001da, 5'd12, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c1, 5'd4, 27'h00000063, 5'd22, 27'h00000101, 32'h00000400,
  1'd1,  5'd9, 27'h000000a2, 5'd13, 27'h00000381, 5'd7, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000146, 5'd11, 27'h00000062, 5'd18, 27'h00000192, 32'h00000400,
  1'd1,  5'd8, 27'h0000038e, 5'd13, 27'h00000369, 5'd30, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000014a, 5'd21, 27'h000002db, 5'd6, 27'h0000022c, 32'h00000400,
  1'd1,  5'd10, 27'h00000080, 5'd24, 27'h00000046, 5'd16, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000013c, 5'd22, 27'h00000105, 5'd29, 27'h00000171, 32'h00000400,
  1'd1,  5'd15, 27'h0000027d, 5'd1, 27'h00000252, 5'd5, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019d, 5'd4, 27'h000000b3, 5'd12, 27'h000000b0, 32'h00000400,
  1'd1,  5'd16, 27'h00000384, 5'd3, 27'h000000ff, 5'd21, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a0, 5'd11, 27'h00000066, 5'd7, 27'h00000059, 32'h00000400,
  1'd1,  5'd19, 27'h000003d9, 5'd14, 27'h0000006e, 5'd20, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000dc, 5'd10, 27'h0000031b, 5'd30, 27'h000000c9, 32'h00000400,
  1'd1,  5'd17, 27'h00000022, 5'd24, 27'h000001e4, 5'd6, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000186, 5'd24, 27'h00000307, 5'd15, 27'h00000203, 32'h00000400,
  1'd1,  5'd19, 27'h00000164, 5'd22, 27'h0000030e, 5'd30, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000009a, 5'd0, 27'h00000189, 5'd9, 27'h000002d7, 32'h00000400,
  1'd1,  5'd27, 27'h000001b7, 5'd4, 27'h000003c9, 5'd18, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000358, 5'd0, 27'h000003ad, 5'd29, 27'h00000100, 32'h00000400,
  1'd1,  5'd28, 27'h00000210, 5'd11, 27'h00000090, 5'd7, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000144, 5'd14, 27'h000003d8, 5'd20, 27'h0000003d, 32'h00000400,
  1'd1,  5'd27, 27'h000003ed, 5'd11, 27'h0000034b, 5'd27, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000281, 5'd23, 27'h00000318, 5'd6, 27'h000000d5, 32'h00000400,
  1'd1,  5'd28, 27'h0000019e, 5'd21, 27'h000002da, 5'd20, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000361, 5'd23, 27'h00000074, 5'd28, 27'h00000231, 32'h00000400,
  1'd1,  5'd7, 27'h000000ab, 5'd9, 27'h0000031b, 5'd0, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000032, 5'd9, 27'h000001c0, 5'd10, 27'h00000302, 32'h00000400,
  1'd1,  5'd6, 27'h00000332, 5'd8, 27'h000003b6, 5'd21, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003fe, 5'd16, 27'h00000273, 5'd1, 27'h00000289, 32'h00000400,
  1'd1,  5'd10, 27'h0000013f, 5'd17, 27'h00000295, 5'd10, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000173, 5'd17, 27'h000003c4, 5'd22, 27'h00000228, 32'h00000400,
  1'd1,  5'd8, 27'h0000029c, 5'd28, 27'h00000068, 5'd4, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001bc, 5'd27, 27'h00000332, 5'd13, 27'h000003e4, 32'h00000400,
  1'd1,  5'd7, 27'h0000012b, 5'd30, 27'h000003b2, 5'd20, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000006c, 5'd6, 27'h000002a5, 5'd0, 27'h00000136, 32'h00000400,
  1'd1,  5'd19, 27'h0000028b, 5'd5, 27'h00000110, 5'd13, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f6, 5'd6, 27'h0000004e, 5'd25, 27'h0000000c, 32'h00000400,
  1'd1,  5'd19, 27'h00000378, 5'd16, 27'h00000117, 5'd2, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000373, 5'd16, 27'h00000276, 5'd13, 27'h00000289, 32'h00000400,
  1'd1,  5'd18, 27'h0000034b, 5'd19, 27'h0000014b, 5'd23, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000127, 5'd26, 27'h00000123, 5'd2, 27'h000001a5, 32'h00000400,
  1'd1,  5'd20, 27'h00000249, 5'd30, 27'h000003c1, 5'd12, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003fc, 5'd28, 27'h00000150, 5'd21, 27'h000000f6, 32'h00000400,
  1'd1,  5'd30, 27'h000000c5, 5'd9, 27'h000003de, 5'd2, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012b, 5'd7, 27'h00000294, 5'd11, 27'h0000025b, 32'h00000400,
  1'd1,  5'd27, 27'h000002c3, 5'd7, 27'h00000309, 5'd20, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000030d, 5'd15, 27'h0000033a, 5'd3, 27'h0000038e, 32'h00000400,
  1'd1,  5'd30, 27'h00000064, 5'd19, 27'h000002a0, 5'd11, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003ea, 5'd18, 27'h00000063, 5'd25, 27'h00000321, 32'h00000400,
  1'd1,  5'd26, 27'h00000061, 5'd29, 27'h000001f6, 5'd3, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ff, 5'd25, 27'h00000362, 5'd10, 27'h000001e1, 32'h00000400,
  1'd1,  5'd30, 27'h000003c4, 5'd27, 27'h000003f0, 5'd23, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000024a, 5'd7, 27'h0000009b, 5'd8, 27'h000003c5, 32'h00000400,
  1'd1,  5'd5, 27'h00000230, 5'd5, 27'h0000030b, 5'd18, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000114, 5'd6, 27'h000000ed, 5'd27, 27'h00000015, 32'h00000400,
  1'd1,  5'd6, 27'h0000010c, 5'd20, 27'h000001ec, 5'd9, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e7, 5'd16, 27'h0000034f, 5'd17, 27'h000001fa, 32'h00000400,
  1'd1,  5'd9, 27'h00000110, 5'd16, 27'h000000fa, 5'd30, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000296, 5'd30, 27'h0000015f, 5'd7, 27'h00000037, 32'h00000400,
  1'd1,  5'd7, 27'h00000305, 5'd27, 27'h000002ae, 5'd20, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000fd, 5'd28, 27'h00000300, 5'd30, 27'h000002ad, 32'h00000400,
  1'd1,  5'd19, 27'h0000004d, 5'd5, 27'h000002c6, 5'd6, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000006c, 5'd9, 27'h00000076, 5'd17, 27'h0000016d, 32'h00000400,
  1'd1,  5'd19, 27'h00000185, 5'd10, 27'h00000025, 5'd29, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ca, 5'd18, 27'h00000087, 5'd5, 27'h000001b4, 32'h00000400,
  1'd1,  5'd18, 27'h000000bb, 5'd17, 27'h000003f5, 5'd19, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000186, 5'd18, 27'h00000369, 5'd30, 27'h000002b7, 32'h00000400,
  1'd1,  5'd15, 27'h000003d4, 5'd26, 27'h000003bd, 5'd7, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000346, 5'd30, 27'h000000db, 5'd18, 27'h00000355, 32'h00000400,
  1'd1,  5'd16, 27'h0000029b, 5'd27, 27'h00000289, 5'd30, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ce, 5'd9, 27'h00000334, 5'd9, 27'h000001e3, 32'h00000400,
  1'd1,  5'd28, 27'h0000023c, 5'd8, 27'h0000022e, 5'd15, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b2, 5'd9, 27'h00000147, 5'd30, 27'h0000018a, 32'h00000400,
  1'd1,  5'd28, 27'h00000249, 5'd16, 27'h000003b1, 5'd5, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003bc, 5'd18, 27'h000002ae, 5'd20, 27'h000001ce, 32'h00000400,
  1'd1,  5'd27, 27'h000001cf, 5'd18, 27'h00000312, 5'd29, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000219, 5'd27, 27'h000002c5, 5'd8, 27'h00000222, 32'h00000400,
  1'd1,  5'd28, 27'h0000011c, 5'd29, 27'h0000019c, 5'd20, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000d4, 5'd28, 27'h00000075, 5'd28, 27'h00000063, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000002f9, 5'd2, 27'h00000361, 5'd5, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000049, 5'd1, 27'h0000026d, 5'd13, 27'h0000022c, 32'h00000400,
  1'd1,  5'd0, 27'h000002cc, 5'd2, 27'h00000380, 5'd24, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e1, 5'd11, 27'h000003a9, 5'd3, 27'h00000317, 32'h00000400,
  1'd1,  5'd4, 27'h0000005d, 5'd11, 27'h0000015b, 5'd11, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000345, 5'd11, 27'h00000006, 5'd25, 27'h000001fe, 32'h00000400,
  1'd1,  5'd2, 27'h00000372, 5'd21, 27'h0000035e, 5'd3, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000300, 5'd25, 27'h00000108, 5'd13, 27'h000000ab, 32'h00000400,
  1'd1,  5'd2, 27'h00000133, 5'd24, 27'h000001ff, 5'd21, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f6, 5'd1, 27'h00000294, 5'd1, 27'h0000011f, 32'h00000400,
  1'd1,  5'd14, 27'h00000043, 5'd4, 27'h000000fc, 5'd13, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000271, 5'd0, 27'h0000014d, 5'd20, 27'h000002ff, 32'h00000400,
  1'd1,  5'd10, 27'h0000035e, 5'd10, 27'h000002a5, 5'd4, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d0, 5'd14, 27'h00000377, 5'd13, 27'h0000018a, 32'h00000400,
  1'd1,  5'd10, 27'h0000039e, 5'd15, 27'h00000171, 5'd21, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003cb, 5'd24, 27'h000002b0, 5'd4, 27'h00000122, 32'h00000400,
  1'd1,  5'd13, 27'h000000ec, 5'd22, 27'h000000f4, 5'd10, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000049, 5'd21, 27'h000000ce, 5'd22, 27'h000001d7, 32'h00000400,
  1'd1,  5'd24, 27'h000001f0, 5'd3, 27'h000003a2, 5'd1, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000340, 5'd0, 27'h00000375, 5'd12, 27'h000002e8, 32'h00000400,
  1'd1,  5'd24, 27'h000001fc, 5'd2, 27'h00000372, 5'd25, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ae, 5'd11, 27'h00000326, 5'd4, 27'h00000058, 32'h00000400,
  1'd1,  5'd23, 27'h000000b4, 5'd15, 27'h00000089, 5'd14, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f8, 5'd10, 27'h00000319, 5'd25, 27'h00000252, 32'h00000400,
  1'd1,  5'd21, 27'h0000019d, 5'd21, 27'h000002a5, 5'd5, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000057, 5'd21, 27'h00000207, 5'd11, 27'h000002c1, 32'h00000400,
  1'd1,  5'd24, 27'h0000033c, 5'd24, 27'h000001db, 5'd25, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022d, 5'd1, 27'h000003f3, 5'd8, 27'h00000017, 32'h00000400,
  1'd1,  5'd2, 27'h00000284, 5'd0, 27'h000001e2, 5'd16, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000009d, 5'd2, 27'h000000a4, 5'd26, 27'h00000142, 32'h00000400,
  1'd1,  5'd3, 27'h00000298, 5'd12, 27'h000000c2, 5'd8, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f2, 5'd13, 27'h000003ce, 5'd18, 27'h00000163, 32'h00000400,
  1'd1,  5'd1, 27'h000003c5, 5'd12, 27'h0000009f, 5'd29, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039b, 5'd25, 27'h000000fc, 5'd9, 27'h00000100, 32'h00000400,
  1'd1,  5'd0, 27'h00000365, 5'd21, 27'h00000070, 5'd16, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000282, 5'd21, 27'h0000031a, 5'd29, 27'h000001c8, 32'h00000400,
  1'd1,  5'd11, 27'h00000278, 5'd0, 27'h00000189, 5'd6, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000182, 5'd2, 27'h000001c2, 5'd18, 27'h000003d6, 32'h00000400,
  1'd1,  5'd12, 27'h00000225, 5'd0, 27'h00000040, 5'd26, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000036a, 5'd13, 27'h00000360, 5'd7, 27'h00000149, 32'h00000400,
  1'd1,  5'd12, 27'h00000207, 5'd13, 27'h000000ef, 5'd19, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f6, 5'd13, 27'h00000234, 5'd29, 27'h000002e2, 32'h00000400,
  1'd1,  5'd14, 27'h000000dd, 5'd24, 27'h000002a6, 5'd10, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ec, 5'd22, 27'h000002bc, 5'd17, 27'h000003cc, 32'h00000400,
  1'd1,  5'd11, 27'h000001f1, 5'd21, 27'h000001fc, 5'd27, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000025, 5'd2, 27'h00000194, 5'd6, 27'h00000015, 32'h00000400,
  1'd1,  5'd24, 27'h000001ed, 5'd1, 27'h00000099, 5'd18, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000019, 5'd3, 27'h0000009a, 5'd29, 27'h00000388, 32'h00000400,
  1'd1,  5'd24, 27'h00000087, 5'd13, 27'h00000287, 5'd6, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a1, 5'd13, 27'h0000034d, 5'd19, 27'h00000223, 32'h00000400,
  1'd1,  5'd24, 27'h00000153, 5'd15, 27'h000000a0, 5'd27, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003b3, 5'd25, 27'h00000109, 5'd6, 27'h00000066, 32'h00000400,
  1'd1,  5'd21, 27'h000002b6, 5'd23, 27'h000003d6, 5'd17, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f5, 5'd22, 27'h0000024a, 5'd27, 27'h00000084, 32'h00000400,
  1'd1,  5'd4, 27'h00000101, 5'd8, 27'h0000010e, 5'd1, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000136, 5'd5, 27'h00000238, 5'd11, 27'h0000012b, 32'h00000400,
  1'd1,  5'd1, 27'h000000c3, 5'd7, 27'h00000224, 5'd25, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000019b, 5'd20, 27'h00000262, 5'd3, 27'h0000038d, 32'h00000400,
  1'd1,  5'd2, 27'h0000013d, 5'd19, 27'h000003bc, 5'd13, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036d, 5'd16, 27'h00000235, 5'd22, 27'h00000348, 32'h00000400,
  1'd1,  5'd0, 27'h000003e2, 5'd29, 27'h00000253, 5'd4, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d4, 5'd27, 27'h00000341, 5'd10, 27'h000003be, 32'h00000400,
  1'd1,  5'd0, 27'h000002d1, 5'd26, 27'h000000c8, 5'd25, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000022f, 5'd10, 27'h0000000a, 5'd4, 27'h00000202, 32'h00000400,
  1'd1,  5'd13, 27'h00000261, 5'd8, 27'h0000025c, 5'd11, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000294, 5'd8, 27'h000003b8, 5'd25, 27'h0000023e, 32'h00000400,
  1'd1,  5'd12, 27'h00000256, 5'd18, 27'h0000030e, 5'd0, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003fa, 5'd18, 27'h000001e1, 5'd14, 27'h000000dd, 32'h00000400,
  1'd1,  5'd12, 27'h0000011c, 5'd17, 27'h0000018d, 5'd25, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000167, 5'd26, 27'h000002fd, 5'd3, 27'h0000023c, 32'h00000400,
  1'd1,  5'd13, 27'h00000291, 5'd26, 27'h00000075, 5'd14, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fe, 5'd28, 27'h000002e9, 5'd24, 27'h000001d5, 32'h00000400,
  1'd1,  5'd22, 27'h0000001a, 5'd5, 27'h000003a9, 5'd0, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000053, 5'd9, 27'h00000051, 5'd13, 27'h000001dc, 32'h00000400,
  1'd1,  5'd23, 27'h00000271, 5'd8, 27'h00000199, 5'd24, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002aa, 5'd15, 27'h000002c9, 5'd3, 27'h000002ec, 32'h00000400,
  1'd1,  5'd22, 27'h000000d5, 5'd18, 27'h000002f6, 5'd10, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000329, 5'd18, 27'h0000005f, 5'd24, 27'h00000083, 32'h00000400,
  1'd1,  5'd22, 27'h00000306, 5'd26, 27'h000003a9, 5'd0, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ac, 5'd29, 27'h00000233, 5'd15, 27'h00000076, 32'h00000400,
  1'd1,  5'd25, 27'h00000186, 5'd28, 27'h00000396, 5'd20, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000285, 5'd5, 27'h00000102, 5'd5, 27'h00000115, 32'h00000400,
  1'd1,  5'd2, 27'h000003c4, 5'd6, 27'h00000033, 5'd17, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b3, 5'd5, 27'h000002b9, 5'd30, 27'h000003d6, 32'h00000400,
  1'd1,  5'd1, 27'h0000011a, 5'd15, 27'h00000215, 5'd7, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f2, 5'd16, 27'h000002f0, 5'd17, 27'h00000289, 32'h00000400,
  1'd1,  5'd3, 27'h00000317, 5'd20, 27'h00000032, 5'd28, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002be, 5'd30, 27'h00000040, 5'd6, 27'h00000032, 32'h00000400,
  1'd1,  5'd2, 27'h00000247, 5'd28, 27'h0000021f, 5'd17, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000147, 5'd30, 27'h0000038c, 5'd26, 27'h00000074, 32'h00000400,
  1'd1,  5'd12, 27'h000000e6, 5'd5, 27'h000003b8, 5'd8, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000004f, 5'd9, 27'h000003ee, 5'd17, 27'h00000092, 32'h00000400,
  1'd1,  5'd14, 27'h0000034a, 5'd9, 27'h00000344, 5'd30, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a0, 5'd17, 27'h000002f7, 5'd6, 27'h00000331, 32'h00000400,
  1'd1,  5'd14, 27'h00000293, 5'd16, 27'h0000008e, 5'd16, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000186, 5'd17, 27'h000001f3, 5'd28, 27'h000000e6, 32'h00000400,
  1'd1,  5'd12, 27'h000001ed, 5'd25, 27'h000003f2, 5'd10, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000033a, 5'd25, 27'h0000037b, 5'd19, 27'h00000202, 32'h00000400,
  1'd1,  5'd13, 27'h000001b7, 5'd30, 27'h00000027, 5'd30, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000186, 5'd9, 27'h000001e9, 5'd9, 27'h000001f4, 32'h00000400,
  1'd1,  5'd21, 27'h00000378, 5'd6, 27'h0000030f, 5'd19, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000009b, 5'd7, 27'h000003d3, 5'd30, 27'h0000035b, 32'h00000400,
  1'd1,  5'd24, 27'h000000fb, 5'd20, 27'h00000139, 5'd9, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000317, 5'd19, 27'h000000cf, 5'd18, 27'h0000017b, 32'h00000400,
  1'd1,  5'd24, 27'h00000298, 5'd20, 27'h000001ad, 5'd29, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000c7, 5'd30, 27'h000003b8, 5'd9, 27'h00000113, 32'h00000400,
  1'd1,  5'd23, 27'h0000011b, 5'd27, 27'h00000100, 5'd19, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c8, 5'd29, 27'h00000306, 5'd30, 27'h0000008b, 32'h00000400,
  1'd1,  5'd8, 27'h00000220, 5'd2, 27'h00000160, 5'd8, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000079, 5'd4, 27'h000001a6, 5'd15, 27'h00000373, 32'h00000400,
  1'd1,  5'd10, 27'h000000bd, 5'd3, 27'h00000326, 5'd29, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ef, 5'd11, 27'h00000174, 5'd3, 27'h00000134, 32'h00000400,
  1'd1,  5'd5, 27'h000002bf, 5'd14, 27'h000002cf, 5'd12, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000236, 5'd14, 27'h00000176, 5'd23, 27'h0000016e, 32'h00000400,
  1'd1,  5'd9, 27'h00000242, 5'd22, 27'h0000014d, 5'd3, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f2, 5'd24, 27'h0000018a, 5'd13, 27'h000003f2, 32'h00000400,
  1'd1,  5'd5, 27'h0000026c, 5'd21, 27'h0000007f, 5'd23, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025c, 5'd1, 27'h000001ea, 5'd5, 27'h0000015d, 32'h00000400,
  1'd1,  5'd17, 27'h000000be, 5'd0, 27'h00000147, 5'd20, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a5, 5'd3, 27'h00000146, 5'd28, 27'h00000057, 32'h00000400,
  1'd1,  5'd19, 27'h00000069, 5'd10, 27'h000001d9, 5'd3, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000188, 5'd10, 27'h0000020f, 5'd15, 27'h0000014c, 32'h00000400,
  1'd1,  5'd17, 27'h00000396, 5'd12, 27'h00000280, 5'd23, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ea, 5'd25, 27'h0000003a, 5'd2, 27'h00000161, 32'h00000400,
  1'd1,  5'd18, 27'h000002dc, 5'd24, 27'h000003a8, 5'd15, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000322, 5'd21, 27'h00000235, 5'd24, 27'h0000009f, 32'h00000400,
  1'd1,  5'd28, 27'h000002da, 5'd0, 27'h0000008d, 5'd3, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001e1, 5'd1, 27'h0000002b, 5'd15, 27'h00000131, 32'h00000400,
  1'd1,  5'd26, 27'h00000222, 5'd0, 27'h00000107, 5'd21, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000050, 5'd13, 27'h000003cb, 5'd0, 27'h000003b0, 32'h00000400,
  1'd1,  5'd30, 27'h00000084, 5'd10, 27'h000003cc, 5'd11, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000075, 5'd10, 27'h00000342, 5'd25, 27'h00000319, 32'h00000400,
  1'd1,  5'd30, 27'h000003a1, 5'd21, 27'h0000014e, 5'd0, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000218, 5'd21, 27'h0000031c, 5'd12, 27'h00000189, 32'h00000400,
  1'd1,  5'd27, 27'h000001a9, 5'd25, 27'h000002a2, 5'd23, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000039b, 5'd0, 27'h00000273, 5'd1, 27'h00000157, 32'h00000400,
  1'd1,  5'd5, 27'h000000e1, 5'd2, 27'h0000013b, 5'd10, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d9, 5'd2, 27'h000000eb, 5'd21, 27'h00000216, 32'h00000400,
  1'd1,  5'd7, 27'h0000022d, 5'd14, 27'h0000026b, 5'd5, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e9, 5'd14, 27'h0000000f, 5'd17, 27'h000000ab, 32'h00000400,
  1'd1,  5'd8, 27'h00000204, 5'd12, 27'h00000216, 5'd29, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000009a, 5'd21, 27'h000003c9, 5'd6, 27'h00000147, 32'h00000400,
  1'd1,  5'd8, 27'h000002bf, 5'd23, 27'h0000029a, 5'd15, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a0, 5'd24, 27'h000003cc, 5'd27, 27'h0000016d, 32'h00000400,
  1'd1,  5'd17, 27'h0000035b, 5'd0, 27'h00000155, 5'd5, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003ab, 5'd0, 27'h00000393, 5'd11, 27'h0000021a, 32'h00000400,
  1'd1,  5'd18, 27'h00000163, 5'd1, 27'h00000078, 5'd24, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000345, 5'd14, 27'h000003c6, 5'd5, 27'h00000106, 32'h00000400,
  1'd1,  5'd15, 27'h00000398, 5'd14, 27'h0000001f, 5'd18, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000f0, 5'd13, 27'h000000b2, 5'd26, 27'h00000308, 32'h00000400,
  1'd1,  5'd19, 27'h000003b5, 5'd25, 27'h000001e6, 5'd8, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000df, 5'd25, 27'h00000000, 5'd20, 27'h00000136, 32'h00000400,
  1'd1,  5'd17, 27'h0000012b, 5'd25, 27'h00000311, 5'd28, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001ca, 5'd1, 27'h000002ff, 5'd7, 27'h000001f3, 32'h00000400,
  1'd1,  5'd30, 27'h00000322, 5'd3, 27'h00000309, 5'd19, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000248, 5'd4, 27'h000002cf, 5'd30, 27'h00000053, 32'h00000400,
  1'd1,  5'd26, 27'h000002df, 5'd13, 27'h00000132, 5'd10, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000382, 5'd14, 27'h00000296, 5'd19, 27'h0000015f, 32'h00000400,
  1'd1,  5'd28, 27'h000003eb, 5'd15, 27'h00000109, 5'd30, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e8, 5'd24, 27'h0000025b, 5'd6, 27'h000002bf, 32'h00000400,
  1'd1,  5'd26, 27'h0000024c, 5'd21, 27'h000003bd, 5'd19, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000098, 5'd21, 27'h0000011e, 5'd26, 27'h00000396, 32'h00000400,
  1'd1,  5'd5, 27'h00000327, 5'd5, 27'h0000015c, 5'd0, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012e, 5'd5, 27'h00000186, 5'd14, 27'h00000329, 32'h00000400,
  1'd1,  5'd9, 27'h00000286, 5'd5, 27'h000002db, 5'd21, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000196, 5'd19, 27'h0000024f, 5'd1, 27'h00000358, 32'h00000400,
  1'd1,  5'd8, 27'h0000039c, 5'd15, 27'h000002bb, 5'd11, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c9, 5'd19, 27'h0000002b, 5'd24, 27'h000001a7, 32'h00000400,
  1'd1,  5'd8, 27'h000002ff, 5'd29, 27'h000003b3, 5'd3, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000018c, 5'd26, 27'h0000018c, 5'd14, 27'h00000267, 32'h00000400,
  1'd1,  5'd9, 27'h0000018d, 5'd30, 27'h00000246, 5'd23, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000024e, 5'd6, 27'h00000216, 5'd0, 27'h00000229, 32'h00000400,
  1'd1,  5'd18, 27'h000002c9, 5'd9, 27'h000002ad, 5'd15, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000024f, 5'd8, 27'h000001d1, 5'd24, 27'h0000039f, 32'h00000400,
  1'd1,  5'd20, 27'h0000000a, 5'd17, 27'h000003d6, 5'd4, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000b1, 5'd19, 27'h00000267, 5'd13, 27'h0000019b, 32'h00000400,
  1'd1,  5'd17, 27'h000003a7, 5'd18, 27'h000000c3, 5'd21, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000309, 5'd27, 27'h00000160, 5'd3, 27'h0000008a, 32'h00000400,
  1'd1,  5'd17, 27'h000000d4, 5'd26, 27'h000002c4, 5'd15, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032d, 5'd30, 27'h000002f2, 5'd24, 27'h0000034e, 32'h00000400,
  1'd1,  5'd27, 27'h000000f0, 5'd7, 27'h00000170, 5'd4, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000212, 5'd10, 27'h0000003b, 5'd15, 27'h00000078, 32'h00000400,
  1'd1,  5'd28, 27'h00000385, 5'd7, 27'h000001af, 5'd20, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000386, 5'd19, 27'h000000b5, 5'd4, 27'h000003f4, 32'h00000400,
  1'd1,  5'd26, 27'h0000002a, 5'd20, 27'h00000207, 5'd14, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d6, 5'd17, 27'h00000043, 5'd21, 27'h00000133, 32'h00000400,
  1'd1,  5'd27, 27'h00000289, 5'd27, 27'h00000063, 5'd0, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a9, 5'd30, 27'h000002fa, 5'd15, 27'h00000086, 32'h00000400,
  1'd1,  5'd28, 27'h0000013b, 5'd26, 27'h0000013e, 5'd25, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000029e, 5'd9, 27'h0000011d, 5'd8, 27'h00000005, 32'h00000400,
  1'd1,  5'd8, 27'h00000017, 5'd10, 27'h000000f8, 5'd18, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f3, 5'd7, 27'h000001b8, 5'd29, 27'h000002ad, 32'h00000400,
  1'd1,  5'd7, 27'h00000277, 5'd18, 27'h0000033c, 5'd9, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b5, 5'd20, 27'h00000257, 5'd20, 27'h0000017a, 32'h00000400,
  1'd1,  5'd9, 27'h000003d1, 5'd19, 27'h000003d4, 5'd26, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000362, 5'd27, 27'h00000244, 5'd5, 27'h00000199, 32'h00000400,
  1'd1,  5'd9, 27'h000003a4, 5'd30, 27'h0000012d, 5'd16, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000135, 5'd29, 27'h00000324, 5'd27, 27'h00000386, 32'h00000400,
  1'd1,  5'd20, 27'h000001c7, 5'd7, 27'h0000031e, 5'd8, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006a, 5'd6, 27'h00000225, 5'd17, 27'h00000354, 32'h00000400,
  1'd1,  5'd18, 27'h0000029a, 5'd9, 27'h00000200, 5'd26, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000005, 5'd18, 27'h0000016c, 5'd8, 27'h000002fa, 32'h00000400,
  1'd1,  5'd15, 27'h000002d6, 5'd19, 27'h00000268, 5'd20, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000012c, 5'd20, 27'h00000208, 5'd26, 27'h0000025f, 32'h00000400,
  1'd1,  5'd17, 27'h00000253, 5'd29, 27'h0000036c, 5'd8, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000345, 5'd26, 27'h0000006f, 5'd18, 27'h000002b1, 32'h00000400,
  1'd1,  5'd19, 27'h0000025f, 5'd28, 27'h00000218, 5'd29, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000033c, 5'd6, 27'h000000f5, 5'd8, 27'h00000137, 32'h00000400,
  1'd1,  5'd30, 27'h0000035f, 5'd7, 27'h00000268, 5'd16, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021d, 5'd8, 27'h0000037f, 5'd26, 27'h00000371, 32'h00000400,
  1'd1,  5'd28, 27'h00000330, 5'd16, 27'h0000036b, 5'd8, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000201, 5'd16, 27'h0000018e, 5'd20, 27'h00000028, 32'h00000400,
  1'd1,  5'd29, 27'h00000160, 5'd18, 27'h00000209, 5'd27, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003c4, 5'd27, 27'h0000016e, 5'd7, 27'h000002c2, 32'h00000400,
  1'd1,  5'd29, 27'h0000000d, 5'd27, 27'h000000ac, 5'd19, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000057, 5'd30, 27'h0000016c, 5'd27, 27'h00000153, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h0000001e, 5'd2, 27'h00000045, 5'd2, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028c, 5'd4, 27'h00000155, 5'd13, 27'h00000059, 32'h00000400,
  1'd1,  5'd4, 27'h000002c5, 5'd2, 27'h000003f5, 5'd22, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000029e, 5'd14, 27'h000003a2, 5'd0, 27'h000000d6, 32'h00000400,
  1'd1,  5'd2, 27'h000002d5, 5'd14, 27'h00000154, 5'd13, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003df, 5'd11, 27'h0000022b, 5'd22, 27'h000003d5, 32'h00000400,
  1'd1,  5'd2, 27'h00000300, 5'd23, 27'h00000356, 5'd2, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000059, 5'd24, 27'h00000261, 5'd12, 27'h00000320, 32'h00000400,
  1'd1,  5'd3, 27'h0000037c, 5'd20, 27'h0000033a, 5'd22, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029c, 5'd3, 27'h000000c3, 5'd3, 27'h0000030b, 32'h00000400,
  1'd1,  5'd13, 27'h0000005a, 5'd0, 27'h0000023d, 5'd13, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000270, 5'd5, 27'h00000088, 5'd23, 27'h000002ad, 32'h00000400,
  1'd1,  5'd10, 27'h0000033b, 5'd14, 27'h00000052, 5'd1, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002b9, 5'd11, 27'h000002e0, 5'd13, 27'h00000353, 32'h00000400,
  1'd1,  5'd12, 27'h0000011f, 5'd10, 27'h00000395, 5'd25, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000fd, 5'd24, 27'h0000025b, 5'd1, 27'h000001a6, 32'h00000400,
  1'd1,  5'd10, 27'h00000298, 5'd21, 27'h0000031c, 5'd13, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c0, 5'd25, 27'h0000028e, 5'd25, 27'h000001a3, 32'h00000400,
  1'd1,  5'd24, 27'h000002a4, 5'd4, 27'h000001a9, 5'd3, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d0, 5'd2, 27'h000002ea, 5'd13, 27'h00000225, 32'h00000400,
  1'd1,  5'd24, 27'h000003f1, 5'd4, 27'h0000000a, 5'd21, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d2, 5'd14, 27'h00000130, 5'd0, 27'h000003e5, 32'h00000400,
  1'd1,  5'd24, 27'h000001fe, 5'd12, 27'h00000122, 5'd12, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003a2, 5'd14, 27'h0000024d, 5'd24, 27'h0000011b, 32'h00000400,
  1'd1,  5'd21, 27'h00000097, 5'd21, 27'h00000101, 5'd1, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000081, 5'd23, 27'h00000307, 5'd14, 27'h00000282, 32'h00000400,
  1'd1,  5'd23, 27'h000003be, 5'd21, 27'h000001f3, 5'd23, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f2, 5'd2, 27'h0000008f, 5'd7, 27'h0000033e, 32'h00000400,
  1'd1,  5'd2, 27'h000002c4, 5'd1, 27'h0000009a, 5'd19, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ff, 5'd4, 27'h00000117, 5'd28, 27'h000003cb, 32'h00000400,
  1'd1,  5'd4, 27'h000000c5, 5'd13, 27'h000001fa, 5'd7, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000082, 5'd13, 27'h000000ff, 5'd16, 27'h0000000d, 32'h00000400,
  1'd1,  5'd2, 27'h00000258, 5'd11, 27'h000003d7, 5'd28, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002c4, 5'd24, 27'h000002ce, 5'd8, 27'h0000003b, 32'h00000400,
  1'd1,  5'd3, 27'h000001c3, 5'd22, 27'h00000275, 5'd17, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000184, 5'd25, 27'h0000013b, 5'd25, 27'h000003d6, 32'h00000400,
  1'd1,  5'd11, 27'h0000009c, 5'd4, 27'h00000244, 5'd9, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b9, 5'd2, 27'h00000310, 5'd16, 27'h0000035b, 32'h00000400,
  1'd1,  5'd13, 27'h000000b2, 5'd4, 27'h00000378, 5'd26, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000179, 5'd12, 27'h00000298, 5'd5, 27'h00000215, 32'h00000400,
  1'd1,  5'd12, 27'h00000366, 5'd12, 27'h000001b0, 5'd18, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000193, 5'd13, 27'h000000ff, 5'd29, 27'h0000002c, 32'h00000400,
  1'd1,  5'd13, 27'h00000001, 5'd25, 27'h00000294, 5'd8, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021c, 5'd25, 27'h000001d3, 5'd16, 27'h000002e9, 32'h00000400,
  1'd1,  5'd10, 27'h0000021b, 5'd25, 27'h000002be, 5'd26, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003aa, 5'd0, 27'h00000211, 5'd9, 27'h00000108, 32'h00000400,
  1'd1,  5'd21, 27'h000003ef, 5'd2, 27'h00000339, 5'd18, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019c, 5'd3, 27'h00000193, 5'd26, 27'h000001a0, 32'h00000400,
  1'd1,  5'd24, 27'h0000034b, 5'd10, 27'h000001e8, 5'd6, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a7, 5'd15, 27'h000001db, 5'd18, 27'h000001e5, 32'h00000400,
  1'd1,  5'd25, 27'h00000171, 5'd15, 27'h000000d8, 5'd26, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000003e, 5'd22, 27'h0000036e, 5'd6, 27'h0000036a, 32'h00000400,
  1'd1,  5'd23, 27'h000003cb, 5'd23, 27'h00000264, 5'd19, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000038a, 5'd21, 27'h000003ba, 5'd27, 27'h00000170, 32'h00000400,
  1'd1,  5'd0, 27'h000002de, 5'd8, 27'h0000016c, 5'd4, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d9, 5'd7, 27'h000002b8, 5'd15, 27'h00000121, 32'h00000400,
  1'd1,  5'd4, 27'h000000a9, 5'd9, 27'h00000398, 5'd22, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000140, 5'd18, 27'h000002da, 5'd0, 27'h00000340, 32'h00000400,
  1'd1,  5'd2, 27'h000003fd, 5'd16, 27'h00000134, 5'd11, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000392, 5'd16, 27'h00000022, 5'd22, 27'h000003ec, 32'h00000400,
  1'd1,  5'd0, 27'h00000019, 5'd29, 27'h00000317, 5'd0, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000026b, 5'd27, 27'h000000df, 5'd10, 27'h00000312, 32'h00000400,
  1'd1,  5'd1, 27'h000000e3, 5'd28, 27'h000001c4, 5'd25, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000036d, 5'd5, 27'h000001ad, 5'd1, 27'h0000035e, 32'h00000400,
  1'd1,  5'd14, 27'h0000015b, 5'd5, 27'h000000d1, 5'd14, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000009c, 5'd9, 27'h0000012d, 5'd24, 27'h000001ef, 32'h00000400,
  1'd1,  5'd15, 27'h00000181, 5'd18, 27'h00000239, 5'd4, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000005, 5'd19, 27'h000001c0, 5'd11, 27'h0000022f, 32'h00000400,
  1'd1,  5'd13, 27'h000003ff, 5'd18, 27'h000000b2, 5'd23, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000023, 5'd25, 27'h000003f4, 5'd4, 27'h000002e7, 32'h00000400,
  1'd1,  5'd13, 27'h000003ba, 5'd28, 27'h0000036b, 5'd11, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000210, 5'd26, 27'h00000226, 5'd25, 27'h00000210, 32'h00000400,
  1'd1,  5'd24, 27'h00000037, 5'd8, 27'h000001be, 5'd1, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000014f, 5'd7, 27'h0000002e, 5'd11, 27'h00000113, 32'h00000400,
  1'd1,  5'd23, 27'h0000010e, 5'd5, 27'h000002ca, 5'd23, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000311, 5'd16, 27'h000000e8, 5'd4, 27'h00000075, 32'h00000400,
  1'd1,  5'd25, 27'h0000017d, 5'd16, 27'h0000016e, 5'd15, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001f9, 5'd20, 27'h000000b1, 5'd21, 27'h000003fb, 32'h00000400,
  1'd1,  5'd23, 27'h000003ac, 5'd28, 27'h000002cd, 5'd3, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000014e, 5'd27, 27'h00000158, 5'd14, 27'h0000037a, 32'h00000400,
  1'd1,  5'd21, 27'h000003a4, 5'd26, 27'h000003cc, 5'd20, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000018f, 5'd9, 27'h00000336, 5'd5, 27'h000002f5, 32'h00000400,
  1'd1,  5'd3, 27'h00000284, 5'd7, 27'h00000018, 5'd15, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000355, 5'd9, 27'h0000000f, 5'd28, 27'h00000052, 32'h00000400,
  1'd1,  5'd3, 27'h000000c2, 5'd20, 27'h000000e3, 5'd6, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000038a, 5'd16, 27'h00000355, 5'd17, 27'h00000381, 32'h00000400,
  1'd1,  5'd3, 27'h00000257, 5'd16, 27'h00000190, 5'd28, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000165, 5'd30, 27'h00000382, 5'd7, 27'h000000b4, 32'h00000400,
  1'd1,  5'd0, 27'h00000057, 5'd28, 27'h000002a9, 5'd18, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000cd, 5'd29, 27'h000000be, 5'd27, 27'h00000022, 32'h00000400,
  1'd1,  5'd12, 27'h0000002b, 5'd9, 27'h00000248, 5'd8, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000006b, 5'd8, 27'h000001fb, 5'd19, 27'h000001a7, 32'h00000400,
  1'd1,  5'd11, 27'h000000bd, 5'd7, 27'h000003e4, 5'd28, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000266, 5'd15, 27'h00000252, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd14, 27'h000003fa, 5'd19, 27'h00000035, 5'd17, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000238, 5'd16, 27'h000002ca, 5'd26, 27'h000002b6, 32'h00000400,
  1'd1,  5'd11, 27'h00000073, 5'd29, 27'h00000195, 5'd7, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000009a, 5'd29, 27'h00000240, 5'd15, 27'h0000030c, 32'h00000400,
  1'd1,  5'd10, 27'h00000272, 5'd29, 27'h00000045, 5'd30, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000cb, 5'd6, 27'h00000044, 5'd9, 27'h00000373, 32'h00000400,
  1'd1,  5'd23, 27'h00000288, 5'd7, 27'h00000098, 5'd20, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001d6, 5'd8, 27'h00000211, 5'd30, 27'h000000bd, 32'h00000400,
  1'd1,  5'd22, 27'h000002db, 5'd17, 27'h00000069, 5'd7, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ed, 5'd16, 27'h0000035e, 5'd17, 27'h00000006, 32'h00000400,
  1'd1,  5'd23, 27'h000000a0, 5'd18, 27'h00000270, 5'd26, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000fc, 5'd28, 27'h00000182, 5'd8, 27'h000001ea, 32'h00000400,
  1'd1,  5'd25, 27'h0000000a, 5'd28, 27'h000000e0, 5'd15, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000187, 5'd30, 27'h0000002a, 5'd30, 27'h00000060, 32'h00000400,
  1'd1,  5'd8, 27'h00000198, 5'd2, 27'h00000329, 5'd6, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000033a, 5'd0, 27'h000003b2, 5'd20, 27'h00000011, 32'h00000400,
  1'd1,  5'd9, 27'h00000025, 5'd2, 27'h00000101, 5'd30, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000074, 5'd11, 27'h00000343, 5'd1, 27'h00000298, 32'h00000400,
  1'd1,  5'd5, 27'h00000325, 5'd13, 27'h00000152, 5'd15, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001e1, 5'd11, 27'h00000197, 5'd25, 27'h00000155, 32'h00000400,
  1'd1,  5'd8, 27'h000001ac, 5'd23, 27'h00000344, 5'd3, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000010f, 5'd25, 27'h000002f9, 5'd14, 27'h0000015e, 32'h00000400,
  1'd1,  5'd9, 27'h00000106, 5'd23, 27'h00000105, 5'd25, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e1, 5'd3, 27'h00000322, 5'd6, 27'h000002ad, 32'h00000400,
  1'd1,  5'd19, 27'h00000126, 5'd2, 27'h00000251, 5'd19, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030a, 5'd4, 27'h00000393, 5'd27, 27'h000002f4, 32'h00000400,
  1'd1,  5'd17, 27'h000001b5, 5'd11, 27'h000003cf, 5'd4, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e8, 5'd15, 27'h000000b5, 5'd14, 27'h0000003f, 32'h00000400,
  1'd1,  5'd18, 27'h00000230, 5'd12, 27'h000001cd, 5'd23, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002d6, 5'd24, 27'h00000343, 5'd4, 27'h000002df, 32'h00000400,
  1'd1,  5'd16, 27'h00000062, 5'd24, 27'h000000d1, 5'd13, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ad, 5'd23, 27'h00000343, 5'd23, 27'h00000332, 32'h00000400,
  1'd1,  5'd28, 27'h00000018, 5'd4, 27'h0000005d, 5'd4, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023c, 5'd3, 27'h00000273, 5'd13, 27'h00000253, 32'h00000400,
  1'd1,  5'd29, 27'h000001f1, 5'd0, 27'h00000159, 5'd23, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000028c, 5'd10, 27'h00000363, 5'd0, 27'h000003bc, 32'h00000400,
  1'd1,  5'd30, 27'h000001cd, 5'd12, 27'h0000030b, 5'd11, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000180, 5'd10, 27'h00000356, 5'd21, 27'h0000033f, 32'h00000400,
  1'd1,  5'd28, 27'h00000222, 5'd23, 27'h0000006d, 5'd3, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000365, 5'd22, 27'h000000b3, 5'd15, 27'h000000fb, 32'h00000400,
  1'd1,  5'd30, 27'h00000285, 5'd22, 27'h000003d5, 5'd23, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000356, 5'd0, 27'h00000122, 5'd2, 27'h000000cd, 32'h00000400,
  1'd1,  5'd9, 27'h0000039f, 5'd1, 27'h000002ad, 5'd12, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000018, 5'd0, 27'h0000036d, 5'd21, 27'h00000282, 32'h00000400,
  1'd1,  5'd6, 27'h00000286, 5'd15, 27'h00000087, 5'd5, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ab, 5'd11, 27'h0000001b, 5'd16, 27'h0000024d, 32'h00000400,
  1'd1,  5'd7, 27'h00000024, 5'd13, 27'h0000003c, 5'd27, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000238, 5'd21, 27'h000003be, 5'd5, 27'h00000135, 32'h00000400,
  1'd1,  5'd7, 27'h000002ca, 5'd25, 27'h0000026a, 5'd20, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000379, 5'd22, 27'h00000200, 5'd26, 27'h00000146, 32'h00000400,
  1'd1,  5'd15, 27'h00000202, 5'd4, 27'h000000c0, 5'd0, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000005b, 5'd3, 27'h00000115, 5'd14, 27'h000002ad, 32'h00000400,
  1'd1,  5'd18, 27'h0000006b, 5'd4, 27'h000001ae, 5'd21, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000125, 5'd14, 27'h000003c8, 5'd7, 27'h0000039e, 32'h00000400,
  1'd1,  5'd19, 27'h00000353, 5'd11, 27'h00000245, 5'd19, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000103, 5'd10, 27'h00000283, 5'd29, 27'h00000017, 32'h00000400,
  1'd1,  5'd20, 27'h000001f1, 5'd22, 27'h0000018b, 5'd5, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000366, 5'd23, 27'h000002df, 5'd19, 27'h000000f0, 32'h00000400,
  1'd1,  5'd20, 27'h000000ac, 5'd24, 27'h00000178, 5'd26, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000185, 5'd3, 27'h0000039c, 5'd7, 27'h00000176, 32'h00000400,
  1'd1,  5'd30, 27'h00000381, 5'd0, 27'h0000007b, 5'd17, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000241, 5'd4, 27'h0000024b, 5'd26, 27'h000001af, 32'h00000400,
  1'd1,  5'd29, 27'h00000358, 5'd11, 27'h000003f6, 5'd5, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c4, 5'd14, 27'h000003e2, 5'd18, 27'h00000379, 32'h00000400,
  1'd1,  5'd27, 27'h0000011f, 5'd11, 27'h00000095, 5'd30, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025b, 5'd24, 27'h000002bc, 5'd7, 27'h000001a1, 32'h00000400,
  1'd1,  5'd26, 27'h0000029f, 5'd21, 27'h00000121, 5'd17, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d0, 5'd23, 27'h00000396, 5'd30, 27'h000000c0, 32'h00000400,
  1'd1,  5'd9, 27'h000001e1, 5'd9, 27'h00000395, 5'd4, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000104, 5'd6, 27'h000002a7, 5'd14, 27'h0000030d, 32'h00000400,
  1'd1,  5'd6, 27'h0000008a, 5'd9, 27'h00000365, 5'd22, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000013, 5'd16, 27'h000002da, 5'd0, 27'h00000252, 32'h00000400,
  1'd1,  5'd5, 27'h000000bf, 5'd17, 27'h000001b8, 5'd13, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032e, 5'd20, 27'h00000145, 5'd21, 27'h00000055, 32'h00000400,
  1'd1,  5'd9, 27'h00000167, 5'd28, 27'h00000317, 5'd4, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005c, 5'd29, 27'h00000331, 5'd11, 27'h00000227, 32'h00000400,
  1'd1,  5'd8, 27'h00000183, 5'd25, 27'h0000035c, 5'd21, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000172, 5'd10, 27'h000000e3, 5'd0, 27'h00000286, 32'h00000400,
  1'd1,  5'd16, 27'h0000038b, 5'd5, 27'h00000215, 5'd14, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000021, 5'd9, 27'h0000015e, 5'd21, 27'h00000085, 32'h00000400,
  1'd1,  5'd19, 27'h000001b1, 5'd16, 27'h000002c7, 5'd1, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000016c, 5'd17, 27'h000003d7, 5'd14, 27'h0000011a, 32'h00000400,
  1'd1,  5'd17, 27'h000000a3, 5'd19, 27'h000001be, 5'd21, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000082, 5'd30, 27'h000000a6, 5'd4, 27'h000002d5, 32'h00000400,
  1'd1,  5'd17, 27'h00000371, 5'd30, 27'h00000154, 5'd13, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000008e, 5'd26, 27'h000002bf, 5'd25, 27'h000000d1, 32'h00000400,
  1'd1,  5'd30, 27'h00000063, 5'd7, 27'h000003bf, 5'd1, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e1, 5'd9, 27'h000003ff, 5'd12, 27'h00000275, 32'h00000400,
  1'd1,  5'd29, 27'h00000071, 5'd6, 27'h0000012d, 5'd22, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000e4, 5'd20, 27'h0000004f, 5'd0, 27'h0000026f, 32'h00000400,
  1'd1,  5'd28, 27'h00000370, 5'd20, 27'h00000295, 5'd11, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000172, 5'd19, 27'h00000364, 5'd25, 27'h00000171, 32'h00000400,
  1'd1,  5'd30, 27'h0000033e, 5'd29, 27'h0000009a, 5'd0, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d4, 5'd28, 27'h000000d7, 5'd11, 27'h00000259, 32'h00000400,
  1'd1,  5'd27, 27'h0000006b, 5'd30, 27'h000001c1, 5'd23, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c0, 5'd7, 27'h000000b6, 5'd8, 27'h00000097, 32'h00000400,
  1'd1,  5'd9, 27'h00000216, 5'd6, 27'h000001c3, 5'd19, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001a3, 5'd5, 27'h00000208, 5'd26, 27'h0000005e, 32'h00000400,
  1'd1,  5'd10, 27'h00000088, 5'd17, 27'h000000e8, 5'd9, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a6, 5'd20, 27'h00000005, 5'd18, 27'h00000344, 32'h00000400,
  1'd1,  5'd7, 27'h00000229, 5'd19, 27'h00000038, 5'd28, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d0, 5'd26, 27'h00000166, 5'd7, 27'h00000372, 32'h00000400,
  1'd1,  5'd6, 27'h0000021a, 5'd30, 27'h000001f8, 5'd17, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003f5, 5'd28, 27'h000000c8, 5'd27, 27'h000001aa, 32'h00000400,
  1'd1,  5'd16, 27'h00000352, 5'd5, 27'h000003ad, 5'd7, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d3, 5'd6, 27'h0000000a, 5'd17, 27'h000000a3, 32'h00000400,
  1'd1,  5'd16, 27'h000002ec, 5'd5, 27'h000003c7, 5'd30, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000009b, 5'd19, 27'h000001c4, 5'd7, 27'h0000023e, 32'h00000400,
  1'd1,  5'd17, 27'h000002c6, 5'd16, 27'h000000c7, 5'd17, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b3, 5'd20, 27'h00000280, 5'd27, 27'h00000037, 32'h00000400,
  1'd1,  5'd15, 27'h000002c7, 5'd26, 27'h000002dd, 5'd6, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000358, 5'd25, 27'h00000386, 5'd20, 27'h00000160, 32'h00000400,
  1'd1,  5'd17, 27'h00000041, 5'd26, 27'h00000218, 5'd26, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000027, 5'd5, 27'h000003e9, 5'd7, 27'h000001ab, 32'h00000400,
  1'd1,  5'd27, 27'h00000385, 5'd6, 27'h0000002f, 5'd16, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000278, 5'd9, 27'h000003f0, 5'd29, 27'h000003e8, 32'h00000400,
  1'd1,  5'd27, 27'h00000165, 5'd16, 27'h00000233, 5'd8, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000164, 5'd20, 27'h00000062, 5'd18, 27'h000002e4, 32'h00000400,
  1'd1,  5'd27, 27'h00000130, 5'd18, 27'h00000204, 5'd26, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001ed, 5'd29, 27'h0000008c, 5'd10, 27'h00000135, 32'h00000400,
  1'd1,  5'd27, 27'h00000234, 5'd29, 27'h00000146, 5'd16, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000143, 5'd28, 27'h0000006a, 5'd26, 27'h000003c4, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h0000026c, 5'd3, 27'h0000036f, 5'd3, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003bb, 5'd2, 27'h00000231, 5'd13, 27'h000001d0, 32'h00000400,
  1'd1,  5'd2, 27'h00000262, 5'd3, 27'h00000205, 5'd21, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000002, 5'd12, 27'h000001b0, 5'd3, 27'h0000011e, 32'h00000400,
  1'd1,  5'd0, 27'h0000014a, 5'd10, 27'h00000218, 5'd12, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000390, 5'd14, 27'h0000027b, 5'd20, 27'h0000033c, 32'h00000400,
  1'd1,  5'd0, 27'h00000290, 5'd23, 27'h00000197, 5'd1, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000249, 5'd24, 27'h000000b1, 5'd14, 27'h00000184, 32'h00000400,
  1'd1,  5'd1, 27'h0000031f, 5'd25, 27'h000000c1, 5'd22, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000246, 5'd4, 27'h0000008d, 5'd2, 27'h000000ee, 32'h00000400,
  1'd1,  5'd13, 27'h0000027f, 5'd2, 27'h0000013c, 5'd12, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017d, 5'd3, 27'h00000093, 5'd21, 27'h000002bf, 32'h00000400,
  1'd1,  5'd11, 27'h00000117, 5'd15, 27'h0000002a, 5'd0, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b4, 5'd12, 27'h0000007c, 5'd14, 27'h00000245, 32'h00000400,
  1'd1,  5'd15, 27'h00000184, 5'd11, 27'h000002f8, 5'd23, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000158, 5'd24, 27'h0000007a, 5'd3, 27'h000003f4, 32'h00000400,
  1'd1,  5'd11, 27'h0000013a, 5'd21, 27'h0000010f, 5'd11, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001b9, 5'd25, 27'h0000001c, 5'd23, 27'h0000030c, 32'h00000400,
  1'd1,  5'd21, 27'h0000036e, 5'd2, 27'h0000014c, 5'd1, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ef, 5'd3, 27'h000003c0, 5'd11, 27'h000002e0, 32'h00000400,
  1'd1,  5'd24, 27'h000003e3, 5'd5, 27'h00000014, 5'd25, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000118, 5'd15, 27'h00000186, 5'd2, 27'h000003ec, 32'h00000400,
  1'd1,  5'd25, 27'h00000309, 5'd14, 27'h00000293, 5'd14, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034b, 5'd13, 27'h000001f4, 5'd22, 27'h000003c9, 32'h00000400,
  1'd1,  5'd23, 27'h000003de, 5'd23, 27'h0000010c, 5'd1, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000398, 5'd21, 27'h000001e2, 5'd12, 27'h0000037f, 32'h00000400,
  1'd1,  5'd23, 27'h00000059, 5'd20, 27'h000003bb, 5'd21, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f5, 5'd0, 27'h0000014d, 5'd6, 27'h000001a2, 32'h00000400,
  1'd1,  5'd3, 27'h00000082, 5'd0, 27'h000001f4, 5'd19, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005b, 5'd2, 27'h000001de, 5'd28, 27'h000002b5, 32'h00000400,
  1'd1,  5'd3, 27'h0000020b, 5'd11, 27'h0000001d, 5'd6, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000c9, 5'd15, 27'h00000143, 5'd15, 27'h000002e1, 32'h00000400,
  1'd1,  5'd4, 27'h00000246, 5'd15, 27'h00000075, 5'd26, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e4, 5'd23, 27'h000003ff, 5'd7, 27'h0000039c, 32'h00000400,
  1'd1,  5'd2, 27'h0000026d, 5'd25, 27'h0000020f, 5'd17, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000023b, 5'd22, 27'h00000101, 5'd30, 27'h000002ab, 32'h00000400,
  1'd1,  5'd11, 27'h00000225, 5'd2, 27'h000002bf, 5'd5, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003dc, 5'd2, 27'h000000e9, 5'd20, 27'h000001f5, 32'h00000400,
  1'd1,  5'd13, 27'h0000000b, 5'd4, 27'h000000fc, 5'd30, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002c7, 5'd13, 27'h00000371, 5'd9, 27'h000000d0, 32'h00000400,
  1'd1,  5'd13, 27'h0000012a, 5'd13, 27'h0000036c, 5'd15, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000399, 5'd15, 27'h00000067, 5'd28, 27'h00000343, 32'h00000400,
  1'd1,  5'd12, 27'h0000006e, 5'd25, 27'h00000102, 5'd6, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000003e, 5'd25, 27'h00000062, 5'd19, 27'h000000b8, 32'h00000400,
  1'd1,  5'd14, 27'h00000306, 5'd22, 27'h000000cb, 5'd30, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000016b, 5'd1, 27'h000002d7, 5'd8, 27'h0000001d, 32'h00000400,
  1'd1,  5'd21, 27'h000003d0, 5'd0, 27'h00000321, 5'd16, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ed, 5'd0, 27'h0000039e, 5'd27, 27'h00000149, 32'h00000400,
  1'd1,  5'd23, 27'h000003aa, 5'd11, 27'h000002b0, 5'd5, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e0, 5'd12, 27'h00000206, 5'd16, 27'h000003b5, 32'h00000400,
  1'd1,  5'd25, 27'h0000027f, 5'd13, 27'h00000218, 5'd30, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000008e, 5'd21, 27'h00000016, 5'd8, 27'h0000032f, 32'h00000400,
  1'd1,  5'd22, 27'h0000031a, 5'd22, 27'h00000315, 5'd19, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f6, 5'd23, 27'h0000007c, 5'd27, 27'h00000023, 32'h00000400,
  1'd1,  5'd2, 27'h00000044, 5'd5, 27'h0000018d, 5'd0, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003fe, 5'd8, 27'h000003d9, 5'd13, 27'h00000225, 32'h00000400,
  1'd1,  5'd3, 27'h00000243, 5'd9, 27'h000000a4, 5'd25, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032b, 5'd17, 27'h00000314, 5'd0, 27'h00000259, 32'h00000400,
  1'd1,  5'd4, 27'h00000387, 5'd18, 27'h00000176, 5'd12, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000378, 5'd18, 27'h00000200, 5'd23, 27'h00000080, 32'h00000400,
  1'd1,  5'd3, 27'h00000190, 5'd27, 27'h00000264, 5'd3, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000009, 5'd29, 27'h000003ff, 5'd14, 27'h000003f7, 32'h00000400,
  1'd1,  5'd0, 27'h00000185, 5'd29, 27'h0000008e, 5'd23, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000290, 5'd7, 27'h000001a2, 5'd2, 27'h0000039b, 32'h00000400,
  1'd1,  5'd12, 27'h0000011f, 5'd6, 27'h0000006b, 5'd13, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c3, 5'd7, 27'h000001d0, 5'd21, 27'h00000077, 32'h00000400,
  1'd1,  5'd10, 27'h000003a2, 5'd16, 27'h000000a1, 5'd3, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000001f, 5'd16, 27'h000001aa, 5'd10, 27'h00000284, 32'h00000400,
  1'd1,  5'd13, 27'h000001ae, 5'd18, 27'h000000bc, 5'd22, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f0, 5'd30, 27'h0000005d, 5'd4, 27'h0000023c, 32'h00000400,
  1'd1,  5'd15, 27'h000000d4, 5'd29, 27'h00000218, 5'd14, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000027c, 5'd28, 27'h00000285, 5'd21, 27'h000000e0, 32'h00000400,
  1'd1,  5'd24, 27'h00000247, 5'd7, 27'h00000030, 5'd3, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000001, 5'd9, 27'h00000094, 5'd10, 27'h000002aa, 32'h00000400,
  1'd1,  5'd25, 27'h000002e9, 5'd8, 27'h0000004a, 5'd22, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f3, 5'd17, 27'h0000014d, 5'd1, 27'h00000196, 32'h00000400,
  1'd1,  5'd23, 27'h0000006d, 5'd17, 27'h0000008e, 5'd11, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000292, 5'd17, 27'h00000047, 5'd21, 27'h00000379, 32'h00000400,
  1'd1,  5'd22, 27'h00000201, 5'd30, 27'h00000156, 5'd2, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001d4, 5'd29, 27'h00000378, 5'd12, 27'h00000215, 32'h00000400,
  1'd1,  5'd23, 27'h00000061, 5'd28, 27'h0000008c, 5'd23, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ce, 5'd7, 27'h000002a4, 5'd9, 27'h00000269, 32'h00000400,
  1'd1,  5'd3, 27'h0000010f, 5'd6, 27'h00000339, 5'd16, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000086, 5'd9, 27'h00000268, 5'd30, 27'h000000f0, 32'h00000400,
  1'd1,  5'd0, 27'h000001eb, 5'd18, 27'h00000282, 5'd7, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020b, 5'd17, 27'h0000019c, 5'd18, 27'h000003be, 32'h00000400,
  1'd1,  5'd2, 27'h00000361, 5'd18, 27'h000000e0, 5'd29, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000076, 5'd27, 27'h0000011d, 5'd10, 27'h000000aa, 32'h00000400,
  1'd1,  5'd4, 27'h000002e5, 5'd30, 27'h000002f1, 5'd16, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000004c, 5'd25, 27'h000003f0, 5'd29, 27'h000002b7, 32'h00000400,
  1'd1,  5'd11, 27'h0000020b, 5'd6, 27'h00000204, 5'd8, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000318, 5'd8, 27'h000002af, 5'd15, 27'h00000384, 32'h00000400,
  1'd1,  5'd14, 27'h000001f3, 5'd7, 27'h000002c5, 5'd26, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000017e, 5'd18, 27'h000002cc, 5'd6, 27'h00000194, 32'h00000400,
  1'd1,  5'd13, 27'h00000022, 5'd19, 27'h00000257, 5'd17, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b5, 5'd17, 27'h00000288, 5'd28, 27'h000000e6, 32'h00000400,
  1'd1,  5'd13, 27'h0000020c, 5'd29, 27'h000002a5, 5'd6, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003a7, 5'd30, 27'h0000004c, 5'd18, 27'h0000027d, 32'h00000400,
  1'd1,  5'd12, 27'h00000120, 5'd25, 27'h000003a5, 5'd26, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000001, 5'd7, 27'h00000014, 5'd7, 27'h000002f4, 32'h00000400,
  1'd1,  5'd20, 27'h000003cd, 5'd6, 27'h0000008c, 5'd18, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000195, 5'd9, 27'h00000332, 5'd28, 27'h00000216, 32'h00000400,
  1'd1,  5'd23, 27'h000002b8, 5'd18, 27'h000002bd, 5'd6, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001fb, 5'd17, 27'h00000065, 5'd19, 27'h0000024c, 32'h00000400,
  1'd1,  5'd25, 27'h00000077, 5'd19, 27'h0000005e, 5'd28, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d2, 5'd27, 27'h0000025b, 5'd10, 27'h0000008f, 32'h00000400,
  1'd1,  5'd24, 27'h00000307, 5'd30, 27'h000003bc, 5'd16, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001fa, 5'd29, 27'h000001c5, 5'd28, 27'h000003a9, 32'h00000400,
  1'd1,  5'd6, 27'h00000030, 5'd4, 27'h00000339, 5'd7, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000d9, 5'd3, 27'h0000029e, 5'd17, 27'h00000268, 32'h00000400,
  1'd1,  5'd8, 27'h000003d9, 5'd0, 27'h00000349, 5'd27, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e3, 5'd13, 27'h000002be, 5'd1, 27'h00000049, 32'h00000400,
  1'd1,  5'd9, 27'h000002ab, 5'd13, 27'h00000351, 5'd14, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000229, 5'd14, 27'h0000009f, 5'd23, 27'h00000047, 32'h00000400,
  1'd1,  5'd6, 27'h00000162, 5'd24, 27'h000001db, 5'd1, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000303, 5'd23, 27'h00000220, 5'd11, 27'h000001b8, 32'h00000400,
  1'd1,  5'd5, 27'h000000e6, 5'd22, 27'h00000282, 5'd24, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000350, 5'd4, 27'h0000025e, 5'd5, 27'h00000358, 32'h00000400,
  1'd1,  5'd19, 27'h000001c5, 5'd2, 27'h000003bb, 5'd19, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000239, 5'd0, 27'h0000039c, 5'd26, 27'h00000306, 32'h00000400,
  1'd1,  5'd19, 27'h000002a2, 5'd14, 27'h00000295, 5'd2, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000160, 5'd12, 27'h000000ef, 5'd13, 27'h000001fa, 32'h00000400,
  1'd1,  5'd16, 27'h000000f9, 5'd15, 27'h00000096, 5'd21, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000014c, 5'd22, 27'h00000289, 5'd1, 27'h00000318, 32'h00000400,
  1'd1,  5'd16, 27'h000000e2, 5'd24, 27'h000001c5, 5'd12, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000367, 5'd21, 27'h00000005, 5'd25, 27'h000000c1, 32'h00000400,
  1'd1,  5'd28, 27'h000000db, 5'd2, 27'h0000015d, 5'd5, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000365, 5'd2, 27'h0000034b, 5'd13, 27'h0000025c, 32'h00000400,
  1'd1,  5'd28, 27'h000000d8, 5'd0, 27'h0000036c, 5'd25, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000330, 5'd12, 27'h000003ad, 5'd2, 27'h000000a0, 32'h00000400,
  1'd1,  5'd27, 27'h0000013d, 5'd12, 27'h000002bb, 5'd13, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001ee, 5'd14, 27'h00000205, 5'd24, 27'h00000108, 32'h00000400,
  1'd1,  5'd29, 27'h0000014d, 5'd22, 27'h000000ac, 5'd2, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002fa, 5'd20, 27'h0000031e, 5'd14, 27'h000003ee, 32'h00000400,
  1'd1,  5'd27, 27'h000001f7, 5'd21, 27'h000003f5, 5'd21, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000115, 5'd2, 27'h00000326, 5'd3, 27'h00000304, 32'h00000400,
  1'd1,  5'd9, 27'h000002c4, 5'd3, 27'h00000129, 5'd11, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000012, 5'd1, 27'h000002f5, 5'd24, 27'h00000006, 32'h00000400,
  1'd1,  5'd9, 27'h000000e9, 5'd12, 27'h00000334, 5'd6, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ce, 5'd13, 27'h0000014a, 5'd15, 27'h00000292, 32'h00000400,
  1'd1,  5'd9, 27'h0000003a, 5'd15, 27'h00000052, 5'd30, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000030, 5'd25, 27'h000000a1, 5'd8, 27'h00000239, 32'h00000400,
  1'd1,  5'd5, 27'h000002c1, 5'd22, 27'h000003fc, 5'd19, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000368, 5'd24, 27'h000002a7, 5'd30, 27'h00000318, 32'h00000400,
  1'd1,  5'd16, 27'h00000008, 5'd4, 27'h0000012e, 5'd2, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001d2, 5'd3, 27'h000002e4, 5'd12, 27'h00000169, 32'h00000400,
  1'd1,  5'd17, 27'h0000018c, 5'd5, 27'h00000055, 5'd22, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ef, 5'd12, 27'h00000323, 5'd5, 27'h0000026d, 32'h00000400,
  1'd1,  5'd16, 27'h00000090, 5'd14, 27'h0000004a, 5'd18, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000347, 5'd10, 27'h0000019e, 5'd28, 27'h00000365, 32'h00000400,
  1'd1,  5'd15, 27'h000003e7, 5'd25, 27'h00000263, 5'd10, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e5, 5'd23, 27'h000000c0, 5'd18, 27'h0000020a, 32'h00000400,
  1'd1,  5'd19, 27'h0000003c, 5'd23, 27'h0000038e, 5'd29, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a5, 5'd3, 27'h000001af, 5'd5, 27'h000003ef, 32'h00000400,
  1'd1,  5'd30, 27'h00000312, 5'd0, 27'h00000024, 5'd19, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000015f, 5'd2, 27'h00000305, 5'd27, 27'h00000299, 32'h00000400,
  1'd1,  5'd29, 27'h00000071, 5'd11, 27'h0000006d, 5'd9, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b2, 5'd14, 27'h000003d5, 5'd18, 27'h00000060, 32'h00000400,
  1'd1,  5'd28, 27'h0000007a, 5'd11, 27'h00000167, 5'd27, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ef, 5'd22, 27'h00000324, 5'd8, 27'h00000128, 32'h00000400,
  1'd1,  5'd27, 27'h00000113, 5'd24, 27'h00000390, 5'd18, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f7, 5'd21, 27'h00000353, 5'd28, 27'h00000107, 32'h00000400,
  1'd1,  5'd6, 27'h00000324, 5'd6, 27'h000000cd, 5'd0, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000039b, 5'd6, 27'h0000009e, 5'd12, 27'h00000315, 32'h00000400,
  1'd1,  5'd8, 27'h000000d6, 5'd5, 27'h0000032e, 5'd21, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000348, 5'd20, 27'h0000023a, 5'd2, 27'h00000078, 32'h00000400,
  1'd1,  5'd9, 27'h00000077, 5'd19, 27'h0000024e, 5'd12, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ec, 5'd15, 27'h0000037f, 5'd24, 27'h000001b5, 32'h00000400,
  1'd1,  5'd6, 27'h00000081, 5'd30, 27'h00000238, 5'd3, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f5, 5'd26, 27'h0000012a, 5'd12, 27'h000000f7, 32'h00000400,
  1'd1,  5'd7, 27'h0000020d, 5'd26, 27'h0000005a, 5'd23, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000004e, 5'd6, 27'h000003e2, 5'd0, 27'h0000036c, 32'h00000400,
  1'd1,  5'd16, 27'h0000031c, 5'd9, 27'h00000325, 5'd10, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035f, 5'd9, 27'h00000138, 5'd20, 27'h000003b8, 32'h00000400,
  1'd1,  5'd20, 27'h00000149, 5'd19, 27'h00000269, 5'd3, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000203, 5'd17, 27'h00000367, 5'd13, 27'h000000d2, 32'h00000400,
  1'd1,  5'd19, 27'h00000131, 5'd20, 27'h00000256, 5'd25, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034d, 5'd28, 27'h00000250, 5'd3, 27'h0000030c, 32'h00000400,
  1'd1,  5'd16, 27'h000000d5, 5'd27, 27'h000002db, 5'd10, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002eb, 5'd29, 27'h0000016b, 5'd21, 27'h00000366, 32'h00000400,
  1'd1,  5'd30, 27'h000001f2, 5'd5, 27'h000000ae, 5'd2, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017f, 5'd10, 27'h000000b3, 5'd11, 27'h000003e5, 32'h00000400,
  1'd1,  5'd29, 27'h000003b9, 5'd7, 27'h00000070, 5'd21, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000085, 5'd17, 27'h000001b4, 5'd4, 27'h000002e1, 32'h00000400,
  1'd1,  5'd28, 27'h000001cd, 5'd17, 27'h000001c2, 5'd12, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012c, 5'd15, 27'h00000299, 5'd21, 27'h00000113, 32'h00000400,
  1'd1,  5'd29, 27'h00000378, 5'd26, 27'h0000039b, 5'd4, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000039c, 5'd26, 27'h000003e0, 5'd11, 27'h000002e6, 32'h00000400,
  1'd1,  5'd29, 27'h000003bb, 5'd27, 27'h0000029e, 5'd24, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000022b, 5'd5, 27'h000002de, 5'd5, 27'h00000384, 32'h00000400,
  1'd1,  5'd6, 27'h00000084, 5'd7, 27'h000002f6, 5'd18, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e7, 5'd7, 27'h000001f4, 5'd26, 27'h0000015c, 32'h00000400,
  1'd1,  5'd10, 27'h000000dc, 5'd16, 27'h00000097, 5'd8, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003a6, 5'd15, 27'h000002f3, 5'd17, 27'h000000bc, 32'h00000400,
  1'd1,  5'd5, 27'h000001d5, 5'd16, 27'h00000314, 5'd30, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000013a, 5'd28, 27'h000001d2, 5'd5, 27'h000000c8, 32'h00000400,
  1'd1,  5'd10, 27'h00000111, 5'd25, 27'h000003d7, 5'd16, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003d8, 5'd29, 27'h0000027c, 5'd25, 27'h00000394, 32'h00000400,
  1'd1,  5'd20, 27'h0000026d, 5'd9, 27'h00000177, 5'd6, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000037c, 5'd9, 27'h000000c6, 5'd19, 27'h000002df, 32'h00000400,
  1'd1,  5'd18, 27'h000002c3, 5'd5, 27'h000001a5, 5'd27, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001cb, 5'd17, 27'h0000016a, 5'd5, 27'h00000359, 32'h00000400,
  1'd1,  5'd17, 27'h00000209, 5'd17, 27'h00000063, 5'd16, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e0, 5'd19, 27'h00000071, 5'd30, 27'h000002e5, 32'h00000400,
  1'd1,  5'd15, 27'h000002d1, 5'd30, 27'h000000d5, 5'd9, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e7, 5'd27, 27'h00000138, 5'd16, 27'h00000357, 32'h00000400,
  1'd1,  5'd19, 27'h000001e5, 5'd27, 27'h0000027a, 5'd27, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003f5, 5'd9, 27'h00000163, 5'd9, 27'h000002f1, 32'h00000400,
  1'd1,  5'd29, 27'h00000353, 5'd6, 27'h0000013c, 5'd17, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007a, 5'd7, 27'h000002fc, 5'd29, 27'h000000f7, 32'h00000400,
  1'd1,  5'd29, 27'h000000d3, 5'd15, 27'h0000025d, 5'd5, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000251, 5'd16, 27'h00000253, 5'd19, 27'h00000118, 32'h00000400,
  1'd1,  5'd30, 27'h0000017b, 5'd16, 27'h00000355, 5'd29, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000037e, 5'd26, 27'h00000022, 5'd7, 27'h00000396, 32'h00000400,
  1'd1,  5'd27, 27'h000001d8, 5'd28, 27'h000003f4, 5'd17, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c3, 5'd27, 27'h00000314, 5'd29, 27'h000002f0, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000001b0, 5'd0, 27'h000001bb, 5'd2, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002e6, 5'd3, 27'h00000123, 5'd14, 27'h000000ee, 32'h00000400,
  1'd1,  5'd0, 27'h000001e9, 5'd0, 27'h000001aa, 5'd24, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000169, 5'd10, 27'h00000246, 5'd3, 27'h000001c8, 32'h00000400,
  1'd1,  5'd0, 27'h0000017c, 5'd10, 27'h00000197, 5'd11, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000036, 5'd14, 27'h0000039a, 5'd22, 27'h000003d5, 32'h00000400,
  1'd1,  5'd2, 27'h0000026f, 5'd21, 27'h0000009b, 5'd3, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003c9, 5'd25, 27'h000000af, 5'd11, 27'h000001e9, 32'h00000400,
  1'd1,  5'd3, 27'h000003a8, 5'd22, 27'h000002ea, 5'd25, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000366, 5'd0, 27'h00000378, 5'd1, 27'h00000196, 32'h00000400,
  1'd1,  5'd11, 27'h000000c1, 5'd4, 27'h000002b7, 5'd15, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001f4, 5'd0, 27'h0000014d, 5'd20, 27'h000002d0, 32'h00000400,
  1'd1,  5'd12, 27'h0000000d, 5'd14, 27'h00000364, 5'd0, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000350, 5'd11, 27'h00000255, 5'd12, 27'h0000038b, 32'h00000400,
  1'd1,  5'd10, 27'h00000200, 5'd11, 27'h0000001a, 5'd25, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000017e, 5'd24, 27'h000002d1, 5'd2, 27'h00000198, 32'h00000400,
  1'd1,  5'd12, 27'h0000035e, 5'd20, 27'h00000346, 5'd11, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000cf, 5'd21, 27'h00000153, 5'd21, 27'h00000048, 32'h00000400,
  1'd1,  5'd23, 27'h00000164, 5'd0, 27'h0000032f, 5'd3, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000015b, 5'd3, 27'h0000037c, 5'd12, 27'h00000017, 32'h00000400,
  1'd1,  5'd24, 27'h00000382, 5'd1, 27'h00000189, 5'd22, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000010e, 5'd11, 27'h000002dd, 5'd0, 27'h00000210, 32'h00000400,
  1'd1,  5'd25, 27'h000002a8, 5'd14, 27'h0000036d, 5'd14, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001b, 5'd12, 27'h0000030c, 5'd21, 27'h00000003, 32'h00000400,
  1'd1,  5'd25, 27'h000002e4, 5'd24, 27'h00000145, 5'd4, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a5, 5'd24, 27'h00000062, 5'd13, 27'h0000001f, 32'h00000400,
  1'd1,  5'd24, 27'h00000267, 5'd24, 27'h000000d1, 5'd24, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000236, 5'd0, 27'h00000358, 5'd8, 27'h000001c3, 32'h00000400,
  1'd1,  5'd0, 27'h000000f1, 5'd4, 27'h0000005e, 5'd16, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001e2, 5'd1, 27'h000000e0, 5'd27, 27'h00000100, 32'h00000400,
  1'd1,  5'd1, 27'h00000076, 5'd13, 27'h000000e5, 5'd9, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000126, 5'd15, 27'h00000147, 5'd19, 27'h000001df, 32'h00000400,
  1'd1,  5'd3, 27'h00000178, 5'd14, 27'h00000247, 5'd27, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000170, 5'd24, 27'h00000191, 5'd7, 27'h000001dd, 32'h00000400,
  1'd1,  5'd2, 27'h0000000c, 5'd22, 27'h00000280, 5'd17, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000021f, 5'd24, 27'h0000028b, 5'd25, 27'h0000037a, 32'h00000400,
  1'd1,  5'd15, 27'h00000195, 5'd2, 27'h0000018c, 5'd10, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000033d, 5'd0, 27'h00000302, 5'd17, 27'h00000105, 32'h00000400,
  1'd1,  5'd13, 27'h0000024e, 5'd1, 27'h00000146, 5'd28, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000d4, 5'd12, 27'h00000100, 5'd7, 27'h000002a0, 32'h00000400,
  1'd1,  5'd12, 27'h00000381, 5'd14, 27'h00000343, 5'd20, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ac, 5'd14, 27'h000000c7, 5'd28, 27'h000000e9, 32'h00000400,
  1'd1,  5'd12, 27'h00000017, 5'd21, 27'h000002eb, 5'd6, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000225, 5'd24, 27'h0000011b, 5'd15, 27'h00000330, 32'h00000400,
  1'd1,  5'd11, 27'h00000194, 5'd22, 27'h00000123, 5'd28, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000130, 5'd2, 27'h000003ba, 5'd7, 27'h0000004a, 32'h00000400,
  1'd1,  5'd22, 27'h00000048, 5'd0, 27'h00000143, 5'd16, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000115, 5'd2, 27'h00000210, 5'd27, 27'h000002d4, 32'h00000400,
  1'd1,  5'd22, 27'h00000099, 5'd12, 27'h00000399, 5'd6, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000033a, 5'd11, 27'h00000316, 5'd16, 27'h0000009e, 32'h00000400,
  1'd1,  5'd21, 27'h000000de, 5'd14, 27'h000002f7, 5'd26, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a8, 5'd22, 27'h000002c2, 5'd6, 27'h0000020e, 32'h00000400,
  1'd1,  5'd23, 27'h000001fb, 5'd22, 27'h0000011b, 5'd18, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a1, 5'd25, 27'h00000286, 5'd30, 27'h00000223, 32'h00000400,
  1'd1,  5'd1, 27'h00000299, 5'd7, 27'h00000239, 5'd1, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000026, 5'd9, 27'h0000011f, 5'd11, 27'h0000021d, 32'h00000400,
  1'd1,  5'd0, 27'h00000350, 5'd7, 27'h00000138, 5'd23, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000004, 5'd19, 27'h000000b8, 5'd1, 27'h000000e5, 32'h00000400,
  1'd1,  5'd4, 27'h000000a2, 5'd18, 27'h0000021c, 5'd10, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000ea, 5'd18, 27'h0000036a, 5'd25, 27'h00000167, 32'h00000400,
  1'd1,  5'd4, 27'h000002d8, 5'd29, 27'h0000016a, 5'd4, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000373, 5'd27, 27'h000002cd, 5'd12, 27'h00000328, 32'h00000400,
  1'd1,  5'd3, 27'h00000023, 5'd27, 27'h00000328, 5'd25, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ef, 5'd8, 27'h00000338, 5'd4, 27'h00000270, 32'h00000400,
  1'd1,  5'd12, 27'h00000057, 5'd5, 27'h000001b4, 5'd10, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003a5, 5'd8, 27'h000002d0, 5'd24, 27'h000003bd, 32'h00000400,
  1'd1,  5'd15, 27'h0000003b, 5'd15, 27'h00000229, 5'd2, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ec, 5'd15, 27'h000002ee, 5'd13, 27'h0000007e, 32'h00000400,
  1'd1,  5'd11, 27'h000002fe, 5'd16, 27'h0000003c, 5'd24, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001de, 5'd30, 27'h000000b8, 5'd1, 27'h000000ae, 32'h00000400,
  1'd1,  5'd13, 27'h000000d3, 5'd29, 27'h0000025e, 5'd14, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038a, 5'd27, 27'h00000389, 5'd24, 27'h00000326, 32'h00000400,
  1'd1,  5'd25, 27'h000002ee, 5'd5, 27'h0000039c, 5'd4, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c8, 5'd8, 27'h000001f4, 5'd11, 27'h00000335, 32'h00000400,
  1'd1,  5'd24, 27'h00000132, 5'd5, 27'h00000371, 5'd23, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a6, 5'd16, 27'h000001bf, 5'd1, 27'h00000345, 32'h00000400,
  1'd1,  5'd22, 27'h00000095, 5'd17, 27'h0000039d, 5'd11, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000032a, 5'd16, 27'h000003dd, 5'd25, 27'h000000e5, 32'h00000400,
  1'd1,  5'd25, 27'h00000240, 5'd27, 27'h00000078, 5'd4, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000230, 5'd28, 27'h00000216, 5'd11, 27'h00000086, 32'h00000400,
  1'd1,  5'd25, 27'h00000182, 5'd28, 27'h00000291, 5'd25, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000024c, 5'd6, 27'h00000305, 5'd8, 27'h00000002, 32'h00000400,
  1'd1,  5'd4, 27'h000003de, 5'd5, 27'h00000321, 5'd18, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f4, 5'd8, 27'h000003bc, 5'd30, 27'h000000bf, 32'h00000400,
  1'd1,  5'd1, 27'h000002cd, 5'd17, 27'h0000011c, 5'd7, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023d, 5'd15, 27'h00000244, 5'd20, 27'h00000194, 32'h00000400,
  1'd1,  5'd3, 27'h0000008b, 5'd17, 27'h0000012e, 5'd27, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000033e, 5'd29, 27'h00000175, 5'd8, 27'h00000049, 32'h00000400,
  1'd1,  5'd4, 27'h000003a4, 5'd27, 27'h0000001e, 5'd20, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e9, 5'd28, 27'h00000271, 5'd27, 27'h00000399, 32'h00000400,
  1'd1,  5'd12, 27'h00000226, 5'd10, 27'h00000122, 5'd7, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000336, 5'd9, 27'h00000333, 5'd18, 27'h000003e5, 32'h00000400,
  1'd1,  5'd14, 27'h000002f4, 5'd5, 27'h000001c1, 5'd26, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b0, 5'd18, 27'h00000119, 5'd9, 27'h00000311, 32'h00000400,
  1'd1,  5'd13, 27'h0000029d, 5'd19, 27'h0000016c, 5'd19, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000074, 5'd17, 27'h00000123, 5'd28, 27'h0000007a, 32'h00000400,
  1'd1,  5'd10, 27'h000002a0, 5'd27, 27'h00000101, 5'd9, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003a5, 5'd28, 27'h000003f8, 5'd19, 27'h00000258, 32'h00000400,
  1'd1,  5'd10, 27'h000002d6, 5'd29, 27'h0000024c, 5'd28, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000010e, 5'd5, 27'h00000105, 5'd7, 27'h0000034d, 32'h00000400,
  1'd1,  5'd24, 27'h000003ab, 5'd8, 27'h00000208, 5'd18, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000373, 5'd5, 27'h0000039d, 5'd26, 27'h00000008, 32'h00000400,
  1'd1,  5'd25, 27'h000000b0, 5'd17, 27'h00000002, 5'd5, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000248, 5'd19, 27'h00000339, 5'd17, 27'h000002f1, 32'h00000400,
  1'd1,  5'd24, 27'h00000377, 5'd16, 27'h00000162, 5'd27, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000356, 5'd29, 27'h000002de, 5'd5, 27'h000001e5, 32'h00000400,
  1'd1,  5'd21, 27'h0000008b, 5'd29, 27'h00000308, 5'd19, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000339, 5'd28, 27'h00000273, 5'd28, 27'h0000001d, 32'h00000400,
  1'd1,  5'd6, 27'h00000082, 5'd1, 27'h000002b6, 5'd8, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002c7, 5'd5, 27'h00000035, 5'd19, 27'h000001d1, 32'h00000400,
  1'd1,  5'd5, 27'h0000012d, 5'd3, 27'h000003db, 5'd29, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000221, 5'd14, 27'h0000034c, 5'd0, 27'h0000024e, 32'h00000400,
  1'd1,  5'd6, 27'h00000173, 5'd11, 27'h0000015a, 5'd12, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000245, 5'd15, 27'h000001c1, 5'd24, 27'h000003d3, 32'h00000400,
  1'd1,  5'd5, 27'h0000017f, 5'd21, 27'h0000015d, 5'd4, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000162, 5'd23, 27'h00000140, 5'd11, 27'h0000011a, 32'h00000400,
  1'd1,  5'd9, 27'h00000378, 5'd21, 27'h000003f4, 5'd21, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000079, 5'd3, 27'h000003bc, 5'd8, 27'h00000088, 32'h00000400,
  1'd1,  5'd19, 27'h0000037a, 5'd3, 27'h00000037, 5'd18, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000b2, 5'd4, 27'h000001f7, 5'd29, 27'h00000010, 32'h00000400,
  1'd1,  5'd17, 27'h00000240, 5'd10, 27'h00000224, 5'd3, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000028b, 5'd14, 27'h00000065, 5'd12, 27'h00000389, 32'h00000400,
  1'd1,  5'd18, 27'h000003eb, 5'd13, 27'h0000033c, 5'd23, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000335, 5'd23, 27'h000003dc, 5'd1, 27'h00000069, 32'h00000400,
  1'd1,  5'd17, 27'h000000df, 5'd24, 27'h00000293, 5'd11, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000148, 5'd21, 27'h0000000e, 5'd22, 27'h000003b3, 32'h00000400,
  1'd1,  5'd30, 27'h00000050, 5'd3, 27'h000001a0, 5'd1, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000197, 5'd5, 27'h0000008c, 5'd13, 27'h00000270, 32'h00000400,
  1'd1,  5'd30, 27'h000003bf, 5'd4, 27'h000003cb, 5'd23, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000011b, 5'd14, 27'h000003d6, 5'd0, 27'h00000083, 32'h00000400,
  1'd1,  5'd27, 27'h0000002b, 5'd12, 27'h00000058, 5'd11, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000023b, 5'd13, 27'h00000357, 5'd21, 27'h000001ff, 32'h00000400,
  1'd1,  5'd28, 27'h000001e2, 5'd21, 27'h00000191, 5'd2, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000158, 5'd24, 27'h0000001b, 5'd11, 27'h000002bf, 32'h00000400,
  1'd1,  5'd30, 27'h0000004f, 5'd24, 27'h000003c3, 5'd23, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003f0, 5'd0, 27'h00000304, 5'd3, 27'h000003cb, 32'h00000400,
  1'd1,  5'd8, 27'h000003eb, 5'd1, 27'h000001c4, 5'd11, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ce, 5'd0, 27'h000002eb, 5'd21, 27'h00000008, 32'h00000400,
  1'd1,  5'd7, 27'h000003ec, 5'd13, 27'h00000187, 5'd8, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ec, 5'd11, 27'h000001ba, 5'd15, 27'h000002d7, 32'h00000400,
  1'd1,  5'd9, 27'h00000377, 5'd15, 27'h00000107, 5'd30, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e9, 5'd23, 27'h0000035e, 5'd7, 27'h000001bc, 32'h00000400,
  1'd1,  5'd7, 27'h000002df, 5'd24, 27'h000001a4, 5'd19, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000365, 5'd25, 27'h000002e2, 5'd27, 27'h00000323, 32'h00000400,
  1'd1,  5'd16, 27'h00000318, 5'd4, 27'h000001c4, 5'd0, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000088, 5'd1, 27'h000003d0, 5'd10, 27'h000002a3, 32'h00000400,
  1'd1,  5'd16, 27'h000001bc, 5'd3, 27'h000002d3, 5'd22, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000009b, 5'd13, 27'h0000020b, 5'd5, 27'h00000225, 32'h00000400,
  1'd1,  5'd18, 27'h00000097, 5'd10, 27'h000001d5, 5'd17, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009a, 5'd11, 27'h000000a8, 5'd29, 27'h00000080, 32'h00000400,
  1'd1,  5'd16, 27'h000001bf, 5'd22, 27'h0000037d, 5'd5, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000a6, 5'd21, 27'h0000018c, 5'd17, 27'h000001e6, 32'h00000400,
  1'd1,  5'd19, 27'h00000201, 5'd21, 27'h000000c6, 5'd26, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000183, 5'd1, 27'h00000134, 5'd9, 27'h000000ba, 32'h00000400,
  1'd1,  5'd28, 27'h0000018a, 5'd2, 27'h000000d8, 5'd20, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000018d, 5'd4, 27'h0000010d, 5'd29, 27'h00000021, 32'h00000400,
  1'd1,  5'd27, 27'h000000f1, 5'd14, 27'h000001a1, 5'd6, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000178, 5'd13, 27'h0000002e, 5'd16, 27'h000001e6, 32'h00000400,
  1'd1,  5'd29, 27'h0000037b, 5'd12, 27'h00000106, 5'd27, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003d1, 5'd21, 27'h000003c7, 5'd6, 27'h0000020a, 32'h00000400,
  1'd1,  5'd27, 27'h000001db, 5'd22, 27'h00000040, 5'd18, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000313, 5'd23, 27'h00000303, 5'd30, 27'h0000038c, 32'h00000400,
  1'd1,  5'd8, 27'h00000192, 5'd10, 27'h0000014e, 5'd3, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ef, 5'd6, 27'h00000284, 5'd14, 27'h000000fd, 32'h00000400,
  1'd1,  5'd6, 27'h00000164, 5'd7, 27'h0000000e, 5'd22, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000021f, 5'd20, 27'h00000034, 5'd3, 27'h0000023d, 32'h00000400,
  1'd1,  5'd8, 27'h0000013c, 5'd20, 27'h000000bb, 5'd13, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002bd, 5'd17, 27'h000001e6, 5'd22, 27'h00000172, 32'h00000400,
  1'd1,  5'd8, 27'h000000c6, 5'd25, 27'h00000377, 5'd3, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000141, 5'd29, 27'h00000189, 5'd15, 27'h00000046, 32'h00000400,
  1'd1,  5'd6, 27'h00000274, 5'd30, 27'h000002ec, 5'd21, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000064, 5'd6, 27'h00000049, 5'd1, 27'h0000037b, 32'h00000400,
  1'd1,  5'd17, 27'h00000256, 5'd7, 27'h0000002e, 5'd13, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000007f, 5'd9, 27'h0000039f, 5'd23, 27'h00000374, 32'h00000400,
  1'd1,  5'd15, 27'h00000234, 5'd20, 27'h00000026, 5'd0, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d1, 5'd15, 27'h00000257, 5'd14, 27'h000003e0, 32'h00000400,
  1'd1,  5'd17, 27'h0000017e, 5'd18, 27'h000002b9, 5'd21, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000249, 5'd28, 27'h000000a3, 5'd4, 27'h00000223, 32'h00000400,
  1'd1,  5'd16, 27'h0000034f, 5'd29, 27'h0000034f, 5'd15, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000001f, 5'd27, 27'h00000345, 5'd21, 27'h00000338, 32'h00000400,
  1'd1,  5'd26, 27'h00000128, 5'd6, 27'h0000009c, 5'd2, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000269, 5'd9, 27'h000001f7, 5'd14, 27'h0000000f, 32'h00000400,
  1'd1,  5'd30, 27'h000000ca, 5'd6, 27'h0000016f, 5'd24, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000339, 5'd19, 27'h0000019f, 5'd3, 27'h000001f8, 32'h00000400,
  1'd1,  5'd28, 27'h0000033a, 5'd18, 27'h0000004d, 5'd11, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000021d, 5'd18, 27'h00000107, 5'd25, 27'h000001b4, 32'h00000400,
  1'd1,  5'd28, 27'h00000185, 5'd26, 27'h000002e0, 5'd4, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000379, 5'd30, 27'h000003a0, 5'd13, 27'h000003f7, 32'h00000400,
  1'd1,  5'd29, 27'h00000116, 5'd29, 27'h0000026f, 5'd21, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001b9, 5'd8, 27'h000001cb, 5'd6, 27'h00000146, 32'h00000400,
  1'd1,  5'd5, 27'h000000f5, 5'd8, 27'h000000c8, 5'd16, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000002e, 5'd9, 27'h0000030f, 5'd30, 27'h0000025e, 32'h00000400,
  1'd1,  5'd7, 27'h0000023b, 5'd15, 27'h0000037b, 5'd5, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000063, 5'd17, 27'h000003c0, 5'd19, 27'h0000005e, 32'h00000400,
  1'd1,  5'd9, 27'h0000025d, 5'd15, 27'h00000216, 5'd26, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ac, 5'd27, 27'h000002cb, 5'd6, 27'h0000026d, 32'h00000400,
  1'd1,  5'd5, 27'h0000013c, 5'd30, 27'h000003ce, 5'd19, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000001c, 5'd27, 27'h000003b8, 5'd28, 27'h00000225, 32'h00000400,
  1'd1,  5'd16, 27'h00000330, 5'd10, 27'h000000d3, 5'd6, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000276, 5'd5, 27'h00000273, 5'd17, 27'h00000248, 32'h00000400,
  1'd1,  5'd15, 27'h00000210, 5'd8, 27'h000000b7, 5'd26, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ba, 5'd17, 27'h00000304, 5'd8, 27'h00000309, 32'h00000400,
  1'd1,  5'd16, 27'h000000ff, 5'd20, 27'h0000004c, 5'd20, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000044, 5'd16, 27'h000002cb, 5'd30, 27'h00000392, 32'h00000400,
  1'd1,  5'd18, 27'h000002b5, 5'd26, 27'h00000288, 5'd9, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a5, 5'd26, 27'h00000188, 5'd15, 27'h000002a7, 32'h00000400,
  1'd1,  5'd17, 27'h00000082, 5'd27, 27'h000001b4, 5'd26, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002da, 5'd5, 27'h0000031e, 5'd10, 27'h000000b7, 32'h00000400,
  1'd1,  5'd28, 27'h00000237, 5'd6, 27'h000001d7, 5'd16, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000004b, 5'd9, 27'h000001f4, 5'd28, 27'h0000037d, 32'h00000400,
  1'd1,  5'd26, 27'h0000003f, 5'd20, 27'h00000113, 5'd10, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000079, 5'd15, 27'h000003c3, 5'd20, 27'h000001a1, 32'h00000400,
  1'd1,  5'd28, 27'h0000036e, 5'd18, 27'h000003ec, 5'd26, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000297, 5'd27, 27'h000001f3, 5'd10, 27'h0000007c, 32'h00000400,
  1'd1,  5'd25, 27'h000003c6, 5'd29, 27'h0000001d, 5'd20, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001cf, 5'd29, 27'h000000ff, 5'd29, 27'h00000267, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000028, 5'd4, 27'h00000158, 5'd1, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000044, 5'd1, 27'h00000370, 5'd13, 27'h000000a9, 32'h00000400,
  1'd1,  5'd3, 27'h00000200, 5'd1, 27'h000003be, 5'd23, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000056, 5'd12, 27'h00000145, 5'd3, 27'h0000018a, 32'h00000400,
  1'd1,  5'd0, 27'h00000335, 5'd13, 27'h00000245, 5'd12, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001a2, 5'd10, 27'h00000165, 5'd23, 27'h000002d0, 32'h00000400,
  1'd1,  5'd3, 27'h000000a0, 5'd22, 27'h00000025, 5'd2, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000fc, 5'd22, 27'h00000005, 5'd11, 27'h00000063, 32'h00000400,
  1'd1,  5'd4, 27'h00000378, 5'd21, 27'h0000010d, 5'd23, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f2, 5'd2, 27'h00000245, 5'd1, 27'h00000247, 32'h00000400,
  1'd1,  5'd13, 27'h000000b5, 5'd3, 27'h000001ed, 5'd12, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002fe, 5'd4, 27'h000003cf, 5'd22, 27'h00000291, 32'h00000400,
  1'd1,  5'd11, 27'h00000009, 5'd13, 27'h00000282, 5'd3, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000280, 5'd15, 27'h000001f5, 5'd10, 27'h00000241, 32'h00000400,
  1'd1,  5'd12, 27'h0000035d, 5'd13, 27'h000003b5, 5'd21, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c7, 5'd21, 27'h000002be, 5'd4, 27'h00000128, 32'h00000400,
  1'd1,  5'd11, 27'h000001fa, 5'd24, 27'h00000201, 5'd14, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000029d, 5'd22, 27'h00000114, 5'd25, 27'h0000022f, 32'h00000400,
  1'd1,  5'd23, 27'h00000025, 5'd0, 27'h00000313, 5'd3, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003f8, 5'd4, 27'h000000d5, 5'd15, 27'h00000033, 32'h00000400,
  1'd1,  5'd23, 27'h00000392, 5'd3, 27'h00000345, 5'd20, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000368, 5'd12, 27'h000001e1, 5'd2, 27'h00000082, 32'h00000400,
  1'd1,  5'd23, 27'h00000121, 5'd14, 27'h0000039b, 5'd13, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000199, 5'd10, 27'h0000032f, 5'd24, 27'h00000136, 32'h00000400,
  1'd1,  5'd25, 27'h0000011a, 5'd25, 27'h00000326, 5'd4, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000320, 5'd24, 27'h000000d9, 5'd10, 27'h000001ce, 32'h00000400,
  1'd1,  5'd21, 27'h00000314, 5'd22, 27'h000003cc, 5'd24, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000ac, 5'd3, 27'h0000010b, 5'd8, 27'h000003b7, 32'h00000400,
  1'd1,  5'd4, 27'h00000374, 5'd3, 27'h00000083, 5'd20, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002bf, 5'd3, 27'h00000309, 5'd27, 27'h00000251, 32'h00000400,
  1'd1,  5'd3, 27'h000002ec, 5'd11, 27'h0000011e, 5'd9, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000005d, 5'd13, 27'h000003d1, 5'd20, 27'h0000027e, 32'h00000400,
  1'd1,  5'd0, 27'h000000e1, 5'd13, 27'h000002f9, 5'd28, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000cd, 5'd22, 27'h0000012d, 5'd10, 27'h000000ce, 32'h00000400,
  1'd1,  5'd4, 27'h000001d3, 5'd20, 27'h000002c9, 5'd20, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000016c, 5'd25, 27'h0000007d, 5'd30, 27'h0000016e, 32'h00000400,
  1'd1,  5'd15, 27'h00000070, 5'd4, 27'h0000014e, 5'd7, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000151, 5'd0, 27'h000002d7, 5'd19, 27'h00000128, 32'h00000400,
  1'd1,  5'd10, 27'h00000176, 5'd4, 27'h000000d7, 5'd29, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000008c, 5'd12, 27'h0000025f, 5'd9, 27'h000000a7, 32'h00000400,
  1'd1,  5'd14, 27'h00000154, 5'd10, 27'h000001a2, 5'd17, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000357, 5'd10, 27'h000001eb, 5'd30, 27'h00000092, 32'h00000400,
  1'd1,  5'd10, 27'h00000370, 5'd25, 27'h000002e1, 5'd5, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000001d, 5'd24, 27'h0000004c, 5'd17, 27'h0000021c, 32'h00000400,
  1'd1,  5'd14, 27'h00000060, 5'd24, 27'h000003d9, 5'd28, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000198, 5'd2, 27'h000001ba, 5'd8, 27'h000003dc, 32'h00000400,
  1'd1,  5'd21, 27'h000000ab, 5'd3, 27'h000001ca, 5'd18, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000018c, 5'd0, 27'h00000166, 5'd27, 27'h00000217, 32'h00000400,
  1'd1,  5'd22, 27'h00000136, 5'd11, 27'h00000003, 5'd7, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000038d, 5'd12, 27'h00000007, 5'd17, 27'h00000281, 32'h00000400,
  1'd1,  5'd21, 27'h000003ef, 5'd10, 27'h000002d6, 5'd30, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000332, 5'd24, 27'h000000cb, 5'd7, 27'h0000012b, 32'h00000400,
  1'd1,  5'd23, 27'h000001db, 5'd25, 27'h000002e2, 5'd19, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001af, 5'd24, 27'h000003cb, 5'd27, 27'h0000021b, 32'h00000400,
  1'd1,  5'd1, 27'h00000357, 5'd7, 27'h0000011e, 5'd0, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000020a, 5'd6, 27'h0000019e, 5'd11, 27'h000000ee, 32'h00000400,
  1'd1,  5'd5, 27'h0000006e, 5'd8, 27'h00000045, 5'd20, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036d, 5'd17, 27'h00000194, 5'd3, 27'h00000228, 32'h00000400,
  1'd1,  5'd2, 27'h000000d0, 5'd16, 27'h00000091, 5'd10, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000270, 5'd17, 27'h000003b6, 5'd24, 27'h000003a7, 32'h00000400,
  1'd1,  5'd4, 27'h00000110, 5'd27, 27'h00000207, 5'd2, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000353, 5'd28, 27'h000002ee, 5'd12, 27'h0000021f, 32'h00000400,
  1'd1,  5'd3, 27'h0000030e, 5'd26, 27'h0000026f, 5'd22, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b6, 5'd8, 27'h000001f1, 5'd2, 27'h00000249, 32'h00000400,
  1'd1,  5'd14, 27'h000001fa, 5'd5, 27'h00000216, 5'd13, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000308, 5'd8, 27'h00000133, 5'd24, 27'h00000209, 32'h00000400,
  1'd1,  5'd10, 27'h0000027c, 5'd17, 27'h00000112, 5'd3, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002be, 5'd19, 27'h000002c7, 5'd12, 27'h000002a1, 32'h00000400,
  1'd1,  5'd15, 27'h000000da, 5'd16, 27'h0000037a, 5'd22, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000007f, 5'd27, 27'h000002b8, 5'd3, 27'h00000094, 32'h00000400,
  1'd1,  5'd10, 27'h00000230, 5'd25, 27'h000003c8, 5'd13, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000cd, 5'd26, 27'h0000004f, 5'd21, 27'h00000295, 32'h00000400,
  1'd1,  5'd20, 27'h00000382, 5'd8, 27'h0000028b, 5'd4, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000202, 5'd6, 27'h000000b7, 5'd11, 27'h0000016f, 32'h00000400,
  1'd1,  5'd20, 27'h0000033e, 5'd5, 27'h000000dd, 5'd20, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032b, 5'd17, 27'h00000325, 5'd1, 27'h000000d6, 32'h00000400,
  1'd1,  5'd22, 27'h000003ca, 5'd18, 27'h00000229, 5'd12, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002cc, 5'd18, 27'h000001fe, 5'd24, 27'h000001f0, 32'h00000400,
  1'd1,  5'd24, 27'h00000267, 5'd26, 27'h00000046, 5'd2, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001a6, 5'd28, 27'h00000144, 5'd12, 27'h000002d6, 32'h00000400,
  1'd1,  5'd21, 27'h00000080, 5'd26, 27'h0000029a, 5'd24, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000017d, 5'd8, 27'h00000094, 5'd6, 27'h0000028c, 32'h00000400,
  1'd1,  5'd3, 27'h00000385, 5'd9, 27'h00000389, 5'd17, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003da, 5'd8, 27'h000002eb, 5'd26, 27'h000000bc, 32'h00000400,
  1'd1,  5'd3, 27'h0000037d, 5'd19, 27'h0000026c, 5'd6, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000059, 5'd19, 27'h0000012f, 5'd18, 27'h000000b1, 32'h00000400,
  1'd1,  5'd3, 27'h00000250, 5'd20, 27'h0000015c, 5'd30, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000035, 5'd29, 27'h00000205, 5'd6, 27'h0000001b, 32'h00000400,
  1'd1,  5'd0, 27'h00000113, 5'd28, 27'h000002ad, 5'd15, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d9, 5'd26, 27'h000000f8, 5'd30, 27'h00000086, 32'h00000400,
  1'd1,  5'd14, 27'h00000119, 5'd5, 27'h0000011b, 5'd9, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000070, 5'd7, 27'h0000003a, 5'd15, 27'h000003d4, 32'h00000400,
  1'd1,  5'd14, 27'h00000027, 5'd9, 27'h000003a7, 5'd29, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000be, 5'd17, 27'h00000138, 5'd10, 27'h00000030, 32'h00000400,
  1'd1,  5'd12, 27'h0000037e, 5'd16, 27'h00000391, 5'd15, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001e0, 5'd16, 27'h0000032f, 5'd29, 27'h000001a6, 32'h00000400,
  1'd1,  5'd13, 27'h00000384, 5'd27, 27'h000003f9, 5'd8, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000175, 5'd29, 27'h00000379, 5'd18, 27'h000000e2, 32'h00000400,
  1'd1,  5'd12, 27'h00000394, 5'd30, 27'h000000c6, 5'd30, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000081, 5'd10, 27'h00000052, 5'd7, 27'h0000037d, 32'h00000400,
  1'd1,  5'd22, 27'h00000287, 5'd8, 27'h000002d5, 5'd16, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006c, 5'd9, 27'h000001fe, 5'd26, 27'h00000180, 32'h00000400,
  1'd1,  5'd22, 27'h00000116, 5'd19, 27'h0000023b, 5'd9, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e7, 5'd19, 27'h000003f3, 5'd18, 27'h0000023e, 32'h00000400,
  1'd1,  5'd23, 27'h00000246, 5'd20, 27'h00000036, 5'd30, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000110, 5'd25, 27'h0000039e, 5'd7, 27'h00000050, 32'h00000400,
  1'd1,  5'd22, 27'h00000080, 5'd29, 27'h000003e2, 5'd18, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000340, 5'd30, 27'h000001df, 5'd26, 27'h000000ae, 32'h00000400,
  1'd1,  5'd8, 27'h000000a7, 5'd0, 27'h00000233, 5'd9, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b1, 5'd4, 27'h00000121, 5'd16, 27'h0000002d, 32'h00000400,
  1'd1,  5'd9, 27'h00000133, 5'd1, 27'h00000216, 5'd28, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e8, 5'd13, 27'h000003d4, 5'd4, 27'h00000235, 32'h00000400,
  1'd1,  5'd8, 27'h00000365, 5'd10, 27'h0000020d, 5'd14, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000228, 5'd11, 27'h000000e8, 5'd25, 27'h00000063, 32'h00000400,
  1'd1,  5'd5, 27'h00000381, 5'd22, 27'h000001dd, 5'd4, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001db, 5'd24, 27'h0000030f, 5'd14, 27'h000001a7, 32'h00000400,
  1'd1,  5'd10, 27'h000000f5, 5'd21, 27'h000000b3, 5'd25, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000f1, 5'd2, 27'h000001f5, 5'd5, 27'h0000010c, 32'h00000400,
  1'd1,  5'd17, 27'h00000229, 5'd0, 27'h0000035f, 5'd17, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000007d, 5'd0, 27'h0000009c, 5'd29, 27'h000000d9, 32'h00000400,
  1'd1,  5'd15, 27'h0000037d, 5'd14, 27'h0000012c, 5'd2, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000286, 5'd12, 27'h000002c0, 5'd11, 27'h000002d5, 32'h00000400,
  1'd1,  5'd17, 27'h000000d1, 5'd12, 27'h00000028, 5'd23, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000011c, 5'd22, 27'h0000025e, 5'd0, 27'h000001f0, 32'h00000400,
  1'd1,  5'd19, 27'h0000025c, 5'd25, 27'h0000019a, 5'd14, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c6, 5'd24, 27'h0000005c, 5'd22, 27'h000003e2, 32'h00000400,
  1'd1,  5'd27, 27'h0000016d, 5'd1, 27'h00000017, 5'd4, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000013f, 5'd2, 27'h0000007e, 5'd11, 27'h000002f7, 32'h00000400,
  1'd1,  5'd26, 27'h00000206, 5'd3, 27'h000003fe, 5'd21, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002ee, 5'd12, 27'h0000021d, 5'd4, 27'h0000024e, 32'h00000400,
  1'd1,  5'd27, 27'h00000382, 5'd14, 27'h00000174, 5'd12, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000317, 5'd10, 27'h000001ec, 5'd22, 27'h00000240, 32'h00000400,
  1'd1,  5'd29, 27'h000002e4, 5'd21, 27'h000002f4, 5'd3, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012b, 5'd23, 27'h00000218, 5'd11, 27'h00000344, 32'h00000400,
  1'd1,  5'd29, 27'h00000090, 5'd22, 27'h0000034f, 5'd22, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000a4, 5'd2, 27'h0000003f, 5'd2, 27'h000002e3, 32'h00000400,
  1'd1,  5'd5, 27'h00000312, 5'd3, 27'h000003d9, 5'd14, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000011, 5'd2, 27'h0000022c, 5'd24, 27'h000001cf, 32'h00000400,
  1'd1,  5'd6, 27'h000002bb, 5'd11, 27'h00000278, 5'd10, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c2, 5'd10, 27'h000001a9, 5'd15, 27'h00000395, 32'h00000400,
  1'd1,  5'd6, 27'h000003b7, 5'd14, 27'h0000038b, 5'd30, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000312, 5'd25, 27'h00000308, 5'd10, 27'h0000011a, 32'h00000400,
  1'd1,  5'd7, 27'h00000006, 5'd21, 27'h00000378, 5'd15, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ea, 5'd23, 27'h0000007e, 5'd26, 27'h00000377, 32'h00000400,
  1'd1,  5'd19, 27'h000001b1, 5'd2, 27'h0000013e, 5'd2, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000339, 5'd4, 27'h000000f5, 5'd11, 27'h0000000a, 32'h00000400,
  1'd1,  5'd18, 27'h000000fb, 5'd1, 27'h00000180, 5'd25, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d3, 5'd15, 27'h00000084, 5'd10, 27'h00000023, 32'h00000400,
  1'd1,  5'd17, 27'h0000010f, 5'd15, 27'h00000078, 5'd16, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000cc, 5'd14, 27'h00000279, 5'd27, 27'h000000e7, 32'h00000400,
  1'd1,  5'd15, 27'h00000207, 5'd24, 27'h0000013e, 5'd9, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000235, 5'd24, 27'h00000367, 5'd18, 27'h0000005a, 32'h00000400,
  1'd1,  5'd20, 27'h0000027f, 5'd22, 27'h000001b5, 5'd27, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002f4, 5'd0, 27'h0000011f, 5'd10, 27'h000000fe, 32'h00000400,
  1'd1,  5'd26, 27'h00000242, 5'd0, 27'h000000d2, 5'd17, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000391, 5'd2, 27'h0000039e, 5'd26, 27'h000002ff, 32'h00000400,
  1'd1,  5'd27, 27'h0000011d, 5'd12, 27'h000002c4, 5'd5, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002eb, 5'd14, 27'h0000000d, 5'd15, 27'h00000265, 32'h00000400,
  1'd1,  5'd27, 27'h0000027e, 5'd14, 27'h00000168, 5'd30, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000f1, 5'd24, 27'h000003f2, 5'd7, 27'h00000022, 32'h00000400,
  1'd1,  5'd27, 27'h00000286, 5'd23, 27'h0000025f, 5'd17, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000c0, 5'd23, 27'h000002b0, 5'd30, 27'h000002e2, 32'h00000400,
  1'd1,  5'd6, 27'h00000165, 5'd5, 27'h000001fd, 5'd2, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000011d, 5'd6, 27'h0000028a, 5'd13, 27'h0000013a, 32'h00000400,
  1'd1,  5'd8, 27'h000003d8, 5'd7, 27'h000000b1, 5'd22, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031e, 5'd17, 27'h00000287, 5'd3, 27'h0000013e, 32'h00000400,
  1'd1,  5'd9, 27'h000001c7, 5'd18, 27'h000003dd, 5'd11, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020f, 5'd19, 27'h00000038, 5'd23, 27'h000001ae, 32'h00000400,
  1'd1,  5'd7, 27'h0000021c, 5'd29, 27'h00000391, 5'd0, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000123, 5'd29, 27'h00000245, 5'd11, 27'h00000391, 32'h00000400,
  1'd1,  5'd7, 27'h0000036f, 5'd27, 27'h00000237, 5'd24, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000178, 5'd8, 27'h00000312, 5'd4, 27'h000000a8, 32'h00000400,
  1'd1,  5'd18, 27'h00000117, 5'd8, 27'h000001dd, 5'd13, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000119, 5'd7, 27'h0000001b, 5'd21, 27'h00000117, 32'h00000400,
  1'd1,  5'd19, 27'h00000057, 5'd18, 27'h000002ab, 5'd4, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003d8, 5'd18, 27'h00000237, 5'd12, 27'h000003e5, 32'h00000400,
  1'd1,  5'd16, 27'h00000122, 5'd20, 27'h0000006e, 5'd23, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000301, 5'd27, 27'h000003d6, 5'd2, 27'h00000367, 32'h00000400,
  1'd1,  5'd18, 27'h00000317, 5'd28, 27'h000001da, 5'd12, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000014b, 5'd27, 27'h0000002a, 5'd22, 27'h00000386, 32'h00000400,
  1'd1,  5'd30, 27'h000000bb, 5'd9, 27'h0000007d, 5'd0, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e8, 5'd6, 27'h000003dc, 5'd10, 27'h00000313, 32'h00000400,
  1'd1,  5'd27, 27'h00000181, 5'd10, 27'h00000124, 5'd21, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000322, 5'd18, 27'h000001eb, 5'd1, 27'h00000021, 32'h00000400,
  1'd1,  5'd30, 27'h0000002f, 5'd18, 27'h0000016b, 5'd11, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000018c, 5'd19, 27'h000001a1, 5'd24, 27'h0000020f, 32'h00000400,
  1'd1,  5'd30, 27'h000003dc, 5'd27, 27'h000003ed, 5'd0, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000240, 5'd28, 27'h000002b0, 5'd12, 27'h000001e7, 32'h00000400,
  1'd1,  5'd29, 27'h000001b3, 5'd30, 27'h00000006, 5'd24, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d4, 5'd8, 27'h00000219, 5'd10, 27'h0000008f, 32'h00000400,
  1'd1,  5'd9, 27'h00000351, 5'd7, 27'h00000136, 5'd18, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000155, 5'd6, 27'h00000349, 5'd30, 27'h00000007, 32'h00000400,
  1'd1,  5'd5, 27'h000002d0, 5'd18, 27'h00000219, 5'd8, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000199, 5'd19, 27'h00000399, 5'd17, 27'h00000029, 32'h00000400,
  1'd1,  5'd8, 27'h00000109, 5'd20, 27'h0000026f, 5'd27, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000271, 5'd28, 27'h00000243, 5'd5, 27'h00000399, 32'h00000400,
  1'd1,  5'd7, 27'h00000272, 5'd26, 27'h00000138, 5'd17, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000022a, 5'd28, 27'h000000c8, 5'd30, 27'h000000cb, 32'h00000400,
  1'd1,  5'd15, 27'h00000301, 5'd7, 27'h000003b1, 5'd6, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e6, 5'd6, 27'h000001d3, 5'd15, 27'h00000309, 32'h00000400,
  1'd1,  5'd20, 27'h000001a2, 5'd9, 27'h000003ad, 5'd29, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000010b, 5'd20, 27'h00000290, 5'd8, 27'h00000212, 32'h00000400,
  1'd1,  5'd15, 27'h00000399, 5'd17, 27'h00000195, 5'd19, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000341, 5'd17, 27'h00000283, 5'd26, 27'h00000287, 32'h00000400,
  1'd1,  5'd17, 27'h000003aa, 5'd29, 27'h00000329, 5'd7, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025c, 5'd30, 27'h0000032c, 5'd17, 27'h0000012b, 32'h00000400,
  1'd1,  5'd15, 27'h0000024f, 5'd28, 27'h00000167, 5'd26, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a6, 5'd8, 27'h000002f1, 5'd8, 27'h000000fb, 32'h00000400,
  1'd1,  5'd30, 27'h00000336, 5'd6, 27'h00000354, 5'd17, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000046, 5'd10, 27'h000000f2, 5'd27, 27'h00000271, 32'h00000400,
  1'd1,  5'd30, 27'h00000221, 5'd18, 27'h00000075, 5'd8, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000028, 5'd20, 27'h00000049, 5'd20, 27'h0000018b, 32'h00000400,
  1'd1,  5'd28, 27'h00000176, 5'd18, 27'h000002be, 5'd30, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e1, 5'd29, 27'h0000038f, 5'd8, 27'h000002f9, 32'h00000400,
  1'd1,  5'd27, 27'h000000ac, 5'd29, 27'h0000033c, 5'd19, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000103, 5'd30, 27'h00000308, 5'd27, 27'h00000310, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000188, 5'd1, 27'h00000212, 5'd1, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000245, 5'd2, 27'h00000236, 5'd13, 27'h00000238, 32'h00000400,
  1'd1,  5'd2, 27'h000002ff, 5'd4, 27'h00000222, 5'd23, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d3, 5'd13, 27'h000001e0, 5'd3, 27'h00000241, 32'h00000400,
  1'd1,  5'd1, 27'h00000109, 5'd11, 27'h000001fd, 5'd13, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ce, 5'd14, 27'h0000008f, 5'd22, 27'h0000030f, 32'h00000400,
  1'd1,  5'd0, 27'h00000351, 5'd25, 27'h0000013b, 5'd1, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000282, 5'd22, 27'h0000006d, 5'd11, 27'h00000244, 32'h00000400,
  1'd1,  5'd3, 27'h0000033d, 5'd20, 27'h000002d7, 5'd22, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000c8, 5'd3, 27'h0000025f, 5'd2, 27'h0000002a, 32'h00000400,
  1'd1,  5'd10, 27'h000002fa, 5'd2, 27'h00000186, 5'd10, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002ae, 5'd1, 27'h0000000b, 5'd23, 27'h000000e0, 32'h00000400,
  1'd1,  5'd10, 27'h000003df, 5'd11, 27'h000000af, 5'd1, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000373, 5'd11, 27'h000001b0, 5'd12, 27'h0000030d, 32'h00000400,
  1'd1,  5'd10, 27'h00000253, 5'd14, 27'h000000a0, 5'd20, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000021, 5'd21, 27'h000003b2, 5'd1, 27'h000001e5, 32'h00000400,
  1'd1,  5'd12, 27'h00000066, 5'd25, 27'h000000a2, 5'd14, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000069, 5'd24, 27'h00000346, 5'd22, 27'h00000267, 32'h00000400,
  1'd1,  5'd22, 27'h000003b3, 5'd0, 27'h00000006, 5'd1, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002bb, 5'd0, 27'h00000162, 5'd12, 27'h00000328, 32'h00000400,
  1'd1,  5'd20, 27'h000002ff, 5'd1, 27'h000001a7, 5'd23, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002dc, 5'd11, 27'h00000378, 5'd1, 27'h00000058, 32'h00000400,
  1'd1,  5'd24, 27'h000001d6, 5'd10, 27'h00000242, 5'd13, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000112, 5'd12, 27'h000000c5, 5'd24, 27'h000000b0, 32'h00000400,
  1'd1,  5'd20, 27'h000003bc, 5'd25, 27'h000000a7, 5'd4, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b4, 5'd21, 27'h00000292, 5'd13, 27'h00000366, 32'h00000400,
  1'd1,  5'd21, 27'h000000c1, 5'd24, 27'h00000069, 5'd23, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000048, 5'd2, 27'h00000150, 5'd8, 27'h000001b5, 32'h00000400,
  1'd1,  5'd4, 27'h00000094, 5'd3, 27'h000001fb, 5'd19, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000258, 5'd4, 27'h00000126, 5'd28, 27'h00000050, 32'h00000400,
  1'd1,  5'd2, 27'h00000148, 5'd14, 27'h00000161, 5'd6, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000250, 5'd10, 27'h0000035b, 5'd15, 27'h00000321, 32'h00000400,
  1'd1,  5'd4, 27'h000001eb, 5'd11, 27'h00000223, 5'd28, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000329, 5'd20, 27'h00000339, 5'd9, 27'h0000005d, 32'h00000400,
  1'd1,  5'd1, 27'h000000d0, 5'd24, 27'h00000344, 5'd16, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000255, 5'd24, 27'h000002c6, 5'd30, 27'h00000298, 32'h00000400,
  1'd1,  5'd14, 27'h0000032f, 5'd4, 27'h0000004c, 5'd5, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000245, 5'd3, 27'h00000081, 5'd16, 27'h0000032c, 32'h00000400,
  1'd1,  5'd11, 27'h000001f6, 5'd2, 27'h000001bf, 5'd30, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000225, 5'd12, 27'h0000038d, 5'd7, 27'h000002c4, 32'h00000400,
  1'd1,  5'd11, 27'h000002a9, 5'd13, 27'h000001ba, 5'd19, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000306, 5'd15, 27'h0000005d, 5'd28, 27'h00000310, 32'h00000400,
  1'd1,  5'd11, 27'h00000135, 5'd23, 27'h00000318, 5'd9, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f8, 5'd22, 27'h00000085, 5'd16, 27'h0000006f, 32'h00000400,
  1'd1,  5'd10, 27'h000002cb, 5'd25, 27'h00000017, 5'd28, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e0, 5'd3, 27'h000000fb, 5'd9, 27'h000003f4, 32'h00000400,
  1'd1,  5'd21, 27'h0000019f, 5'd5, 27'h0000009b, 5'd15, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ac, 5'd2, 27'h0000037a, 5'd27, 27'h00000308, 32'h00000400,
  1'd1,  5'd22, 27'h00000149, 5'd13, 27'h000003b3, 5'd7, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000015b, 5'd15, 27'h00000044, 5'd17, 27'h000001fe, 32'h00000400,
  1'd1,  5'd23, 27'h000002cc, 5'd12, 27'h00000242, 5'd30, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d3, 5'd21, 27'h000000fb, 5'd8, 27'h0000023f, 32'h00000400,
  1'd1,  5'd22, 27'h000000ad, 5'd22, 27'h000002a2, 5'd16, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000065, 5'd24, 27'h00000112, 5'd30, 27'h000003d5, 32'h00000400,
  1'd1,  5'd1, 27'h000003f2, 5'd8, 27'h0000021e, 5'd1, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003e5, 5'd7, 27'h000000ac, 5'd12, 27'h00000245, 32'h00000400,
  1'd1,  5'd2, 27'h000003c2, 5'd9, 27'h000000f9, 5'd24, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000006b, 5'd17, 27'h0000005f, 5'd4, 27'h00000166, 32'h00000400,
  1'd1,  5'd0, 27'h0000009d, 5'd20, 27'h0000017b, 5'd14, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000015, 5'd16, 27'h000003ed, 5'd21, 27'h00000376, 32'h00000400,
  1'd1,  5'd4, 27'h000003f0, 5'd27, 27'h000000da, 5'd2, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000006e, 5'd28, 27'h00000292, 5'd14, 27'h00000164, 32'h00000400,
  1'd1,  5'd0, 27'h00000200, 5'd29, 27'h000002e8, 5'd22, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000004d, 5'd7, 27'h000000bf, 5'd4, 27'h0000032b, 32'h00000400,
  1'd1,  5'd15, 27'h0000013c, 5'd9, 27'h000001ff, 5'd14, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000039f, 5'd7, 27'h0000009d, 5'd23, 27'h00000327, 32'h00000400,
  1'd1,  5'd10, 27'h000002c4, 5'd17, 27'h00000355, 5'd2, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002bf, 5'd20, 27'h00000220, 5'd13, 27'h0000003f, 32'h00000400,
  1'd1,  5'd10, 27'h00000395, 5'd20, 27'h0000005a, 5'd24, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000293, 5'd27, 27'h00000008, 5'd4, 27'h00000244, 32'h00000400,
  1'd1,  5'd12, 27'h000000de, 5'd27, 27'h000002f1, 5'd14, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000039d, 5'd29, 27'h000000f3, 5'd24, 27'h000003ec, 32'h00000400,
  1'd1,  5'd21, 27'h000003f6, 5'd7, 27'h000002b6, 5'd4, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000327, 5'd8, 27'h0000037b, 5'd12, 27'h000002e1, 32'h00000400,
  1'd1,  5'd24, 27'h00000187, 5'd7, 27'h000001f6, 5'd24, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001cb, 5'd19, 27'h00000383, 5'd2, 27'h0000013e, 32'h00000400,
  1'd1,  5'd21, 27'h000000c3, 5'd18, 27'h00000148, 5'd12, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022c, 5'd15, 27'h000003d1, 5'd23, 27'h0000023e, 32'h00000400,
  1'd1,  5'd21, 27'h00000087, 5'd26, 27'h00000124, 5'd1, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000155, 5'd29, 27'h000002c7, 5'd10, 27'h00000281, 32'h00000400,
  1'd1,  5'd22, 27'h00000082, 5'd30, 27'h000003b5, 5'd25, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002cc, 5'd9, 27'h0000001e, 5'd8, 27'h000000be, 32'h00000400,
  1'd1,  5'd3, 27'h00000132, 5'd6, 27'h00000389, 5'd19, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018f, 5'd7, 27'h000001f6, 5'd26, 27'h0000023b, 32'h00000400,
  1'd1,  5'd2, 27'h00000089, 5'd20, 27'h000000b1, 5'd5, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a2, 5'd19, 27'h000003bc, 5'd18, 27'h00000257, 32'h00000400,
  1'd1,  5'd1, 27'h0000011b, 5'd18, 27'h000003e2, 5'd29, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000352, 5'd25, 27'h000003ff, 5'd5, 27'h0000015c, 32'h00000400,
  1'd1,  5'd1, 27'h000001a9, 5'd26, 27'h000002b5, 5'd19, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d6, 5'd26, 27'h00000199, 5'd27, 27'h000001e1, 32'h00000400,
  1'd1,  5'd14, 27'h00000161, 5'd8, 27'h00000309, 5'd10, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000040, 5'd8, 27'h0000001c, 5'd20, 27'h0000021e, 32'h00000400,
  1'd1,  5'd14, 27'h00000073, 5'd8, 27'h000001da, 5'd29, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003cd, 5'd19, 27'h000000b0, 5'd9, 27'h00000084, 32'h00000400,
  1'd1,  5'd11, 27'h000001d6, 5'd18, 27'h00000032, 5'd18, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000113, 5'd18, 27'h0000011a, 5'd26, 27'h000003ec, 32'h00000400,
  1'd1,  5'd14, 27'h000003eb, 5'd27, 27'h0000011b, 5'd9, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000262, 5'd30, 27'h00000045, 5'd16, 27'h00000330, 32'h00000400,
  1'd1,  5'd12, 27'h0000017c, 5'd26, 27'h000001a4, 5'd29, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000165, 5'd8, 27'h000001f4, 5'd5, 27'h00000229, 32'h00000400,
  1'd1,  5'd24, 27'h0000037b, 5'd6, 27'h00000316, 5'd18, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000109, 5'd10, 27'h00000123, 5'd28, 27'h000000ec, 32'h00000400,
  1'd1,  5'd22, 27'h000001e7, 5'd19, 27'h0000015b, 5'd9, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000012, 5'd19, 27'h0000001f, 5'd17, 27'h00000353, 32'h00000400,
  1'd1,  5'd24, 27'h00000222, 5'd20, 27'h000000e7, 5'd27, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000030b, 5'd26, 27'h00000374, 5'd5, 27'h000000ea, 32'h00000400,
  1'd1,  5'd23, 27'h00000269, 5'd28, 27'h000002e2, 5'd20, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000046, 5'd30, 27'h00000056, 5'd27, 27'h000000fc, 32'h00000400,
  1'd1,  5'd7, 27'h000001a8, 5'd2, 27'h0000010d, 5'd9, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003b5, 5'd2, 27'h000001a0, 5'd16, 27'h000000ae, 32'h00000400,
  1'd1,  5'd6, 27'h00000119, 5'd4, 27'h00000346, 5'd30, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000032d, 5'd15, 27'h0000017d, 5'd4, 27'h000000ad, 32'h00000400,
  1'd1,  5'd7, 27'h000000f0, 5'd14, 27'h00000121, 5'd11, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000203, 5'd11, 27'h0000006e, 5'd21, 27'h0000005e, 32'h00000400,
  1'd1,  5'd6, 27'h00000018, 5'd21, 27'h000000b7, 5'd5, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000006d, 5'd22, 27'h00000217, 5'd14, 27'h0000027f, 32'h00000400,
  1'd1,  5'd6, 27'h000002f5, 5'd21, 27'h000003fd, 5'd25, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000102, 5'd1, 27'h000001be, 5'd7, 27'h00000295, 32'h00000400,
  1'd1,  5'd17, 27'h000002f3, 5'd2, 27'h00000144, 5'd17, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003df, 5'd0, 27'h00000172, 5'd29, 27'h000001b0, 32'h00000400,
  1'd1,  5'd16, 27'h0000035e, 5'd11, 27'h0000011d, 5'd1, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000269, 5'd13, 27'h0000037b, 5'd13, 27'h000003d6, 32'h00000400,
  1'd1,  5'd17, 27'h00000009, 5'd10, 27'h000001d4, 5'd23, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000021e, 5'd20, 27'h0000033c, 5'd3, 27'h000000d2, 32'h00000400,
  1'd1,  5'd15, 27'h00000343, 5'd21, 27'h00000074, 5'd11, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000118, 5'd21, 27'h00000031, 5'd25, 27'h000000a1, 32'h00000400,
  1'd1,  5'd26, 27'h00000358, 5'd1, 27'h00000149, 5'd2, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000050, 5'd2, 27'h0000020e, 5'd12, 27'h000002cb, 32'h00000400,
  1'd1,  5'd26, 27'h00000278, 5'd0, 27'h000000f2, 5'd21, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b8, 5'd15, 27'h000001b4, 5'd2, 27'h0000012b, 32'h00000400,
  1'd1,  5'd29, 27'h00000215, 5'd12, 27'h00000375, 5'd12, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000195, 5'd14, 27'h0000034b, 5'd20, 27'h000002ce, 32'h00000400,
  1'd1,  5'd26, 27'h000000ee, 5'd21, 27'h00000060, 5'd3, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000013b, 5'd22, 27'h0000029c, 5'd11, 27'h0000034d, 32'h00000400,
  1'd1,  5'd28, 27'h00000322, 5'd21, 27'h0000031b, 5'd21, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000329, 5'd2, 27'h000002c8, 5'd1, 27'h00000163, 32'h00000400,
  1'd1,  5'd9, 27'h00000246, 5'd4, 27'h00000152, 5'd13, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ec, 5'd2, 27'h0000009e, 5'd20, 27'h000002f4, 32'h00000400,
  1'd1,  5'd8, 27'h00000244, 5'd10, 27'h000001ca, 5'd5, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003de, 5'd11, 27'h0000003f, 5'd15, 27'h00000386, 32'h00000400,
  1'd1,  5'd10, 27'h00000005, 5'd13, 27'h0000030e, 5'd26, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003c8, 5'd21, 27'h0000011f, 5'd6, 27'h000001c0, 32'h00000400,
  1'd1,  5'd7, 27'h0000036e, 5'd21, 27'h0000007f, 5'd15, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000345, 5'd22, 27'h000001a8, 5'd28, 27'h000000a5, 32'h00000400,
  1'd1,  5'd19, 27'h0000025d, 5'd1, 27'h00000240, 5'd4, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000027c, 5'd4, 27'h0000021f, 5'd10, 27'h00000282, 32'h00000400,
  1'd1,  5'd15, 27'h000003bb, 5'd4, 27'h00000167, 5'd21, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d7, 5'd11, 27'h0000016e, 5'd10, 27'h00000111, 32'h00000400,
  1'd1,  5'd18, 27'h00000155, 5'd10, 27'h00000231, 5'd17, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000095, 5'd13, 27'h00000175, 5'd28, 27'h000000f5, 32'h00000400,
  1'd1,  5'd19, 27'h0000013f, 5'd21, 27'h000002e8, 5'd9, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000350, 5'd24, 27'h000003ae, 5'd18, 27'h0000016e, 32'h00000400,
  1'd1,  5'd19, 27'h000000ce, 5'd24, 27'h000001d8, 5'd27, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000233, 5'd0, 27'h000000b5, 5'd6, 27'h000000c5, 32'h00000400,
  1'd1,  5'd30, 27'h000000a2, 5'd2, 27'h00000367, 5'd16, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000212, 5'd2, 27'h000003e0, 5'd27, 27'h000002aa, 32'h00000400,
  1'd1,  5'd25, 27'h0000036c, 5'd10, 27'h000001f2, 5'd8, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000206, 5'd11, 27'h00000306, 5'd15, 27'h000002eb, 32'h00000400,
  1'd1,  5'd28, 27'h00000023, 5'd13, 27'h0000007c, 5'd26, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000df, 5'd25, 27'h00000125, 5'd6, 27'h0000039e, 32'h00000400,
  1'd1,  5'd26, 27'h0000033b, 5'd23, 27'h0000037d, 5'd16, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000017b, 5'd25, 27'h00000137, 5'd27, 27'h000002d3, 32'h00000400,
  1'd1,  5'd5, 27'h00000343, 5'd6, 27'h000001d7, 5'd4, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000241, 5'd5, 27'h0000036b, 5'd11, 27'h00000148, 32'h00000400,
  1'd1,  5'd7, 27'h00000222, 5'd6, 27'h000002bd, 5'd21, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ea, 5'd17, 27'h00000086, 5'd3, 27'h000003db, 32'h00000400,
  1'd1,  5'd5, 27'h00000176, 5'd17, 27'h000000ab, 5'd13, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b8, 5'd16, 27'h00000148, 5'd23, 27'h00000134, 32'h00000400,
  1'd1,  5'd7, 27'h000000e3, 5'd29, 27'h0000035c, 5'd3, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002fb, 5'd27, 27'h0000035d, 5'd12, 27'h000000b6, 32'h00000400,
  1'd1,  5'd5, 27'h0000038d, 5'd29, 27'h000003aa, 5'd24, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ee, 5'd9, 27'h000003d3, 5'd0, 27'h0000021d, 32'h00000400,
  1'd1,  5'd16, 27'h0000002f, 5'd6, 27'h000001ba, 5'd11, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f3, 5'd10, 27'h00000149, 5'd25, 27'h00000062, 32'h00000400,
  1'd1,  5'd16, 27'h0000016a, 5'd17, 27'h0000000e, 5'd1, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000033, 5'd19, 27'h000000e4, 5'd12, 27'h000002c3, 32'h00000400,
  1'd1,  5'd16, 27'h00000148, 5'd20, 27'h00000009, 5'd25, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000032f, 5'd28, 27'h000000ef, 5'd1, 27'h0000039e, 32'h00000400,
  1'd1,  5'd17, 27'h00000024, 5'd28, 27'h00000313, 5'd12, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000297, 5'd27, 27'h000002c4, 5'd22, 27'h00000149, 32'h00000400,
  1'd1,  5'd28, 27'h0000029d, 5'd9, 27'h000000d3, 5'd4, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000396, 5'd6, 27'h000001e8, 5'd10, 27'h000002f5, 32'h00000400,
  1'd1,  5'd27, 27'h00000110, 5'd9, 27'h000001bb, 5'd23, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000339, 5'd16, 27'h00000330, 5'd2, 27'h00000120, 32'h00000400,
  1'd1,  5'd28, 27'h00000061, 5'd17, 27'h0000011e, 5'd12, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000007a, 5'd19, 27'h000003bc, 5'd22, 27'h00000006, 32'h00000400,
  1'd1,  5'd30, 27'h00000177, 5'd28, 27'h0000031e, 5'd3, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000233, 5'd30, 27'h00000298, 5'd12, 27'h0000039b, 32'h00000400,
  1'd1,  5'd25, 27'h00000373, 5'd26, 27'h000002c1, 5'd21, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e8, 5'd8, 27'h0000037e, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd9, 27'h0000003b, 5'd8, 27'h00000352, 5'd16, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000079, 5'd6, 27'h000000b6, 5'd30, 27'h00000314, 32'h00000400,
  1'd1,  5'd7, 27'h0000003b, 5'd19, 27'h000003d8, 5'd8, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003f, 5'd20, 27'h000001d1, 5'd16, 27'h00000089, 32'h00000400,
  1'd1,  5'd6, 27'h000002ce, 5'd19, 27'h0000001b, 5'd30, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ee, 5'd28, 27'h00000051, 5'd8, 27'h000003cd, 32'h00000400,
  1'd1,  5'd6, 27'h0000006b, 5'd28, 27'h000000c4, 5'd15, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000169, 5'd28, 27'h000002cc, 5'd27, 27'h000003e1, 32'h00000400,
  1'd1,  5'd18, 27'h00000024, 5'd5, 27'h0000026d, 5'd8, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002e6, 5'd10, 27'h00000152, 5'd19, 27'h0000025f, 32'h00000400,
  1'd1,  5'd19, 27'h000001e0, 5'd8, 27'h0000007d, 5'd30, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000138, 5'd20, 27'h000001a1, 5'd8, 27'h00000025, 32'h00000400,
  1'd1,  5'd15, 27'h00000382, 5'd17, 27'h000000e4, 5'd19, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000ba, 5'd15, 27'h000003f3, 5'd29, 27'h00000307, 32'h00000400,
  1'd1,  5'd18, 27'h00000366, 5'd29, 27'h00000146, 5'd7, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000eb, 5'd27, 27'h000000aa, 5'd19, 27'h0000033b, 32'h00000400,
  1'd1,  5'd20, 27'h00000194, 5'd28, 27'h000002b4, 5'd30, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001af, 5'd9, 27'h000002fd, 5'd8, 27'h00000008, 32'h00000400,
  1'd1,  5'd26, 27'h000001ac, 5'd10, 27'h000000f1, 5'd19, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000038f, 5'd5, 27'h000003d6, 5'd28, 27'h000000ba, 32'h00000400,
  1'd1,  5'd29, 27'h00000388, 5'd18, 27'h000000f8, 5'd10, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000005e, 5'd17, 27'h00000110, 5'd15, 27'h00000203, 32'h00000400,
  1'd1,  5'd28, 27'h000003d4, 5'd16, 27'h000003e4, 5'd26, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000035c, 5'd30, 27'h000000b1, 5'd5, 27'h00000323, 32'h00000400,
  1'd1,  5'd28, 27'h00000398, 5'd26, 27'h00000353, 5'd16, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000254, 5'd30, 27'h0000010a, 5'd28, 27'h000001fa, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000005f, 5'd0, 27'h000000a2, 5'd1, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003ae, 5'd1, 27'h00000170, 5'd14, 27'h0000019d, 32'h00000400,
  1'd1,  5'd3, 27'h0000033f, 5'd3, 27'h000001a1, 5'd22, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000279, 5'd11, 27'h00000036, 5'd1, 27'h000001e4, 32'h00000400,
  1'd1,  5'd3, 27'h000001f5, 5'd13, 27'h00000149, 5'd13, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e3, 5'd13, 27'h000000be, 5'd21, 27'h00000025, 32'h00000400,
  1'd1,  5'd2, 27'h000000da, 5'd23, 27'h000003df, 5'd0, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a8, 5'd24, 27'h00000148, 5'd12, 27'h000000b2, 32'h00000400,
  1'd1,  5'd4, 27'h0000002a, 5'd23, 27'h000000e6, 5'd25, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d5, 5'd1, 27'h000001d6, 5'd0, 27'h0000010c, 32'h00000400,
  1'd1,  5'd13, 27'h000001d8, 5'd3, 27'h00000125, 5'd14, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c7, 5'd1, 27'h00000037, 5'd24, 27'h0000008d, 32'h00000400,
  1'd1,  5'd12, 27'h000002b8, 5'd14, 27'h000003f3, 5'd4, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000015, 5'd13, 27'h00000274, 5'd14, 27'h00000079, 32'h00000400,
  1'd1,  5'd10, 27'h000001eb, 5'd11, 27'h00000193, 5'd22, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000039d, 5'd21, 27'h00000232, 5'd3, 27'h000003ac, 32'h00000400,
  1'd1,  5'd13, 27'h000002d1, 5'd20, 27'h00000345, 5'd14, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000020, 5'd22, 27'h00000322, 5'd25, 27'h00000291, 32'h00000400,
  1'd1,  5'd24, 27'h000000e8, 5'd3, 27'h00000380, 5'd4, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000365, 5'd1, 27'h00000186, 5'd12, 27'h000001b0, 32'h00000400,
  1'd1,  5'd23, 27'h000002f6, 5'd2, 27'h00000262, 5'd25, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001d1, 5'd11, 27'h000002d4, 5'd1, 27'h00000043, 32'h00000400,
  1'd1,  5'd21, 27'h00000127, 5'd15, 27'h0000018d, 5'd13, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000379, 5'd12, 27'h0000020b, 5'd20, 27'h0000036a, 32'h00000400,
  1'd1,  5'd21, 27'h000000f9, 5'd20, 27'h000002ce, 5'd0, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000210, 5'd24, 27'h00000188, 5'd15, 27'h000000cb, 32'h00000400,
  1'd1,  5'd22, 27'h000002be, 5'd21, 27'h0000004b, 5'd24, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f1, 5'd4, 27'h000003b7, 5'd6, 27'h0000002a, 32'h00000400,
  1'd1,  5'd3, 27'h000000e3, 5'd3, 27'h0000003a, 5'd17, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000002d, 5'd3, 27'h000003a8, 5'd27, 27'h000000c5, 32'h00000400,
  1'd1,  5'd0, 27'h000001bb, 5'd12, 27'h0000034a, 5'd7, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000240, 5'd10, 27'h000003d6, 5'd16, 27'h0000038c, 32'h00000400,
  1'd1,  5'd1, 27'h00000014, 5'd14, 27'h000000f0, 5'd27, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000342, 5'd21, 27'h00000167, 5'd8, 27'h000001ce, 32'h00000400,
  1'd1,  5'd0, 27'h00000353, 5'd22, 27'h00000100, 5'd16, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000318, 5'd23, 27'h000003d7, 5'd27, 27'h0000000c, 32'h00000400,
  1'd1,  5'd11, 27'h000001a1, 5'd2, 27'h00000034, 5'd6, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000381, 5'd3, 27'h000000f2, 5'd18, 27'h00000197, 32'h00000400,
  1'd1,  5'd13, 27'h0000024f, 5'd2, 27'h0000001f, 5'd26, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000013d, 5'd12, 27'h00000140, 5'd5, 27'h000001c2, 32'h00000400,
  1'd1,  5'd13, 27'h00000381, 5'd15, 27'h0000007a, 5'd15, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000299, 5'd15, 27'h000001fa, 5'd29, 27'h00000167, 32'h00000400,
  1'd1,  5'd10, 27'h0000017e, 5'd22, 27'h000002e0, 5'd9, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c5, 5'd22, 27'h00000313, 5'd16, 27'h00000386, 32'h00000400,
  1'd1,  5'd14, 27'h0000024e, 5'd24, 27'h00000272, 5'd26, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001c9, 5'd2, 27'h000002bc, 5'd8, 27'h0000027c, 32'h00000400,
  1'd1,  5'd24, 27'h0000017b, 5'd3, 27'h000002ea, 5'd16, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000030a, 5'd0, 27'h00000234, 5'd28, 27'h000003e8, 32'h00000400,
  1'd1,  5'd25, 27'h0000008b, 5'd10, 27'h00000292, 5'd7, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d2, 5'd14, 27'h000002db, 5'd18, 27'h000003ab, 32'h00000400,
  1'd1,  5'd21, 27'h0000027f, 5'd11, 27'h00000193, 5'd30, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000360, 5'd21, 27'h0000007b, 5'd9, 27'h000001af, 32'h00000400,
  1'd1,  5'd23, 27'h0000037f, 5'd25, 27'h000001ee, 5'd17, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000009a, 5'd23, 27'h000001ca, 5'd27, 27'h0000031b, 32'h00000400,
  1'd1,  5'd3, 27'h000002bd, 5'd8, 27'h000001b7, 5'd4, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000327, 5'd7, 27'h00000061, 5'd12, 27'h000000e7, 32'h00000400,
  1'd1,  5'd3, 27'h000000eb, 5'd5, 27'h000000ae, 5'd25, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000009c, 5'd17, 27'h0000031b, 5'd1, 27'h000000ce, 32'h00000400,
  1'd1,  5'd3, 27'h00000259, 5'd17, 27'h000000df, 5'd12, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000281, 5'd20, 27'h00000236, 5'd24, 27'h00000359, 32'h00000400,
  1'd1,  5'd2, 27'h000001eb, 5'd28, 27'h00000282, 5'd0, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000019d, 5'd29, 27'h00000190, 5'd12, 27'h0000033d, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd29, 27'h000003c0, 5'd21, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000123, 5'd9, 27'h000003df, 5'd1, 27'h000003f8, 32'h00000400,
  1'd1,  5'd14, 27'h0000000c, 5'd6, 27'h00000233, 5'd10, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000010c, 5'd7, 27'h0000039e, 5'd24, 27'h00000252, 32'h00000400,
  1'd1,  5'd12, 27'h00000356, 5'd16, 27'h0000019b, 5'd4, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001e5, 5'd18, 27'h00000068, 5'd13, 27'h0000002f, 32'h00000400,
  1'd1,  5'd13, 27'h000001d1, 5'd17, 27'h00000220, 5'd24, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000366, 5'd28, 27'h00000209, 5'd0, 27'h0000008d, 32'h00000400,
  1'd1,  5'd12, 27'h000001fe, 5'd28, 27'h000003b3, 5'd11, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e1, 5'd27, 27'h000001d2, 5'd22, 27'h0000003d, 32'h00000400,
  1'd1,  5'd24, 27'h00000059, 5'd9, 27'h00000108, 5'd2, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a6, 5'd8, 27'h000002c2, 5'd13, 27'h000002c8, 32'h00000400,
  1'd1,  5'd24, 27'h0000023e, 5'd6, 27'h000000a9, 5'd25, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000016b, 5'd17, 27'h00000361, 5'd1, 27'h000003db, 32'h00000400,
  1'd1,  5'd23, 27'h000003ec, 5'd15, 27'h000003d2, 5'd11, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000339, 5'd16, 27'h000000e0, 5'd22, 27'h00000196, 32'h00000400,
  1'd1,  5'd21, 27'h00000018, 5'd28, 27'h0000001d, 5'd1, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000276, 5'd26, 27'h000000ed, 5'd13, 27'h0000036d, 32'h00000400,
  1'd1,  5'd20, 27'h0000033c, 5'd25, 27'h000003d4, 5'd24, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000e9, 5'd6, 27'h00000274, 5'd6, 27'h0000038c, 32'h00000400,
  1'd1,  5'd1, 27'h00000112, 5'd6, 27'h00000295, 5'd15, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000eb, 5'd9, 27'h000003fd, 5'd28, 27'h000003c0, 32'h00000400,
  1'd1,  5'd2, 27'h000001ce, 5'd16, 27'h000000e1, 5'd8, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000340, 5'd18, 27'h00000072, 5'd17, 27'h0000016b, 32'h00000400,
  1'd1,  5'd2, 27'h000002ab, 5'd18, 27'h000003f5, 5'd30, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022e, 5'd27, 27'h000000af, 5'd7, 27'h00000397, 32'h00000400,
  1'd1,  5'd3, 27'h000003b8, 5'd29, 27'h00000286, 5'd17, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000022f, 5'd29, 27'h00000256, 5'd28, 27'h00000139, 32'h00000400,
  1'd1,  5'd12, 27'h00000296, 5'd9, 27'h00000097, 5'd7, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001dc, 5'd7, 27'h000000af, 5'd18, 27'h0000007b, 32'h00000400,
  1'd1,  5'd14, 27'h0000014a, 5'd9, 27'h00000328, 5'd28, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000148, 5'd19, 27'h000001d1, 5'd6, 27'h000003a8, 32'h00000400,
  1'd1,  5'd13, 27'h0000009f, 5'd15, 27'h000002bf, 5'd17, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021b, 5'd17, 27'h00000023, 5'd28, 27'h0000034d, 32'h00000400,
  1'd1,  5'd10, 27'h000001ef, 5'd28, 27'h000001ee, 5'd8, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025a, 5'd27, 27'h000002d2, 5'd16, 27'h000002aa, 32'h00000400,
  1'd1,  5'd13, 27'h00000109, 5'd26, 27'h000003e8, 5'd30, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002b2, 5'd9, 27'h000000a7, 5'd6, 27'h00000191, 32'h00000400,
  1'd1,  5'd24, 27'h00000345, 5'd5, 27'h00000139, 5'd17, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000361, 5'd5, 27'h000001e0, 5'd27, 27'h000003be, 32'h00000400,
  1'd1,  5'd25, 27'h00000243, 5'd19, 27'h00000008, 5'd10, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000002b, 5'd16, 27'h00000277, 5'd15, 27'h000003d6, 32'h00000400,
  1'd1,  5'd21, 27'h00000292, 5'd18, 27'h0000027e, 5'd27, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a6, 5'd29, 27'h00000380, 5'd7, 27'h000000e9, 32'h00000400,
  1'd1,  5'd23, 27'h000002d9, 5'd28, 27'h00000132, 5'd19, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001b5, 5'd28, 27'h000002ba, 5'd28, 27'h00000244, 32'h00000400,
  1'd1,  5'd7, 27'h0000002e, 5'd2, 27'h00000288, 5'd9, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e1, 5'd3, 27'h0000021c, 5'd19, 27'h000001d8, 32'h00000400,
  1'd1,  5'd6, 27'h000000b8, 5'd1, 27'h00000292, 5'd30, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000025e, 5'd14, 27'h000003f4, 5'd4, 27'h0000025e, 32'h00000400,
  1'd1,  5'd9, 27'h00000111, 5'd14, 27'h000000eb, 5'd13, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002fa, 5'd14, 27'h00000019, 5'd22, 27'h00000127, 32'h00000400,
  1'd1,  5'd8, 27'h00000189, 5'd20, 27'h00000338, 5'd4, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000008e, 5'd24, 27'h0000011a, 5'd15, 27'h00000033, 32'h00000400,
  1'd1,  5'd5, 27'h000001e5, 5'd22, 27'h00000337, 5'd22, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a8, 5'd3, 27'h000003fc, 5'd6, 27'h00000245, 32'h00000400,
  1'd1,  5'd18, 27'h000000f8, 5'd2, 27'h00000067, 5'd17, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003c3, 5'd4, 27'h000002ee, 5'd27, 27'h00000019, 32'h00000400,
  1'd1,  5'd16, 27'h00000221, 5'd13, 27'h000001da, 5'd3, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003a4, 5'd15, 27'h000001c2, 5'd13, 27'h000001b6, 32'h00000400,
  1'd1,  5'd19, 27'h0000003d, 5'd11, 27'h0000019c, 5'd21, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000334, 5'd25, 27'h000001b5, 5'd3, 27'h0000003f, 32'h00000400,
  1'd1,  5'd17, 27'h000002a6, 5'd24, 27'h000003b3, 5'd11, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000283, 5'd22, 27'h000000a4, 5'd23, 27'h000003a4, 32'h00000400,
  1'd1,  5'd28, 27'h000000e6, 5'd2, 27'h00000165, 5'd1, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000128, 5'd5, 27'h0000007d, 5'd15, 27'h00000167, 32'h00000400,
  1'd1,  5'd25, 27'h000003fa, 5'd1, 27'h000001d0, 5'd23, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b5, 5'd11, 27'h000000ae, 5'd4, 27'h00000007, 32'h00000400,
  1'd1,  5'd29, 27'h00000057, 5'd12, 27'h000000dc, 5'd12, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000378, 5'd13, 27'h0000007a, 5'd24, 27'h0000013e, 32'h00000400,
  1'd1,  5'd26, 27'h0000023b, 5'd25, 27'h000000ae, 5'd2, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000382, 5'd21, 27'h0000013c, 5'd14, 27'h00000114, 32'h00000400,
  1'd1,  5'd28, 27'h00000035, 5'd22, 27'h000000b2, 5'd25, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003de, 5'd4, 27'h000001cf, 5'd3, 27'h000003c9, 32'h00000400,
  1'd1,  5'd8, 27'h000003dc, 5'd2, 27'h0000028c, 5'd12, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002aa, 5'd4, 27'h00000374, 5'd25, 27'h00000276, 32'h00000400,
  1'd1,  5'd8, 27'h0000028a, 5'd10, 27'h00000362, 5'd8, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ca, 5'd15, 27'h00000076, 5'd17, 27'h00000188, 32'h00000400,
  1'd1,  5'd6, 27'h00000241, 5'd13, 27'h0000022a, 5'd27, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000137, 5'd21, 27'h00000100, 5'd7, 27'h0000016f, 32'h00000400,
  1'd1,  5'd9, 27'h00000155, 5'd21, 27'h00000339, 5'd19, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000105, 5'd23, 27'h000001f4, 5'd28, 27'h0000014c, 32'h00000400,
  1'd1,  5'd19, 27'h00000233, 5'd2, 27'h00000293, 5'd2, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000353, 5'd1, 27'h00000138, 5'd10, 27'h0000033e, 32'h00000400,
  1'd1,  5'd16, 27'h0000022b, 5'd0, 27'h000001b2, 5'd22, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000232, 5'd12, 27'h00000376, 5'd6, 27'h0000019e, 32'h00000400,
  1'd1,  5'd18, 27'h0000034b, 5'd11, 27'h0000022b, 5'd15, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000331, 5'd10, 27'h000001b3, 5'd26, 27'h0000007a, 32'h00000400,
  1'd1,  5'd19, 27'h000001c4, 5'd21, 27'h000000b4, 5'd7, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000076, 5'd23, 27'h000000bc, 5'd16, 27'h000001bc, 32'h00000400,
  1'd1,  5'd20, 27'h000001e5, 5'd24, 27'h0000035c, 5'd30, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000258, 5'd0, 27'h0000025d, 5'd6, 27'h000002aa, 32'h00000400,
  1'd1,  5'd26, 27'h000002b4, 5'd4, 27'h0000025c, 5'd15, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f6, 5'd0, 27'h000000e8, 5'd27, 27'h0000004b, 32'h00000400,
  1'd1,  5'd26, 27'h000001b6, 5'd14, 27'h0000027d, 5'd7, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000022b, 5'd11, 27'h000003dd, 5'd20, 27'h000000fb, 32'h00000400,
  1'd1,  5'd25, 27'h0000036d, 5'd12, 27'h00000163, 5'd28, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000019f, 5'd25, 27'h0000003e, 5'd10, 27'h00000112, 32'h00000400,
  1'd1,  5'd29, 27'h000002b2, 5'd20, 27'h000002e7, 5'd18, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a4, 5'd24, 27'h00000134, 5'd30, 27'h0000008b, 32'h00000400,
  1'd1,  5'd9, 27'h00000282, 5'd6, 27'h0000017b, 5'd0, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000013, 5'd7, 27'h000003cd, 5'd13, 27'h000003e7, 32'h00000400,
  1'd1,  5'd7, 27'h00000098, 5'd5, 27'h000000b2, 5'd23, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012f, 5'd16, 27'h0000006d, 5'd0, 27'h000001fa, 32'h00000400,
  1'd1,  5'd9, 27'h0000023f, 5'd16, 27'h00000162, 5'd11, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000017e, 5'd19, 27'h0000012d, 5'd22, 27'h0000000f, 32'h00000400,
  1'd1,  5'd6, 27'h0000037e, 5'd28, 27'h00000309, 5'd4, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000115, 5'd28, 27'h00000247, 5'd10, 27'h00000200, 32'h00000400,
  1'd1,  5'd7, 27'h000002b0, 5'd29, 27'h00000385, 5'd23, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003bd, 5'd10, 27'h00000042, 5'd4, 27'h000001a1, 32'h00000400,
  1'd1,  5'd18, 27'h0000009a, 5'd9, 27'h00000098, 5'd12, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000011a, 5'd9, 27'h00000156, 5'd23, 27'h0000016d, 32'h00000400,
  1'd1,  5'd18, 27'h00000215, 5'd19, 27'h0000039d, 5'd0, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ed, 5'd18, 27'h0000032d, 5'd10, 27'h0000038f, 32'h00000400,
  1'd1,  5'd15, 27'h00000374, 5'd20, 27'h00000204, 5'd22, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003f6, 5'd27, 27'h000001b5, 5'd1, 27'h0000021a, 32'h00000400,
  1'd1,  5'd18, 27'h0000020b, 5'd27, 27'h00000168, 5'd11, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000199, 5'd29, 27'h000000d5, 5'd22, 27'h000003f8, 32'h00000400,
  1'd1,  5'd29, 27'h00000113, 5'd6, 27'h00000116, 5'd2, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d6, 5'd10, 27'h0000007f, 5'd11, 27'h00000351, 32'h00000400,
  1'd1,  5'd30, 27'h000003fd, 5'd9, 27'h00000293, 5'd22, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003e9, 5'd17, 27'h0000011a, 5'd0, 27'h0000021e, 32'h00000400,
  1'd1,  5'd27, 27'h0000033f, 5'd19, 27'h000003e7, 5'd13, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000036, 5'd20, 27'h0000016a, 5'd24, 27'h000000e1, 32'h00000400,
  1'd1,  5'd29, 27'h00000004, 5'd30, 27'h00000364, 5'd3, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000257, 5'd29, 27'h00000018, 5'd10, 27'h000002fb, 32'h00000400,
  1'd1,  5'd29, 27'h00000113, 5'd28, 27'h000001c3, 5'd24, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a5, 5'd6, 27'h000001e2, 5'd9, 27'h00000076, 32'h00000400,
  1'd1,  5'd8, 27'h00000352, 5'd9, 27'h000002b4, 5'd18, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000013e, 5'd9, 27'h00000287, 5'd25, 27'h00000392, 32'h00000400,
  1'd1,  5'd10, 27'h00000039, 5'd17, 27'h0000001d, 5'd6, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000096, 5'd20, 27'h000001d3, 5'd17, 27'h0000002f, 32'h00000400,
  1'd1,  5'd9, 27'h000001fd, 5'd17, 27'h000000c7, 5'd27, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000020b, 5'd30, 27'h000002d9, 5'd8, 27'h0000026e, 32'h00000400,
  1'd1,  5'd6, 27'h00000138, 5'd26, 27'h000001ce, 5'd16, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001c8, 5'd27, 27'h0000030d, 5'd29, 27'h00000006, 32'h00000400,
  1'd1,  5'd17, 27'h0000033a, 5'd6, 27'h000002a8, 5'd9, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000261, 5'd8, 27'h000002da, 5'd17, 27'h00000189, 32'h00000400,
  1'd1,  5'd18, 27'h00000270, 5'd6, 27'h000000b0, 5'd27, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000191, 5'd20, 27'h00000033, 5'd10, 27'h00000045, 32'h00000400,
  1'd1,  5'd20, 27'h00000216, 5'd19, 27'h000000ea, 5'd19, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003e1, 5'd19, 27'h0000038c, 5'd26, 27'h0000010b, 32'h00000400,
  1'd1,  5'd16, 27'h00000116, 5'd26, 27'h00000196, 5'd6, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000244, 5'd27, 27'h000000c0, 5'd19, 27'h0000003d, 32'h00000400,
  1'd1,  5'd16, 27'h000001f5, 5'd28, 27'h000003ba, 5'd29, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000226, 5'd7, 27'h00000394, 5'd6, 27'h000000de, 32'h00000400,
  1'd1,  5'd28, 27'h0000017b, 5'd5, 27'h000001f7, 5'd15, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002af, 5'd8, 27'h00000008, 5'd26, 27'h000002eb, 32'h00000400,
  1'd1,  5'd28, 27'h000001ce, 5'd19, 27'h0000030d, 5'd7, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000034e, 5'd16, 27'h000001c0, 5'd19, 27'h0000013d, 32'h00000400,
  1'd1,  5'd26, 27'h000002e1, 5'd18, 27'h00000027, 5'd26, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000005d, 5'd26, 27'h00000188, 5'd6, 27'h00000326, 32'h00000400,
  1'd1,  5'd30, 27'h0000019d, 5'd27, 27'h00000193, 5'd18, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000017c, 5'd29, 27'h00000253, 5'd28, 27'h0000006d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000085, 5'd1, 27'h000001f4, 5'd2, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000178, 5'd2, 27'h00000034, 5'd13, 27'h000002b2, 32'h00000400,
  1'd1,  5'd0, 27'h00000277, 5'd2, 27'h000002fd, 5'd24, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000013e, 5'd13, 27'h000001ce, 5'd0, 27'h00000291, 32'h00000400,
  1'd1,  5'd2, 27'h00000065, 5'd11, 27'h00000170, 5'd10, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000388, 5'd10, 27'h000003e6, 5'd24, 27'h00000330, 32'h00000400,
  1'd1,  5'd0, 27'h00000275, 5'd20, 27'h000003ba, 5'd0, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017e, 5'd25, 27'h000000a7, 5'd15, 27'h00000136, 32'h00000400,
  1'd1,  5'd4, 27'h000001e3, 5'd25, 27'h000000a8, 5'd24, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c4, 5'd2, 27'h00000057, 5'd2, 27'h00000187, 32'h00000400,
  1'd1,  5'd14, 27'h00000351, 5'd1, 27'h00000066, 5'd10, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000030f, 5'd1, 27'h000003cf, 5'd24, 27'h0000011d, 32'h00000400,
  1'd1,  5'd11, 27'h00000245, 5'd15, 27'h0000015f, 5'd2, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c7, 5'd11, 27'h00000051, 5'd12, 27'h0000020f, 32'h00000400,
  1'd1,  5'd14, 27'h00000025, 5'd13, 27'h00000232, 5'd20, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000016, 5'd24, 27'h000001df, 5'd4, 27'h00000382, 32'h00000400,
  1'd1,  5'd14, 27'h000001a0, 5'd21, 27'h000001b1, 5'd14, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ae, 5'd22, 27'h0000009a, 5'd25, 27'h000001a2, 32'h00000400,
  1'd1,  5'd22, 27'h0000026a, 5'd3, 27'h000000cd, 5'd3, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ec, 5'd1, 27'h00000007, 5'd14, 27'h00000052, 32'h00000400,
  1'd1,  5'd25, 27'h00000341, 5'd0, 27'h00000160, 5'd22, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000f7, 5'd13, 27'h00000390, 5'd3, 27'h00000047, 32'h00000400,
  1'd1,  5'd22, 27'h000002f2, 5'd14, 27'h00000396, 5'd10, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b1, 5'd14, 27'h000000ff, 5'd22, 27'h0000008c, 32'h00000400,
  1'd1,  5'd20, 27'h000003a5, 5'd24, 27'h0000005b, 5'd4, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a5, 5'd24, 27'h000000c9, 5'd15, 27'h0000012d, 32'h00000400,
  1'd1,  5'd24, 27'h0000023a, 5'd20, 27'h00000317, 5'd22, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000348, 5'd0, 27'h00000322, 5'd9, 27'h000001b0, 32'h00000400,
  1'd1,  5'd5, 27'h00000069, 5'd2, 27'h0000039f, 5'd16, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ab, 5'd2, 27'h00000322, 5'd25, 27'h00000376, 32'h00000400,
  1'd1,  5'd1, 27'h00000339, 5'd12, 27'h0000039d, 5'd7, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000039, 5'd11, 27'h00000307, 5'd17, 27'h000000e4, 32'h00000400,
  1'd1,  5'd3, 27'h0000003c, 5'd12, 27'h000001dd, 5'd29, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000019e, 5'd23, 27'h00000259, 5'd8, 27'h0000039f, 32'h00000400,
  1'd1,  5'd4, 27'h0000016d, 5'd21, 27'h00000338, 5'd20, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000008d, 5'd21, 27'h0000018d, 5'd29, 27'h0000016a, 32'h00000400,
  1'd1,  5'd10, 27'h000003ac, 5'd0, 27'h0000008f, 5'd7, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000025e, 5'd1, 27'h000002a1, 5'd17, 27'h00000274, 32'h00000400,
  1'd1,  5'd15, 27'h0000013a, 5'd2, 27'h00000363, 5'd27, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000d0, 5'd13, 27'h0000028e, 5'd9, 27'h00000282, 32'h00000400,
  1'd1,  5'd11, 27'h000003ed, 5'd12, 27'h0000006d, 5'd19, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000175, 5'd13, 27'h0000025d, 5'd28, 27'h00000215, 32'h00000400,
  1'd1,  5'd13, 27'h00000331, 5'd25, 27'h00000191, 5'd7, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003a7, 5'd21, 27'h000001eb, 5'd17, 27'h0000035e, 32'h00000400,
  1'd1,  5'd14, 27'h000001b0, 5'd23, 27'h000002dd, 5'd27, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d6, 5'd2, 27'h000003a4, 5'd7, 27'h000000cc, 32'h00000400,
  1'd1,  5'd25, 27'h000001ea, 5'd4, 27'h00000304, 5'd20, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000240, 5'd0, 27'h000001ac, 5'd27, 27'h0000015b, 32'h00000400,
  1'd1,  5'd22, 27'h0000038a, 5'd12, 27'h00000107, 5'd10, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b3, 5'd13, 27'h000003ee, 5'd18, 27'h00000165, 32'h00000400,
  1'd1,  5'd22, 27'h000003a4, 5'd12, 27'h0000014c, 5'd26, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000024b, 5'd21, 27'h000003ac, 5'd7, 27'h00000275, 32'h00000400,
  1'd1,  5'd20, 27'h000002ac, 5'd25, 27'h00000325, 5'd18, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001eb, 5'd22, 27'h000002e3, 5'd25, 27'h000003a1, 32'h00000400,
  1'd1,  5'd3, 27'h000003ec, 5'd5, 27'h000000fe, 5'd2, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000002a, 5'd8, 27'h00000042, 5'd13, 27'h000000d0, 32'h00000400,
  1'd1,  5'd1, 27'h00000037, 5'd5, 27'h000002aa, 5'd21, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000275, 5'd15, 27'h00000241, 5'd3, 27'h000000fe, 32'h00000400,
  1'd1,  5'd1, 27'h0000035a, 5'd16, 27'h000002cb, 5'd13, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000013c, 5'd17, 27'h000001fe, 5'd21, 27'h000000c0, 32'h00000400,
  1'd1,  5'd3, 27'h0000023c, 5'd28, 27'h0000020a, 5'd1, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002cc, 5'd27, 27'h0000009e, 5'd10, 27'h000002ca, 32'h00000400,
  1'd1,  5'd0, 27'h0000025d, 5'd29, 27'h0000029e, 5'd21, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000102, 5'd5, 27'h00000155, 5'd2, 27'h000002dc, 32'h00000400,
  1'd1,  5'd10, 27'h0000028b, 5'd8, 27'h00000195, 5'd12, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000037a, 5'd7, 27'h0000031d, 5'd23, 27'h0000026f, 32'h00000400,
  1'd1,  5'd15, 27'h000000a8, 5'd19, 27'h00000394, 5'd1, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001a9, 5'd18, 27'h00000207, 5'd13, 27'h00000104, 32'h00000400,
  1'd1,  5'd12, 27'h00000262, 5'd19, 27'h00000041, 5'd23, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000253, 5'd29, 27'h000001bb, 5'd3, 27'h0000001a, 32'h00000400,
  1'd1,  5'd10, 27'h00000193, 5'd28, 27'h00000305, 5'd12, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000031, 5'd29, 27'h000003fb, 5'd23, 27'h0000038b, 32'h00000400,
  1'd1,  5'd21, 27'h0000026b, 5'd9, 27'h0000005f, 5'd3, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000fa, 5'd6, 27'h00000335, 5'd14, 27'h00000218, 32'h00000400,
  1'd1,  5'd21, 27'h0000000c, 5'd8, 27'h000002d2, 5'd21, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000037f, 5'd19, 27'h000003ff, 5'd4, 27'h0000016a, 32'h00000400,
  1'd1,  5'd22, 27'h00000227, 5'd20, 27'h00000124, 5'd11, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001b9, 5'd16, 27'h000001e9, 5'd25, 27'h00000082, 32'h00000400,
  1'd1,  5'd22, 27'h00000097, 5'd28, 27'h000003cb, 5'd4, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000331, 5'd26, 27'h00000100, 5'd11, 27'h000003f2, 32'h00000400,
  1'd1,  5'd23, 27'h0000007c, 5'd28, 27'h0000008c, 5'd25, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000210, 5'd8, 27'h00000185, 5'd8, 27'h000001bc, 32'h00000400,
  1'd1,  5'd4, 27'h0000008a, 5'd6, 27'h000003bd, 5'd17, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b5, 5'd6, 27'h00000243, 5'd30, 27'h0000020b, 32'h00000400,
  1'd1,  5'd2, 27'h000002d5, 5'd16, 27'h00000385, 5'd9, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e1, 5'd18, 27'h0000030f, 5'd19, 27'h000001f8, 32'h00000400,
  1'd1,  5'd2, 27'h000000ba, 5'd18, 27'h000003a9, 5'd26, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000161, 5'd27, 27'h000001df, 5'd5, 27'h00000362, 32'h00000400,
  1'd1,  5'd1, 27'h000003f5, 5'd25, 27'h00000374, 5'd15, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000fa, 5'd27, 27'h00000075, 5'd27, 27'h0000023e, 32'h00000400,
  1'd1,  5'd15, 27'h000001d1, 5'd10, 27'h00000130, 5'd9, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000246, 5'd10, 27'h0000004b, 5'd18, 27'h00000002, 32'h00000400,
  1'd1,  5'd12, 27'h0000005f, 5'd9, 27'h000000b5, 5'd28, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011d, 5'd19, 27'h00000003, 5'd7, 27'h00000040, 32'h00000400,
  1'd1,  5'd13, 27'h000000a8, 5'd19, 27'h0000032a, 5'd19, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ca, 5'd16, 27'h00000378, 5'd30, 27'h0000009b, 32'h00000400,
  1'd1,  5'd14, 27'h0000030f, 5'd30, 27'h00000324, 5'd8, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d8, 5'd30, 27'h000001cf, 5'd17, 27'h000000f6, 32'h00000400,
  1'd1,  5'd14, 27'h0000015b, 5'd30, 27'h00000292, 5'd26, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c8, 5'd9, 27'h00000184, 5'd8, 27'h00000165, 32'h00000400,
  1'd1,  5'd21, 27'h000002ae, 5'd5, 27'h000002c7, 5'd15, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f7, 5'd5, 27'h00000127, 5'd28, 27'h00000228, 32'h00000400,
  1'd1,  5'd23, 27'h000002af, 5'd17, 27'h00000063, 5'd6, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000021f, 5'd17, 27'h00000231, 5'd19, 27'h00000017, 32'h00000400,
  1'd1,  5'd23, 27'h0000005e, 5'd17, 27'h00000073, 5'd26, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e4, 5'd30, 27'h000001c5, 5'd9, 27'h00000163, 32'h00000400,
  1'd1,  5'd23, 27'h00000047, 5'd26, 27'h0000018a, 5'd19, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ff, 5'd29, 27'h00000159, 5'd28, 27'h00000211, 32'h00000400,
  1'd1,  5'd9, 27'h0000016c, 5'd3, 27'h0000019c, 5'd6, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000007b, 5'd3, 27'h000003f4, 5'd19, 27'h00000113, 32'h00000400,
  1'd1,  5'd8, 27'h00000110, 5'd1, 27'h00000068, 5'd30, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d7, 5'd10, 27'h00000263, 5'd2, 27'h000003e3, 32'h00000400,
  1'd1,  5'd9, 27'h000000e0, 5'd12, 27'h00000056, 5'd11, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000018d, 5'd11, 27'h00000302, 5'd25, 27'h00000048, 32'h00000400,
  1'd1,  5'd5, 27'h000003e6, 5'd24, 27'h000000cb, 5'd4, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000022d, 5'd24, 27'h000001fe, 5'd12, 27'h0000013b, 32'h00000400,
  1'd1,  5'd6, 27'h00000227, 5'd21, 27'h000002fd, 5'd22, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f7, 5'd4, 27'h000001a5, 5'd8, 27'h000002c0, 32'h00000400,
  1'd1,  5'd16, 27'h000000b8, 5'd4, 27'h000000d3, 5'd15, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ef, 5'd2, 27'h0000017a, 5'd26, 27'h000002a9, 32'h00000400,
  1'd1,  5'd20, 27'h00000025, 5'd12, 27'h000002b5, 5'd4, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000be, 5'd13, 27'h000003f1, 5'd15, 27'h0000005d, 32'h00000400,
  1'd1,  5'd20, 27'h0000008c, 5'd14, 27'h000002ce, 5'd21, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000104, 5'd25, 27'h000001bf, 5'd1, 27'h000002aa, 32'h00000400,
  1'd1,  5'd20, 27'h000001b2, 5'd21, 27'h0000015e, 5'd11, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000074, 5'd20, 27'h000003a1, 5'd23, 27'h00000392, 32'h00000400,
  1'd1,  5'd28, 27'h00000377, 5'd3, 27'h0000002b, 5'd2, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000277, 5'd5, 27'h00000013, 5'd15, 27'h0000011f, 32'h00000400,
  1'd1,  5'd26, 27'h000002b9, 5'd1, 27'h0000019d, 5'd23, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000315, 5'd11, 27'h000001a7, 5'd2, 27'h00000154, 32'h00000400,
  1'd1,  5'd29, 27'h000002fe, 5'd12, 27'h000002ed, 5'd11, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000079, 5'd12, 27'h00000377, 5'd25, 27'h00000348, 32'h00000400,
  1'd1,  5'd27, 27'h0000037a, 5'd21, 27'h000002ae, 5'd3, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000063, 5'd24, 27'h000001b3, 5'd14, 27'h000000a6, 32'h00000400,
  1'd1,  5'd28, 27'h0000001b, 5'd24, 27'h0000017f, 5'd24, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000038d, 5'd4, 27'h000000d0, 5'd1, 27'h0000023a, 32'h00000400,
  1'd1,  5'd10, 27'h000000e5, 5'd0, 27'h000003a4, 5'd11, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e1, 5'd4, 27'h000000ee, 5'd22, 27'h00000037, 32'h00000400,
  1'd1,  5'd7, 27'h000001bf, 5'd14, 27'h00000056, 5'd7, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a3, 5'd15, 27'h00000189, 5'd16, 27'h000000cb, 32'h00000400,
  1'd1,  5'd10, 27'h00000144, 5'd14, 27'h00000201, 5'd30, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e2, 5'd24, 27'h00000370, 5'd9, 27'h000002b5, 32'h00000400,
  1'd1,  5'd6, 27'h000002bd, 5'd24, 27'h000003c1, 5'd17, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000a5, 5'd23, 27'h00000065, 5'd27, 27'h000000d7, 32'h00000400,
  1'd1,  5'd15, 27'h0000031a, 5'd4, 27'h00000070, 5'd4, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000157, 5'd3, 27'h00000090, 5'd10, 27'h00000308, 32'h00000400,
  1'd1,  5'd20, 27'h00000091, 5'd2, 27'h0000034d, 5'd21, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000092, 5'd12, 27'h000002b5, 5'd9, 27'h0000013d, 32'h00000400,
  1'd1,  5'd19, 27'h000002b4, 5'd13, 27'h000001b0, 5'd18, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000266, 5'd11, 27'h00000170, 5'd30, 27'h00000354, 32'h00000400,
  1'd1,  5'd18, 27'h0000006f, 5'd25, 27'h0000025e, 5'd8, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000038, 5'd22, 27'h000001bb, 5'd20, 27'h0000009e, 32'h00000400,
  1'd1,  5'd19, 27'h0000005c, 5'd22, 27'h00000152, 5'd26, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d4, 5'd2, 27'h0000035a, 5'd6, 27'h000001f7, 32'h00000400,
  1'd1,  5'd27, 27'h0000011b, 5'd2, 27'h00000044, 5'd19, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000063, 5'd2, 27'h0000007f, 5'd26, 27'h000002ce, 32'h00000400,
  1'd1,  5'd27, 27'h000003c3, 5'd11, 27'h00000376, 5'd8, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003cd, 5'd10, 27'h000002dd, 5'd18, 27'h00000078, 32'h00000400,
  1'd1,  5'd26, 27'h0000032e, 5'd11, 27'h00000092, 5'd29, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ee, 5'd24, 27'h00000052, 5'd9, 27'h0000016e, 32'h00000400,
  1'd1,  5'd26, 27'h000001c1, 5'd20, 27'h000002e7, 5'd15, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000248, 5'd25, 27'h00000135, 5'd30, 27'h00000145, 32'h00000400,
  1'd1,  5'd10, 27'h00000007, 5'd8, 27'h00000396, 5'd0, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001aa, 5'd10, 27'h00000010, 5'd14, 27'h000000cc, 32'h00000400,
  1'd1,  5'd10, 27'h00000138, 5'd7, 27'h0000011b, 5'd22, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c4, 5'd17, 27'h000003e1, 5'd4, 27'h000002be, 32'h00000400,
  1'd1,  5'd9, 27'h0000028d, 5'd17, 27'h0000012f, 5'd14, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000093, 5'd16, 27'h00000023, 5'd24, 27'h000003c8, 32'h00000400,
  1'd1,  5'd10, 27'h00000052, 5'd28, 27'h00000318, 5'd1, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000212, 5'd30, 27'h000002f3, 5'd15, 27'h000000de, 32'h00000400,
  1'd1,  5'd7, 27'h0000002c, 5'd26, 27'h000000d1, 5'd25, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003b0, 5'd9, 27'h00000327, 5'd4, 27'h000003a0, 32'h00000400,
  1'd1,  5'd16, 27'h0000030f, 5'd5, 27'h00000274, 5'd11, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000232, 5'd7, 27'h00000312, 5'd24, 27'h0000023b, 32'h00000400,
  1'd1,  5'd18, 27'h00000342, 5'd18, 27'h00000102, 5'd2, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000db, 5'd19, 27'h000001d3, 5'd14, 27'h00000291, 32'h00000400,
  1'd1,  5'd20, 27'h00000088, 5'd19, 27'h00000101, 5'd21, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f7, 5'd27, 27'h000002e2, 5'd1, 27'h0000034b, 32'h00000400,
  1'd1,  5'd16, 27'h00000279, 5'd29, 27'h00000367, 5'd10, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000027, 5'd29, 27'h00000050, 5'd22, 27'h000002d0, 32'h00000400,
  1'd1,  5'd27, 27'h0000030b, 5'd10, 27'h00000058, 5'd4, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000011f, 5'd8, 27'h0000001f, 5'd15, 27'h00000055, 32'h00000400,
  1'd1,  5'd26, 27'h000003e7, 5'd7, 27'h0000034e, 5'd23, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000fa, 5'd16, 27'h000001d9, 5'd3, 27'h00000072, 32'h00000400,
  1'd1,  5'd27, 27'h00000236, 5'd19, 27'h0000030a, 5'd12, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000013b, 5'd15, 27'h00000307, 5'd25, 27'h000002e3, 32'h00000400,
  1'd1,  5'd27, 27'h0000017a, 5'd27, 27'h0000012f, 5'd3, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000fa, 5'd28, 27'h000000d4, 5'd14, 27'h00000262, 32'h00000400,
  1'd1,  5'd30, 27'h0000013c, 5'd30, 27'h00000247, 5'd22, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000296, 5'd6, 27'h000002fb, 5'd8, 27'h0000010e, 32'h00000400,
  1'd1,  5'd8, 27'h0000016e, 5'd7, 27'h000003aa, 5'd20, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000212, 5'd5, 27'h0000020b, 5'd25, 27'h0000037a, 32'h00000400,
  1'd1,  5'd6, 27'h0000028f, 5'd20, 27'h000000f5, 5'd7, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c9, 5'd18, 27'h0000016a, 5'd17, 27'h000003ac, 32'h00000400,
  1'd1,  5'd9, 27'h000003cc, 5'd16, 27'h00000080, 5'd29, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000009d, 5'd27, 27'h000001a7, 5'd10, 27'h0000013b, 32'h00000400,
  1'd1,  5'd8, 27'h00000359, 5'd26, 27'h000002e5, 5'd18, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a5, 5'd27, 27'h00000029, 5'd27, 27'h000002c8, 32'h00000400,
  1'd1,  5'd19, 27'h00000184, 5'd10, 27'h00000044, 5'd6, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039d, 5'd9, 27'h000003ca, 5'd15, 27'h00000233, 32'h00000400,
  1'd1,  5'd18, 27'h000003d6, 5'd7, 27'h0000007f, 5'd28, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000152, 5'd15, 27'h00000269, 5'd6, 27'h000000c0, 32'h00000400,
  1'd1,  5'd19, 27'h00000282, 5'd16, 27'h00000074, 5'd18, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000018c, 5'd17, 27'h000002a4, 5'd26, 27'h0000005e, 32'h00000400,
  1'd1,  5'd17, 27'h00000259, 5'd26, 27'h000003d6, 5'd7, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a9, 5'd28, 27'h000000b5, 5'd20, 27'h0000024e, 32'h00000400,
  1'd1,  5'd19, 27'h000000e7, 5'd27, 27'h00000086, 5'd28, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000205, 5'd6, 27'h00000295, 5'd7, 27'h000000fd, 32'h00000400,
  1'd1,  5'd28, 27'h00000346, 5'd6, 27'h000001be, 5'd17, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c7, 5'd9, 27'h00000142, 5'd25, 27'h000003a8, 32'h00000400,
  1'd1,  5'd29, 27'h000001e7, 5'd17, 27'h00000231, 5'd6, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001db, 5'd16, 27'h00000315, 5'd20, 27'h0000028c, 32'h00000400,
  1'd1,  5'd27, 27'h0000010e, 5'd15, 27'h00000286, 5'd29, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000c7, 5'd29, 27'h000003f4, 5'd8, 27'h0000020e, 32'h00000400,
  1'd1,  5'd25, 27'h000003f5, 5'd30, 27'h000000d3, 5'd19, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000149, 5'd27, 27'h00000278, 5'd26, 27'h0000001a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000187, 5'd4, 27'h0000032c, 5'd2, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000002, 5'd2, 27'h00000212, 5'd12, 27'h0000006b, 32'h00000400,
  1'd1,  5'd2, 27'h00000259, 5'd2, 27'h000003cb, 5'd22, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000106, 5'd12, 27'h000003b1, 5'd3, 27'h000003aa, 32'h00000400,
  1'd1,  5'd2, 27'h000003cb, 5'd12, 27'h000000e2, 5'd12, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a8, 5'd11, 27'h0000021a, 5'd21, 27'h00000119, 32'h00000400,
  1'd1,  5'd4, 27'h000002e7, 5'd23, 27'h000001c7, 5'd1, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000033, 5'd20, 27'h000002dd, 5'd12, 27'h00000010, 32'h00000400,
  1'd1,  5'd2, 27'h00000218, 5'd21, 27'h0000039a, 5'd24, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000351, 5'd2, 27'h0000009c, 5'd3, 27'h0000037c, 32'h00000400,
  1'd1,  5'd15, 27'h0000000b, 5'd3, 27'h00000232, 5'd11, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000281, 5'd2, 27'h0000033e, 5'd22, 27'h000001ec, 32'h00000400,
  1'd1,  5'd14, 27'h00000144, 5'd12, 27'h0000030e, 5'd1, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000009e, 5'd13, 27'h0000002a, 5'd11, 27'h000003ff, 32'h00000400,
  1'd1,  5'd11, 27'h0000032c, 5'd14, 27'h00000103, 5'd22, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f8, 5'd25, 27'h00000298, 5'd4, 27'h0000039f, 32'h00000400,
  1'd1,  5'd10, 27'h000003b8, 5'd23, 27'h000003b0, 5'd14, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001d0, 5'd24, 27'h00000314, 5'd23, 27'h000001d4, 32'h00000400,
  1'd1,  5'd25, 27'h00000160, 5'd0, 27'h00000059, 5'd3, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000375, 5'd3, 27'h00000264, 5'd15, 27'h00000127, 32'h00000400,
  1'd1,  5'd23, 27'h000000ed, 5'd3, 27'h00000324, 5'd22, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000359, 5'd14, 27'h000000d7, 5'd0, 27'h00000102, 32'h00000400,
  1'd1,  5'd22, 27'h000003bb, 5'd15, 27'h000000e6, 5'd13, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003b1, 5'd15, 27'h00000128, 5'd25, 27'h0000002a, 32'h00000400,
  1'd1,  5'd23, 27'h0000002d, 5'd21, 27'h00000285, 5'd0, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000016, 5'd21, 27'h00000103, 5'd14, 27'h000000ff, 32'h00000400,
  1'd1,  5'd21, 27'h0000002e, 5'd24, 27'h00000074, 5'd24, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000287, 5'd0, 27'h0000006a, 5'd5, 27'h0000033a, 32'h00000400,
  1'd1,  5'd4, 27'h00000113, 5'd3, 27'h000002bd, 5'd19, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000279, 5'd1, 27'h0000007e, 5'd26, 27'h000000fb, 32'h00000400,
  1'd1,  5'd2, 27'h00000248, 5'd10, 27'h00000163, 5'd5, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000006e, 5'd13, 27'h000003aa, 5'd20, 27'h0000007b, 32'h00000400,
  1'd1,  5'd1, 27'h0000035b, 5'd11, 27'h000001b9, 5'd28, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029e, 5'd25, 27'h00000077, 5'd5, 27'h000000ae, 32'h00000400,
  1'd1,  5'd3, 27'h000000d7, 5'd21, 27'h0000018c, 5'd15, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ec, 5'd25, 27'h000001e2, 5'd28, 27'h000003cc, 32'h00000400,
  1'd1,  5'd11, 27'h0000021d, 5'd3, 27'h000003be, 5'd7, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000392, 5'd2, 27'h0000034e, 5'd17, 27'h0000009c, 32'h00000400,
  1'd1,  5'd13, 27'h00000144, 5'd1, 27'h000003d4, 5'd27, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000022b, 5'd14, 27'h000001cd, 5'd6, 27'h000002ee, 32'h00000400,
  1'd1,  5'd14, 27'h0000034d, 5'd11, 27'h00000230, 5'd16, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000156, 5'd12, 27'h000001ce, 5'd29, 27'h0000011d, 32'h00000400,
  1'd1,  5'd14, 27'h0000027e, 5'd24, 27'h0000001b, 5'd7, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000030c, 5'd22, 27'h00000128, 5'd20, 27'h000000c2, 32'h00000400,
  1'd1,  5'd11, 27'h00000285, 5'd24, 27'h000001c0, 5'd30, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019c, 5'd4, 27'h000002bf, 5'd7, 27'h000002df, 32'h00000400,
  1'd1,  5'd21, 27'h00000017, 5'd3, 27'h00000397, 5'd18, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e6, 5'd1, 27'h0000024f, 5'd29, 27'h0000007b, 32'h00000400,
  1'd1,  5'd24, 27'h00000363, 5'd11, 27'h000000f4, 5'd6, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000278, 5'd12, 27'h00000181, 5'd18, 27'h000000ae, 32'h00000400,
  1'd1,  5'd22, 27'h000001e2, 5'd10, 27'h000003f3, 5'd30, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000107, 5'd20, 27'h000003f3, 5'd7, 27'h0000014f, 32'h00000400,
  1'd1,  5'd21, 27'h000001b3, 5'd21, 27'h00000201, 5'd18, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002f3, 5'd23, 27'h0000001a, 5'd30, 27'h00000259, 32'h00000400,
  1'd1,  5'd2, 27'h0000031d, 5'd7, 27'h00000065, 5'd1, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029a, 5'd10, 27'h00000080, 5'd11, 27'h000001a3, 32'h00000400,
  1'd1,  5'd4, 27'h0000010b, 5'd7, 27'h00000167, 5'd24, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000032, 5'd16, 27'h000001bf, 5'd3, 27'h00000380, 32'h00000400,
  1'd1,  5'd3, 27'h000002d3, 5'd18, 27'h00000259, 5'd14, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000182, 5'd20, 27'h00000149, 5'd25, 27'h000002e0, 32'h00000400,
  1'd1,  5'd2, 27'h0000015f, 5'd26, 27'h0000017d, 5'd1, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000030b, 5'd28, 27'h00000305, 5'd11, 27'h000002e2, 32'h00000400,
  1'd1,  5'd0, 27'h000000c4, 5'd27, 27'h00000241, 5'd20, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000167, 5'd9, 27'h00000221, 5'd4, 27'h0000003f, 32'h00000400,
  1'd1,  5'd13, 27'h00000100, 5'd10, 27'h00000086, 5'd14, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000039f, 5'd8, 27'h000000ce, 5'd24, 27'h0000031c, 32'h00000400,
  1'd1,  5'd11, 27'h000001c7, 5'd18, 27'h000000db, 5'd0, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000037b, 5'd16, 27'h00000332, 5'd14, 27'h000000ed, 32'h00000400,
  1'd1,  5'd12, 27'h000003c3, 5'd18, 27'h000000f2, 5'd25, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001dc, 5'd28, 27'h0000036d, 5'd0, 27'h0000031a, 32'h00000400,
  1'd1,  5'd12, 27'h00000076, 5'd27, 27'h00000162, 5'd13, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000150, 5'd27, 27'h0000032c, 5'd22, 27'h0000006a, 32'h00000400,
  1'd1,  5'd23, 27'h000003e5, 5'd5, 27'h0000035d, 5'd4, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d4, 5'd5, 27'h0000027c, 5'd10, 27'h0000038e, 32'h00000400,
  1'd1,  5'd25, 27'h00000204, 5'd7, 27'h00000056, 5'd22, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000391, 5'd19, 27'h0000039d, 5'd2, 27'h00000356, 32'h00000400,
  1'd1,  5'd23, 27'h00000020, 5'd19, 27'h0000014c, 5'd12, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000019f, 5'd15, 27'h00000346, 5'd24, 27'h000002a9, 32'h00000400,
  1'd1,  5'd21, 27'h00000121, 5'd26, 27'h000001c8, 5'd0, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000011, 5'd30, 27'h00000036, 5'd14, 27'h00000279, 32'h00000400,
  1'd1,  5'd21, 27'h00000259, 5'd30, 27'h00000284, 5'd23, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002b8, 5'd5, 27'h000002cc, 5'd7, 27'h000000c4, 32'h00000400,
  1'd1,  5'd5, 27'h0000000e, 5'd7, 27'h00000159, 5'd19, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000393, 5'd7, 27'h00000275, 5'd28, 27'h0000000c, 32'h00000400,
  1'd1,  5'd4, 27'h000000c9, 5'd20, 27'h000000b1, 5'd7, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000033, 5'd19, 27'h000000f9, 5'd18, 27'h000001a8, 32'h00000400,
  1'd1,  5'd0, 27'h000001aa, 5'd17, 27'h000002e4, 5'd28, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000277, 5'd28, 27'h00000266, 5'd10, 27'h000000b4, 32'h00000400,
  1'd1,  5'd3, 27'h000000c4, 5'd30, 27'h000002cc, 5'd16, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000190, 5'd30, 27'h00000058, 5'd29, 27'h0000026f, 32'h00000400,
  1'd1,  5'd14, 27'h00000227, 5'd9, 27'h000003fa, 5'd9, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000016f, 5'd5, 27'h0000017d, 5'd18, 27'h0000019c, 32'h00000400,
  1'd1,  5'd15, 27'h00000014, 5'd9, 27'h00000365, 5'd30, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000171, 5'd18, 27'h00000177, 5'd10, 27'h00000064, 32'h00000400,
  1'd1,  5'd13, 27'h000001d0, 5'd20, 27'h0000000d, 5'd18, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f6, 5'd19, 27'h00000215, 5'd27, 27'h00000065, 32'h00000400,
  1'd1,  5'd11, 27'h000000de, 5'd26, 27'h000001f1, 5'd10, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d0, 5'd30, 27'h00000036, 5'd18, 27'h0000029a, 32'h00000400,
  1'd1,  5'd14, 27'h000000ed, 5'd30, 27'h00000079, 5'd27, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b7, 5'd5, 27'h00000330, 5'd8, 27'h000003fb, 32'h00000400,
  1'd1,  5'd25, 27'h000000f6, 5'd6, 27'h00000341, 5'd18, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a4, 5'd10, 27'h000000e2, 5'd29, 27'h000003d3, 32'h00000400,
  1'd1,  5'd24, 27'h00000331, 5'd19, 27'h000001fd, 5'd5, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000020b, 5'd17, 27'h00000343, 5'd15, 27'h0000033a, 32'h00000400,
  1'd1,  5'd22, 27'h0000032e, 5'd15, 27'h0000038b, 5'd29, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b8, 5'd26, 27'h00000396, 5'd7, 27'h000002f3, 32'h00000400,
  1'd1,  5'd23, 27'h0000013f, 5'd30, 27'h000003cd, 5'd15, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000037, 5'd27, 27'h000002ef, 5'd27, 27'h00000052, 32'h00000400,
  1'd1,  5'd9, 27'h00000293, 5'd2, 27'h00000090, 5'd8, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000023a, 5'd4, 27'h00000131, 5'd16, 27'h0000014d, 32'h00000400,
  1'd1,  5'd8, 27'h000000e9, 5'd0, 27'h000001e0, 5'd30, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000e7, 5'd14, 27'h00000041, 5'd2, 27'h00000040, 32'h00000400,
  1'd1,  5'd6, 27'h000001e1, 5'd13, 27'h000001b8, 5'd13, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000262, 5'd12, 27'h00000325, 5'd20, 27'h000003d8, 32'h00000400,
  1'd1,  5'd9, 27'h0000000e, 5'd24, 27'h00000366, 5'd0, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000343, 5'd25, 27'h00000009, 5'd15, 27'h00000065, 32'h00000400,
  1'd1,  5'd5, 27'h000003ef, 5'd23, 27'h00000121, 5'd24, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d3, 5'd1, 27'h000003f3, 5'd7, 27'h000000f6, 32'h00000400,
  1'd1,  5'd16, 27'h0000033d, 5'd0, 27'h00000281, 5'd17, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ce, 5'd0, 27'h0000021e, 5'd25, 27'h000003a4, 32'h00000400,
  1'd1,  5'd17, 27'h00000199, 5'd12, 27'h00000259, 5'd2, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000246, 5'd10, 27'h000002c8, 5'd13, 27'h0000008e, 32'h00000400,
  1'd1,  5'd19, 27'h000002f2, 5'd11, 27'h000002e8, 5'd24, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ae, 5'd22, 27'h00000373, 5'd1, 27'h00000277, 32'h00000400,
  1'd1,  5'd16, 27'h0000003c, 5'd24, 27'h0000022a, 5'd14, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d4, 5'd21, 27'h00000315, 5'd20, 27'h000003f1, 32'h00000400,
  1'd1,  5'd29, 27'h0000036e, 5'd3, 27'h000003a8, 5'd1, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000250, 5'd3, 27'h000000d7, 5'd11, 27'h00000210, 32'h00000400,
  1'd1,  5'd30, 27'h00000160, 5'd2, 27'h00000165, 5'd21, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000271, 5'd13, 27'h00000075, 5'd1, 27'h0000025a, 32'h00000400,
  1'd1,  5'd27, 27'h0000021c, 5'd11, 27'h00000146, 5'd15, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000fc, 5'd14, 27'h00000078, 5'd21, 27'h000002d9, 32'h00000400,
  1'd1,  5'd29, 27'h000000d3, 5'd22, 27'h00000164, 5'd2, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ee, 5'd20, 27'h00000386, 5'd14, 27'h0000014e, 32'h00000400,
  1'd1,  5'd28, 27'h00000109, 5'd22, 27'h0000003a, 5'd22, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000351, 5'd1, 27'h000001b3, 5'd0, 27'h000002cb, 32'h00000400,
  1'd1,  5'd10, 27'h0000002e, 5'd5, 27'h0000004a, 5'd14, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000008e, 5'd4, 27'h0000012a, 5'd25, 27'h00000077, 32'h00000400,
  1'd1,  5'd9, 27'h00000312, 5'd12, 27'h000000ed, 5'd9, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ac, 5'd12, 27'h000002ad, 5'd19, 27'h00000233, 32'h00000400,
  1'd1,  5'd9, 27'h0000030b, 5'd15, 27'h000001a5, 5'd27, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002af, 5'd21, 27'h00000001, 5'd7, 27'h000000e8, 32'h00000400,
  1'd1,  5'd8, 27'h00000169, 5'd24, 27'h000003d0, 5'd16, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001f0, 5'd22, 27'h000001b3, 5'd26, 27'h0000022f, 32'h00000400,
  1'd1,  5'd18, 27'h00000103, 5'd1, 27'h000002b0, 5'd3, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000243, 5'd1, 27'h0000022c, 5'd10, 27'h000001da, 32'h00000400,
  1'd1,  5'd18, 27'h00000366, 5'd0, 27'h000000f0, 5'd23, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000352, 5'd13, 27'h00000003, 5'd8, 27'h0000033b, 32'h00000400,
  1'd1,  5'd18, 27'h000001d6, 5'd10, 27'h00000230, 5'd16, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000287, 5'd11, 27'h000000c5, 5'd26, 27'h00000047, 32'h00000400,
  1'd1,  5'd20, 27'h000000cf, 5'd23, 27'h000000c0, 5'd5, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003f6, 5'd23, 27'h000000c8, 5'd17, 27'h000000b9, 32'h00000400,
  1'd1,  5'd20, 27'h00000029, 5'd22, 27'h00000012, 5'd28, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003fa, 5'd1, 27'h00000293, 5'd6, 27'h00000276, 32'h00000400,
  1'd1,  5'd29, 27'h000001bd, 5'd3, 27'h0000029e, 5'd20, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001b8, 5'd2, 27'h00000228, 5'd28, 27'h000003f2, 32'h00000400,
  1'd1,  5'd29, 27'h000003b4, 5'd15, 27'h00000013, 5'd5, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e6, 5'd14, 27'h000002f2, 5'd16, 27'h000003f7, 32'h00000400,
  1'd1,  5'd26, 27'h0000034c, 5'd12, 27'h00000088, 5'd27, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000188, 5'd25, 27'h00000149, 5'd8, 27'h00000329, 32'h00000400,
  1'd1,  5'd29, 27'h000000c5, 5'd25, 27'h0000010e, 5'd17, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000170, 5'd25, 27'h000002e4, 5'd26, 27'h000001da, 32'h00000400,
  1'd1,  5'd5, 27'h000001c3, 5'd7, 27'h00000037, 5'd3, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000019a, 5'd9, 27'h000003e8, 5'd12, 27'h00000082, 32'h00000400,
  1'd1,  5'd8, 27'h000000e9, 5'd6, 27'h00000356, 5'd24, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000014c, 5'd16, 27'h00000148, 5'd0, 27'h00000038, 32'h00000400,
  1'd1,  5'd9, 27'h00000375, 5'd16, 27'h0000008a, 5'd12, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003c2, 5'd17, 27'h00000165, 5'd23, 27'h0000014f, 32'h00000400,
  1'd1,  5'd10, 27'h000000b6, 5'd26, 27'h0000020b, 5'd3, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000016c, 5'd29, 27'h00000365, 5'd10, 27'h000003a3, 32'h00000400,
  1'd1,  5'd7, 27'h000003fe, 5'd30, 27'h00000286, 5'd22, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000072, 5'd8, 27'h00000259, 5'd1, 27'h000000e0, 32'h00000400,
  1'd1,  5'd19, 27'h0000029d, 5'd5, 27'h0000035a, 5'd15, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000340, 5'd5, 27'h000003c8, 5'd20, 27'h00000353, 32'h00000400,
  1'd1,  5'd17, 27'h00000135, 5'd18, 27'h000002af, 5'd3, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000333, 5'd20, 27'h00000010, 5'd13, 27'h00000245, 32'h00000400,
  1'd1,  5'd19, 27'h00000342, 5'd17, 27'h000001da, 5'd22, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000359, 5'd26, 27'h00000369, 5'd4, 27'h000001c3, 32'h00000400,
  1'd1,  5'd19, 27'h000001ea, 5'd28, 27'h00000100, 5'd10, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000217, 5'd29, 27'h00000231, 5'd22, 27'h0000021c, 32'h00000400,
  1'd1,  5'd27, 27'h00000192, 5'd9, 27'h00000247, 5'd0, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000057, 5'd6, 27'h00000235, 5'd11, 27'h000003cb, 32'h00000400,
  1'd1,  5'd28, 27'h000003f5, 5'd7, 27'h00000219, 5'd25, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003d8, 5'd17, 27'h0000001e, 5'd0, 27'h000001da, 32'h00000400,
  1'd1,  5'd30, 27'h00000006, 5'd19, 27'h000003ea, 5'd10, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003cf, 5'd18, 27'h00000271, 5'd24, 27'h0000016f, 32'h00000400,
  1'd1,  5'd27, 27'h0000000b, 5'd26, 27'h00000371, 5'd2, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000039f, 5'd29, 27'h000001ea, 5'd13, 27'h00000349, 32'h00000400,
  1'd1,  5'd30, 27'h00000252, 5'd30, 27'h000003a5, 5'd22, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000012a, 5'd8, 27'h00000142, 5'd8, 27'h00000375, 32'h00000400,
  1'd1,  5'd8, 27'h000000c6, 5'd6, 27'h000000ff, 5'd20, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000044, 5'd7, 27'h00000113, 5'd28, 27'h000003d1, 32'h00000400,
  1'd1,  5'd8, 27'h00000101, 5'd16, 27'h000002e8, 5'd9, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000310, 5'd16, 27'h000001e5, 5'd17, 27'h00000160, 32'h00000400,
  1'd1,  5'd8, 27'h000000d8, 5'd16, 27'h000003af, 5'd30, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032c, 5'd29, 27'h0000007e, 5'd6, 27'h00000056, 32'h00000400,
  1'd1,  5'd9, 27'h00000400, 5'd30, 27'h0000037c, 5'd19, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e7, 5'd27, 27'h00000301, 5'd28, 27'h000003f5, 32'h00000400,
  1'd1,  5'd18, 27'h00000371, 5'd8, 27'h000002d0, 5'd9, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002d6, 5'd7, 27'h000000e1, 5'd19, 27'h000002f7, 32'h00000400,
  1'd1,  5'd18, 27'h0000028e, 5'd8, 27'h00000075, 5'd30, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ea, 5'd16, 27'h0000003a, 5'd6, 27'h000001fc, 32'h00000400,
  1'd1,  5'd15, 27'h000003b2, 5'd20, 27'h00000127, 5'd17, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000030f, 5'd16, 27'h00000346, 5'd26, 27'h000002fd, 32'h00000400,
  1'd1,  5'd17, 27'h000000ed, 5'd26, 27'h000000a3, 5'd5, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000019e, 5'd26, 27'h0000024f, 5'd19, 27'h00000127, 32'h00000400,
  1'd1,  5'd16, 27'h00000001, 5'd25, 27'h000003b2, 5'd29, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000038, 5'd5, 27'h00000289, 5'd9, 27'h00000190, 32'h00000400,
  1'd1,  5'd29, 27'h000002f8, 5'd6, 27'h000000ad, 5'd16, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000e0, 5'd6, 27'h000003bc, 5'd26, 27'h00000326, 32'h00000400,
  1'd1,  5'd26, 27'h000000ed, 5'd20, 27'h0000026f, 5'd5, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000180, 5'd17, 27'h0000024f, 5'd15, 27'h000003aa, 32'h00000400,
  1'd1,  5'd30, 27'h0000039f, 5'd17, 27'h0000028f, 5'd29, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000117, 5'd29, 27'h0000018a, 5'd8, 27'h000001f3, 32'h00000400,
  1'd1,  5'd30, 27'h00000123, 5'd26, 27'h00000018, 5'd20, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003cf, 5'd27, 27'h0000029e, 5'd26, 27'h000003f6, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000002ba, 5'd3, 27'h0000005a, 5'd3, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a2, 5'd5, 27'h00000083, 5'd15, 27'h00000192, 32'h00000400,
  1'd1,  5'd2, 27'h000002d4, 5'd4, 27'h000002c1, 5'd23, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000181, 5'd11, 27'h0000036d, 5'd2, 27'h00000134, 32'h00000400,
  1'd1,  5'd3, 27'h000002a7, 5'd11, 27'h00000223, 5'd14, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000133, 5'd15, 27'h0000019d, 5'd25, 27'h000000e9, 32'h00000400,
  1'd1,  5'd2, 27'h00000275, 5'd22, 27'h000003ad, 5'd2, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002ad, 5'd24, 27'h00000381, 5'd11, 27'h0000004f, 32'h00000400,
  1'd1,  5'd4, 27'h000002e0, 5'd22, 27'h00000280, 5'd22, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000034a, 5'd2, 27'h00000206, 5'd3, 27'h000001e5, 32'h00000400,
  1'd1,  5'd12, 27'h0000037f, 5'd2, 27'h00000343, 5'd13, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000283, 5'd4, 27'h0000008d, 5'd21, 27'h00000141, 32'h00000400,
  1'd1,  5'd12, 27'h000002f7, 5'd15, 27'h000001bf, 5'd3, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000018d, 5'd11, 27'h0000010a, 5'd13, 27'h00000038, 32'h00000400,
  1'd1,  5'd11, 27'h00000030, 5'd10, 27'h000001fd, 5'd21, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003af, 5'd21, 27'h00000226, 5'd2, 27'h000003df, 32'h00000400,
  1'd1,  5'd12, 27'h00000087, 5'd24, 27'h00000232, 5'd11, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000085, 5'd24, 27'h000001c4, 5'd20, 27'h000002d6, 32'h00000400,
  1'd1,  5'd25, 27'h00000339, 5'd3, 27'h000001c1, 5'd2, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000273, 5'd4, 27'h000002d5, 5'd10, 27'h000003e2, 32'h00000400,
  1'd1,  5'd24, 27'h000002ce, 5'd4, 27'h000001c7, 5'd22, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002cf, 5'd11, 27'h00000305, 5'd1, 27'h0000003d, 32'h00000400,
  1'd1,  5'd25, 27'h0000002a, 5'd14, 27'h0000005d, 5'd15, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000035d, 5'd15, 27'h000000a8, 5'd23, 27'h0000014a, 32'h00000400,
  1'd1,  5'd22, 27'h000002f8, 5'd25, 27'h0000015a, 5'd3, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000171, 5'd22, 27'h00000047, 5'd10, 27'h000003d6, 32'h00000400,
  1'd1,  5'd25, 27'h0000007a, 5'd23, 27'h000000aa, 5'd25, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000004a, 5'd4, 27'h00000178, 5'd5, 27'h0000013e, 32'h00000400,
  1'd1,  5'd4, 27'h000002e6, 5'd4, 27'h00000011, 5'd18, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000035, 5'd1, 27'h000003fb, 5'd28, 27'h00000252, 32'h00000400,
  1'd1,  5'd3, 27'h00000292, 5'd11, 27'h000003c1, 5'd9, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000003c, 5'd12, 27'h000002a5, 5'd15, 27'h00000241, 32'h00000400,
  1'd1,  5'd4, 27'h000003d8, 5'd11, 27'h0000016d, 5'd30, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000214, 5'd22, 27'h000002df, 5'd7, 27'h000003b4, 32'h00000400,
  1'd1,  5'd0, 27'h00000173, 5'd25, 27'h00000350, 5'd18, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000265, 5'd22, 27'h00000079, 5'd26, 27'h000003b9, 32'h00000400,
  1'd1,  5'd13, 27'h000000c5, 5'd3, 27'h00000208, 5'd9, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000a2, 5'd1, 27'h00000027, 5'd16, 27'h0000013a, 32'h00000400,
  1'd1,  5'd11, 27'h000002cd, 5'd0, 27'h000002fe, 5'd28, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000216, 5'd13, 27'h00000351, 5'd10, 27'h000000a7, 32'h00000400,
  1'd1,  5'd12, 27'h0000011d, 5'd13, 27'h00000123, 5'd17, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003be, 5'd13, 27'h000001aa, 5'd27, 27'h00000375, 32'h00000400,
  1'd1,  5'd13, 27'h00000377, 5'd20, 27'h000003aa, 5'd7, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000307, 5'd21, 27'h000003f8, 5'd15, 27'h0000021c, 32'h00000400,
  1'd1,  5'd11, 27'h000003a5, 5'd25, 27'h0000000e, 5'd29, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000034e, 5'd3, 27'h000002fe, 5'd7, 27'h000002f8, 32'h00000400,
  1'd1,  5'd23, 27'h00000168, 5'd0, 27'h0000035a, 5'd20, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002c1, 5'd2, 27'h00000237, 5'd27, 27'h000000cf, 32'h00000400,
  1'd1,  5'd24, 27'h000002bb, 5'd13, 27'h00000100, 5'd9, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000031c, 5'd12, 27'h00000176, 5'd19, 27'h00000180, 32'h00000400,
  1'd1,  5'd21, 27'h00000231, 5'd12, 27'h00000376, 5'd25, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000015e, 5'd24, 27'h00000210, 5'd8, 27'h00000105, 32'h00000400,
  1'd1,  5'd23, 27'h000002f2, 5'd23, 27'h000002ad, 5'd16, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a0, 5'd24, 27'h000001da, 5'd26, 27'h00000128, 32'h00000400,
  1'd1,  5'd3, 27'h00000328, 5'd7, 27'h0000016f, 5'd2, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000000a, 5'd9, 27'h00000173, 5'd14, 27'h0000036c, 32'h00000400,
  1'd1,  5'd3, 27'h000002e3, 5'd6, 27'h000001d8, 5'd24, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f1, 5'd19, 27'h000002da, 5'd4, 27'h000003f5, 32'h00000400,
  1'd1,  5'd1, 27'h00000125, 5'd20, 27'h0000010e, 5'd11, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e5, 5'd20, 27'h00000284, 5'd25, 27'h00000037, 32'h00000400,
  1'd1,  5'd4, 27'h00000229, 5'd30, 27'h00000145, 5'd2, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001dd, 5'd29, 27'h0000035b, 5'd14, 27'h000000aa, 32'h00000400,
  1'd1,  5'd4, 27'h00000274, 5'd27, 27'h00000350, 5'd25, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000016c, 5'd9, 27'h00000052, 5'd5, 27'h00000098, 32'h00000400,
  1'd1,  5'd15, 27'h000001ff, 5'd9, 27'h000000b9, 5'd10, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000034e, 5'd9, 27'h00000147, 5'd22, 27'h00000045, 32'h00000400,
  1'd1,  5'd15, 27'h0000010e, 5'd16, 27'h0000023a, 5'd0, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003e9, 5'd17, 27'h00000322, 5'd12, 27'h0000008a, 32'h00000400,
  1'd1,  5'd14, 27'h0000000b, 5'd19, 27'h0000015c, 5'd25, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002c2, 5'd29, 27'h00000006, 5'd1, 27'h000001b7, 32'h00000400,
  1'd1,  5'd14, 27'h00000334, 5'd28, 27'h000001a3, 5'd10, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e2, 5'd27, 27'h0000037b, 5'd21, 27'h000000e7, 32'h00000400,
  1'd1,  5'd24, 27'h00000318, 5'd9, 27'h000002c5, 5'd4, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003c3, 5'd9, 27'h000003ad, 5'd15, 27'h000000e6, 32'h00000400,
  1'd1,  5'd23, 27'h00000261, 5'd7, 27'h00000389, 5'd23, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000fa, 5'd18, 27'h000001ae, 5'd2, 27'h0000018c, 32'h00000400,
  1'd1,  5'd25, 27'h0000009f, 5'd15, 27'h0000021f, 5'd10, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000016b, 5'd19, 27'h00000026, 5'd22, 27'h00000124, 32'h00000400,
  1'd1,  5'd24, 27'h00000339, 5'd29, 27'h00000289, 5'd5, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b7, 5'd29, 27'h0000026f, 5'd14, 27'h00000050, 32'h00000400,
  1'd1,  5'd24, 27'h00000140, 5'd26, 27'h00000099, 5'd25, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000bd, 5'd8, 27'h00000191, 5'd7, 27'h00000113, 32'h00000400,
  1'd1,  5'd0, 27'h00000023, 5'd9, 27'h000003bc, 5'd16, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000209, 5'd8, 27'h00000298, 5'd29, 27'h000003ca, 32'h00000400,
  1'd1,  5'd3, 27'h00000349, 5'd16, 27'h00000279, 5'd7, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000400, 5'd16, 27'h00000397, 5'd19, 27'h000003d4, 32'h00000400,
  1'd1,  5'd3, 27'h000002c5, 5'd18, 27'h00000104, 5'd26, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d0, 5'd26, 27'h0000031a, 5'd5, 27'h0000018c, 32'h00000400,
  1'd1,  5'd4, 27'h00000258, 5'd27, 27'h00000097, 5'd19, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b3, 5'd27, 27'h0000033a, 5'd26, 27'h0000021b, 32'h00000400,
  1'd1,  5'd10, 27'h0000039b, 5'd5, 27'h00000245, 5'd6, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001c6, 5'd5, 27'h000002aa, 5'd17, 27'h000002da, 32'h00000400,
  1'd1,  5'd12, 27'h000002da, 5'd8, 27'h00000301, 5'd26, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000aa, 5'd16, 27'h0000023d, 5'd7, 27'h0000029e, 32'h00000400,
  1'd1,  5'd15, 27'h0000002d, 5'd15, 27'h00000322, 5'd19, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002a0, 5'd18, 27'h00000042, 5'd28, 27'h0000016b, 32'h00000400,
  1'd1,  5'd10, 27'h0000032f, 5'd28, 27'h000000f6, 5'd5, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000295, 5'd29, 27'h00000239, 5'd20, 27'h00000112, 32'h00000400,
  1'd1,  5'd13, 27'h00000188, 5'd28, 27'h0000014a, 5'd26, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000051, 5'd6, 27'h0000033f, 5'd6, 27'h0000009b, 32'h00000400,
  1'd1,  5'd21, 27'h000002fc, 5'd5, 27'h00000387, 5'd15, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000244, 5'd6, 27'h000003c4, 5'd28, 27'h00000070, 32'h00000400,
  1'd1,  5'd23, 27'h00000380, 5'd20, 27'h000002a1, 5'd6, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000169, 5'd19, 27'h000002ca, 5'd18, 27'h00000312, 32'h00000400,
  1'd1,  5'd23, 27'h000003b5, 5'd16, 27'h000001e2, 5'd29, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000007f, 5'd26, 27'h000000ac, 5'd9, 27'h00000129, 32'h00000400,
  1'd1,  5'd22, 27'h00000033, 5'd26, 27'h00000132, 5'd17, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000399, 5'd30, 27'h000001da, 5'd30, 27'h000003b3, 32'h00000400,
  1'd1,  5'd9, 27'h00000088, 5'd4, 27'h000003b0, 5'd6, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000018d, 5'd1, 27'h00000242, 5'd19, 27'h00000159, 32'h00000400,
  1'd1,  5'd6, 27'h0000019d, 5'd1, 27'h000003f8, 5'd28, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000017e, 5'd14, 27'h00000325, 5'd4, 27'h000000e6, 32'h00000400,
  1'd1,  5'd5, 27'h000001c3, 5'd10, 27'h000003b3, 5'd13, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000fb, 5'd11, 27'h00000245, 5'd22, 27'h0000035d, 32'h00000400,
  1'd1,  5'd9, 27'h000001c9, 5'd24, 27'h00000107, 5'd3, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ef, 5'd23, 27'h0000002e, 5'd13, 27'h000002a8, 32'h00000400,
  1'd1,  5'd9, 27'h000000ec, 5'd25, 27'h000000dc, 5'd22, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002d1, 5'd2, 27'h00000266, 5'd6, 27'h0000001e, 32'h00000400,
  1'd1,  5'd15, 27'h000003d5, 5'd3, 27'h00000328, 5'd19, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000217, 5'd0, 27'h00000007, 5'd29, 27'h00000087, 32'h00000400,
  1'd1,  5'd20, 27'h000001c1, 5'd10, 27'h00000289, 5'd0, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000049, 5'd10, 27'h0000021a, 5'd15, 27'h0000009f, 32'h00000400,
  1'd1,  5'd20, 27'h000000ce, 5'd11, 27'h000000cc, 5'd25, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000310, 5'd25, 27'h00000074, 5'd0, 27'h000000e9, 32'h00000400,
  1'd1,  5'd16, 27'h000000f6, 5'd24, 27'h000003b4, 5'd11, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000299, 5'd23, 27'h000002be, 5'd21, 27'h0000025b, 32'h00000400,
  1'd1,  5'd29, 27'h000000f6, 5'd5, 27'h00000057, 5'd3, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000004a, 5'd4, 27'h000000af, 5'd14, 27'h000001f4, 32'h00000400,
  1'd1,  5'd28, 27'h0000012d, 5'd2, 27'h000002b7, 5'd23, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002bf, 5'd15, 27'h0000006a, 5'd2, 27'h00000297, 32'h00000400,
  1'd1,  5'd28, 27'h0000037d, 5'd11, 27'h00000198, 5'd10, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000198, 5'd10, 27'h00000399, 5'd20, 27'h000003fd, 32'h00000400,
  1'd1,  5'd29, 27'h0000034b, 5'd24, 27'h000001f9, 5'd2, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000018f, 5'd25, 27'h0000009c, 5'd13, 27'h00000093, 32'h00000400,
  1'd1,  5'd27, 27'h00000040, 5'd21, 27'h00000026, 5'd25, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001cf, 5'd2, 27'h00000280, 5'd3, 27'h000001bd, 32'h00000400,
  1'd1,  5'd5, 27'h00000247, 5'd2, 27'h000000cc, 5'd13, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c4, 5'd1, 27'h000002ef, 5'd21, 27'h000000a8, 32'h00000400,
  1'd1,  5'd7, 27'h000002a2, 5'd13, 27'h00000394, 5'd8, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000013b, 5'd11, 27'h00000342, 5'd20, 27'h000001a7, 32'h00000400,
  1'd1,  5'd6, 27'h00000097, 5'd10, 27'h00000227, 5'd28, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000056, 5'd22, 27'h000003eb, 5'd8, 27'h000003e4, 32'h00000400,
  1'd1,  5'd6, 27'h0000012a, 5'd25, 27'h0000016e, 5'd20, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000024c, 5'd24, 27'h00000277, 5'd26, 27'h0000039f, 32'h00000400,
  1'd1,  5'd18, 27'h00000098, 5'd0, 27'h0000029e, 5'd5, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c2, 5'd0, 27'h00000008, 5'd12, 27'h0000011a, 32'h00000400,
  1'd1,  5'd16, 27'h000003c2, 5'd1, 27'h00000228, 5'd24, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025e, 5'd12, 27'h00000241, 5'd8, 27'h0000029e, 32'h00000400,
  1'd1,  5'd15, 27'h000003ed, 5'd15, 27'h000001d9, 5'd17, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000015d, 5'd10, 27'h00000271, 5'd28, 27'h000002ab, 32'h00000400,
  1'd1,  5'd18, 27'h00000354, 5'd22, 27'h00000194, 5'd5, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000039d, 5'd24, 27'h000000f5, 5'd20, 27'h00000178, 32'h00000400,
  1'd1,  5'd18, 27'h000000d5, 5'd23, 27'h0000016c, 5'd29, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b5, 5'd3, 27'h000002fe, 5'd7, 27'h0000005a, 32'h00000400,
  1'd1,  5'd26, 27'h00000309, 5'd4, 27'h000001f8, 5'd19, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000152, 5'd5, 27'h00000097, 5'd27, 27'h000002e9, 32'h00000400,
  1'd1,  5'd26, 27'h0000003a, 5'd14, 27'h000002f2, 5'd9, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d6, 5'd12, 27'h0000006d, 5'd20, 27'h00000034, 32'h00000400,
  1'd1,  5'd27, 27'h0000007c, 5'd14, 27'h00000272, 5'd26, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000eb, 5'd25, 27'h000000ee, 5'd6, 27'h00000202, 32'h00000400,
  1'd1,  5'd29, 27'h000003d9, 5'd24, 27'h00000378, 5'd16, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000221, 5'd20, 27'h00000387, 5'd30, 27'h00000314, 32'h00000400,
  1'd1,  5'd6, 27'h0000020a, 5'd7, 27'h00000184, 5'd1, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d7, 5'd7, 27'h0000009a, 5'd14, 27'h0000010c, 32'h00000400,
  1'd1,  5'd5, 27'h000001a6, 5'd5, 27'h0000028c, 5'd25, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e3, 5'd19, 27'h000001ce, 5'd3, 27'h000001c6, 32'h00000400,
  1'd1,  5'd7, 27'h0000018c, 5'd19, 27'h00000176, 5'd11, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000033d, 5'd17, 27'h0000026c, 5'd21, 27'h000003bc, 32'h00000400,
  1'd1,  5'd8, 27'h000003f7, 5'd28, 27'h000002f7, 5'd0, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b3, 5'd28, 27'h00000271, 5'd11, 27'h0000025b, 32'h00000400,
  1'd1,  5'd7, 27'h000001f3, 5'd28, 27'h000001cc, 5'd22, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000157, 5'd7, 27'h0000005a, 5'd1, 27'h0000013b, 32'h00000400,
  1'd1,  5'd18, 27'h00000337, 5'd6, 27'h00000183, 5'd15, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001a1, 5'd8, 27'h00000177, 5'd22, 27'h000003a0, 32'h00000400,
  1'd1,  5'd17, 27'h0000011d, 5'd16, 27'h000000bb, 5'd0, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e3, 5'd20, 27'h000000f1, 5'd10, 27'h00000224, 32'h00000400,
  1'd1,  5'd16, 27'h0000009f, 5'd19, 27'h0000011d, 5'd22, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003ec, 5'd28, 27'h00000043, 5'd2, 27'h0000007e, 32'h00000400,
  1'd1,  5'd17, 27'h00000124, 5'd29, 27'h000002dd, 5'd11, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001fb, 5'd28, 27'h000002a5, 5'd23, 27'h000000ff, 32'h00000400,
  1'd1,  5'd27, 27'h00000369, 5'd6, 27'h00000017, 5'd5, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000014f, 5'd6, 27'h00000274, 5'd13, 27'h000000cd, 32'h00000400,
  1'd1,  5'd30, 27'h000001fa, 5'd9, 27'h00000164, 5'd25, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000072, 5'd19, 27'h000001fc, 5'd0, 27'h000001fc, 32'h00000400,
  1'd1,  5'd27, 27'h0000015c, 5'd16, 27'h000001e9, 5'd12, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000020a, 5'd18, 27'h000001b1, 5'd25, 27'h0000028f, 32'h00000400,
  1'd1,  5'd27, 27'h00000287, 5'd30, 27'h00000242, 5'd1, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000281, 5'd26, 27'h00000384, 5'd11, 27'h00000366, 32'h00000400,
  1'd1,  5'd29, 27'h00000215, 5'd28, 27'h0000022e, 5'd22, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000031c, 5'd5, 27'h0000012e, 5'd6, 27'h00000055, 32'h00000400,
  1'd1,  5'd8, 27'h00000089, 5'd5, 27'h000002fd, 5'd20, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000013b, 5'd8, 27'h000002d2, 5'd28, 27'h000000e2, 32'h00000400,
  1'd1,  5'd5, 27'h000003bd, 5'd16, 27'h000003c4, 5'd8, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000093, 5'd17, 27'h000000aa, 5'd19, 27'h000000f4, 32'h00000400,
  1'd1,  5'd9, 27'h00000080, 5'd18, 27'h00000173, 5'd27, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001f1, 5'd29, 27'h000000e8, 5'd6, 27'h0000026a, 32'h00000400,
  1'd1,  5'd6, 27'h00000251, 5'd28, 27'h0000018c, 5'd15, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cf, 5'd30, 27'h000000e9, 5'd27, 27'h00000306, 32'h00000400,
  1'd1,  5'd16, 27'h00000043, 5'd9, 27'h0000034c, 5'd9, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000ac, 5'd8, 27'h0000038f, 5'd18, 27'h00000324, 32'h00000400,
  1'd1,  5'd19, 27'h00000338, 5'd6, 27'h00000037, 5'd30, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a3, 5'd17, 27'h000001f7, 5'd7, 27'h000000ea, 32'h00000400,
  1'd1,  5'd16, 27'h0000017e, 5'd15, 27'h00000250, 5'd19, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a5, 5'd18, 27'h00000050, 5'd28, 27'h000003b0, 32'h00000400,
  1'd1,  5'd20, 27'h00000067, 5'd27, 27'h000000af, 5'd6, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b1, 5'd27, 27'h00000120, 5'd17, 27'h00000121, 32'h00000400,
  1'd1,  5'd18, 27'h000003fb, 5'd26, 27'h00000043, 5'd26, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000346, 5'd5, 27'h0000033c, 5'd5, 27'h00000309, 32'h00000400,
  1'd1,  5'd29, 27'h00000200, 5'd8, 27'h0000016a, 5'd18, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000391, 5'd8, 27'h000001d9, 5'd28, 27'h00000041, 32'h00000400,
  1'd1,  5'd29, 27'h0000028f, 5'd16, 27'h0000021e, 5'd6, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000117, 5'd17, 27'h000003de, 5'd15, 27'h0000038c, 32'h00000400,
  1'd1,  5'd29, 27'h00000089, 5'd17, 27'h000000dc, 5'd27, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000356, 5'd28, 27'h0000010a, 5'd6, 27'h000002a6, 32'h00000400,
  1'd1,  5'd26, 27'h00000066, 5'd30, 27'h0000014b, 5'd18, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000014, 5'd30, 27'h00000283, 5'd29, 27'h00000272, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000000de, 5'd0, 27'h000000fc, 5'd1, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000015b, 5'd2, 27'h000001dc, 5'd12, 27'h00000337, 32'h00000400,
  1'd1,  5'd4, 27'h000003c5, 5'd4, 27'h00000275, 5'd24, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ad, 5'd11, 27'h00000113, 5'd2, 27'h0000015a, 32'h00000400,
  1'd1,  5'd1, 27'h000001f0, 5'd11, 27'h000001d7, 5'd11, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000ca, 5'd10, 27'h00000170, 5'd21, 27'h000003a6, 32'h00000400,
  1'd1,  5'd3, 27'h0000020b, 5'd25, 27'h00000121, 5'd0, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000029d, 5'd25, 27'h000002f9, 5'd10, 27'h00000168, 32'h00000400,
  1'd1,  5'd4, 27'h0000030a, 5'd22, 27'h0000034d, 5'd21, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000254, 5'd3, 27'h000002c0, 5'd3, 27'h000003be, 32'h00000400,
  1'd1,  5'd13, 27'h00000040, 5'd0, 27'h00000094, 5'd14, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000031b, 5'd1, 27'h00000001, 5'd21, 27'h00000248, 32'h00000400,
  1'd1,  5'd13, 27'h0000008c, 5'd15, 27'h0000000c, 5'd0, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000140, 5'd15, 27'h000000f9, 5'd14, 27'h000003e0, 32'h00000400,
  1'd1,  5'd10, 27'h00000381, 5'd14, 27'h0000016d, 5'd23, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000271, 5'd25, 27'h000001f7, 5'd3, 27'h00000199, 32'h00000400,
  1'd1,  5'd13, 27'h00000337, 5'd25, 27'h00000019, 5'd14, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002af, 5'd21, 27'h000002af, 5'd24, 27'h00000377, 32'h00000400,
  1'd1,  5'd24, 27'h0000037b, 5'd4, 27'h00000330, 5'd4, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d8, 5'd2, 27'h00000011, 5'd11, 27'h000003ab, 32'h00000400,
  1'd1,  5'd20, 27'h000002fe, 5'd2, 27'h0000009c, 5'd20, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000017b, 5'd14, 27'h000001bd, 5'd3, 27'h00000315, 32'h00000400,
  1'd1,  5'd22, 27'h000001fd, 5'd14, 27'h0000038f, 5'd14, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000370, 5'd10, 27'h000003de, 5'd21, 27'h0000006d, 32'h00000400,
  1'd1,  5'd23, 27'h0000012c, 5'd24, 27'h000000e7, 5'd2, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b6, 5'd24, 27'h00000345, 5'd14, 27'h00000005, 32'h00000400,
  1'd1,  5'd22, 27'h000002eb, 5'd25, 27'h00000078, 5'd23, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000385, 5'd0, 27'h00000317, 5'd8, 27'h000002d9, 32'h00000400,
  1'd1,  5'd2, 27'h0000024c, 5'd3, 27'h00000326, 5'd20, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000014, 5'd1, 27'h000000a6, 5'd27, 27'h0000012f, 32'h00000400,
  1'd1,  5'd2, 27'h000002b9, 5'd11, 27'h000003d8, 5'd8, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000272, 5'd11, 27'h000000e0, 5'd16, 27'h000003c1, 32'h00000400,
  1'd1,  5'd0, 27'h000002ad, 5'd11, 27'h000000c5, 5'd29, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000161, 5'd24, 27'h00000242, 5'd7, 27'h000003e2, 32'h00000400,
  1'd1,  5'd5, 27'h0000001e, 5'd21, 27'h0000010f, 5'd15, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000295, 5'd24, 27'h00000217, 5'd30, 27'h000002c3, 32'h00000400,
  1'd1,  5'd10, 27'h0000035e, 5'd3, 27'h000001ae, 5'd6, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b7, 5'd2, 27'h000001e6, 5'd16, 27'h000002bb, 32'h00000400,
  1'd1,  5'd10, 27'h00000347, 5'd0, 27'h0000022a, 5'd29, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009f, 5'd10, 27'h0000024d, 5'd8, 27'h0000010c, 32'h00000400,
  1'd1,  5'd11, 27'h00000157, 5'd12, 27'h00000347, 5'd15, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001a7, 5'd13, 27'h000001d3, 5'd29, 27'h00000313, 32'h00000400,
  1'd1,  5'd11, 27'h00000253, 5'd22, 27'h0000019f, 5'd6, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000133, 5'd25, 27'h000001fe, 5'd20, 27'h000000c6, 32'h00000400,
  1'd1,  5'd13, 27'h00000183, 5'd24, 27'h000003b8, 5'd28, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000de, 5'd0, 27'h00000137, 5'd5, 27'h000003d4, 32'h00000400,
  1'd1,  5'd25, 27'h0000025d, 5'd3, 27'h000000bf, 5'd19, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000011c, 5'd5, 27'h00000027, 5'd26, 27'h00000344, 32'h00000400,
  1'd1,  5'd23, 27'h000003ed, 5'd12, 27'h00000142, 5'd6, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000312, 5'd10, 27'h0000015b, 5'd17, 27'h000001f5, 32'h00000400,
  1'd1,  5'd21, 27'h0000020f, 5'd13, 27'h000002bf, 5'd25, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000165, 5'd25, 27'h000001d4, 5'd8, 27'h0000035d, 32'h00000400,
  1'd1,  5'd21, 27'h000003bb, 5'd23, 27'h00000381, 5'd15, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003be, 5'd25, 27'h00000217, 5'd27, 27'h00000215, 32'h00000400,
  1'd1,  5'd4, 27'h000002b6, 5'd9, 27'h000002cb, 5'd3, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000264, 5'd8, 27'h000003ac, 5'd14, 27'h000000c9, 32'h00000400,
  1'd1,  5'd1, 27'h0000028d, 5'd6, 27'h0000031e, 5'd25, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000150, 5'd17, 27'h00000102, 5'd4, 27'h00000284, 32'h00000400,
  1'd1,  5'd1, 27'h00000091, 5'd16, 27'h000001c1, 5'd13, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000157, 5'd16, 27'h0000019c, 5'd22, 27'h000000df, 32'h00000400,
  1'd1,  5'd0, 27'h00000358, 5'd27, 27'h000002ca, 5'd2, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000099, 5'd30, 27'h00000354, 5'd11, 27'h00000039, 32'h00000400,
  1'd1,  5'd0, 27'h00000260, 5'd27, 27'h0000031f, 5'd23, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001d7, 5'd9, 27'h000000f2, 5'd4, 27'h00000331, 32'h00000400,
  1'd1,  5'd12, 27'h0000022c, 5'd7, 27'h000003b9, 5'd15, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ae, 5'd8, 27'h000003ac, 5'd24, 27'h0000004e, 32'h00000400,
  1'd1,  5'd11, 27'h000002ae, 5'd16, 27'h00000374, 5'd0, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000080, 5'd15, 27'h0000020c, 5'd13, 27'h00000159, 32'h00000400,
  1'd1,  5'd13, 27'h00000270, 5'd18, 27'h00000117, 5'd25, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000035a, 5'd26, 27'h000001c2, 5'd3, 27'h0000031e, 32'h00000400,
  1'd1,  5'd14, 27'h000002e2, 5'd26, 27'h000000bc, 5'd11, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000062, 5'd28, 27'h000001d5, 5'd25, 27'h0000002a, 32'h00000400,
  1'd1,  5'd21, 27'h00000171, 5'd6, 27'h0000001d, 5'd1, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000026f, 5'd8, 27'h000003e5, 5'd13, 27'h000003c0, 32'h00000400,
  1'd1,  5'd25, 27'h000001ab, 5'd5, 27'h0000021d, 5'd21, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b0, 5'd15, 27'h0000023f, 5'd0, 27'h000002dd, 32'h00000400,
  1'd1,  5'd22, 27'h00000041, 5'd18, 27'h00000010, 5'd12, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000024c, 5'd16, 27'h000001d1, 5'd21, 27'h00000006, 32'h00000400,
  1'd1,  5'd24, 27'h0000006c, 5'd30, 27'h00000092, 5'd0, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001c1, 5'd29, 27'h0000006a, 5'd13, 27'h00000129, 32'h00000400,
  1'd1,  5'd21, 27'h00000123, 5'd27, 27'h0000039d, 5'd24, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003df, 5'd9, 27'h00000290, 5'd9, 27'h000003c6, 32'h00000400,
  1'd1,  5'd2, 27'h000001d0, 5'd5, 27'h0000030b, 5'd18, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000076, 5'd7, 27'h000002d7, 5'd29, 27'h000000f3, 32'h00000400,
  1'd1,  5'd0, 27'h00000235, 5'd17, 27'h000003ac, 5'd9, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b0, 5'd18, 27'h0000016e, 5'd19, 27'h000001b4, 32'h00000400,
  1'd1,  5'd2, 27'h00000141, 5'd17, 27'h0000016a, 5'd28, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000111, 5'd28, 27'h00000353, 5'd10, 27'h000000d7, 32'h00000400,
  1'd1,  5'd2, 27'h00000048, 5'd26, 27'h0000022b, 5'd20, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000000b, 5'd27, 27'h0000038a, 5'd27, 27'h000000dc, 32'h00000400,
  1'd1,  5'd15, 27'h0000008b, 5'd6, 27'h0000033c, 5'd6, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000275, 5'd5, 27'h000003a9, 5'd19, 27'h000003f0, 32'h00000400,
  1'd1,  5'd12, 27'h000000c6, 5'd10, 27'h0000010d, 5'd30, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000178, 5'd18, 27'h00000056, 5'd6, 27'h000003e8, 32'h00000400,
  1'd1,  5'd11, 27'h000001ce, 5'd16, 27'h000001de, 5'd18, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000033c, 5'd20, 27'h0000029f, 5'd27, 27'h00000227, 32'h00000400,
  1'd1,  5'd14, 27'h000001fe, 5'd29, 27'h000000a8, 5'd8, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000032a, 5'd27, 27'h00000194, 5'd15, 27'h0000023e, 32'h00000400,
  1'd1,  5'd11, 27'h0000017e, 5'd29, 27'h000003a0, 5'd29, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000254, 5'd7, 27'h00000249, 5'd7, 27'h000003f5, 32'h00000400,
  1'd1,  5'd23, 27'h00000185, 5'd6, 27'h00000312, 5'd19, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ec, 5'd6, 27'h000003f0, 5'd27, 27'h000000ec, 32'h00000400,
  1'd1,  5'd23, 27'h00000344, 5'd17, 27'h000000b2, 5'd8, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000009b, 5'd16, 27'h00000015, 5'd19, 27'h00000104, 32'h00000400,
  1'd1,  5'd23, 27'h000000a9, 5'd16, 27'h00000327, 5'd26, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000017e, 5'd30, 27'h000002e1, 5'd5, 27'h000003a3, 32'h00000400,
  1'd1,  5'd25, 27'h00000234, 5'd30, 27'h00000341, 5'd20, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000198, 5'd26, 27'h000002f3, 5'd29, 27'h00000334, 32'h00000400,
  1'd1,  5'd10, 27'h000000fb, 5'd3, 27'h00000353, 5'd6, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000011d, 5'd0, 27'h00000122, 5'd17, 27'h00000398, 32'h00000400,
  1'd1,  5'd9, 27'h0000022f, 5'd0, 27'h0000004c, 5'd26, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003fd, 5'd12, 27'h000003a6, 5'd2, 27'h000002c0, 32'h00000400,
  1'd1,  5'd6, 27'h0000008d, 5'd13, 27'h000001f0, 5'd11, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000135, 5'd10, 27'h000002ef, 5'd25, 27'h0000033a, 32'h00000400,
  1'd1,  5'd9, 27'h00000005, 5'd21, 27'h0000028b, 5'd2, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000013a, 5'd24, 27'h0000024b, 5'd10, 27'h00000247, 32'h00000400,
  1'd1,  5'd7, 27'h000001e5, 5'd20, 27'h000003ae, 5'd22, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d4, 5'd4, 27'h00000189, 5'd5, 27'h000003c1, 32'h00000400,
  1'd1,  5'd19, 27'h000003ff, 5'd4, 27'h000002f3, 5'd16, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a5, 5'd4, 27'h000002ba, 5'd29, 27'h0000014b, 32'h00000400,
  1'd1,  5'd19, 27'h00000023, 5'd14, 27'h00000004, 5'd1, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f1, 5'd14, 27'h00000362, 5'd13, 27'h000003ce, 32'h00000400,
  1'd1,  5'd19, 27'h00000207, 5'd11, 27'h000001d4, 5'd22, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000031d, 5'd24, 27'h000003c8, 5'd0, 27'h00000071, 32'h00000400,
  1'd1,  5'd15, 27'h000003f6, 5'd23, 27'h00000100, 5'd14, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000193, 5'd22, 27'h0000020c, 5'd23, 27'h0000032f, 32'h00000400,
  1'd1,  5'd27, 27'h000002bb, 5'd4, 27'h000000e1, 5'd3, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000008, 5'd2, 27'h00000206, 5'd15, 27'h0000014c, 32'h00000400,
  1'd1,  5'd28, 27'h000001b6, 5'd2, 27'h0000025b, 5'd24, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002cf, 5'd10, 27'h00000369, 5'd1, 27'h000001b3, 32'h00000400,
  1'd1,  5'd29, 27'h0000039d, 5'd15, 27'h000001a3, 5'd10, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000fc, 5'd13, 27'h00000240, 5'd20, 27'h0000030c, 32'h00000400,
  1'd1,  5'd26, 27'h00000041, 5'd24, 27'h00000390, 5'd3, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002af, 5'd22, 27'h00000137, 5'd14, 27'h0000026f, 32'h00000400,
  1'd1,  5'd29, 27'h000001d7, 5'd25, 27'h000000fb, 5'd25, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003df, 5'd0, 27'h000000a1, 5'd3, 27'h000001c5, 32'h00000400,
  1'd1,  5'd6, 27'h0000019b, 5'd0, 27'h000001e0, 5'd14, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000005e, 5'd5, 27'h0000008e, 5'd22, 27'h000001c5, 32'h00000400,
  1'd1,  5'd9, 27'h000000cc, 5'd12, 27'h00000203, 5'd9, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000039e, 5'd12, 27'h000003fb, 5'd16, 27'h00000197, 32'h00000400,
  1'd1,  5'd7, 27'h0000027c, 5'd12, 27'h0000023e, 5'd28, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000028e, 5'd23, 27'h000002ea, 5'd9, 27'h0000010c, 32'h00000400,
  1'd1,  5'd7, 27'h00000358, 5'd25, 27'h000001d8, 5'd19, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007c, 5'd21, 27'h0000026a, 5'd28, 27'h0000030c, 32'h00000400,
  1'd1,  5'd20, 27'h00000164, 5'd1, 27'h00000109, 5'd3, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000133, 5'd3, 27'h00000337, 5'd11, 27'h00000309, 32'h00000400,
  1'd1,  5'd19, 27'h000001bc, 5'd0, 27'h00000201, 5'd20, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000023a, 5'd15, 27'h00000191, 5'd7, 27'h000003e6, 32'h00000400,
  1'd1,  5'd15, 27'h000003ca, 5'd11, 27'h00000305, 5'd18, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000034b, 5'd12, 27'h00000183, 5'd29, 27'h0000008f, 32'h00000400,
  1'd1,  5'd16, 27'h000000d0, 5'd22, 27'h00000123, 5'd8, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000352, 5'd24, 27'h00000177, 5'd17, 27'h0000005a, 32'h00000400,
  1'd1,  5'd17, 27'h000002c6, 5'd24, 27'h00000317, 5'd29, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000036, 5'd5, 27'h0000005a, 5'd7, 27'h00000214, 32'h00000400,
  1'd1,  5'd29, 27'h0000012e, 5'd4, 27'h00000001, 5'd16, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000300, 5'd2, 27'h000002b3, 5'd30, 27'h00000140, 32'h00000400,
  1'd1,  5'd29, 27'h000003e1, 5'd11, 27'h000002e4, 5'd9, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000155, 5'd12, 27'h00000374, 5'd19, 27'h0000011e, 32'h00000400,
  1'd1,  5'd30, 27'h00000367, 5'd13, 27'h00000035, 5'd28, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000011d, 5'd21, 27'h00000111, 5'd8, 27'h00000377, 32'h00000400,
  1'd1,  5'd30, 27'h00000085, 5'd24, 27'h00000192, 5'd17, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ef, 5'd22, 27'h00000394, 5'd29, 27'h0000035a, 32'h00000400,
  1'd1,  5'd8, 27'h0000022c, 5'd7, 27'h000002bc, 5'd2, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000158, 5'd10, 27'h0000007f, 5'd15, 27'h00000098, 32'h00000400,
  1'd1,  5'd5, 27'h000002b7, 5'd9, 27'h00000230, 5'd23, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000351, 5'd16, 27'h00000220, 5'd1, 27'h0000010e, 32'h00000400,
  1'd1,  5'd8, 27'h00000023, 5'd17, 27'h0000038e, 5'd14, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000009a, 5'd18, 27'h000001f4, 5'd23, 27'h000002c9, 32'h00000400,
  1'd1,  5'd6, 27'h000000d3, 5'd27, 27'h00000026, 5'd2, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001cd, 5'd28, 27'h00000051, 5'd12, 27'h00000333, 32'h00000400,
  1'd1,  5'd8, 27'h0000003c, 5'd29, 27'h000000f5, 5'd22, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000023f, 5'd9, 27'h000000b4, 5'd0, 27'h00000233, 32'h00000400,
  1'd1,  5'd17, 27'h000003f3, 5'd6, 27'h00000172, 5'd11, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000023d, 5'd6, 27'h00000016, 5'd24, 27'h00000044, 32'h00000400,
  1'd1,  5'd17, 27'h00000230, 5'd17, 27'h00000341, 5'd0, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ba, 5'd19, 27'h000000a5, 5'd13, 27'h000003a9, 32'h00000400,
  1'd1,  5'd16, 27'h000002cd, 5'd20, 27'h000000ce, 5'd22, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032c, 5'd27, 27'h0000008e, 5'd0, 27'h000002fc, 32'h00000400,
  1'd1,  5'd17, 27'h000001af, 5'd26, 27'h00000277, 5'd12, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000010b, 5'd28, 27'h00000177, 5'd24, 27'h000003c4, 32'h00000400,
  1'd1,  5'd28, 27'h0000024b, 5'd8, 27'h00000196, 5'd4, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d7, 5'd7, 27'h0000037b, 5'd11, 27'h000002fc, 32'h00000400,
  1'd1,  5'd26, 27'h000001d5, 5'd7, 27'h0000030c, 5'd22, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017c, 5'd16, 27'h00000164, 5'd2, 27'h0000027f, 32'h00000400,
  1'd1,  5'd29, 27'h00000067, 5'd19, 27'h00000123, 5'd12, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000007f, 5'd18, 27'h00000354, 5'd21, 27'h00000151, 32'h00000400,
  1'd1,  5'd25, 27'h0000035b, 5'd29, 27'h00000236, 5'd4, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a8, 5'd29, 27'h000002a4, 5'd10, 27'h000001b5, 32'h00000400,
  1'd1,  5'd27, 27'h0000021f, 5'd26, 27'h0000000e, 5'd25, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000212, 5'd8, 27'h00000119, 5'd7, 27'h00000343, 32'h00000400,
  1'd1,  5'd6, 27'h000001ad, 5'd8, 27'h00000120, 5'd18, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001cd, 5'd5, 27'h00000227, 5'd29, 27'h000001b6, 32'h00000400,
  1'd1,  5'd6, 27'h0000022f, 5'd15, 27'h0000036b, 5'd7, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000131, 5'd19, 27'h00000055, 5'd19, 27'h00000344, 32'h00000400,
  1'd1,  5'd5, 27'h00000387, 5'd16, 27'h00000198, 5'd27, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000df, 5'd26, 27'h000001c5, 5'd9, 27'h00000078, 32'h00000400,
  1'd1,  5'd6, 27'h000003c8, 5'd28, 27'h00000183, 5'd16, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000024d, 5'd29, 27'h0000000c, 5'd26, 27'h0000003a, 32'h00000400,
  1'd1,  5'd18, 27'h00000296, 5'd9, 27'h00000359, 5'd6, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000016b, 5'd9, 27'h0000035d, 5'd15, 27'h000003b1, 32'h00000400,
  1'd1,  5'd20, 27'h000001a7, 5'd7, 27'h00000319, 5'd25, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f8, 5'd18, 27'h00000122, 5'd5, 27'h0000018f, 32'h00000400,
  1'd1,  5'd15, 27'h0000033a, 5'd19, 27'h00000022, 5'd20, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000074, 5'd17, 27'h0000003a, 5'd27, 27'h000002ce, 32'h00000400,
  1'd1,  5'd18, 27'h0000002a, 5'd29, 27'h0000013f, 5'd5, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000102, 5'd27, 27'h0000028f, 5'd19, 27'h000000fe, 32'h00000400,
  1'd1,  5'd16, 27'h00000164, 5'd26, 27'h0000035b, 5'd27, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000018c, 5'd7, 27'h00000301, 5'd8, 27'h000003e7, 32'h00000400,
  1'd1,  5'd29, 27'h00000265, 5'd6, 27'h00000144, 5'd19, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000176, 5'd7, 27'h0000017e, 5'd26, 27'h00000275, 32'h00000400,
  1'd1,  5'd29, 27'h00000101, 5'd19, 27'h00000264, 5'd5, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000037, 5'd19, 27'h00000153, 5'd19, 27'h0000015a, 32'h00000400,
  1'd1,  5'd29, 27'h000000b8, 5'd16, 27'h000003fd, 5'd27, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a3, 5'd29, 27'h0000020e, 5'd8, 27'h00000380, 32'h00000400,
  1'd1,  5'd30, 27'h0000007d, 5'd27, 27'h000001f5, 5'd20, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000036c, 5'd27, 27'h00000215, 5'd29, 27'h000003a9, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000000d8, 5'd3, 27'h00000100, 5'd3, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000220, 5'd3, 27'h000003f7, 5'd14, 27'h000003c9, 32'h00000400,
  1'd1,  5'd4, 27'h00000066, 5'd4, 27'h000002c4, 5'd21, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f0, 5'd14, 27'h0000037e, 5'd4, 27'h00000206, 32'h00000400,
  1'd1,  5'd3, 27'h000002f8, 5'd14, 27'h000003f7, 5'd13, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000c0, 5'd14, 27'h00000287, 5'd21, 27'h0000026f, 32'h00000400,
  1'd1,  5'd4, 27'h00000132, 5'd25, 27'h000000cc, 5'd3, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ea, 5'd23, 27'h000000bf, 5'd13, 27'h00000026, 32'h00000400,
  1'd1,  5'd0, 27'h0000010e, 5'd23, 27'h0000026f, 5'd25, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000270, 5'd1, 27'h0000004b, 5'd1, 27'h00000178, 32'h00000400,
  1'd1,  5'd14, 27'h000000f8, 5'd2, 27'h0000018f, 5'd12, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000364, 5'd2, 27'h000000d7, 5'd25, 27'h00000009, 32'h00000400,
  1'd1,  5'd13, 27'h000002b4, 5'd10, 27'h000002aa, 5'd4, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f1, 5'd11, 27'h000003f1, 5'd11, 27'h0000039a, 32'h00000400,
  1'd1,  5'd10, 27'h0000015a, 5'd13, 27'h000002b1, 5'd25, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000012e, 5'd22, 27'h00000302, 5'd4, 27'h000000ce, 32'h00000400,
  1'd1,  5'd12, 27'h00000381, 5'd25, 27'h0000001a, 5'd12, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002f7, 5'd22, 27'h00000117, 5'd23, 27'h000003f5, 32'h00000400,
  1'd1,  5'd24, 27'h00000237, 5'd1, 27'h00000135, 5'd4, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000035b, 5'd0, 27'h000002c8, 5'd11, 27'h00000227, 32'h00000400,
  1'd1,  5'd25, 27'h000000a2, 5'd3, 27'h000000e3, 5'd22, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b9, 5'd12, 27'h00000077, 5'd4, 27'h00000152, 32'h00000400,
  1'd1,  5'd21, 27'h00000268, 5'd12, 27'h00000028, 5'd14, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000026c, 5'd11, 27'h00000321, 5'd21, 27'h000001e8, 32'h00000400,
  1'd1,  5'd22, 27'h00000120, 5'd24, 27'h000002e2, 5'd1, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000367, 5'd25, 27'h000000c1, 5'd13, 27'h0000003b, 32'h00000400,
  1'd1,  5'd22, 27'h0000019f, 5'd24, 27'h0000004c, 5'd21, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000309, 5'd5, 27'h00000098, 5'd5, 27'h000002f9, 32'h00000400,
  1'd1,  5'd1, 27'h000003e3, 5'd4, 27'h00000111, 5'd15, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000033, 5'd1, 27'h000000af, 5'd30, 27'h000001f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000163, 5'd10, 27'h0000024d, 5'd6, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000388, 5'd15, 27'h000000a7, 5'd20, 27'h0000019a, 32'h00000400,
  1'd1,  5'd2, 27'h00000275, 5'd10, 27'h00000170, 5'd28, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000306, 5'd22, 27'h00000074, 5'd8, 27'h000002e4, 32'h00000400,
  1'd1,  5'd4, 27'h00000314, 5'd22, 27'h000000bc, 5'd17, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017c, 5'd23, 27'h0000001a, 5'd26, 27'h00000387, 32'h00000400,
  1'd1,  5'd14, 27'h0000000c, 5'd4, 27'h00000200, 5'd6, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f1, 5'd1, 27'h000003e4, 5'd19, 27'h000001a0, 32'h00000400,
  1'd1,  5'd12, 27'h0000029f, 5'd0, 27'h000003cf, 5'd27, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000162, 5'd11, 27'h00000030, 5'd9, 27'h000001d5, 32'h00000400,
  1'd1,  5'd11, 27'h00000168, 5'd11, 27'h000002e7, 5'd19, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000006a, 5'd10, 27'h0000034c, 5'd26, 27'h000000ba, 32'h00000400,
  1'd1,  5'd11, 27'h00000316, 5'd23, 27'h0000030d, 5'd9, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001b0, 5'd22, 27'h00000062, 5'd18, 27'h00000342, 32'h00000400,
  1'd1,  5'd14, 27'h000001e9, 5'd24, 27'h00000012, 5'd28, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c5, 5'd3, 27'h0000012a, 5'd7, 27'h000003f7, 32'h00000400,
  1'd1,  5'd23, 27'h00000075, 5'd4, 27'h00000077, 5'd20, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ab, 5'd1, 27'h000000fb, 5'd28, 27'h0000014d, 32'h00000400,
  1'd1,  5'd24, 27'h000001bc, 5'd10, 27'h000002d0, 5'd7, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000028a, 5'd14, 27'h00000091, 5'd18, 27'h00000214, 32'h00000400,
  1'd1,  5'd24, 27'h00000298, 5'd13, 27'h000001e0, 5'd29, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002fa, 5'd24, 27'h000001e1, 5'd7, 27'h0000008b, 32'h00000400,
  1'd1,  5'd20, 27'h00000361, 5'd25, 27'h000001e8, 5'd17, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000001b, 5'd21, 27'h000003ce, 5'd26, 27'h000000a2, 32'h00000400,
  1'd1,  5'd2, 27'h000002a6, 5'd10, 27'h00000065, 5'd3, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000166, 5'd6, 27'h00000301, 5'd11, 27'h000000f7, 32'h00000400,
  1'd1,  5'd2, 27'h000003d9, 5'd8, 27'h00000221, 5'd21, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000014b, 5'd19, 27'h0000015c, 5'd4, 27'h000000ba, 32'h00000400,
  1'd1,  5'd4, 27'h000003db, 5'd19, 27'h000003aa, 5'd14, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002e1, 5'd16, 27'h000003b8, 5'd23, 27'h000003bb, 32'h00000400,
  1'd1,  5'd2, 27'h0000037c, 5'd29, 27'h0000029c, 5'd2, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000212, 5'd26, 27'h00000128, 5'd15, 27'h0000008a, 32'h00000400,
  1'd1,  5'd3, 27'h00000059, 5'd26, 27'h000003c9, 5'd24, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000197, 5'd8, 27'h00000188, 5'd4, 27'h000003d2, 32'h00000400,
  1'd1,  5'd15, 27'h0000009a, 5'd8, 27'h0000002f, 5'd13, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000216, 5'd6, 27'h000003be, 5'd25, 27'h000001d7, 32'h00000400,
  1'd1,  5'd10, 27'h0000036d, 5'd15, 27'h00000305, 5'd1, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000268, 5'd17, 27'h0000019e, 5'd12, 27'h00000263, 32'h00000400,
  1'd1,  5'd13, 27'h000002d0, 5'd16, 27'h000003a7, 5'd25, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000af, 5'd26, 27'h00000316, 5'd3, 27'h0000021a, 32'h00000400,
  1'd1,  5'd13, 27'h000001c1, 5'd26, 27'h000000b6, 5'd11, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000178, 5'd27, 27'h00000103, 5'd23, 27'h0000015a, 32'h00000400,
  1'd1,  5'd25, 27'h0000007c, 5'd5, 27'h000001c2, 5'd2, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000003, 5'd7, 27'h000003b4, 5'd11, 27'h000000a5, 32'h00000400,
  1'd1,  5'd23, 27'h000002ea, 5'd6, 27'h00000225, 5'd23, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001cf, 5'd16, 27'h00000102, 5'd0, 27'h00000243, 32'h00000400,
  1'd1,  5'd21, 27'h00000076, 5'd19, 27'h0000033e, 5'd15, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000002d, 5'd19, 27'h0000013e, 5'd23, 27'h000001e2, 32'h00000400,
  1'd1,  5'd22, 27'h0000024a, 5'd30, 27'h0000027f, 5'd0, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000055, 5'd27, 27'h0000011c, 5'd11, 27'h000000e1, 32'h00000400,
  1'd1,  5'd24, 27'h00000244, 5'd27, 27'h000000e4, 5'd25, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f9, 5'd5, 27'h000003e4, 5'd10, 27'h00000099, 32'h00000400,
  1'd1,  5'd4, 27'h00000108, 5'd6, 27'h00000074, 5'd17, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001f4, 5'd10, 27'h000000cd, 5'd28, 27'h00000313, 32'h00000400,
  1'd1,  5'd3, 27'h0000015b, 5'd16, 27'h0000005a, 5'd8, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b2, 5'd18, 27'h00000102, 5'd16, 27'h00000325, 32'h00000400,
  1'd1,  5'd0, 27'h000001a5, 5'd19, 27'h0000002a, 5'd28, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018a, 5'd30, 27'h000002fa, 5'd5, 27'h0000017a, 32'h00000400,
  1'd1,  5'd0, 27'h00000050, 5'd26, 27'h00000122, 5'd16, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000178, 5'd30, 27'h0000001e, 5'd29, 27'h000002c6, 32'h00000400,
  1'd1,  5'd12, 27'h000002f0, 5'd9, 27'h000002a7, 5'd8, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ac, 5'd6, 27'h0000020d, 5'd16, 27'h000003fe, 32'h00000400,
  1'd1,  5'd10, 27'h000001c2, 5'd10, 27'h00000150, 5'd26, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ce, 5'd19, 27'h0000039f, 5'd7, 27'h000002f6, 32'h00000400,
  1'd1,  5'd10, 27'h000003c8, 5'd18, 27'h00000383, 5'd16, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035f, 5'd15, 27'h00000275, 5'd27, 27'h000001a4, 32'h00000400,
  1'd1,  5'd10, 27'h000003f1, 5'd28, 27'h0000031c, 5'd7, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000319, 5'd27, 27'h00000095, 5'd17, 27'h000003f8, 32'h00000400,
  1'd1,  5'd14, 27'h0000029a, 5'd30, 27'h00000060, 5'd30, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000185, 5'd7, 27'h00000069, 5'd6, 27'h000003c9, 32'h00000400,
  1'd1,  5'd24, 27'h0000023d, 5'd7, 27'h0000007c, 5'd17, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000000c, 5'd8, 27'h0000035e, 5'd28, 27'h00000050, 32'h00000400,
  1'd1,  5'd22, 27'h00000363, 5'd18, 27'h000002b6, 5'd6, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f8, 5'd18, 27'h000002f0, 5'd16, 27'h000003c3, 32'h00000400,
  1'd1,  5'd24, 27'h0000018f, 5'd15, 27'h00000287, 5'd29, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000022f, 5'd27, 27'h00000004, 5'd7, 27'h00000161, 32'h00000400,
  1'd1,  5'd25, 27'h000001be, 5'd28, 27'h000001ce, 5'd17, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ab, 5'd26, 27'h0000028d, 5'd27, 27'h0000023a, 32'h00000400,
  1'd1,  5'd8, 27'h000001b6, 5'd1, 27'h0000036f, 5'd7, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021c, 5'd3, 27'h00000333, 5'd17, 27'h0000024c, 32'h00000400,
  1'd1,  5'd7, 27'h000001b4, 5'd4, 27'h00000340, 5'd29, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000226, 5'd11, 27'h00000243, 5'd1, 27'h00000254, 32'h00000400,
  1'd1,  5'd6, 27'h000001b1, 5'd14, 27'h00000099, 5'd12, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cf, 5'd12, 27'h0000013a, 5'd23, 27'h000001fa, 32'h00000400,
  1'd1,  5'd7, 27'h00000342, 5'd24, 27'h0000039d, 5'd0, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000027, 5'd24, 27'h000001d5, 5'd11, 27'h000000f9, 32'h00000400,
  1'd1,  5'd9, 27'h00000326, 5'd23, 27'h000001d3, 5'd21, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000114, 5'd3, 27'h0000031e, 5'd8, 27'h000001bf, 32'h00000400,
  1'd1,  5'd19, 27'h00000028, 5'd4, 27'h000002b9, 5'd17, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000023a, 5'd4, 27'h00000016, 5'd28, 27'h0000023a, 32'h00000400,
  1'd1,  5'd16, 27'h000001dd, 5'd13, 27'h0000012f, 5'd2, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001fb, 5'd13, 27'h000002da, 5'd15, 27'h0000016a, 32'h00000400,
  1'd1,  5'd19, 27'h00000390, 5'd12, 27'h00000095, 5'd24, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029d, 5'd23, 27'h000001a0, 5'd4, 27'h0000035c, 32'h00000400,
  1'd1,  5'd17, 27'h000003c3, 5'd23, 27'h0000005d, 5'd13, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000019d, 5'd22, 27'h000003a8, 5'd24, 27'h000003dd, 32'h00000400,
  1'd1,  5'd30, 27'h000002f6, 5'd0, 27'h000001da, 5'd1, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b2, 5'd3, 27'h0000025d, 5'd11, 27'h0000011d, 32'h00000400,
  1'd1,  5'd28, 27'h000001c3, 5'd4, 27'h0000023e, 5'd22, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000f7, 5'd13, 27'h0000019f, 5'd1, 27'h0000002c, 32'h00000400,
  1'd1,  5'd29, 27'h0000015e, 5'd14, 27'h000001f3, 5'd10, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000378, 5'd14, 27'h00000388, 5'd23, 27'h000003a9, 32'h00000400,
  1'd1,  5'd25, 27'h000003c5, 5'd20, 27'h0000036e, 5'd4, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e9, 5'd25, 27'h00000080, 5'd14, 27'h0000039a, 32'h00000400,
  1'd1,  5'd27, 27'h00000330, 5'd20, 27'h000003e1, 5'd22, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000014b, 5'd0, 27'h000001ff, 5'd2, 27'h000002c8, 32'h00000400,
  1'd1,  5'd5, 27'h0000016e, 5'd4, 27'h000001af, 5'd12, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e7, 5'd4, 27'h0000020c, 5'd24, 27'h0000022c, 32'h00000400,
  1'd1,  5'd9, 27'h00000113, 5'd13, 27'h000001d8, 5'd8, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000007d, 5'd14, 27'h000001f6, 5'd17, 27'h000000bc, 32'h00000400,
  1'd1,  5'd8, 27'h00000179, 5'd15, 27'h000000ba, 5'd27, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000024, 5'd25, 27'h00000241, 5'd6, 27'h000003db, 32'h00000400,
  1'd1,  5'd9, 27'h000000d4, 5'd24, 27'h000001ef, 5'd19, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001ab, 5'd24, 27'h000002f1, 5'd25, 27'h00000371, 32'h00000400,
  1'd1,  5'd19, 27'h0000033e, 5'd0, 27'h000000de, 5'd2, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000129, 5'd2, 27'h00000318, 5'd13, 27'h000003d5, 32'h00000400,
  1'd1,  5'd18, 27'h000003cd, 5'd1, 27'h00000099, 5'd24, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000171, 5'd12, 27'h0000004d, 5'd9, 27'h000003b4, 32'h00000400,
  1'd1,  5'd19, 27'h00000257, 5'd11, 27'h00000299, 5'd16, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f5, 5'd13, 27'h0000024a, 5'd30, 27'h0000007c, 32'h00000400,
  1'd1,  5'd20, 27'h000001d7, 5'd23, 27'h0000031a, 5'd9, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000011c, 5'd23, 27'h000001e2, 5'd18, 27'h00000117, 32'h00000400,
  1'd1,  5'd16, 27'h000000da, 5'd24, 27'h00000380, 5'd29, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017d, 5'd0, 27'h00000063, 5'd7, 27'h0000026a, 32'h00000400,
  1'd1,  5'd27, 27'h000000a7, 5'd2, 27'h0000021b, 5'd16, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000018a, 5'd2, 27'h0000001f, 5'd30, 27'h0000000e, 32'h00000400,
  1'd1,  5'd29, 27'h00000053, 5'd12, 27'h0000033d, 5'd5, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000165, 5'd11, 27'h000001c2, 5'd18, 27'h000001d7, 32'h00000400,
  1'd1,  5'd30, 27'h0000002f, 5'd14, 27'h00000396, 5'd27, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a5, 5'd22, 27'h000001f9, 5'd6, 27'h0000037f, 32'h00000400,
  1'd1,  5'd30, 27'h0000022e, 5'd25, 27'h00000045, 5'd16, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003c3, 5'd22, 27'h000001fe, 5'd29, 27'h00000079, 32'h00000400,
  1'd1,  5'd5, 27'h00000272, 5'd7, 27'h0000012e, 5'd4, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000000c, 5'd8, 27'h00000099, 5'd11, 27'h00000057, 32'h00000400,
  1'd1,  5'd10, 27'h0000014a, 5'd6, 27'h000001f1, 5'd22, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000189, 5'd15, 27'h0000034e, 5'd2, 27'h000000c1, 32'h00000400,
  1'd1,  5'd5, 27'h000003cc, 5'd16, 27'h00000149, 5'd14, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c3, 5'd19, 27'h00000153, 5'd24, 27'h000003db, 32'h00000400,
  1'd1,  5'd5, 27'h0000018d, 5'd29, 27'h0000006d, 5'd1, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b3, 5'd27, 27'h000003fa, 5'd15, 27'h0000015f, 32'h00000400,
  1'd1,  5'd6, 27'h0000023d, 5'd28, 27'h000002c5, 5'd23, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e9, 5'd7, 27'h0000028f, 5'd4, 27'h00000352, 32'h00000400,
  1'd1,  5'd20, 27'h000001d9, 5'd9, 27'h000001d9, 5'd11, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c0, 5'd7, 27'h000000f7, 5'd21, 27'h00000368, 32'h00000400,
  1'd1,  5'd19, 27'h00000347, 5'd16, 27'h000001f8, 5'd3, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000037d, 5'd15, 27'h00000296, 5'd11, 27'h000000f4, 32'h00000400,
  1'd1,  5'd19, 27'h00000014, 5'd16, 27'h00000121, 5'd21, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000182, 5'd30, 27'h000000d5, 5'd4, 27'h00000394, 32'h00000400,
  1'd1,  5'd19, 27'h00000223, 5'd27, 27'h000001bc, 5'd11, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000005f, 5'd30, 27'h00000094, 5'd22, 27'h00000069, 32'h00000400,
  1'd1,  5'd29, 27'h000002cb, 5'd8, 27'h000002f0, 5'd1, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000007d, 5'd10, 27'h000000aa, 5'd12, 27'h00000312, 32'h00000400,
  1'd1,  5'd30, 27'h00000365, 5'd5, 27'h00000378, 5'd24, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003bb, 5'd18, 27'h00000008, 5'd0, 27'h000000ae, 32'h00000400,
  1'd1,  5'd27, 27'h00000159, 5'd17, 27'h00000256, 5'd12, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002b9, 5'd20, 27'h000000b3, 5'd21, 27'h000002e7, 32'h00000400,
  1'd1,  5'd29, 27'h00000181, 5'd28, 27'h00000273, 5'd4, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001f5, 5'd26, 27'h000003ad, 5'd15, 27'h00000147, 32'h00000400,
  1'd1,  5'd25, 27'h0000039e, 5'd26, 27'h00000041, 5'd22, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000218, 5'd6, 27'h00000123, 5'd5, 27'h000001c9, 32'h00000400,
  1'd1,  5'd9, 27'h00000136, 5'd9, 27'h000000fb, 5'd19, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000123, 5'd6, 27'h0000001c, 5'd29, 27'h00000055, 32'h00000400,
  1'd1,  5'd5, 27'h00000119, 5'd16, 27'h00000360, 5'd8, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000038f, 5'd18, 27'h00000192, 5'd20, 27'h0000012a, 32'h00000400,
  1'd1,  5'd5, 27'h00000187, 5'd18, 27'h000001e0, 5'd27, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000364, 5'd30, 27'h00000394, 5'd7, 27'h0000006c, 32'h00000400,
  1'd1,  5'd8, 27'h0000038b, 5'd28, 27'h00000022, 5'd16, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002c9, 5'd30, 27'h00000083, 5'd30, 27'h0000033c, 32'h00000400,
  1'd1,  5'd17, 27'h0000031f, 5'd6, 27'h000002f9, 5'd6, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000004, 5'd7, 27'h000002c5, 5'd18, 27'h000000e8, 32'h00000400,
  1'd1,  5'd17, 27'h00000235, 5'd7, 27'h00000365, 5'd28, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d1, 5'd16, 27'h000002fd, 5'd5, 27'h000000f6, 32'h00000400,
  1'd1,  5'd20, 27'h00000085, 5'd19, 27'h0000006e, 5'd17, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000008d, 5'd18, 27'h00000168, 5'd28, 27'h00000196, 32'h00000400,
  1'd1,  5'd17, 27'h00000366, 5'd26, 27'h000002e0, 5'd6, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000039f, 5'd27, 27'h00000257, 5'd17, 27'h00000215, 32'h00000400,
  1'd1,  5'd16, 27'h00000203, 5'd25, 27'h00000399, 5'd27, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000258, 5'd8, 27'h0000031c, 5'd7, 27'h00000247, 32'h00000400,
  1'd1,  5'd30, 27'h00000310, 5'd9, 27'h000002ae, 5'd16, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001cf, 5'd5, 27'h000003eb, 5'd29, 27'h00000105, 32'h00000400,
  1'd1,  5'd29, 27'h00000126, 5'd15, 27'h00000269, 5'd8, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000bd, 5'd17, 27'h000003c0, 5'd18, 27'h0000010d, 32'h00000400,
  1'd1,  5'd27, 27'h000001fe, 5'd17, 27'h0000009b, 5'd29, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034c, 5'd27, 27'h0000030e, 5'd6, 27'h00000213, 32'h00000400,
  1'd1,  5'd28, 27'h000000e8, 5'd27, 27'h000001f3, 5'd20, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000172, 5'd27, 27'h000002c2, 5'd26, 27'h00000121, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003e4, 5'd1, 27'h000001c0, 5'd0, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000002a, 5'd0, 27'h0000018b, 5'd14, 27'h000002b6, 32'h00000400,
  1'd1,  5'd0, 27'h00000177, 5'd4, 27'h000002ce, 5'd23, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000268, 5'd13, 27'h0000007d, 5'd2, 27'h000001a4, 32'h00000400,
  1'd1,  5'd2, 27'h00000132, 5'd11, 27'h00000376, 5'd12, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000097, 5'd10, 27'h000002eb, 5'd25, 27'h0000033e, 32'h00000400,
  1'd1,  5'd0, 27'h000002b7, 5'd22, 27'h000000e1, 5'd4, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000286, 5'd21, 27'h00000363, 5'd10, 27'h000001d5, 32'h00000400,
  1'd1,  5'd5, 27'h00000009, 5'd23, 27'h0000019a, 5'd23, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000054, 5'd2, 27'h000001a5, 5'd0, 27'h000001ab, 32'h00000400,
  1'd1,  5'd14, 27'h0000033c, 5'd5, 27'h0000004d, 5'd11, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000373, 5'd1, 27'h000000ac, 5'd24, 27'h00000356, 32'h00000400,
  1'd1,  5'd13, 27'h0000012a, 5'd11, 27'h00000009, 5'd4, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001fa, 5'd10, 27'h000001b0, 5'd11, 27'h00000118, 32'h00000400,
  1'd1,  5'd10, 27'h00000332, 5'd13, 27'h0000038d, 5'd24, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000bc, 5'd25, 27'h000002d9, 5'd3, 27'h0000012f, 32'h00000400,
  1'd1,  5'd14, 27'h00000095, 5'd23, 27'h0000002a, 5'd13, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000373, 5'd23, 27'h000003c9, 5'd25, 27'h00000109, 32'h00000400,
  1'd1,  5'd24, 27'h00000204, 5'd4, 27'h000003e7, 5'd1, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000021f, 5'd0, 27'h00000174, 5'd15, 27'h00000101, 32'h00000400,
  1'd1,  5'd20, 27'h0000039b, 5'd2, 27'h000003a0, 5'd24, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000130, 5'd12, 27'h00000331, 5'd4, 27'h0000000d, 32'h00000400,
  1'd1,  5'd24, 27'h00000367, 5'd12, 27'h0000008d, 5'd15, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000020, 5'd11, 27'h0000032a, 5'd21, 27'h000001cc, 32'h00000400,
  1'd1,  5'd21, 27'h00000239, 5'd23, 27'h00000005, 5'd3, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000375, 5'd20, 27'h000002eb, 5'd13, 27'h0000004c, 32'h00000400,
  1'd1,  5'd24, 27'h00000313, 5'd24, 27'h0000010d, 5'd21, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a6, 5'd3, 27'h00000172, 5'd7, 27'h000000e4, 32'h00000400,
  1'd1,  5'd1, 27'h00000033, 5'd2, 27'h00000083, 5'd18, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000db, 5'd4, 27'h000002fc, 5'd29, 27'h000001d2, 32'h00000400,
  1'd1,  5'd4, 27'h000003ff, 5'd11, 27'h0000028d, 5'd5, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000031a, 5'd13, 27'h00000243, 5'd17, 27'h000001c2, 32'h00000400,
  1'd1,  5'd2, 27'h000001fc, 5'd11, 27'h0000017b, 5'd27, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c0, 5'd24, 27'h000002f2, 5'd8, 27'h000001bf, 32'h00000400,
  1'd1,  5'd4, 27'h000003c0, 5'd25, 27'h00000159, 5'd19, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000056, 5'd21, 27'h0000033b, 5'd28, 27'h0000026b, 32'h00000400,
  1'd1,  5'd11, 27'h00000083, 5'd2, 27'h000001ed, 5'd8, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000148, 5'd1, 27'h00000346, 5'd20, 27'h00000196, 32'h00000400,
  1'd1,  5'd12, 27'h000000c7, 5'd1, 27'h00000089, 5'd26, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000291, 5'd12, 27'h00000099, 5'd8, 27'h00000276, 32'h00000400,
  1'd1,  5'd12, 27'h00000192, 5'd10, 27'h00000248, 5'd19, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000112, 5'd11, 27'h0000026f, 5'd29, 27'h00000100, 32'h00000400,
  1'd1,  5'd12, 27'h000003f0, 5'd21, 27'h00000024, 5'd6, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002cd, 5'd21, 27'h000002bb, 5'd18, 27'h00000296, 32'h00000400,
  1'd1,  5'd15, 27'h000001ea, 5'd23, 27'h00000352, 5'd30, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000022c, 5'd5, 27'h00000003, 5'd7, 27'h000002c0, 32'h00000400,
  1'd1,  5'd21, 27'h00000349, 5'd0, 27'h00000106, 5'd20, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000230, 5'd1, 27'h0000005f, 5'd26, 27'h000002fa, 32'h00000400,
  1'd1,  5'd22, 27'h000000cb, 5'd13, 27'h000000e4, 5'd7, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000039d, 5'd11, 27'h00000358, 5'd18, 27'h00000001, 32'h00000400,
  1'd1,  5'd21, 27'h00000212, 5'd10, 27'h00000360, 5'd26, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000352, 5'd21, 27'h00000072, 5'd9, 27'h00000347, 32'h00000400,
  1'd1,  5'd21, 27'h0000023a, 5'd24, 27'h00000377, 5'd19, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000182, 5'd25, 27'h000002b7, 5'd27, 27'h0000008d, 32'h00000400,
  1'd1,  5'd3, 27'h000001a0, 5'd7, 27'h0000032e, 5'd3, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000005c, 5'd7, 27'h0000038a, 5'd10, 27'h00000266, 32'h00000400,
  1'd1,  5'd2, 27'h00000024, 5'd9, 27'h000002e1, 5'd22, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000310, 5'd18, 27'h0000018a, 5'd0, 27'h00000119, 32'h00000400,
  1'd1,  5'd3, 27'h00000013, 5'd16, 27'h0000029f, 5'd13, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d0, 5'd17, 27'h0000021c, 5'd22, 27'h0000018a, 32'h00000400,
  1'd1,  5'd0, 27'h0000013a, 5'd27, 27'h00000102, 5'd4, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d3, 5'd30, 27'h00000243, 5'd13, 27'h00000018, 32'h00000400,
  1'd1,  5'd2, 27'h000000bd, 5'd29, 27'h0000013f, 5'd24, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000045, 5'd8, 27'h000001ba, 5'd4, 27'h000000d5, 32'h00000400,
  1'd1,  5'd12, 27'h000001b6, 5'd9, 27'h00000162, 5'd11, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000326, 5'd8, 27'h000002c8, 5'd23, 27'h000000be, 32'h00000400,
  1'd1,  5'd11, 27'h00000354, 5'd16, 27'h0000008e, 5'd4, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000013c, 5'd16, 27'h00000237, 5'd14, 27'h0000022d, 32'h00000400,
  1'd1,  5'd14, 27'h0000030f, 5'd18, 27'h00000116, 5'd21, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001cd, 5'd27, 27'h00000260, 5'd2, 27'h00000171, 32'h00000400,
  1'd1,  5'd11, 27'h0000025c, 5'd29, 27'h00000373, 5'd14, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ef, 5'd30, 27'h00000045, 5'd25, 27'h000000c2, 32'h00000400,
  1'd1,  5'd22, 27'h00000248, 5'd7, 27'h00000346, 5'd3, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000236, 5'd5, 27'h000001ea, 5'd11, 27'h00000369, 32'h00000400,
  1'd1,  5'd22, 27'h00000038, 5'd5, 27'h000003f5, 5'd23, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032a, 5'd17, 27'h000001c6, 5'd4, 27'h00000359, 32'h00000400,
  1'd1,  5'd25, 27'h00000241, 5'd19, 27'h000000b3, 5'd13, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000400, 5'd17, 27'h0000026e, 5'd23, 27'h0000021c, 32'h00000400,
  1'd1,  5'd21, 27'h000003c5, 5'd26, 27'h0000005c, 5'd0, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001cc, 5'd28, 27'h000002a4, 5'd12, 27'h000001b3, 32'h00000400,
  1'd1,  5'd21, 27'h00000074, 5'd29, 27'h000003ee, 5'd23, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038c, 5'd7, 27'h0000014d, 5'd9, 27'h00000099, 32'h00000400,
  1'd1,  5'd2, 27'h0000006a, 5'd10, 27'h00000089, 5'd17, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000200, 5'd8, 27'h00000320, 5'd27, 27'h000001af, 32'h00000400,
  1'd1,  5'd3, 27'h000000bb, 5'd17, 27'h00000382, 5'd7, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b4, 5'd17, 27'h00000224, 5'd20, 27'h00000145, 32'h00000400,
  1'd1,  5'd3, 27'h000001e1, 5'd17, 27'h0000039c, 5'd28, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001fe, 5'd29, 27'h00000083, 5'd9, 27'h0000037b, 32'h00000400,
  1'd1,  5'd4, 27'h000001a1, 5'd26, 27'h000000f5, 5'd16, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000034, 5'd27, 27'h00000034, 5'd28, 27'h000000fa, 32'h00000400,
  1'd1,  5'd11, 27'h00000322, 5'd6, 27'h00000180, 5'd5, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c0, 5'd6, 27'h00000058, 5'd15, 27'h00000255, 32'h00000400,
  1'd1,  5'd13, 27'h0000008e, 5'd9, 27'h000002a9, 5'd30, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d0, 5'd20, 27'h00000219, 5'd7, 27'h00000399, 32'h00000400,
  1'd1,  5'd11, 27'h00000246, 5'd15, 27'h0000026e, 5'd15, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000046, 5'd19, 27'h00000237, 5'd28, 27'h000000a6, 32'h00000400,
  1'd1,  5'd11, 27'h000000f9, 5'd30, 27'h000003df, 5'd6, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e9, 5'd27, 27'h000003f3, 5'd19, 27'h0000035f, 32'h00000400,
  1'd1,  5'd13, 27'h00000012, 5'd25, 27'h000003eb, 5'd27, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000011b, 5'd8, 27'h0000023f, 5'd7, 27'h000002bf, 32'h00000400,
  1'd1,  5'd23, 27'h0000008c, 5'd7, 27'h000002ac, 5'd20, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000367, 5'd6, 27'h0000002c, 5'd28, 27'h00000079, 32'h00000400,
  1'd1,  5'd23, 27'h0000016c, 5'd19, 27'h00000156, 5'd9, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000023e, 5'd19, 27'h00000055, 5'd20, 27'h00000264, 32'h00000400,
  1'd1,  5'd23, 27'h00000043, 5'd18, 27'h00000008, 5'd28, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000021c, 5'd30, 27'h0000039a, 5'd6, 27'h0000006f, 32'h00000400,
  1'd1,  5'd24, 27'h000001dc, 5'd27, 27'h000003d1, 5'd17, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a5, 5'd30, 27'h000001bd, 5'd25, 27'h00000376, 32'h00000400,
  1'd1,  5'd6, 27'h000001de, 5'd2, 27'h000001ea, 5'd5, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000092, 5'd4, 27'h000001a3, 5'd18, 27'h000002a4, 32'h00000400,
  1'd1,  5'd9, 27'h00000093, 5'd5, 27'h0000001d, 5'd30, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000258, 5'd12, 27'h000000d0, 5'd0, 27'h0000007a, 32'h00000400,
  1'd1,  5'd5, 27'h0000037b, 5'd11, 27'h00000077, 5'd12, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034d, 5'd13, 27'h000001fb, 5'd23, 27'h0000001a, 32'h00000400,
  1'd1,  5'd8, 27'h00000381, 5'd22, 27'h0000017b, 5'd4, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000341, 5'd22, 27'h00000186, 5'd10, 27'h00000287, 32'h00000400,
  1'd1,  5'd5, 27'h00000120, 5'd25, 27'h00000255, 5'd24, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000170, 5'd1, 27'h00000378, 5'd7, 27'h0000032f, 32'h00000400,
  1'd1,  5'd18, 27'h00000019, 5'd1, 27'h000001cf, 5'd18, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000323, 5'd3, 27'h00000252, 5'd27, 27'h0000028b, 32'h00000400,
  1'd1,  5'd19, 27'h00000092, 5'd10, 27'h000002d9, 5'd5, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002be, 5'd12, 27'h000002ad, 5'd14, 27'h00000389, 32'h00000400,
  1'd1,  5'd19, 27'h00000295, 5'd13, 27'h00000039, 5'd24, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b4, 5'd23, 27'h000002aa, 5'd3, 27'h00000330, 32'h00000400,
  1'd1,  5'd19, 27'h000002b4, 5'd22, 27'h00000073, 5'd10, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b7, 5'd23, 27'h00000004, 5'd22, 27'h0000027d, 32'h00000400,
  1'd1,  5'd27, 27'h0000021c, 5'd0, 27'h00000004, 5'd2, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ee, 5'd1, 27'h00000020, 5'd13, 27'h0000022d, 32'h00000400,
  1'd1,  5'd28, 27'h0000028f, 5'd4, 27'h00000310, 5'd21, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000016, 5'd12, 27'h000000d8, 5'd0, 27'h000002ad, 32'h00000400,
  1'd1,  5'd28, 27'h00000264, 5'd14, 27'h000001aa, 5'd14, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ff, 5'd11, 27'h000001cd, 5'd23, 27'h00000100, 32'h00000400,
  1'd1,  5'd28, 27'h000002be, 5'd24, 27'h000002cc, 5'd1, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000046, 5'd23, 27'h0000004b, 5'd11, 27'h000003f2, 32'h00000400,
  1'd1,  5'd29, 27'h000002d8, 5'd22, 27'h00000224, 5'd21, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000036a, 5'd2, 27'h00000071, 5'd1, 27'h00000170, 32'h00000400,
  1'd1,  5'd6, 27'h00000352, 5'd0, 27'h00000024, 5'd10, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000016c, 5'd3, 27'h00000219, 5'd25, 27'h000000df, 32'h00000400,
  1'd1,  5'd6, 27'h00000227, 5'd12, 27'h000002cb, 5'd9, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000016, 5'd13, 27'h00000127, 5'd16, 27'h000000cd, 32'h00000400,
  1'd1,  5'd6, 27'h000003d7, 5'd10, 27'h000003c0, 5'd28, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000251, 5'd21, 27'h00000217, 5'd6, 27'h000002e9, 32'h00000400,
  1'd1,  5'd8, 27'h0000038a, 5'd24, 27'h00000294, 5'd16, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000035a, 5'd25, 27'h000001be, 5'd29, 27'h000001c7, 32'h00000400,
  1'd1,  5'd17, 27'h00000261, 5'd1, 27'h000000d2, 5'd5, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000047, 5'd3, 27'h00000345, 5'd12, 27'h000001e8, 32'h00000400,
  1'd1,  5'd19, 27'h0000025a, 5'd4, 27'h0000030d, 5'd23, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000351, 5'd10, 27'h0000037f, 5'd10, 27'h000000c9, 32'h00000400,
  1'd1,  5'd15, 27'h00000290, 5'd13, 27'h00000365, 5'd19, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039e, 5'd12, 27'h000001b1, 5'd28, 27'h0000035f, 32'h00000400,
  1'd1,  5'd19, 27'h00000193, 5'd24, 27'h000000c8, 5'd6, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b4, 5'd24, 27'h0000014e, 5'd19, 27'h0000033f, 32'h00000400,
  1'd1,  5'd19, 27'h0000034d, 5'd24, 27'h00000258, 5'd30, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002bf, 5'd1, 27'h000002c9, 5'd9, 27'h000001df, 32'h00000400,
  1'd1,  5'd30, 27'h00000025, 5'd1, 27'h0000037d, 5'd19, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000030a, 5'd2, 27'h0000020a, 5'd27, 27'h0000029f, 32'h00000400,
  1'd1,  5'd26, 27'h000000a9, 5'd10, 27'h000002e1, 5'd6, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000200, 5'd13, 27'h000000a0, 5'd16, 27'h00000040, 32'h00000400,
  1'd1,  5'd28, 27'h00000334, 5'd10, 27'h000002f0, 5'd30, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000010e, 5'd20, 27'h000003d8, 5'd5, 27'h00000316, 32'h00000400,
  1'd1,  5'd29, 27'h000001f4, 5'd22, 27'h00000015, 5'd15, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ed, 5'd22, 27'h000000e1, 5'd26, 27'h000003a3, 32'h00000400,
  1'd1,  5'd7, 27'h000000cc, 5'd7, 27'h000000e4, 5'd2, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000130, 5'd8, 27'h0000031a, 5'd13, 27'h0000008b, 32'h00000400,
  1'd1,  5'd8, 27'h00000174, 5'd7, 27'h000003c7, 5'd22, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000033c, 5'd19, 27'h000002a1, 5'd2, 27'h00000015, 32'h00000400,
  1'd1,  5'd5, 27'h00000223, 5'd18, 27'h000000a0, 5'd11, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000120, 5'd17, 27'h0000004a, 5'd22, 27'h00000090, 32'h00000400,
  1'd1,  5'd6, 27'h00000120, 5'd29, 27'h000002a0, 5'd4, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000080, 5'd27, 27'h0000001b, 5'd10, 27'h000002dd, 32'h00000400,
  1'd1,  5'd7, 27'h000003ed, 5'd29, 27'h00000132, 5'd23, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000007a, 5'd5, 27'h000003fb, 5'd3, 27'h000003ff, 32'h00000400,
  1'd1,  5'd17, 27'h00000183, 5'd6, 27'h000000c0, 5'd13, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a2, 5'd6, 27'h0000035f, 5'd22, 27'h000003cd, 32'h00000400,
  1'd1,  5'd16, 27'h000002cf, 5'd19, 27'h00000144, 5'd3, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001f4, 5'd16, 27'h00000055, 5'd14, 27'h00000339, 32'h00000400,
  1'd1,  5'd20, 27'h000000f7, 5'd20, 27'h000002a0, 5'd23, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000294, 5'd28, 27'h00000008, 5'd1, 27'h000003a6, 32'h00000400,
  1'd1,  5'd17, 27'h00000255, 5'd27, 27'h00000218, 5'd13, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000077, 5'd26, 27'h00000035, 5'd25, 27'h0000022f, 32'h00000400,
  1'd1,  5'd27, 27'h00000027, 5'd5, 27'h0000030b, 5'd2, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b6, 5'd8, 27'h000001a5, 5'd11, 27'h00000209, 32'h00000400,
  1'd1,  5'd27, 27'h000003d8, 5'd5, 27'h00000142, 5'd24, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f7, 5'd19, 27'h000000c0, 5'd2, 27'h000003ce, 32'h00000400,
  1'd1,  5'd30, 27'h00000351, 5'd18, 27'h000001b7, 5'd14, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000037, 5'd16, 27'h0000003d, 5'd24, 27'h0000011d, 32'h00000400,
  1'd1,  5'd30, 27'h00000332, 5'd28, 27'h0000008b, 5'd1, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000187, 5'd27, 27'h000000da, 5'd10, 27'h0000021c, 32'h00000400,
  1'd1,  5'd27, 27'h000002e8, 5'd27, 27'h00000335, 5'd21, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000009, 5'd6, 27'h000002c4, 5'd5, 27'h0000032c, 32'h00000400,
  1'd1,  5'd6, 27'h000003d5, 5'd6, 27'h0000024d, 5'd16, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003f8, 5'd6, 27'h000001a4, 5'd28, 27'h000003eb, 32'h00000400,
  1'd1,  5'd5, 27'h000001cf, 5'd18, 27'h000000e7, 5'd9, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000007c, 5'd16, 27'h000002b1, 5'd18, 27'h00000104, 32'h00000400,
  1'd1,  5'd10, 27'h0000010e, 5'd15, 27'h000002fc, 5'd30, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000020a, 5'd28, 27'h00000121, 5'd7, 27'h0000002f, 32'h00000400,
  1'd1,  5'd7, 27'h00000318, 5'd30, 27'h000003e8, 5'd20, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000233, 5'd26, 27'h0000029a, 5'd26, 27'h000003af, 32'h00000400,
  1'd1,  5'd16, 27'h000003c0, 5'd9, 27'h0000015b, 5'd6, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000040, 5'd10, 27'h0000001c, 5'd16, 27'h00000055, 32'h00000400,
  1'd1,  5'd16, 27'h00000371, 5'd7, 27'h00000048, 5'd28, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000356, 5'd16, 27'h00000078, 5'd9, 27'h00000303, 32'h00000400,
  1'd1,  5'd19, 27'h000002c9, 5'd15, 27'h00000286, 5'd19, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b4, 5'd18, 27'h000003cd, 5'd26, 27'h000000f2, 32'h00000400,
  1'd1,  5'd16, 27'h00000027, 5'd28, 27'h00000310, 5'd7, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000107, 5'd29, 27'h0000022f, 5'd16, 27'h00000069, 32'h00000400,
  1'd1,  5'd16, 27'h0000024e, 5'd27, 27'h0000035a, 5'd27, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000122, 5'd8, 27'h0000023f, 5'd6, 27'h000002b7, 32'h00000400,
  1'd1,  5'd26, 27'h000000cf, 5'd7, 27'h0000010d, 5'd17, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000067, 5'd5, 27'h000002f9, 5'd25, 27'h0000039a, 32'h00000400,
  1'd1,  5'd30, 27'h000002cb, 5'd19, 27'h0000027a, 5'd6, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a5, 5'd19, 27'h000003fe, 5'd16, 27'h0000003f, 32'h00000400,
  1'd1,  5'd29, 27'h00000174, 5'd19, 27'h00000203, 5'd30, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000be, 5'd27, 27'h000001f5, 5'd7, 27'h00000375, 32'h00000400,
  1'd1,  5'd30, 27'h00000185, 5'd27, 27'h00000269, 5'd16, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000358, 5'd28, 27'h0000015d, 5'd30, 27'h0000037f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h0000031e, 5'd1, 27'h00000039, 5'd1, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000a8, 5'd2, 27'h000000a5, 5'd10, 27'h0000021f, 32'h00000400,
  1'd1,  5'd3, 27'h00000031, 5'd0, 27'h0000007f, 5'd25, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000240, 5'd10, 27'h000003fb, 5'd1, 27'h00000267, 32'h00000400,
  1'd1,  5'd1, 27'h00000375, 5'd13, 27'h0000039b, 5'd12, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001b6, 5'd10, 27'h0000029e, 5'd24, 27'h000003b9, 32'h00000400,
  1'd1,  5'd4, 27'h000001ef, 5'd23, 27'h00000126, 5'd1, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000371, 5'd20, 27'h000003ed, 5'd11, 27'h00000249, 32'h00000400,
  1'd1,  5'd0, 27'h00000109, 5'd21, 27'h00000085, 5'd23, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000049, 5'd0, 27'h00000267, 5'd3, 27'h0000035c, 32'h00000400,
  1'd1,  5'd13, 27'h000002c2, 5'd4, 27'h00000188, 5'd12, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003eb, 5'd2, 27'h000003b6, 5'd21, 27'h00000324, 32'h00000400,
  1'd1,  5'd10, 27'h000002d9, 5'd13, 27'h00000365, 5'd1, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000022, 5'd13, 27'h00000069, 5'd14, 27'h0000009d, 32'h00000400,
  1'd1,  5'd11, 27'h000003fb, 5'd13, 27'h00000264, 5'd22, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000016b, 5'd25, 27'h0000030e, 5'd4, 27'h00000234, 32'h00000400,
  1'd1,  5'd11, 27'h00000159, 5'd22, 27'h000002be, 5'd10, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000135, 5'd22, 27'h00000128, 5'd20, 27'h000003c9, 32'h00000400,
  1'd1,  5'd24, 27'h00000290, 5'd3, 27'h000001b8, 5'd3, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000052, 5'd3, 27'h00000005, 5'd14, 27'h000001a3, 32'h00000400,
  1'd1,  5'd24, 27'h0000008e, 5'd4, 27'h00000304, 5'd21, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000063, 5'd13, 27'h0000024e, 5'd4, 27'h0000016e, 32'h00000400,
  1'd1,  5'd21, 27'h00000005, 5'd15, 27'h000001f9, 5'd12, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000156, 5'd12, 27'h000002d7, 5'd24, 27'h000002e5, 32'h00000400,
  1'd1,  5'd21, 27'h000003ef, 5'd24, 27'h000001e9, 5'd3, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000062, 5'd22, 27'h00000183, 5'd10, 27'h00000330, 32'h00000400,
  1'd1,  5'd25, 27'h000001f8, 5'd25, 27'h0000003d, 5'd20, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000103, 5'd3, 27'h00000331, 5'd6, 27'h0000010d, 32'h00000400,
  1'd1,  5'd3, 27'h000002cd, 5'd4, 27'h000003ce, 5'd17, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000396, 5'd4, 27'h000002c9, 5'd27, 27'h0000035d, 32'h00000400,
  1'd1,  5'd1, 27'h0000016d, 5'd14, 27'h00000098, 5'd7, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000278, 5'd12, 27'h00000009, 5'd16, 27'h00000067, 32'h00000400,
  1'd1,  5'd0, 27'h000002b0, 5'd13, 27'h00000222, 5'd27, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038a, 5'd25, 27'h00000071, 5'd8, 27'h000003bc, 32'h00000400,
  1'd1,  5'd3, 27'h000003f6, 5'd25, 27'h0000006f, 5'd18, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000198, 5'd24, 27'h000001cf, 5'd27, 27'h0000037e, 32'h00000400,
  1'd1,  5'd13, 27'h00000069, 5'd0, 27'h000002b2, 5'd5, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000233, 5'd0, 27'h000000a0, 5'd17, 27'h00000167, 32'h00000400,
  1'd1,  5'd14, 27'h0000022f, 5'd0, 27'h00000222, 5'd26, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001de, 5'd12, 27'h00000310, 5'd8, 27'h00000005, 32'h00000400,
  1'd1,  5'd13, 27'h00000061, 5'd11, 27'h00000227, 5'd18, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000e6, 5'd12, 27'h000000fe, 5'd30, 27'h0000033a, 32'h00000400,
  1'd1,  5'd13, 27'h000001a1, 5'd21, 27'h00000205, 5'd10, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000050, 5'd21, 27'h000000f8, 5'd17, 27'h000001bc, 32'h00000400,
  1'd1,  5'd12, 27'h00000067, 5'd25, 27'h00000268, 5'd30, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003c4, 5'd4, 27'h00000140, 5'd6, 27'h00000192, 32'h00000400,
  1'd1,  5'd22, 27'h000001b0, 5'd1, 27'h000002f8, 5'd18, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000033c, 5'd4, 27'h000000a9, 5'd27, 27'h000000f2, 32'h00000400,
  1'd1,  5'd22, 27'h000002ce, 5'd12, 27'h00000362, 5'd6, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000028c, 5'd14, 27'h00000371, 5'd19, 27'h00000155, 32'h00000400,
  1'd1,  5'd22, 27'h0000010b, 5'd14, 27'h0000036b, 5'd27, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000106, 5'd22, 27'h00000378, 5'd5, 27'h0000039d, 32'h00000400,
  1'd1,  5'd24, 27'h0000028b, 5'd22, 27'h00000323, 5'd19, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002e3, 5'd21, 27'h00000221, 5'd28, 27'h00000397, 32'h00000400,
  1'd1,  5'd0, 27'h00000060, 5'd8, 27'h00000281, 5'd0, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000387, 5'd7, 27'h00000384, 5'd14, 27'h00000148, 32'h00000400,
  1'd1,  5'd2, 27'h0000008d, 5'd9, 27'h00000154, 5'd24, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d3, 5'd18, 27'h000003ef, 5'd3, 27'h0000024c, 32'h00000400,
  1'd1,  5'd0, 27'h00000189, 5'd20, 27'h0000010f, 5'd13, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b0, 5'd17, 27'h000002fc, 5'd24, 27'h000001bf, 32'h00000400,
  1'd1,  5'd3, 27'h0000037c, 5'd28, 27'h000003b2, 5'd1, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000393, 5'd30, 27'h000002b3, 5'd11, 27'h000002dc, 32'h00000400,
  1'd1,  5'd4, 27'h00000177, 5'd26, 27'h000002f2, 5'd23, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001a5, 5'd9, 27'h0000004f, 5'd2, 27'h000003ee, 32'h00000400,
  1'd1,  5'd13, 27'h00000332, 5'd9, 27'h000000de, 5'd13, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000021, 5'd9, 27'h00000029, 5'd22, 27'h0000031d, 32'h00000400,
  1'd1,  5'd11, 27'h0000027b, 5'd19, 27'h000002f2, 5'd2, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003fd, 5'd18, 27'h0000013b, 5'd13, 27'h00000289, 32'h00000400,
  1'd1,  5'd14, 27'h00000175, 5'd19, 27'h0000006c, 5'd22, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000014a, 5'd30, 27'h0000029d, 5'd1, 27'h00000331, 32'h00000400,
  1'd1,  5'd11, 27'h0000014b, 5'd30, 27'h00000368, 5'd10, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e0, 5'd27, 27'h00000069, 5'd24, 27'h000000c9, 32'h00000400,
  1'd1,  5'd21, 27'h0000006b, 5'd5, 27'h000001df, 5'd0, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000219, 5'd8, 27'h0000012d, 5'd15, 27'h00000136, 32'h00000400,
  1'd1,  5'd22, 27'h000000c7, 5'd6, 27'h0000002e, 5'd21, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001d0, 5'd17, 27'h000003ea, 5'd3, 27'h00000267, 32'h00000400,
  1'd1,  5'd22, 27'h00000225, 5'd18, 27'h00000053, 5'd15, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000102, 5'd16, 27'h0000012d, 5'd22, 27'h000001d3, 32'h00000400,
  1'd1,  5'd23, 27'h00000378, 5'd25, 27'h0000038c, 5'd3, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000a0, 5'd26, 27'h000001d5, 5'd13, 27'h0000006f, 32'h00000400,
  1'd1,  5'd24, 27'h0000024d, 5'd29, 27'h0000011f, 5'd24, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000367, 5'd6, 27'h00000388, 5'd8, 27'h000000d0, 32'h00000400,
  1'd1,  5'd1, 27'h000000dd, 5'd5, 27'h00000286, 5'd18, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002c6, 5'd7, 27'h00000077, 5'd30, 27'h000001fc, 32'h00000400,
  1'd1,  5'd2, 27'h000000af, 5'd15, 27'h000002fa, 5'd5, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000043, 5'd17, 27'h00000011, 5'd19, 27'h0000034d, 32'h00000400,
  1'd1,  5'd3, 27'h0000006b, 5'd19, 27'h000000ca, 5'd30, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000021d, 5'd28, 27'h0000015d, 5'd10, 27'h00000014, 32'h00000400,
  1'd1,  5'd1, 27'h00000017, 5'd27, 27'h000001df, 5'd15, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029d, 5'd26, 27'h00000107, 5'd26, 27'h0000037e, 32'h00000400,
  1'd1,  5'd11, 27'h000002bb, 5'd9, 27'h000003a1, 5'd7, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000a3, 5'd8, 27'h0000000e, 5'd18, 27'h000002ec, 32'h00000400,
  1'd1,  5'd14, 27'h000000bd, 5'd5, 27'h000003bd, 5'd29, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d0, 5'd18, 27'h00000174, 5'd8, 27'h00000357, 32'h00000400,
  1'd1,  5'd10, 27'h00000347, 5'd16, 27'h00000281, 5'd18, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000149, 5'd19, 27'h00000368, 5'd28, 27'h0000005b, 32'h00000400,
  1'd1,  5'd10, 27'h00000200, 5'd27, 27'h0000036f, 5'd7, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f1, 5'd26, 27'h00000269, 5'd17, 27'h0000003b, 32'h00000400,
  1'd1,  5'd14, 27'h000000a9, 5'd27, 27'h00000321, 5'd30, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000035f, 5'd6, 27'h000001de, 5'd9, 27'h0000003f, 32'h00000400,
  1'd1,  5'd22, 27'h000003b3, 5'd7, 27'h0000000e, 5'd16, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000222, 5'd8, 27'h00000136, 5'd27, 27'h000001a8, 32'h00000400,
  1'd1,  5'd22, 27'h00000016, 5'd18, 27'h00000358, 5'd9, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000031, 5'd19, 27'h00000278, 5'd17, 27'h00000324, 32'h00000400,
  1'd1,  5'd22, 27'h000002f5, 5'd17, 27'h000003c8, 5'd28, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000289, 5'd29, 27'h00000131, 5'd6, 27'h000001a0, 32'h00000400,
  1'd1,  5'd24, 27'h00000302, 5'd27, 27'h0000039b, 5'd16, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000329, 5'd27, 27'h00000154, 5'd27, 27'h0000028e, 32'h00000400,
  1'd1,  5'd5, 27'h000001da, 5'd2, 27'h00000094, 5'd7, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000026a, 5'd4, 27'h000002ef, 5'd15, 27'h000003e9, 32'h00000400,
  1'd1,  5'd9, 27'h000000ee, 5'd2, 27'h00000298, 5'd27, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000020, 5'd11, 27'h000000c6, 5'd4, 27'h00000167, 32'h00000400,
  1'd1,  5'd7, 27'h00000365, 5'd11, 27'h000002b2, 5'd15, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000332, 5'd10, 27'h00000219, 5'd23, 27'h00000293, 32'h00000400,
  1'd1,  5'd8, 27'h00000270, 5'd24, 27'h00000199, 5'd0, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000197, 5'd21, 27'h000002e3, 5'd11, 27'h00000294, 32'h00000400,
  1'd1,  5'd9, 27'h00000269, 5'd25, 27'h00000193, 5'd25, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001e6, 5'd3, 27'h000002ef, 5'd5, 27'h000003c7, 32'h00000400,
  1'd1,  5'd18, 27'h000000d1, 5'd3, 27'h00000300, 5'd19, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000270, 5'd1, 27'h00000360, 5'd28, 27'h000003c1, 32'h00000400,
  1'd1,  5'd19, 27'h00000178, 5'd13, 27'h0000001a, 5'd2, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000043, 5'd14, 27'h000000c5, 5'd14, 27'h0000020e, 32'h00000400,
  1'd1,  5'd17, 27'h00000361, 5'd13, 27'h00000213, 5'd23, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000240, 5'd23, 27'h00000342, 5'd3, 27'h0000029c, 32'h00000400,
  1'd1,  5'd16, 27'h000003fe, 5'd23, 27'h000002ee, 5'd11, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000017f, 5'd25, 27'h0000026b, 5'd22, 27'h000000a2, 32'h00000400,
  1'd1,  5'd27, 27'h000003c7, 5'd2, 27'h00000128, 5'd2, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000242, 5'd3, 27'h000000cc, 5'd13, 27'h0000021d, 32'h00000400,
  1'd1,  5'd27, 27'h00000017, 5'd2, 27'h0000002d, 5'd25, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a7, 5'd15, 27'h0000018d, 5'd3, 27'h00000060, 32'h00000400,
  1'd1,  5'd29, 27'h00000273, 5'd14, 27'h000000b9, 5'd14, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001f2, 5'd13, 27'h000000c4, 5'd22, 27'h00000340, 32'h00000400,
  1'd1,  5'd25, 27'h000003f6, 5'd25, 27'h000002c6, 5'd3, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003da, 5'd22, 27'h000002f6, 5'd10, 27'h00000312, 32'h00000400,
  1'd1,  5'd29, 27'h00000269, 5'd25, 27'h0000017f, 5'd23, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000029b, 5'd0, 27'h000003b9, 5'd4, 27'h0000002b, 32'h00000400,
  1'd1,  5'd6, 27'h00000200, 5'd1, 27'h000001e0, 5'd13, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000004c, 5'd2, 27'h00000149, 5'd25, 27'h00000112, 32'h00000400,
  1'd1,  5'd10, 27'h00000072, 5'd10, 27'h000003fc, 5'd7, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a7, 5'd13, 27'h000000f5, 5'd20, 27'h00000284, 32'h00000400,
  1'd1,  5'd8, 27'h0000023f, 5'd13, 27'h00000148, 5'd27, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023d, 5'd21, 27'h000000fd, 5'd5, 27'h000003c0, 32'h00000400,
  1'd1,  5'd8, 27'h000000dd, 5'd21, 27'h000002d6, 5'd16, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a5, 5'd20, 27'h000002c2, 5'd30, 27'h00000015, 32'h00000400,
  1'd1,  5'd17, 27'h000001dd, 5'd2, 27'h00000043, 5'd2, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cb, 5'd3, 27'h0000020d, 5'd14, 27'h00000213, 32'h00000400,
  1'd1,  5'd15, 27'h00000212, 5'd3, 27'h000001ae, 5'd24, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000384, 5'd12, 27'h000002af, 5'd7, 27'h000001b8, 32'h00000400,
  1'd1,  5'd20, 27'h00000156, 5'd13, 27'h000003c9, 5'd15, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c3, 5'd11, 27'h000000b0, 5'd26, 27'h000002ea, 32'h00000400,
  1'd1,  5'd17, 27'h00000055, 5'd20, 27'h000003de, 5'd8, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000073, 5'd25, 27'h0000033f, 5'd15, 27'h000002c3, 32'h00000400,
  1'd1,  5'd17, 27'h00000153, 5'd21, 27'h00000258, 5'd29, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000037b, 5'd4, 27'h000003c2, 5'd8, 27'h000002d8, 32'h00000400,
  1'd1,  5'd28, 27'h00000235, 5'd0, 27'h000003df, 5'd18, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000018a, 5'd2, 27'h00000249, 5'd27, 27'h00000265, 32'h00000400,
  1'd1,  5'd27, 27'h00000254, 5'd13, 27'h000001a7, 5'd7, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000017f, 5'd10, 27'h00000400, 5'd20, 27'h00000223, 32'h00000400,
  1'd1,  5'd26, 27'h00000034, 5'd10, 27'h00000184, 5'd29, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a3, 5'd21, 27'h00000380, 5'd5, 27'h00000273, 32'h00000400,
  1'd1,  5'd27, 27'h00000287, 5'd23, 27'h0000002d, 5'd17, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000016e, 5'd25, 27'h00000121, 5'd29, 27'h0000038d, 32'h00000400,
  1'd1,  5'd8, 27'h000002d8, 5'd6, 27'h000002ae, 5'd1, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000c7, 5'd8, 27'h000000d3, 5'd14, 27'h000000f1, 32'h00000400,
  1'd1,  5'd7, 27'h00000103, 5'd5, 27'h0000034b, 5'd23, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000187, 5'd17, 27'h0000014e, 5'd1, 27'h00000009, 32'h00000400,
  1'd1,  5'd8, 27'h000000a8, 5'd16, 27'h00000196, 5'd15, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000113, 5'd16, 27'h00000037, 5'd24, 27'h000001c3, 32'h00000400,
  1'd1,  5'd5, 27'h000000d5, 5'd28, 27'h00000135, 5'd0, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020c, 5'd27, 27'h00000132, 5'd15, 27'h0000014f, 32'h00000400,
  1'd1,  5'd9, 27'h0000008c, 5'd28, 27'h00000169, 5'd25, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000013d, 5'd5, 27'h00000296, 5'd2, 27'h0000015c, 32'h00000400,
  1'd1,  5'd17, 27'h000003ad, 5'd6, 27'h0000003c, 5'd10, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ed, 5'd9, 27'h000001a9, 5'd23, 27'h0000031c, 32'h00000400,
  1'd1,  5'd20, 27'h000001cb, 5'd15, 27'h000003c1, 5'd1, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000026f, 5'd18, 27'h0000015b, 5'd13, 27'h00000268, 32'h00000400,
  1'd1,  5'd16, 27'h000002db, 5'd19, 27'h000003db, 5'd23, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000374, 5'd27, 27'h000003e9, 5'd0, 27'h0000016c, 32'h00000400,
  1'd1,  5'd17, 27'h00000370, 5'd27, 27'h0000000e, 5'd11, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039c, 5'd27, 27'h000001ea, 5'd21, 27'h000003f5, 32'h00000400,
  1'd1,  5'd29, 27'h0000007b, 5'd5, 27'h00000253, 5'd3, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000231, 5'd7, 27'h0000002d, 5'd15, 27'h0000014c, 32'h00000400,
  1'd1,  5'd27, 27'h000003d5, 5'd9, 27'h0000017a, 5'd25, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000024c, 5'd20, 27'h00000207, 5'd3, 27'h00000164, 32'h00000400,
  1'd1,  5'd27, 27'h00000388, 5'd17, 27'h000000f8, 5'd12, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000100, 5'd19, 27'h00000139, 5'd20, 27'h00000329, 32'h00000400,
  1'd1,  5'd27, 27'h00000339, 5'd30, 27'h000000b0, 5'd2, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000008, 5'd30, 27'h00000291, 5'd13, 27'h000003b6, 32'h00000400,
  1'd1,  5'd28, 27'h00000338, 5'd28, 27'h000002af, 5'd23, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000269, 5'd8, 27'h00000074, 5'd5, 27'h0000024d, 32'h00000400,
  1'd1,  5'd9, 27'h000002d6, 5'd8, 27'h0000008b, 5'd18, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c2, 5'd8, 27'h000002ee, 5'd29, 27'h000003c0, 32'h00000400,
  1'd1,  5'd5, 27'h000001e9, 5'd18, 27'h000001ad, 5'd6, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000247, 5'd16, 27'h00000192, 5'd19, 27'h0000008b, 32'h00000400,
  1'd1,  5'd7, 27'h000001bf, 5'd16, 27'h000003c5, 5'd28, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000006a, 5'd30, 27'h000002b7, 5'd9, 27'h00000086, 32'h00000400,
  1'd1,  5'd8, 27'h000002cc, 5'd26, 27'h000000ec, 5'd17, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002d3, 5'd26, 27'h000001f3, 5'd30, 27'h00000101, 32'h00000400,
  1'd1,  5'd20, 27'h00000013, 5'd5, 27'h00000175, 5'd6, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000134, 5'd9, 27'h00000158, 5'd20, 27'h0000004b, 32'h00000400,
  1'd1,  5'd17, 27'h00000399, 5'd5, 27'h00000393, 5'd28, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ae, 5'd17, 27'h000002c1, 5'd5, 27'h0000038a, 32'h00000400,
  1'd1,  5'd17, 27'h00000008, 5'd18, 27'h000000b1, 5'd16, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000023b, 5'd16, 27'h00000121, 5'd30, 27'h0000022c, 32'h00000400,
  1'd1,  5'd16, 27'h000000b9, 5'd26, 27'h00000358, 5'd5, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000057, 5'd29, 27'h00000221, 5'd18, 27'h00000390, 32'h00000400,
  1'd1,  5'd20, 27'h0000010b, 5'd26, 27'h000000c9, 5'd25, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000357, 5'd6, 27'h000002f0, 5'd7, 27'h000000d5, 32'h00000400,
  1'd1,  5'd29, 27'h0000009c, 5'd5, 27'h000001a0, 5'd16, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006e, 5'd7, 27'h00000114, 5'd28, 27'h00000257, 32'h00000400,
  1'd1,  5'd30, 27'h00000042, 5'd20, 27'h00000181, 5'd10, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000039f, 5'd17, 27'h000003f2, 5'd17, 27'h00000034, 32'h00000400,
  1'd1,  5'd26, 27'h00000233, 5'd15, 27'h000002e4, 5'd26, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000052, 5'd29, 27'h000002f1, 5'd5, 27'h0000026f, 32'h00000400,
  1'd1,  5'd28, 27'h00000058, 5'd29, 27'h0000008c, 5'd16, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000257, 5'd30, 27'h00000379, 5'd30, 27'h00000276, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000393, 5'd3, 27'h000000f2, 5'd2, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000241, 5'd1, 27'h000002b5, 5'd12, 27'h00000017, 32'h00000400,
  1'd1,  5'd0, 27'h00000145, 5'd4, 27'h00000359, 5'd24, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000105, 5'd12, 27'h000001e0, 5'd2, 27'h00000280, 32'h00000400,
  1'd1,  5'd1, 27'h00000354, 5'd12, 27'h0000036d, 5'd14, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000006b, 5'd13, 27'h0000029e, 5'd21, 27'h0000039d, 32'h00000400,
  1'd1,  5'd3, 27'h00000321, 5'd24, 27'h00000396, 5'd0, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000092, 5'd22, 27'h000002e5, 5'd14, 27'h0000011b, 32'h00000400,
  1'd1,  5'd4, 27'h0000031c, 5'd20, 27'h00000391, 5'd24, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e5, 5'd2, 27'h000001b0, 5'd0, 27'h00000187, 32'h00000400,
  1'd1,  5'd14, 27'h000003be, 5'd4, 27'h000000fa, 5'd10, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000185, 5'd2, 27'h0000033b, 5'd22, 27'h00000388, 32'h00000400,
  1'd1,  5'd12, 27'h0000025f, 5'd12, 27'h000003b8, 5'd2, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000188, 5'd13, 27'h0000004e, 5'd11, 27'h000002e2, 32'h00000400,
  1'd1,  5'd12, 27'h0000015d, 5'd10, 27'h00000182, 5'd22, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000388, 5'd22, 27'h000003e5, 5'd3, 27'h000002f0, 32'h00000400,
  1'd1,  5'd13, 27'h0000028f, 5'd22, 27'h000000e5, 5'd11, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c5, 5'd24, 27'h0000026f, 5'd21, 27'h0000031d, 32'h00000400,
  1'd1,  5'd25, 27'h0000013a, 5'd0, 27'h000002e9, 5'd0, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ad, 5'd1, 27'h000000eb, 5'd11, 27'h0000029e, 32'h00000400,
  1'd1,  5'd23, 27'h00000011, 5'd1, 27'h000002ea, 5'd24, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000374, 5'd12, 27'h000002a5, 5'd4, 27'h00000379, 32'h00000400,
  1'd1,  5'd22, 27'h00000132, 5'd15, 27'h000001bf, 5'd13, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000264, 5'd15, 27'h00000191, 5'd21, 27'h00000388, 32'h00000400,
  1'd1,  5'd22, 27'h0000033f, 5'd20, 27'h000002fa, 5'd0, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c8, 5'd22, 27'h00000113, 5'd11, 27'h000001ce, 32'h00000400,
  1'd1,  5'd24, 27'h00000012, 5'd24, 27'h0000032f, 5'd24, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005c, 5'd1, 27'h0000037a, 5'd8, 27'h00000360, 32'h00000400,
  1'd1,  5'd2, 27'h00000362, 5'd3, 27'h000000f0, 5'd20, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000010a, 5'd3, 27'h000000d0, 5'd29, 27'h000000f2, 32'h00000400,
  1'd1,  5'd4, 27'h000000d7, 5'd11, 27'h000001e2, 5'd9, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c3, 5'd11, 27'h0000011e, 5'd16, 27'h000002f3, 32'h00000400,
  1'd1,  5'd0, 27'h000002c1, 5'd14, 27'h0000027f, 5'd28, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001d9, 5'd25, 27'h00000069, 5'd6, 27'h000000d1, 32'h00000400,
  1'd1,  5'd1, 27'h00000141, 5'd22, 27'h000003a9, 5'd18, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000315, 5'd20, 27'h00000358, 5'd26, 27'h000003cc, 32'h00000400,
  1'd1,  5'd13, 27'h000002ec, 5'd3, 27'h000000f3, 5'd10, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000203, 5'd3, 27'h0000016f, 5'd19, 27'h000001f1, 32'h00000400,
  1'd1,  5'd11, 27'h00000028, 5'd3, 27'h00000130, 5'd28, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000031b, 5'd12, 27'h0000025b, 5'd7, 27'h0000024f, 32'h00000400,
  1'd1,  5'd14, 27'h00000278, 5'd12, 27'h00000256, 5'd20, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000071, 5'd11, 27'h0000014e, 5'd30, 27'h000001c1, 32'h00000400,
  1'd1,  5'd12, 27'h00000314, 5'd23, 27'h0000011b, 5'd8, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000e6, 5'd25, 27'h0000016c, 5'd18, 27'h00000164, 32'h00000400,
  1'd1,  5'd13, 27'h000001e5, 5'd22, 27'h0000032a, 5'd30, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002f1, 5'd2, 27'h000000d0, 5'd5, 27'h00000392, 32'h00000400,
  1'd1,  5'd21, 27'h00000113, 5'd3, 27'h00000374, 5'd18, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000010e, 5'd4, 27'h0000012b, 5'd27, 27'h0000037d, 32'h00000400,
  1'd1,  5'd24, 27'h00000177, 5'd12, 27'h000000f6, 5'd6, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000354, 5'd11, 27'h00000131, 5'd15, 27'h000002c8, 32'h00000400,
  1'd1,  5'd23, 27'h0000022b, 5'd11, 27'h0000025d, 5'd28, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000051, 5'd22, 27'h0000014f, 5'd6, 27'h0000039d, 32'h00000400,
  1'd1,  5'd23, 27'h00000103, 5'd23, 27'h00000358, 5'd18, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000164, 5'd23, 27'h0000028f, 5'd25, 27'h00000373, 32'h00000400,
  1'd1,  5'd3, 27'h0000027b, 5'd7, 27'h0000017b, 5'd1, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c3, 5'd10, 27'h00000131, 5'd13, 27'h000002ef, 32'h00000400,
  1'd1,  5'd3, 27'h000002a9, 5'd6, 27'h0000007c, 5'd24, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000028, 5'd15, 27'h000002ff, 5'd4, 27'h00000154, 32'h00000400,
  1'd1,  5'd5, 27'h0000008f, 5'd19, 27'h000003d9, 5'd12, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001db, 5'd16, 27'h00000124, 5'd23, 27'h000000e6, 32'h00000400,
  1'd1,  5'd5, 27'h00000068, 5'd27, 27'h00000161, 5'd4, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001ea, 5'd29, 27'h000000ff, 5'd13, 27'h00000124, 32'h00000400,
  1'd1,  5'd1, 27'h0000006d, 5'd28, 27'h00000359, 5'd24, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000359, 5'd5, 27'h0000029b, 5'd1, 27'h0000008e, 32'h00000400,
  1'd1,  5'd12, 27'h0000030a, 5'd5, 27'h0000036b, 5'd13, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001af, 5'd6, 27'h00000287, 5'd25, 27'h000000ca, 32'h00000400,
  1'd1,  5'd15, 27'h00000125, 5'd16, 27'h000002d4, 5'd2, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000215, 5'd16, 27'h00000203, 5'd11, 27'h000000e2, 32'h00000400,
  1'd1,  5'd14, 27'h000001b1, 5'd17, 27'h0000019e, 5'd21, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000012d, 5'd25, 27'h0000037e, 5'd3, 27'h00000393, 32'h00000400,
  1'd1,  5'd15, 27'h0000004f, 5'd29, 27'h00000190, 5'd13, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000034d, 5'd28, 27'h00000020, 5'd21, 27'h00000365, 32'h00000400,
  1'd1,  5'd21, 27'h000003e3, 5'd8, 27'h0000030e, 5'd2, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000066, 5'd9, 27'h00000082, 5'd11, 27'h000002fe, 32'h00000400,
  1'd1,  5'd22, 27'h0000037d, 5'd7, 27'h000000d7, 5'd24, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002dd, 5'd19, 27'h000001aa, 5'd2, 27'h0000039a, 32'h00000400,
  1'd1,  5'd20, 27'h00000344, 5'd19, 27'h00000226, 5'd11, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000081, 5'd20, 27'h000001a7, 5'd24, 27'h000001cd, 32'h00000400,
  1'd1,  5'd25, 27'h000000d2, 5'd28, 27'h00000110, 5'd4, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000036e, 5'd26, 27'h00000195, 5'd13, 27'h000000d4, 32'h00000400,
  1'd1,  5'd21, 27'h00000106, 5'd25, 27'h0000038f, 5'd25, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ce, 5'd6, 27'h00000154, 5'd5, 27'h000002c0, 32'h00000400,
  1'd1,  5'd2, 27'h00000186, 5'd9, 27'h00000372, 5'd19, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000120, 5'd7, 27'h0000020d, 5'd27, 27'h000002ac, 32'h00000400,
  1'd1,  5'd1, 27'h000002c8, 5'd18, 27'h00000339, 5'd9, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000023f, 5'd17, 27'h000003bb, 5'd20, 27'h000000ab, 32'h00000400,
  1'd1,  5'd0, 27'h0000013f, 5'd18, 27'h00000261, 5'd27, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000119, 5'd30, 27'h000000a8, 5'd9, 27'h0000016e, 32'h00000400,
  1'd1,  5'd3, 27'h000003cf, 5'd27, 27'h0000015c, 5'd17, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002fb, 5'd30, 27'h00000342, 5'd27, 27'h0000006e, 32'h00000400,
  1'd1,  5'd11, 27'h000000fb, 5'd10, 27'h000000d3, 5'd6, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001d3, 5'd5, 27'h00000222, 5'd15, 27'h000002ca, 32'h00000400,
  1'd1,  5'd12, 27'h00000275, 5'd9, 27'h00000046, 5'd26, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000290, 5'd20, 27'h00000112, 5'd10, 27'h000000ed, 32'h00000400,
  1'd1,  5'd10, 27'h00000286, 5'd17, 27'h00000099, 5'd20, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000073, 5'd15, 27'h00000202, 5'd30, 27'h00000267, 32'h00000400,
  1'd1,  5'd10, 27'h0000028f, 5'd27, 27'h0000026a, 5'd8, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000009c, 5'd30, 27'h0000031b, 5'd16, 27'h000001ae, 32'h00000400,
  1'd1,  5'd11, 27'h0000012e, 5'd27, 27'h0000011d, 5'd26, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000273, 5'd9, 27'h000001b9, 5'd5, 27'h0000025f, 32'h00000400,
  1'd1,  5'd22, 27'h000003ec, 5'd8, 27'h000000d9, 5'd16, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000292, 5'd9, 27'h000000c5, 5'd29, 27'h000000a0, 32'h00000400,
  1'd1,  5'd23, 27'h00000146, 5'd18, 27'h00000168, 5'd8, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000243, 5'd19, 27'h000000f4, 5'd16, 27'h000000e4, 32'h00000400,
  1'd1,  5'd21, 27'h0000038a, 5'd19, 27'h000001c8, 5'd29, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000034b, 5'd30, 27'h00000172, 5'd9, 27'h000001d9, 32'h00000400,
  1'd1,  5'd25, 27'h00000203, 5'd26, 27'h00000201, 5'd18, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000142, 5'd29, 27'h0000036d, 5'd26, 27'h0000001e, 32'h00000400,
  1'd1,  5'd7, 27'h000001c6, 5'd4, 27'h00000082, 5'd5, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000150, 5'd2, 27'h000002e2, 5'd19, 27'h000000a6, 32'h00000400,
  1'd1,  5'd5, 27'h00000295, 5'd0, 27'h00000218, 5'd26, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001b4, 5'd14, 27'h000003f2, 5'd1, 27'h00000275, 32'h00000400,
  1'd1,  5'd8, 27'h00000251, 5'd11, 27'h00000362, 5'd15, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000255, 5'd13, 27'h0000019d, 5'd24, 27'h000002ff, 32'h00000400,
  1'd1,  5'd5, 27'h000000ee, 5'd24, 27'h0000038d, 5'd3, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000020, 5'd21, 27'h0000037b, 5'd13, 27'h0000024b, 32'h00000400,
  1'd1,  5'd8, 27'h000002fa, 5'd23, 27'h00000353, 5'd24, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035a, 5'd0, 27'h000000a4, 5'd6, 27'h000001fe, 32'h00000400,
  1'd1,  5'd17, 27'h00000071, 5'd1, 27'h000003a7, 5'd16, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000037, 5'd3, 27'h000001b4, 5'd29, 27'h00000270, 32'h00000400,
  1'd1,  5'd19, 27'h0000006c, 5'd13, 27'h000002ce, 5'd1, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b6, 5'd12, 27'h000001c1, 5'd10, 27'h000001c9, 32'h00000400,
  1'd1,  5'd15, 27'h000003df, 5'd14, 27'h00000162, 5'd25, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001f7, 5'd23, 27'h00000302, 5'd2, 27'h000003ae, 32'h00000400,
  1'd1,  5'd18, 27'h0000023f, 5'd24, 27'h0000002f, 5'd13, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000074, 5'd22, 27'h000001c1, 5'd25, 27'h000000b9, 32'h00000400,
  1'd1,  5'd26, 27'h00000170, 5'd1, 27'h00000256, 5'd2, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000e, 5'd2, 27'h00000124, 5'd13, 27'h0000010f, 32'h00000400,
  1'd1,  5'd26, 27'h000002c6, 5'd1, 27'h000003f0, 5'd21, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000289, 5'd14, 27'h00000003, 5'd0, 27'h0000020c, 32'h00000400,
  1'd1,  5'd26, 27'h0000039e, 5'd14, 27'h000002ac, 5'd14, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000039b, 5'd15, 27'h00000010, 5'd22, 27'h0000017d, 32'h00000400,
  1'd1,  5'd30, 27'h00000229, 5'd24, 27'h000002f8, 5'd3, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f8, 5'd24, 27'h0000037c, 5'd11, 27'h000003e9, 32'h00000400,
  1'd1,  5'd29, 27'h00000213, 5'd25, 27'h00000206, 5'd21, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000173, 5'd3, 27'h000002da, 5'd4, 27'h00000051, 32'h00000400,
  1'd1,  5'd5, 27'h000001bc, 5'd3, 27'h0000012a, 5'd14, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001cd, 5'd4, 27'h000001bd, 5'd24, 27'h00000075, 32'h00000400,
  1'd1,  5'd9, 27'h00000036, 5'd14, 27'h000002d7, 5'd7, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000116, 5'd10, 27'h00000220, 5'd18, 27'h000003cb, 32'h00000400,
  1'd1,  5'd8, 27'h000003ba, 5'd14, 27'h00000163, 5'd29, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000031e, 5'd25, 27'h000001bd, 5'd5, 27'h0000029d, 32'h00000400,
  1'd1,  5'd6, 27'h00000080, 5'd21, 27'h0000027a, 5'd16, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002a9, 5'd24, 27'h000003f3, 5'd26, 27'h000000fa, 32'h00000400,
  1'd1,  5'd17, 27'h000003d2, 5'd2, 27'h00000306, 5'd3, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000246, 5'd4, 27'h00000169, 5'd13, 27'h00000072, 32'h00000400,
  1'd1,  5'd16, 27'h000003ba, 5'd0, 27'h000003ad, 5'd22, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000009b, 5'd15, 27'h00000140, 5'd9, 27'h00000100, 32'h00000400,
  1'd1,  5'd18, 27'h0000012f, 5'd14, 27'h00000174, 5'd17, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000016f, 5'd11, 27'h000002cf, 5'd28, 27'h00000207, 32'h00000400,
  1'd1,  5'd17, 27'h000000be, 5'd25, 27'h00000143, 5'd8, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000076, 5'd23, 27'h00000012, 5'd19, 27'h000001d6, 32'h00000400,
  1'd1,  5'd17, 27'h000003d7, 5'd25, 27'h0000000b, 5'd28, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000005f, 5'd2, 27'h00000295, 5'd7, 27'h000000e0, 32'h00000400,
  1'd1,  5'd28, 27'h0000038e, 5'd5, 27'h00000047, 5'd17, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000021, 5'd4, 27'h00000265, 5'd26, 27'h000001ca, 32'h00000400,
  1'd1,  5'd27, 27'h000002a8, 5'd13, 27'h000001af, 5'd6, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000288, 5'd11, 27'h0000002f, 5'd15, 27'h000003ba, 32'h00000400,
  1'd1,  5'd28, 27'h000003cf, 5'd15, 27'h00000189, 5'd26, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000157, 5'd21, 27'h00000326, 5'd8, 27'h0000003d, 32'h00000400,
  1'd1,  5'd26, 27'h00000347, 5'd23, 27'h0000008b, 5'd16, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000228, 5'd23, 27'h0000014d, 5'd30, 27'h00000381, 32'h00000400,
  1'd1,  5'd7, 27'h00000036, 5'd8, 27'h00000101, 5'd0, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ad, 5'd5, 27'h000001b7, 5'd13, 27'h000003be, 32'h00000400,
  1'd1,  5'd7, 27'h0000039a, 5'd6, 27'h000002c2, 5'd21, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000000b, 5'd15, 27'h0000034d, 5'd4, 27'h00000313, 32'h00000400,
  1'd1,  5'd9, 27'h00000369, 5'd17, 27'h0000001d, 5'd11, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007c, 5'd16, 27'h000002fd, 5'd25, 27'h00000117, 32'h00000400,
  1'd1,  5'd7, 27'h000000c0, 5'd27, 27'h00000221, 5'd1, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000359, 5'd26, 27'h000003a9, 5'd12, 27'h0000037d, 32'h00000400,
  1'd1,  5'd5, 27'h0000031f, 5'd27, 27'h00000386, 5'd21, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000285, 5'd10, 27'h0000002c, 5'd1, 27'h00000324, 32'h00000400,
  1'd1,  5'd19, 27'h000003c3, 5'd9, 27'h0000000f, 5'd13, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000017b, 5'd6, 27'h000002d3, 5'd23, 27'h00000093, 32'h00000400,
  1'd1,  5'd18, 27'h000000df, 5'd16, 27'h000000b5, 5'd1, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000012e, 5'd19, 27'h0000026c, 5'd10, 27'h00000216, 32'h00000400,
  1'd1,  5'd15, 27'h00000359, 5'd18, 27'h0000004c, 5'd21, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000207, 5'd27, 27'h00000327, 5'd2, 27'h000000e0, 32'h00000400,
  1'd1,  5'd16, 27'h000000a4, 5'd26, 27'h000000a4, 5'd15, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000085, 5'd28, 27'h00000339, 5'd21, 27'h00000268, 32'h00000400,
  1'd1,  5'd27, 27'h00000046, 5'd5, 27'h00000243, 5'd2, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a7, 5'd8, 27'h000000e8, 5'd15, 27'h000000ee, 32'h00000400,
  1'd1,  5'd30, 27'h0000024b, 5'd7, 27'h0000016d, 5'd20, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001f4, 5'd19, 27'h0000023c, 5'd4, 27'h000001b6, 32'h00000400,
  1'd1,  5'd28, 27'h000003cf, 5'd18, 27'h000002b2, 5'd10, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000014, 5'd20, 27'h000000c3, 5'd21, 27'h00000326, 32'h00000400,
  1'd1,  5'd30, 27'h0000039e, 5'd29, 27'h0000039c, 5'd0, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000378, 5'd27, 27'h000002c1, 5'd11, 27'h00000091, 32'h00000400,
  1'd1,  5'd27, 27'h00000320, 5'd30, 27'h00000338, 5'd24, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013d, 5'd5, 27'h000002f6, 5'd6, 27'h000001ed, 32'h00000400,
  1'd1,  5'd6, 27'h00000184, 5'd7, 27'h00000100, 5'd18, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000039b, 5'd10, 27'h000000fc, 5'd30, 27'h00000236, 32'h00000400,
  1'd1,  5'd8, 27'h000000e6, 5'd16, 27'h00000345, 5'd7, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000015e, 5'd20, 27'h0000025d, 5'd18, 27'h000001dc, 32'h00000400,
  1'd1,  5'd5, 27'h0000010f, 5'd19, 27'h000003a0, 5'd26, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000003e, 5'd26, 27'h000002f1, 5'd8, 27'h00000191, 32'h00000400,
  1'd1,  5'd9, 27'h0000008e, 5'd28, 27'h000003ff, 5'd16, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003b6, 5'd29, 27'h000001bf, 5'd30, 27'h0000026d, 32'h00000400,
  1'd1,  5'd18, 27'h000003c8, 5'd9, 27'h000001c5, 5'd10, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000183, 5'd5, 27'h000000c3, 5'd19, 27'h00000352, 32'h00000400,
  1'd1,  5'd15, 27'h00000206, 5'd9, 27'h00000080, 5'd29, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000016e, 5'd18, 27'h000002d0, 5'd8, 27'h000001f4, 32'h00000400,
  1'd1,  5'd16, 27'h000001dc, 5'd20, 27'h0000004b, 5'd16, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000012a, 5'd17, 27'h000003e2, 5'd30, 27'h000003dd, 32'h00000400,
  1'd1,  5'd15, 27'h0000034f, 5'd29, 27'h00000126, 5'd8, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000008f, 5'd29, 27'h000001bf, 5'd20, 27'h0000017f, 32'h00000400,
  1'd1,  5'd20, 27'h0000010c, 5'd29, 27'h000001cb, 5'd28, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a1, 5'd8, 27'h00000119, 5'd8, 27'h00000003, 32'h00000400,
  1'd1,  5'd26, 27'h000001ae, 5'd9, 27'h000001f3, 5'd20, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c1, 5'd6, 27'h0000001f, 5'd29, 27'h000003e8, 32'h00000400,
  1'd1,  5'd26, 27'h00000180, 5'd18, 27'h0000035f, 5'd10, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ca, 5'd16, 27'h00000022, 5'd19, 27'h00000384, 32'h00000400,
  1'd1,  5'd29, 27'h00000321, 5'd18, 27'h000001f6, 5'd30, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001bd, 5'd26, 27'h00000003, 5'd8, 27'h000001db, 32'h00000400,
  1'd1,  5'd28, 27'h0000021e, 5'd26, 27'h0000003a, 5'd19, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000262, 5'd30, 27'h0000003e, 5'd29, 27'h000001f7, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000001a7, 5'd0, 27'h00000307, 5'd4, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d0, 5'd5, 27'h00000037, 5'd12, 27'h0000025d, 32'h00000400,
  1'd1,  5'd2, 27'h00000065, 5'd0, 27'h000000ac, 5'd24, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039b, 5'd13, 27'h000001c1, 5'd3, 27'h000000de, 32'h00000400,
  1'd1,  5'd0, 27'h000001d2, 5'd13, 27'h00000137, 5'd14, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d5, 5'd10, 27'h00000313, 5'd20, 27'h000003a5, 32'h00000400,
  1'd1,  5'd2, 27'h00000182, 5'd22, 27'h0000002a, 5'd4, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002bc, 5'd25, 27'h000001b1, 5'd12, 27'h000001a4, 32'h00000400,
  1'd1,  5'd3, 27'h00000005, 5'd21, 27'h000002e8, 5'd24, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a9, 5'd3, 27'h00000262, 5'd2, 27'h00000398, 32'h00000400,
  1'd1,  5'd15, 27'h00000001, 5'd1, 27'h00000387, 5'd14, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000031d, 5'd0, 27'h0000039a, 5'd22, 27'h000003e9, 32'h00000400,
  1'd1,  5'd12, 27'h00000218, 5'd15, 27'h00000018, 5'd5, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000368, 5'd11, 27'h0000015c, 5'd15, 27'h000001e3, 32'h00000400,
  1'd1,  5'd12, 27'h00000342, 5'd13, 27'h00000008, 5'd23, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c4, 5'd23, 27'h00000193, 5'd1, 27'h0000011e, 32'h00000400,
  1'd1,  5'd11, 27'h000003ba, 5'd22, 27'h00000217, 5'd12, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038e, 5'd24, 27'h00000397, 5'd25, 27'h000000f7, 32'h00000400,
  1'd1,  5'd23, 27'h00000302, 5'd3, 27'h000003e3, 5'd1, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000159, 5'd3, 27'h00000030, 5'd12, 27'h00000299, 32'h00000400,
  1'd1,  5'd21, 27'h00000022, 5'd0, 27'h0000005c, 5'd25, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000004c, 5'd12, 27'h0000004b, 5'd4, 27'h0000016e, 32'h00000400,
  1'd1,  5'd22, 27'h0000026b, 5'd13, 27'h00000052, 5'd11, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002f0, 5'd11, 27'h00000156, 5'd23, 27'h000002c2, 32'h00000400,
  1'd1,  5'd22, 27'h00000160, 5'd24, 27'h00000371, 5'd2, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ff, 5'd22, 27'h0000028c, 5'd14, 27'h000001e6, 32'h00000400,
  1'd1,  5'd23, 27'h00000286, 5'd22, 27'h0000000c, 5'd22, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000121, 5'd3, 27'h0000020c, 5'd9, 27'h0000036d, 32'h00000400,
  1'd1,  5'd2, 27'h00000070, 5'd1, 27'h0000018a, 5'd17, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001aa, 5'd2, 27'h00000252, 5'd30, 27'h000001c4, 32'h00000400,
  1'd1,  5'd5, 27'h00000028, 5'd11, 27'h000002c9, 5'd6, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ee, 5'd12, 27'h00000389, 5'd16, 27'h0000026a, 32'h00000400,
  1'd1,  5'd0, 27'h000000c3, 5'd11, 27'h00000191, 5'd29, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ea, 5'd24, 27'h0000010c, 5'd9, 27'h000002aa, 32'h00000400,
  1'd1,  5'd0, 27'h000003e7, 5'd24, 27'h000001de, 5'd17, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014a, 5'd24, 27'h000003d0, 5'd30, 27'h00000144, 32'h00000400,
  1'd1,  5'd10, 27'h000002b3, 5'd3, 27'h0000014a, 5'd9, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000246, 5'd5, 27'h0000007d, 5'd19, 27'h000001ee, 32'h00000400,
  1'd1,  5'd15, 27'h000000ab, 5'd2, 27'h00000146, 5'd30, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000045, 5'd11, 27'h0000030e, 5'd8, 27'h000003b5, 32'h00000400,
  1'd1,  5'd14, 27'h00000106, 5'd14, 27'h000000c1, 5'd17, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fe, 5'd11, 27'h000003ff, 5'd25, 27'h0000036f, 32'h00000400,
  1'd1,  5'd10, 27'h00000386, 5'd24, 27'h000002c4, 5'd8, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e6, 5'd20, 27'h00000310, 5'd18, 27'h00000059, 32'h00000400,
  1'd1,  5'd11, 27'h000002e6, 5'd24, 27'h00000253, 5'd30, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000347, 5'd1, 27'h00000298, 5'd10, 27'h0000008b, 32'h00000400,
  1'd1,  5'd20, 27'h00000390, 5'd3, 27'h000000d4, 5'd20, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000025a, 5'd4, 27'h000003dc, 5'd28, 27'h000002b8, 32'h00000400,
  1'd1,  5'd23, 27'h0000039d, 5'd10, 27'h00000276, 5'd8, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c1, 5'd12, 27'h0000014c, 5'd19, 27'h000000dd, 32'h00000400,
  1'd1,  5'd21, 27'h000002ba, 5'd13, 27'h00000065, 5'd28, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000005d, 5'd24, 27'h0000004d, 5'd7, 27'h0000022d, 32'h00000400,
  1'd1,  5'd25, 27'h00000307, 5'd25, 27'h00000061, 5'd18, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000140, 5'd24, 27'h000002b6, 5'd27, 27'h00000356, 32'h00000400,
  1'd1,  5'd3, 27'h00000192, 5'd9, 27'h000001bf, 5'd2, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032c, 5'd5, 27'h000002be, 5'd11, 27'h000003ca, 32'h00000400,
  1'd1,  5'd2, 27'h000002e3, 5'd6, 27'h00000105, 5'd20, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000021a, 5'd18, 27'h0000020e, 5'd4, 27'h000000e3, 32'h00000400,
  1'd1,  5'd3, 27'h0000015c, 5'd18, 27'h000000be, 5'd13, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000153, 5'd19, 27'h000002f2, 5'd21, 27'h0000028e, 32'h00000400,
  1'd1,  5'd4, 27'h00000388, 5'd30, 27'h000000c0, 5'd0, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000009, 5'd27, 27'h0000034b, 5'd13, 27'h0000036b, 32'h00000400,
  1'd1,  5'd4, 27'h00000353, 5'd26, 27'h000003d7, 5'd23, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000122, 5'd6, 27'h000002bf, 5'd4, 27'h00000227, 32'h00000400,
  1'd1,  5'd10, 27'h0000017c, 5'd8, 27'h000003aa, 5'd14, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000287, 5'd9, 27'h00000129, 5'd21, 27'h00000374, 32'h00000400,
  1'd1,  5'd12, 27'h000001cb, 5'd20, 27'h000000a4, 5'd3, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000025c, 5'd17, 27'h00000143, 5'd14, 27'h000000ee, 32'h00000400,
  1'd1,  5'd12, 27'h00000101, 5'd17, 27'h000000b0, 5'd22, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000fd, 5'd28, 27'h0000024b, 5'd4, 27'h00000156, 32'h00000400,
  1'd1,  5'd14, 27'h0000003f, 5'd26, 27'h00000364, 5'd14, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000038c, 5'd29, 27'h00000318, 5'd21, 27'h0000021f, 32'h00000400,
  1'd1,  5'd22, 27'h00000177, 5'd8, 27'h00000062, 5'd1, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f0, 5'd6, 27'h000002af, 5'd15, 27'h00000172, 32'h00000400,
  1'd1,  5'd23, 27'h000000bd, 5'd5, 27'h0000018c, 5'd22, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a0, 5'd15, 27'h000003fa, 5'd2, 27'h0000010e, 32'h00000400,
  1'd1,  5'd22, 27'h00000211, 5'd19, 27'h000001a9, 5'd11, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000185, 5'd19, 27'h000003f5, 5'd21, 27'h00000004, 32'h00000400,
  1'd1,  5'd22, 27'h000002b3, 5'd26, 27'h00000238, 5'd0, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b9, 5'd30, 27'h0000011d, 5'd13, 27'h00000355, 32'h00000400,
  1'd1,  5'd23, 27'h000001f5, 5'd29, 27'h000003e6, 5'd22, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000170, 5'd9, 27'h00000010, 5'd6, 27'h00000063, 32'h00000400,
  1'd1,  5'd0, 27'h00000065, 5'd8, 27'h000003a8, 5'd19, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000207, 5'd5, 27'h0000039d, 5'd26, 27'h000000a6, 32'h00000400,
  1'd1,  5'd0, 27'h0000012d, 5'd19, 27'h000001dc, 5'd10, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001a8, 5'd19, 27'h00000058, 5'd18, 27'h000001da, 32'h00000400,
  1'd1,  5'd1, 27'h0000012f, 5'd17, 27'h00000081, 5'd30, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000009f, 5'd28, 27'h000003ba, 5'd7, 27'h00000133, 32'h00000400,
  1'd1,  5'd1, 27'h0000033b, 5'd29, 27'h00000140, 5'd16, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000235, 5'd30, 27'h000003d9, 5'd26, 27'h000002e9, 32'h00000400,
  1'd1,  5'd11, 27'h00000260, 5'd5, 27'h000001e7, 5'd7, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d5, 5'd6, 27'h00000028, 5'd17, 27'h00000133, 32'h00000400,
  1'd1,  5'd14, 27'h000000c3, 5'd8, 27'h000000ee, 5'd29, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c2, 5'd16, 27'h000002ce, 5'd8, 27'h00000366, 32'h00000400,
  1'd1,  5'd14, 27'h00000048, 5'd17, 27'h00000309, 5'd19, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000099, 5'd20, 27'h00000152, 5'd27, 27'h00000338, 32'h00000400,
  1'd1,  5'd13, 27'h00000375, 5'd30, 27'h000000aa, 5'd5, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e2, 5'd27, 27'h0000009d, 5'd17, 27'h000003f7, 32'h00000400,
  1'd1,  5'd12, 27'h000000c8, 5'd29, 27'h000001cd, 5'd30, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001cc, 5'd9, 27'h00000275, 5'd6, 27'h0000004c, 32'h00000400,
  1'd1,  5'd22, 27'h000002c2, 5'd5, 27'h0000025f, 5'd18, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000154, 5'd8, 27'h00000267, 5'd28, 27'h000000c5, 32'h00000400,
  1'd1,  5'd21, 27'h00000171, 5'd18, 27'h000003f0, 5'd9, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000030b, 5'd16, 27'h000002d7, 5'd17, 27'h00000191, 32'h00000400,
  1'd1,  5'd22, 27'h000001c4, 5'd16, 27'h000003d5, 5'd28, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000016e, 5'd27, 27'h000003c5, 5'd9, 27'h0000000d, 32'h00000400,
  1'd1,  5'd23, 27'h000003be, 5'd27, 27'h000001a3, 5'd16, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e9, 5'd28, 27'h0000026f, 5'd30, 27'h00000107, 32'h00000400,
  1'd1,  5'd9, 27'h000002bc, 5'd4, 27'h0000029a, 5'd7, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000322, 5'd2, 27'h00000108, 5'd16, 27'h00000266, 32'h00000400,
  1'd1,  5'd5, 27'h00000107, 5'd1, 27'h0000015a, 5'd28, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000044, 5'd15, 27'h000001d7, 5'd2, 27'h000003b7, 32'h00000400,
  1'd1,  5'd7, 27'h00000143, 5'd12, 27'h00000072, 5'd11, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002c5, 5'd12, 27'h000003bd, 5'd21, 27'h00000325, 32'h00000400,
  1'd1,  5'd10, 27'h000000c8, 5'd22, 27'h0000002c, 5'd2, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000378, 5'd21, 27'h000002c1, 5'd13, 27'h000002cc, 32'h00000400,
  1'd1,  5'd9, 27'h0000024b, 5'd20, 27'h0000039b, 5'd22, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003ef, 5'd2, 27'h0000015d, 5'd8, 27'h0000039b, 32'h00000400,
  1'd1,  5'd17, 27'h00000005, 5'd2, 27'h0000026c, 5'd20, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000023, 5'd0, 27'h00000292, 5'd27, 27'h0000022e, 32'h00000400,
  1'd1,  5'd16, 27'h000002e3, 5'd15, 27'h00000111, 5'd2, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ee, 5'd11, 27'h0000001c, 5'd11, 27'h000001dc, 32'h00000400,
  1'd1,  5'd18, 27'h00000251, 5'd11, 27'h0000024d, 5'd25, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003fe, 5'd23, 27'h000001ce, 5'd2, 27'h00000032, 32'h00000400,
  1'd1,  5'd19, 27'h00000019, 5'd21, 27'h0000009f, 5'd12, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a9, 5'd24, 27'h00000278, 5'd22, 27'h000000fa, 32'h00000400,
  1'd1,  5'd28, 27'h000003e3, 5'd4, 27'h000003cc, 5'd4, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001b5, 5'd3, 27'h000000ae, 5'd13, 27'h0000008a, 32'h00000400,
  1'd1,  5'd30, 27'h0000011e, 5'd4, 27'h00000156, 5'd22, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001c3, 5'd13, 27'h000003b0, 5'd3, 27'h0000007f, 32'h00000400,
  1'd1,  5'd30, 27'h00000333, 5'd13, 27'h00000128, 5'd11, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000016f, 5'd13, 27'h000001a3, 5'd23, 27'h00000215, 32'h00000400,
  1'd1,  5'd29, 27'h0000000a, 5'd23, 27'h0000027c, 5'd4, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000dc, 5'd20, 27'h00000337, 5'd12, 27'h00000097, 32'h00000400,
  1'd1,  5'd27, 27'h0000022e, 5'd23, 27'h0000003f, 5'd23, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002d8, 5'd0, 27'h000000a1, 5'd3, 27'h00000106, 32'h00000400,
  1'd1,  5'd7, 27'h0000011b, 5'd4, 27'h00000082, 5'd14, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000126, 5'd0, 27'h000003d3, 5'd22, 27'h00000359, 32'h00000400,
  1'd1,  5'd8, 27'h000000cc, 5'd11, 27'h000002e8, 5'd6, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000383, 5'd12, 27'h00000328, 5'd17, 27'h0000011c, 32'h00000400,
  1'd1,  5'd8, 27'h0000019d, 5'd12, 27'h0000011b, 5'd30, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000005f, 5'd22, 27'h00000183, 5'd8, 27'h00000004, 32'h00000400,
  1'd1,  5'd6, 27'h000001d1, 5'd24, 27'h000000c1, 5'd18, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000301, 5'd22, 27'h00000310, 5'd28, 27'h000003d7, 32'h00000400,
  1'd1,  5'd18, 27'h000000d2, 5'd1, 27'h000000bc, 5'd1, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000123, 5'd1, 27'h00000388, 5'd10, 27'h000001ea, 32'h00000400,
  1'd1,  5'd17, 27'h000002b2, 5'd2, 27'h000001b4, 5'd21, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e6, 5'd12, 27'h0000026c, 5'd6, 27'h00000317, 32'h00000400,
  1'd1,  5'd19, 27'h000002ff, 5'd15, 27'h00000172, 5'd19, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000034f, 5'd14, 27'h000001a8, 5'd28, 27'h000001d6, 32'h00000400,
  1'd1,  5'd19, 27'h0000001f, 5'd23, 27'h00000162, 5'd9, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003f4, 5'd24, 27'h00000123, 5'd19, 27'h000001f3, 32'h00000400,
  1'd1,  5'd15, 27'h00000332, 5'd24, 27'h0000024a, 5'd30, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000282, 5'd0, 27'h0000001c, 5'd5, 27'h000000b7, 32'h00000400,
  1'd1,  5'd26, 27'h000003ad, 5'd4, 27'h00000135, 5'd19, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000078, 5'd3, 27'h00000230, 5'd29, 27'h000000ed, 32'h00000400,
  1'd1,  5'd27, 27'h000002f0, 5'd13, 27'h0000016e, 5'd10, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f1, 5'd13, 27'h00000002, 5'd18, 27'h00000300, 32'h00000400,
  1'd1,  5'd29, 27'h00000016, 5'd13, 27'h000001b0, 5'd29, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007c, 5'd20, 27'h00000313, 5'd6, 27'h00000267, 32'h00000400,
  1'd1,  5'd28, 27'h00000167, 5'd25, 27'h0000002a, 5'd15, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000029e, 5'd22, 27'h000002c6, 5'd28, 27'h0000018d, 32'h00000400,
  1'd1,  5'd8, 27'h00000170, 5'd6, 27'h00000257, 5'd1, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001b6, 5'd7, 27'h000002b5, 5'd14, 27'h00000284, 32'h00000400,
  1'd1,  5'd10, 27'h0000012c, 5'd9, 27'h000003d6, 5'd20, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000363, 5'd16, 27'h000001e7, 5'd0, 27'h00000002, 32'h00000400,
  1'd1,  5'd9, 27'h0000037f, 5'd20, 27'h0000016a, 5'd11, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000188, 5'd19, 27'h000001eb, 5'd22, 27'h0000032d, 32'h00000400,
  1'd1,  5'd5, 27'h00000279, 5'd29, 27'h00000225, 5'd4, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000153, 5'd30, 27'h000002ec, 5'd13, 27'h0000016c, 32'h00000400,
  1'd1,  5'd7, 27'h000000de, 5'd27, 27'h00000364, 5'd21, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000123, 5'd7, 27'h000003c8, 5'd0, 27'h000001b0, 32'h00000400,
  1'd1,  5'd16, 27'h000003d5, 5'd10, 27'h00000101, 5'd11, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021e, 5'd10, 27'h00000093, 5'd22, 27'h0000033c, 32'h00000400,
  1'd1,  5'd19, 27'h00000118, 5'd20, 27'h000001eb, 5'd0, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003cc, 5'd16, 27'h00000060, 5'd11, 27'h000002b2, 32'h00000400,
  1'd1,  5'd16, 27'h000003b9, 5'd20, 27'h0000010f, 5'd23, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000007f, 5'd29, 27'h00000014, 5'd2, 27'h0000032e, 32'h00000400,
  1'd1,  5'd17, 27'h000003d3, 5'd26, 27'h000002e6, 5'd11, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ac, 5'd27, 27'h0000022b, 5'd24, 27'h000003a4, 32'h00000400,
  1'd1,  5'd27, 27'h00000333, 5'd5, 27'h000003bf, 5'd1, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000226, 5'd8, 27'h00000262, 5'd12, 27'h000002ac, 32'h00000400,
  1'd1,  5'd28, 27'h0000022d, 5'd8, 27'h000000ee, 5'd21, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000007, 5'd20, 27'h00000284, 5'd0, 27'h0000027b, 32'h00000400,
  1'd1,  5'd27, 27'h00000348, 5'd15, 27'h0000025e, 5'd10, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025c, 5'd16, 27'h000002e0, 5'd24, 27'h000001be, 32'h00000400,
  1'd1,  5'd26, 27'h000002ea, 5'd28, 27'h000000c9, 5'd1, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c8, 5'd26, 27'h000002de, 5'd12, 27'h000001bd, 32'h00000400,
  1'd1,  5'd30, 27'h00000279, 5'd27, 27'h000000f3, 5'd23, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f6, 5'd9, 27'h000003e0, 5'd7, 27'h00000354, 32'h00000400,
  1'd1,  5'd7, 27'h00000110, 5'd9, 27'h000000d5, 5'd15, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002cd, 5'd8, 27'h00000164, 5'd27, 27'h000003e1, 32'h00000400,
  1'd1,  5'd7, 27'h000002a0, 5'd20, 27'h000000cf, 5'd5, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000154, 5'd19, 27'h00000269, 5'd17, 27'h00000342, 32'h00000400,
  1'd1,  5'd5, 27'h00000391, 5'd20, 27'h000001f4, 5'd29, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000340, 5'd26, 27'h00000227, 5'd9, 27'h00000275, 32'h00000400,
  1'd1,  5'd7, 27'h000000d0, 5'd28, 27'h0000030c, 5'd18, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000d5, 5'd26, 27'h00000365, 5'd29, 27'h000002ac, 32'h00000400,
  1'd1,  5'd15, 27'h0000025a, 5'd6, 27'h000002f9, 5'd7, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000034, 5'd6, 27'h0000003a, 5'd16, 27'h00000395, 32'h00000400,
  1'd1,  5'd19, 27'h000002ca, 5'd8, 27'h0000029e, 5'd29, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000005c, 5'd18, 27'h00000010, 5'd5, 27'h0000013a, 32'h00000400,
  1'd1,  5'd15, 27'h00000217, 5'd19, 27'h0000003a, 5'd18, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003be, 5'd16, 27'h0000009d, 5'd27, 27'h000002c2, 32'h00000400,
  1'd1,  5'd16, 27'h000000e0, 5'd30, 27'h000003e2, 5'd8, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000190, 5'd29, 27'h000000a1, 5'd18, 27'h0000039c, 32'h00000400,
  1'd1,  5'd18, 27'h0000027d, 5'd26, 27'h00000268, 5'd28, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000e5, 5'd9, 27'h00000251, 5'd5, 27'h00000221, 32'h00000400,
  1'd1,  5'd27, 27'h000000e7, 5'd9, 27'h000003f3, 5'd15, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000226, 5'd9, 27'h000000e2, 5'd30, 27'h00000348, 32'h00000400,
  1'd1,  5'd29, 27'h000002df, 5'd19, 27'h000003b5, 5'd8, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000003b, 5'd16, 27'h000001ef, 5'd18, 27'h00000234, 32'h00000400,
  1'd1,  5'd27, 27'h0000035d, 5'd17, 27'h00000076, 5'd29, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000011b, 5'd26, 27'h00000019, 5'd5, 27'h0000020a, 32'h00000400,
  1'd1,  5'd27, 27'h00000162, 5'd28, 27'h00000234, 5'd16, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000255, 5'd28, 27'h000001fe, 5'd29, 27'h000002a8, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000000d7, 5'd0, 27'h0000021c, 5'd2, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000399, 5'd2, 27'h00000035, 5'd15, 27'h00000040, 32'h00000400,
  1'd1,  5'd3, 27'h0000037e, 5'd2, 27'h000002f3, 5'd23, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000208, 5'd11, 27'h00000256, 5'd1, 27'h00000238, 32'h00000400,
  1'd1,  5'd0, 27'h00000020, 5'd14, 27'h000001ae, 5'd11, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000010, 5'd13, 27'h000003cf, 5'd21, 27'h000000b6, 32'h00000400,
  1'd1,  5'd4, 27'h0000022d, 5'd24, 27'h00000256, 5'd1, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000030f, 5'd25, 27'h0000030b, 5'd12, 27'h0000005f, 32'h00000400,
  1'd1,  5'd0, 27'h00000240, 5'd23, 27'h00000181, 5'd23, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020f, 5'd0, 27'h0000032b, 5'd1, 27'h00000309, 32'h00000400,
  1'd1,  5'd13, 27'h000001a0, 5'd1, 27'h000003fd, 5'd14, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f3, 5'd1, 27'h00000398, 5'd21, 27'h000000cd, 32'h00000400,
  1'd1,  5'd10, 27'h00000205, 5'd11, 27'h0000017f, 5'd2, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000249, 5'd14, 27'h000000cc, 5'd10, 27'h00000305, 32'h00000400,
  1'd1,  5'd14, 27'h000003fc, 5'd13, 27'h000003db, 5'd21, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000013f, 5'd22, 27'h0000003d, 5'd4, 27'h000001e2, 32'h00000400,
  1'd1,  5'd12, 27'h000001b0, 5'd24, 27'h000001c6, 5'd13, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000039c, 5'd21, 27'h00000156, 5'd23, 27'h00000041, 32'h00000400,
  1'd1,  5'd22, 27'h00000074, 5'd1, 27'h00000066, 5'd5, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000026a, 5'd4, 27'h00000204, 5'd14, 27'h00000024, 32'h00000400,
  1'd1,  5'd20, 27'h0000032e, 5'd4, 27'h00000348, 5'd25, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000022a, 5'd12, 27'h000000e6, 5'd3, 27'h00000283, 32'h00000400,
  1'd1,  5'd20, 27'h000003f8, 5'd13, 27'h00000383, 5'd10, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000012c, 5'd15, 27'h00000074, 5'd20, 27'h000003cf, 32'h00000400,
  1'd1,  5'd23, 27'h000002a5, 5'd20, 27'h0000030e, 5'd1, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000032, 5'd21, 27'h00000105, 5'd12, 27'h00000209, 32'h00000400,
  1'd1,  5'd24, 27'h000003c6, 5'd20, 27'h000003f1, 5'd23, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c0, 5'd4, 27'h00000374, 5'd8, 27'h000003df, 32'h00000400,
  1'd1,  5'd3, 27'h0000035d, 5'd0, 27'h00000242, 5'd19, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000300, 5'd3, 27'h000000a9, 5'd30, 27'h0000018c, 32'h00000400,
  1'd1,  5'd0, 27'h000001a7, 5'd10, 27'h000003e6, 5'd7, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000194, 5'd11, 27'h0000007e, 5'd17, 27'h000000d1, 32'h00000400,
  1'd1,  5'd2, 27'h0000012a, 5'd11, 27'h00000318, 5'd29, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000017b, 5'd22, 27'h000000af, 5'd6, 27'h00000118, 32'h00000400,
  1'd1,  5'd2, 27'h00000392, 5'd23, 27'h00000372, 5'd19, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000016, 5'd24, 27'h00000033, 5'd28, 27'h0000031a, 32'h00000400,
  1'd1,  5'd11, 27'h0000003e, 5'd3, 27'h000003d3, 5'd7, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000006d, 5'd0, 27'h00000321, 5'd18, 27'h0000030a, 32'h00000400,
  1'd1,  5'd11, 27'h00000097, 5'd0, 27'h0000006b, 5'd27, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d8, 5'd15, 27'h0000014a, 5'd9, 27'h00000364, 32'h00000400,
  1'd1,  5'd11, 27'h00000156, 5'd11, 27'h0000007c, 5'd16, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001bf, 5'd13, 27'h00000162, 5'd26, 27'h000003b5, 32'h00000400,
  1'd1,  5'd12, 27'h0000013f, 5'd20, 27'h00000378, 5'd7, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000088, 5'd23, 27'h00000102, 5'd16, 27'h00000375, 32'h00000400,
  1'd1,  5'd13, 27'h000003c4, 5'd22, 27'h000001d5, 5'd28, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e6, 5'd3, 27'h00000308, 5'd10, 27'h0000012b, 32'h00000400,
  1'd1,  5'd23, 27'h000001e5, 5'd1, 27'h00000110, 5'd19, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000026b, 5'd0, 27'h000002af, 5'd28, 27'h00000175, 32'h00000400,
  1'd1,  5'd22, 27'h00000193, 5'd11, 27'h000002be, 5'd5, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002f3, 5'd12, 27'h000003f6, 5'd17, 27'h00000308, 32'h00000400,
  1'd1,  5'd24, 27'h000003f9, 5'd11, 27'h00000294, 5'd29, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002af, 5'd20, 27'h000003ce, 5'd7, 27'h00000121, 32'h00000400,
  1'd1,  5'd22, 27'h00000377, 5'd23, 27'h0000003f, 5'd18, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000020a, 5'd25, 27'h00000003, 5'd30, 27'h00000155, 32'h00000400,
  1'd1,  5'd3, 27'h000000f3, 5'd5, 27'h0000013b, 5'd0, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002d, 5'd9, 27'h0000014e, 5'd15, 27'h00000044, 32'h00000400,
  1'd1,  5'd1, 27'h0000016e, 5'd8, 27'h000000c1, 5'd21, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000035e, 5'd18, 27'h000003b8, 5'd1, 27'h0000034f, 32'h00000400,
  1'd1,  5'd1, 27'h0000010f, 5'd18, 27'h00000088, 5'd13, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000269, 5'd16, 27'h00000161, 5'd21, 27'h0000016e, 32'h00000400,
  1'd1,  5'd3, 27'h000003c9, 5'd26, 27'h00000305, 5'd0, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017d, 5'd30, 27'h0000006e, 5'd12, 27'h00000312, 32'h00000400,
  1'd1,  5'd2, 27'h000000c4, 5'd30, 27'h00000066, 5'd22, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003d4, 5'd9, 27'h0000020f, 5'd1, 27'h0000027c, 32'h00000400,
  1'd1,  5'd15, 27'h0000013b, 5'd5, 27'h00000183, 5'd14, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000369, 5'd6, 27'h00000075, 5'd23, 27'h000001ff, 32'h00000400,
  1'd1,  5'd12, 27'h000001ba, 5'd16, 27'h000001da, 5'd0, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000dd, 5'd19, 27'h00000201, 5'd14, 27'h00000152, 32'h00000400,
  1'd1,  5'd10, 27'h000001f8, 5'd19, 27'h000002e3, 5'd25, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000279, 5'd27, 27'h000002e3, 5'd3, 27'h0000001a, 32'h00000400,
  1'd1,  5'd12, 27'h000000ba, 5'd25, 27'h00000375, 5'd10, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000149, 5'd29, 27'h000002e3, 5'd25, 27'h00000088, 32'h00000400,
  1'd1,  5'd24, 27'h000002fd, 5'd6, 27'h0000038a, 5'd4, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000364, 5'd10, 27'h0000013e, 5'd11, 27'h000001f9, 32'h00000400,
  1'd1,  5'd25, 27'h00000084, 5'd8, 27'h000000ae, 5'd21, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000bc, 5'd15, 27'h0000030a, 5'd4, 27'h0000020a, 32'h00000400,
  1'd1,  5'd20, 27'h00000322, 5'd20, 27'h000000a1, 5'd11, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000260, 5'd15, 27'h000002ef, 5'd23, 27'h0000013d, 32'h00000400,
  1'd1,  5'd21, 27'h000000ba, 5'd29, 27'h0000030f, 5'd1, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000225, 5'd27, 27'h000000ec, 5'd10, 27'h00000282, 32'h00000400,
  1'd1,  5'd22, 27'h00000077, 5'd27, 27'h00000351, 5'd21, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000033d, 5'd5, 27'h00000337, 5'd8, 27'h000002d8, 32'h00000400,
  1'd1,  5'd0, 27'h00000264, 5'd6, 27'h000003fd, 5'd18, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000360, 5'd8, 27'h000000a0, 5'd28, 27'h00000285, 32'h00000400,
  1'd1,  5'd5, 27'h00000008, 5'd19, 27'h00000161, 5'd5, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e9, 5'd15, 27'h00000276, 5'd16, 27'h00000060, 32'h00000400,
  1'd1,  5'd4, 27'h0000013d, 5'd15, 27'h0000023b, 5'd28, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000019, 5'd29, 27'h00000298, 5'd6, 27'h000001f7, 32'h00000400,
  1'd1,  5'd2, 27'h00000373, 5'd28, 27'h000003b2, 5'd15, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000187, 5'd28, 27'h000000b8, 5'd25, 27'h000003b5, 32'h00000400,
  1'd1,  5'd12, 27'h00000042, 5'd6, 27'h000002d5, 5'd9, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000340, 5'd6, 27'h000003ac, 5'd18, 27'h0000015d, 32'h00000400,
  1'd1,  5'd11, 27'h000002ce, 5'd8, 27'h000000ac, 5'd25, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000151, 5'd19, 27'h0000012e, 5'd5, 27'h0000033e, 32'h00000400,
  1'd1,  5'd13, 27'h000000d3, 5'd16, 27'h00000038, 5'd16, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000013, 5'd18, 27'h000001d2, 5'd29, 27'h000002b2, 32'h00000400,
  1'd1,  5'd15, 27'h0000019f, 5'd28, 27'h0000007b, 5'd9, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002b8, 5'd28, 27'h000002a4, 5'd20, 27'h00000031, 32'h00000400,
  1'd1,  5'd10, 27'h00000382, 5'd29, 27'h000001c7, 5'd26, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d5, 5'd6, 27'h0000029a, 5'd5, 27'h000001b7, 32'h00000400,
  1'd1,  5'd23, 27'h00000248, 5'd6, 27'h0000032f, 5'd20, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003eb, 5'd9, 27'h000001e6, 5'd30, 27'h0000005c, 32'h00000400,
  1'd1,  5'd24, 27'h000002a9, 5'd16, 27'h000003c8, 5'd6, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ce, 5'd19, 27'h00000244, 5'd20, 27'h00000060, 32'h00000400,
  1'd1,  5'd23, 27'h00000382, 5'd20, 27'h000001a1, 5'd30, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000070, 5'd26, 27'h00000262, 5'd10, 27'h000000af, 32'h00000400,
  1'd1,  5'd24, 27'h0000006b, 5'd28, 27'h00000069, 5'd18, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000316, 5'd29, 27'h00000013, 5'd28, 27'h00000005, 32'h00000400,
  1'd1,  5'd6, 27'h0000014f, 5'd3, 27'h00000256, 5'd9, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000034e, 5'd4, 27'h000002bd, 5'd19, 27'h00000103, 32'h00000400,
  1'd1,  5'd5, 27'h0000028a, 5'd0, 27'h00000267, 5'd26, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000175, 5'd14, 27'h000000b1, 5'd1, 27'h0000006b, 32'h00000400,
  1'd1,  5'd9, 27'h0000020d, 5'd14, 27'h000002a8, 5'd14, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000237, 5'd14, 27'h000001e4, 5'd23, 27'h000002f4, 32'h00000400,
  1'd1,  5'd9, 27'h0000033c, 5'd24, 27'h0000002e, 5'd1, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012d, 5'd24, 27'h000001a1, 5'd11, 27'h0000007e, 32'h00000400,
  1'd1,  5'd8, 27'h00000008, 5'd24, 27'h000002d3, 5'd24, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000111, 5'd0, 27'h00000356, 5'd8, 27'h000000c5, 32'h00000400,
  1'd1,  5'd15, 27'h000002cb, 5'd4, 27'h0000013c, 5'd19, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ad, 5'd4, 27'h00000036, 5'd29, 27'h000001ca, 32'h00000400,
  1'd1,  5'd20, 27'h000000e4, 5'd11, 27'h0000014b, 5'd3, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025a, 5'd10, 27'h000002cd, 5'd13, 27'h000000f9, 32'h00000400,
  1'd1,  5'd17, 27'h000003a0, 5'd12, 27'h00000034, 5'd20, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000370, 5'd21, 27'h00000068, 5'd4, 27'h0000004b, 32'h00000400,
  1'd1,  5'd18, 27'h000003b4, 5'd21, 27'h000003fd, 5'd15, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003c7, 5'd25, 27'h00000243, 5'd21, 27'h000002c9, 32'h00000400,
  1'd1,  5'd26, 27'h000003a7, 5'd0, 27'h00000050, 5'd0, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000166, 5'd3, 27'h00000377, 5'd11, 27'h000002a1, 32'h00000400,
  1'd1,  5'd28, 27'h000002aa, 5'd4, 27'h00000146, 5'd21, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d2, 5'd14, 27'h000000c9, 5'd3, 27'h000000b6, 32'h00000400,
  1'd1,  5'd26, 27'h000000e1, 5'd10, 27'h00000193, 5'd12, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000390, 5'd10, 27'h00000216, 5'd25, 27'h00000050, 32'h00000400,
  1'd1,  5'd29, 27'h0000013f, 5'd22, 27'h0000006c, 5'd2, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000275, 5'd20, 27'h000003e5, 5'd10, 27'h000003b2, 32'h00000400,
  1'd1,  5'd30, 27'h000001b0, 5'd24, 27'h000001df, 5'd24, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e1, 5'd3, 27'h00000397, 5'd2, 27'h00000168, 32'h00000400,
  1'd1,  5'd6, 27'h00000020, 5'd1, 27'h0000029a, 5'd15, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001df, 5'd2, 27'h000002fd, 5'd23, 27'h00000329, 32'h00000400,
  1'd1,  5'd7, 27'h00000197, 5'd13, 27'h000003be, 5'd7, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002a8, 5'd14, 27'h000003e2, 5'd19, 27'h0000019e, 32'h00000400,
  1'd1,  5'd9, 27'h0000006a, 5'd14, 27'h000002aa, 5'd26, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001de, 5'd23, 27'h00000374, 5'd9, 27'h0000008c, 32'h00000400,
  1'd1,  5'd9, 27'h00000365, 5'd23, 27'h000000cd, 5'd18, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013a, 5'd21, 27'h00000330, 5'd26, 27'h000001d0, 32'h00000400,
  1'd1,  5'd17, 27'h000003e8, 5'd2, 27'h0000027a, 5'd0, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ee, 5'd3, 27'h0000030c, 5'd10, 27'h00000268, 32'h00000400,
  1'd1,  5'd18, 27'h0000036d, 5'd3, 27'h000001b4, 5'd25, 27'h00000257, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000022, 5'd12, 27'h00000316, 5'd8, 27'h000000c0, 32'h00000400,
  1'd1,  5'd19, 27'h00000387, 5'd13, 27'h00000060, 5'd15, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e8, 5'd12, 27'h00000019, 5'd28, 27'h0000031e, 32'h00000400,
  1'd1,  5'd18, 27'h00000299, 5'd24, 27'h00000150, 5'd7, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000014c, 5'd24, 27'h0000025b, 5'd17, 27'h000003d8, 32'h00000400,
  1'd1,  5'd19, 27'h000000f4, 5'd22, 27'h00000055, 5'd26, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000214, 5'd2, 27'h00000238, 5'd8, 27'h00000031, 32'h00000400,
  1'd1,  5'd28, 27'h0000008f, 5'd0, 27'h00000308, 5'd19, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ce, 5'd2, 27'h000000fd, 5'd25, 27'h00000372, 32'h00000400,
  1'd1,  5'd26, 27'h000001fa, 5'd12, 27'h000003a6, 5'd6, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000366, 5'd14, 27'h00000336, 5'd18, 27'h0000035b, 32'h00000400,
  1'd1,  5'd28, 27'h000003d5, 5'd14, 27'h0000005e, 5'd28, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001f5, 5'd24, 27'h0000039f, 5'd9, 27'h000000dd, 32'h00000400,
  1'd1,  5'd27, 27'h000001a9, 5'd25, 27'h000002e5, 5'd16, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e2, 5'd23, 27'h00000372, 5'd27, 27'h000001da, 32'h00000400,
  1'd1,  5'd6, 27'h000001f8, 5'd6, 27'h000003a1, 5'd1, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a3, 5'd8, 27'h000001e7, 5'd13, 27'h00000154, 32'h00000400,
  1'd1,  5'd7, 27'h000002ba, 5'd8, 27'h000003af, 5'd21, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000092, 5'd18, 27'h000001cc, 5'd0, 27'h0000024a, 32'h00000400,
  1'd1,  5'd5, 27'h000003cf, 5'd17, 27'h00000138, 5'd10, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032e, 5'd20, 27'h00000004, 5'd22, 27'h00000045, 32'h00000400,
  1'd1,  5'd8, 27'h000001d3, 5'd27, 27'h00000248, 5'd4, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000369, 5'd26, 27'h00000179, 5'd13, 27'h000000d8, 32'h00000400,
  1'd1,  5'd5, 27'h000003f5, 5'd25, 27'h000003d7, 5'd21, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f2, 5'd8, 27'h00000396, 5'd1, 27'h000003f5, 32'h00000400,
  1'd1,  5'd16, 27'h000000ac, 5'd6, 27'h000001a9, 5'd13, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b5, 5'd8, 27'h000003ed, 5'd21, 27'h000003d5, 32'h00000400,
  1'd1,  5'd16, 27'h0000020a, 5'd17, 27'h0000003a, 5'd2, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001fa, 5'd17, 27'h00000225, 5'd15, 27'h000001da, 32'h00000400,
  1'd1,  5'd20, 27'h0000024d, 5'd17, 27'h0000018a, 5'd22, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000395, 5'd30, 27'h00000327, 5'd2, 27'h0000039f, 32'h00000400,
  1'd1,  5'd16, 27'h000003fe, 5'd28, 27'h000002af, 5'd12, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ec, 5'd29, 27'h000002e2, 5'd24, 27'h000001e4, 32'h00000400,
  1'd1,  5'd27, 27'h000002e0, 5'd8, 27'h000000c6, 5'd2, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e7, 5'd9, 27'h000003d4, 5'd13, 27'h0000024a, 32'h00000400,
  1'd1,  5'd29, 27'h00000149, 5'd7, 27'h00000180, 5'd21, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000150, 5'd19, 27'h000000ef, 5'd1, 27'h00000307, 32'h00000400,
  1'd1,  5'd28, 27'h000000f0, 5'd15, 27'h000002c3, 5'd12, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001e0, 5'd18, 27'h00000119, 5'd25, 27'h00000222, 32'h00000400,
  1'd1,  5'd30, 27'h00000244, 5'd29, 27'h00000367, 5'd2, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000015b, 5'd30, 27'h00000363, 5'd11, 27'h00000097, 32'h00000400,
  1'd1,  5'd30, 27'h00000114, 5'd28, 27'h000000ad, 5'd24, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000287, 5'd6, 27'h0000027e, 5'd6, 27'h0000015e, 32'h00000400,
  1'd1,  5'd6, 27'h0000033c, 5'd7, 27'h00000079, 5'd19, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000240, 5'd9, 27'h0000038a, 5'd26, 27'h0000028c, 32'h00000400,
  1'd1,  5'd9, 27'h000003c1, 5'd17, 27'h00000036, 5'd6, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c0, 5'd15, 27'h00000392, 5'd18, 27'h000003bc, 32'h00000400,
  1'd1,  5'd9, 27'h00000236, 5'd20, 27'h00000089, 5'd29, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000293, 5'd30, 27'h000001b3, 5'd8, 27'h00000190, 32'h00000400,
  1'd1,  5'd8, 27'h00000247, 5'd27, 27'h000001a9, 5'd20, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b9, 5'd26, 27'h00000383, 5'd26, 27'h000000ce, 32'h00000400,
  1'd1,  5'd17, 27'h000002e4, 5'd7, 27'h000002b5, 5'd9, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f5, 5'd9, 27'h00000228, 5'd16, 27'h0000017f, 32'h00000400,
  1'd1,  5'd20, 27'h000001a1, 5'd6, 27'h00000010, 5'd27, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000023c, 5'd18, 27'h0000013d, 5'd6, 27'h0000023e, 32'h00000400,
  1'd1,  5'd19, 27'h000003ec, 5'd18, 27'h00000183, 5'd18, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002be, 5'd15, 27'h00000225, 5'd27, 27'h0000010e, 32'h00000400,
  1'd1,  5'd19, 27'h00000083, 5'd30, 27'h00000088, 5'd6, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b5, 5'd29, 27'h00000137, 5'd17, 27'h00000323, 32'h00000400,
  1'd1,  5'd17, 27'h00000319, 5'd25, 27'h00000376, 5'd26, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000007b, 5'd6, 27'h000000d2, 5'd6, 27'h00000370, 32'h00000400,
  1'd1,  5'd26, 27'h0000001b, 5'd7, 27'h00000278, 5'd20, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000033f, 5'd9, 27'h000003d2, 5'd29, 27'h00000188, 32'h00000400,
  1'd1,  5'd27, 27'h0000010a, 5'd19, 27'h000001c7, 5'd7, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000150, 5'd15, 27'h000003e8, 5'd17, 27'h0000006c, 32'h00000400,
  1'd1,  5'd30, 27'h000003d3, 5'd18, 27'h00000296, 5'd28, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000000a, 5'd26, 27'h000001e9, 5'd6, 27'h00000084, 32'h00000400,
  1'd1,  5'd30, 27'h00000108, 5'd26, 27'h00000305, 5'd18, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000019d, 5'd27, 27'h00000287, 5'd30, 27'h00000351, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000054, 5'd2, 27'h0000031b, 5'd1, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000381, 5'd1, 27'h00000290, 5'd14, 27'h000002d7, 32'h00000400,
  1'd1,  5'd1, 27'h000003f3, 5'd4, 27'h000000b3, 5'd21, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000001d, 5'd15, 27'h00000130, 5'd2, 27'h000003b0, 32'h00000400,
  1'd1,  5'd0, 27'h000003c5, 5'd13, 27'h00000258, 5'd11, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001f6, 5'd14, 27'h000000a0, 5'd25, 27'h000002b3, 32'h00000400,
  1'd1,  5'd0, 27'h00000318, 5'd23, 27'h0000006a, 5'd4, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a7, 5'd22, 27'h00000266, 5'd13, 27'h000003ee, 32'h00000400,
  1'd1,  5'd4, 27'h00000396, 5'd22, 27'h000000ca, 5'd24, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c7, 5'd4, 27'h000000fc, 5'd0, 27'h00000067, 32'h00000400,
  1'd1,  5'd15, 27'h000000c4, 5'd3, 27'h000000dc, 5'd14, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000028e, 5'd4, 27'h0000022c, 5'd23, 27'h00000347, 32'h00000400,
  1'd1,  5'd11, 27'h000002df, 5'd11, 27'h0000005d, 5'd3, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000371, 5'd13, 27'h00000327, 5'd14, 27'h000000b7, 32'h00000400,
  1'd1,  5'd14, 27'h0000009d, 5'd13, 27'h0000032c, 5'd23, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000390, 5'd24, 27'h00000095, 5'd4, 27'h00000350, 32'h00000400,
  1'd1,  5'd15, 27'h000000ef, 5'd24, 27'h00000261, 5'd11, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000015f, 5'd22, 27'h000003e8, 5'd23, 27'h000002fc, 32'h00000400,
  1'd1,  5'd25, 27'h000002a3, 5'd1, 27'h000001a8, 5'd2, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000033a, 5'd4, 27'h00000103, 5'd15, 27'h000001dd, 32'h00000400,
  1'd1,  5'd25, 27'h00000209, 5'd0, 27'h0000037c, 5'd24, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000af, 5'd12, 27'h00000324, 5'd2, 27'h00000023, 32'h00000400,
  1'd1,  5'd22, 27'h000000a4, 5'd13, 27'h000001c3, 5'd10, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000208, 5'd14, 27'h000002a9, 5'd22, 27'h000002cb, 32'h00000400,
  1'd1,  5'd21, 27'h000001ba, 5'd21, 27'h00000235, 5'd0, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001cc, 5'd25, 27'h00000256, 5'd10, 27'h0000016e, 32'h00000400,
  1'd1,  5'd21, 27'h000001e9, 5'd23, 27'h0000010b, 5'd23, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d8, 5'd1, 27'h000003dd, 5'd7, 27'h000003f9, 32'h00000400,
  1'd1,  5'd4, 27'h000003a6, 5'd3, 27'h0000021c, 5'd20, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000037b, 5'd1, 27'h0000001d, 5'd27, 27'h00000122, 32'h00000400,
  1'd1,  5'd4, 27'h0000010a, 5'd15, 27'h0000014d, 5'd8, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000035a, 5'd10, 27'h000002d9, 5'd17, 27'h00000324, 32'h00000400,
  1'd1,  5'd2, 27'h000002b3, 5'd11, 27'h000002c6, 5'd30, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000134, 5'd25, 27'h0000034b, 5'd6, 27'h000003bb, 32'h00000400,
  1'd1,  5'd2, 27'h0000017a, 5'd24, 27'h00000112, 5'd16, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000366, 5'd21, 27'h0000006b, 5'd27, 27'h0000000a, 32'h00000400,
  1'd1,  5'd12, 27'h000000fe, 5'd2, 27'h000003fc, 5'd9, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000229, 5'd0, 27'h000000c1, 5'd19, 27'h00000359, 32'h00000400,
  1'd1,  5'd13, 27'h00000133, 5'd5, 27'h0000002d, 5'd29, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000032d, 5'd11, 27'h00000153, 5'd9, 27'h00000323, 32'h00000400,
  1'd1,  5'd13, 27'h000000b9, 5'd13, 27'h000001eb, 5'd20, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002bc, 5'd12, 27'h0000006a, 5'd29, 27'h000000ae, 32'h00000400,
  1'd1,  5'd11, 27'h000000c7, 5'd21, 27'h00000261, 5'd8, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008a, 5'd22, 27'h0000019e, 5'd19, 27'h000003a8, 32'h00000400,
  1'd1,  5'd12, 27'h000000e6, 5'd22, 27'h000003aa, 5'd28, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000325, 5'd2, 27'h00000130, 5'd5, 27'h000001fb, 32'h00000400,
  1'd1,  5'd25, 27'h00000112, 5'd2, 27'h00000146, 5'd16, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000023, 5'd2, 27'h000003bc, 5'd30, 27'h000003a4, 32'h00000400,
  1'd1,  5'd23, 27'h0000015a, 5'd12, 27'h00000035, 5'd7, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000017b, 5'd11, 27'h000000f2, 5'd18, 27'h00000221, 32'h00000400,
  1'd1,  5'd20, 27'h0000038d, 5'd12, 27'h0000019b, 5'd29, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000256, 5'd24, 27'h0000001c, 5'd7, 27'h00000010, 32'h00000400,
  1'd1,  5'd21, 27'h00000399, 5'd24, 27'h000002d2, 5'd16, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003de, 5'd23, 27'h000000f7, 5'd30, 27'h00000127, 32'h00000400,
  1'd1,  5'd4, 27'h00000263, 5'd9, 27'h000002ab, 5'd4, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000285, 5'd9, 27'h00000241, 5'd11, 27'h00000149, 32'h00000400,
  1'd1,  5'd3, 27'h000000db, 5'd9, 27'h00000165, 5'd24, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000315, 5'd19, 27'h00000302, 5'd0, 27'h00000378, 32'h00000400,
  1'd1,  5'd4, 27'h000002d8, 5'd19, 27'h000000a3, 5'd11, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027b, 5'd17, 27'h00000318, 5'd21, 27'h0000026b, 32'h00000400,
  1'd1,  5'd0, 27'h00000062, 5'd27, 27'h00000141, 5'd3, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000014, 5'd28, 27'h00000059, 5'd11, 27'h000002d5, 32'h00000400,
  1'd1,  5'd3, 27'h0000035d, 5'd27, 27'h00000114, 5'd24, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e1, 5'd7, 27'h00000169, 5'd4, 27'h000001ef, 32'h00000400,
  1'd1,  5'd14, 27'h0000006b, 5'd8, 27'h0000019d, 5'd13, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002be, 5'd6, 27'h000001e8, 5'd21, 27'h000000c5, 32'h00000400,
  1'd1,  5'd12, 27'h000003e8, 5'd20, 27'h000000ba, 5'd2, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000cd, 5'd17, 27'h000000c2, 5'd12, 27'h0000035a, 32'h00000400,
  1'd1,  5'd10, 27'h000001d1, 5'd19, 27'h00000038, 5'd22, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000260, 5'd29, 27'h000000a9, 5'd2, 27'h00000081, 32'h00000400,
  1'd1,  5'd12, 27'h0000018a, 5'd27, 27'h00000369, 5'd11, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000022c, 5'd28, 27'h00000185, 5'd23, 27'h0000014d, 32'h00000400,
  1'd1,  5'd21, 27'h000000ca, 5'd6, 27'h000002a6, 5'd1, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031b, 5'd6, 27'h00000386, 5'd13, 27'h00000249, 32'h00000400,
  1'd1,  5'd21, 27'h00000334, 5'd10, 27'h00000044, 5'd23, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000090, 5'd18, 27'h0000022c, 5'd2, 27'h0000030b, 32'h00000400,
  1'd1,  5'd21, 27'h00000391, 5'd18, 27'h000002f6, 5'd13, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000255, 5'd20, 27'h0000003c, 5'd22, 27'h00000315, 32'h00000400,
  1'd1,  5'd22, 27'h0000032c, 5'd27, 27'h000000fb, 5'd2, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000012c, 5'd28, 27'h00000278, 5'd11, 27'h0000012a, 32'h00000400,
  1'd1,  5'd23, 27'h000001ca, 5'd27, 27'h000000a3, 5'd24, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000243, 5'd8, 27'h00000265, 5'd6, 27'h000000d1, 32'h00000400,
  1'd1,  5'd3, 27'h000002e8, 5'd8, 27'h000000f7, 5'd16, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000246, 5'd9, 27'h000001ee, 5'd28, 27'h00000005, 32'h00000400,
  1'd1,  5'd1, 27'h000001ca, 5'd20, 27'h0000018d, 5'd6, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000a3, 5'd20, 27'h0000020c, 5'd17, 27'h00000342, 32'h00000400,
  1'd1,  5'd2, 27'h000003eb, 5'd18, 27'h00000154, 5'd30, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000018, 5'd26, 27'h0000009e, 5'd9, 27'h0000011a, 32'h00000400,
  1'd1,  5'd5, 27'h00000010, 5'd29, 27'h0000029a, 5'd17, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a2, 5'd30, 27'h00000123, 5'd26, 27'h00000111, 32'h00000400,
  1'd1,  5'd14, 27'h0000018f, 5'd7, 27'h000003d7, 5'd8, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000007, 5'd7, 27'h00000189, 5'd17, 27'h000001a4, 32'h00000400,
  1'd1,  5'd13, 27'h00000180, 5'd8, 27'h000000e3, 5'd27, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020d, 5'd20, 27'h00000132, 5'd5, 27'h0000025b, 32'h00000400,
  1'd1,  5'd12, 27'h000001e9, 5'd16, 27'h000003ac, 5'd17, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000017f, 5'd20, 27'h000001a8, 5'd26, 27'h00000063, 32'h00000400,
  1'd1,  5'd13, 27'h000000eb, 5'd28, 27'h000002cd, 5'd6, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000161, 5'd28, 27'h0000022e, 5'd19, 27'h0000000d, 32'h00000400,
  1'd1,  5'd12, 27'h000001b5, 5'd26, 27'h000003fb, 5'd27, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001b5, 5'd8, 27'h000001ca, 5'd7, 27'h0000007d, 32'h00000400,
  1'd1,  5'd21, 27'h000002fc, 5'd10, 27'h0000001c, 5'd20, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003bf, 5'd5, 27'h00000250, 5'd26, 27'h000002a6, 32'h00000400,
  1'd1,  5'd23, 27'h00000107, 5'd16, 27'h0000000d, 5'd7, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f8, 5'd20, 27'h000001a2, 5'd15, 27'h0000031f, 32'h00000400,
  1'd1,  5'd20, 27'h00000309, 5'd20, 27'h000001e3, 5'd26, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000143, 5'd30, 27'h0000013b, 5'd9, 27'h000002e6, 32'h00000400,
  1'd1,  5'd25, 27'h000001aa, 5'd30, 27'h0000039d, 5'd17, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000008, 5'd29, 27'h0000002b, 5'd29, 27'h000000cc, 32'h00000400,
  1'd1,  5'd8, 27'h000000eb, 5'd3, 27'h00000265, 5'd5, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f4, 5'd2, 27'h00000344, 5'd16, 27'h000002c0, 32'h00000400,
  1'd1,  5'd6, 27'h0000038d, 5'd4, 27'h000002f0, 5'd28, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000016d, 5'd11, 27'h000000c5, 5'd5, 27'h00000057, 32'h00000400,
  1'd1,  5'd6, 27'h00000377, 5'd12, 27'h00000249, 5'd13, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000359, 5'd10, 27'h0000038d, 5'd24, 27'h000003f4, 32'h00000400,
  1'd1,  5'd7, 27'h000000c8, 5'd25, 27'h00000045, 5'd0, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a5, 5'd24, 27'h0000011c, 5'd11, 27'h00000294, 32'h00000400,
  1'd1,  5'd6, 27'h000003c1, 5'd21, 27'h000001b0, 5'd22, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000013e, 5'd0, 27'h00000247, 5'd8, 27'h000003b5, 32'h00000400,
  1'd1,  5'd19, 27'h0000001f, 5'd1, 27'h0000026a, 5'd17, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001d2, 5'd2, 27'h00000382, 5'd29, 27'h0000021f, 32'h00000400,
  1'd1,  5'd20, 27'h000001ae, 5'd11, 27'h000003a5, 5'd3, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000020c, 5'd10, 27'h000001a4, 5'd14, 27'h000003be, 32'h00000400,
  1'd1,  5'd18, 27'h000003eb, 5'd11, 27'h000003c0, 5'd23, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a2, 5'd23, 27'h0000004d, 5'd1, 27'h000002cf, 32'h00000400,
  1'd1,  5'd18, 27'h00000333, 5'd21, 27'h000000e9, 5'd12, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011c, 5'd23, 27'h000003e4, 5'd21, 27'h0000015d, 32'h00000400,
  1'd1,  5'd30, 27'h000002c2, 5'd2, 27'h000002d3, 5'd1, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000131, 5'd3, 27'h000000fd, 5'd13, 27'h0000029d, 32'h00000400,
  1'd1,  5'd26, 27'h000003f9, 5'd4, 27'h00000100, 5'd20, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000138, 5'd12, 27'h0000002f, 5'd0, 27'h000001ab, 32'h00000400,
  1'd1,  5'd27, 27'h000000b4, 5'd13, 27'h0000019a, 5'd14, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000117, 5'd15, 27'h00000050, 5'd22, 27'h000002d0, 32'h00000400,
  1'd1,  5'd29, 27'h00000095, 5'd22, 27'h000002db, 5'd2, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000df, 5'd24, 27'h0000028a, 5'd15, 27'h0000018b, 32'h00000400,
  1'd1,  5'd30, 27'h0000020f, 5'd21, 27'h00000237, 5'd24, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000289, 5'd2, 27'h0000029a, 5'd3, 27'h00000285, 32'h00000400,
  1'd1,  5'd5, 27'h00000144, 5'd1, 27'h000000d0, 5'd15, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000113, 5'd2, 27'h000002da, 5'd23, 27'h00000334, 32'h00000400,
  1'd1,  5'd7, 27'h0000027c, 5'd13, 27'h000003d8, 5'd7, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000033a, 5'd15, 27'h00000115, 5'd20, 27'h00000263, 32'h00000400,
  1'd1,  5'd5, 27'h000000f1, 5'd11, 27'h000003de, 5'd29, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000147, 5'd25, 27'h000002d7, 5'd6, 27'h000003d3, 32'h00000400,
  1'd1,  5'd8, 27'h000000fd, 5'd22, 27'h00000186, 5'd16, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000140, 5'd22, 27'h0000006b, 5'd26, 27'h00000131, 32'h00000400,
  1'd1,  5'd17, 27'h0000029c, 5'd0, 27'h000002cd, 5'd4, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ff, 5'd3, 27'h000002c8, 5'd12, 27'h00000371, 32'h00000400,
  1'd1,  5'd16, 27'h00000059, 5'd0, 27'h00000319, 5'd25, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000328, 5'd12, 27'h000003e9, 5'd7, 27'h00000137, 32'h00000400,
  1'd1,  5'd19, 27'h000000a4, 5'd10, 27'h00000280, 5'd17, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034a, 5'd10, 27'h00000302, 5'd28, 27'h00000075, 32'h00000400,
  1'd1,  5'd16, 27'h00000132, 5'd24, 27'h00000166, 5'd5, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003b7, 5'd21, 27'h000000e6, 5'd20, 27'h00000284, 32'h00000400,
  1'd1,  5'd16, 27'h00000062, 5'd21, 27'h000003f2, 5'd29, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000137, 5'd4, 27'h000000d3, 5'd8, 27'h0000018c, 32'h00000400,
  1'd1,  5'd30, 27'h000001ce, 5'd0, 27'h00000214, 5'd17, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002b7, 5'd5, 27'h00000099, 5'd28, 27'h000001a1, 32'h00000400,
  1'd1,  5'd29, 27'h00000397, 5'd11, 27'h0000010a, 5'd6, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000114, 5'd10, 27'h000003e5, 5'd17, 27'h00000242, 32'h00000400,
  1'd1,  5'd29, 27'h0000037d, 5'd14, 27'h00000218, 5'd29, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024a, 5'd24, 27'h000003cd, 5'd7, 27'h000003ab, 32'h00000400,
  1'd1,  5'd27, 27'h00000142, 5'd24, 27'h00000195, 5'd18, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000345, 5'd24, 27'h000003ed, 5'd30, 27'h00000021, 32'h00000400,
  1'd1,  5'd7, 27'h000003e0, 5'd9, 27'h00000190, 5'd3, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000001f, 5'd7, 27'h00000013, 5'd15, 27'h00000132, 32'h00000400,
  1'd1,  5'd5, 27'h00000111, 5'd7, 27'h000001f5, 5'd23, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000036f, 5'd19, 27'h000002fc, 5'd4, 27'h000000e7, 32'h00000400,
  1'd1,  5'd8, 27'h000000ed, 5'd16, 27'h00000072, 5'd10, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000211, 5'd18, 27'h000003cd, 5'd24, 27'h0000037f, 32'h00000400,
  1'd1,  5'd8, 27'h000002e5, 5'd25, 27'h000003dc, 5'd0, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001b6, 5'd27, 27'h00000075, 5'd14, 27'h000000fc, 32'h00000400,
  1'd1,  5'd8, 27'h000003e6, 5'd29, 27'h00000394, 5'd22, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000015e, 5'd9, 27'h00000231, 5'd1, 27'h000002e9, 32'h00000400,
  1'd1,  5'd19, 27'h000001bb, 5'd9, 27'h0000027a, 5'd11, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a3, 5'd6, 27'h000003dd, 5'd24, 27'h000003e7, 32'h00000400,
  1'd1,  5'd18, 27'h0000018b, 5'd18, 27'h0000002e, 5'd4, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000a4, 5'd19, 27'h00000373, 5'd14, 27'h00000165, 32'h00000400,
  1'd1,  5'd18, 27'h000003d8, 5'd20, 27'h0000014c, 5'd24, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000382, 5'd27, 27'h0000011a, 5'd1, 27'h00000211, 32'h00000400,
  1'd1,  5'd15, 27'h000002d3, 5'd26, 27'h000003ff, 5'd12, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e9, 5'd27, 27'h00000342, 5'd24, 27'h000001d0, 32'h00000400,
  1'd1,  5'd26, 27'h00000322, 5'd7, 27'h000000c3, 5'd0, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000022, 5'd8, 27'h00000201, 5'd11, 27'h0000022d, 32'h00000400,
  1'd1,  5'd27, 27'h000000c3, 5'd7, 27'h0000023c, 5'd24, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000019c, 5'd18, 27'h00000360, 5'd2, 27'h000000f2, 32'h00000400,
  1'd1,  5'd27, 27'h0000001c, 5'd16, 27'h000002d6, 5'd13, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000036b, 5'd17, 27'h00000201, 5'd25, 27'h00000186, 32'h00000400,
  1'd1,  5'd26, 27'h000003e9, 5'd30, 27'h00000140, 5'd3, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002b1, 5'd29, 27'h000003fc, 5'd12, 27'h00000264, 32'h00000400,
  1'd1,  5'd30, 27'h000001ca, 5'd29, 27'h00000209, 5'd22, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000033b, 5'd8, 27'h000001c3, 5'd9, 27'h000003d9, 32'h00000400,
  1'd1,  5'd5, 27'h000000c9, 5'd8, 27'h0000009c, 5'd17, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a5, 5'd9, 27'h00000028, 5'd29, 27'h0000003a, 32'h00000400,
  1'd1,  5'd8, 27'h00000148, 5'd17, 27'h0000002d, 5'd9, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c8, 5'd18, 27'h000002b9, 5'd18, 27'h000002c9, 32'h00000400,
  1'd1,  5'd7, 27'h000001a8, 5'd19, 27'h00000353, 5'd30, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ed, 5'd29, 27'h000000e9, 5'd6, 27'h00000181, 32'h00000400,
  1'd1,  5'd7, 27'h0000001a, 5'd29, 27'h00000019, 5'd19, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cd, 5'd27, 27'h000002f4, 5'd27, 27'h0000018f, 32'h00000400,
  1'd1,  5'd17, 27'h0000010f, 5'd7, 27'h00000062, 5'd7, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000259, 5'd5, 27'h0000022a, 5'd18, 27'h0000022e, 32'h00000400,
  1'd1,  5'd18, 27'h00000322, 5'd9, 27'h00000273, 5'd30, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a3, 5'd20, 27'h0000018f, 5'd10, 27'h000000c0, 32'h00000400,
  1'd1,  5'd18, 27'h00000359, 5'd19, 27'h000000ca, 5'd19, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000325, 5'd18, 27'h0000023c, 5'd27, 27'h000000a0, 32'h00000400,
  1'd1,  5'd19, 27'h00000345, 5'd27, 27'h0000026f, 5'd5, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000235, 5'd28, 27'h000000b6, 5'd17, 27'h000000a8, 32'h00000400,
  1'd1,  5'd18, 27'h0000026d, 5'd26, 27'h000002df, 5'd26, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000013d, 5'd8, 27'h000001be, 5'd7, 27'h0000002d, 32'h00000400,
  1'd1,  5'd27, 27'h0000018b, 5'd8, 27'h0000032a, 5'd15, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b3, 5'd6, 27'h000001a5, 5'd27, 27'h00000360, 32'h00000400,
  1'd1,  5'd27, 27'h000003e4, 5'd19, 27'h000000ad, 5'd7, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000396, 5'd19, 27'h0000033f, 5'd15, 27'h00000248, 32'h00000400,
  1'd1,  5'd27, 27'h00000269, 5'd16, 27'h0000021b, 5'd28, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000063, 5'd26, 27'h000000e4, 5'd6, 27'h0000021f, 32'h00000400,
  1'd1,  5'd28, 27'h00000220, 5'd29, 27'h00000097, 5'd16, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000091, 5'd28, 27'h000002a0, 5'd30, 27'h00000239, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000001b0, 5'd0, 27'h000003a6, 5'd3, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000373, 5'd3, 27'h000002f8, 5'd11, 27'h000001d6, 32'h00000400,
  1'd1,  5'd4, 27'h000003c9, 5'd4, 27'h000001f7, 5'd22, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001e8, 5'd11, 27'h000003be, 5'd5, 27'h0000002d, 32'h00000400,
  1'd1,  5'd2, 27'h00000343, 5'd13, 27'h00000182, 5'd13, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000170, 5'd14, 27'h000002db, 5'd22, 27'h00000089, 32'h00000400,
  1'd1,  5'd3, 27'h000002dd, 5'd24, 27'h0000039a, 5'd1, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000331, 5'd22, 27'h0000028a, 5'd12, 27'h00000030, 32'h00000400,
  1'd1,  5'd0, 27'h00000334, 5'd22, 27'h00000034, 5'd20, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001b9, 5'd4, 27'h0000026f, 5'd2, 27'h00000317, 32'h00000400,
  1'd1,  5'd11, 27'h00000371, 5'd5, 27'h000000a1, 5'd15, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e4, 5'd0, 27'h00000052, 5'd20, 27'h0000031f, 32'h00000400,
  1'd1,  5'd10, 27'h00000241, 5'd15, 27'h00000077, 5'd1, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000014f, 5'd12, 27'h00000001, 5'd13, 27'h00000067, 32'h00000400,
  1'd1,  5'd11, 27'h0000021c, 5'd13, 27'h00000052, 5'd22, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000395, 5'd22, 27'h000000b5, 5'd1, 27'h000003c2, 32'h00000400,
  1'd1,  5'd11, 27'h0000031a, 5'd22, 27'h00000330, 5'd14, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e4, 5'd25, 27'h0000025e, 5'd23, 27'h000000e0, 32'h00000400,
  1'd1,  5'd24, 27'h000002d0, 5'd3, 27'h0000034f, 5'd4, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000059, 5'd3, 27'h000002ee, 5'd13, 27'h0000007d, 32'h00000400,
  1'd1,  5'd25, 27'h00000129, 5'd1, 27'h000002b2, 5'd23, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000138, 5'd15, 27'h000001fd, 5'd1, 27'h000003ee, 32'h00000400,
  1'd1,  5'd24, 27'h00000397, 5'd13, 27'h00000086, 5'd11, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d5, 5'd14, 27'h00000368, 5'd25, 27'h000001e2, 32'h00000400,
  1'd1,  5'd23, 27'h0000004c, 5'd23, 27'h000003d2, 5'd3, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ac, 5'd24, 27'h000001b9, 5'd12, 27'h00000030, 32'h00000400,
  1'd1,  5'd20, 27'h000002c6, 5'd21, 27'h0000000d, 5'd21, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d6, 5'd3, 27'h0000023c, 5'd8, 27'h000002f8, 32'h00000400,
  1'd1,  5'd3, 27'h00000266, 5'd3, 27'h000000fa, 5'd18, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ed, 5'd0, 27'h000000aa, 5'd30, 27'h000001f0, 32'h00000400,
  1'd1,  5'd0, 27'h0000015b, 5'd12, 27'h00000193, 5'd5, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000074, 5'd10, 27'h000002bc, 5'd15, 27'h00000390, 32'h00000400,
  1'd1,  5'd4, 27'h00000114, 5'd13, 27'h0000013b, 5'd29, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003a7, 5'd25, 27'h000001dc, 5'd6, 27'h0000018a, 32'h00000400,
  1'd1,  5'd1, 27'h000003fe, 5'd24, 27'h00000087, 5'd20, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ed, 5'd23, 27'h00000020, 5'd30, 27'h00000143, 32'h00000400,
  1'd1,  5'd14, 27'h000002f8, 5'd2, 27'h000002bd, 5'd8, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000107, 5'd1, 27'h000000ee, 5'd16, 27'h000000bb, 32'h00000400,
  1'd1,  5'd15, 27'h000000ff, 5'd1, 27'h00000272, 5'd30, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000010d, 5'd10, 27'h0000016a, 5'd9, 27'h000001d7, 32'h00000400,
  1'd1,  5'd14, 27'h00000101, 5'd12, 27'h00000068, 5'd16, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f8, 5'd15, 27'h00000193, 5'd26, 27'h0000006a, 32'h00000400,
  1'd1,  5'd12, 27'h0000034e, 5'd22, 27'h00000177, 5'd6, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ba, 5'd20, 27'h0000036e, 5'd17, 27'h00000188, 32'h00000400,
  1'd1,  5'd11, 27'h0000003c, 5'd24, 27'h0000026d, 5'd28, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000087, 5'd3, 27'h0000032c, 5'd7, 27'h000003f6, 32'h00000400,
  1'd1,  5'd22, 27'h000001ac, 5'd2, 27'h00000246, 5'd19, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000317, 5'd1, 27'h00000079, 5'd27, 27'h000001d3, 32'h00000400,
  1'd1,  5'd22, 27'h0000009d, 5'd11, 27'h0000035b, 5'd5, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000384, 5'd10, 27'h0000037c, 5'd19, 27'h000002ed, 32'h00000400,
  1'd1,  5'd22, 27'h00000045, 5'd13, 27'h000000d9, 5'd29, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000303, 5'd23, 27'h00000381, 5'd7, 27'h00000225, 32'h00000400,
  1'd1,  5'd25, 27'h000002d8, 5'd21, 27'h00000113, 5'd18, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fc, 5'd25, 27'h00000306, 5'd28, 27'h0000039e, 32'h00000400,
  1'd1,  5'd2, 27'h000002fa, 5'd8, 27'h00000290, 5'd1, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000036, 5'd10, 27'h00000124, 5'd12, 27'h000001db, 32'h00000400,
  1'd1,  5'd3, 27'h00000104, 5'd9, 27'h000001fa, 5'd21, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000236, 5'd19, 27'h0000006b, 5'd3, 27'h000001b2, 32'h00000400,
  1'd1,  5'd2, 27'h000003aa, 5'd20, 27'h00000109, 5'd14, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000154, 5'd17, 27'h000002ed, 5'd21, 27'h00000058, 32'h00000400,
  1'd1,  5'd1, 27'h00000082, 5'd27, 27'h0000020a, 5'd0, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a3, 5'd26, 27'h00000380, 5'd10, 27'h0000026c, 32'h00000400,
  1'd1,  5'd2, 27'h00000135, 5'd30, 27'h0000028e, 5'd23, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000237, 5'd8, 27'h00000175, 5'd0, 27'h00000365, 32'h00000400,
  1'd1,  5'd14, 27'h000000a6, 5'd7, 27'h00000225, 5'd10, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002cc, 5'd8, 27'h0000030d, 5'd22, 27'h00000158, 32'h00000400,
  1'd1,  5'd15, 27'h000000e5, 5'd20, 27'h00000092, 5'd1, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e7, 5'd16, 27'h00000097, 5'd11, 27'h000003a3, 32'h00000400,
  1'd1,  5'd12, 27'h000002a2, 5'd19, 27'h00000105, 5'd22, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029f, 5'd26, 27'h00000052, 5'd3, 27'h00000010, 32'h00000400,
  1'd1,  5'd13, 27'h00000055, 5'd29, 27'h00000140, 5'd12, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d2, 5'd30, 27'h000000c7, 5'd22, 27'h000001ff, 32'h00000400,
  1'd1,  5'd20, 27'h000003e1, 5'd10, 27'h00000144, 5'd4, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000135, 5'd6, 27'h000000b7, 5'd14, 27'h0000023b, 32'h00000400,
  1'd1,  5'd21, 27'h000002f9, 5'd7, 27'h00000265, 5'd24, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b8, 5'd17, 27'h00000339, 5'd3, 27'h0000011d, 32'h00000400,
  1'd1,  5'd22, 27'h000001c5, 5'd19, 27'h0000023f, 5'd12, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003b8, 5'd16, 27'h00000164, 5'd21, 27'h0000034b, 32'h00000400,
  1'd1,  5'd24, 27'h00000087, 5'd30, 27'h000003a3, 5'd3, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000358, 5'd27, 27'h00000070, 5'd12, 27'h0000026a, 32'h00000400,
  1'd1,  5'd25, 27'h000001ca, 5'd28, 27'h0000008d, 5'd22, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000011c, 5'd8, 27'h00000199, 5'd5, 27'h00000298, 32'h00000400,
  1'd1,  5'd4, 27'h00000386, 5'd5, 27'h00000198, 5'd18, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000355, 5'd9, 27'h00000043, 5'd29, 27'h0000011b, 32'h00000400,
  1'd1,  5'd3, 27'h0000031e, 5'd19, 27'h00000215, 5'd7, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002b9, 5'd20, 27'h00000217, 5'd19, 27'h00000360, 32'h00000400,
  1'd1,  5'd1, 27'h00000042, 5'd19, 27'h0000010f, 5'd29, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000384, 5'd29, 27'h000000a6, 5'd9, 27'h00000076, 32'h00000400,
  1'd1,  5'd0, 27'h000001c7, 5'd27, 27'h000000c6, 5'd16, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002b6, 5'd30, 27'h000002ae, 5'd26, 27'h00000199, 32'h00000400,
  1'd1,  5'd12, 27'h0000001b, 5'd8, 27'h00000116, 5'd8, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b5, 5'd8, 27'h00000354, 5'd18, 27'h00000157, 32'h00000400,
  1'd1,  5'd10, 27'h0000027f, 5'd9, 27'h0000007f, 5'd29, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002dc, 5'd16, 27'h000000cb, 5'd10, 27'h000000c0, 32'h00000400,
  1'd1,  5'd14, 27'h000000a9, 5'd17, 27'h00000226, 5'd18, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000174, 5'd17, 27'h0000009c, 5'd30, 27'h00000072, 32'h00000400,
  1'd1,  5'd12, 27'h00000205, 5'd26, 27'h0000039f, 5'd5, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000037e, 5'd27, 27'h0000031d, 5'd19, 27'h000000ce, 32'h00000400,
  1'd1,  5'd14, 27'h0000030d, 5'd29, 27'h000001f9, 5'd26, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000cb, 5'd9, 27'h000000e5, 5'd5, 27'h00000331, 32'h00000400,
  1'd1,  5'd24, 27'h00000185, 5'd9, 27'h0000039f, 5'd18, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000032f, 5'd7, 27'h00000082, 5'd27, 27'h0000031b, 32'h00000400,
  1'd1,  5'd23, 27'h0000004b, 5'd15, 27'h000002c6, 5'd9, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000002, 5'd18, 27'h00000245, 5'd17, 27'h000000f2, 32'h00000400,
  1'd1,  5'd23, 27'h00000132, 5'd20, 27'h00000297, 5'd26, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001d4, 5'd30, 27'h00000246, 5'd6, 27'h000000cd, 32'h00000400,
  1'd1,  5'd24, 27'h000002f0, 5'd27, 27'h000001c5, 5'd18, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000c2, 5'd26, 27'h00000165, 5'd30, 27'h000003aa, 32'h00000400,
  1'd1,  5'd9, 27'h00000177, 5'd0, 27'h0000027b, 5'd9, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000cc, 5'd4, 27'h00000312, 5'd16, 27'h0000004d, 32'h00000400,
  1'd1,  5'd9, 27'h00000052, 5'd3, 27'h000003e3, 5'd29, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000259, 5'd13, 27'h0000034d, 5'd3, 27'h000002c2, 32'h00000400,
  1'd1,  5'd9, 27'h00000106, 5'd10, 27'h0000023b, 5'd12, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002aa, 5'd12, 27'h0000038a, 5'd22, 27'h00000361, 32'h00000400,
  1'd1,  5'd8, 27'h00000380, 5'd23, 27'h00000298, 5'd1, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002c0, 5'd20, 27'h000002d0, 5'd12, 27'h00000362, 32'h00000400,
  1'd1,  5'd9, 27'h00000269, 5'd24, 27'h0000012c, 5'd22, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000033e, 5'd4, 27'h0000019b, 5'd6, 27'h000002b2, 32'h00000400,
  1'd1,  5'd17, 27'h0000001c, 5'd0, 27'h00000102, 5'd18, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000346, 5'd1, 27'h0000033e, 5'd26, 27'h000000e8, 32'h00000400,
  1'd1,  5'd16, 27'h00000161, 5'd15, 27'h0000006e, 5'd0, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e0, 5'd15, 27'h000000f9, 5'd10, 27'h00000342, 32'h00000400,
  1'd1,  5'd19, 27'h0000018b, 5'd12, 27'h000000a6, 5'd22, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000015f, 5'd25, 27'h0000011b, 5'd3, 27'h000000c3, 32'h00000400,
  1'd1,  5'd16, 27'h000002e0, 5'd24, 27'h00000059, 5'd12, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001b, 5'd25, 27'h00000176, 5'd25, 27'h000000d1, 32'h00000400,
  1'd1,  5'd30, 27'h000001f1, 5'd1, 27'h0000014e, 5'd1, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000272, 5'd1, 27'h0000004a, 5'd15, 27'h00000147, 32'h00000400,
  1'd1,  5'd27, 27'h000003be, 5'd2, 27'h00000088, 5'd22, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000021, 5'd13, 27'h00000025, 5'd4, 27'h0000020d, 32'h00000400,
  1'd1,  5'd28, 27'h00000124, 5'd10, 27'h00000333, 5'd15, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000019c, 5'd11, 27'h00000199, 5'd20, 27'h000002ae, 32'h00000400,
  1'd1,  5'd30, 27'h000000f5, 5'd24, 27'h00000349, 5'd3, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003e4, 5'd24, 27'h000001a3, 5'd14, 27'h0000006d, 32'h00000400,
  1'd1,  5'd26, 27'h00000028, 5'd21, 27'h000002c9, 5'd24, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000082, 5'd4, 27'h0000032b, 5'd4, 27'h00000162, 32'h00000400,
  1'd1,  5'd5, 27'h00000198, 5'd4, 27'h000000ca, 5'd13, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032d, 5'd3, 27'h0000005f, 5'd20, 27'h000002c7, 32'h00000400,
  1'd1,  5'd6, 27'h000001c9, 5'd13, 27'h000000c8, 5'd5, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000020a, 5'd11, 27'h000002fb, 5'd17, 27'h000001e6, 32'h00000400,
  1'd1,  5'd5, 27'h000003c8, 5'd12, 27'h0000024b, 5'd30, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001b5, 5'd21, 27'h000003aa, 5'd7, 27'h00000088, 32'h00000400,
  1'd1,  5'd8, 27'h000003f5, 5'd24, 27'h00000236, 5'd16, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003cd, 5'd24, 27'h0000017f, 5'd28, 27'h00000114, 32'h00000400,
  1'd1,  5'd19, 27'h000002a9, 5'd1, 27'h0000035a, 5'd4, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029c, 5'd1, 27'h00000126, 5'd12, 27'h0000015a, 32'h00000400,
  1'd1,  5'd17, 27'h000000a6, 5'd1, 27'h000001d0, 5'd24, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000170, 5'd10, 27'h0000022d, 5'd8, 27'h0000008b, 32'h00000400,
  1'd1,  5'd16, 27'h0000007e, 5'd12, 27'h000000c6, 5'd17, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025f, 5'd13, 27'h000000b6, 5'd28, 27'h000002e8, 32'h00000400,
  1'd1,  5'd19, 27'h000002f0, 5'd23, 27'h000002bd, 5'd6, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ac, 5'd23, 27'h000001a5, 5'd18, 27'h00000093, 32'h00000400,
  1'd1,  5'd15, 27'h00000209, 5'd25, 27'h0000034e, 5'd27, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000014d, 5'd3, 27'h00000021, 5'd7, 27'h000000f3, 32'h00000400,
  1'd1,  5'd28, 27'h000002cf, 5'd3, 27'h000000a3, 5'd19, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000196, 5'd4, 27'h000002d1, 5'd27, 27'h0000036c, 32'h00000400,
  1'd1,  5'd26, 27'h000002be, 5'd12, 27'h00000299, 5'd7, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000157, 5'd14, 27'h000002b0, 5'd20, 27'h00000208, 32'h00000400,
  1'd1,  5'd27, 27'h0000015a, 5'd12, 27'h00000204, 5'd27, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003f0, 5'd24, 27'h00000030, 5'd9, 27'h00000176, 32'h00000400,
  1'd1,  5'd27, 27'h000003f8, 5'd22, 27'h00000126, 5'd17, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000021, 5'd23, 27'h0000006c, 5'd26, 27'h0000039f, 32'h00000400,
  1'd1,  5'd5, 27'h00000184, 5'd8, 27'h0000006f, 5'd2, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a9, 5'd8, 27'h00000281, 5'd12, 27'h0000010d, 32'h00000400,
  1'd1,  5'd6, 27'h000003e3, 5'd7, 27'h0000033a, 5'd24, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000012e, 5'd18, 27'h00000194, 5'd3, 27'h0000010b, 32'h00000400,
  1'd1,  5'd10, 27'h000000ad, 5'd19, 27'h000003e2, 5'd13, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003fe, 5'd20, 27'h00000137, 5'd24, 27'h000002e7, 32'h00000400,
  1'd1,  5'd6, 27'h00000356, 5'd28, 27'h00000243, 5'd3, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ab, 5'd27, 27'h00000365, 5'd12, 27'h000002ad, 32'h00000400,
  1'd1,  5'd7, 27'h000001f9, 5'd30, 27'h0000028e, 5'd22, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000035f, 5'd9, 27'h00000337, 5'd0, 27'h00000026, 32'h00000400,
  1'd1,  5'd17, 27'h000002f8, 5'd6, 27'h00000227, 5'd11, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000229, 5'd8, 27'h00000060, 5'd20, 27'h000002c6, 32'h00000400,
  1'd1,  5'd16, 27'h00000395, 5'd19, 27'h0000002b, 5'd1, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e5, 5'd16, 27'h0000005a, 5'd14, 27'h0000016a, 32'h00000400,
  1'd1,  5'd19, 27'h0000008b, 5'd17, 27'h000001fe, 5'd21, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000073, 5'd28, 27'h0000038d, 5'd4, 27'h000003b8, 32'h00000400,
  1'd1,  5'd16, 27'h00000080, 5'd25, 27'h0000035c, 5'd14, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000067, 5'd28, 27'h000000a4, 5'd25, 27'h00000147, 32'h00000400,
  1'd1,  5'd27, 27'h00000103, 5'd7, 27'h00000057, 5'd2, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000374, 5'd5, 27'h0000014d, 5'd13, 27'h000000d5, 32'h00000400,
  1'd1,  5'd27, 27'h00000357, 5'd9, 27'h000001f9, 5'd22, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000172, 5'd20, 27'h000001f0, 5'd2, 27'h0000031a, 32'h00000400,
  1'd1,  5'd26, 27'h000001b5, 5'd19, 27'h000000df, 5'd13, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000377, 5'd18, 27'h000003ac, 5'd23, 27'h0000011c, 32'h00000400,
  1'd1,  5'd29, 27'h000002da, 5'd26, 27'h000002c7, 5'd0, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000336, 5'd25, 27'h000003cd, 5'd15, 27'h000000ce, 32'h00000400,
  1'd1,  5'd27, 27'h000001f8, 5'd29, 27'h00000294, 5'd25, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000037a, 5'd7, 27'h00000304, 5'd8, 27'h00000152, 32'h00000400,
  1'd1,  5'd5, 27'h0000022c, 5'd8, 27'h0000019a, 5'd19, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000242, 5'd9, 27'h00000275, 5'd30, 27'h00000138, 32'h00000400,
  1'd1,  5'd6, 27'h0000038d, 5'd16, 27'h00000311, 5'd7, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003e, 5'd20, 27'h00000117, 5'd17, 27'h00000000, 32'h00000400,
  1'd1,  5'd9, 27'h000003e5, 5'd18, 27'h0000008f, 5'd28, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f9, 5'd28, 27'h000000e2, 5'd6, 27'h0000001a, 32'h00000400,
  1'd1,  5'd6, 27'h000000da, 5'd30, 27'h0000003a, 5'd20, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000041, 5'd30, 27'h00000047, 5'd29, 27'h00000007, 32'h00000400,
  1'd1,  5'd17, 27'h000003bd, 5'd7, 27'h00000245, 5'd7, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e5, 5'd5, 27'h000001f8, 5'd16, 27'h00000242, 32'h00000400,
  1'd1,  5'd18, 27'h0000008c, 5'd7, 27'h00000283, 5'd27, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002e3, 5'd18, 27'h00000028, 5'd6, 27'h000000b1, 32'h00000400,
  1'd1,  5'd18, 27'h000001f7, 5'd17, 27'h000000d0, 5'd18, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f0, 5'd19, 27'h000001ca, 5'd28, 27'h000003e0, 32'h00000400,
  1'd1,  5'd20, 27'h000000dc, 5'd29, 27'h000001c2, 5'd7, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000242, 5'd29, 27'h000003b9, 5'd19, 27'h000002f2, 32'h00000400,
  1'd1,  5'd16, 27'h0000005b, 5'd26, 27'h00000134, 5'd27, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002bd, 5'd10, 27'h00000085, 5'd9, 27'h000001cc, 32'h00000400,
  1'd1,  5'd28, 27'h00000008, 5'd8, 27'h00000299, 5'd17, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000021d, 5'd5, 27'h000000d3, 5'd28, 27'h0000030f, 32'h00000400,
  1'd1,  5'd29, 27'h00000225, 5'd15, 27'h0000020b, 5'd8, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000010f, 5'd18, 27'h00000280, 5'd18, 27'h000000e6, 32'h00000400,
  1'd1,  5'd27, 27'h000001dd, 5'd16, 27'h0000019b, 5'd26, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021f, 5'd29, 27'h000001a7, 5'd7, 27'h000001fc, 32'h00000400,
  1'd1,  5'd27, 27'h000001f4, 5'd27, 27'h00000156, 5'd15, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000256, 5'd27, 27'h0000025d, 5'd28, 27'h0000002d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000245, 5'd2, 27'h000001c0, 5'd2, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000d8, 5'd2, 27'h00000302, 5'd14, 27'h00000134, 32'h00000400,
  1'd1,  5'd4, 27'h000001dd, 5'd3, 27'h000000d1, 5'd21, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002b0, 5'd15, 27'h0000004e, 5'd0, 27'h00000323, 32'h00000400,
  1'd1,  5'd0, 27'h00000196, 5'd10, 27'h000002a8, 5'd14, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000323, 5'd14, 27'h00000179, 5'd23, 27'h00000256, 32'h00000400,
  1'd1,  5'd4, 27'h00000169, 5'd20, 27'h000003dd, 5'd0, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000165, 5'd24, 27'h00000338, 5'd12, 27'h00000381, 32'h00000400,
  1'd1,  5'd0, 27'h000003a9, 5'd20, 27'h000002cb, 5'd22, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ee, 5'd4, 27'h00000266, 5'd2, 27'h0000025a, 32'h00000400,
  1'd1,  5'd12, 27'h00000041, 5'd0, 27'h0000037f, 5'd12, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003c3, 5'd3, 27'h000002df, 5'd24, 27'h0000020b, 32'h00000400,
  1'd1,  5'd13, 27'h00000338, 5'd11, 27'h000001ad, 5'd2, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c5, 5'd10, 27'h000003e7, 5'd12, 27'h000003a7, 32'h00000400,
  1'd1,  5'd12, 27'h00000398, 5'd11, 27'h0000038b, 5'd22, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000260, 5'd22, 27'h00000048, 5'd0, 27'h00000355, 32'h00000400,
  1'd1,  5'd11, 27'h00000328, 5'd23, 27'h000002c8, 5'd13, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000238, 5'd20, 27'h000002e4, 5'd20, 27'h000002ab, 32'h00000400,
  1'd1,  5'd25, 27'h00000093, 5'd1, 27'h00000278, 5'd2, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000016c, 5'd0, 27'h00000026, 5'd11, 27'h000002e6, 32'h00000400,
  1'd1,  5'd25, 27'h000001c0, 5'd0, 27'h000003ec, 5'd20, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002c9, 5'd11, 27'h000002c2, 5'd0, 27'h00000136, 32'h00000400,
  1'd1,  5'd21, 27'h000000be, 5'd11, 27'h000001b2, 5'd14, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000229, 5'd15, 27'h0000014d, 5'd22, 27'h00000351, 32'h00000400,
  1'd1,  5'd25, 27'h0000012e, 5'd24, 27'h00000057, 5'd3, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000372, 5'd23, 27'h000000d8, 5'd13, 27'h0000039d, 32'h00000400,
  1'd1,  5'd24, 27'h00000126, 5'd25, 27'h0000018f, 5'd23, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000169, 5'd4, 27'h000003bb, 5'd7, 27'h00000128, 32'h00000400,
  1'd1,  5'd0, 27'h000003bd, 5'd3, 27'h000000ee, 5'd18, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000329, 5'd3, 27'h00000080, 5'd30, 27'h0000000f, 32'h00000400,
  1'd1,  5'd2, 27'h00000119, 5'd11, 27'h00000159, 5'd5, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000035d, 5'd10, 27'h0000039d, 5'd17, 27'h000002c4, 32'h00000400,
  1'd1,  5'd3, 27'h00000167, 5'd12, 27'h0000029c, 5'd29, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000cc, 5'd21, 27'h00000368, 5'd6, 27'h0000039a, 32'h00000400,
  1'd1,  5'd2, 27'h0000005d, 5'd22, 27'h00000241, 5'd17, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028b, 5'd21, 27'h000002fd, 5'd26, 27'h000000c0, 32'h00000400,
  1'd1,  5'd12, 27'h0000027d, 5'd0, 27'h00000341, 5'd8, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d4, 5'd3, 27'h0000022f, 5'd19, 27'h00000234, 32'h00000400,
  1'd1,  5'd11, 27'h0000025f, 5'd1, 27'h000003e0, 5'd28, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003d6, 5'd14, 27'h0000009a, 5'd8, 27'h000003e8, 32'h00000400,
  1'd1,  5'd11, 27'h00000099, 5'd15, 27'h000000dd, 5'd19, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f4, 5'd12, 27'h00000234, 5'd25, 27'h000003c1, 32'h00000400,
  1'd1,  5'd13, 27'h00000117, 5'd21, 27'h000002f2, 5'd8, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b1, 5'd25, 27'h000001ac, 5'd20, 27'h00000047, 32'h00000400,
  1'd1,  5'd11, 27'h00000043, 5'd24, 27'h0000007e, 5'd27, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000b9, 5'd4, 27'h00000270, 5'd5, 27'h000002b1, 32'h00000400,
  1'd1,  5'd24, 27'h0000006b, 5'd4, 27'h0000025c, 5'd19, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d0, 5'd0, 27'h0000024b, 5'd28, 27'h000001c7, 32'h00000400,
  1'd1,  5'd23, 27'h000001fe, 5'd13, 27'h00000232, 5'd6, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001b7, 5'd12, 27'h00000081, 5'd16, 27'h000000b0, 32'h00000400,
  1'd1,  5'd23, 27'h00000315, 5'd12, 27'h00000239, 5'd26, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001b6, 5'd24, 27'h0000033b, 5'd7, 27'h000002a0, 32'h00000400,
  1'd1,  5'd25, 27'h000002e0, 5'd22, 27'h00000228, 5'd16, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001d9, 5'd21, 27'h000003df, 5'd30, 27'h00000303, 32'h00000400,
  1'd1,  5'd4, 27'h0000025f, 5'd6, 27'h000001ae, 5'd0, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000359, 5'd8, 27'h0000010c, 5'd11, 27'h00000309, 32'h00000400,
  1'd1,  5'd2, 27'h00000196, 5'd6, 27'h000001c1, 5'd24, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b0, 5'd18, 27'h000002d1, 5'd2, 27'h0000017b, 32'h00000400,
  1'd1,  5'd2, 27'h000002d8, 5'd15, 27'h0000022c, 5'd14, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000321, 5'd19, 27'h00000141, 5'd21, 27'h0000033b, 32'h00000400,
  1'd1,  5'd4, 27'h000003fb, 5'd29, 27'h000002c3, 5'd3, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b1, 5'd26, 27'h00000015, 5'd15, 27'h00000141, 32'h00000400,
  1'd1,  5'd0, 27'h000002c2, 5'd30, 27'h00000003, 5'd25, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003cd, 5'd6, 27'h0000027a, 5'd1, 27'h000000ff, 32'h00000400,
  1'd1,  5'd12, 27'h00000161, 5'd6, 27'h00000394, 5'd15, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003bc, 5'd8, 27'h000000cb, 5'd23, 27'h000001fc, 32'h00000400,
  1'd1,  5'd11, 27'h0000033d, 5'd19, 27'h00000102, 5'd3, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000213, 5'd16, 27'h000001ff, 5'd11, 27'h00000184, 32'h00000400,
  1'd1,  5'd12, 27'h00000220, 5'd19, 27'h000002a5, 5'd21, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003da, 5'd28, 27'h000002fe, 5'd2, 27'h00000271, 32'h00000400,
  1'd1,  5'd13, 27'h0000024e, 5'd26, 27'h00000199, 5'd13, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000274, 5'd27, 27'h00000343, 5'd25, 27'h0000002c, 32'h00000400,
  1'd1,  5'd20, 27'h000002ae, 5'd10, 27'h00000090, 5'd0, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000039e, 5'd8, 27'h000000ec, 5'd13, 27'h00000191, 32'h00000400,
  1'd1,  5'd24, 27'h00000114, 5'd6, 27'h000001c1, 5'd24, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002be, 5'd16, 27'h000002fe, 5'd2, 27'h0000022e, 32'h00000400,
  1'd1,  5'd22, 27'h000002a3, 5'd19, 27'h000002f2, 5'd14, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000213, 5'd19, 27'h0000003c, 5'd24, 27'h00000370, 32'h00000400,
  1'd1,  5'd22, 27'h00000061, 5'd26, 27'h0000038f, 5'd3, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000041, 5'd29, 27'h0000011d, 5'd12, 27'h0000003c, 32'h00000400,
  1'd1,  5'd21, 27'h00000348, 5'd29, 27'h000003cc, 5'd21, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000035b, 5'd9, 27'h00000080, 5'd6, 27'h000003b5, 32'h00000400,
  1'd1,  5'd1, 27'h000001d9, 5'd5, 27'h000003a3, 5'd18, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000045, 5'd7, 27'h00000322, 5'd28, 27'h00000248, 32'h00000400,
  1'd1,  5'd3, 27'h000003bd, 5'd18, 27'h00000045, 5'd5, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002e2, 5'd18, 27'h00000258, 5'd20, 27'h00000080, 32'h00000400,
  1'd1,  5'd0, 27'h000002a1, 5'd16, 27'h0000012f, 5'd28, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b9, 5'd27, 27'h00000210, 5'd9, 27'h0000021d, 32'h00000400,
  1'd1,  5'd0, 27'h000000d9, 5'd26, 27'h0000016f, 5'd20, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000296, 5'd27, 27'h00000342, 5'd26, 27'h000002b3, 32'h00000400,
  1'd1,  5'd13, 27'h000000e2, 5'd6, 27'h00000023, 5'd8, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000222, 5'd9, 27'h000001b2, 5'd20, 27'h00000008, 32'h00000400,
  1'd1,  5'd11, 27'h0000034c, 5'd9, 27'h000002cd, 5'd28, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000215, 5'd19, 27'h0000018e, 5'd9, 27'h000000e8, 32'h00000400,
  1'd1,  5'd15, 27'h0000011c, 5'd16, 27'h00000035, 5'd17, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000320, 5'd17, 27'h00000016, 5'd25, 27'h000003e4, 32'h00000400,
  1'd1,  5'd14, 27'h0000017d, 5'd27, 27'h000002b3, 5'd5, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ae, 5'd25, 27'h00000382, 5'd18, 27'h000000a1, 32'h00000400,
  1'd1,  5'd12, 27'h000001cc, 5'd29, 27'h0000015d, 5'd28, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003e8, 5'd5, 27'h000002b0, 5'd6, 27'h00000152, 32'h00000400,
  1'd1,  5'd22, 27'h0000023c, 5'd9, 27'h000003ee, 5'd18, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000036f, 5'd6, 27'h00000350, 5'd29, 27'h00000022, 32'h00000400,
  1'd1,  5'd21, 27'h000000a9, 5'd16, 27'h000003ea, 5'd9, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000ce, 5'd17, 27'h0000020f, 5'd18, 27'h00000046, 32'h00000400,
  1'd1,  5'd23, 27'h000001ef, 5'd19, 27'h00000366, 5'd30, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000178, 5'd25, 27'h0000039d, 5'd8, 27'h000002e9, 32'h00000400,
  1'd1,  5'd23, 27'h0000003b, 5'd28, 27'h00000282, 5'd17, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000037e, 5'd27, 27'h000001d6, 5'd28, 27'h0000013f, 32'h00000400,
  1'd1,  5'd8, 27'h00000073, 5'd3, 27'h000003a6, 5'd10, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b3, 5'd4, 27'h0000027c, 5'd19, 27'h00000281, 32'h00000400,
  1'd1,  5'd8, 27'h00000384, 5'd1, 27'h00000282, 5'd28, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000003f, 5'd12, 27'h000002ed, 5'd2, 27'h000002b3, 32'h00000400,
  1'd1,  5'd6, 27'h000002c8, 5'd15, 27'h000001db, 5'd11, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d7, 5'd12, 27'h000000d8, 5'd23, 27'h000002e8, 32'h00000400,
  1'd1,  5'd9, 27'h0000022d, 5'd23, 27'h0000039d, 5'd1, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000031d, 5'd23, 27'h000002e8, 5'd10, 27'h000003c8, 32'h00000400,
  1'd1,  5'd9, 27'h0000019e, 5'd22, 27'h00000291, 5'd25, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000ca, 5'd2, 27'h00000194, 5'd9, 27'h000003b1, 32'h00000400,
  1'd1,  5'd19, 27'h000000b5, 5'd1, 27'h0000010c, 5'd20, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003a6, 5'd0, 27'h000003ce, 5'd27, 27'h000003df, 32'h00000400,
  1'd1,  5'd19, 27'h0000015d, 5'd12, 27'h000003ee, 5'd3, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002dd, 5'd11, 27'h00000100, 5'd11, 27'h00000018, 32'h00000400,
  1'd1,  5'd17, 27'h0000008b, 5'd14, 27'h00000162, 5'd25, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000024c, 5'd23, 27'h000001c9, 5'd2, 27'h00000072, 32'h00000400,
  1'd1,  5'd17, 27'h00000344, 5'd22, 27'h00000091, 5'd12, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d1, 5'd22, 27'h0000035d, 5'd25, 27'h00000195, 32'h00000400,
  1'd1,  5'd27, 27'h000000b3, 5'd3, 27'h00000214, 5'd0, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000216, 5'd2, 27'h00000160, 5'd13, 27'h000003b2, 32'h00000400,
  1'd1,  5'd27, 27'h0000019a, 5'd3, 27'h000003a9, 5'd22, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000eb, 5'd10, 27'h0000023e, 5'd3, 27'h00000142, 32'h00000400,
  1'd1,  5'd29, 27'h00000309, 5'd13, 27'h000002d7, 5'd10, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007b, 5'd12, 27'h000002e7, 5'd24, 27'h000002b3, 32'h00000400,
  1'd1,  5'd30, 27'h0000034c, 5'd22, 27'h00000345, 5'd3, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a5, 5'd25, 27'h000000f9, 5'd13, 27'h00000148, 32'h00000400,
  1'd1,  5'd29, 27'h00000134, 5'd21, 27'h000003bc, 5'd23, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a2, 5'd2, 27'h000000d6, 5'd3, 27'h00000108, 32'h00000400,
  1'd1,  5'd8, 27'h00000016, 5'd0, 27'h0000033b, 5'd14, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003fc, 5'd5, 27'h00000053, 5'd20, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h0000014f, 5'd14, 27'h000002e1, 5'd8, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a7, 5'd14, 27'h00000304, 5'd16, 27'h0000033c, 32'h00000400,
  1'd1,  5'd8, 27'h000003df, 5'd12, 27'h000000bb, 5'd26, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000244, 5'd22, 27'h000002e1, 5'd8, 27'h000000ff, 32'h00000400,
  1'd1,  5'd8, 27'h00000114, 5'd24, 27'h000003d7, 5'd17, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003e8, 5'd24, 27'h00000057, 5'd28, 27'h0000024c, 32'h00000400,
  1'd1,  5'd19, 27'h00000033, 5'd3, 27'h000003b0, 5'd4, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001f3, 5'd4, 27'h00000184, 5'd13, 27'h00000203, 32'h00000400,
  1'd1,  5'd19, 27'h00000091, 5'd1, 27'h000003ad, 5'd23, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000000, 5'd12, 27'h00000042, 5'd7, 27'h0000033b, 32'h00000400,
  1'd1,  5'd16, 27'h000002b6, 5'd12, 27'h0000036a, 5'd18, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000022e, 5'd13, 27'h000001b5, 5'd26, 27'h00000028, 32'h00000400,
  1'd1,  5'd19, 27'h000002f5, 5'd21, 27'h000000eb, 5'd9, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000395, 5'd24, 27'h0000016e, 5'd17, 27'h0000037b, 32'h00000400,
  1'd1,  5'd16, 27'h000002ef, 5'd22, 27'h00000240, 5'd26, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000015d, 5'd0, 27'h0000014c, 5'd7, 27'h000002f5, 32'h00000400,
  1'd1,  5'd29, 27'h000002c2, 5'd4, 27'h00000295, 5'd15, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000055, 5'd2, 27'h0000017c, 5'd25, 27'h00000364, 32'h00000400,
  1'd1,  5'd26, 27'h00000093, 5'd15, 27'h00000035, 5'd6, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001fb, 5'd10, 27'h000002ce, 5'd20, 27'h00000149, 32'h00000400,
  1'd1,  5'd28, 27'h000001e3, 5'd12, 27'h000003e8, 5'd28, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000039, 5'd24, 27'h0000008b, 5'd10, 27'h00000146, 32'h00000400,
  1'd1,  5'd27, 27'h00000253, 5'd24, 27'h00000305, 5'd17, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000cb, 5'd20, 27'h00000346, 5'd29, 27'h00000064, 32'h00000400,
  1'd1,  5'd6, 27'h00000082, 5'd9, 27'h000001f3, 5'd2, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000209, 5'd10, 27'h00000070, 5'd14, 27'h00000116, 32'h00000400,
  1'd1,  5'd7, 27'h00000253, 5'd7, 27'h00000179, 5'd22, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000af, 5'd17, 27'h0000015a, 5'd4, 27'h00000090, 32'h00000400,
  1'd1,  5'd10, 27'h00000058, 5'd17, 27'h000000e7, 5'd11, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000291, 5'd16, 27'h00000091, 5'd22, 27'h0000027a, 32'h00000400,
  1'd1,  5'd7, 27'h00000170, 5'd28, 27'h00000117, 5'd3, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c1, 5'd28, 27'h000001d5, 5'd12, 27'h000002f6, 32'h00000400,
  1'd1,  5'd6, 27'h000002b3, 5'd26, 27'h00000265, 5'd24, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000222, 5'd5, 27'h00000289, 5'd0, 27'h0000025e, 32'h00000400,
  1'd1,  5'd15, 27'h0000023a, 5'd7, 27'h000001c5, 5'd14, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000269, 5'd9, 27'h00000022, 5'd21, 27'h00000070, 32'h00000400,
  1'd1,  5'd20, 27'h000000aa, 5'd20, 27'h00000067, 5'd2, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000037a, 5'd15, 27'h000002da, 5'd11, 27'h00000391, 32'h00000400,
  1'd1,  5'd18, 27'h000000eb, 5'd20, 27'h000001a7, 5'd21, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c8, 5'd28, 27'h0000039a, 5'd3, 27'h000002bc, 32'h00000400,
  1'd1,  5'd16, 27'h000003a4, 5'd27, 27'h000002c8, 5'd10, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000179, 5'd26, 27'h00000081, 5'd23, 27'h000002d0, 32'h00000400,
  1'd1,  5'd26, 27'h0000020d, 5'd6, 27'h000000ef, 5'd5, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000185, 5'd5, 27'h000001dd, 5'd14, 27'h000001ca, 32'h00000400,
  1'd1,  5'd29, 27'h000000a4, 5'd9, 27'h000001ee, 5'd24, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000022c, 5'd19, 27'h0000004d, 5'd4, 27'h0000029e, 32'h00000400,
  1'd1,  5'd26, 27'h000000d9, 5'd16, 27'h00000259, 5'd12, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000006b, 5'd16, 27'h0000011d, 5'd25, 27'h0000022d, 32'h00000400,
  1'd1,  5'd26, 27'h00000240, 5'd29, 27'h00000196, 5'd2, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012b, 5'd27, 27'h000000a9, 5'd12, 27'h00000350, 32'h00000400,
  1'd1,  5'd29, 27'h00000221, 5'd29, 27'h000001ca, 5'd23, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000347, 5'd6, 27'h000002d0, 5'd5, 27'h00000132, 32'h00000400,
  1'd1,  5'd8, 27'h0000021a, 5'd10, 27'h0000014b, 5'd19, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000004b, 5'd5, 27'h00000286, 5'd30, 27'h0000037e, 32'h00000400,
  1'd1,  5'd9, 27'h000002ea, 5'd20, 27'h000000b1, 5'd5, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002de, 5'd15, 27'h00000369, 5'd19, 27'h00000246, 32'h00000400,
  1'd1,  5'd9, 27'h00000300, 5'd16, 27'h000002df, 5'd26, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000246, 5'd29, 27'h00000030, 5'd7, 27'h00000360, 32'h00000400,
  1'd1,  5'd6, 27'h00000008, 5'd29, 27'h00000219, 5'd17, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000144, 5'd27, 27'h00000132, 5'd29, 27'h00000035, 32'h00000400,
  1'd1,  5'd18, 27'h000000d8, 5'd10, 27'h000000cb, 5'd5, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000021, 5'd8, 27'h000003ec, 5'd16, 27'h000001e7, 32'h00000400,
  1'd1,  5'd17, 27'h00000079, 5'd8, 27'h00000355, 5'd28, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025c, 5'd18, 27'h000000e6, 5'd8, 27'h000003b2, 32'h00000400,
  1'd1,  5'd16, 27'h00000140, 5'd16, 27'h0000008c, 5'd15, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021d, 5'd18, 27'h000003a4, 5'd29, 27'h0000001b, 32'h00000400,
  1'd1,  5'd19, 27'h000003ee, 5'd28, 27'h00000236, 5'd6, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a8, 5'd28, 27'h000000f3, 5'd17, 27'h000003ee, 32'h00000400,
  1'd1,  5'd20, 27'h00000016, 5'd28, 27'h000002cd, 5'd29, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001a1, 5'd6, 27'h0000026b, 5'd7, 27'h0000009b, 32'h00000400,
  1'd1,  5'd27, 27'h000001a4, 5'd7, 27'h00000251, 5'd17, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000052, 5'd9, 27'h000003a9, 5'd26, 27'h000000fe, 32'h00000400,
  1'd1,  5'd29, 27'h00000133, 5'd18, 27'h000003c3, 5'd10, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003cc, 5'd15, 27'h0000037d, 5'd15, 27'h00000398, 32'h00000400,
  1'd1,  5'd26, 27'h000000fc, 5'd20, 27'h00000092, 5'd28, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000130, 5'd28, 27'h00000099, 5'd9, 27'h0000036e, 32'h00000400,
  1'd1,  5'd28, 27'h00000289, 5'd30, 27'h00000233, 5'd16, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000006, 5'd27, 27'h000003f3, 5'd27, 27'h000001f9, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000378, 5'd2, 27'h000000f7, 5'd0, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000034a, 5'd3, 27'h000001d4, 5'd14, 27'h0000031e, 32'h00000400,
  1'd1,  5'd3, 27'h0000007e, 5'd2, 27'h0000034d, 5'd25, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a7, 5'd13, 27'h000000fe, 5'd3, 27'h00000070, 32'h00000400,
  1'd1,  5'd4, 27'h000001ff, 5'd15, 27'h0000001e, 5'd10, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000033d, 5'd11, 27'h000002d2, 5'd21, 27'h00000338, 32'h00000400,
  1'd1,  5'd0, 27'h000003c0, 5'd24, 27'h000003c9, 5'd1, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000322, 5'd24, 27'h000000aa, 5'd13, 27'h000002c1, 32'h00000400,
  1'd1,  5'd2, 27'h00000110, 5'd23, 27'h000002df, 5'd22, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000290, 5'd3, 27'h0000017f, 5'd0, 27'h00000216, 32'h00000400,
  1'd1,  5'd14, 27'h0000028a, 5'd3, 27'h0000029b, 5'd14, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000012a, 5'd1, 27'h0000019a, 5'd22, 27'h000003ab, 32'h00000400,
  1'd1,  5'd12, 27'h000002b4, 5'd14, 27'h000003ad, 5'd3, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000206, 5'd12, 27'h00000231, 5'd11, 27'h00000330, 32'h00000400,
  1'd1,  5'd13, 27'h00000325, 5'd15, 27'h00000025, 5'd21, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000382, 5'd21, 27'h000001a7, 5'd4, 27'h0000023a, 32'h00000400,
  1'd1,  5'd10, 27'h0000034e, 5'd24, 27'h00000235, 5'd12, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000354, 5'd22, 27'h00000070, 5'd23, 27'h000003d9, 32'h00000400,
  1'd1,  5'd23, 27'h0000020b, 5'd3, 27'h000000b5, 5'd0, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000342, 5'd1, 27'h00000036, 5'd15, 27'h000001d5, 32'h00000400,
  1'd1,  5'd22, 27'h0000034a, 5'd2, 27'h00000212, 5'd21, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000011, 5'd15, 27'h000001b4, 5'd3, 27'h00000382, 32'h00000400,
  1'd1,  5'd24, 27'h0000036f, 5'd14, 27'h000002b7, 5'd14, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ea, 5'd11, 27'h00000109, 5'd24, 27'h000001c0, 32'h00000400,
  1'd1,  5'd20, 27'h000003b5, 5'd22, 27'h000000c7, 5'd1, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000248, 5'd24, 27'h0000006b, 5'd12, 27'h0000015e, 32'h00000400,
  1'd1,  5'd22, 27'h000003ea, 5'd20, 27'h000003b7, 5'd24, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000019f, 5'd2, 27'h000003e1, 5'd8, 27'h00000362, 32'h00000400,
  1'd1,  5'd1, 27'h000002be, 5'd1, 27'h000002fd, 5'd18, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000034f, 5'd4, 27'h00000232, 5'd27, 27'h00000246, 32'h00000400,
  1'd1,  5'd3, 27'h00000091, 5'd12, 27'h000003f1, 5'd6, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003f1, 5'd15, 27'h000001d3, 5'd20, 27'h0000003a, 32'h00000400,
  1'd1,  5'd2, 27'h00000345, 5'd13, 27'h00000223, 5'd27, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001e1, 5'd20, 27'h000002dc, 5'd8, 27'h00000107, 32'h00000400,
  1'd1,  5'd3, 27'h00000187, 5'd24, 27'h00000077, 5'd15, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000112, 5'd21, 27'h0000009e, 5'd28, 27'h0000000f, 32'h00000400,
  1'd1,  5'd13, 27'h000001c6, 5'd5, 27'h00000046, 5'd7, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003c1, 5'd0, 27'h000002a3, 5'd18, 27'h0000004e, 32'h00000400,
  1'd1,  5'd12, 27'h0000014a, 5'd2, 27'h000003cb, 5'd27, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000359, 5'd14, 27'h00000269, 5'd5, 27'h00000133, 32'h00000400,
  1'd1,  5'd15, 27'h00000052, 5'd10, 27'h000003c6, 5'd18, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000013a, 5'd10, 27'h000003ee, 5'd29, 27'h000002d8, 32'h00000400,
  1'd1,  5'd10, 27'h00000179, 5'd22, 27'h000003db, 5'd7, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001cf, 5'd22, 27'h0000029f, 5'd15, 27'h000002bf, 32'h00000400,
  1'd1,  5'd14, 27'h00000131, 5'd23, 27'h000003ff, 5'd28, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000027f, 5'd4, 27'h0000027b, 5'd5, 27'h0000036f, 32'h00000400,
  1'd1,  5'd22, 27'h0000037a, 5'd2, 27'h000003a0, 5'd17, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000240, 5'd1, 27'h00000010, 5'd26, 27'h0000028e, 32'h00000400,
  1'd1,  5'd21, 27'h00000089, 5'd11, 27'h000003e6, 5'd9, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ca, 5'd13, 27'h0000034e, 5'd15, 27'h0000024a, 32'h00000400,
  1'd1,  5'd25, 27'h00000010, 5'd11, 27'h000001e2, 5'd26, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000160, 5'd22, 27'h0000012d, 5'd5, 27'h00000269, 32'h00000400,
  1'd1,  5'd24, 27'h0000024b, 5'd21, 27'h0000032b, 5'd15, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b8, 5'd23, 27'h0000018f, 5'd30, 27'h000003e5, 32'h00000400,
  1'd1,  5'd3, 27'h00000329, 5'd6, 27'h00000008, 5'd4, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a7, 5'd9, 27'h00000038, 5'd14, 27'h000000ff, 32'h00000400,
  1'd1,  5'd1, 27'h000002af, 5'd8, 27'h00000108, 5'd24, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000189, 5'd16, 27'h000000bd, 5'd4, 27'h000002ca, 32'h00000400,
  1'd1,  5'd2, 27'h00000369, 5'd19, 27'h000003d4, 5'd13, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000014d, 5'd16, 27'h000002e1, 5'd21, 27'h00000108, 32'h00000400,
  1'd1,  5'd2, 27'h0000003d, 5'd25, 27'h000003e5, 5'd1, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000012f, 5'd26, 27'h00000048, 5'd14, 27'h00000248, 32'h00000400,
  1'd1,  5'd1, 27'h00000141, 5'd28, 27'h00000297, 5'd21, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002a2, 5'd6, 27'h0000019b, 5'd2, 27'h0000009d, 32'h00000400,
  1'd1,  5'd14, 27'h0000007d, 5'd5, 27'h0000021f, 5'd14, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001da, 5'd6, 27'h000003cf, 5'd20, 27'h0000031c, 32'h00000400,
  1'd1,  5'd12, 27'h0000016b, 5'd20, 27'h00000164, 5'd2, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b6, 5'd16, 27'h000002ad, 5'd12, 27'h0000030f, 32'h00000400,
  1'd1,  5'd11, 27'h00000387, 5'd15, 27'h00000248, 5'd21, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000375, 5'd26, 27'h000001eb, 5'd2, 27'h00000169, 32'h00000400,
  1'd1,  5'd11, 27'h00000345, 5'd29, 27'h00000245, 5'd13, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a7, 5'd27, 27'h00000352, 5'd24, 27'h00000063, 32'h00000400,
  1'd1,  5'd24, 27'h0000035f, 5'd7, 27'h00000171, 5'd1, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002fc, 5'd6, 27'h00000010, 5'd14, 27'h00000251, 32'h00000400,
  1'd1,  5'd24, 27'h000001e6, 5'd6, 27'h00000176, 5'd25, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003dd, 5'd16, 27'h00000095, 5'd0, 27'h0000017d, 32'h00000400,
  1'd1,  5'd22, 27'h00000107, 5'd15, 27'h00000298, 5'd12, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000313, 5'd19, 27'h0000004a, 5'd22, 27'h000001d4, 32'h00000400,
  1'd1,  5'd25, 27'h000001c9, 5'd28, 27'h000001cc, 5'd1, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000098, 5'd25, 27'h0000038f, 5'd14, 27'h0000020e, 32'h00000400,
  1'd1,  5'd22, 27'h0000019e, 5'd26, 27'h000001e0, 5'd20, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001fd, 5'd9, 27'h00000292, 5'd7, 27'h000002a8, 32'h00000400,
  1'd1,  5'd4, 27'h00000166, 5'd8, 27'h00000126, 5'd19, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000002d, 5'd6, 27'h000001c8, 5'd28, 27'h00000278, 32'h00000400,
  1'd1,  5'd2, 27'h0000014b, 5'd18, 27'h00000090, 5'd8, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000271, 5'd20, 27'h000000b7, 5'd16, 27'h000001c1, 32'h00000400,
  1'd1,  5'd1, 27'h0000008c, 5'd16, 27'h00000170, 5'd29, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000013b, 5'd25, 27'h000003a0, 5'd8, 27'h000000b5, 32'h00000400,
  1'd1,  5'd0, 27'h000001cf, 5'd29, 27'h0000025f, 5'd20, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001cc, 5'd26, 27'h000003b2, 5'd30, 27'h00000106, 32'h00000400,
  1'd1,  5'd12, 27'h00000155, 5'd8, 27'h000000ed, 5'd5, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000030a, 5'd5, 27'h00000145, 5'd18, 27'h00000373, 32'h00000400,
  1'd1,  5'd14, 27'h00000368, 5'd8, 27'h000000e2, 5'd26, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000000d, 5'd17, 27'h00000314, 5'd9, 27'h000002a2, 32'h00000400,
  1'd1,  5'd14, 27'h00000365, 5'd17, 27'h0000029f, 5'd19, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000171, 5'd19, 27'h0000019b, 5'd26, 27'h0000025c, 32'h00000400,
  1'd1,  5'd12, 27'h000003d8, 5'd30, 27'h00000336, 5'd8, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003db, 5'd28, 27'h000003ff, 5'd16, 27'h00000277, 32'h00000400,
  1'd1,  5'd14, 27'h0000035b, 5'd27, 27'h000001ae, 5'd25, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006a, 5'd6, 27'h0000012b, 5'd6, 27'h000003ac, 32'h00000400,
  1'd1,  5'd22, 27'h0000024a, 5'd9, 27'h000002f6, 5'd18, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000016a, 5'd8, 27'h00000354, 5'd30, 27'h00000049, 32'h00000400,
  1'd1,  5'd24, 27'h000002ff, 5'd19, 27'h000001ce, 5'd5, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000024, 5'd17, 27'h00000372, 5'd18, 27'h0000031b, 32'h00000400,
  1'd1,  5'd21, 27'h000000de, 5'd17, 27'h0000017e, 5'd28, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000027c, 5'd30, 27'h0000005c, 5'd5, 27'h00000257, 32'h00000400,
  1'd1,  5'd24, 27'h000000d8, 5'd29, 27'h00000305, 5'd20, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000023b, 5'd27, 27'h000001b5, 5'd28, 27'h000000ed, 32'h00000400,
  1'd1,  5'd6, 27'h00000050, 5'd4, 27'h000001df, 5'd6, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000072, 5'd2, 27'h0000034d, 5'd18, 27'h000003a3, 32'h00000400,
  1'd1,  5'd8, 27'h000002a3, 5'd0, 27'h00000400, 5'd26, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000196, 5'd15, 27'h000000b0, 5'd0, 27'h00000157, 32'h00000400,
  1'd1,  5'd7, 27'h00000106, 5'd15, 27'h00000074, 5'd13, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ec, 5'd13, 27'h000000bb, 5'd24, 27'h000002bb, 32'h00000400,
  1'd1,  5'd9, 27'h000001f8, 5'd25, 27'h0000025e, 5'd0, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000243, 5'd21, 27'h0000025b, 5'd14, 27'h00000350, 32'h00000400,
  1'd1,  5'd6, 27'h00000207, 5'd23, 27'h0000015d, 5'd21, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000025e, 5'd0, 27'h0000013d, 5'd6, 27'h00000137, 32'h00000400,
  1'd1,  5'd18, 27'h00000381, 5'd1, 27'h000001da, 5'd18, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c1, 5'd4, 27'h00000318, 5'd29, 27'h000003f6, 32'h00000400,
  1'd1,  5'd20, 27'h000000a5, 5'd15, 27'h000001ba, 5'd3, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001bd, 5'd14, 27'h000003bd, 5'd14, 27'h000003c6, 32'h00000400,
  1'd1,  5'd16, 27'h0000016a, 5'd13, 27'h00000115, 5'd21, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000000f, 5'd24, 27'h00000299, 5'd1, 27'h00000105, 32'h00000400,
  1'd1,  5'd15, 27'h000003cb, 5'd22, 27'h00000322, 5'd12, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000175, 5'd21, 27'h00000396, 5'd23, 27'h00000088, 32'h00000400,
  1'd1,  5'd29, 27'h0000034e, 5'd3, 27'h00000164, 5'd2, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000f0, 5'd4, 27'h00000139, 5'd15, 27'h0000011b, 32'h00000400,
  1'd1,  5'd26, 27'h000000a6, 5'd5, 27'h00000096, 5'd23, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000007e, 5'd12, 27'h0000027d, 5'd1, 27'h000001a8, 32'h00000400,
  1'd1,  5'd26, 27'h0000030c, 5'd14, 27'h0000009e, 5'd14, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000033e, 5'd12, 27'h000001a8, 5'd22, 27'h000000e6, 32'h00000400,
  1'd1,  5'd29, 27'h00000139, 5'd22, 27'h00000319, 5'd4, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002b6, 5'd21, 27'h00000209, 5'd12, 27'h000003bf, 32'h00000400,
  1'd1,  5'd27, 27'h00000169, 5'd21, 27'h000002b7, 5'd25, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000204, 5'd0, 27'h00000251, 5'd0, 27'h00000140, 32'h00000400,
  1'd1,  5'd9, 27'h00000047, 5'd5, 27'h00000007, 5'd13, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003cf, 5'd4, 27'h00000077, 5'd23, 27'h00000089, 32'h00000400,
  1'd1,  5'd7, 27'h000000e7, 5'd13, 27'h0000011a, 5'd9, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000046, 5'd11, 27'h00000118, 5'd15, 27'h0000033e, 32'h00000400,
  1'd1,  5'd8, 27'h0000014f, 5'd12, 27'h0000005d, 5'd30, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000003d, 5'd20, 27'h0000034d, 5'd6, 27'h00000076, 32'h00000400,
  1'd1,  5'd10, 27'h0000008a, 5'd22, 27'h0000035d, 5'd19, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000bb, 5'd23, 27'h00000118, 5'd28, 27'h0000023d, 32'h00000400,
  1'd1,  5'd16, 27'h00000102, 5'd3, 27'h000001bb, 5'd4, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000031c, 5'd0, 27'h000001be, 5'd14, 27'h00000117, 32'h00000400,
  1'd1,  5'd19, 27'h0000037d, 5'd2, 27'h0000024c, 5'd22, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000008d, 5'd14, 27'h0000031b, 5'd5, 27'h000001ac, 32'h00000400,
  1'd1,  5'd16, 27'h0000029e, 5'd15, 27'h000001d7, 5'd16, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000023e, 5'd13, 27'h00000128, 5'd30, 27'h00000153, 32'h00000400,
  1'd1,  5'd20, 27'h00000071, 5'd21, 27'h00000154, 5'd8, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001d3, 5'd25, 27'h0000014c, 5'd17, 27'h0000007f, 32'h00000400,
  1'd1,  5'd18, 27'h00000139, 5'd22, 27'h000002a4, 5'd28, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e7, 5'd3, 27'h00000113, 5'd6, 27'h0000038c, 32'h00000400,
  1'd1,  5'd29, 27'h000001db, 5'd3, 27'h0000011c, 5'd16, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000236, 5'd0, 27'h000002c1, 5'd26, 27'h0000035d, 32'h00000400,
  1'd1,  5'd30, 27'h00000226, 5'd15, 27'h00000032, 5'd9, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000000c, 5'd13, 27'h00000122, 5'd16, 27'h000001b1, 32'h00000400,
  1'd1,  5'd27, 27'h00000030, 5'd14, 27'h00000268, 5'd25, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003e2, 5'd25, 27'h000000c3, 5'd8, 27'h00000305, 32'h00000400,
  1'd1,  5'd29, 27'h00000111, 5'd25, 27'h00000040, 5'd15, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000027d, 5'd20, 27'h000003a1, 5'd30, 27'h000002df, 32'h00000400,
  1'd1,  5'd10, 27'h00000071, 5'd9, 27'h0000039d, 5'd4, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002dc, 5'd6, 27'h000001ec, 5'd14, 27'h00000067, 32'h00000400,
  1'd1,  5'd8, 27'h00000375, 5'd9, 27'h00000077, 5'd20, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ab, 5'd17, 27'h000003c9, 5'd0, 27'h00000194, 32'h00000400,
  1'd1,  5'd5, 27'h0000033d, 5'd17, 27'h00000273, 5'd12, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000204, 5'd17, 27'h0000030b, 5'd21, 27'h00000157, 32'h00000400,
  1'd1,  5'd7, 27'h00000037, 5'd27, 27'h00000192, 5'd2, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d2, 5'd30, 27'h000001c7, 5'd14, 27'h0000026f, 32'h00000400,
  1'd1,  5'd8, 27'h00000386, 5'd26, 27'h0000038e, 5'd25, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000222, 5'd9, 27'h00000008, 5'd4, 27'h00000334, 32'h00000400,
  1'd1,  5'd20, 27'h00000233, 5'd9, 27'h000003cb, 5'd13, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ca, 5'd5, 27'h000000dc, 5'd24, 27'h000001ed, 32'h00000400,
  1'd1,  5'd17, 27'h00000130, 5'd17, 27'h00000383, 5'd0, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000018f, 5'd18, 27'h00000152, 5'd10, 27'h000002b4, 32'h00000400,
  1'd1,  5'd16, 27'h00000349, 5'd17, 27'h000000ca, 5'd24, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000216, 5'd29, 27'h00000202, 5'd0, 27'h000001b3, 32'h00000400,
  1'd1,  5'd19, 27'h00000329, 5'd27, 27'h000001bd, 5'd11, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c3, 5'd26, 27'h00000166, 5'd23, 27'h0000035d, 32'h00000400,
  1'd1,  5'd29, 27'h0000035f, 5'd9, 27'h000001e3, 5'd0, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000031c, 5'd9, 27'h000000d7, 5'd10, 27'h00000277, 32'h00000400,
  1'd1,  5'd28, 27'h000003d7, 5'd6, 27'h000003f4, 5'd20, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003b4, 5'd15, 27'h00000225, 5'd1, 27'h00000151, 32'h00000400,
  1'd1,  5'd26, 27'h000003be, 5'd17, 27'h00000104, 5'd11, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003d6, 5'd17, 27'h00000193, 5'd23, 27'h00000190, 32'h00000400,
  1'd1,  5'd29, 27'h000001cf, 5'd26, 27'h0000007f, 5'd0, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000de, 5'd30, 27'h000003de, 5'd10, 27'h0000034b, 32'h00000400,
  1'd1,  5'd28, 27'h00000112, 5'd28, 27'h0000029e, 5'd22, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000bb, 5'd5, 27'h000000d3, 5'd8, 27'h0000007f, 32'h00000400,
  1'd1,  5'd6, 27'h000000e1, 5'd8, 27'h000003c4, 5'd18, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001fc, 5'd9, 27'h00000314, 5'd28, 27'h00000132, 32'h00000400,
  1'd1,  5'd6, 27'h000001e4, 5'd17, 27'h0000016b, 5'd6, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000185, 5'd17, 27'h0000007f, 5'd18, 27'h00000358, 32'h00000400,
  1'd1,  5'd7, 27'h000002f7, 5'd19, 27'h0000028d, 5'd30, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000214, 5'd30, 27'h0000019f, 5'd5, 27'h000001e6, 32'h00000400,
  1'd1,  5'd7, 27'h000003fd, 5'd30, 27'h000002b2, 5'd15, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000206, 5'd25, 27'h000003f6, 5'd27, 27'h0000025d, 32'h00000400,
  1'd1,  5'd17, 27'h00000299, 5'd8, 27'h000003ac, 5'd6, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000027c, 5'd5, 27'h00000227, 5'd19, 27'h00000131, 32'h00000400,
  1'd1,  5'd19, 27'h0000035f, 5'd6, 27'h000001f0, 5'd27, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000138, 5'd19, 27'h0000035b, 5'd5, 27'h000003b0, 32'h00000400,
  1'd1,  5'd19, 27'h0000037d, 5'd19, 27'h000003b7, 5'd16, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000239, 5'd20, 27'h000001f9, 5'd29, 27'h000000be, 32'h00000400,
  1'd1,  5'd20, 27'h000001eb, 5'd26, 27'h000001d9, 5'd8, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003da, 5'd26, 27'h0000039b, 5'd17, 27'h000000ea, 32'h00000400,
  1'd1,  5'd20, 27'h00000180, 5'd30, 27'h0000039c, 5'd26, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d8, 5'd9, 27'h000001b2, 5'd8, 27'h000001e5, 32'h00000400,
  1'd1,  5'd26, 27'h0000026d, 5'd7, 27'h000002fb, 5'd19, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000bc, 5'd8, 27'h00000207, 5'd29, 27'h000000c4, 32'h00000400,
  1'd1,  5'd30, 27'h000003eb, 5'd20, 27'h000001e2, 5'd5, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003be, 5'd18, 27'h00000029, 5'd15, 27'h0000029a, 32'h00000400,
  1'd1,  5'd26, 27'h000000f8, 5'd20, 27'h00000012, 5'd29, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a9, 5'd30, 27'h0000031e, 5'd5, 27'h00000346, 32'h00000400,
  1'd1,  5'd28, 27'h000002ec, 5'd26, 27'h0000026c, 5'd17, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000000d, 5'd28, 27'h000003cd, 5'd27, 27'h000003bc, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000192, 5'd4, 27'h00000251, 5'd1, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000018c, 5'd4, 27'h000001e2, 5'd10, 27'h0000030e, 32'h00000400,
  1'd1,  5'd1, 27'h0000005b, 5'd4, 27'h00000369, 5'd24, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000343, 5'd14, 27'h00000074, 5'd3, 27'h000003ac, 32'h00000400,
  1'd1,  5'd2, 27'h000003b6, 5'd10, 27'h0000024e, 5'd10, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000046, 5'd15, 27'h000000f9, 5'd25, 27'h000001a9, 32'h00000400,
  1'd1,  5'd0, 27'h000000cd, 5'd24, 27'h0000023c, 5'd1, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000023b, 5'd21, 27'h00000130, 5'd14, 27'h000000ba, 32'h00000400,
  1'd1,  5'd2, 27'h00000085, 5'd23, 27'h00000145, 5'd22, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000b7, 5'd1, 27'h0000009f, 5'd1, 27'h000002ca, 32'h00000400,
  1'd1,  5'd13, 27'h000002f8, 5'd5, 27'h00000048, 5'd10, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003c3, 5'd4, 27'h00000002, 5'd24, 27'h00000201, 32'h00000400,
  1'd1,  5'd11, 27'h000000b5, 5'd14, 27'h00000278, 5'd2, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f5, 5'd10, 27'h000001e5, 5'd13, 27'h000002bb, 32'h00000400,
  1'd1,  5'd10, 27'h0000029d, 5'd15, 27'h00000024, 5'd21, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000016, 5'd23, 27'h00000281, 5'd2, 27'h0000019c, 32'h00000400,
  1'd1,  5'd13, 27'h00000174, 5'd23, 27'h00000054, 5'd12, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000275, 5'd22, 27'h0000038c, 5'd23, 27'h00000120, 32'h00000400,
  1'd1,  5'd23, 27'h00000392, 5'd0, 27'h00000204, 5'd2, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000327, 5'd4, 27'h0000038c, 5'd12, 27'h000002b4, 32'h00000400,
  1'd1,  5'd21, 27'h00000211, 5'd1, 27'h00000349, 5'd23, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000230, 5'd10, 27'h00000326, 5'd3, 27'h0000033a, 32'h00000400,
  1'd1,  5'd24, 27'h0000033c, 5'd12, 27'h00000048, 5'd14, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c6, 5'd11, 27'h00000177, 5'd24, 27'h000002b5, 32'h00000400,
  1'd1,  5'd22, 27'h000003a2, 5'd21, 27'h00000125, 5'd3, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002e4, 5'd24, 27'h000002c9, 5'd13, 27'h0000000f, 32'h00000400,
  1'd1,  5'd24, 27'h000000b3, 5'd24, 27'h0000032b, 5'd21, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a8, 5'd4, 27'h0000025c, 5'd7, 27'h000002bc, 32'h00000400,
  1'd1,  5'd2, 27'h0000016f, 5'd2, 27'h0000035b, 5'd15, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000160, 5'd4, 27'h0000037d, 5'd28, 27'h000002a6, 32'h00000400,
  1'd1,  5'd1, 27'h0000001c, 5'd13, 27'h00000175, 5'd9, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000057, 5'd14, 27'h000001cb, 5'd19, 27'h0000009d, 32'h00000400,
  1'd1,  5'd1, 27'h0000008c, 5'd11, 27'h0000034f, 5'd28, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000033c, 5'd21, 27'h00000388, 5'd10, 27'h000000a3, 32'h00000400,
  1'd1,  5'd3, 27'h000001ec, 5'd24, 27'h000000da, 5'd17, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000013d, 5'd22, 27'h00000136, 5'd30, 27'h000002e8, 32'h00000400,
  1'd1,  5'd13, 27'h000003ba, 5'd2, 27'h00000210, 5'd7, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002c5, 5'd1, 27'h000003f6, 5'd18, 27'h0000008d, 32'h00000400,
  1'd1,  5'd14, 27'h000001ef, 5'd2, 27'h00000151, 5'd30, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f9, 5'd15, 27'h0000018b, 5'd7, 27'h000003a4, 32'h00000400,
  1'd1,  5'd15, 27'h0000009c, 5'd12, 27'h0000015b, 5'd16, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000030, 5'd12, 27'h00000192, 5'd26, 27'h000000a6, 32'h00000400,
  1'd1,  5'd13, 27'h0000030f, 5'd21, 27'h000003a8, 5'd9, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018b, 5'd22, 27'h0000012f, 5'd18, 27'h000001ce, 32'h00000400,
  1'd1,  5'd14, 27'h000003ee, 5'd23, 27'h00000368, 5'd27, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000035, 5'd0, 27'h0000007a, 5'd6, 27'h00000084, 32'h00000400,
  1'd1,  5'd25, 27'h00000316, 5'd0, 27'h00000005, 5'd17, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000176, 5'd2, 27'h00000262, 5'd30, 27'h00000223, 32'h00000400,
  1'd1,  5'd23, 27'h00000157, 5'd14, 27'h0000029b, 5'd5, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000180, 5'd13, 27'h00000329, 5'd19, 27'h00000051, 32'h00000400,
  1'd1,  5'd25, 27'h00000193, 5'd12, 27'h000001cb, 5'd27, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003c7, 5'd25, 27'h00000235, 5'd10, 27'h0000012e, 32'h00000400,
  1'd1,  5'd21, 27'h000003d7, 5'd24, 27'h000001cb, 5'd16, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001bd, 5'd21, 27'h0000028a, 5'd27, 27'h0000003e, 32'h00000400,
  1'd1,  5'd0, 27'h000000bc, 5'd7, 27'h00000005, 5'd1, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f2, 5'd9, 27'h000002ff, 5'd15, 27'h00000020, 32'h00000400,
  1'd1,  5'd0, 27'h00000318, 5'd9, 27'h00000355, 5'd24, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000033d, 5'd19, 27'h00000233, 5'd4, 27'h000003fc, 32'h00000400,
  1'd1,  5'd0, 27'h000002f5, 5'd18, 27'h000003e0, 5'd10, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002cf, 5'd16, 27'h000002e2, 5'd25, 27'h000000cd, 32'h00000400,
  1'd1,  5'd4, 27'h000003f6, 5'd29, 27'h0000031c, 5'd5, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000082, 5'd30, 27'h00000386, 5'd10, 27'h000002db, 32'h00000400,
  1'd1,  5'd0, 27'h00000266, 5'd26, 27'h000003a3, 5'd21, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001a3, 5'd8, 27'h0000014b, 5'd0, 27'h0000012e, 32'h00000400,
  1'd1,  5'd13, 27'h00000138, 5'd7, 27'h000002cc, 5'd13, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000065, 5'd5, 27'h0000013a, 5'd25, 27'h0000028d, 32'h00000400,
  1'd1,  5'd12, 27'h00000039, 5'd18, 27'h00000105, 5'd0, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f6, 5'd19, 27'h00000392, 5'd14, 27'h00000287, 32'h00000400,
  1'd1,  5'd11, 27'h00000139, 5'd20, 27'h0000029f, 5'd23, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000006e, 5'd27, 27'h000003ad, 5'd1, 27'h000000ec, 32'h00000400,
  1'd1,  5'd11, 27'h00000266, 5'd27, 27'h000003a5, 5'd11, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000025a, 5'd27, 27'h00000226, 5'd25, 27'h00000163, 32'h00000400,
  1'd1,  5'd22, 27'h00000321, 5'd10, 27'h000000d1, 5'd0, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000008a, 5'd9, 27'h000000e7, 5'd10, 27'h000002c6, 32'h00000400,
  1'd1,  5'd23, 27'h0000034e, 5'd7, 27'h00000356, 5'd23, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001a7, 5'd17, 27'h000001ee, 5'd3, 27'h000001a8, 32'h00000400,
  1'd1,  5'd25, 27'h00000147, 5'd19, 27'h00000160, 5'd11, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001c6, 5'd18, 27'h00000317, 5'd25, 27'h00000224, 32'h00000400,
  1'd1,  5'd25, 27'h000000e3, 5'd26, 27'h000002e3, 5'd2, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000074, 5'd30, 27'h00000165, 5'd10, 27'h00000384, 32'h00000400,
  1'd1,  5'd21, 27'h0000008c, 5'd26, 27'h00000197, 5'd24, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000069, 5'd7, 27'h0000000a, 5'd9, 27'h000002cb, 32'h00000400,
  1'd1,  5'd1, 27'h0000039b, 5'd6, 27'h000001de, 5'd20, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d8, 5'd7, 27'h000002ab, 5'd30, 27'h000000fd, 32'h00000400,
  1'd1,  5'd2, 27'h00000128, 5'd16, 27'h00000128, 5'd8, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002e3, 5'd15, 27'h00000247, 5'd18, 27'h0000001d, 32'h00000400,
  1'd1,  5'd4, 27'h000002b7, 5'd16, 27'h0000032d, 5'd30, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000300, 5'd26, 27'h00000237, 5'd6, 27'h00000191, 32'h00000400,
  1'd1,  5'd3, 27'h000000bb, 5'd30, 27'h00000388, 5'd18, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000001b, 5'd27, 27'h000003e7, 5'd28, 27'h000002e0, 32'h00000400,
  1'd1,  5'd11, 27'h000001bb, 5'd6, 27'h00000039, 5'd8, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000370, 5'd9, 27'h000003b7, 5'd18, 27'h0000033c, 32'h00000400,
  1'd1,  5'd10, 27'h000003e8, 5'd10, 27'h00000115, 5'd26, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000009c, 5'd16, 27'h00000294, 5'd5, 27'h000003bf, 32'h00000400,
  1'd1,  5'd12, 27'h000001e1, 5'd16, 27'h00000337, 5'd16, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000154, 5'd19, 27'h000000c4, 5'd29, 27'h0000017f, 32'h00000400,
  1'd1,  5'd14, 27'h000001ae, 5'd29, 27'h000001a2, 5'd5, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e5, 5'd28, 27'h0000034e, 5'd17, 27'h000002b2, 32'h00000400,
  1'd1,  5'd12, 27'h00000296, 5'd27, 27'h00000251, 5'd28, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000371, 5'd8, 27'h0000032e, 5'd9, 27'h000001d4, 32'h00000400,
  1'd1,  5'd24, 27'h0000015c, 5'd6, 27'h0000022d, 5'd18, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000060, 5'd5, 27'h000003b1, 5'd27, 27'h000001bf, 32'h00000400,
  1'd1,  5'd20, 27'h00000372, 5'd18, 27'h0000025f, 5'd5, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000116, 5'd15, 27'h000002e4, 5'd18, 27'h0000013d, 32'h00000400,
  1'd1,  5'd23, 27'h0000022d, 5'd19, 27'h000000ce, 5'd30, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000201, 5'd30, 27'h0000035b, 5'd6, 27'h000002bd, 32'h00000400,
  1'd1,  5'd24, 27'h0000033f, 5'd30, 27'h000001da, 5'd17, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000158, 5'd30, 27'h00000038, 5'd29, 27'h00000359, 32'h00000400,
  1'd1,  5'd9, 27'h000000ac, 5'd1, 27'h00000153, 5'd7, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000315, 5'd4, 27'h000001d7, 5'd19, 27'h000001a9, 32'h00000400,
  1'd1,  5'd6, 27'h0000030a, 5'd2, 27'h00000189, 5'd30, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000269, 5'd13, 27'h00000390, 5'd2, 27'h000003e4, 32'h00000400,
  1'd1,  5'd10, 27'h00000049, 5'd12, 27'h00000232, 5'd10, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000309, 5'd10, 27'h000001cd, 5'd25, 27'h00000296, 32'h00000400,
  1'd1,  5'd8, 27'h00000107, 5'd22, 27'h000001ae, 5'd1, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000027f, 5'd21, 27'h0000020d, 5'd10, 27'h00000229, 32'h00000400,
  1'd1,  5'd9, 27'h000000cf, 5'd25, 27'h00000312, 5'd21, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001d5, 5'd0, 27'h00000288, 5'd8, 27'h00000363, 32'h00000400,
  1'd1,  5'd20, 27'h000000ac, 5'd0, 27'h000000ca, 5'd17, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000337, 5'd2, 27'h000001ad, 5'd25, 27'h00000366, 32'h00000400,
  1'd1,  5'd18, 27'h0000004b, 5'd13, 27'h0000014a, 5'd0, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b8, 5'd11, 27'h00000297, 5'd12, 27'h0000027d, 32'h00000400,
  1'd1,  5'd18, 27'h000002a9, 5'd10, 27'h00000248, 5'd24, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000025e, 5'd23, 27'h00000243, 5'd0, 27'h000002f9, 32'h00000400,
  1'd1,  5'd15, 27'h0000033f, 5'd23, 27'h000001ba, 5'd14, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002d, 5'd24, 27'h000001fe, 5'd25, 27'h000001dd, 32'h00000400,
  1'd1,  5'd27, 27'h000002f1, 5'd4, 27'h00000341, 5'd5, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000181, 5'd0, 27'h00000250, 5'd12, 27'h000002d6, 32'h00000400,
  1'd1,  5'd27, 27'h000002b7, 5'd3, 27'h000001ae, 5'd21, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b9, 5'd10, 27'h000001fd, 5'd3, 27'h00000005, 32'h00000400,
  1'd1,  5'd30, 27'h00000135, 5'd12, 27'h0000017c, 5'd13, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000039d, 5'd12, 27'h00000166, 5'd25, 27'h0000021d, 32'h00000400,
  1'd1,  5'd28, 27'h000003dd, 5'd25, 27'h00000088, 5'd0, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000347, 5'd24, 27'h00000042, 5'd11, 27'h00000398, 32'h00000400,
  1'd1,  5'd28, 27'h00000024, 5'd22, 27'h000003be, 5'd22, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000213, 5'd3, 27'h0000016d, 5'd2, 27'h00000060, 32'h00000400,
  1'd1,  5'd8, 27'h00000121, 5'd1, 27'h00000334, 5'd11, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e7, 5'd2, 27'h000001ef, 5'd23, 27'h0000031a, 32'h00000400,
  1'd1,  5'd6, 27'h00000331, 5'd12, 27'h000001c9, 5'd5, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000029e, 5'd11, 27'h000003ee, 5'd16, 27'h00000208, 32'h00000400,
  1'd1,  5'd6, 27'h000003c8, 5'd14, 27'h000003e1, 5'd26, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000091, 5'd24, 27'h00000223, 5'd9, 27'h0000007c, 32'h00000400,
  1'd1,  5'd9, 27'h00000337, 5'd23, 27'h0000037e, 5'd16, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000029c, 5'd21, 27'h000003a4, 5'd26, 27'h0000037d, 32'h00000400,
  1'd1,  5'd16, 27'h00000348, 5'd2, 27'h00000077, 5'd1, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002be, 5'd1, 27'h00000294, 5'd12, 27'h0000006f, 32'h00000400,
  1'd1,  5'd16, 27'h000003e1, 5'd0, 27'h00000075, 5'd21, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003b9, 5'd13, 27'h00000057, 5'd7, 27'h000003de, 32'h00000400,
  1'd1,  5'd15, 27'h0000028a, 5'd12, 27'h000001d3, 5'd18, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000004f, 5'd13, 27'h0000006b, 5'd30, 27'h0000022b, 32'h00000400,
  1'd1,  5'd20, 27'h00000213, 5'd21, 27'h00000057, 5'd7, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e1, 5'd24, 27'h000000d1, 5'd17, 27'h00000083, 32'h00000400,
  1'd1,  5'd15, 27'h0000033d, 5'd20, 27'h000003da, 5'd29, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000184, 5'd0, 27'h0000028b, 5'd5, 27'h000000c6, 32'h00000400,
  1'd1,  5'd29, 27'h0000016b, 5'd4, 27'h000002c4, 5'd19, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000bf, 5'd5, 27'h00000098, 5'd29, 27'h00000156, 32'h00000400,
  1'd1,  5'd26, 27'h00000010, 5'd14, 27'h000003dd, 5'd7, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000249, 5'd10, 27'h00000309, 5'd16, 27'h00000337, 32'h00000400,
  1'd1,  5'd30, 27'h00000369, 5'd12, 27'h000003e4, 5'd29, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000035d, 5'd20, 27'h000003d0, 5'd5, 27'h000000d3, 32'h00000400,
  1'd1,  5'd26, 27'h000003d4, 5'd21, 27'h000000a6, 5'd15, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e5, 5'd21, 27'h00000214, 5'd26, 27'h000000fd, 32'h00000400,
  1'd1,  5'd10, 27'h0000004a, 5'd7, 27'h000000c7, 5'd4, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000317, 5'd8, 27'h00000241, 5'd11, 27'h00000086, 32'h00000400,
  1'd1,  5'd7, 27'h000002d2, 5'd6, 27'h0000014d, 5'd24, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000007d, 5'd20, 27'h00000232, 5'd4, 27'h00000129, 32'h00000400,
  1'd1,  5'd5, 27'h000000f4, 5'd16, 27'h000003c8, 5'd14, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000102, 5'd16, 27'h00000325, 5'd21, 27'h00000081, 32'h00000400,
  1'd1,  5'd8, 27'h00000191, 5'd30, 27'h00000068, 5'd1, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000071, 5'd26, 27'h00000174, 5'd13, 27'h0000006e, 32'h00000400,
  1'd1,  5'd5, 27'h00000180, 5'd30, 27'h000000f1, 5'd24, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000127, 5'd9, 27'h0000023d, 5'd3, 27'h000003fa, 32'h00000400,
  1'd1,  5'd16, 27'h0000022f, 5'd9, 27'h000003be, 5'd14, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000026, 5'd7, 27'h00000310, 5'd22, 27'h000001a5, 32'h00000400,
  1'd1,  5'd16, 27'h000000da, 5'd19, 27'h00000179, 5'd4, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000102, 5'd18, 27'h000003fc, 5'd13, 27'h000000be, 32'h00000400,
  1'd1,  5'd18, 27'h00000003, 5'd20, 27'h0000027d, 5'd21, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c7, 5'd27, 27'h000002d2, 5'd3, 27'h0000032b, 32'h00000400,
  1'd1,  5'd19, 27'h00000218, 5'd26, 27'h00000114, 5'd11, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000009d, 5'd29, 27'h00000136, 5'd21, 27'h00000236, 32'h00000400,
  1'd1,  5'd26, 27'h000000f2, 5'd10, 27'h0000004c, 5'd1, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000bc, 5'd9, 27'h000000fe, 5'd13, 27'h0000022e, 32'h00000400,
  1'd1,  5'd28, 27'h0000021d, 5'd7, 27'h000003bf, 5'd24, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003ab, 5'd18, 27'h00000386, 5'd0, 27'h00000299, 32'h00000400,
  1'd1,  5'd28, 27'h000000d0, 5'd17, 27'h00000242, 5'd11, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002be, 5'd17, 27'h00000023, 5'd20, 27'h00000320, 32'h00000400,
  1'd1,  5'd26, 27'h0000003c, 5'd28, 27'h00000086, 5'd4, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000a0, 5'd29, 27'h000000e2, 5'd12, 27'h000003de, 32'h00000400,
  1'd1,  5'd26, 27'h000000a3, 5'd25, 27'h000003e8, 5'd23, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000044, 5'd5, 27'h00000212, 5'd5, 27'h00000371, 32'h00000400,
  1'd1,  5'd9, 27'h00000141, 5'd5, 27'h00000400, 5'd16, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000100, 5'd6, 27'h000003f3, 5'd30, 27'h00000344, 32'h00000400,
  1'd1,  5'd9, 27'h000002ee, 5'd17, 27'h0000009b, 5'd10, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ac, 5'd17, 27'h0000003d, 5'd17, 27'h00000024, 32'h00000400,
  1'd1,  5'd9, 27'h000002ab, 5'd20, 27'h00000257, 5'd29, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000199, 5'd27, 27'h00000261, 5'd8, 27'h00000385, 32'h00000400,
  1'd1,  5'd5, 27'h000000ed, 5'd30, 27'h000003eb, 5'd16, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000016e, 5'd28, 27'h000003e7, 5'd28, 27'h000003e0, 32'h00000400,
  1'd1,  5'd16, 27'h0000010d, 5'd6, 27'h000003df, 5'd7, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000156, 5'd9, 27'h000000a1, 5'd16, 27'h000003d9, 32'h00000400,
  1'd1,  5'd20, 27'h00000290, 5'd9, 27'h0000016c, 5'd29, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ee, 5'd17, 27'h00000091, 5'd7, 27'h000003b3, 32'h00000400,
  1'd1,  5'd18, 27'h00000013, 5'd20, 27'h000001a8, 5'd15, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000151, 5'd15, 27'h000003d1, 5'd25, 27'h00000379, 32'h00000400,
  1'd1,  5'd20, 27'h0000018c, 5'd27, 27'h00000068, 5'd9, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003a5, 5'd29, 27'h0000004f, 5'd17, 27'h0000011e, 32'h00000400,
  1'd1,  5'd17, 27'h000001da, 5'd29, 27'h00000083, 5'd28, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000194, 5'd6, 27'h0000032f, 5'd6, 27'h0000009e, 32'h00000400,
  1'd1,  5'd30, 27'h0000007f, 5'd7, 27'h00000296, 5'd17, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000037c, 5'd8, 27'h000002ca, 5'd27, 27'h0000031f, 32'h00000400,
  1'd1,  5'd30, 27'h00000223, 5'd18, 27'h0000014d, 5'd10, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000006b, 5'd17, 27'h00000042, 5'd16, 27'h0000013f, 32'h00000400,
  1'd1,  5'd30, 27'h00000137, 5'd16, 27'h00000365, 5'd28, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000025f, 5'd27, 27'h00000292, 5'd7, 27'h00000131, 32'h00000400,
  1'd1,  5'd27, 27'h000001bf, 5'd25, 27'h000003e0, 5'd15, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001c7, 5'd26, 27'h000003b5, 5'd28, 27'h0000024e, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000322, 5'd2, 27'h00000135, 5'd3, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000032, 5'd0, 27'h000001a5, 5'd12, 27'h0000029f, 32'h00000400,
  1'd1,  5'd4, 27'h000002b4, 5'd1, 27'h00000340, 5'd25, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038b, 5'd14, 27'h00000108, 5'd2, 27'h000000a7, 32'h00000400,
  1'd1,  5'd2, 27'h00000311, 5'd12, 27'h0000010b, 5'd14, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000025f, 5'd15, 27'h00000105, 5'd21, 27'h00000255, 32'h00000400,
  1'd1,  5'd4, 27'h0000009e, 5'd22, 27'h00000317, 5'd1, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b8, 5'd21, 27'h000000c2, 5'd11, 27'h00000219, 32'h00000400,
  1'd1,  5'd0, 27'h00000191, 5'd23, 27'h000000c1, 5'd25, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ba, 5'd4, 27'h00000157, 5'd4, 27'h000001a2, 32'h00000400,
  1'd1,  5'd15, 27'h00000139, 5'd4, 27'h000001a9, 5'd10, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002c7, 5'd1, 27'h0000039c, 5'd24, 27'h00000205, 32'h00000400,
  1'd1,  5'd14, 27'h000003f5, 5'd12, 27'h000000cc, 5'd2, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001cb, 5'd14, 27'h00000194, 5'd13, 27'h000001c5, 32'h00000400,
  1'd1,  5'd10, 27'h00000390, 5'd12, 27'h00000135, 5'd25, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d3, 5'd24, 27'h000003ec, 5'd0, 27'h000001ca, 32'h00000400,
  1'd1,  5'd11, 27'h0000034a, 5'd20, 27'h00000314, 5'd12, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000017a, 5'd23, 27'h00000069, 5'd24, 27'h000003e0, 32'h00000400,
  1'd1,  5'd25, 27'h00000180, 5'd3, 27'h0000007f, 5'd0, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000297, 5'd2, 27'h00000229, 5'd14, 27'h000003c0, 32'h00000400,
  1'd1,  5'd20, 27'h000002b4, 5'd0, 27'h00000291, 5'd24, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001e2, 5'd12, 27'h0000036c, 5'd2, 27'h000000ea, 32'h00000400,
  1'd1,  5'd24, 27'h00000243, 5'd11, 27'h0000024c, 5'd10, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000019b, 5'd13, 27'h00000186, 5'd24, 27'h000001dc, 32'h00000400,
  1'd1,  5'd25, 27'h00000239, 5'd21, 27'h000002b4, 5'd4, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000014, 5'd23, 27'h000000fc, 5'd12, 27'h00000302, 32'h00000400,
  1'd1,  5'd23, 27'h0000001e, 5'd24, 27'h00000305, 5'd21, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002aa, 5'd3, 27'h000001d1, 5'd5, 27'h000002b6, 32'h00000400,
  1'd1,  5'd4, 27'h00000113, 5'd3, 27'h0000002c, 5'd17, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000181, 5'd4, 27'h000001ea, 5'd27, 27'h00000296, 32'h00000400,
  1'd1,  5'd3, 27'h00000150, 5'd15, 27'h000000e1, 5'd10, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002b8, 5'd15, 27'h00000031, 5'd17, 27'h00000347, 32'h00000400,
  1'd1,  5'd1, 27'h0000014c, 5'd15, 27'h00000188, 5'd26, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000377, 5'd22, 27'h000000c5, 5'd9, 27'h000000fd, 32'h00000400,
  1'd1,  5'd0, 27'h000002fa, 5'd24, 27'h000002a7, 5'd16, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000375, 5'd23, 27'h000000c2, 5'd28, 27'h000000d1, 32'h00000400,
  1'd1,  5'd14, 27'h0000014f, 5'd4, 27'h000003bd, 5'd7, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000028a, 5'd1, 27'h000001a6, 5'd17, 27'h0000019d, 32'h00000400,
  1'd1,  5'd10, 27'h00000251, 5'd3, 27'h000001da, 5'd30, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000015d, 5'd10, 27'h0000020f, 5'd8, 27'h00000084, 32'h00000400,
  1'd1,  5'd13, 27'h00000243, 5'd13, 27'h0000015b, 5'd18, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000016c, 5'd10, 27'h000003b2, 5'd27, 27'h000001cc, 32'h00000400,
  1'd1,  5'd11, 27'h00000400, 5'd25, 27'h000000cf, 5'd10, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000136, 5'd24, 27'h0000037c, 5'd20, 27'h000001c0, 32'h00000400,
  1'd1,  5'd14, 27'h000002b9, 5'd25, 27'h00000145, 5'd30, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002f0, 5'd3, 27'h000001ba, 5'd6, 27'h000003cb, 32'h00000400,
  1'd1,  5'd25, 27'h000001ca, 5'd0, 27'h00000225, 5'd16, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000109, 5'd0, 27'h00000251, 5'd26, 27'h0000027c, 32'h00000400,
  1'd1,  5'd25, 27'h0000017d, 5'd13, 27'h000002b4, 5'd9, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ac, 5'd15, 27'h000000c9, 5'd19, 27'h000000e2, 32'h00000400,
  1'd1,  5'd21, 27'h00000300, 5'd11, 27'h00000075, 5'd27, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000205, 5'd23, 27'h00000191, 5'd7, 27'h0000013e, 32'h00000400,
  1'd1,  5'd22, 27'h000001a8, 5'd23, 27'h000002a9, 5'd16, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001be, 5'd23, 27'h0000036a, 5'd26, 27'h00000033, 32'h00000400,
  1'd1,  5'd1, 27'h0000027e, 5'd7, 27'h00000183, 5'd0, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000036, 5'd8, 27'h00000105, 5'd10, 27'h00000273, 32'h00000400,
  1'd1,  5'd2, 27'h000002ee, 5'd8, 27'h00000101, 5'd23, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000084, 5'd18, 27'h0000010d, 5'd4, 27'h00000343, 32'h00000400,
  1'd1,  5'd2, 27'h000002b7, 5'd15, 27'h000003a2, 5'd10, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000208, 5'd18, 27'h00000123, 5'd25, 27'h00000268, 32'h00000400,
  1'd1,  5'd4, 27'h0000032e, 5'd26, 27'h00000324, 5'd0, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000296, 5'd26, 27'h0000033b, 5'd13, 27'h000003d4, 32'h00000400,
  1'd1,  5'd2, 27'h0000021d, 5'd29, 27'h000000ea, 5'd25, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000243, 5'd6, 27'h00000359, 5'd4, 27'h00000184, 32'h00000400,
  1'd1,  5'd12, 27'h000000f0, 5'd8, 27'h000002d2, 5'd13, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001d9, 5'd5, 27'h000000b8, 5'd24, 27'h000002cd, 32'h00000400,
  1'd1,  5'd11, 27'h000000a0, 5'd15, 27'h000002a7, 5'd4, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000196, 5'd18, 27'h0000000c, 5'd14, 27'h00000018, 32'h00000400,
  1'd1,  5'd14, 27'h00000147, 5'd15, 27'h000002e2, 5'd20, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002bc, 5'd30, 27'h000001d6, 5'd3, 27'h00000385, 32'h00000400,
  1'd1,  5'd14, 27'h00000378, 5'd30, 27'h000003f1, 5'd15, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000383, 5'd30, 27'h00000030, 5'd25, 27'h000002bb, 32'h00000400,
  1'd1,  5'd23, 27'h00000320, 5'd7, 27'h00000076, 5'd1, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001ab, 5'd5, 27'h00000367, 5'd12, 27'h000001e8, 32'h00000400,
  1'd1,  5'd25, 27'h00000147, 5'd9, 27'h00000236, 5'd25, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000103, 5'd17, 27'h000002ee, 5'd3, 27'h0000006f, 32'h00000400,
  1'd1,  5'd21, 27'h000002c7, 5'd15, 27'h00000231, 5'd12, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e2, 5'd20, 27'h0000008f, 5'd25, 27'h00000290, 32'h00000400,
  1'd1,  5'd25, 27'h000002c7, 5'd27, 27'h00000290, 5'd1, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000023c, 5'd26, 27'h0000027f, 5'd10, 27'h000002a6, 32'h00000400,
  1'd1,  5'd24, 27'h000002a7, 5'd27, 27'h000003a8, 5'd21, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000021, 5'd9, 27'h00000076, 5'd6, 27'h000002dd, 32'h00000400,
  1'd1,  5'd4, 27'h000003ae, 5'd8, 27'h0000017a, 5'd17, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ca, 5'd10, 27'h0000011c, 5'd26, 27'h000002f4, 32'h00000400,
  1'd1,  5'd0, 27'h000003cc, 5'd15, 27'h000002ee, 5'd6, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000036e, 5'd16, 27'h000003f6, 5'd20, 27'h0000013e, 32'h00000400,
  1'd1,  5'd0, 27'h0000014b, 5'd17, 27'h00000164, 5'd29, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000253, 5'd30, 27'h000001c5, 5'd8, 27'h000001f2, 32'h00000400,
  1'd1,  5'd1, 27'h0000015c, 5'd29, 27'h000001c0, 5'd18, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000004c, 5'd30, 27'h00000058, 5'd30, 27'h000000d9, 32'h00000400,
  1'd1,  5'd14, 27'h00000050, 5'd7, 27'h000000f9, 5'd5, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000018e, 5'd9, 27'h00000338, 5'd16, 27'h000003b6, 32'h00000400,
  1'd1,  5'd11, 27'h000000d2, 5'd8, 27'h0000015d, 5'd26, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f0, 5'd15, 27'h000003de, 5'd5, 27'h000002aa, 32'h00000400,
  1'd1,  5'd14, 27'h0000021b, 5'd19, 27'h00000158, 5'd16, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000063, 5'd18, 27'h00000045, 5'd26, 27'h000003f6, 32'h00000400,
  1'd1,  5'd14, 27'h00000185, 5'd26, 27'h0000011f, 5'd7, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f9, 5'd29, 27'h000001b1, 5'd17, 27'h0000001e, 32'h00000400,
  1'd1,  5'd12, 27'h000000a2, 5'd28, 27'h00000248, 5'd27, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000009d, 5'd9, 27'h000001a7, 5'd7, 27'h000001b4, 32'h00000400,
  1'd1,  5'd22, 27'h00000309, 5'd7, 27'h000001dd, 5'd17, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001e6, 5'd5, 27'h00000332, 5'd26, 27'h0000004d, 32'h00000400,
  1'd1,  5'd25, 27'h00000209, 5'd18, 27'h000003d0, 5'd7, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000021e, 5'd16, 27'h000000e4, 5'd18, 27'h00000027, 32'h00000400,
  1'd1,  5'd20, 27'h00000395, 5'd19, 27'h000002fb, 5'd30, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000aa, 5'd27, 27'h000002f5, 5'd8, 27'h0000008a, 32'h00000400,
  1'd1,  5'd24, 27'h0000024a, 5'd28, 27'h000003a6, 5'd17, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000008e, 5'd27, 27'h0000008e, 5'd29, 27'h00000035, 32'h00000400,
  1'd1,  5'd6, 27'h000000cf, 5'd2, 27'h000001a1, 5'd8, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000020c, 5'd3, 27'h00000102, 5'd19, 27'h00000215, 32'h00000400,
  1'd1,  5'd5, 27'h000001ac, 5'd2, 27'h000002bd, 5'd29, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000032d, 5'd15, 27'h000001f9, 5'd0, 27'h00000032, 32'h00000400,
  1'd1,  5'd6, 27'h000002a9, 5'd13, 27'h0000010c, 5'd15, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000338, 5'd11, 27'h000002e5, 5'd24, 27'h0000027c, 32'h00000400,
  1'd1,  5'd8, 27'h0000004d, 5'd22, 27'h00000241, 5'd1, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023f, 5'd22, 27'h0000000d, 5'd11, 27'h00000165, 32'h00000400,
  1'd1,  5'd8, 27'h0000028e, 5'd25, 27'h0000004f, 5'd21, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000251, 5'd4, 27'h00000332, 5'd5, 27'h000000fc, 32'h00000400,
  1'd1,  5'd18, 27'h000000a5, 5'd4, 27'h0000035f, 5'd18, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000012b, 5'd2, 27'h000001c6, 5'd27, 27'h00000024, 32'h00000400,
  1'd1,  5'd19, 27'h00000236, 5'd15, 27'h0000009f, 5'd4, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000024e, 5'd11, 27'h000003c8, 5'd11, 27'h000003da, 32'h00000400,
  1'd1,  5'd18, 27'h00000207, 5'd13, 27'h000001ac, 5'd24, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000003e, 5'd24, 27'h000002a9, 5'd2, 27'h0000001b, 32'h00000400,
  1'd1,  5'd19, 27'h000000af, 5'd21, 27'h000002f7, 5'd10, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000370, 5'd21, 27'h00000216, 5'd23, 27'h00000276, 32'h00000400,
  1'd1,  5'd28, 27'h000000cb, 5'd3, 27'h00000384, 5'd3, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001f7, 5'd2, 27'h00000285, 5'd14, 27'h000000ce, 32'h00000400,
  1'd1,  5'd30, 27'h000001b1, 5'd4, 27'h0000018b, 5'd23, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003fe, 5'd13, 27'h000000c3, 5'd4, 27'h000000d4, 32'h00000400,
  1'd1,  5'd30, 27'h0000016b, 5'd13, 27'h00000080, 5'd11, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001db, 5'd15, 27'h0000007f, 5'd20, 27'h000002fd, 32'h00000400,
  1'd1,  5'd26, 27'h000000d9, 5'd24, 27'h000002ec, 5'd2, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000002f, 5'd20, 27'h00000349, 5'd14, 27'h000002fc, 32'h00000400,
  1'd1,  5'd25, 27'h00000375, 5'd25, 27'h0000029f, 5'd23, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a2, 5'd0, 27'h00000188, 5'd0, 27'h000002a1, 32'h00000400,
  1'd1,  5'd7, 27'h00000305, 5'd0, 27'h000002ac, 5'd12, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000026e, 5'd0, 27'h000003c6, 5'd25, 27'h00000269, 32'h00000400,
  1'd1,  5'd7, 27'h00000254, 5'd12, 27'h00000164, 5'd10, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000245, 5'd11, 27'h000002d2, 5'd19, 27'h000001dd, 32'h00000400,
  1'd1,  5'd5, 27'h000001a9, 5'd15, 27'h00000102, 5'd27, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000d8, 5'd23, 27'h000001ef, 5'd9, 27'h0000039e, 32'h00000400,
  1'd1,  5'd7, 27'h000003e1, 5'd24, 27'h000000e1, 5'd17, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002fb, 5'd20, 27'h00000310, 5'd26, 27'h0000036b, 32'h00000400,
  1'd1,  5'd17, 27'h000003fb, 5'd0, 27'h000003b8, 5'd0, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002f1, 5'd0, 27'h00000041, 5'd13, 27'h00000099, 32'h00000400,
  1'd1,  5'd16, 27'h0000006a, 5'd0, 27'h000003ec, 5'd24, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ae, 5'd14, 27'h0000027d, 5'd5, 27'h000003e2, 32'h00000400,
  1'd1,  5'd19, 27'h00000162, 5'd13, 27'h000000ae, 5'd18, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000006d, 5'd10, 27'h000002fb, 5'd29, 27'h000003e2, 32'h00000400,
  1'd1,  5'd16, 27'h000003ef, 5'd21, 27'h000003a9, 5'd8, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000037a, 5'd21, 27'h000002ae, 5'd15, 27'h000003b1, 32'h00000400,
  1'd1,  5'd15, 27'h00000277, 5'd25, 27'h0000032d, 5'd28, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002db, 5'd4, 27'h000003fc, 5'd5, 27'h00000358, 32'h00000400,
  1'd1,  5'd30, 27'h000002a1, 5'd2, 27'h000002e0, 5'd20, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003fe, 5'd1, 27'h00000224, 5'd28, 27'h0000022f, 32'h00000400,
  1'd1,  5'd29, 27'h000001fc, 5'd14, 27'h000002fb, 5'd8, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000db, 5'd10, 27'h000002b2, 5'd19, 27'h00000043, 32'h00000400,
  1'd1,  5'd27, 27'h0000014b, 5'd11, 27'h0000022f, 5'd28, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000368, 5'd22, 27'h000003d1, 5'd8, 27'h0000009b, 32'h00000400,
  1'd1,  5'd26, 27'h00000043, 5'd23, 27'h00000151, 5'd16, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000039c, 5'd22, 27'h0000038f, 5'd29, 27'h00000171, 32'h00000400,
  1'd1,  5'd7, 27'h000003f8, 5'd9, 27'h00000166, 5'd3, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002d9, 5'd8, 27'h000003e4, 5'd14, 27'h00000316, 32'h00000400,
  1'd1,  5'd7, 27'h0000024e, 5'd9, 27'h00000105, 5'd25, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000151, 5'd20, 27'h000001e1, 5'd4, 27'h00000367, 32'h00000400,
  1'd1,  5'd7, 27'h000003f4, 5'd15, 27'h000002a4, 5'd10, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000194, 5'd17, 27'h00000130, 5'd22, 27'h000001fd, 32'h00000400,
  1'd1,  5'd6, 27'h00000115, 5'd29, 27'h000001f3, 5'd1, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000003e, 5'd27, 27'h00000090, 5'd11, 27'h00000246, 32'h00000400,
  1'd1,  5'd7, 27'h00000342, 5'd26, 27'h00000306, 5'd20, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000260, 5'd7, 27'h000002eb, 5'd4, 27'h0000024b, 32'h00000400,
  1'd1,  5'd17, 27'h00000161, 5'd9, 27'h00000396, 5'd11, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002d7, 5'd6, 27'h000000b0, 5'd21, 27'h00000062, 32'h00000400,
  1'd1,  5'd18, 27'h00000010, 5'd19, 27'h000001e0, 5'd3, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000273, 5'd18, 27'h000001f3, 5'd14, 27'h00000006, 32'h00000400,
  1'd1,  5'd18, 27'h00000159, 5'd16, 27'h000002e9, 5'd21, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001bb, 5'd29, 27'h0000020a, 5'd1, 27'h00000356, 32'h00000400,
  1'd1,  5'd17, 27'h000002bd, 5'd30, 27'h000001e7, 5'd10, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ed, 5'd28, 27'h000000cb, 5'd21, 27'h000002d4, 32'h00000400,
  1'd1,  5'd28, 27'h000000ab, 5'd6, 27'h000002a4, 5'd2, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000206, 5'd7, 27'h00000258, 5'd14, 27'h00000358, 32'h00000400,
  1'd1,  5'd29, 27'h00000260, 5'd9, 27'h000002cb, 5'd22, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000277, 5'd18, 27'h0000031b, 5'd1, 27'h000003eb, 32'h00000400,
  1'd1,  5'd27, 27'h0000004c, 5'd19, 27'h00000227, 5'd12, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000067, 5'd17, 27'h00000047, 5'd21, 27'h000001a2, 32'h00000400,
  1'd1,  5'd29, 27'h0000022d, 5'd27, 27'h00000359, 5'd3, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000035e, 5'd30, 27'h00000012, 5'd10, 27'h000001ef, 32'h00000400,
  1'd1,  5'd27, 27'h00000329, 5'd26, 27'h000001c9, 5'd22, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000373, 5'd9, 27'h0000030f, 5'd6, 27'h00000292, 32'h00000400,
  1'd1,  5'd8, 27'h00000300, 5'd6, 27'h0000012f, 5'd15, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000105, 5'd9, 27'h0000018a, 5'd26, 27'h000000c0, 32'h00000400,
  1'd1,  5'd6, 27'h00000248, 5'd19, 27'h00000322, 5'd9, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000065, 5'd17, 27'h00000208, 5'd17, 27'h0000007c, 32'h00000400,
  1'd1,  5'd5, 27'h0000033e, 5'd16, 27'h0000033d, 5'd29, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000355, 5'd30, 27'h00000285, 5'd8, 27'h0000028a, 32'h00000400,
  1'd1,  5'd9, 27'h00000189, 5'd27, 27'h00000374, 5'd18, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000121, 5'd27, 27'h000002ec, 5'd27, 27'h000002a6, 32'h00000400,
  1'd1,  5'd16, 27'h000001fb, 5'd7, 27'h000000ef, 5'd6, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000132, 5'd7, 27'h00000180, 5'd18, 27'h00000394, 32'h00000400,
  1'd1,  5'd20, 27'h000000a1, 5'd10, 27'h00000103, 5'd26, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001cf, 5'd18, 27'h00000199, 5'd8, 27'h00000199, 32'h00000400,
  1'd1,  5'd18, 27'h000003a6, 5'd15, 27'h00000384, 5'd15, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d5, 5'd20, 27'h0000025f, 5'd27, 27'h0000014e, 32'h00000400,
  1'd1,  5'd15, 27'h0000023b, 5'd26, 27'h0000012d, 5'd7, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034c, 5'd29, 27'h00000236, 5'd19, 27'h000001ed, 32'h00000400,
  1'd1,  5'd20, 27'h00000151, 5'd30, 27'h00000333, 5'd26, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002a5, 5'd6, 27'h0000032b, 5'd9, 27'h000003ca, 32'h00000400,
  1'd1,  5'd29, 27'h000001b0, 5'd5, 27'h0000021b, 5'd17, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000087, 5'd8, 27'h00000278, 5'd26, 27'h00000124, 32'h00000400,
  1'd1,  5'd26, 27'h00000173, 5'd16, 27'h0000032a, 5'd9, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000029a, 5'd18, 27'h000002c7, 5'd18, 27'h00000121, 32'h00000400,
  1'd1,  5'd29, 27'h000003aa, 5'd17, 27'h00000012, 5'd25, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000146, 5'd26, 27'h000001a5, 5'd8, 27'h000003eb, 32'h00000400,
  1'd1,  5'd30, 27'h000002ea, 5'd27, 27'h00000006, 5'd19, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000df, 5'd30, 27'h0000014c, 5'd28, 27'h00000016, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000001be, 5'd0, 27'h000000e6, 5'd4, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000150, 5'd4, 27'h0000009b, 5'd13, 27'h000001a0, 32'h00000400,
  1'd1,  5'd1, 27'h00000172, 5'd2, 27'h0000004f, 5'd21, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b6, 5'd15, 27'h00000127, 5'd4, 27'h00000023, 32'h00000400,
  1'd1,  5'd0, 27'h000002d6, 5'd15, 27'h000000c6, 5'd12, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e5, 5'd10, 27'h00000305, 5'd21, 27'h00000169, 32'h00000400,
  1'd1,  5'd4, 27'h00000270, 5'd24, 27'h00000284, 5'd4, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000085, 5'd22, 27'h000003e0, 5'd14, 27'h0000036d, 32'h00000400,
  1'd1,  5'd5, 27'h00000050, 5'd22, 27'h000002c0, 5'd22, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000012c, 5'd2, 27'h000003c2, 5'd2, 27'h0000017e, 32'h00000400,
  1'd1,  5'd14, 27'h0000014e, 5'd1, 27'h00000270, 5'd12, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000179, 5'd0, 27'h0000000b, 5'd22, 27'h0000037f, 32'h00000400,
  1'd1,  5'd13, 27'h000002c5, 5'd13, 27'h000000e8, 5'd2, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000283, 5'd11, 27'h00000082, 5'd11, 27'h00000334, 32'h00000400,
  1'd1,  5'd10, 27'h0000027c, 5'd11, 27'h000000c8, 5'd25, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000342, 5'd25, 27'h0000007f, 5'd1, 27'h00000004, 32'h00000400,
  1'd1,  5'd14, 27'h0000029f, 5'd23, 27'h0000022f, 5'd11, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000043, 5'd23, 27'h0000025a, 5'd21, 27'h000001aa, 32'h00000400,
  1'd1,  5'd24, 27'h00000174, 5'd2, 27'h0000030c, 5'd0, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000144, 5'd0, 27'h000000c4, 5'd12, 27'h000001cf, 32'h00000400,
  1'd1,  5'd21, 27'h0000026a, 5'd1, 27'h000000e1, 5'd23, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000164, 5'd15, 27'h000000f7, 5'd3, 27'h00000253, 32'h00000400,
  1'd1,  5'd24, 27'h00000375, 5'd14, 27'h00000122, 5'd12, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000027c, 5'd14, 27'h000000fe, 5'd21, 27'h000003a5, 32'h00000400,
  1'd1,  5'd24, 27'h0000017c, 5'd21, 27'h00000222, 5'd0, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000219, 5'd25, 27'h000000d0, 5'd11, 27'h000000eb, 32'h00000400,
  1'd1,  5'd22, 27'h000002f1, 5'd23, 27'h0000003b, 5'd25, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001bb, 5'd4, 27'h0000006e, 5'd8, 27'h00000088, 32'h00000400,
  1'd1,  5'd3, 27'h0000031e, 5'd4, 27'h0000031c, 5'd16, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001a9, 5'd4, 27'h0000011a, 5'd28, 27'h000003f1, 32'h00000400,
  1'd1,  5'd3, 27'h0000000b, 5'd14, 27'h00000400, 5'd8, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f8, 5'd11, 27'h00000246, 5'd16, 27'h00000191, 32'h00000400,
  1'd1,  5'd1, 27'h000001bb, 5'd12, 27'h0000017a, 5'd26, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000281, 5'd23, 27'h00000170, 5'd10, 27'h0000009e, 32'h00000400,
  1'd1,  5'd0, 27'h00000240, 5'd25, 27'h0000017e, 5'd15, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d0, 5'd22, 27'h00000143, 5'd30, 27'h00000211, 32'h00000400,
  1'd1,  5'd11, 27'h0000000f, 5'd4, 27'h00000200, 5'd5, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000279, 5'd1, 27'h0000008e, 5'd15, 27'h000002db, 32'h00000400,
  1'd1,  5'd13, 27'h0000038f, 5'd1, 27'h00000066, 5'd26, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000e1, 5'd13, 27'h000001f2, 5'd7, 27'h000001d0, 32'h00000400,
  1'd1,  5'd13, 27'h0000018d, 5'd11, 27'h000003f3, 5'd18, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000078, 5'd14, 27'h00000017, 5'd28, 27'h000001ed, 32'h00000400,
  1'd1,  5'd14, 27'h0000003c, 5'd21, 27'h00000116, 5'd7, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000001a, 5'd25, 27'h00000025, 5'd20, 27'h00000120, 32'h00000400,
  1'd1,  5'd10, 27'h0000030d, 5'd22, 27'h000003d8, 5'd27, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001f4, 5'd4, 27'h00000055, 5'd8, 27'h0000024c, 32'h00000400,
  1'd1,  5'd21, 27'h00000003, 5'd1, 27'h00000305, 5'd16, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000020a, 5'd4, 27'h000001f1, 5'd28, 27'h0000006d, 32'h00000400,
  1'd1,  5'd24, 27'h0000027d, 5'd14, 27'h00000345, 5'd6, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000140, 5'd14, 27'h00000206, 5'd20, 27'h0000004b, 32'h00000400,
  1'd1,  5'd24, 27'h000002ee, 5'd11, 27'h00000006, 5'd30, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022a, 5'd23, 27'h0000035c, 5'd7, 27'h0000005b, 32'h00000400,
  1'd1,  5'd24, 27'h0000018c, 5'd23, 27'h0000007b, 5'd15, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035f, 5'd22, 27'h00000193, 5'd30, 27'h000003a9, 32'h00000400,
  1'd1,  5'd4, 27'h00000116, 5'd9, 27'h00000185, 5'd2, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000018c, 5'd9, 27'h0000022a, 5'd13, 27'h00000068, 32'h00000400,
  1'd1,  5'd3, 27'h000000d8, 5'd8, 27'h00000357, 5'd21, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000015d, 5'd16, 27'h00000363, 5'd2, 27'h000001c8, 32'h00000400,
  1'd1,  5'd4, 27'h0000009a, 5'd16, 27'h00000352, 5'd13, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001ee, 5'd17, 27'h00000306, 5'd24, 27'h000000ec, 32'h00000400,
  1'd1,  5'd4, 27'h0000020c, 5'd27, 27'h0000015f, 5'd2, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000277, 5'd27, 27'h000002df, 5'd14, 27'h000003fa, 32'h00000400,
  1'd1,  5'd2, 27'h00000133, 5'd27, 27'h000002a5, 5'd20, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000013d, 5'd9, 27'h0000020c, 5'd1, 27'h000002e8, 32'h00000400,
  1'd1,  5'd13, 27'h00000279, 5'd9, 27'h000001a9, 5'd12, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001cd, 5'd9, 27'h000000d8, 5'd25, 27'h00000211, 32'h00000400,
  1'd1,  5'd13, 27'h000002b3, 5'd17, 27'h0000032a, 5'd1, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e2, 5'd19, 27'h00000173, 5'd15, 27'h000001b8, 32'h00000400,
  1'd1,  5'd15, 27'h000000da, 5'd16, 27'h00000290, 5'd25, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000114, 5'd26, 27'h00000229, 5'd4, 27'h000002f6, 32'h00000400,
  1'd1,  5'd10, 27'h00000231, 5'd30, 27'h000003a0, 5'd14, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ec, 5'd27, 27'h000001db, 5'd20, 27'h000003e5, 32'h00000400,
  1'd1,  5'd22, 27'h000003c2, 5'd9, 27'h000002c8, 5'd0, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000296, 5'd9, 27'h00000289, 5'd11, 27'h0000032e, 32'h00000400,
  1'd1,  5'd25, 27'h00000193, 5'd7, 27'h00000012, 5'd25, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000029d, 5'd18, 27'h00000287, 5'd3, 27'h00000084, 32'h00000400,
  1'd1,  5'd22, 27'h00000040, 5'd20, 27'h000000a0, 5'd11, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000036b, 5'd19, 27'h000003bf, 5'd23, 27'h00000140, 32'h00000400,
  1'd1,  5'd20, 27'h000002e4, 5'd26, 27'h00000232, 5'd4, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002e1, 5'd29, 27'h0000039c, 5'd10, 27'h000003fb, 32'h00000400,
  1'd1,  5'd25, 27'h000002b0, 5'd26, 27'h00000182, 5'd25, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000b8, 5'd5, 27'h0000021a, 5'd6, 27'h000001e4, 32'h00000400,
  1'd1,  5'd0, 27'h0000003a, 5'd5, 27'h00000240, 5'd17, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000238, 5'd6, 27'h00000124, 5'd27, 27'h00000313, 32'h00000400,
  1'd1,  5'd0, 27'h000003da, 5'd19, 27'h00000192, 5'd6, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000005c, 5'd15, 27'h0000022c, 5'd16, 27'h00000300, 32'h00000400,
  1'd1,  5'd0, 27'h000003ff, 5'd16, 27'h0000001f, 5'd28, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000115, 5'd29, 27'h000003b6, 5'd5, 27'h000002e5, 32'h00000400,
  1'd1,  5'd0, 27'h00000258, 5'd28, 27'h0000007d, 5'd19, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000024f, 5'd30, 27'h0000029d, 5'd26, 27'h0000005c, 32'h00000400,
  1'd1,  5'd15, 27'h0000001c, 5'd6, 27'h000003f3, 5'd5, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000325, 5'd10, 27'h000000a8, 5'd18, 27'h00000255, 32'h00000400,
  1'd1,  5'd12, 27'h00000223, 5'd5, 27'h000002a3, 5'd28, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000000d, 5'd19, 27'h000003d7, 5'd7, 27'h0000015e, 32'h00000400,
  1'd1,  5'd12, 27'h000002d3, 5'd15, 27'h00000247, 5'd16, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001aa, 5'd18, 27'h0000011f, 5'd28, 27'h00000083, 32'h00000400,
  1'd1,  5'd10, 27'h000003e2, 5'd30, 27'h00000059, 5'd7, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000197, 5'd27, 27'h000002a3, 5'd16, 27'h000002f9, 32'h00000400,
  1'd1,  5'd14, 27'h000003d0, 5'd26, 27'h00000049, 5'd26, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002fc, 5'd7, 27'h000002ee, 5'd7, 27'h00000235, 32'h00000400,
  1'd1,  5'd23, 27'h00000277, 5'd9, 27'h000003ce, 5'd18, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000350, 5'd8, 27'h00000039, 5'd27, 27'h0000027e, 32'h00000400,
  1'd1,  5'd23, 27'h00000143, 5'd19, 27'h00000097, 5'd6, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000263, 5'd18, 27'h000000e0, 5'd18, 27'h00000254, 32'h00000400,
  1'd1,  5'd23, 27'h00000110, 5'd19, 27'h000002b6, 5'd28, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000026d, 5'd25, 27'h00000398, 5'd8, 27'h000002ed, 32'h00000400,
  1'd1,  5'd24, 27'h0000024c, 5'd27, 27'h000003c5, 5'd16, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000005e, 5'd30, 27'h00000172, 5'd28, 27'h0000010e, 32'h00000400,
  1'd1,  5'd5, 27'h000000d5, 5'd3, 27'h0000003a, 5'd5, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000140, 5'd2, 27'h000002d1, 5'd20, 27'h00000281, 32'h00000400,
  1'd1,  5'd8, 27'h0000039f, 5'd1, 27'h00000201, 5'd30, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000185, 5'd15, 27'h00000178, 5'd4, 27'h000002d6, 32'h00000400,
  1'd1,  5'd6, 27'h000000ae, 5'd11, 27'h00000345, 5'd14, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001d5, 5'd14, 27'h0000007f, 5'd20, 27'h00000319, 32'h00000400,
  1'd1,  5'd9, 27'h00000061, 5'd25, 27'h00000096, 5'd1, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000179, 5'd24, 27'h000001ec, 5'd14, 27'h00000310, 32'h00000400,
  1'd1,  5'd8, 27'h0000039d, 5'd20, 27'h000003fa, 5'd25, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002e8, 5'd0, 27'h00000189, 5'd5, 27'h00000106, 32'h00000400,
  1'd1,  5'd18, 27'h0000034f, 5'd4, 27'h000002e6, 5'd17, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021e, 5'd0, 27'h0000012c, 5'd25, 27'h00000359, 32'h00000400,
  1'd1,  5'd15, 27'h000003f7, 5'd12, 27'h0000001a, 5'd4, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000282, 5'd10, 27'h00000313, 5'd10, 27'h000001b0, 32'h00000400,
  1'd1,  5'd17, 27'h00000099, 5'd14, 27'h000003b4, 5'd25, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ea, 5'd24, 27'h0000020a, 5'd0, 27'h000002f6, 32'h00000400,
  1'd1,  5'd18, 27'h000002dd, 5'd23, 27'h00000066, 5'd10, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000010f, 5'd22, 27'h00000236, 5'd24, 27'h000001eb, 32'h00000400,
  1'd1,  5'd30, 27'h00000286, 5'd3, 27'h00000307, 5'd2, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000a6, 5'd2, 27'h00000191, 5'd14, 27'h0000030c, 32'h00000400,
  1'd1,  5'd28, 27'h000000eb, 5'd1, 27'h00000100, 5'd22, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ea, 5'd13, 27'h000002ef, 5'd1, 27'h000002fb, 32'h00000400,
  1'd1,  5'd27, 27'h0000005b, 5'd12, 27'h0000011a, 5'd12, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f3, 5'd13, 27'h000003cb, 5'd23, 27'h00000333, 32'h00000400,
  1'd1,  5'd28, 27'h000002dc, 5'd22, 27'h0000014b, 5'd3, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000032d, 5'd20, 27'h00000391, 5'd10, 27'h00000392, 32'h00000400,
  1'd1,  5'd26, 27'h000003f0, 5'd23, 27'h000002dd, 5'd22, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003eb, 5'd0, 27'h000000cf, 5'd2, 27'h00000154, 32'h00000400,
  1'd1,  5'd8, 27'h000002e7, 5'd4, 27'h0000028b, 5'd13, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000264, 5'd1, 27'h000001b7, 5'd20, 27'h000002f6, 32'h00000400,
  1'd1,  5'd5, 27'h000003c6, 5'd11, 27'h0000030c, 5'd9, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000012, 5'd14, 27'h00000280, 5'd19, 27'h00000056, 32'h00000400,
  1'd1,  5'd5, 27'h0000019b, 5'd12, 27'h000000d4, 5'd29, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003bc, 5'd22, 27'h000003ac, 5'd9, 27'h000001e9, 32'h00000400,
  1'd1,  5'd5, 27'h00000345, 5'd24, 27'h0000011e, 5'd20, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000311, 5'd23, 27'h000000f7, 5'd26, 27'h000002a3, 32'h00000400,
  1'd1,  5'd17, 27'h00000087, 5'd4, 27'h00000391, 5'd4, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000025c, 5'd1, 27'h0000016c, 5'd11, 27'h000003d4, 32'h00000400,
  1'd1,  5'd18, 27'h000001cb, 5'd2, 27'h000000c5, 5'd25, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000298, 5'd11, 27'h000002b3, 5'd8, 27'h000003d2, 32'h00000400,
  1'd1,  5'd20, 27'h000000a2, 5'd10, 27'h000003ac, 5'd20, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000186, 5'd10, 27'h000003a6, 5'd30, 27'h00000378, 32'h00000400,
  1'd1,  5'd17, 27'h000002e4, 5'd25, 27'h0000009f, 5'd8, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000c8, 5'd24, 27'h000000b7, 5'd19, 27'h00000312, 32'h00000400,
  1'd1,  5'd16, 27'h000002ec, 5'd24, 27'h00000163, 5'd30, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000007d, 5'd3, 27'h00000089, 5'd9, 27'h00000318, 32'h00000400,
  1'd1,  5'd28, 27'h00000108, 5'd3, 27'h0000009f, 5'd15, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000393, 5'd1, 27'h00000339, 5'd26, 27'h000001f5, 32'h00000400,
  1'd1,  5'd28, 27'h0000011b, 5'd14, 27'h0000031e, 5'd5, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000016b, 5'd10, 27'h000002be, 5'd20, 27'h0000021d, 32'h00000400,
  1'd1,  5'd26, 27'h00000379, 5'd15, 27'h00000135, 5'd26, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003df, 5'd22, 27'h000000f1, 5'd7, 27'h00000035, 32'h00000400,
  1'd1,  5'd30, 27'h000003c6, 5'd23, 27'h000001e5, 5'd16, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000037a, 5'd24, 27'h00000133, 5'd28, 27'h000001bb, 32'h00000400,
  1'd1,  5'd6, 27'h00000315, 5'd10, 27'h00000069, 5'd3, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a5, 5'd9, 27'h000001d6, 5'd11, 27'h0000004d, 32'h00000400,
  1'd1,  5'd9, 27'h00000305, 5'd9, 27'h0000020e, 5'd22, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000301, 5'd18, 27'h0000012c, 5'd2, 27'h0000006f, 32'h00000400,
  1'd1,  5'd7, 27'h0000006c, 5'd18, 27'h0000018e, 5'd10, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000047, 5'd20, 27'h000001f0, 5'd25, 27'h0000000d, 32'h00000400,
  1'd1,  5'd9, 27'h00000306, 5'd27, 27'h000000e1, 5'd1, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f5, 5'd27, 27'h000000b3, 5'd12, 27'h00000259, 32'h00000400,
  1'd1,  5'd6, 27'h00000336, 5'd30, 27'h00000239, 5'd20, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000068, 5'd6, 27'h00000049, 5'd0, 27'h00000062, 32'h00000400,
  1'd1,  5'd17, 27'h0000020e, 5'd9, 27'h000002a9, 5'd14, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b2, 5'd7, 27'h000000b8, 5'd24, 27'h00000202, 32'h00000400,
  1'd1,  5'd20, 27'h0000020f, 5'd16, 27'h000002d8, 5'd1, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000095, 5'd19, 27'h000002b3, 5'd13, 27'h00000376, 32'h00000400,
  1'd1,  5'd17, 27'h000001af, 5'd17, 27'h000002c6, 5'd23, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000339, 5'd30, 27'h000003de, 5'd4, 27'h0000026b, 32'h00000400,
  1'd1,  5'd16, 27'h00000200, 5'd28, 27'h0000001f, 5'd11, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ef, 5'd26, 27'h0000004c, 5'd24, 27'h000001a8, 32'h00000400,
  1'd1,  5'd26, 27'h0000005d, 5'd7, 27'h00000178, 5'd4, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c8, 5'd10, 27'h00000034, 5'd11, 27'h0000004f, 32'h00000400,
  1'd1,  5'd28, 27'h000001e8, 5'd6, 27'h00000398, 5'd24, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001fc, 5'd17, 27'h00000111, 5'd4, 27'h0000036e, 32'h00000400,
  1'd1,  5'd30, 27'h00000078, 5'd17, 27'h000003b3, 5'd10, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003f0, 5'd19, 27'h00000100, 5'd23, 27'h000003d2, 32'h00000400,
  1'd1,  5'd28, 27'h00000188, 5'd30, 27'h000003ff, 5'd0, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000033e, 5'd27, 27'h00000117, 5'd10, 27'h000002f0, 32'h00000400,
  1'd1,  5'd29, 27'h0000015a, 5'd27, 27'h000001a6, 5'd23, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000247, 5'd5, 27'h0000011e, 5'd10, 27'h00000054, 32'h00000400,
  1'd1,  5'd7, 27'h0000037a, 5'd5, 27'h000003e6, 5'd20, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000002e, 5'd6, 27'h00000032, 5'd27, 27'h000000b7, 32'h00000400,
  1'd1,  5'd8, 27'h00000369, 5'd17, 27'h00000302, 5'd6, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000018d, 5'd19, 27'h000001d1, 5'd18, 27'h00000043, 32'h00000400,
  1'd1,  5'd9, 27'h00000356, 5'd15, 27'h0000025d, 5'd30, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a8, 5'd27, 27'h000003f3, 5'd9, 27'h00000371, 32'h00000400,
  1'd1,  5'd7, 27'h000001f3, 5'd28, 27'h0000039d, 5'd17, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000181, 5'd30, 27'h000001f0, 5'd30, 27'h000000b4, 32'h00000400,
  1'd1,  5'd17, 27'h00000002, 5'd7, 27'h000003a1, 5'd6, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000308, 5'd5, 27'h000000ee, 5'd20, 27'h000001b1, 32'h00000400,
  1'd1,  5'd19, 27'h00000289, 5'd9, 27'h000003b8, 5'd27, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000019f, 5'd17, 27'h000003ee, 5'd5, 27'h0000035c, 32'h00000400,
  1'd1,  5'd16, 27'h0000001a, 5'd17, 27'h00000254, 5'd19, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000024e, 5'd19, 27'h0000002f, 5'd29, 27'h00000108, 32'h00000400,
  1'd1,  5'd19, 27'h00000202, 5'd29, 27'h00000286, 5'd8, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ad, 5'd28, 27'h000000f5, 5'd18, 27'h0000033b, 32'h00000400,
  1'd1,  5'd20, 27'h0000011d, 5'd28, 27'h0000020f, 5'd26, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000dd, 5'd9, 27'h0000016d, 5'd10, 27'h0000004d, 32'h00000400,
  1'd1,  5'd26, 27'h000000f9, 5'd8, 27'h0000031d, 5'd17, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000175, 5'd9, 27'h000001dc, 5'd26, 27'h0000033b, 32'h00000400,
  1'd1,  5'd30, 27'h0000007a, 5'd18, 27'h00000388, 5'd9, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003c3, 5'd15, 27'h00000397, 5'd18, 27'h000002d8, 32'h00000400,
  1'd1,  5'd29, 27'h0000030b, 5'd15, 27'h000003b8, 5'd28, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002b1, 5'd29, 27'h00000102, 5'd7, 27'h0000036a, 32'h00000400,
  1'd1,  5'd26, 27'h000000e1, 5'd27, 27'h00000035, 5'd17, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000348, 5'd29, 27'h00000252, 5'd26, 27'h000002e6, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000211, 5'd2, 27'h000000fa, 5'd4, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000008f, 5'd2, 27'h0000028c, 5'd12, 27'h000001a1, 32'h00000400,
  1'd1,  5'd4, 27'h000002e7, 5'd1, 27'h000001c9, 5'd21, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000129, 5'd14, 27'h0000024d, 5'd0, 27'h000000e4, 32'h00000400,
  1'd1,  5'd1, 27'h00000269, 5'd12, 27'h000003bc, 5'd11, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000235, 5'd12, 27'h000003e0, 5'd20, 27'h0000030a, 32'h00000400,
  1'd1,  5'd0, 27'h00000139, 5'd25, 27'h00000300, 5'd5, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000031a, 5'd24, 27'h0000026a, 5'd14, 27'h000002c6, 32'h00000400,
  1'd1,  5'd1, 27'h0000015a, 5'd25, 27'h0000009c, 5'd20, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000156, 5'd2, 27'h000001ae, 5'd2, 27'h0000022b, 32'h00000400,
  1'd1,  5'd10, 27'h000003d0, 5'd4, 27'h00000023, 5'd14, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000b2, 5'd0, 27'h00000093, 5'd20, 27'h00000343, 32'h00000400,
  1'd1,  5'd13, 27'h00000144, 5'd14, 27'h000001ce, 5'd2, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000007a, 5'd12, 27'h0000023a, 5'd11, 27'h0000028f, 32'h00000400,
  1'd1,  5'd14, 27'h0000008b, 5'd12, 27'h0000011b, 5'd25, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f3, 5'd23, 27'h00000307, 5'd0, 27'h00000047, 32'h00000400,
  1'd1,  5'd15, 27'h00000086, 5'd24, 27'h000000fd, 5'd14, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008d, 5'd21, 27'h000003af, 5'd25, 27'h000000ab, 32'h00000400,
  1'd1,  5'd22, 27'h0000035c, 5'd0, 27'h00000049, 5'd1, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000331, 5'd1, 27'h00000164, 5'd14, 27'h00000349, 32'h00000400,
  1'd1,  5'd25, 27'h00000058, 5'd4, 27'h000001b7, 5'd21, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000031f, 5'd13, 27'h00000175, 5'd2, 27'h0000012e, 32'h00000400,
  1'd1,  5'd22, 27'h000001ba, 5'd12, 27'h00000137, 5'd12, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000034c, 5'd14, 27'h00000008, 5'd23, 27'h0000000d, 32'h00000400,
  1'd1,  5'd24, 27'h0000017c, 5'd24, 27'h000000b8, 5'd1, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000309, 5'd22, 27'h000003e5, 5'd15, 27'h0000009a, 32'h00000400,
  1'd1,  5'd21, 27'h00000327, 5'd24, 27'h000001b0, 5'd21, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000003a, 5'd2, 27'h0000033e, 5'd10, 27'h00000035, 32'h00000400,
  1'd1,  5'd4, 27'h00000078, 5'd0, 27'h0000031e, 5'd18, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e9, 5'd0, 27'h0000032f, 5'd28, 27'h00000263, 32'h00000400,
  1'd1,  5'd4, 27'h00000250, 5'd12, 27'h00000317, 5'd7, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000130, 5'd15, 27'h000000b9, 5'd17, 27'h000000d9, 32'h00000400,
  1'd1,  5'd2, 27'h000001ea, 5'd13, 27'h000002fc, 5'd29, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000031a, 5'd21, 27'h00000384, 5'd5, 27'h000003a9, 32'h00000400,
  1'd1,  5'd0, 27'h00000386, 5'd24, 27'h00000124, 5'd16, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000043, 5'd20, 27'h0000039c, 5'd30, 27'h0000017e, 32'h00000400,
  1'd1,  5'd12, 27'h000001fe, 5'd0, 27'h00000237, 5'd10, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003c4, 5'd0, 27'h000000f1, 5'd18, 27'h000002fb, 32'h00000400,
  1'd1,  5'd13, 27'h00000163, 5'd4, 27'h00000376, 5'd28, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d3, 5'd11, 27'h00000080, 5'd9, 27'h000001ac, 32'h00000400,
  1'd1,  5'd11, 27'h00000378, 5'd13, 27'h000001cf, 5'd16, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000fd, 5'd10, 27'h00000156, 5'd27, 27'h000001b2, 32'h00000400,
  1'd1,  5'd14, 27'h000000d5, 5'd21, 27'h000001ac, 5'd10, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029c, 5'd21, 27'h000003cb, 5'd20, 27'h000000d6, 32'h00000400,
  1'd1,  5'd13, 27'h0000027e, 5'd24, 27'h00000110, 5'd30, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000014, 5'd4, 27'h000003f1, 5'd10, 27'h00000023, 32'h00000400,
  1'd1,  5'd23, 27'h000000da, 5'd1, 27'h00000298, 5'd17, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000343, 5'd2, 27'h000000ae, 5'd27, 27'h0000007e, 32'h00000400,
  1'd1,  5'd21, 27'h00000359, 5'd13, 27'h0000026f, 5'd7, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000009a, 5'd11, 27'h00000232, 5'd17, 27'h00000178, 32'h00000400,
  1'd1,  5'd25, 27'h00000049, 5'd10, 27'h00000263, 5'd27, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000037e, 5'd25, 27'h00000136, 5'd9, 27'h000000a7, 32'h00000400,
  1'd1,  5'd25, 27'h0000018b, 5'd22, 27'h000003ae, 5'd19, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000007c, 5'd21, 27'h0000023e, 5'd27, 27'h00000371, 32'h00000400,
  1'd1,  5'd0, 27'h000003c0, 5'd6, 27'h000000b6, 5'd2, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000038b, 5'd5, 27'h000001d9, 5'd11, 27'h000000cb, 32'h00000400,
  1'd1,  5'd2, 27'h000002aa, 5'd9, 27'h0000000b, 5'd22, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000233, 5'd15, 27'h0000039e, 5'd3, 27'h00000189, 32'h00000400,
  1'd1,  5'd3, 27'h000001bd, 5'd16, 27'h000001d4, 5'd12, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003bb, 5'd20, 27'h000001f8, 5'd23, 27'h000002a8, 32'h00000400,
  1'd1,  5'd2, 27'h0000011f, 5'd30, 27'h000002b5, 5'd4, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e2, 5'd30, 27'h00000204, 5'd11, 27'h000000d6, 32'h00000400,
  1'd1,  5'd3, 27'h00000373, 5'd30, 27'h000002d2, 5'd22, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000118, 5'd6, 27'h00000290, 5'd2, 27'h00000368, 32'h00000400,
  1'd1,  5'd13, 27'h000002db, 5'd7, 27'h00000142, 5'd12, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000119, 5'd7, 27'h000003a6, 5'd24, 27'h000001a3, 32'h00000400,
  1'd1,  5'd13, 27'h00000098, 5'd18, 27'h0000032f, 5'd1, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000282, 5'd19, 27'h00000317, 5'd11, 27'h000002fd, 32'h00000400,
  1'd1,  5'd13, 27'h00000248, 5'd17, 27'h00000146, 5'd24, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000061, 5'd26, 27'h0000015d, 5'd5, 27'h00000087, 32'h00000400,
  1'd1,  5'd11, 27'h0000019d, 5'd27, 27'h0000036b, 5'd15, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000035e, 5'd27, 27'h00000106, 5'd20, 27'h00000369, 32'h00000400,
  1'd1,  5'd21, 27'h000002c4, 5'd8, 27'h00000379, 5'd1, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000042, 5'd8, 27'h00000177, 5'd11, 27'h000000a9, 32'h00000400,
  1'd1,  5'd23, 27'h000003cb, 5'd10, 27'h000000b7, 5'd22, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002bd, 5'd16, 27'h00000057, 5'd3, 27'h000003ae, 32'h00000400,
  1'd1,  5'd21, 27'h00000399, 5'd15, 27'h00000390, 5'd14, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000249, 5'd18, 27'h000003de, 5'd22, 27'h000001eb, 32'h00000400,
  1'd1,  5'd25, 27'h000001bf, 5'd26, 27'h000001f9, 5'd2, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000030e, 5'd26, 27'h00000350, 5'd14, 27'h000000a1, 32'h00000400,
  1'd1,  5'd25, 27'h0000018e, 5'd26, 27'h000002cd, 5'd23, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000023e, 5'd9, 27'h0000011c, 5'd6, 27'h000000e0, 32'h00000400,
  1'd1,  5'd2, 27'h00000113, 5'd7, 27'h000000d5, 5'd19, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e2, 5'd9, 27'h0000039f, 5'd30, 27'h00000071, 32'h00000400,
  1'd1,  5'd4, 27'h00000002, 5'd16, 27'h00000071, 5'd8, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000261, 5'd16, 27'h0000019e, 5'd20, 27'h0000012e, 32'h00000400,
  1'd1,  5'd0, 27'h000000dc, 5'd20, 27'h000001f0, 5'd30, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000023a, 5'd27, 27'h000000bb, 5'd7, 27'h000003de, 32'h00000400,
  1'd1,  5'd1, 27'h00000152, 5'd28, 27'h0000013d, 5'd19, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000031e, 5'd26, 27'h0000028e, 5'd30, 27'h00000298, 32'h00000400,
  1'd1,  5'd13, 27'h000000d7, 5'd8, 27'h00000257, 5'd8, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ff, 5'd5, 27'h000001f7, 5'd20, 27'h00000114, 32'h00000400,
  1'd1,  5'd10, 27'h00000174, 5'd8, 27'h00000208, 5'd30, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000019e, 5'd17, 27'h0000032c, 5'd10, 27'h00000097, 32'h00000400,
  1'd1,  5'd10, 27'h000001e0, 5'd19, 27'h0000008b, 5'd19, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001cb, 5'd19, 27'h0000010a, 5'd26, 27'h00000157, 32'h00000400,
  1'd1,  5'd12, 27'h00000089, 5'd28, 27'h00000102, 5'd10, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000217, 5'd27, 27'h00000351, 5'd18, 27'h00000061, 32'h00000400,
  1'd1,  5'd12, 27'h000002ae, 5'd25, 27'h0000037f, 5'd27, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000021c, 5'd9, 27'h00000293, 5'd6, 27'h000001cb, 32'h00000400,
  1'd1,  5'd21, 27'h0000029a, 5'd6, 27'h00000290, 5'd19, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000bf, 5'd7, 27'h000001c7, 5'd29, 27'h000002ff, 32'h00000400,
  1'd1,  5'd25, 27'h000002a3, 5'd17, 27'h0000016b, 5'd9, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001fd, 5'd16, 27'h000002fc, 5'd16, 27'h0000007c, 32'h00000400,
  1'd1,  5'd22, 27'h00000118, 5'd20, 27'h000000d0, 5'd27, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000e9, 5'd30, 27'h0000027b, 5'd9, 27'h000003ae, 32'h00000400,
  1'd1,  5'd24, 27'h0000035e, 5'd28, 27'h000000d3, 5'd17, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000ce, 5'd30, 27'h000003d7, 5'd27, 27'h0000025e, 32'h00000400,
  1'd1,  5'd7, 27'h00000311, 5'd3, 27'h0000013c, 5'd10, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ff, 5'd0, 27'h000003b7, 5'd17, 27'h00000064, 32'h00000400,
  1'd1,  5'd9, 27'h00000147, 5'd4, 27'h000000b7, 5'd27, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000027d, 5'd12, 27'h000003bf, 5'd1, 27'h0000001d, 32'h00000400,
  1'd1,  5'd5, 27'h0000027e, 5'd12, 27'h00000251, 5'd13, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000163, 5'd10, 27'h0000034e, 5'd21, 27'h000003cf, 32'h00000400,
  1'd1,  5'd8, 27'h00000397, 5'd24, 27'h000003d3, 5'd2, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000038a, 5'd23, 27'h00000148, 5'd14, 27'h0000037c, 32'h00000400,
  1'd1,  5'd7, 27'h0000009d, 5'd24, 27'h0000024a, 5'd24, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000021e, 5'd3, 27'h00000078, 5'd7, 27'h000003ad, 32'h00000400,
  1'd1,  5'd19, 27'h0000013b, 5'd4, 27'h00000013, 5'd18, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000036c, 5'd3, 27'h0000038e, 5'd29, 27'h00000040, 32'h00000400,
  1'd1,  5'd16, 27'h000001e3, 5'd12, 27'h000000ee, 5'd2, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000383, 5'd11, 27'h00000191, 5'd14, 27'h000000ca, 32'h00000400,
  1'd1,  5'd15, 27'h0000034b, 5'd10, 27'h00000311, 5'd21, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000010b, 5'd22, 27'h000003d5, 5'd3, 27'h000003ee, 32'h00000400,
  1'd1,  5'd15, 27'h00000358, 5'd22, 27'h000001b8, 5'd15, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000338, 5'd21, 27'h000000c2, 5'd23, 27'h00000245, 32'h00000400,
  1'd1,  5'd27, 27'h0000031d, 5'd3, 27'h00000282, 5'd3, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c8, 5'd3, 27'h00000355, 5'd13, 27'h0000028a, 32'h00000400,
  1'd1,  5'd29, 27'h0000009a, 5'd0, 27'h0000004f, 5'd23, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000314, 5'd11, 27'h000000ba, 5'd0, 27'h0000034a, 32'h00000400,
  1'd1,  5'd27, 27'h0000008e, 5'd14, 27'h00000319, 5'd14, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000016d, 5'd14, 27'h000001d8, 5'd25, 27'h000001f2, 32'h00000400,
  1'd1,  5'd26, 27'h0000012c, 5'd20, 27'h000002e9, 5'd5, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000c4, 5'd22, 27'h0000011f, 5'd12, 27'h000003b9, 32'h00000400,
  1'd1,  5'd29, 27'h000000bc, 5'd25, 27'h000002ce, 5'd23, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b8, 5'd1, 27'h000002b0, 5'd1, 27'h00000156, 32'h00000400,
  1'd1,  5'd7, 27'h000003c9, 5'd1, 27'h00000051, 5'd11, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000024c, 5'd3, 27'h000002f3, 5'd21, 27'h00000314, 32'h00000400,
  1'd1,  5'd9, 27'h00000049, 5'd13, 27'h00000109, 5'd6, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000280, 5'd10, 27'h000001b4, 5'd18, 27'h0000012b, 32'h00000400,
  1'd1,  5'd9, 27'h00000341, 5'd13, 27'h00000187, 5'd29, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003da, 5'd21, 27'h000002a8, 5'd8, 27'h00000097, 32'h00000400,
  1'd1,  5'd5, 27'h00000167, 5'd25, 27'h00000222, 5'd16, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ad, 5'd24, 27'h0000029d, 5'd27, 27'h0000008e, 32'h00000400,
  1'd1,  5'd16, 27'h0000026b, 5'd2, 27'h000003b2, 5'd1, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000184, 5'd4, 27'h00000021, 5'd14, 27'h0000039a, 32'h00000400,
  1'd1,  5'd17, 27'h00000173, 5'd1, 27'h000003dd, 5'd22, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000298, 5'd13, 27'h000001a8, 5'd10, 27'h0000011f, 32'h00000400,
  1'd1,  5'd16, 27'h000002b6, 5'd14, 27'h00000078, 5'd19, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000128, 5'd13, 27'h00000201, 5'd27, 27'h00000139, 32'h00000400,
  1'd1,  5'd17, 27'h000001c4, 5'd22, 27'h000000e4, 5'd5, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000224, 5'd23, 27'h0000010b, 5'd18, 27'h0000039e, 32'h00000400,
  1'd1,  5'd18, 27'h0000030b, 5'd21, 27'h000003ab, 5'd30, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000114, 5'd0, 27'h00000378, 5'd10, 27'h000000d4, 32'h00000400,
  1'd1,  5'd29, 27'h00000087, 5'd5, 27'h00000085, 5'd20, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b0, 5'd1, 27'h0000005e, 5'd27, 27'h00000014, 32'h00000400,
  1'd1,  5'd29, 27'h00000232, 5'd10, 27'h00000284, 5'd7, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000af, 5'd12, 27'h00000150, 5'd18, 27'h00000156, 32'h00000400,
  1'd1,  5'd27, 27'h0000010c, 5'd14, 27'h00000069, 5'd30, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000102, 5'd23, 27'h000000ca, 5'd6, 27'h000003fb, 32'h00000400,
  1'd1,  5'd26, 27'h000000de, 5'd24, 27'h00000192, 5'd18, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000035f, 5'd24, 27'h000002f4, 5'd27, 27'h00000013, 32'h00000400,
  1'd1,  5'd8, 27'h00000269, 5'd7, 27'h00000215, 5'd3, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000172, 5'd7, 27'h00000154, 5'd14, 27'h0000025c, 32'h00000400,
  1'd1,  5'd6, 27'h00000146, 5'd6, 27'h000003b4, 5'd25, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001b4, 5'd17, 27'h00000035, 5'd1, 27'h0000017a, 32'h00000400,
  1'd1,  5'd9, 27'h00000120, 5'd19, 27'h00000141, 5'd13, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000083, 5'd19, 27'h000002fd, 5'd23, 27'h00000371, 32'h00000400,
  1'd1,  5'd7, 27'h00000001, 5'd28, 27'h000002c2, 5'd1, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000368, 5'd29, 27'h000002fa, 5'd13, 27'h000002a6, 32'h00000400,
  1'd1,  5'd9, 27'h0000010b, 5'd26, 27'h000002cb, 5'd22, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000007a, 5'd10, 27'h00000061, 5'd0, 27'h000000b2, 32'h00000400,
  1'd1,  5'd16, 27'h0000021e, 5'd8, 27'h000002bb, 5'd12, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d7, 5'd5, 27'h00000372, 5'd21, 27'h000002e6, 32'h00000400,
  1'd1,  5'd16, 27'h00000178, 5'd17, 27'h00000367, 5'd5, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f9, 5'd19, 27'h000000f1, 5'd10, 27'h000003ee, 32'h00000400,
  1'd1,  5'd17, 27'h00000337, 5'd16, 27'h000000f9, 5'd22, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000253, 5'd28, 27'h000003e1, 5'd4, 27'h00000044, 32'h00000400,
  1'd1,  5'd18, 27'h000003db, 5'd26, 27'h00000191, 5'd13, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000300, 5'd30, 27'h00000237, 5'd21, 27'h00000370, 32'h00000400,
  1'd1,  5'd25, 27'h00000357, 5'd6, 27'h00000300, 5'd3, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001f8, 5'd10, 27'h000000c7, 5'd15, 27'h000001ab, 32'h00000400,
  1'd1,  5'd29, 27'h000001c7, 5'd7, 27'h00000252, 5'd23, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000010, 5'd16, 27'h0000010f, 5'd4, 27'h0000034e, 32'h00000400,
  1'd1,  5'd30, 27'h0000035c, 5'd17, 27'h000001d3, 5'd15, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000383, 5'd19, 27'h00000309, 5'd25, 27'h000000a2, 32'h00000400,
  1'd1,  5'd28, 27'h000003eb, 5'd28, 27'h00000284, 5'd1, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000014b, 5'd26, 27'h000001cb, 5'd11, 27'h00000225, 32'h00000400,
  1'd1,  5'd28, 27'h0000034a, 5'd26, 27'h00000216, 5'd25, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000364, 5'd7, 27'h000001e7, 5'd9, 27'h00000333, 32'h00000400,
  1'd1,  5'd9, 27'h00000197, 5'd7, 27'h0000011d, 5'd15, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001fc, 5'd10, 27'h0000003f, 5'd30, 27'h00000181, 32'h00000400,
  1'd1,  5'd7, 27'h000003a4, 5'd17, 27'h000000e9, 5'd7, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031b, 5'd16, 27'h00000335, 5'd17, 27'h0000000c, 32'h00000400,
  1'd1,  5'd7, 27'h000000e8, 5'd16, 27'h000003c0, 5'd28, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001dc, 5'd27, 27'h000003f2, 5'd6, 27'h000001cd, 32'h00000400,
  1'd1,  5'd9, 27'h0000024d, 5'd26, 27'h000003e9, 5'd17, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000259, 5'd27, 27'h0000006d, 5'd30, 27'h0000002e, 32'h00000400,
  1'd1,  5'd15, 27'h000003e6, 5'd6, 27'h000001bb, 5'd6, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e0, 5'd8, 27'h0000012a, 5'd19, 27'h00000081, 32'h00000400,
  1'd1,  5'd18, 27'h0000010f, 5'd5, 27'h0000020e, 5'd29, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000bc, 5'd18, 27'h0000024e, 5'd7, 27'h00000131, 32'h00000400,
  1'd1,  5'd20, 27'h0000024b, 5'd15, 27'h00000270, 5'd15, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c5, 5'd15, 27'h000003cf, 5'd26, 27'h0000021c, 32'h00000400,
  1'd1,  5'd16, 27'h000000ca, 5'd30, 27'h00000040, 5'd7, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000fb, 5'd28, 27'h000001cb, 5'd18, 27'h0000032a, 32'h00000400,
  1'd1,  5'd17, 27'h000003ad, 5'd28, 27'h000003b8, 5'd26, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000190, 5'd8, 27'h00000106, 5'd5, 27'h000002d7, 32'h00000400,
  1'd1,  5'd27, 27'h0000033b, 5'd9, 27'h0000028e, 5'd19, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000030a, 5'd9, 27'h000003bb, 5'd28, 27'h000000bc, 32'h00000400,
  1'd1,  5'd29, 27'h0000002a, 5'd16, 27'h00000128, 5'd5, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f2, 5'd16, 27'h00000155, 5'd17, 27'h00000184, 32'h00000400,
  1'd1,  5'd28, 27'h000002be, 5'd17, 27'h000000a6, 5'd29, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f4, 5'd30, 27'h0000039b, 5'd8, 27'h00000042, 32'h00000400,
  1'd1,  5'd27, 27'h000001c9, 5'd27, 27'h0000000c, 5'd20, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000373, 5'd27, 27'h00000080, 5'd30, 27'h000003d9, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h0000026c, 5'd2, 27'h000002cb, 5'd3, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000230, 5'd2, 27'h000001e9, 5'd11, 27'h000001f3, 32'h00000400,
  1'd1,  5'd2, 27'h000000ac, 5'd2, 27'h00000103, 5'd22, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000062, 5'd13, 27'h0000026d, 5'd1, 27'h00000336, 32'h00000400,
  1'd1,  5'd4, 27'h0000031a, 5'd12, 27'h00000017, 5'd15, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000241, 5'd12, 27'h00000035, 5'd23, 27'h00000184, 32'h00000400,
  1'd1,  5'd2, 27'h00000020, 5'd21, 27'h000002e9, 5'd0, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000007, 5'd24, 27'h000003b5, 5'd13, 27'h00000168, 32'h00000400,
  1'd1,  5'd1, 27'h0000039b, 5'd25, 27'h00000137, 5'd23, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001da, 5'd2, 27'h00000336, 5'd3, 27'h000001b1, 32'h00000400,
  1'd1,  5'd13, 27'h0000010e, 5'd3, 27'h00000341, 5'd14, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d1, 5'd0, 27'h00000312, 5'd25, 27'h000001cd, 32'h00000400,
  1'd1,  5'd10, 27'h00000302, 5'd15, 27'h0000013f, 5'd3, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000002, 5'd10, 27'h00000191, 5'd14, 27'h00000039, 32'h00000400,
  1'd1,  5'd15, 27'h00000004, 5'd15, 27'h00000108, 5'd21, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000024b, 5'd23, 27'h000002ad, 5'd2, 27'h0000034e, 32'h00000400,
  1'd1,  5'd11, 27'h000003bf, 5'd21, 27'h00000338, 5'd11, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000307, 5'd22, 27'h0000032e, 5'd23, 27'h00000094, 32'h00000400,
  1'd1,  5'd23, 27'h00000258, 5'd0, 27'h000003ce, 5'd1, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000030f, 5'd2, 27'h00000220, 5'd12, 27'h000000f0, 32'h00000400,
  1'd1,  5'd23, 27'h00000198, 5'd0, 27'h0000018d, 5'd20, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000004, 5'd11, 27'h000000c6, 5'd0, 27'h000000bc, 32'h00000400,
  1'd1,  5'd23, 27'h000000ec, 5'd13, 27'h000003b1, 5'd14, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000002f, 5'd13, 27'h00000085, 5'd24, 27'h0000004e, 32'h00000400,
  1'd1,  5'd20, 27'h0000035a, 5'd21, 27'h00000007, 5'd2, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000002f, 5'd21, 27'h00000102, 5'd13, 27'h00000138, 32'h00000400,
  1'd1,  5'd22, 27'h000000cc, 5'd23, 27'h00000301, 5'd22, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002bd, 5'd1, 27'h000003ef, 5'd7, 27'h000000db, 32'h00000400,
  1'd1,  5'd5, 27'h0000006a, 5'd4, 27'h000002fe, 5'd15, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e1, 5'd3, 27'h000001b7, 5'd26, 27'h00000016, 32'h00000400,
  1'd1,  5'd3, 27'h00000303, 5'd14, 27'h00000176, 5'd10, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000012d, 5'd12, 27'h0000029a, 5'd16, 27'h00000309, 32'h00000400,
  1'd1,  5'd0, 27'h00000074, 5'd12, 27'h00000121, 5'd28, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b6, 5'd23, 27'h000000c1, 5'd5, 27'h0000035c, 32'h00000400,
  1'd1,  5'd2, 27'h00000019, 5'd24, 27'h000001f7, 5'd19, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017f, 5'd22, 27'h00000168, 5'd28, 27'h000002c9, 32'h00000400,
  1'd1,  5'd10, 27'h0000035d, 5'd3, 27'h0000007d, 5'd9, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ae, 5'd0, 27'h0000033b, 5'd20, 27'h00000275, 32'h00000400,
  1'd1,  5'd12, 27'h00000368, 5'd0, 27'h00000045, 5'd28, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000083, 5'd12, 27'h00000293, 5'd5, 27'h00000277, 32'h00000400,
  1'd1,  5'd14, 27'h000002e4, 5'd11, 27'h00000063, 5'd19, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000027a, 5'd12, 27'h00000086, 5'd28, 27'h0000039d, 32'h00000400,
  1'd1,  5'd11, 27'h000003fc, 5'd22, 27'h00000034, 5'd7, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000239, 5'd22, 27'h00000347, 5'd20, 27'h00000212, 32'h00000400,
  1'd1,  5'd14, 27'h00000108, 5'd22, 27'h0000029f, 5'd29, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001af, 5'd0, 27'h00000156, 5'd8, 27'h000002b6, 32'h00000400,
  1'd1,  5'd21, 27'h0000035b, 5'd2, 27'h000003f8, 5'd19, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000023f, 5'd0, 27'h00000077, 5'd29, 27'h000000df, 32'h00000400,
  1'd1,  5'd23, 27'h00000260, 5'd14, 27'h000000e6, 5'd5, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000242, 5'd14, 27'h0000027d, 5'd19, 27'h0000031f, 32'h00000400,
  1'd1,  5'd24, 27'h00000385, 5'd11, 27'h000002e3, 5'd28, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a5, 5'd21, 27'h00000389, 5'd8, 27'h0000016b, 32'h00000400,
  1'd1,  5'd25, 27'h00000201, 5'd25, 27'h000001d5, 5'd16, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000093, 5'd21, 27'h000002f9, 5'd28, 27'h00000272, 32'h00000400,
  1'd1,  5'd1, 27'h0000021b, 5'd6, 27'h000003c0, 5'd0, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000010f, 5'd7, 27'h000002ed, 5'd13, 27'h000000ad, 32'h00000400,
  1'd1,  5'd4, 27'h00000156, 5'd8, 27'h000003d8, 5'd20, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000320, 5'd17, 27'h00000162, 5'd4, 27'h000001ab, 32'h00000400,
  1'd1,  5'd2, 27'h00000193, 5'd19, 27'h00000264, 5'd11, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027a, 5'd17, 27'h00000330, 5'd25, 27'h00000259, 32'h00000400,
  1'd1,  5'd0, 27'h000000d7, 5'd29, 27'h000002a6, 5'd3, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000d2, 5'd28, 27'h000002cb, 5'd10, 27'h00000216, 32'h00000400,
  1'd1,  5'd1, 27'h000000e9, 5'd29, 27'h0000028e, 5'd20, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f9, 5'd9, 27'h0000010e, 5'd2, 27'h00000119, 32'h00000400,
  1'd1,  5'd12, 27'h000000b9, 5'd9, 27'h0000031e, 5'd12, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000373, 5'd10, 27'h0000014c, 5'd23, 27'h000003fb, 32'h00000400,
  1'd1,  5'd13, 27'h0000029f, 5'd19, 27'h000001b1, 5'd4, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000014f, 5'd19, 27'h0000017f, 5'd12, 27'h00000227, 32'h00000400,
  1'd1,  5'd13, 27'h00000183, 5'd17, 27'h000003a0, 5'd22, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000018b, 5'd27, 27'h00000309, 5'd0, 27'h0000034d, 32'h00000400,
  1'd1,  5'd14, 27'h00000119, 5'd29, 27'h00000333, 5'd13, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000140, 5'd29, 27'h000000f0, 5'd23, 27'h000002b4, 32'h00000400,
  1'd1,  5'd20, 27'h000003cf, 5'd10, 27'h00000073, 5'd0, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000004e, 5'd8, 27'h0000034c, 5'd11, 27'h000002fa, 32'h00000400,
  1'd1,  5'd24, 27'h000000b6, 5'd9, 27'h0000019d, 5'd23, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000374, 5'd19, 27'h000000a0, 5'd1, 27'h00000116, 32'h00000400,
  1'd1,  5'd24, 27'h0000029e, 5'd15, 27'h0000020c, 5'd10, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000010b, 5'd17, 27'h00000244, 5'd22, 27'h0000021f, 32'h00000400,
  1'd1,  5'd25, 27'h00000118, 5'd29, 27'h0000016f, 5'd2, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000008, 5'd27, 27'h00000290, 5'd12, 27'h0000029f, 32'h00000400,
  1'd1,  5'd24, 27'h000001d7, 5'd27, 27'h00000032, 5'd24, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000018, 5'd9, 27'h000001d0, 5'd6, 27'h00000396, 32'h00000400,
  1'd1,  5'd0, 27'h0000037b, 5'd8, 27'h0000030f, 5'd20, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000014, 5'd9, 27'h00000000, 5'd29, 27'h00000224, 32'h00000400,
  1'd1,  5'd3, 27'h00000175, 5'd19, 27'h000003be, 5'd5, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000038a, 5'd19, 27'h000000cc, 5'd16, 27'h00000025, 32'h00000400,
  1'd1,  5'd3, 27'h00000085, 5'd16, 27'h0000006e, 5'd29, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003a3, 5'd26, 27'h0000015d, 5'd8, 27'h00000037, 32'h00000400,
  1'd1,  5'd4, 27'h0000009e, 5'd29, 27'h000003a4, 5'd16, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000001, 5'd30, 27'h0000012e, 5'd30, 27'h00000191, 32'h00000400,
  1'd1,  5'd14, 27'h000002ad, 5'd6, 27'h00000201, 5'd9, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003c1, 5'd6, 27'h00000304, 5'd16, 27'h0000015b, 32'h00000400,
  1'd1,  5'd11, 27'h0000022d, 5'd6, 27'h0000020a, 5'd30, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ad, 5'd18, 27'h00000182, 5'd9, 27'h000001f9, 32'h00000400,
  1'd1,  5'd13, 27'h00000123, 5'd19, 27'h000002cd, 5'd17, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ea, 5'd19, 27'h0000023c, 5'd30, 27'h000003ad, 32'h00000400,
  1'd1,  5'd10, 27'h000002c2, 5'd29, 27'h000000a8, 5'd5, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017b, 5'd28, 27'h000002f4, 5'd17, 27'h00000238, 32'h00000400,
  1'd1,  5'd11, 27'h00000321, 5'd27, 27'h000003f2, 5'd27, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000d3, 5'd7, 27'h000000c3, 5'd7, 27'h00000124, 32'h00000400,
  1'd1,  5'd22, 27'h00000156, 5'd8, 27'h00000253, 5'd20, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f3, 5'd9, 27'h000002bb, 5'd27, 27'h00000220, 32'h00000400,
  1'd1,  5'd25, 27'h000002f1, 5'd19, 27'h000001d9, 5'd8, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000219, 5'd16, 27'h00000071, 5'd16, 27'h00000205, 32'h00000400,
  1'd1,  5'd22, 27'h000003a5, 5'd17, 27'h00000397, 5'd30, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000032, 5'd30, 27'h0000007c, 5'd6, 27'h000003c4, 32'h00000400,
  1'd1,  5'd23, 27'h000000a8, 5'd26, 27'h00000261, 5'd19, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000228, 5'd27, 27'h00000068, 5'd28, 27'h000003c4, 32'h00000400,
  1'd1,  5'd7, 27'h00000345, 5'd0, 27'h000000c2, 5'd8, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e4, 5'd4, 27'h00000305, 5'd18, 27'h000003fe, 32'h00000400,
  1'd1,  5'd9, 27'h000002c2, 5'd3, 27'h00000278, 5'd30, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000135, 5'd11, 27'h0000004b, 5'd4, 27'h00000239, 32'h00000400,
  1'd1,  5'd6, 27'h000002fc, 5'd12, 27'h00000318, 5'd15, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000329, 5'd14, 27'h0000021d, 5'd25, 27'h0000015d, 32'h00000400,
  1'd1,  5'd6, 27'h000003db, 5'd25, 27'h00000076, 5'd4, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ff, 5'd23, 27'h00000099, 5'd10, 27'h00000343, 32'h00000400,
  1'd1,  5'd5, 27'h0000032f, 5'd24, 27'h00000138, 5'd22, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000dd, 5'd3, 27'h000001d7, 5'd7, 27'h0000009c, 32'h00000400,
  1'd1,  5'd20, 27'h00000141, 5'd2, 27'h0000019e, 5'd19, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000017, 5'd0, 27'h000000a2, 5'd26, 27'h000000a9, 32'h00000400,
  1'd1,  5'd18, 27'h000003b4, 5'd11, 27'h00000272, 5'd4, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000003a, 5'd12, 27'h00000046, 5'd14, 27'h000000c3, 32'h00000400,
  1'd1,  5'd15, 27'h0000032c, 5'd12, 27'h00000065, 5'd23, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000010c, 5'd21, 27'h0000022e, 5'd4, 27'h00000273, 32'h00000400,
  1'd1,  5'd15, 27'h00000320, 5'd23, 27'h0000031a, 5'd14, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002f5, 5'd23, 27'h000000d7, 5'd22, 27'h0000013c, 32'h00000400,
  1'd1,  5'd27, 27'h0000011b, 5'd3, 27'h000002a8, 5'd2, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000271, 5'd4, 27'h000001ca, 5'd13, 27'h00000133, 32'h00000400,
  1'd1,  5'd26, 27'h00000119, 5'd4, 27'h000000e0, 5'd21, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001d9, 5'd10, 27'h000002a7, 5'd2, 27'h00000037, 32'h00000400,
  1'd1,  5'd26, 27'h0000022d, 5'd10, 27'h00000273, 5'd10, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000001, 5'd13, 27'h00000353, 5'd22, 27'h000002d5, 32'h00000400,
  1'd1,  5'd26, 27'h0000017a, 5'd23, 27'h0000039b, 5'd4, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000206, 5'd21, 27'h00000147, 5'd14, 27'h00000339, 32'h00000400,
  1'd1,  5'd26, 27'h0000022d, 5'd21, 27'h00000017, 5'd25, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c3, 5'd1, 27'h00000384, 5'd2, 27'h000002ae, 32'h00000400,
  1'd1,  5'd5, 27'h00000379, 5'd1, 27'h0000011b, 5'd11, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000236, 5'd1, 27'h00000084, 5'd23, 27'h00000055, 32'h00000400,
  1'd1,  5'd6, 27'h0000013b, 5'd15, 27'h000000a4, 5'd9, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000014, 5'd11, 27'h00000315, 5'd20, 27'h000000b9, 32'h00000400,
  1'd1,  5'd9, 27'h0000028a, 5'd11, 27'h0000031c, 5'd30, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ba, 5'd24, 27'h00000310, 5'd8, 27'h0000027f, 32'h00000400,
  1'd1,  5'd7, 27'h00000191, 5'd25, 27'h00000301, 5'd18, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000278, 5'd21, 27'h0000002c, 5'd27, 27'h000001e3, 32'h00000400,
  1'd1,  5'd19, 27'h000000fe, 5'd2, 27'h0000038a, 5'd1, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000012a, 5'd0, 27'h000001b7, 5'd12, 27'h00000332, 32'h00000400,
  1'd1,  5'd15, 27'h00000359, 5'd0, 27'h00000375, 5'd23, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003b8, 5'd14, 27'h0000016f, 5'd6, 27'h000000a5, 32'h00000400,
  1'd1,  5'd16, 27'h000003fa, 5'd11, 27'h00000174, 5'd18, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000022a, 5'd14, 27'h000001d5, 5'd28, 27'h0000030d, 32'h00000400,
  1'd1,  5'd18, 27'h0000035f, 5'd23, 27'h0000029e, 5'd8, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000014e, 5'd22, 27'h00000038, 5'd17, 27'h000001c7, 32'h00000400,
  1'd1,  5'd19, 27'h00000056, 5'd23, 27'h000001a6, 5'd29, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023c, 5'd3, 27'h00000255, 5'd8, 27'h000002c3, 32'h00000400,
  1'd1,  5'd26, 27'h000003e3, 5'd2, 27'h0000011e, 5'd18, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000268, 5'd4, 27'h00000320, 5'd30, 27'h000003d3, 32'h00000400,
  1'd1,  5'd28, 27'h000000e0, 5'd12, 27'h000001c7, 5'd7, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007b, 5'd14, 27'h00000255, 5'd17, 27'h000002cd, 32'h00000400,
  1'd1,  5'd30, 27'h0000008c, 5'd13, 27'h00000059, 5'd28, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024b, 5'd25, 27'h000000db, 5'd5, 27'h00000399, 32'h00000400,
  1'd1,  5'd27, 27'h000000bc, 5'd20, 27'h00000361, 5'd18, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000133, 5'd25, 27'h000002c5, 5'd29, 27'h0000001b, 32'h00000400,
  1'd1,  5'd7, 27'h0000003e, 5'd7, 27'h00000307, 5'd2, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002e2, 5'd10, 27'h00000154, 5'd13, 27'h00000161, 32'h00000400,
  1'd1,  5'd9, 27'h000000f1, 5'd5, 27'h000002e8, 5'd22, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000018, 5'd19, 27'h00000346, 5'd3, 27'h000000db, 32'h00000400,
  1'd1,  5'd5, 27'h00000131, 5'd20, 27'h00000270, 5'd12, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000e7, 5'd19, 27'h0000007a, 5'd21, 27'h00000131, 32'h00000400,
  1'd1,  5'd8, 27'h00000214, 5'd29, 27'h00000049, 5'd0, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000dd, 5'd29, 27'h000000aa, 5'd13, 27'h0000018d, 32'h00000400,
  1'd1,  5'd9, 27'h00000193, 5'd27, 27'h000003e5, 5'd20, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003b2, 5'd8, 27'h0000009d, 5'd4, 27'h000003d5, 32'h00000400,
  1'd1,  5'd17, 27'h000002ce, 5'd5, 27'h0000039a, 5'd12, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000139, 5'd9, 27'h00000395, 5'd25, 27'h00000134, 32'h00000400,
  1'd1,  5'd19, 27'h000003a2, 5'd19, 27'h000001aa, 5'd2, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000223, 5'd20, 27'h00000059, 5'd12, 27'h00000085, 32'h00000400,
  1'd1,  5'd16, 27'h0000017f, 5'd16, 27'h0000003f, 5'd24, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001e8, 5'd30, 27'h0000020a, 5'd3, 27'h00000349, 32'h00000400,
  1'd1,  5'd15, 27'h000003fc, 5'd27, 27'h000000ef, 5'd14, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001bd, 5'd29, 27'h000003b5, 5'd25, 27'h00000258, 32'h00000400,
  1'd1,  5'd26, 27'h00000294, 5'd9, 27'h00000386, 5'd0, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000278, 5'd8, 27'h00000192, 5'd10, 27'h00000245, 32'h00000400,
  1'd1,  5'd27, 27'h0000012a, 5'd6, 27'h000002d8, 5'd23, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000396, 5'd16, 27'h000003fe, 5'd1, 27'h000000a8, 32'h00000400,
  1'd1,  5'd28, 27'h000001e6, 5'd19, 27'h00000328, 5'd12, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f5, 5'd20, 27'h00000172, 5'd22, 27'h00000344, 32'h00000400,
  1'd1,  5'd26, 27'h00000169, 5'd30, 27'h000003f9, 5'd3, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b8, 5'd27, 27'h000000e3, 5'd11, 27'h00000390, 32'h00000400,
  1'd1,  5'd27, 27'h00000046, 5'd28, 27'h00000037, 5'd21, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000364, 5'd6, 27'h000003c9, 5'd9, 27'h000003d3, 32'h00000400,
  1'd1,  5'd6, 27'h0000033b, 5'd9, 27'h00000056, 5'd20, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000003b, 5'd5, 27'h00000320, 5'd25, 27'h000003ce, 32'h00000400,
  1'd1,  5'd6, 27'h000001b6, 5'd17, 27'h000000dd, 5'd10, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003a7, 5'd19, 27'h000002bd, 5'd19, 27'h000001a2, 32'h00000400,
  1'd1,  5'd10, 27'h000000ea, 5'd19, 27'h00000147, 5'd26, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000002c, 5'd26, 27'h0000012f, 5'd5, 27'h00000137, 32'h00000400,
  1'd1,  5'd7, 27'h00000381, 5'd29, 27'h00000179, 5'd16, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000396, 5'd27, 27'h000000d3, 5'd29, 27'h0000036d, 32'h00000400,
  1'd1,  5'd15, 27'h0000038d, 5'd6, 27'h000001ca, 5'd10, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034f, 5'd5, 27'h00000208, 5'd18, 27'h0000037c, 32'h00000400,
  1'd1,  5'd18, 27'h000002ad, 5'd7, 27'h000000e6, 5'd29, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000223, 5'd17, 27'h00000305, 5'd5, 27'h00000343, 32'h00000400,
  1'd1,  5'd19, 27'h0000018f, 5'd17, 27'h00000135, 5'd16, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000036a, 5'd20, 27'h00000268, 5'd27, 27'h00000259, 32'h00000400,
  1'd1,  5'd18, 27'h00000093, 5'd27, 27'h0000009b, 5'd10, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000002c, 5'd26, 27'h0000028b, 5'd17, 27'h00000208, 32'h00000400,
  1'd1,  5'd19, 27'h000003ac, 5'd29, 27'h00000098, 5'd29, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000357, 5'd8, 27'h000002a0, 5'd5, 27'h000003d2, 32'h00000400,
  1'd1,  5'd30, 27'h00000150, 5'd6, 27'h0000009b, 5'd17, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b9, 5'd8, 27'h00000364, 5'd28, 27'h0000026a, 32'h00000400,
  1'd1,  5'd29, 27'h0000020f, 5'd15, 27'h0000024e, 5'd7, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000d8, 5'd17, 27'h0000017d, 5'd18, 27'h0000037c, 32'h00000400,
  1'd1,  5'd27, 27'h00000238, 5'd18, 27'h00000393, 5'd30, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000de, 5'd30, 27'h000001fc, 5'd7, 27'h00000335, 32'h00000400,
  1'd1,  5'd28, 27'h000001c9, 5'd29, 27'h00000144, 5'd17, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000139, 5'd29, 27'h0000018b, 5'd29, 27'h000003fd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000296, 5'd0, 27'h00000246, 5'd0, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000030b, 5'd4, 27'h0000012c, 5'd11, 27'h000002a2, 32'h00000400,
  1'd1,  5'd0, 27'h0000001a, 5'd2, 27'h0000022b, 5'd22, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000069, 5'd12, 27'h00000026, 5'd2, 27'h00000391, 32'h00000400,
  1'd1,  5'd0, 27'h00000246, 5'd13, 27'h00000206, 5'd12, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000163, 5'd14, 27'h00000364, 5'd20, 27'h00000338, 32'h00000400,
  1'd1,  5'd2, 27'h000002ca, 5'd25, 27'h00000040, 5'd0, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000084, 5'd22, 27'h000001c5, 5'd13, 27'h000003a0, 32'h00000400,
  1'd1,  5'd1, 27'h00000229, 5'd25, 27'h0000019f, 5'd21, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025f, 5'd1, 27'h0000005d, 5'd1, 27'h00000322, 32'h00000400,
  1'd1,  5'd14, 27'h0000035e, 5'd3, 27'h000003d4, 5'd12, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001c4, 5'd4, 27'h000000e5, 5'd25, 27'h00000172, 32'h00000400,
  1'd1,  5'd12, 27'h000002d2, 5'd14, 27'h000003f2, 5'd4, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000029d, 5'd14, 27'h000001e9, 5'd11, 27'h00000164, 32'h00000400,
  1'd1,  5'd13, 27'h0000008f, 5'd12, 27'h00000269, 5'd23, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000032e, 5'd21, 27'h0000011f, 5'd2, 27'h000000c8, 32'h00000400,
  1'd1,  5'd12, 27'h0000037b, 5'd25, 27'h000000bd, 5'd13, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000271, 5'd24, 27'h000003ed, 5'd24, 27'h00000350, 32'h00000400,
  1'd1,  5'd22, 27'h0000013f, 5'd4, 27'h0000029a, 5'd0, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000038a, 5'd2, 27'h0000026d, 5'd12, 27'h000003b4, 32'h00000400,
  1'd1,  5'd25, 27'h00000324, 5'd5, 27'h00000096, 5'd21, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000005d, 5'd10, 27'h000002b3, 5'd1, 27'h000001a4, 32'h00000400,
  1'd1,  5'd25, 27'h00000325, 5'd14, 27'h000001ae, 5'd10, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000151, 5'd14, 27'h000000c0, 5'd24, 27'h000001f3, 32'h00000400,
  1'd1,  5'd22, 27'h000000f3, 5'd22, 27'h00000370, 5'd4, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000027f, 5'd25, 27'h0000013b, 5'd10, 27'h000001e7, 32'h00000400,
  1'd1,  5'd24, 27'h000003e9, 5'd23, 27'h00000229, 5'd24, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000033f, 5'd2, 27'h0000027a, 5'd5, 27'h00000245, 32'h00000400,
  1'd1,  5'd3, 27'h00000372, 5'd3, 27'h0000038c, 5'd17, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000399, 5'd0, 27'h000001ea, 5'd29, 27'h00000142, 32'h00000400,
  1'd1,  5'd1, 27'h00000081, 5'd10, 27'h000001d6, 5'd8, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000400, 5'd13, 27'h0000019d, 5'd20, 27'h0000006f, 32'h00000400,
  1'd1,  5'd1, 27'h000001fb, 5'd15, 27'h0000007f, 5'd29, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000259, 5'd20, 27'h0000033e, 5'd5, 27'h00000294, 32'h00000400,
  1'd1,  5'd4, 27'h00000123, 5'd23, 27'h00000176, 5'd17, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001bd, 5'd21, 27'h0000027e, 5'd29, 27'h00000015, 32'h00000400,
  1'd1,  5'd13, 27'h0000010f, 5'd0, 27'h0000025a, 5'd9, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d0, 5'd3, 27'h000000b6, 5'd18, 27'h00000067, 32'h00000400,
  1'd1,  5'd14, 27'h000003f2, 5'd3, 27'h000003f5, 5'd27, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f4, 5'd14, 27'h00000285, 5'd6, 27'h000003a2, 32'h00000400,
  1'd1,  5'd12, 27'h0000009a, 5'd11, 27'h00000137, 5'd16, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002d2, 5'd12, 27'h000000c8, 5'd27, 27'h000001d1, 32'h00000400,
  1'd1,  5'd14, 27'h000003b8, 5'd21, 27'h000000fd, 5'd9, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c0, 5'd25, 27'h00000071, 5'd18, 27'h000000db, 32'h00000400,
  1'd1,  5'd12, 27'h00000275, 5'd21, 27'h000003da, 5'd29, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000197, 5'd2, 27'h00000177, 5'd6, 27'h0000011d, 32'h00000400,
  1'd1,  5'd22, 27'h000001dd, 5'd1, 27'h000000dc, 5'd19, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000171, 5'd4, 27'h00000159, 5'd28, 27'h00000055, 32'h00000400,
  1'd1,  5'd25, 27'h000000f9, 5'd14, 27'h00000190, 5'd8, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000390, 5'd11, 27'h000002c4, 5'd15, 27'h000003fa, 32'h00000400,
  1'd1,  5'd23, 27'h0000001e, 5'd15, 27'h00000030, 5'd30, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000138, 5'd24, 27'h00000241, 5'd6, 27'h00000371, 32'h00000400,
  1'd1,  5'd20, 27'h000002c6, 5'd24, 27'h000002d4, 5'd17, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003ab, 5'd24, 27'h00000268, 5'd26, 27'h000000a4, 32'h00000400,
  1'd1,  5'd1, 27'h000000bb, 5'd9, 27'h0000003b, 5'd0, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005a, 5'd7, 27'h00000053, 5'd13, 27'h000003eb, 32'h00000400,
  1'd1,  5'd4, 27'h00000384, 5'd7, 27'h00000020, 5'd21, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000315, 5'd20, 27'h000000db, 5'd5, 27'h000000a0, 32'h00000400,
  1'd1,  5'd1, 27'h000003c0, 5'd16, 27'h0000039a, 5'd10, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002c0, 5'd18, 27'h00000254, 5'd23, 27'h00000263, 32'h00000400,
  1'd1,  5'd4, 27'h0000011b, 5'd28, 27'h00000311, 5'd0, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000096, 5'd26, 27'h00000014, 5'd14, 27'h00000104, 32'h00000400,
  1'd1,  5'd4, 27'h000001ce, 5'd26, 27'h000003ae, 5'd22, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000033c, 5'd7, 27'h00000371, 5'd0, 27'h0000026d, 32'h00000400,
  1'd1,  5'd13, 27'h000000c9, 5'd10, 27'h0000003e, 5'd11, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000392, 5'd7, 27'h000001b2, 5'd22, 27'h00000271, 32'h00000400,
  1'd1,  5'd11, 27'h000003a5, 5'd20, 27'h0000005c, 5'd3, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000094, 5'd18, 27'h000000ac, 5'd13, 27'h00000348, 32'h00000400,
  1'd1,  5'd10, 27'h00000229, 5'd18, 27'h00000168, 5'd20, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000001f, 5'd28, 27'h00000205, 5'd0, 27'h000002b4, 32'h00000400,
  1'd1,  5'd11, 27'h000002ca, 5'd29, 27'h00000258, 5'd11, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000252, 5'd27, 27'h000000ee, 5'd23, 27'h00000134, 32'h00000400,
  1'd1,  5'd25, 27'h000001b3, 5'd6, 27'h0000019b, 5'd1, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000024b, 5'd9, 27'h00000283, 5'd11, 27'h00000082, 32'h00000400,
  1'd1,  5'd21, 27'h00000274, 5'd7, 27'h0000015a, 5'd25, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000391, 5'd20, 27'h000000ee, 5'd4, 27'h0000033d, 32'h00000400,
  1'd1,  5'd22, 27'h000000a9, 5'd19, 27'h000001e9, 5'd14, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000251, 5'd19, 27'h00000336, 5'd22, 27'h000000cd, 32'h00000400,
  1'd1,  5'd25, 27'h00000246, 5'd29, 27'h0000035b, 5'd4, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000039c, 5'd29, 27'h0000031c, 5'd11, 27'h00000357, 32'h00000400,
  1'd1,  5'd24, 27'h000001b5, 5'd29, 27'h0000015b, 5'd25, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000257, 5'd6, 27'h00000300, 5'd8, 27'h000003b5, 32'h00000400,
  1'd1,  5'd2, 27'h00000020, 5'd7, 27'h000000d8, 5'd19, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001cd, 5'd8, 27'h00000387, 5'd30, 27'h00000275, 32'h00000400,
  1'd1,  5'd0, 27'h0000002a, 5'd18, 27'h000003a1, 5'd5, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000066, 5'd19, 27'h00000139, 5'd17, 27'h00000339, 32'h00000400,
  1'd1,  5'd3, 27'h000002b8, 5'd19, 27'h00000150, 5'd26, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003e3, 5'd28, 27'h000001a1, 5'd8, 27'h0000028f, 32'h00000400,
  1'd1,  5'd4, 27'h000002ac, 5'd25, 27'h000003ee, 5'd17, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000086, 5'd28, 27'h000003c2, 5'd30, 27'h00000281, 32'h00000400,
  1'd1,  5'd12, 27'h000002b0, 5'd6, 27'h00000109, 5'd8, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000133, 5'd6, 27'h00000219, 5'd19, 27'h000001f2, 32'h00000400,
  1'd1,  5'd12, 27'h000002a1, 5'd9, 27'h00000165, 5'd29, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000309, 5'd18, 27'h00000170, 5'd7, 27'h000002a6, 32'h00000400,
  1'd1,  5'd12, 27'h00000108, 5'd20, 27'h00000257, 5'd18, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f1, 5'd20, 27'h0000010d, 5'd30, 27'h000001c2, 32'h00000400,
  1'd1,  5'd13, 27'h000003dc, 5'd29, 27'h00000302, 5'd6, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000018a, 5'd28, 27'h0000012b, 5'd15, 27'h00000353, 32'h00000400,
  1'd1,  5'd13, 27'h00000033, 5'd30, 27'h0000006e, 5'd29, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000040, 5'd10, 27'h000000aa, 5'd8, 27'h0000004c, 32'h00000400,
  1'd1,  5'd23, 27'h0000001a, 5'd9, 27'h00000297, 5'd15, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ed, 5'd8, 27'h0000027e, 5'd26, 27'h0000023b, 32'h00000400,
  1'd1,  5'd22, 27'h000001e3, 5'd17, 27'h00000292, 5'd7, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003e4, 5'd16, 27'h000003ac, 5'd19, 27'h00000295, 32'h00000400,
  1'd1,  5'd25, 27'h00000109, 5'd18, 27'h0000018e, 5'd26, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000018f, 5'd28, 27'h000001f8, 5'd5, 27'h000002db, 32'h00000400,
  1'd1,  5'd21, 27'h000000a7, 5'd28, 27'h000003c3, 5'd18, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e0, 5'd30, 27'h0000019e, 5'd30, 27'h0000011a, 32'h00000400,
  1'd1,  5'd9, 27'h00000002, 5'd2, 27'h0000017c, 5'd9, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000021d, 5'd0, 27'h0000022d, 5'd16, 27'h00000057, 32'h00000400,
  1'd1,  5'd5, 27'h000001bf, 5'd2, 27'h000001ec, 5'd26, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d7, 5'd12, 27'h0000005f, 5'd2, 27'h0000032b, 32'h00000400,
  1'd1,  5'd9, 27'h000002ba, 5'd14, 27'h0000012a, 5'd14, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000169, 5'd10, 27'h0000037d, 5'd21, 27'h000002a5, 32'h00000400,
  1'd1,  5'd7, 27'h00000176, 5'd21, 27'h0000023e, 5'd2, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000af, 5'd24, 27'h00000332, 5'd12, 27'h0000031f, 32'h00000400,
  1'd1,  5'd10, 27'h00000130, 5'd24, 27'h0000014e, 5'd21, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002a3, 5'd3, 27'h00000221, 5'd8, 27'h000001fb, 32'h00000400,
  1'd1,  5'd17, 27'h0000036c, 5'd0, 27'h000002b6, 5'd18, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000011a, 5'd1, 27'h0000014e, 5'd26, 27'h00000269, 32'h00000400,
  1'd1,  5'd20, 27'h0000007f, 5'd12, 27'h00000322, 5'd1, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000aa, 5'd10, 27'h00000174, 5'd11, 27'h0000033d, 32'h00000400,
  1'd1,  5'd15, 27'h0000028c, 5'd13, 27'h0000012f, 5'd25, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000094, 5'd24, 27'h000001de, 5'd4, 27'h00000186, 32'h00000400,
  1'd1,  5'd17, 27'h00000352, 5'd22, 27'h0000008c, 5'd14, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c7, 5'd23, 27'h000001d7, 5'd23, 27'h00000080, 32'h00000400,
  1'd1,  5'd27, 27'h000001eb, 5'd3, 27'h00000156, 5'd0, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000136, 5'd4, 27'h00000282, 5'd12, 27'h00000088, 32'h00000400,
  1'd1,  5'd26, 27'h00000088, 5'd2, 27'h00000056, 5'd22, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a8, 5'd15, 27'h00000009, 5'd3, 27'h00000282, 32'h00000400,
  1'd1,  5'd27, 27'h000003ac, 5'd10, 27'h000001eb, 5'd13, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021a, 5'd12, 27'h000001d3, 5'd25, 27'h00000049, 32'h00000400,
  1'd1,  5'd28, 27'h00000376, 5'd20, 27'h00000389, 5'd4, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001e7, 5'd25, 27'h0000011c, 5'd15, 27'h000001fd, 32'h00000400,
  1'd1,  5'd30, 27'h000000ee, 5'd24, 27'h00000342, 5'd25, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c1, 5'd3, 27'h0000002e, 5'd2, 27'h00000328, 32'h00000400,
  1'd1,  5'd7, 27'h000001bc, 5'd1, 27'h0000038d, 5'd10, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001bc, 5'd1, 27'h000001fe, 5'd24, 27'h000002de, 32'h00000400,
  1'd1,  5'd8, 27'h000000ad, 5'd12, 27'h00000260, 5'd10, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000009a, 5'd12, 27'h000002ba, 5'd16, 27'h000003c0, 32'h00000400,
  1'd1,  5'd6, 27'h000001ba, 5'd14, 27'h00000241, 5'd27, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000050, 5'd22, 27'h000001ea, 5'd5, 27'h000000bb, 32'h00000400,
  1'd1,  5'd8, 27'h000003fd, 5'd23, 27'h00000347, 5'd15, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000053, 5'd24, 27'h00000105, 5'd29, 27'h000003de, 32'h00000400,
  1'd1,  5'd20, 27'h0000014d, 5'd5, 27'h00000034, 5'd0, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a8, 5'd3, 27'h000002ee, 5'd11, 27'h000003e8, 32'h00000400,
  1'd1,  5'd16, 27'h00000279, 5'd3, 27'h00000132, 5'd24, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000253, 5'd11, 27'h000002aa, 5'd5, 27'h000001ce, 32'h00000400,
  1'd1,  5'd16, 27'h000000af, 5'd14, 27'h0000019d, 5'd16, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000002, 5'd14, 27'h0000031b, 5'd28, 27'h000000e0, 32'h00000400,
  1'd1,  5'd19, 27'h00000263, 5'd21, 27'h000000df, 5'd9, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000363, 5'd23, 27'h000003f1, 5'd17, 27'h00000085, 32'h00000400,
  1'd1,  5'd19, 27'h000002f3, 5'd21, 27'h00000121, 5'd28, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019d, 5'd0, 27'h0000018a, 5'd9, 27'h000001ee, 32'h00000400,
  1'd1,  5'd29, 27'h00000399, 5'd1, 27'h000002bb, 5'd19, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000010e, 5'd4, 27'h000002e7, 5'd26, 27'h00000259, 32'h00000400,
  1'd1,  5'd30, 27'h00000267, 5'd13, 27'h000000db, 5'd7, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f7, 5'd11, 27'h000001f7, 5'd16, 27'h000000cb, 32'h00000400,
  1'd1,  5'd26, 27'h000000ed, 5'd11, 27'h0000003d, 5'd26, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000013, 5'd23, 27'h000003dc, 5'd8, 27'h00000069, 32'h00000400,
  1'd1,  5'd26, 27'h0000011b, 5'd21, 27'h00000202, 5'd19, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000087, 5'd24, 27'h00000121, 5'd30, 27'h00000192, 32'h00000400,
  1'd1,  5'd5, 27'h0000026d, 5'd6, 27'h000001b3, 5'd1, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ac, 5'd8, 27'h00000373, 5'd13, 27'h00000185, 32'h00000400,
  1'd1,  5'd7, 27'h0000032a, 5'd6, 27'h00000313, 5'd25, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000065, 5'd20, 27'h00000279, 5'd0, 27'h00000070, 32'h00000400,
  1'd1,  5'd9, 27'h00000240, 5'd18, 27'h000000f9, 5'd11, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000014b, 5'd16, 27'h0000010f, 5'd21, 27'h00000224, 32'h00000400,
  1'd1,  5'd9, 27'h000001f4, 5'd29, 27'h000003ba, 5'd1, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000395, 5'd26, 27'h00000264, 5'd14, 27'h0000030a, 32'h00000400,
  1'd1,  5'd6, 27'h00000143, 5'd28, 27'h000000e9, 5'd22, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a0, 5'd8, 27'h00000108, 5'd2, 27'h000001cc, 32'h00000400,
  1'd1,  5'd15, 27'h00000231, 5'd9, 27'h000003f3, 5'd13, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001cc, 5'd6, 27'h0000036c, 5'd22, 27'h00000395, 32'h00000400,
  1'd1,  5'd17, 27'h0000025b, 5'd15, 27'h000003e8, 5'd3, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000090, 5'd17, 27'h0000000c, 5'd13, 27'h0000022e, 32'h00000400,
  1'd1,  5'd15, 27'h00000275, 5'd15, 27'h00000371, 5'd23, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001cf, 5'd27, 27'h0000003a, 5'd1, 27'h000000c4, 32'h00000400,
  1'd1,  5'd16, 27'h000001fe, 5'd25, 27'h000003e9, 5'd15, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000321, 5'd30, 27'h00000312, 5'd25, 27'h00000087, 32'h00000400,
  1'd1,  5'd30, 27'h0000020f, 5'd8, 27'h00000260, 5'd2, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002b8, 5'd6, 27'h0000001c, 5'd14, 27'h0000009a, 32'h00000400,
  1'd1,  5'd26, 27'h000000d2, 5'd8, 27'h00000247, 5'd23, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000285, 5'd15, 27'h00000391, 5'd0, 27'h00000218, 32'h00000400,
  1'd1,  5'd27, 27'h000001c5, 5'd16, 27'h000001e6, 5'd11, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000015b, 5'd16, 27'h000000eb, 5'd22, 27'h0000008d, 32'h00000400,
  1'd1,  5'd27, 27'h0000036d, 5'd29, 27'h00000264, 5'd2, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ea, 5'd27, 27'h0000013c, 5'd14, 27'h00000029, 32'h00000400,
  1'd1,  5'd26, 27'h00000076, 5'd27, 27'h00000030, 5'd25, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000d6, 5'd9, 27'h000002b7, 5'd9, 27'h000001f1, 32'h00000400,
  1'd1,  5'd6, 27'h00000221, 5'd6, 27'h00000026, 5'd16, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000184, 5'd6, 27'h000003d8, 5'd29, 27'h00000356, 32'h00000400,
  1'd1,  5'd9, 27'h0000016c, 5'd16, 27'h0000015b, 5'd5, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000028c, 5'd20, 27'h0000002c, 5'd17, 27'h00000131, 32'h00000400,
  1'd1,  5'd5, 27'h0000037e, 5'd15, 27'h000002bd, 5'd28, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003ad, 5'd29, 27'h00000104, 5'd9, 27'h000002a1, 32'h00000400,
  1'd1,  5'd6, 27'h0000007c, 5'd27, 27'h000003f4, 5'd17, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000203, 5'd26, 27'h0000024b, 5'd29, 27'h00000050, 32'h00000400,
  1'd1,  5'd19, 27'h000002ee, 5'd5, 27'h000003f2, 5'd7, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000338, 5'd8, 27'h000000a3, 5'd15, 27'h000002bd, 32'h00000400,
  1'd1,  5'd15, 27'h00000220, 5'd7, 27'h000001c2, 5'd26, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031d, 5'd19, 27'h000002ab, 5'd10, 27'h00000091, 32'h00000400,
  1'd1,  5'd17, 27'h00000186, 5'd19, 27'h0000020e, 5'd20, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003fa, 5'd20, 27'h00000009, 5'd27, 27'h0000006f, 32'h00000400,
  1'd1,  5'd17, 27'h000000b9, 5'd26, 27'h000002d3, 5'd10, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ef, 5'd26, 27'h000000e7, 5'd20, 27'h0000026f, 32'h00000400,
  1'd1,  5'd19, 27'h0000017a, 5'd27, 27'h000003d8, 5'd27, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000172, 5'd7, 27'h000001da, 5'd6, 27'h00000214, 32'h00000400,
  1'd1,  5'd29, 27'h00000054, 5'd9, 27'h000000b4, 5'd16, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000233, 5'd9, 27'h00000090, 5'd28, 27'h000003f0, 32'h00000400,
  1'd1,  5'd27, 27'h00000072, 5'd16, 27'h000000e4, 5'd10, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000272, 5'd17, 27'h0000019f, 5'd17, 27'h00000090, 32'h00000400,
  1'd1,  5'd27, 27'h00000216, 5'd18, 27'h0000026e, 5'd27, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000029, 5'd29, 27'h0000027d, 5'd9, 27'h000002b4, 32'h00000400,
  1'd1,  5'd29, 27'h00000103, 5'd29, 27'h0000015a, 5'd20, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000065, 5'd27, 27'h0000027d, 5'd30, 27'h00000365, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000000b7, 5'd1, 27'h00000145, 5'd1, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000ae, 5'd0, 27'h000001fa, 5'd13, 27'h000002bd, 32'h00000400,
  1'd1,  5'd3, 27'h000001a5, 5'd0, 27'h000002c5, 5'd20, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000279, 5'd12, 27'h0000011e, 5'd4, 27'h000003ee, 32'h00000400,
  1'd1,  5'd1, 27'h000000ab, 5'd14, 27'h0000030c, 5'd10, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003cd, 5'd12, 27'h00000143, 5'd25, 27'h000000d7, 32'h00000400,
  1'd1,  5'd1, 27'h0000018c, 5'd23, 27'h000002c0, 5'd4, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000041, 5'd25, 27'h00000282, 5'd13, 27'h00000179, 32'h00000400,
  1'd1,  5'd3, 27'h000003fa, 5'd22, 27'h000000ef, 5'd22, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000129, 5'd3, 27'h000003ec, 5'd3, 27'h0000031f, 32'h00000400,
  1'd1,  5'd14, 27'h00000272, 5'd2, 27'h000001ec, 5'd12, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000093, 5'd0, 27'h0000012e, 5'd22, 27'h00000266, 32'h00000400,
  1'd1,  5'd10, 27'h00000211, 5'd10, 27'h00000254, 5'd2, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011f, 5'd12, 27'h000000ae, 5'd14, 27'h0000038d, 32'h00000400,
  1'd1,  5'd13, 27'h000000bc, 5'd13, 27'h0000009a, 5'd21, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000038a, 5'd22, 27'h000001ac, 5'd4, 27'h0000005e, 32'h00000400,
  1'd1,  5'd10, 27'h0000026d, 5'd22, 27'h00000338, 5'd12, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003fb, 5'd23, 27'h00000021, 5'd23, 27'h000002a8, 32'h00000400,
  1'd1,  5'd23, 27'h000003c7, 5'd4, 27'h000002f0, 5'd4, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000d9, 5'd2, 27'h0000023a, 5'd12, 27'h000001be, 32'h00000400,
  1'd1,  5'd25, 27'h00000092, 5'd2, 27'h000002e8, 5'd22, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000070, 5'd14, 27'h000003f4, 5'd4, 27'h000001ea, 32'h00000400,
  1'd1,  5'd24, 27'h00000043, 5'd11, 27'h0000010c, 5'd12, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000bf, 5'd11, 27'h000000bd, 5'd24, 27'h0000007e, 32'h00000400,
  1'd1,  5'd22, 27'h000003ac, 5'd25, 27'h00000133, 5'd5, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ab, 5'd21, 27'h000000bd, 5'd11, 27'h00000051, 32'h00000400,
  1'd1,  5'd21, 27'h0000028e, 5'd20, 27'h000003d2, 5'd22, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003c5, 5'd3, 27'h00000194, 5'd10, 27'h00000071, 32'h00000400,
  1'd1,  5'd4, 27'h00000344, 5'd2, 27'h00000148, 5'd18, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c3, 5'd4, 27'h000002a0, 5'd25, 27'h000003a1, 32'h00000400,
  1'd1,  5'd2, 27'h00000347, 5'd12, 27'h00000382, 5'd9, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032a, 5'd14, 27'h000003b4, 5'd17, 27'h0000018d, 32'h00000400,
  1'd1,  5'd1, 27'h000001a9, 5'd12, 27'h000002cc, 5'd28, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000360, 5'd23, 27'h00000051, 5'd9, 27'h0000017d, 32'h00000400,
  1'd1,  5'd0, 27'h00000370, 5'd22, 27'h00000014, 5'd20, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000bb, 5'd21, 27'h0000016f, 5'd30, 27'h0000010d, 32'h00000400,
  1'd1,  5'd10, 27'h0000018e, 5'd1, 27'h00000192, 5'd7, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002da, 5'd3, 27'h00000131, 5'd15, 27'h0000038d, 32'h00000400,
  1'd1,  5'd13, 27'h0000027b, 5'd4, 27'h000001b9, 5'd27, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002da, 5'd11, 27'h00000016, 5'd10, 27'h0000004f, 32'h00000400,
  1'd1,  5'd11, 27'h0000005f, 5'd14, 27'h00000348, 5'd17, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f0, 5'd11, 27'h00000380, 5'd28, 27'h000002a6, 32'h00000400,
  1'd1,  5'd13, 27'h00000360, 5'd22, 27'h00000133, 5'd7, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f1, 5'd21, 27'h000003b7, 5'd16, 27'h0000029e, 32'h00000400,
  1'd1,  5'd15, 27'h00000176, 5'd23, 27'h00000103, 5'd28, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003a5, 5'd3, 27'h00000388, 5'd5, 27'h00000366, 32'h00000400,
  1'd1,  5'd24, 27'h0000017f, 5'd2, 27'h000001e0, 5'd19, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000205, 5'd0, 27'h00000280, 5'd30, 27'h00000037, 32'h00000400,
  1'd1,  5'd24, 27'h00000160, 5'd12, 27'h00000119, 5'd5, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000187, 5'd13, 27'h0000039a, 5'd19, 27'h0000024e, 32'h00000400,
  1'd1,  5'd21, 27'h000002bf, 5'd12, 27'h0000008e, 5'd29, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000014d, 5'd22, 27'h0000029d, 5'd9, 27'h0000033f, 32'h00000400,
  1'd1,  5'd21, 27'h0000032b, 5'd25, 27'h00000174, 5'd19, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000365, 5'd23, 27'h00000320, 5'd25, 27'h00000378, 32'h00000400,
  1'd1,  5'd1, 27'h000001c7, 5'd9, 27'h00000324, 5'd0, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000356, 5'd9, 27'h0000016f, 5'd12, 27'h000003ca, 32'h00000400,
  1'd1,  5'd3, 27'h000003df, 5'd8, 27'h000000d6, 5'd22, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ca, 5'd16, 27'h00000120, 5'd5, 27'h00000021, 32'h00000400,
  1'd1,  5'd4, 27'h00000063, 5'd16, 27'h000003e7, 5'd10, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000089, 5'd20, 27'h00000045, 5'd21, 27'h00000335, 32'h00000400,
  1'd1,  5'd2, 27'h000003be, 5'd25, 27'h00000366, 5'd1, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028a, 5'd27, 27'h00000289, 5'd13, 27'h0000018e, 32'h00000400,
  1'd1,  5'd2, 27'h000001ae, 5'd29, 27'h0000011e, 5'd23, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003af, 5'd9, 27'h000003e8, 5'd0, 27'h000002ce, 32'h00000400,
  1'd1,  5'd12, 27'h00000251, 5'd8, 27'h00000274, 5'd15, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d0, 5'd5, 27'h000003a7, 5'd24, 27'h000001b0, 32'h00000400,
  1'd1,  5'd10, 27'h0000017a, 5'd18, 27'h0000009c, 5'd2, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001a0, 5'd16, 27'h0000019f, 5'd12, 27'h00000378, 32'h00000400,
  1'd1,  5'd12, 27'h0000002f, 5'd15, 27'h00000315, 5'd21, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009f, 5'd28, 27'h0000036b, 5'd0, 27'h00000178, 32'h00000400,
  1'd1,  5'd10, 27'h00000394, 5'd28, 27'h00000169, 5'd13, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f9, 5'd30, 27'h0000027d, 5'd20, 27'h00000382, 32'h00000400,
  1'd1,  5'd22, 27'h000003f5, 5'd9, 27'h000001ee, 5'd3, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002b5, 5'd5, 27'h000002a0, 5'd10, 27'h00000210, 32'h00000400,
  1'd1,  5'd24, 27'h000003cc, 5'd8, 27'h0000036f, 5'd23, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000204, 5'd20, 27'h0000012d, 5'd0, 27'h00000020, 32'h00000400,
  1'd1,  5'd25, 27'h000000d2, 5'd18, 27'h00000264, 5'd15, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000010, 5'd18, 27'h0000021d, 5'd23, 27'h000001ab, 32'h00000400,
  1'd1,  5'd23, 27'h000001e0, 5'd28, 27'h0000024b, 5'd4, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000361, 5'd30, 27'h000000dc, 5'd10, 27'h00000370, 32'h00000400,
  1'd1,  5'd23, 27'h000002e5, 5'd30, 27'h000001e4, 5'd25, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000256, 5'd10, 27'h00000101, 5'd7, 27'h00000353, 32'h00000400,
  1'd1,  5'd0, 27'h00000150, 5'd9, 27'h00000128, 5'd17, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000069, 5'd6, 27'h000002f4, 5'd29, 27'h00000234, 32'h00000400,
  1'd1,  5'd3, 27'h000001aa, 5'd17, 27'h000001f8, 5'd6, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d3, 5'd20, 27'h00000106, 5'd16, 27'h000000c0, 32'h00000400,
  1'd1,  5'd2, 27'h000000dd, 5'd16, 27'h000001e4, 5'd26, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000343, 5'd30, 27'h00000087, 5'd10, 27'h00000089, 32'h00000400,
  1'd1,  5'd3, 27'h000002e2, 5'd29, 27'h0000028d, 5'd20, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000cf, 5'd26, 27'h00000090, 5'd28, 27'h0000016d, 32'h00000400,
  1'd1,  5'd10, 27'h0000031a, 5'd7, 27'h0000017d, 5'd9, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c5, 5'd9, 27'h000002a5, 5'd17, 27'h00000352, 32'h00000400,
  1'd1,  5'd14, 27'h00000264, 5'd7, 27'h000002c9, 5'd27, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000383, 5'd18, 27'h0000014f, 5'd6, 27'h000000fa, 32'h00000400,
  1'd1,  5'd11, 27'h0000028b, 5'd16, 27'h00000074, 5'd16, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000010f, 5'd17, 27'h000001ed, 5'd26, 27'h000002cc, 32'h00000400,
  1'd1,  5'd13, 27'h000002cb, 5'd29, 27'h00000236, 5'd6, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003df, 5'd30, 27'h00000042, 5'd17, 27'h000002b6, 32'h00000400,
  1'd1,  5'd14, 27'h00000010, 5'd30, 27'h00000281, 5'd28, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000269, 5'd7, 27'h000000ec, 5'd8, 27'h0000014e, 32'h00000400,
  1'd1,  5'd25, 27'h0000017b, 5'd7, 27'h000003f9, 5'd16, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000236, 5'd9, 27'h000002d9, 5'd30, 27'h0000034c, 32'h00000400,
  1'd1,  5'd23, 27'h0000032e, 5'd16, 27'h00000090, 5'd6, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000098, 5'd15, 27'h00000357, 5'd18, 27'h000000c4, 32'h00000400,
  1'd1,  5'd20, 27'h00000320, 5'd16, 27'h000001a4, 5'd27, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000004, 5'd30, 27'h000002d6, 5'd9, 27'h00000044, 32'h00000400,
  1'd1,  5'd22, 27'h00000239, 5'd30, 27'h0000007f, 5'd16, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000355, 5'd29, 27'h00000019, 5'd29, 27'h00000398, 32'h00000400,
  1'd1,  5'd7, 27'h0000017d, 5'd3, 27'h0000009a, 5'd8, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000019d, 5'd2, 27'h000003a4, 5'd16, 27'h00000079, 32'h00000400,
  1'd1,  5'd7, 27'h00000059, 5'd0, 27'h00000058, 5'd25, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ab, 5'd11, 27'h0000005b, 5'd2, 27'h000001f8, 32'h00000400,
  1'd1,  5'd10, 27'h0000006e, 5'd13, 27'h00000030, 5'd15, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000007d, 5'd11, 27'h0000013c, 5'd21, 27'h00000189, 32'h00000400,
  1'd1,  5'd7, 27'h000000e1, 5'd22, 27'h000003ab, 5'd4, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b0, 5'd21, 27'h00000331, 5'd13, 27'h0000011e, 32'h00000400,
  1'd1,  5'd7, 27'h000003ea, 5'd21, 27'h000001f4, 5'd22, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000030e, 5'd4, 27'h00000158, 5'd8, 27'h0000015e, 32'h00000400,
  1'd1,  5'd17, 27'h000002fe, 5'd3, 27'h000001f5, 5'd20, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000bb, 5'd3, 27'h00000244, 5'd30, 27'h000003a1, 32'h00000400,
  1'd1,  5'd16, 27'h000000f5, 5'd13, 27'h00000146, 5'd2, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ec, 5'd11, 27'h00000269, 5'd11, 27'h00000208, 32'h00000400,
  1'd1,  5'd16, 27'h000001ce, 5'd12, 27'h0000032a, 5'd25, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001cf, 5'd20, 27'h0000031d, 5'd0, 27'h000000bb, 32'h00000400,
  1'd1,  5'd16, 27'h00000123, 5'd24, 27'h000001d8, 5'd11, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000001b, 5'd23, 27'h000003cb, 5'd25, 27'h000001f6, 32'h00000400,
  1'd1,  5'd28, 27'h0000021e, 5'd2, 27'h000000b8, 5'd4, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c6, 5'd4, 27'h0000023a, 5'd12, 27'h000000e4, 32'h00000400,
  1'd1,  5'd27, 27'h000001c5, 5'd0, 27'h000002e5, 5'd20, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002bd, 5'd11, 27'h0000000e, 5'd2, 27'h00000070, 32'h00000400,
  1'd1,  5'd30, 27'h000003f0, 5'd12, 27'h000000c0, 5'd14, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000358, 5'd11, 27'h0000032c, 5'd21, 27'h000003fd, 32'h00000400,
  1'd1,  5'd28, 27'h0000007b, 5'd22, 27'h00000344, 5'd0, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002e3, 5'd21, 27'h0000012f, 5'd11, 27'h0000019e, 32'h00000400,
  1'd1,  5'd26, 27'h0000005d, 5'd22, 27'h000003a3, 5'd24, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d7, 5'd0, 27'h000000ce, 5'd3, 27'h00000322, 32'h00000400,
  1'd1,  5'd8, 27'h0000005b, 5'd0, 27'h00000271, 5'd14, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000028a, 5'd5, 27'h00000090, 5'd21, 27'h000000a9, 32'h00000400,
  1'd1,  5'd10, 27'h000000a9, 5'd13, 27'h0000011d, 5'd5, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000029, 5'd10, 27'h00000339, 5'd19, 27'h000003b9, 32'h00000400,
  1'd1,  5'd7, 27'h00000379, 5'd11, 27'h00000038, 5'd27, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000039d, 5'd21, 27'h00000094, 5'd10, 27'h00000090, 32'h00000400,
  1'd1,  5'd5, 27'h0000035c, 5'd21, 27'h0000005e, 5'd16, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000257, 5'd21, 27'h000002a4, 5'd29, 27'h00000027, 32'h00000400,
  1'd1,  5'd20, 27'h00000114, 5'd4, 27'h0000023a, 5'd3, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d4, 5'd1, 27'h0000000c, 5'd10, 27'h000001f4, 32'h00000400,
  1'd1,  5'd16, 27'h000001bb, 5'd2, 27'h000003b0, 5'd25, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000de, 5'd14, 27'h00000389, 5'd7, 27'h0000039a, 32'h00000400,
  1'd1,  5'd15, 27'h00000253, 5'd11, 27'h00000034, 5'd17, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000037b, 5'd11, 27'h00000372, 5'd29, 27'h00000073, 32'h00000400,
  1'd1,  5'd17, 27'h0000021e, 5'd22, 27'h000000a3, 5'd9, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000022, 5'd23, 27'h00000128, 5'd15, 27'h00000296, 32'h00000400,
  1'd1,  5'd17, 27'h000003e6, 5'd23, 27'h000000ce, 5'd29, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000258, 5'd0, 27'h000003e5, 5'd8, 27'h000003ea, 32'h00000400,
  1'd1,  5'd29, 27'h00000280, 5'd2, 27'h0000035b, 5'd18, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000007, 5'd1, 27'h000002ec, 5'd30, 27'h000001f3, 32'h00000400,
  1'd1,  5'd29, 27'h000001f2, 5'd12, 27'h000003c2, 5'd6, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001f9, 5'd10, 27'h0000033d, 5'd16, 27'h00000147, 32'h00000400,
  1'd1,  5'd27, 27'h000003a7, 5'd13, 27'h0000003d, 5'd29, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000ea, 5'd22, 27'h0000008f, 5'd9, 27'h00000126, 32'h00000400,
  1'd1,  5'd27, 27'h00000329, 5'd21, 27'h0000023e, 5'd19, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000329, 5'd23, 27'h000000ff, 5'd30, 27'h0000028c, 32'h00000400,
  1'd1,  5'd6, 27'h00000018, 5'd6, 27'h00000168, 5'd4, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000172, 5'd5, 27'h0000029c, 5'd14, 27'h00000128, 32'h00000400,
  1'd1,  5'd5, 27'h00000211, 5'd8, 27'h00000034, 5'd25, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ed, 5'd17, 27'h00000354, 5'd1, 27'h00000203, 32'h00000400,
  1'd1,  5'd8, 27'h000003ff, 5'd18, 27'h0000018d, 5'd12, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000006c, 5'd18, 27'h0000016e, 5'd24, 27'h000000fb, 32'h00000400,
  1'd1,  5'd6, 27'h00000200, 5'd26, 27'h000000c9, 5'd2, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000104, 5'd30, 27'h0000028f, 5'd11, 27'h00000318, 32'h00000400,
  1'd1,  5'd5, 27'h000002e9, 5'd27, 27'h00000177, 5'd24, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011e, 5'd5, 27'h000003a2, 5'd3, 27'h000003ed, 32'h00000400,
  1'd1,  5'd19, 27'h000000a0, 5'd9, 27'h00000258, 5'd14, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000028c, 5'd10, 27'h000000f8, 5'd22, 27'h000000da, 32'h00000400,
  1'd1,  5'd18, 27'h000000ce, 5'd16, 27'h000000e8, 5'd2, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000020c, 5'd19, 27'h0000013b, 5'd15, 27'h000000a6, 32'h00000400,
  1'd1,  5'd18, 27'h0000000e, 5'd17, 27'h0000039d, 5'd22, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025b, 5'd30, 27'h00000072, 5'd3, 27'h00000170, 32'h00000400,
  1'd1,  5'd17, 27'h000000d4, 5'd30, 27'h0000000d, 5'd12, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021a, 5'd30, 27'h0000034a, 5'd22, 27'h000001af, 32'h00000400,
  1'd1,  5'd29, 27'h000003b0, 5'd7, 27'h0000022f, 5'd4, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000293, 5'd9, 27'h00000360, 5'd10, 27'h0000022e, 32'h00000400,
  1'd1,  5'd26, 27'h00000364, 5'd8, 27'h000003cc, 5'd21, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000299, 5'd18, 27'h00000389, 5'd2, 27'h000000c4, 32'h00000400,
  1'd1,  5'd30, 27'h0000002d, 5'd16, 27'h00000032, 5'd10, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000005b, 5'd16, 27'h00000025, 5'd23, 27'h00000191, 32'h00000400,
  1'd1,  5'd29, 27'h00000193, 5'd29, 27'h0000014c, 5'd2, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003d0, 5'd29, 27'h00000385, 5'd11, 27'h00000262, 32'h00000400,
  1'd1,  5'd29, 27'h000002f3, 5'd27, 27'h00000149, 5'd21, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000380, 5'd5, 27'h00000141, 5'd9, 27'h00000037, 32'h00000400,
  1'd1,  5'd9, 27'h00000226, 5'd9, 27'h0000016e, 5'd17, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000006d, 5'd8, 27'h000000e7, 5'd26, 27'h0000014a, 32'h00000400,
  1'd1,  5'd8, 27'h0000015f, 5'd19, 27'h0000023c, 5'd9, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009e, 5'd18, 27'h000001dd, 5'd18, 27'h00000078, 32'h00000400,
  1'd1,  5'd6, 27'h0000027a, 5'd19, 27'h0000037e, 5'd27, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001f3, 5'd27, 27'h0000039f, 5'd9, 27'h00000239, 32'h00000400,
  1'd1,  5'd7, 27'h00000019, 5'd29, 27'h000003c5, 5'd16, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000176, 5'd27, 27'h00000272, 5'd29, 27'h0000022d, 32'h00000400,
  1'd1,  5'd15, 27'h000002a5, 5'd8, 27'h0000024b, 5'd9, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b0, 5'd9, 27'h0000024c, 5'd18, 27'h000000f3, 32'h00000400,
  1'd1,  5'd16, 27'h00000314, 5'd5, 27'h0000034d, 5'd30, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ca, 5'd15, 27'h0000036a, 5'd8, 27'h000002e0, 32'h00000400,
  1'd1,  5'd20, 27'h0000016a, 5'd20, 27'h0000000c, 5'd18, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000394, 5'd15, 27'h00000362, 5'd28, 27'h000003ba, 32'h00000400,
  1'd1,  5'd16, 27'h000002a3, 5'd28, 27'h0000034e, 5'd5, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002be, 5'd28, 27'h00000316, 5'd16, 27'h00000074, 32'h00000400,
  1'd1,  5'd18, 27'h000000a9, 5'd27, 27'h000003d0, 5'd28, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000037c, 5'd6, 27'h00000396, 5'd10, 27'h00000139, 32'h00000400,
  1'd1,  5'd27, 27'h0000018a, 5'd6, 27'h0000028e, 5'd15, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f8, 5'd8, 27'h00000199, 5'd25, 27'h000003d9, 32'h00000400,
  1'd1,  5'd27, 27'h00000378, 5'd17, 27'h000001ff, 5'd8, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000033e, 5'd17, 27'h0000019b, 5'd16, 27'h00000338, 32'h00000400,
  1'd1,  5'd28, 27'h000003cd, 5'd19, 27'h000003ca, 5'd30, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000081, 5'd29, 27'h0000038d, 5'd5, 27'h000003de, 32'h00000400,
  1'd1,  5'd30, 27'h000000ef, 5'd30, 27'h00000391, 5'd19, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003aa, 5'd30, 27'h0000004a, 5'd26, 27'h00000251, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h0000008f, 5'd2, 27'h000001be, 5'd2, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029b, 5'd1, 27'h0000025f, 5'd11, 27'h000002b5, 32'h00000400,
  1'd1,  5'd0, 27'h00000083, 5'd2, 27'h00000365, 5'd25, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000030e, 5'd10, 27'h00000341, 5'd4, 27'h00000234, 32'h00000400,
  1'd1,  5'd0, 27'h000000e3, 5'd15, 27'h00000169, 5'd12, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000086, 5'd11, 27'h0000032b, 5'd21, 27'h00000301, 32'h00000400,
  1'd1,  5'd0, 27'h0000003b, 5'd23, 27'h00000391, 5'd4, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ed, 5'd20, 27'h00000356, 5'd13, 27'h00000299, 32'h00000400,
  1'd1,  5'd3, 27'h0000021e, 5'd25, 27'h0000021b, 5'd21, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e3, 5'd1, 27'h00000386, 5'd4, 27'h00000008, 32'h00000400,
  1'd1,  5'd10, 27'h000002f1, 5'd4, 27'h000003e0, 5'd13, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001b3, 5'd1, 27'h00000263, 5'd22, 27'h00000127, 32'h00000400,
  1'd1,  5'd13, 27'h00000158, 5'd13, 27'h00000340, 5'd1, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c9, 5'd13, 27'h000001ae, 5'd12, 27'h000001ff, 32'h00000400,
  1'd1,  5'd13, 27'h000003cb, 5'd15, 27'h0000008b, 5'd23, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000240, 5'd23, 27'h00000261, 5'd3, 27'h000000c8, 32'h00000400,
  1'd1,  5'd10, 27'h000003f1, 5'd21, 27'h0000036e, 5'd12, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003ec, 5'd23, 27'h000000e9, 5'd24, 27'h0000016d, 32'h00000400,
  1'd1,  5'd22, 27'h0000023e, 5'd2, 27'h0000024e, 5'd2, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000f0, 5'd2, 27'h00000200, 5'd12, 27'h000003fc, 32'h00000400,
  1'd1,  5'd22, 27'h00000320, 5'd1, 27'h00000021, 5'd21, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d8, 5'd12, 27'h00000277, 5'd3, 27'h00000087, 32'h00000400,
  1'd1,  5'd23, 27'h000000a8, 5'd13, 27'h000003e4, 5'd12, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000c4, 5'd11, 27'h000001aa, 5'd20, 27'h00000383, 32'h00000400,
  1'd1,  5'd25, 27'h00000218, 5'd23, 27'h00000030, 5'd1, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e1, 5'd24, 27'h000002f0, 5'd13, 27'h00000270, 32'h00000400,
  1'd1,  5'd23, 27'h00000308, 5'd24, 27'h000002bb, 5'd25, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000003c, 5'd4, 27'h00000063, 5'd9, 27'h00000056, 32'h00000400,
  1'd1,  5'd3, 27'h00000133, 5'd4, 27'h00000052, 5'd16, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000024a, 5'd1, 27'h000001ab, 5'd29, 27'h000000ad, 32'h00000400,
  1'd1,  5'd4, 27'h00000371, 5'd10, 27'h000003d6, 5'd5, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000204, 5'd14, 27'h000000c2, 5'd16, 27'h000002a0, 32'h00000400,
  1'd1,  5'd3, 27'h000002ba, 5'd12, 27'h0000011b, 5'd25, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000f8, 5'd24, 27'h00000262, 5'd9, 27'h000000cd, 32'h00000400,
  1'd1,  5'd2, 27'h0000008c, 5'd21, 27'h0000016b, 5'd16, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d0, 5'd21, 27'h000003ce, 5'd28, 27'h000003f9, 32'h00000400,
  1'd1,  5'd11, 27'h000002cd, 5'd0, 27'h00000163, 5'd6, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000186, 5'd1, 27'h000003e1, 5'd20, 27'h00000064, 32'h00000400,
  1'd1,  5'd13, 27'h0000018d, 5'd2, 27'h0000035a, 5'd26, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c8, 5'd15, 27'h000001c5, 5'd5, 27'h000003b8, 32'h00000400,
  1'd1,  5'd14, 27'h00000193, 5'd15, 27'h0000001d, 5'd18, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ea, 5'd11, 27'h000002b3, 5'd30, 27'h0000017d, 32'h00000400,
  1'd1,  5'd13, 27'h0000018a, 5'd25, 27'h00000343, 5'd5, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000ef, 5'd21, 27'h000002e8, 5'd18, 27'h000003aa, 32'h00000400,
  1'd1,  5'd14, 27'h00000036, 5'd23, 27'h000001fb, 5'd26, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000015f, 5'd4, 27'h0000039c, 5'd8, 27'h00000203, 32'h00000400,
  1'd1,  5'd22, 27'h0000031d, 5'd1, 27'h00000061, 5'd17, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d0, 5'd2, 27'h000002ce, 5'd29, 27'h00000365, 32'h00000400,
  1'd1,  5'd23, 27'h0000039c, 5'd12, 27'h00000333, 5'd9, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ef, 5'd15, 27'h000000fa, 5'd17, 27'h000001b8, 32'h00000400,
  1'd1,  5'd23, 27'h00000012, 5'd10, 27'h000003ac, 5'd28, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000276, 5'd22, 27'h0000026d, 5'd10, 27'h00000077, 32'h00000400,
  1'd1,  5'd23, 27'h00000094, 5'd20, 27'h000002e7, 5'd19, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000012b, 5'd21, 27'h00000379, 5'd29, 27'h000001b8, 32'h00000400,
  1'd1,  5'd3, 27'h0000018a, 5'd9, 27'h0000039a, 5'd2, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000251, 5'd7, 27'h000000b9, 5'd14, 27'h000002b4, 32'h00000400,
  1'd1,  5'd2, 27'h0000021d, 5'd5, 27'h000003bc, 5'd23, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001e3, 5'd20, 27'h00000054, 5'd1, 27'h000000e9, 32'h00000400,
  1'd1,  5'd0, 27'h000001e3, 5'd20, 27'h000000d3, 5'd11, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000090, 5'd15, 27'h000002de, 5'd24, 27'h00000391, 32'h00000400,
  1'd1,  5'd0, 27'h00000001, 5'd28, 27'h00000136, 5'd0, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001cf, 5'd29, 27'h00000089, 5'd11, 27'h00000208, 32'h00000400,
  1'd1,  5'd3, 27'h0000017b, 5'd27, 27'h0000007c, 5'd24, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000011b, 5'd6, 27'h00000061, 5'd3, 27'h00000193, 32'h00000400,
  1'd1,  5'd15, 27'h000001df, 5'd10, 27'h0000002b, 5'd15, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000216, 5'd5, 27'h0000024a, 5'd22, 27'h00000256, 32'h00000400,
  1'd1,  5'd11, 27'h00000338, 5'd18, 27'h0000003b, 5'd2, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000022, 5'd17, 27'h000003ba, 5'd14, 27'h0000024e, 32'h00000400,
  1'd1,  5'd13, 27'h000000ba, 5'd16, 27'h000003a2, 5'd25, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038e, 5'd26, 27'h000001f7, 5'd1, 27'h00000211, 32'h00000400,
  1'd1,  5'd12, 27'h000000c2, 5'd29, 27'h0000039d, 5'd15, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002c8, 5'd26, 27'h000002c2, 5'd24, 27'h0000005f, 32'h00000400,
  1'd1,  5'd22, 27'h0000034f, 5'd8, 27'h000003de, 5'd0, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a0, 5'd5, 27'h000000d1, 5'd14, 27'h0000029a, 32'h00000400,
  1'd1,  5'd21, 27'h0000005a, 5'd9, 27'h0000022a, 5'd25, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003db, 5'd16, 27'h00000026, 5'd1, 27'h000003ae, 32'h00000400,
  1'd1,  5'd24, 27'h00000225, 5'd15, 27'h00000323, 5'd15, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000046, 5'd16, 27'h00000110, 5'd21, 27'h0000029c, 32'h00000400,
  1'd1,  5'd21, 27'h00000398, 5'd29, 27'h000001a6, 5'd2, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000253, 5'd28, 27'h00000392, 5'd12, 27'h00000041, 32'h00000400,
  1'd1,  5'd24, 27'h000000a8, 5'd30, 27'h00000245, 5'd21, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000367, 5'd5, 27'h00000399, 5'd9, 27'h00000281, 32'h00000400,
  1'd1,  5'd4, 27'h000000ca, 5'd7, 27'h00000129, 5'd15, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012e, 5'd9, 27'h00000335, 5'd28, 27'h000000cf, 32'h00000400,
  1'd1,  5'd1, 27'h00000097, 5'd19, 27'h0000016c, 5'd6, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000180, 5'd15, 27'h00000330, 5'd18, 27'h0000028b, 32'h00000400,
  1'd1,  5'd0, 27'h00000110, 5'd19, 27'h000000df, 5'd30, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022c, 5'd29, 27'h000000e5, 5'd7, 27'h00000012, 32'h00000400,
  1'd1,  5'd0, 27'h00000146, 5'd28, 27'h00000083, 5'd17, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005d, 5'd28, 27'h000001d7, 5'd26, 27'h000001a3, 32'h00000400,
  1'd1,  5'd15, 27'h0000005a, 5'd6, 27'h000002b5, 5'd7, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000d8, 5'd9, 27'h00000029, 5'd15, 27'h000002ac, 32'h00000400,
  1'd1,  5'd10, 27'h000002b8, 5'd8, 27'h00000263, 5'd29, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000018c, 5'd18, 27'h00000385, 5'd7, 27'h0000012f, 32'h00000400,
  1'd1,  5'd12, 27'h000002ca, 5'd18, 27'h000000d4, 5'd15, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000372, 5'd17, 27'h00000362, 5'd28, 27'h0000000d, 32'h00000400,
  1'd1,  5'd14, 27'h00000193, 5'd27, 27'h000003ed, 5'd5, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000167, 5'd29, 27'h000002e9, 5'd15, 27'h000002f3, 32'h00000400,
  1'd1,  5'd14, 27'h0000028f, 5'd28, 27'h0000001c, 5'd28, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000076, 5'd6, 27'h000001a6, 5'd9, 27'h00000341, 32'h00000400,
  1'd1,  5'd21, 27'h0000026b, 5'd5, 27'h000002e5, 5'd17, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000023b, 5'd9, 27'h000000bc, 5'd27, 27'h000002f6, 32'h00000400,
  1'd1,  5'd22, 27'h000003cc, 5'd17, 27'h00000296, 5'd8, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ad, 5'd18, 27'h00000022, 5'd19, 27'h000002af, 32'h00000400,
  1'd1,  5'd20, 27'h000002ff, 5'd15, 27'h0000028a, 5'd28, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001c2, 5'd26, 27'h000001d1, 5'd6, 27'h000001e5, 32'h00000400,
  1'd1,  5'd21, 27'h00000248, 5'd29, 27'h000000fc, 5'd17, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b7, 5'd30, 27'h0000020d, 5'd29, 27'h000003e2, 32'h00000400,
  1'd1,  5'd8, 27'h00000031, 5'd2, 27'h0000015d, 5'd9, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002db, 5'd3, 27'h000003e1, 5'd19, 27'h00000214, 32'h00000400,
  1'd1,  5'd8, 27'h0000013b, 5'd0, 27'h0000032f, 5'd26, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000fd, 5'd10, 27'h000001e6, 5'd2, 27'h000001cc, 32'h00000400,
  1'd1,  5'd9, 27'h00000319, 5'd11, 27'h000002d4, 5'd12, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000038a, 5'd11, 27'h0000034e, 5'd21, 27'h0000018d, 32'h00000400,
  1'd1,  5'd9, 27'h0000015f, 5'd22, 27'h00000148, 5'd1, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000014c, 5'd25, 27'h00000035, 5'd14, 27'h00000075, 32'h00000400,
  1'd1,  5'd5, 27'h00000133, 5'd23, 27'h0000020b, 5'd25, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000311, 5'd1, 27'h000003f7, 5'd8, 27'h000000cb, 32'h00000400,
  1'd1,  5'd16, 27'h0000033f, 5'd2, 27'h00000211, 5'd15, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000b1, 5'd2, 27'h0000019a, 5'd29, 27'h000000b8, 32'h00000400,
  1'd1,  5'd16, 27'h00000243, 5'd12, 27'h00000115, 5'd4, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000199, 5'd11, 27'h00000329, 5'd13, 27'h00000045, 32'h00000400,
  1'd1,  5'd15, 27'h000003c6, 5'd15, 27'h00000111, 5'd24, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002fd, 5'd23, 27'h00000201, 5'd1, 27'h00000084, 32'h00000400,
  1'd1,  5'd16, 27'h00000120, 5'd21, 27'h000002be, 5'd15, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000015a, 5'd23, 27'h00000393, 5'd22, 27'h000002bd, 32'h00000400,
  1'd1,  5'd26, 27'h000001ab, 5'd1, 27'h000003a2, 5'd3, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d5, 5'd1, 27'h000002fe, 5'd13, 27'h00000222, 32'h00000400,
  1'd1,  5'd29, 27'h0000034d, 5'd4, 27'h000003f2, 5'd21, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000363, 5'd13, 27'h00000079, 5'd0, 27'h0000029c, 32'h00000400,
  1'd1,  5'd29, 27'h00000126, 5'd14, 27'h00000027, 5'd11, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001da, 5'd13, 27'h00000316, 5'd21, 27'h0000023e, 32'h00000400,
  1'd1,  5'd27, 27'h000003a9, 5'd23, 27'h0000020b, 5'd3, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000026f, 5'd24, 27'h00000079, 5'd14, 27'h00000333, 32'h00000400,
  1'd1,  5'd28, 27'h0000016e, 5'd23, 27'h000003b4, 5'd25, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000011, 5'd0, 27'h00000159, 5'd0, 27'h00000013, 32'h00000400,
  1'd1,  5'd9, 27'h00000383, 5'd4, 27'h0000028b, 5'd13, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020d, 5'd1, 27'h0000002f, 5'd22, 27'h0000005b, 32'h00000400,
  1'd1,  5'd8, 27'h00000234, 5'd11, 27'h000000e4, 5'd5, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000301, 5'd13, 27'h000003eb, 5'd16, 27'h0000000f, 32'h00000400,
  1'd1,  5'd5, 27'h0000025c, 5'd15, 27'h00000197, 5'd27, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000233, 5'd24, 27'h000003bd, 5'd10, 27'h00000128, 32'h00000400,
  1'd1,  5'd5, 27'h000002b7, 5'd25, 27'h00000069, 5'd17, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000135, 5'd21, 27'h00000369, 5'd26, 27'h00000179, 32'h00000400,
  1'd1,  5'd20, 27'h0000018a, 5'd4, 27'h00000051, 5'd1, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000008b, 5'd2, 27'h0000004c, 5'd14, 27'h0000038f, 32'h00000400,
  1'd1,  5'd15, 27'h00000320, 5'd3, 27'h0000020d, 5'd24, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000086, 5'd13, 27'h00000220, 5'd6, 27'h0000028f, 32'h00000400,
  1'd1,  5'd19, 27'h00000019, 5'd12, 27'h0000035d, 5'd19, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000097, 5'd10, 27'h0000020f, 5'd27, 27'h000003fe, 32'h00000400,
  1'd1,  5'd20, 27'h0000019e, 5'd20, 27'h000003db, 5'd9, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b3, 5'd23, 27'h0000035f, 5'd16, 27'h0000019d, 32'h00000400,
  1'd1,  5'd20, 27'h0000028b, 5'd21, 27'h00000353, 5'd26, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003f6, 5'd2, 27'h00000034, 5'd8, 27'h000001f8, 32'h00000400,
  1'd1,  5'd26, 27'h00000064, 5'd1, 27'h000002dd, 5'd16, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000007f, 5'd2, 27'h00000377, 5'd28, 27'h0000001a, 32'h00000400,
  1'd1,  5'd29, 27'h00000078, 5'd12, 27'h000001ac, 5'd9, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000bc, 5'd13, 27'h00000049, 5'd18, 27'h00000171, 32'h00000400,
  1'd1,  5'd26, 27'h00000364, 5'd11, 27'h0000034d, 5'd30, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000003, 5'd21, 27'h00000031, 5'd10, 27'h000000e2, 32'h00000400,
  1'd1,  5'd25, 27'h000003da, 5'd24, 27'h00000255, 5'd17, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003d1, 5'd25, 27'h000000f2, 5'd28, 27'h00000103, 32'h00000400,
  1'd1,  5'd8, 27'h000001df, 5'd6, 27'h000001f9, 5'd4, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002cd, 5'd9, 27'h000001a3, 5'd12, 27'h000001dc, 32'h00000400,
  1'd1,  5'd5, 27'h0000033d, 5'd6, 27'h00000389, 5'd23, 27'h00000242, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000152, 5'd17, 27'h000003c8, 5'd5, 27'h00000039, 32'h00000400,
  1'd1,  5'd9, 27'h000003e3, 5'd20, 27'h0000027e, 5'd10, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000157, 5'd20, 27'h0000013e, 5'd23, 27'h000002ba, 32'h00000400,
  1'd1,  5'd5, 27'h000001ea, 5'd29, 27'h00000399, 5'd0, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000018a, 5'd28, 27'h0000037a, 5'd14, 27'h000000c9, 32'h00000400,
  1'd1,  5'd7, 27'h00000115, 5'd29, 27'h00000151, 5'd25, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001eb, 5'd9, 27'h000003bc, 5'd2, 27'h00000180, 32'h00000400,
  1'd1,  5'd17, 27'h000001f3, 5'd8, 27'h000003b6, 5'd13, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d4, 5'd8, 27'h000000dc, 5'd21, 27'h00000090, 32'h00000400,
  1'd1,  5'd15, 27'h000003fc, 5'd16, 27'h00000195, 5'd3, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001bf, 5'd18, 27'h000001f3, 5'd14, 27'h00000285, 32'h00000400,
  1'd1,  5'd15, 27'h00000366, 5'd18, 27'h000000fd, 5'd21, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000090, 5'd27, 27'h00000140, 5'd4, 27'h0000011b, 32'h00000400,
  1'd1,  5'd15, 27'h000003fc, 5'd26, 27'h00000020, 5'd12, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d0, 5'd30, 27'h000002db, 5'd23, 27'h000001d1, 32'h00000400,
  1'd1,  5'd26, 27'h000002d8, 5'd8, 27'h000000e9, 5'd2, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000136, 5'd9, 27'h000001b9, 5'd10, 27'h0000031e, 32'h00000400,
  1'd1,  5'd30, 27'h000003d2, 5'd5, 27'h000001c8, 5'd22, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000316, 5'd20, 27'h000000d4, 5'd3, 27'h000003db, 32'h00000400,
  1'd1,  5'd27, 27'h00000041, 5'd16, 27'h00000233, 5'd15, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001aa, 5'd16, 27'h000002d7, 5'd25, 27'h000000e7, 32'h00000400,
  1'd1,  5'd28, 27'h0000002f, 5'd29, 27'h000003bb, 5'd4, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000040, 5'd27, 27'h000000eb, 5'd13, 27'h00000397, 32'h00000400,
  1'd1,  5'd30, 27'h000002f7, 5'd27, 27'h000000f7, 5'd21, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000338, 5'd6, 27'h00000324, 5'd6, 27'h000003dc, 32'h00000400,
  1'd1,  5'd10, 27'h0000009f, 5'd10, 27'h000000a2, 5'd20, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ef, 5'd9, 27'h000001ec, 5'd26, 27'h0000012a, 32'h00000400,
  1'd1,  5'd9, 27'h000002eb, 5'd17, 27'h00000004, 5'd9, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000009b, 5'd16, 27'h00000004, 5'd16, 27'h00000219, 32'h00000400,
  1'd1,  5'd6, 27'h000001d8, 5'd17, 27'h0000008c, 5'd28, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b0, 5'd29, 27'h000001e8, 5'd6, 27'h000003e8, 32'h00000400,
  1'd1,  5'd10, 27'h000000dc, 5'd27, 27'h00000106, 5'd18, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e4, 5'd28, 27'h000003d5, 5'd27, 27'h0000011b, 32'h00000400,
  1'd1,  5'd18, 27'h0000014d, 5'd7, 27'h0000030c, 5'd7, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000029d, 5'd6, 27'h000003b7, 5'd18, 27'h00000338, 32'h00000400,
  1'd1,  5'd17, 27'h00000147, 5'd8, 27'h000003e2, 5'd28, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000122, 5'd18, 27'h0000025c, 5'd7, 27'h0000039e, 32'h00000400,
  1'd1,  5'd18, 27'h00000073, 5'd17, 27'h000002b8, 5'd18, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000026e, 5'd18, 27'h000002c4, 5'd27, 27'h0000002e, 32'h00000400,
  1'd1,  5'd18, 27'h00000301, 5'd30, 27'h000002aa, 5'd7, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000039f, 5'd25, 27'h000003e3, 5'd17, 27'h00000265, 32'h00000400,
  1'd1,  5'd18, 27'h0000037b, 5'd28, 27'h000002d9, 5'd27, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000366, 5'd8, 27'h00000373, 5'd5, 27'h00000359, 32'h00000400,
  1'd1,  5'd29, 27'h000002e3, 5'd5, 27'h000003d6, 5'd18, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003d6, 5'd5, 27'h000001d5, 5'd28, 27'h00000051, 32'h00000400,
  1'd1,  5'd30, 27'h00000001, 5'd16, 27'h0000018f, 5'd7, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000023d, 5'd18, 27'h000001bc, 5'd19, 27'h00000184, 32'h00000400,
  1'd1,  5'd28, 27'h00000099, 5'd15, 27'h00000209, 5'd27, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002a2, 5'd28, 27'h00000005, 5'd5, 27'h00000325, 32'h00000400,
  1'd1,  5'd30, 27'h00000275, 5'd27, 27'h0000035d, 5'd16, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000185, 5'd27, 27'h00000281, 5'd29, 27'h00000291, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000002a6, 5'd0, 27'h000003ac, 5'd0, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a6, 5'd1, 27'h00000132, 5'd13, 27'h0000021b, 32'h00000400,
  1'd1,  5'd4, 27'h00000051, 5'd4, 27'h0000031e, 5'd23, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000244, 5'd14, 27'h0000011d, 5'd1, 27'h00000379, 32'h00000400,
  1'd1,  5'd1, 27'h00000378, 5'd13, 27'h000001fc, 5'd14, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000017a, 5'd10, 27'h00000373, 5'd25, 27'h000002d0, 32'h00000400,
  1'd1,  5'd1, 27'h00000130, 5'd23, 27'h00000233, 5'd2, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029b, 5'd21, 27'h00000105, 5'd10, 27'h00000342, 32'h00000400,
  1'd1,  5'd1, 27'h000001a6, 5'd25, 27'h0000000b, 5'd24, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000322, 5'd2, 27'h00000066, 5'd4, 27'h000003e0, 32'h00000400,
  1'd1,  5'd12, 27'h000003f1, 5'd4, 27'h00000389, 5'd14, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000038e, 5'd0, 27'h0000024c, 5'd24, 27'h0000008c, 32'h00000400,
  1'd1,  5'd11, 27'h000003ea, 5'd15, 27'h0000019f, 5'd0, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000212, 5'd13, 27'h00000216, 5'd13, 27'h000002c4, 32'h00000400,
  1'd1,  5'd12, 27'h000002e4, 5'd13, 27'h0000030a, 5'd21, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001c2, 5'd25, 27'h000001ae, 5'd1, 27'h00000130, 32'h00000400,
  1'd1,  5'd10, 27'h00000207, 5'd24, 27'h00000017, 5'd11, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000008b, 5'd24, 27'h000002db, 5'd25, 27'h00000151, 32'h00000400,
  1'd1,  5'd20, 27'h00000397, 5'd5, 27'h00000024, 5'd0, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000008, 5'd1, 27'h000003d0, 5'd12, 27'h00000057, 32'h00000400,
  1'd1,  5'd24, 27'h000001a9, 5'd3, 27'h000001f4, 5'd23, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a5, 5'd15, 27'h00000063, 5'd1, 27'h0000023f, 32'h00000400,
  1'd1,  5'd21, 27'h00000088, 5'd14, 27'h00000013, 5'd12, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a5, 5'd14, 27'h00000085, 5'd24, 27'h00000033, 32'h00000400,
  1'd1,  5'd21, 27'h00000297, 5'd22, 27'h000003b5, 5'd2, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000328, 5'd24, 27'h000002a0, 5'd11, 27'h00000264, 32'h00000400,
  1'd1,  5'd24, 27'h000003c5, 5'd23, 27'h0000026f, 5'd25, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000024e, 5'd0, 27'h000003a3, 5'd6, 27'h000000a5, 32'h00000400,
  1'd1,  5'd4, 27'h0000031f, 5'd2, 27'h000000ea, 5'd19, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000213, 5'd1, 27'h000000ae, 5'd26, 27'h0000024f, 32'h00000400,
  1'd1,  5'd2, 27'h00000091, 5'd14, 27'h000002da, 5'd6, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000021, 5'd14, 27'h0000016a, 5'd20, 27'h000000f1, 32'h00000400,
  1'd1,  5'd3, 27'h0000030e, 5'd15, 27'h000000fe, 5'd30, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029d, 5'd20, 27'h00000308, 5'd8, 27'h00000002, 32'h00000400,
  1'd1,  5'd3, 27'h00000252, 5'd23, 27'h00000372, 5'd19, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002f8, 5'd21, 27'h0000028d, 5'd30, 27'h0000029e, 32'h00000400,
  1'd1,  5'd10, 27'h0000035f, 5'd4, 27'h0000011b, 5'd7, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000016, 5'd2, 27'h00000035, 5'd20, 27'h00000170, 32'h00000400,
  1'd1,  5'd13, 27'h000001a7, 5'd0, 27'h000001a5, 5'd29, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c1, 5'd13, 27'h0000028a, 5'd5, 27'h0000035f, 32'h00000400,
  1'd1,  5'd13, 27'h00000004, 5'd13, 27'h000000c1, 5'd15, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000a4, 5'd11, 27'h00000245, 5'd30, 27'h00000391, 32'h00000400,
  1'd1,  5'd14, 27'h00000180, 5'd23, 27'h000001c9, 5'd8, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000141, 5'd23, 27'h00000308, 5'd18, 27'h000003d2, 32'h00000400,
  1'd1,  5'd13, 27'h0000025a, 5'd23, 27'h000002d2, 5'd28, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000068, 5'd1, 27'h0000000d, 5'd7, 27'h000003f6, 32'h00000400,
  1'd1,  5'd23, 27'h0000019c, 5'd3, 27'h0000031f, 5'd17, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000055, 5'd0, 27'h000003e7, 5'd30, 27'h0000038f, 32'h00000400,
  1'd1,  5'd24, 27'h0000002f, 5'd15, 27'h00000004, 5'd8, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000026, 5'd12, 27'h000001de, 5'd19, 27'h00000241, 32'h00000400,
  1'd1,  5'd22, 27'h000002db, 5'd13, 27'h00000368, 5'd28, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000003a, 5'd25, 27'h00000074, 5'd6, 27'h000000a3, 32'h00000400,
  1'd1,  5'd25, 27'h000002d8, 5'd25, 27'h00000293, 5'd17, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000252, 5'd22, 27'h0000003b, 5'd30, 27'h000002d2, 32'h00000400,
  1'd1,  5'd3, 27'h00000220, 5'd9, 27'h00000256, 5'd3, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d1, 5'd8, 27'h000003d9, 5'd14, 27'h00000281, 32'h00000400,
  1'd1,  5'd2, 27'h000002df, 5'd5, 27'h000000f7, 5'd25, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001f2, 5'd19, 27'h00000303, 5'd0, 27'h00000112, 32'h00000400,
  1'd1,  5'd2, 27'h00000148, 5'd16, 27'h00000277, 5'd11, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b8, 5'd20, 27'h0000019a, 5'd24, 27'h00000142, 32'h00000400,
  1'd1,  5'd3, 27'h00000356, 5'd27, 27'h0000033d, 5'd2, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000026a, 5'd30, 27'h000001f7, 5'd11, 27'h0000010f, 32'h00000400,
  1'd1,  5'd1, 27'h00000367, 5'd28, 27'h00000385, 5'd21, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000364, 5'd5, 27'h00000136, 5'd5, 27'h000000a5, 32'h00000400,
  1'd1,  5'd14, 27'h000003e8, 5'd5, 27'h00000164, 5'd12, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000079, 5'd9, 27'h000001bc, 5'd23, 27'h000001a6, 32'h00000400,
  1'd1,  5'd12, 27'h0000013c, 5'd15, 27'h0000022b, 5'd0, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ef, 5'd19, 27'h000001d5, 5'd13, 27'h00000379, 32'h00000400,
  1'd1,  5'd14, 27'h000000ba, 5'd15, 27'h00000276, 5'd24, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000a5, 5'd26, 27'h00000388, 5'd3, 27'h00000080, 32'h00000400,
  1'd1,  5'd10, 27'h0000020a, 5'd27, 27'h0000012d, 5'd13, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003fe, 5'd29, 27'h00000291, 5'd23, 27'h00000393, 32'h00000400,
  1'd1,  5'd23, 27'h000003a3, 5'd9, 27'h00000146, 5'd4, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000299, 5'd6, 27'h0000000c, 5'd14, 27'h000000cc, 32'h00000400,
  1'd1,  5'd25, 27'h00000204, 5'd6, 27'h0000022a, 5'd23, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ef, 5'd15, 27'h00000290, 5'd4, 27'h0000012b, 32'h00000400,
  1'd1,  5'd24, 27'h0000031b, 5'd19, 27'h0000011b, 5'd11, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000141, 5'd18, 27'h0000005f, 5'd24, 27'h000002de, 32'h00000400,
  1'd1,  5'd22, 27'h0000030e, 5'd26, 27'h00000394, 5'd2, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000202, 5'd28, 27'h000001a4, 5'd14, 27'h000003af, 32'h00000400,
  1'd1,  5'd23, 27'h000002bf, 5'd30, 27'h0000032d, 5'd21, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000041, 5'd8, 27'h00000378, 5'd8, 27'h00000252, 32'h00000400,
  1'd1,  5'd2, 27'h00000304, 5'd5, 27'h00000170, 5'd15, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000315, 5'd7, 27'h00000121, 5'd27, 27'h0000022a, 32'h00000400,
  1'd1,  5'd4, 27'h0000017e, 5'd16, 27'h000003cb, 5'd8, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000393, 5'd20, 27'h00000072, 5'd17, 27'h00000079, 32'h00000400,
  1'd1,  5'd3, 27'h000002cb, 5'd19, 27'h000002f0, 5'd30, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000038, 5'd30, 27'h00000114, 5'd9, 27'h00000148, 32'h00000400,
  1'd1,  5'd0, 27'h000002dd, 5'd28, 27'h00000179, 5'd16, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002fa, 5'd29, 27'h000001db, 5'd27, 27'h00000059, 32'h00000400,
  1'd1,  5'd11, 27'h00000126, 5'd7, 27'h000000d3, 5'd10, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f5, 5'd6, 27'h0000010d, 5'd18, 27'h00000197, 32'h00000400,
  1'd1,  5'd10, 27'h0000019e, 5'd9, 27'h0000018d, 5'd27, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000031b, 5'd16, 27'h000002db, 5'd7, 27'h0000007c, 32'h00000400,
  1'd1,  5'd14, 27'h0000036a, 5'd17, 27'h000002a6, 5'd18, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000023c, 5'd19, 27'h0000010a, 5'd30, 27'h000003e0, 32'h00000400,
  1'd1,  5'd13, 27'h00000205, 5'd28, 27'h0000015b, 5'd7, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029c, 5'd28, 27'h00000071, 5'd15, 27'h000002b1, 32'h00000400,
  1'd1,  5'd14, 27'h00000111, 5'd27, 27'h000000ee, 5'd28, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d3, 5'd9, 27'h00000266, 5'd7, 27'h00000014, 32'h00000400,
  1'd1,  5'd23, 27'h00000243, 5'd10, 27'h0000007c, 5'd18, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000385, 5'd8, 27'h000001d7, 5'd30, 27'h00000039, 32'h00000400,
  1'd1,  5'd24, 27'h000001e8, 5'd16, 27'h0000024e, 5'd7, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000370, 5'd16, 27'h00000187, 5'd17, 27'h00000027, 32'h00000400,
  1'd1,  5'd25, 27'h0000004c, 5'd20, 27'h0000001e, 5'd26, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000179, 5'd30, 27'h000002ee, 5'd7, 27'h00000094, 32'h00000400,
  1'd1,  5'd25, 27'h000001ec, 5'd28, 27'h00000025, 5'd19, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000128, 5'd29, 27'h0000039c, 5'd27, 27'h000002d1, 32'h00000400,
  1'd1,  5'd6, 27'h000000bb, 5'd2, 27'h00000312, 5'd7, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a5, 5'd3, 27'h00000011, 5'd16, 27'h00000084, 32'h00000400,
  1'd1,  5'd6, 27'h0000005c, 5'd4, 27'h00000273, 5'd25, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a9, 5'd15, 27'h000001aa, 5'd2, 27'h0000024c, 32'h00000400,
  1'd1,  5'd6, 27'h000003ea, 5'd10, 27'h00000246, 5'd11, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000027f, 5'd11, 27'h000000cb, 5'd24, 27'h00000062, 32'h00000400,
  1'd1,  5'd8, 27'h00000234, 5'd23, 27'h00000255, 5'd4, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000124, 5'd23, 27'h00000041, 5'd13, 27'h00000168, 32'h00000400,
  1'd1,  5'd6, 27'h0000039c, 5'd25, 27'h000000b5, 5'd22, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d2, 5'd4, 27'h0000039f, 5'd5, 27'h00000271, 32'h00000400,
  1'd1,  5'd20, 27'h000000e4, 5'd3, 27'h00000279, 5'd20, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000039c, 5'd0, 27'h0000019d, 5'd29, 27'h00000095, 32'h00000400,
  1'd1,  5'd19, 27'h000002fa, 5'd12, 27'h000002c3, 5'd4, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000b7, 5'd13, 27'h0000015a, 5'd13, 27'h00000085, 32'h00000400,
  1'd1,  5'd17, 27'h000000e0, 5'd11, 27'h000001cc, 5'd23, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ec, 5'd22, 27'h00000064, 5'd3, 27'h00000296, 32'h00000400,
  1'd1,  5'd20, 27'h000001ae, 5'd20, 27'h000002d1, 5'd15, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000393, 5'd23, 27'h0000037f, 5'd21, 27'h0000027b, 32'h00000400,
  1'd1,  5'd30, 27'h00000122, 5'd1, 27'h0000030b, 5'd1, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000267, 5'd3, 27'h00000169, 5'd12, 27'h000000a7, 32'h00000400,
  1'd1,  5'd28, 27'h000003f5, 5'd1, 27'h000001d0, 5'd23, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000062, 5'd15, 27'h0000015e, 5'd0, 27'h0000020f, 32'h00000400,
  1'd1,  5'd28, 27'h0000022a, 5'd14, 27'h00000187, 5'd14, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000024b, 5'd15, 27'h000001f7, 5'd24, 27'h00000349, 32'h00000400,
  1'd1,  5'd26, 27'h000000d7, 5'd21, 27'h000003a2, 5'd2, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a4, 5'd20, 27'h00000340, 5'd12, 27'h000002d4, 32'h00000400,
  1'd1,  5'd27, 27'h00000085, 5'd22, 27'h00000241, 5'd21, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000138, 5'd4, 27'h00000252, 5'd3, 27'h000002ca, 32'h00000400,
  1'd1,  5'd7, 27'h00000149, 5'd4, 27'h0000003e, 5'd12, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000011, 5'd3, 27'h00000325, 5'd21, 27'h00000004, 32'h00000400,
  1'd1,  5'd6, 27'h000003ae, 5'd12, 27'h0000032a, 5'd9, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ca, 5'd10, 27'h000002a4, 5'd20, 27'h000001ef, 32'h00000400,
  1'd1,  5'd6, 27'h00000121, 5'd13, 27'h00000002, 5'd26, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fe, 5'd24, 27'h000000a4, 5'd8, 27'h0000027c, 32'h00000400,
  1'd1,  5'd6, 27'h000002f9, 5'd22, 27'h000003c0, 5'd16, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000317, 5'd23, 27'h00000239, 5'd29, 27'h00000125, 32'h00000400,
  1'd1,  5'd18, 27'h00000190, 5'd2, 27'h0000005d, 5'd1, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000147, 5'd1, 27'h000001b4, 5'd15, 27'h0000008b, 32'h00000400,
  1'd1,  5'd16, 27'h0000014e, 5'd3, 27'h000000cb, 5'd25, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000365, 5'd10, 27'h00000398, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd16, 27'h0000039b, 5'd10, 27'h00000304, 5'd16, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039f, 5'd11, 27'h000003b7, 5'd26, 27'h0000015d, 32'h00000400,
  1'd1,  5'd20, 27'h00000022, 5'd20, 27'h000002db, 5'd7, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001d9, 5'd25, 27'h00000332, 5'd16, 27'h0000008c, 32'h00000400,
  1'd1,  5'd18, 27'h000000f1, 5'd25, 27'h00000166, 5'd26, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000211, 5'd1, 27'h000003e7, 5'd8, 27'h00000382, 32'h00000400,
  1'd1,  5'd26, 27'h0000031f, 5'd2, 27'h0000033d, 5'd16, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b0, 5'd1, 27'h0000002c, 5'd28, 27'h00000124, 32'h00000400,
  1'd1,  5'd26, 27'h000002c4, 5'd15, 27'h00000016, 5'd9, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000301, 5'd15, 27'h000001e9, 5'd19, 27'h000003f4, 32'h00000400,
  1'd1,  5'd26, 27'h000001d7, 5'd12, 27'h00000129, 5'd29, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000141, 5'd24, 27'h0000013c, 5'd8, 27'h0000037e, 32'h00000400,
  1'd1,  5'd26, 27'h00000113, 5'd22, 27'h00000148, 5'd18, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007d, 5'd23, 27'h0000037a, 5'd28, 27'h0000034c, 32'h00000400,
  1'd1,  5'd9, 27'h00000341, 5'd6, 27'h0000001f, 5'd2, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003d9, 5'd7, 27'h00000085, 5'd13, 27'h000003ce, 32'h00000400,
  1'd1,  5'd6, 27'h00000006, 5'd9, 27'h00000037, 5'd21, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a9, 5'd20, 27'h0000023c, 5'd3, 27'h000000ce, 32'h00000400,
  1'd1,  5'd5, 27'h00000305, 5'd16, 27'h00000023, 5'd15, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000016e, 5'd15, 27'h000003f2, 5'd23, 27'h00000220, 32'h00000400,
  1'd1,  5'd5, 27'h0000029d, 5'd30, 27'h000003d7, 5'd4, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000278, 5'd27, 27'h000002d3, 5'd14, 27'h0000025a, 32'h00000400,
  1'd1,  5'd7, 27'h0000030f, 5'd30, 27'h000003ed, 5'd23, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d7, 5'd5, 27'h000002d9, 5'd4, 27'h000000bd, 32'h00000400,
  1'd1,  5'd17, 27'h00000132, 5'd5, 27'h000000bb, 5'd14, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ce, 5'd5, 27'h000002e0, 5'd21, 27'h0000031e, 32'h00000400,
  1'd1,  5'd16, 27'h00000125, 5'd20, 27'h00000008, 5'd4, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000132, 5'd16, 27'h00000210, 5'd12, 27'h0000011a, 32'h00000400,
  1'd1,  5'd18, 27'h000003e2, 5'd18, 27'h00000238, 5'd23, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000018b, 5'd27, 27'h00000343, 5'd0, 27'h00000220, 32'h00000400,
  1'd1,  5'd16, 27'h000003a9, 5'd29, 27'h000000a2, 5'd13, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001b1, 5'd26, 27'h0000011e, 5'd24, 27'h000002d3, 32'h00000400,
  1'd1,  5'd26, 27'h0000031d, 5'd6, 27'h00000215, 5'd2, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001bb, 5'd8, 27'h000001f5, 5'd15, 27'h0000014b, 32'h00000400,
  1'd1,  5'd30, 27'h000002cb, 5'd7, 27'h000002a5, 5'd22, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002bd, 5'd19, 27'h0000011b, 5'd1, 27'h0000008c, 32'h00000400,
  1'd1,  5'd29, 27'h0000034c, 5'd16, 27'h00000351, 5'd14, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003cb, 5'd16, 27'h0000019c, 5'd25, 27'h0000022a, 32'h00000400,
  1'd1,  5'd27, 27'h000003af, 5'd30, 27'h00000302, 5'd3, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000347, 5'd30, 27'h000001ab, 5'd14, 27'h000000a6, 32'h00000400,
  1'd1,  5'd29, 27'h00000090, 5'd28, 27'h00000046, 5'd24, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000007, 5'd6, 27'h0000014e, 5'd9, 27'h00000043, 32'h00000400,
  1'd1,  5'd9, 27'h00000190, 5'd8, 27'h00000165, 5'd15, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e3, 5'd7, 27'h000000c8, 5'd30, 27'h000002d8, 32'h00000400,
  1'd1,  5'd9, 27'h00000051, 5'd16, 27'h000002e9, 5'd9, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000030, 5'd16, 27'h0000015c, 5'd16, 27'h00000080, 32'h00000400,
  1'd1,  5'd7, 27'h000001d5, 5'd15, 27'h00000342, 5'd26, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000269, 5'd30, 27'h000001b6, 5'd7, 27'h000002ce, 32'h00000400,
  1'd1,  5'd10, 27'h00000051, 5'd27, 27'h000003de, 5'd16, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e7, 5'd30, 27'h00000211, 5'd28, 27'h000001c0, 32'h00000400,
  1'd1,  5'd17, 27'h00000009, 5'd5, 27'h0000023a, 5'd5, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000025a, 5'd8, 27'h00000004, 5'd17, 27'h000000b6, 32'h00000400,
  1'd1,  5'd20, 27'h0000020a, 5'd6, 27'h000000fe, 5'd30, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000033, 5'd18, 27'h0000009a, 5'd6, 27'h00000338, 32'h00000400,
  1'd1,  5'd16, 27'h00000395, 5'd20, 27'h000000ef, 5'd15, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000039, 5'd19, 27'h000003af, 5'd29, 27'h0000000c, 32'h00000400,
  1'd1,  5'd15, 27'h00000329, 5'd29, 27'h000001ee, 5'd8, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a0, 5'd29, 27'h00000058, 5'd19, 27'h00000272, 32'h00000400,
  1'd1,  5'd18, 27'h0000020d, 5'd26, 27'h00000246, 5'd26, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000129, 5'd8, 27'h000000b4, 5'd6, 27'h00000319, 32'h00000400,
  1'd1,  5'd27, 27'h000002a5, 5'd6, 27'h000000ba, 5'd19, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000374, 5'd7, 27'h000003e9, 5'd27, 27'h000001ad, 32'h00000400,
  1'd1,  5'd29, 27'h000003b8, 5'd16, 27'h00000109, 5'd8, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000197, 5'd20, 27'h0000004c, 5'd20, 27'h00000039, 32'h00000400,
  1'd1,  5'd30, 27'h000000ec, 5'd18, 27'h0000016b, 5'd29, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000031a, 5'd26, 27'h000001c9, 5'd9, 27'h0000035b, 32'h00000400,
  1'd1,  5'd29, 27'h00000365, 5'd30, 27'h0000024b, 5'd18, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000336, 5'd27, 27'h0000017c, 5'd26, 27'h0000038b, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001a4, 5'd0, 27'h000001fb, 5'd1, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ab, 5'd3, 27'h000003e9, 5'd10, 27'h0000016c, 32'h00000400,
  1'd1,  5'd0, 27'h00000055, 5'd3, 27'h00000073, 5'd23, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d5, 5'd14, 27'h0000013f, 5'd2, 27'h00000041, 32'h00000400,
  1'd1,  5'd0, 27'h000002fe, 5'd14, 27'h00000241, 5'd13, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000059, 5'd12, 27'h0000015d, 5'd24, 27'h000001b7, 32'h00000400,
  1'd1,  5'd1, 27'h00000328, 5'd24, 27'h00000010, 5'd5, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d7, 5'd21, 27'h00000273, 5'd13, 27'h00000030, 32'h00000400,
  1'd1,  5'd0, 27'h00000248, 5'd20, 27'h000002c9, 5'd21, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035d, 5'd1, 27'h000000cf, 5'd1, 27'h00000190, 32'h00000400,
  1'd1,  5'd12, 27'h0000024f, 5'd2, 27'h000002b7, 5'd10, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001fb, 5'd1, 27'h0000025f, 5'd22, 27'h00000010, 32'h00000400,
  1'd1,  5'd13, 27'h000002da, 5'd14, 27'h00000225, 5'd1, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ad, 5'd12, 27'h000000ad, 5'd12, 27'h00000146, 32'h00000400,
  1'd1,  5'd12, 27'h00000208, 5'd10, 27'h0000029f, 5'd25, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000033a, 5'd22, 27'h00000136, 5'd2, 27'h000001b1, 32'h00000400,
  1'd1,  5'd12, 27'h00000316, 5'd23, 27'h000001f8, 5'd13, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000371, 5'd25, 27'h00000036, 5'd23, 27'h00000187, 32'h00000400,
  1'd1,  5'd22, 27'h00000237, 5'd4, 27'h0000023a, 5'd2, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000011b, 5'd4, 27'h000002e0, 5'd13, 27'h00000383, 32'h00000400,
  1'd1,  5'd25, 27'h00000049, 5'd5, 27'h0000009b, 5'd25, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000028e, 5'd12, 27'h000003bf, 5'd2, 27'h00000146, 32'h00000400,
  1'd1,  5'd24, 27'h0000012c, 5'd11, 27'h000003ec, 5'd12, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000150, 5'd11, 27'h0000001e, 5'd24, 27'h00000399, 32'h00000400,
  1'd1,  5'd21, 27'h00000280, 5'd25, 27'h00000047, 5'd3, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e3, 5'd23, 27'h00000393, 5'd14, 27'h0000000c, 32'h00000400,
  1'd1,  5'd24, 27'h0000009e, 5'd25, 27'h000000e2, 5'd21, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000308, 5'd4, 27'h0000030e, 5'd9, 27'h000000c0, 32'h00000400,
  1'd1,  5'd0, 27'h00000359, 5'd1, 27'h00000003, 5'd16, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003f0, 5'd2, 27'h000003e1, 5'd26, 27'h0000005b, 32'h00000400,
  1'd1,  5'd4, 27'h00000329, 5'd12, 27'h000003db, 5'd7, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b2, 5'd13, 27'h00000377, 5'd19, 27'h00000106, 32'h00000400,
  1'd1,  5'd4, 27'h000001a5, 5'd11, 27'h000001c0, 5'd28, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000027, 5'd22, 27'h00000203, 5'd7, 27'h00000377, 32'h00000400,
  1'd1,  5'd1, 27'h00000277, 5'd23, 27'h0000006d, 5'd15, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000006e, 5'd22, 27'h00000024, 5'd30, 27'h000001a4, 32'h00000400,
  1'd1,  5'd11, 27'h000000f4, 5'd3, 27'h00000383, 5'd9, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ce, 5'd2, 27'h000003ad, 5'd18, 27'h00000362, 32'h00000400,
  1'd1,  5'd14, 27'h0000006f, 5'd3, 27'h0000012d, 5'd28, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000002f, 5'd14, 27'h000002e0, 5'd8, 27'h000003ed, 32'h00000400,
  1'd1,  5'd10, 27'h000001ed, 5'd14, 27'h000003a5, 5'd18, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000036b, 5'd11, 27'h00000131, 5'd28, 27'h000001a1, 32'h00000400,
  1'd1,  5'd12, 27'h00000106, 5'd21, 27'h00000124, 5'd7, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000206, 5'd25, 27'h0000002f, 5'd18, 27'h00000110, 32'h00000400,
  1'd1,  5'd13, 27'h00000328, 5'd24, 27'h00000210, 5'd29, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000270, 5'd3, 27'h000000d7, 5'd10, 27'h00000075, 32'h00000400,
  1'd1,  5'd21, 27'h0000001b, 5'd3, 27'h0000021f, 5'd16, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003ba, 5'd1, 27'h0000021d, 5'd28, 27'h000001ae, 32'h00000400,
  1'd1,  5'd21, 27'h00000092, 5'd12, 27'h000000c0, 5'd6, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000326, 5'd11, 27'h000000ba, 5'd19, 27'h00000057, 32'h00000400,
  1'd1,  5'd20, 27'h000003d5, 5'd13, 27'h00000318, 5'd25, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000007b, 5'd22, 27'h00000059, 5'd5, 27'h000001f3, 32'h00000400,
  1'd1,  5'd25, 27'h00000096, 5'd20, 27'h00000300, 5'd17, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000023b, 5'd24, 27'h000001a9, 5'd29, 27'h00000124, 32'h00000400,
  1'd1,  5'd0, 27'h0000033d, 5'd10, 27'h0000014b, 5'd5, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000027b, 5'd9, 27'h0000039b, 5'd14, 27'h00000010, 32'h00000400,
  1'd1,  5'd1, 27'h0000017e, 5'd7, 27'h00000079, 5'd22, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002b, 5'd16, 27'h000001b7, 5'd2, 27'h00000115, 32'h00000400,
  1'd1,  5'd0, 27'h00000399, 5'd17, 27'h0000034c, 5'd13, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000016c, 5'd15, 27'h00000281, 5'd22, 27'h000002a0, 32'h00000400,
  1'd1,  5'd1, 27'h0000035f, 5'd26, 27'h00000020, 5'd3, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000297, 5'd27, 27'h00000033, 5'd12, 27'h0000009c, 32'h00000400,
  1'd1,  5'd4, 27'h0000022d, 5'd26, 27'h00000290, 5'd24, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000030, 5'd8, 27'h00000342, 5'd0, 27'h000001b1, 32'h00000400,
  1'd1,  5'd13, 27'h0000007c, 5'd6, 27'h00000313, 5'd14, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003bb, 5'd8, 27'h0000016f, 5'd22, 27'h0000031b, 32'h00000400,
  1'd1,  5'd12, 27'h0000019e, 5'd19, 27'h0000024d, 5'd0, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000000b, 5'd16, 27'h00000093, 5'd13, 27'h000001ee, 32'h00000400,
  1'd1,  5'd13, 27'h0000026a, 5'd19, 27'h00000279, 5'd21, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000012e, 5'd25, 27'h000003af, 5'd2, 27'h0000002e, 32'h00000400,
  1'd1,  5'd13, 27'h0000037e, 5'd30, 27'h0000027f, 5'd11, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000060, 5'd28, 27'h000000a8, 5'd24, 27'h00000270, 32'h00000400,
  1'd1,  5'd20, 27'h000003ff, 5'd10, 27'h000000c6, 5'd4, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000346, 5'd5, 27'h00000300, 5'd13, 27'h000001f3, 32'h00000400,
  1'd1,  5'd23, 27'h00000127, 5'd7, 27'h000002f7, 5'd22, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032d, 5'd18, 27'h00000143, 5'd1, 27'h000002a6, 32'h00000400,
  1'd1,  5'd21, 27'h00000357, 5'd18, 27'h000002e9, 5'd12, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000021b, 5'd19, 27'h0000034e, 5'd24, 27'h00000193, 32'h00000400,
  1'd1,  5'd25, 27'h00000329, 5'd29, 27'h0000017f, 5'd3, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000037d, 5'd30, 27'h000001c2, 5'd13, 27'h00000040, 32'h00000400,
  1'd1,  5'd20, 27'h000002e5, 5'd28, 27'h000002af, 5'd22, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003cc, 5'd9, 27'h000001c9, 5'd7, 27'h00000075, 32'h00000400,
  1'd1,  5'd0, 27'h000002ba, 5'd7, 27'h000003f6, 5'd19, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ba, 5'd7, 27'h0000015e, 5'd27, 27'h000000e4, 32'h00000400,
  1'd1,  5'd1, 27'h00000135, 5'd19, 27'h0000028a, 5'd6, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001b2, 5'd18, 27'h000001e5, 5'd16, 27'h00000360, 32'h00000400,
  1'd1,  5'd4, 27'h000003db, 5'd19, 27'h00000015, 5'd26, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f7, 5'd30, 27'h000003cd, 5'd10, 27'h000000f4, 32'h00000400,
  1'd1,  5'd3, 27'h000002c1, 5'd26, 27'h00000130, 5'd17, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002ca, 5'd26, 27'h0000036d, 5'd29, 27'h00000288, 32'h00000400,
  1'd1,  5'd10, 27'h0000037c, 5'd5, 27'h0000019f, 5'd9, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000306, 5'd6, 27'h000001b3, 5'd18, 27'h000003b5, 32'h00000400,
  1'd1,  5'd13, 27'h00000208, 5'd8, 27'h00000029, 5'd28, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000152, 5'd17, 27'h0000025c, 5'd9, 27'h0000025d, 32'h00000400,
  1'd1,  5'd11, 27'h0000004c, 5'd20, 27'h00000190, 5'd16, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000301, 5'd18, 27'h00000226, 5'd26, 27'h000001a2, 32'h00000400,
  1'd1,  5'd14, 27'h000001c1, 5'd28, 27'h0000036b, 5'd9, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a0, 5'd28, 27'h00000077, 5'd19, 27'h000001ce, 32'h00000400,
  1'd1,  5'd12, 27'h000000cf, 5'd30, 27'h000000e9, 5'd29, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001cb, 5'd7, 27'h00000318, 5'd5, 27'h0000015b, 32'h00000400,
  1'd1,  5'd21, 27'h000000b1, 5'd8, 27'h00000218, 5'd20, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000192, 5'd6, 27'h000003a8, 5'd29, 27'h0000007a, 32'h00000400,
  1'd1,  5'd20, 27'h000002c9, 5'd20, 27'h00000099, 5'd8, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001cf, 5'd20, 27'h00000145, 5'd17, 27'h00000012, 32'h00000400,
  1'd1,  5'd22, 27'h000000a5, 5'd20, 27'h000001f3, 5'd28, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000162, 5'd30, 27'h000001e5, 5'd8, 27'h00000158, 32'h00000400,
  1'd1,  5'd21, 27'h00000168, 5'd28, 27'h00000231, 5'd20, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002c6, 5'd26, 27'h000003e8, 5'd30, 27'h000000f2, 32'h00000400,
  1'd1,  5'd6, 27'h00000399, 5'd4, 27'h0000018d, 5'd6, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032a, 5'd3, 27'h000001fa, 5'd20, 27'h000001fd, 32'h00000400,
  1'd1,  5'd6, 27'h00000216, 5'd3, 27'h000003d9, 5'd30, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000029d, 5'd12, 27'h000000e0, 5'd0, 27'h000002ff, 32'h00000400,
  1'd1,  5'd7, 27'h0000023f, 5'd13, 27'h000002fc, 5'd14, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000025d, 5'd13, 27'h000000ea, 5'd20, 27'h00000335, 32'h00000400,
  1'd1,  5'd7, 27'h0000027f, 5'd23, 27'h000001ca, 5'd0, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001be, 5'd24, 27'h00000056, 5'd13, 27'h000003f1, 32'h00000400,
  1'd1,  5'd5, 27'h00000266, 5'd22, 27'h000002ee, 5'd25, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000044, 5'd1, 27'h000003e7, 5'd8, 27'h00000250, 32'h00000400,
  1'd1,  5'd18, 27'h000003a4, 5'd2, 27'h00000387, 5'd18, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000129, 5'd0, 27'h00000235, 5'd27, 27'h000003ba, 32'h00000400,
  1'd1,  5'd18, 27'h000000e2, 5'd13, 27'h00000368, 5'd3, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000284, 5'd14, 27'h0000005f, 5'd11, 27'h000002e1, 32'h00000400,
  1'd1,  5'd17, 27'h000000a3, 5'd13, 27'h000003c1, 5'd20, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000072, 5'd25, 27'h00000178, 5'd4, 27'h00000315, 32'h00000400,
  1'd1,  5'd16, 27'h0000004c, 5'd23, 27'h000003bc, 5'd12, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000291, 5'd24, 27'h0000034a, 5'd21, 27'h000001f2, 32'h00000400,
  1'd1,  5'd27, 27'h00000369, 5'd4, 27'h000001b9, 5'd3, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002d9, 5'd0, 27'h000000a9, 5'd11, 27'h00000193, 32'h00000400,
  1'd1,  5'd27, 27'h00000171, 5'd0, 27'h0000012e, 5'd23, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002fd, 5'd10, 27'h000001e0, 5'd0, 27'h000000ac, 32'h00000400,
  1'd1,  5'd29, 27'h00000070, 5'd12, 27'h0000003b, 5'd12, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000200, 5'd10, 27'h00000351, 5'd22, 27'h0000023d, 32'h00000400,
  1'd1,  5'd25, 27'h00000399, 5'd24, 27'h00000302, 5'd1, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000209, 5'd23, 27'h000002a2, 5'd13, 27'h00000075, 32'h00000400,
  1'd1,  5'd26, 27'h0000003a, 5'd23, 27'h00000282, 5'd23, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000fa, 5'd0, 27'h000002c7, 5'd2, 27'h00000288, 32'h00000400,
  1'd1,  5'd7, 27'h00000301, 5'd0, 27'h0000027c, 5'd13, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e4, 5'd5, 27'h00000011, 5'd21, 27'h00000223, 32'h00000400,
  1'd1,  5'd6, 27'h00000223, 5'd14, 27'h00000367, 5'd5, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000076, 5'd15, 27'h00000193, 5'd16, 27'h00000253, 32'h00000400,
  1'd1,  5'd8, 27'h000001ed, 5'd11, 27'h000001fd, 5'd27, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000343, 5'd25, 27'h000000dc, 5'd5, 27'h000002e9, 32'h00000400,
  1'd1,  5'd7, 27'h000000b0, 5'd22, 27'h00000261, 5'd18, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003f5, 5'd22, 27'h00000068, 5'd29, 27'h00000189, 32'h00000400,
  1'd1,  5'd15, 27'h000002cb, 5'd2, 27'h000002e1, 5'd2, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002df, 5'd3, 27'h00000151, 5'd14, 27'h0000007c, 32'h00000400,
  1'd1,  5'd19, 27'h0000027d, 5'd0, 27'h00000191, 5'd21, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016c, 5'd12, 27'h000003b5, 5'd8, 27'h000002f8, 32'h00000400,
  1'd1,  5'd18, 27'h000003c1, 5'd13, 27'h000003e7, 5'd16, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a1, 5'd14, 27'h000001ab, 5'd29, 27'h000002e8, 32'h00000400,
  1'd1,  5'd20, 27'h0000010a, 5'd23, 27'h00000377, 5'd7, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000377, 5'd22, 27'h000002cf, 5'd17, 27'h00000372, 32'h00000400,
  1'd1,  5'd18, 27'h0000008a, 5'd23, 27'h0000010d, 5'd28, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003a7, 5'd0, 27'h00000204, 5'd7, 27'h000003c4, 32'h00000400,
  1'd1,  5'd26, 27'h000000e2, 5'd4, 27'h0000027d, 5'd16, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000020, 5'd2, 27'h00000226, 5'd30, 27'h0000010e, 32'h00000400,
  1'd1,  5'd27, 27'h0000036c, 5'd12, 27'h000000f6, 5'd6, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000125, 5'd13, 27'h000000d3, 5'd20, 27'h000001b0, 32'h00000400,
  1'd1,  5'd26, 27'h000002c2, 5'd10, 27'h00000284, 5'd28, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000240, 5'd23, 27'h000002de, 5'd6, 27'h0000039f, 32'h00000400,
  1'd1,  5'd29, 27'h000002fb, 5'd22, 27'h000000e9, 5'd18, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ec, 5'd24, 27'h00000200, 5'd26, 27'h000000b0, 32'h00000400,
  1'd1,  5'd7, 27'h000002d7, 5'd5, 27'h0000028f, 5'd1, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b4, 5'd6, 27'h00000382, 5'd12, 27'h0000005e, 32'h00000400,
  1'd1,  5'd5, 27'h000001bc, 5'd6, 27'h000002b6, 5'd23, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f1, 5'd17, 27'h000002df, 5'd1, 27'h00000240, 32'h00000400,
  1'd1,  5'd10, 27'h00000089, 5'd17, 27'h000001b5, 5'd10, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000bb, 5'd20, 27'h000001d0, 5'd25, 27'h00000019, 32'h00000400,
  1'd1,  5'd9, 27'h00000195, 5'd30, 27'h000002f0, 5'd2, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b0, 5'd27, 27'h00000135, 5'd10, 27'h000003fe, 32'h00000400,
  1'd1,  5'd6, 27'h000003da, 5'd29, 27'h000003f9, 5'd25, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000011, 5'd6, 27'h00000147, 5'd0, 27'h000001a6, 32'h00000400,
  1'd1,  5'd18, 27'h0000004c, 5'd10, 27'h000000c5, 5'd10, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000042, 5'd6, 27'h000001fc, 5'd22, 27'h000003b0, 32'h00000400,
  1'd1,  5'd20, 27'h00000041, 5'd17, 27'h00000313, 5'd2, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000364, 5'd16, 27'h000003d1, 5'd10, 27'h0000023e, 32'h00000400,
  1'd1,  5'd19, 27'h000002e8, 5'd17, 27'h000000f7, 5'd23, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003bb, 5'd29, 27'h00000388, 5'd0, 27'h00000189, 32'h00000400,
  1'd1,  5'd18, 27'h000000ac, 5'd26, 27'h0000019e, 5'd13, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000036, 5'd30, 27'h00000292, 5'd22, 27'h00000372, 32'h00000400,
  1'd1,  5'd28, 27'h00000374, 5'd6, 27'h0000016b, 5'd4, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000017f, 5'd7, 27'h00000307, 5'd13, 27'h000001e6, 32'h00000400,
  1'd1,  5'd30, 27'h00000240, 5'd7, 27'h0000016c, 5'd24, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000238, 5'd19, 27'h00000379, 5'd1, 27'h000002bb, 32'h00000400,
  1'd1,  5'd26, 27'h00000036, 5'd18, 27'h0000013d, 5'd11, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000206, 5'd20, 27'h00000127, 5'd22, 27'h00000132, 32'h00000400,
  1'd1,  5'd29, 27'h00000045, 5'd26, 27'h0000036a, 5'd0, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ed, 5'd26, 27'h000000ac, 5'd14, 27'h00000086, 32'h00000400,
  1'd1,  5'd30, 27'h00000088, 5'd28, 27'h00000111, 5'd24, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000394, 5'd6, 27'h00000251, 5'd5, 27'h000003b3, 32'h00000400,
  1'd1,  5'd6, 27'h00000036, 5'd5, 27'h00000208, 5'd16, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000201, 5'd6, 27'h000000af, 5'd30, 27'h0000031a, 32'h00000400,
  1'd1,  5'd7, 27'h0000021d, 5'd19, 27'h00000298, 5'd9, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b9, 5'd17, 27'h00000187, 5'd19, 27'h00000288, 32'h00000400,
  1'd1,  5'd9, 27'h000002b2, 5'd20, 27'h00000040, 5'd26, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000036a, 5'd26, 27'h00000332, 5'd8, 27'h000000fc, 32'h00000400,
  1'd1,  5'd10, 27'h00000072, 5'd30, 27'h0000007c, 5'd16, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000067, 5'd26, 27'h00000294, 5'd26, 27'h00000130, 32'h00000400,
  1'd1,  5'd18, 27'h000002fb, 5'd10, 27'h00000101, 5'd10, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000302, 5'd9, 27'h00000129, 5'd19, 27'h00000053, 32'h00000400,
  1'd1,  5'd20, 27'h0000026d, 5'd9, 27'h00000062, 5'd28, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000272, 5'd18, 27'h00000316, 5'd9, 27'h0000034b, 32'h00000400,
  1'd1,  5'd16, 27'h000002dd, 5'd18, 27'h00000213, 5'd17, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ef, 5'd17, 27'h0000007e, 5'd27, 27'h000002d6, 32'h00000400,
  1'd1,  5'd19, 27'h00000257, 5'd30, 27'h00000379, 5'd9, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000030f, 5'd26, 27'h000003be, 5'd16, 27'h0000034d, 32'h00000400,
  1'd1,  5'd17, 27'h000000f2, 5'd26, 27'h0000038c, 5'd26, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000036, 5'd9, 27'h000003f3, 5'd9, 27'h000001d0, 32'h00000400,
  1'd1,  5'd28, 27'h00000228, 5'd6, 27'h0000018a, 5'd20, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ce, 5'd7, 27'h00000368, 5'd28, 27'h000003e7, 32'h00000400,
  1'd1,  5'd28, 27'h0000014b, 5'd20, 27'h0000009f, 5'd8, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000198, 5'd19, 27'h00000175, 5'd19, 27'h000000e9, 32'h00000400,
  1'd1,  5'd29, 27'h0000035a, 5'd16, 27'h0000022b, 5'd27, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000190, 5'd26, 27'h0000024b, 5'd9, 27'h00000337, 32'h00000400,
  1'd1,  5'd29, 27'h000003ad, 5'd28, 27'h00000266, 5'd16, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003d3, 5'd28, 27'h000002f4, 5'd27, 27'h00000392, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000000a4, 5'd1, 27'h00000301, 5'd4, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000223, 5'd2, 27'h000002bd, 5'd11, 27'h00000106, 32'h00000400,
  1'd1,  5'd2, 27'h000001d7, 5'd4, 27'h000002e5, 5'd21, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000375, 5'd11, 27'h000001ec, 5'd1, 27'h000001d8, 32'h00000400,
  1'd1,  5'd5, 27'h0000008b, 5'd11, 27'h0000011e, 5'd12, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000011f, 5'd11, 27'h00000262, 5'd24, 27'h00000031, 32'h00000400,
  1'd1,  5'd3, 27'h000001cd, 5'd23, 27'h0000000e, 5'd2, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000006e, 5'd24, 27'h000002d8, 5'd14, 27'h000002a2, 32'h00000400,
  1'd1,  5'd3, 27'h00000136, 5'd25, 27'h000002d9, 5'd21, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000cd, 5'd4, 27'h0000033d, 5'd1, 27'h00000162, 32'h00000400,
  1'd1,  5'd12, 27'h00000151, 5'd1, 27'h00000200, 5'd11, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ee, 5'd3, 27'h0000019f, 5'd21, 27'h000001ea, 32'h00000400,
  1'd1,  5'd10, 27'h00000389, 5'd10, 27'h00000197, 5'd0, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000189, 5'd11, 27'h00000106, 5'd11, 27'h000001a9, 32'h00000400,
  1'd1,  5'd13, 27'h0000012a, 5'd10, 27'h0000022d, 5'd23, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001f4, 5'd23, 27'h0000018f, 5'd2, 27'h000000f0, 32'h00000400,
  1'd1,  5'd12, 27'h000001d1, 5'd24, 27'h000002e8, 5'd14, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000191, 5'd21, 27'h000003c4, 5'd22, 27'h00000014, 32'h00000400,
  1'd1,  5'd24, 27'h00000077, 5'd2, 27'h00000006, 5'd2, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000128, 5'd4, 27'h000000f5, 5'd11, 27'h00000017, 32'h00000400,
  1'd1,  5'd21, 27'h0000023c, 5'd5, 27'h0000008f, 5'd23, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000340, 5'd10, 27'h00000165, 5'd2, 27'h0000003f, 32'h00000400,
  1'd1,  5'd20, 27'h000003ed, 5'd13, 27'h00000191, 5'd14, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000033f, 5'd11, 27'h00000105, 5'd24, 27'h00000321, 32'h00000400,
  1'd1,  5'd23, 27'h0000020c, 5'd23, 27'h000002d3, 5'd0, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038b, 5'd25, 27'h00000211, 5'd10, 27'h00000372, 32'h00000400,
  1'd1,  5'd21, 27'h000000a5, 5'd23, 27'h000003b7, 5'd23, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000016a, 5'd2, 27'h000003c6, 5'd9, 27'h0000004f, 32'h00000400,
  1'd1,  5'd1, 27'h000001ea, 5'd3, 27'h00000005, 5'd20, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d5, 5'd3, 27'h00000361, 5'd26, 27'h000003c1, 32'h00000400,
  1'd1,  5'd4, 27'h0000014e, 5'd10, 27'h000003ca, 5'd5, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000254, 5'd14, 27'h00000121, 5'd17, 27'h00000009, 32'h00000400,
  1'd1,  5'd1, 27'h000000f4, 5'd12, 27'h00000236, 5'd30, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c0, 5'd23, 27'h0000010f, 5'd9, 27'h000001e1, 32'h00000400,
  1'd1,  5'd2, 27'h00000159, 5'd21, 27'h000003b6, 5'd20, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003dd, 5'd24, 27'h00000319, 5'd30, 27'h0000002d, 32'h00000400,
  1'd1,  5'd12, 27'h0000024a, 5'd2, 27'h000002d1, 5'd8, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000184, 5'd2, 27'h000003fa, 5'd20, 27'h0000004c, 32'h00000400,
  1'd1,  5'd11, 27'h0000024b, 5'd0, 27'h00000030, 5'd27, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c2, 5'd12, 27'h000003ea, 5'd6, 27'h000003a5, 32'h00000400,
  1'd1,  5'd12, 27'h0000023e, 5'd11, 27'h000001a6, 5'd17, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000317, 5'd13, 27'h0000027e, 5'd29, 27'h000002b1, 32'h00000400,
  1'd1,  5'd11, 27'h00000115, 5'd24, 27'h000002e5, 5'd6, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000153, 5'd22, 27'h0000017a, 5'd17, 27'h00000004, 32'h00000400,
  1'd1,  5'd11, 27'h00000018, 5'd21, 27'h000000cb, 5'd28, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002e3, 5'd3, 27'h00000207, 5'd7, 27'h000001ad, 32'h00000400,
  1'd1,  5'd21, 27'h00000191, 5'd2, 27'h000001a8, 5'd20, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000056, 5'd4, 27'h00000013, 5'd26, 27'h00000009, 32'h00000400,
  1'd1,  5'd25, 27'h000000ce, 5'd13, 27'h000002f5, 5'd5, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000108, 5'd13, 27'h00000013, 5'd20, 27'h000000be, 32'h00000400,
  1'd1,  5'd23, 27'h0000011e, 5'd14, 27'h000001ba, 5'd28, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b7, 5'd21, 27'h000003f2, 5'd6, 27'h00000016, 32'h00000400,
  1'd1,  5'd22, 27'h00000250, 5'd22, 27'h0000039d, 5'd19, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f3, 5'd23, 27'h000003fa, 5'd28, 27'h000003ff, 32'h00000400,
  1'd1,  5'd0, 27'h0000005d, 5'd9, 27'h000003f0, 5'd2, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000175, 5'd5, 27'h0000010c, 5'd15, 27'h0000003d, 32'h00000400,
  1'd1,  5'd1, 27'h0000013e, 5'd8, 27'h0000009a, 5'd24, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000107, 5'd20, 27'h00000067, 5'd2, 27'h00000298, 32'h00000400,
  1'd1,  5'd4, 27'h0000018e, 5'd17, 27'h00000129, 5'd12, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000381, 5'd16, 27'h000000f3, 5'd24, 27'h000000c1, 32'h00000400,
  1'd1,  5'd2, 27'h0000007b, 5'd29, 27'h000002ab, 5'd0, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000006a, 5'd26, 27'h00000180, 5'd10, 27'h000003c8, 32'h00000400,
  1'd1,  5'd3, 27'h000002ea, 5'd27, 27'h00000041, 5'd22, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000203, 5'd8, 27'h000002bd, 5'd0, 27'h000000a7, 32'h00000400,
  1'd1,  5'd12, 27'h00000223, 5'd8, 27'h00000328, 5'd10, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000204, 5'd9, 27'h00000153, 5'd24, 27'h000003ae, 32'h00000400,
  1'd1,  5'd11, 27'h000000d5, 5'd18, 27'h000003d5, 5'd3, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000258, 5'd19, 27'h000000c4, 5'd12, 27'h000003b3, 32'h00000400,
  1'd1,  5'd12, 27'h0000023b, 5'd18, 27'h000001a2, 5'd21, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000300, 5'd29, 27'h00000175, 5'd2, 27'h000000cb, 32'h00000400,
  1'd1,  5'd15, 27'h0000019c, 5'd25, 27'h00000371, 5'd11, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003fa, 5'd27, 27'h000002e8, 5'd22, 27'h0000014d, 32'h00000400,
  1'd1,  5'd20, 27'h00000316, 5'd6, 27'h0000009d, 5'd2, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000202, 5'd6, 27'h000003ec, 5'd15, 27'h0000009a, 32'h00000400,
  1'd1,  5'd22, 27'h0000025e, 5'd6, 27'h00000264, 5'd25, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000203, 5'd20, 27'h00000192, 5'd4, 27'h0000004d, 32'h00000400,
  1'd1,  5'd25, 27'h000001dd, 5'd19, 27'h000000c6, 5'd11, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f4, 5'd19, 27'h0000002e, 5'd23, 27'h000002b7, 32'h00000400,
  1'd1,  5'd24, 27'h00000046, 5'd28, 27'h00000331, 5'd2, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000003f, 5'd30, 27'h00000239, 5'd11, 27'h000000c0, 32'h00000400,
  1'd1,  5'd22, 27'h00000077, 5'd28, 27'h000002b5, 5'd25, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000235, 5'd7, 27'h00000234, 5'd9, 27'h00000049, 32'h00000400,
  1'd1,  5'd1, 27'h0000027d, 5'd5, 27'h000002ed, 5'd16, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026f, 5'd5, 27'h000000cd, 5'd30, 27'h00000067, 32'h00000400,
  1'd1,  5'd2, 27'h000003c8, 5'd20, 27'h00000044, 5'd10, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002a4, 5'd15, 27'h000002a1, 5'd17, 27'h0000031f, 32'h00000400,
  1'd1,  5'd2, 27'h00000064, 5'd16, 27'h00000379, 5'd26, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000047, 5'd26, 27'h0000020d, 5'd8, 27'h000000b5, 32'h00000400,
  1'd1,  5'd0, 27'h000003a9, 5'd28, 27'h0000020d, 5'd15, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000270, 5'd29, 27'h0000008a, 5'd26, 27'h000003dd, 32'h00000400,
  1'd1,  5'd12, 27'h000000a3, 5'd10, 27'h0000012a, 5'd5, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000040, 5'd6, 27'h00000331, 5'd20, 27'h000000e2, 32'h00000400,
  1'd1,  5'd14, 27'h0000035f, 5'd6, 27'h000003c7, 5'd30, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d0, 5'd20, 27'h00000013, 5'd6, 27'h0000038e, 32'h00000400,
  1'd1,  5'd10, 27'h00000209, 5'd18, 27'h000003d2, 5'd16, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000114, 5'd18, 27'h000001f6, 5'd30, 27'h00000225, 32'h00000400,
  1'd1,  5'd11, 27'h00000021, 5'd26, 27'h00000393, 5'd7, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001ec, 5'd28, 27'h000002d7, 5'd16, 27'h0000034c, 32'h00000400,
  1'd1,  5'd11, 27'h0000037a, 5'd30, 27'h000000e1, 5'd30, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003ae, 5'd9, 27'h0000032c, 5'd8, 27'h000003d1, 32'h00000400,
  1'd1,  5'd22, 27'h000003d9, 5'd9, 27'h0000031c, 5'd17, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000392, 5'd6, 27'h00000225, 5'd25, 27'h000003d8, 32'h00000400,
  1'd1,  5'd25, 27'h0000011b, 5'd19, 27'h00000130, 5'd7, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001f2, 5'd18, 27'h00000234, 5'd15, 27'h0000026d, 32'h00000400,
  1'd1,  5'd24, 27'h0000039f, 5'd15, 27'h0000027d, 5'd27, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001b9, 5'd27, 27'h000003f6, 5'd8, 27'h00000338, 32'h00000400,
  1'd1,  5'd25, 27'h000001d2, 5'd30, 27'h000001f1, 5'd17, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000222, 5'd29, 27'h000001ba, 5'd29, 27'h000002ae, 32'h00000400,
  1'd1,  5'd5, 27'h000001a8, 5'd3, 27'h00000193, 5'd8, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002c8, 5'd2, 27'h000002c2, 5'd17, 27'h00000285, 32'h00000400,
  1'd1,  5'd5, 27'h000001d1, 5'd4, 27'h00000346, 5'd28, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c3, 5'd10, 27'h0000026a, 5'd0, 27'h0000022a, 32'h00000400,
  1'd1,  5'd5, 27'h00000138, 5'd14, 27'h000001ec, 5'd14, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000030a, 5'd10, 27'h00000389, 5'd25, 27'h00000012, 32'h00000400,
  1'd1,  5'd6, 27'h00000240, 5'd23, 27'h00000372, 5'd1, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000067, 5'd24, 27'h000000f6, 5'd14, 27'h0000015d, 32'h00000400,
  1'd1,  5'd6, 27'h0000026e, 5'd21, 27'h00000059, 5'd24, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000ff, 5'd2, 27'h0000001a, 5'd7, 27'h0000006e, 32'h00000400,
  1'd1,  5'd17, 27'h0000004e, 5'd3, 27'h000000cf, 5'd15, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000013a, 5'd2, 27'h000003ea, 5'd26, 27'h00000195, 32'h00000400,
  1'd1,  5'd16, 27'h00000243, 5'd12, 27'h00000259, 5'd1, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000071, 5'd11, 27'h00000240, 5'd11, 27'h0000014a, 32'h00000400,
  1'd1,  5'd17, 27'h000002d2, 5'd11, 27'h00000095, 5'd24, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003cf, 5'd25, 27'h0000015d, 5'd4, 27'h00000166, 32'h00000400,
  1'd1,  5'd15, 27'h000002a4, 5'd22, 27'h000002ee, 5'd12, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000046, 5'd21, 27'h000001b9, 5'd25, 27'h0000022b, 32'h00000400,
  1'd1,  5'd30, 27'h00000353, 5'd3, 27'h0000038e, 5'd1, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000012f, 5'd3, 27'h000003d2, 5'd14, 27'h000000c1, 32'h00000400,
  1'd1,  5'd28, 27'h00000135, 5'd1, 27'h0000005e, 5'd20, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003c3, 5'd12, 27'h0000002c, 5'd1, 27'h000001d4, 32'h00000400,
  1'd1,  5'd28, 27'h000000c8, 5'd11, 27'h000001d4, 5'd13, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000352, 5'd15, 27'h00000054, 5'd21, 27'h0000014e, 32'h00000400,
  1'd1,  5'd27, 27'h0000005c, 5'd21, 27'h00000074, 5'd5, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ae, 5'd25, 27'h000000a3, 5'd12, 27'h0000029f, 32'h00000400,
  1'd1,  5'd28, 27'h00000387, 5'd21, 27'h0000005e, 5'd24, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000390, 5'd1, 27'h0000004b, 5'd2, 27'h000001c2, 32'h00000400,
  1'd1,  5'd7, 27'h00000001, 5'd4, 27'h000002bc, 5'd15, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000391, 5'd3, 27'h00000294, 5'd24, 27'h0000026c, 32'h00000400,
  1'd1,  5'd5, 27'h000001c6, 5'd12, 27'h0000006d, 5'd6, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000004, 5'd12, 27'h00000373, 5'd17, 27'h00000250, 32'h00000400,
  1'd1,  5'd7, 27'h000000e0, 5'd12, 27'h00000041, 5'd29, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000019a, 5'd23, 27'h000002eb, 5'd8, 27'h0000015c, 32'h00000400,
  1'd1,  5'd9, 27'h0000007d, 5'd22, 27'h00000344, 5'd20, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000011, 5'd22, 27'h00000083, 5'd29, 27'h0000037a, 32'h00000400,
  1'd1,  5'd20, 27'h0000013e, 5'd3, 27'h00000012, 5'd2, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000293, 5'd1, 27'h000003c3, 5'd15, 27'h00000008, 32'h00000400,
  1'd1,  5'd15, 27'h00000257, 5'd2, 27'h00000008, 5'd20, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001db, 5'd13, 27'h000001a5, 5'd10, 27'h00000082, 32'h00000400,
  1'd1,  5'd19, 27'h00000084, 5'd14, 27'h00000391, 5'd19, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000370, 5'd12, 27'h000001be, 5'd30, 27'h000000ee, 32'h00000400,
  1'd1,  5'd17, 27'h0000017c, 5'd21, 27'h000000e9, 5'd7, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e1, 5'd22, 27'h000000d3, 5'd16, 27'h00000055, 32'h00000400,
  1'd1,  5'd16, 27'h000002b8, 5'd20, 27'h00000329, 5'd25, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000121, 5'd3, 27'h00000037, 5'd8, 27'h000000d0, 32'h00000400,
  1'd1,  5'd26, 27'h00000031, 5'd0, 27'h000001df, 5'd19, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000321, 5'd3, 27'h000003f5, 5'd27, 27'h00000107, 32'h00000400,
  1'd1,  5'd29, 27'h0000030f, 5'd12, 27'h00000313, 5'd6, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ec, 5'd15, 27'h00000161, 5'd16, 27'h00000097, 32'h00000400,
  1'd1,  5'd30, 27'h000003f2, 5'd12, 27'h000001cf, 5'd30, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003e2, 5'd22, 27'h00000035, 5'd8, 27'h0000035b, 32'h00000400,
  1'd1,  5'd30, 27'h0000028b, 5'd25, 27'h00000054, 5'd18, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000235, 5'd25, 27'h00000067, 5'd29, 27'h000001f0, 32'h00000400,
  1'd1,  5'd6, 27'h00000057, 5'd5, 27'h00000257, 5'd4, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001bd, 5'd10, 27'h000000bd, 5'd10, 27'h00000163, 32'h00000400,
  1'd1,  5'd6, 27'h0000004f, 5'd5, 27'h00000171, 5'd22, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b0, 5'd18, 27'h00000082, 5'd3, 27'h000003ed, 32'h00000400,
  1'd1,  5'd9, 27'h00000308, 5'd18, 27'h000001ce, 5'd12, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000349, 5'd20, 27'h00000102, 5'd23, 27'h0000036b, 32'h00000400,
  1'd1,  5'd9, 27'h00000262, 5'd29, 27'h00000030, 5'd3, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000015d, 5'd26, 27'h00000117, 5'd12, 27'h0000033a, 32'h00000400,
  1'd1,  5'd6, 27'h00000093, 5'd26, 27'h000002a5, 5'd23, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000397, 5'd9, 27'h0000022f, 5'd1, 27'h00000229, 32'h00000400,
  1'd1,  5'd18, 27'h00000003, 5'd9, 27'h00000035, 5'd14, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000017, 5'd6, 27'h000001ca, 5'd21, 27'h00000001, 32'h00000400,
  1'd1,  5'd17, 27'h00000306, 5'd18, 27'h0000018e, 5'd2, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d1, 5'd15, 27'h00000379, 5'd12, 27'h000002e9, 32'h00000400,
  1'd1,  5'd19, 27'h00000334, 5'd17, 27'h000003fd, 5'd23, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000231, 5'd26, 27'h00000031, 5'd3, 27'h00000006, 32'h00000400,
  1'd1,  5'd19, 27'h00000333, 5'd30, 27'h000003f7, 5'd15, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002f7, 5'd29, 27'h00000168, 5'd21, 27'h00000008, 32'h00000400,
  1'd1,  5'd26, 27'h00000079, 5'd9, 27'h000001e4, 5'd2, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000172, 5'd5, 27'h000000fb, 5'd10, 27'h00000381, 32'h00000400,
  1'd1,  5'd30, 27'h00000010, 5'd9, 27'h0000005a, 5'd24, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000022, 5'd16, 27'h000002e5, 5'd3, 27'h0000012d, 32'h00000400,
  1'd1,  5'd27, 27'h00000202, 5'd15, 27'h000002fc, 5'd11, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000289, 5'd19, 27'h000000c8, 5'd22, 27'h000002c1, 32'h00000400,
  1'd1,  5'd30, 27'h0000001a, 5'd29, 27'h0000001c, 5'd2, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000291, 5'd27, 27'h000001f2, 5'd11, 27'h0000024a, 32'h00000400,
  1'd1,  5'd26, 27'h0000036e, 5'd27, 27'h0000011d, 5'd22, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000012d, 5'd5, 27'h00000211, 5'd8, 27'h000002cc, 32'h00000400,
  1'd1,  5'd10, 27'h00000047, 5'd9, 27'h00000343, 5'd17, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000165, 5'd5, 27'h000000c6, 5'd27, 27'h00000186, 32'h00000400,
  1'd1,  5'd8, 27'h0000013d, 5'd18, 27'h000003ac, 5'd7, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e4, 5'd18, 27'h000001d5, 5'd16, 27'h000000ba, 32'h00000400,
  1'd1,  5'd8, 27'h00000341, 5'd18, 27'h00000146, 5'd30, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002ee, 5'd26, 27'h000001e2, 5'd9, 27'h00000060, 32'h00000400,
  1'd1,  5'd9, 27'h000000dd, 5'd27, 27'h0000016a, 5'd16, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000aa, 5'd30, 27'h00000012, 5'd26, 27'h0000009e, 32'h00000400,
  1'd1,  5'd18, 27'h00000087, 5'd8, 27'h000002a4, 5'd9, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000019f, 5'd8, 27'h000000ce, 5'd15, 27'h000002e0, 32'h00000400,
  1'd1,  5'd19, 27'h00000374, 5'd10, 27'h00000103, 5'd28, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a3, 5'd18, 27'h0000025c, 5'd5, 27'h000002f4, 32'h00000400,
  1'd1,  5'd18, 27'h000003f5, 5'd17, 27'h0000002e, 5'd20, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002bd, 5'd16, 27'h00000170, 5'd30, 27'h000002ec, 32'h00000400,
  1'd1,  5'd18, 27'h000003f4, 5'd26, 27'h0000034f, 5'd10, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000164, 5'd29, 27'h000000da, 5'd16, 27'h00000348, 32'h00000400,
  1'd1,  5'd18, 27'h0000003f, 5'd29, 27'h000000c8, 5'd30, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001a0, 5'd9, 27'h00000154, 5'd8, 27'h0000028a, 32'h00000400,
  1'd1,  5'd25, 27'h00000390, 5'd5, 27'h00000303, 5'd18, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000013c, 5'd8, 27'h0000022a, 5'd30, 27'h000002cc, 32'h00000400,
  1'd1,  5'd26, 27'h000002f2, 5'd20, 27'h00000116, 5'd8, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ec, 5'd18, 27'h000001c4, 5'd19, 27'h000003e6, 32'h00000400,
  1'd1,  5'd28, 27'h00000267, 5'd20, 27'h000001b0, 5'd25, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000222, 5'd27, 27'h00000386, 5'd9, 27'h00000293, 32'h00000400,
  1'd1,  5'd27, 27'h000003bc, 5'd30, 27'h00000146, 5'd17, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000032f, 5'd26, 27'h000003f1, 5'd27, 27'h00000370, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000001aa, 5'd3, 27'h000000d4, 5'd0, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002aa, 5'd1, 27'h00000290, 5'd13, 27'h00000106, 32'h00000400,
  1'd1,  5'd1, 27'h0000002e, 5'd3, 27'h0000005b, 5'd21, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000c2, 5'd12, 27'h000001df, 5'd1, 27'h00000095, 32'h00000400,
  1'd1,  5'd0, 27'h000000d1, 5'd13, 27'h00000357, 5'd12, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000204, 5'd13, 27'h00000248, 5'd20, 27'h0000033f, 32'h00000400,
  1'd1,  5'd2, 27'h00000285, 5'd24, 27'h000001d8, 5'd5, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003e7, 5'd24, 27'h0000024e, 5'd14, 27'h00000279, 32'h00000400,
  1'd1,  5'd3, 27'h0000006f, 5'd23, 27'h000003de, 5'd23, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000020d, 5'd3, 27'h00000268, 5'd2, 27'h000000d7, 32'h00000400,
  1'd1,  5'd10, 27'h000002df, 5'd0, 27'h000002fd, 5'd10, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003cf, 5'd2, 27'h00000260, 5'd22, 27'h000003a9, 32'h00000400,
  1'd1,  5'd12, 27'h000003a1, 5'd10, 27'h000002cf, 5'd3, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000016e, 5'd12, 27'h0000009e, 5'd12, 27'h0000030f, 32'h00000400,
  1'd1,  5'd10, 27'h0000019f, 5'd15, 27'h00000188, 5'd22, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000304, 5'd22, 27'h000001d9, 5'd0, 27'h00000245, 32'h00000400,
  1'd1,  5'd10, 27'h0000039e, 5'd22, 27'h0000022a, 5'd10, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000017c, 5'd22, 27'h0000036e, 5'd23, 27'h0000011e, 32'h00000400,
  1'd1,  5'd20, 27'h00000389, 5'd2, 27'h000002e2, 5'd4, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ae, 5'd2, 27'h0000010a, 5'd13, 27'h000000b5, 32'h00000400,
  1'd1,  5'd25, 27'h000000bb, 5'd4, 27'h00000325, 5'd24, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022f, 5'd13, 27'h00000188, 5'd2, 27'h000001d8, 32'h00000400,
  1'd1,  5'd22, 27'h000003a5, 5'd11, 27'h000000f5, 5'd14, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a1, 5'd12, 27'h00000388, 5'd24, 27'h000003f3, 32'h00000400,
  1'd1,  5'd24, 27'h00000139, 5'd22, 27'h00000212, 5'd2, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000099, 5'd24, 27'h00000341, 5'd13, 27'h00000239, 32'h00000400,
  1'd1,  5'd22, 27'h0000029e, 5'd24, 27'h00000080, 5'd25, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000297, 5'd0, 27'h00000316, 5'd9, 27'h00000027, 32'h00000400,
  1'd1,  5'd1, 27'h00000002, 5'd2, 27'h00000203, 5'd17, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000304, 5'd0, 27'h000002b6, 5'd29, 27'h00000037, 32'h00000400,
  1'd1,  5'd0, 27'h000000b9, 5'd14, 27'h00000380, 5'd9, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f3, 5'd12, 27'h0000023e, 5'd17, 27'h00000274, 32'h00000400,
  1'd1,  5'd2, 27'h00000388, 5'd11, 27'h00000038, 5'd29, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000074, 5'd21, 27'h0000005a, 5'd9, 27'h00000331, 32'h00000400,
  1'd1,  5'd0, 27'h0000019f, 5'd22, 27'h000000ee, 5'd19, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000007d, 5'd24, 27'h0000036f, 5'd29, 27'h00000106, 32'h00000400,
  1'd1,  5'd12, 27'h000000d8, 5'd4, 27'h00000243, 5'd6, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003c4, 5'd2, 27'h0000030c, 5'd15, 27'h00000274, 32'h00000400,
  1'd1,  5'd13, 27'h000001c6, 5'd3, 27'h000003f2, 5'd28, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034c, 5'd10, 27'h00000302, 5'd9, 27'h00000215, 32'h00000400,
  1'd1,  5'd12, 27'h00000143, 5'd14, 27'h000002e9, 5'd17, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b1, 5'd14, 27'h000003b4, 5'd26, 27'h0000013b, 32'h00000400,
  1'd1,  5'd14, 27'h0000002b, 5'd23, 27'h0000007c, 5'd5, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c5, 5'd21, 27'h0000024d, 5'd20, 27'h0000025a, 32'h00000400,
  1'd1,  5'd12, 27'h0000007c, 5'd24, 27'h00000012, 5'd30, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002bc, 5'd4, 27'h000003ab, 5'd7, 27'h000003fc, 32'h00000400,
  1'd1,  5'd23, 27'h000002a6, 5'd2, 27'h0000035a, 5'd15, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000008b, 5'd4, 27'h000003eb, 5'd30, 27'h000003fa, 32'h00000400,
  1'd1,  5'd22, 27'h0000030c, 5'd12, 27'h00000306, 5'd7, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000175, 5'd10, 27'h000003be, 5'd15, 27'h00000373, 32'h00000400,
  1'd1,  5'd22, 27'h00000011, 5'd13, 27'h000002ab, 5'd30, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e8, 5'd21, 27'h00000395, 5'd9, 27'h000002d4, 32'h00000400,
  1'd1,  5'd24, 27'h00000162, 5'd24, 27'h000003c7, 5'd16, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003bc, 5'd24, 27'h000003a6, 5'd29, 27'h000000c4, 32'h00000400,
  1'd1,  5'd2, 27'h000003a4, 5'd10, 27'h0000009c, 5'd1, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003fb, 5'd9, 27'h00000116, 5'd14, 27'h000002ba, 32'h00000400,
  1'd1,  5'd0, 27'h000001ee, 5'd9, 27'h00000093, 5'd25, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018d, 5'd19, 27'h00000048, 5'd3, 27'h000002b0, 32'h00000400,
  1'd1,  5'd1, 27'h000001d0, 5'd20, 27'h00000135, 5'd11, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000303, 5'd16, 27'h00000164, 5'd21, 27'h00000031, 32'h00000400,
  1'd1,  5'd4, 27'h00000146, 5'd26, 27'h0000007c, 5'd4, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000107, 5'd26, 27'h000003de, 5'd12, 27'h00000071, 32'h00000400,
  1'd1,  5'd1, 27'h000002ad, 5'd28, 27'h000001ce, 5'd22, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000004, 5'd9, 27'h000001ce, 5'd1, 27'h0000031b, 32'h00000400,
  1'd1,  5'd14, 27'h000002b4, 5'd9, 27'h000001c5, 5'd12, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000021d, 5'd7, 27'h000000ca, 5'd22, 27'h00000199, 32'h00000400,
  1'd1,  5'd13, 27'h00000396, 5'd18, 27'h00000076, 5'd0, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000b3, 5'd19, 27'h0000009b, 5'd13, 27'h00000051, 32'h00000400,
  1'd1,  5'd10, 27'h000001f5, 5'd16, 27'h00000262, 5'd23, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ea, 5'd28, 27'h000003b8, 5'd2, 27'h00000386, 32'h00000400,
  1'd1,  5'd14, 27'h000001c0, 5'd30, 27'h000000a6, 5'd12, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000354, 5'd26, 27'h00000262, 5'd21, 27'h00000099, 32'h00000400,
  1'd1,  5'd25, 27'h0000026f, 5'd8, 27'h0000003c, 5'd4, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000175, 5'd7, 27'h00000051, 5'd10, 27'h00000320, 32'h00000400,
  1'd1,  5'd22, 27'h000001f8, 5'd7, 27'h000001bf, 5'd24, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000ce, 5'd19, 27'h00000257, 5'd1, 27'h0000002c, 32'h00000400,
  1'd1,  5'd20, 27'h0000036d, 5'd17, 27'h000002b0, 5'd12, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000309, 5'd20, 27'h00000036, 5'd22, 27'h0000010a, 32'h00000400,
  1'd1,  5'd22, 27'h000003bd, 5'd29, 27'h0000012e, 5'd3, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000030d, 5'd30, 27'h000000f7, 5'd13, 27'h00000168, 32'h00000400,
  1'd1,  5'd24, 27'h0000026d, 5'd29, 27'h00000149, 5'd23, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000234, 5'd5, 27'h00000231, 5'd8, 27'h000003fd, 32'h00000400,
  1'd1,  5'd4, 27'h000000e4, 5'd8, 27'h00000262, 5'd18, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000024e, 5'd9, 27'h00000040, 5'd25, 27'h000003f9, 32'h00000400,
  1'd1,  5'd3, 27'h000003a1, 5'd18, 27'h000002d5, 5'd8, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036d, 5'd18, 27'h000002ea, 5'd19, 27'h000000a2, 32'h00000400,
  1'd1,  5'd2, 27'h000000e4, 5'd20, 27'h00000209, 5'd28, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000024d, 5'd27, 27'h00000336, 5'd9, 27'h0000038e, 32'h00000400,
  1'd1,  5'd4, 27'h0000002c, 5'd27, 27'h000003d8, 5'd20, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000c3, 5'd27, 27'h00000222, 5'd28, 27'h000000ff, 32'h00000400,
  1'd1,  5'd10, 27'h00000273, 5'd10, 27'h00000063, 5'd6, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000017f, 5'd7, 27'h00000102, 5'd18, 27'h000000d0, 32'h00000400,
  1'd1,  5'd14, 27'h0000000c, 5'd8, 27'h000000da, 5'd28, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000147, 5'd19, 27'h00000273, 5'd6, 27'h0000023e, 32'h00000400,
  1'd1,  5'd12, 27'h000001a8, 5'd16, 27'h0000010e, 5'd16, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000309, 5'd18, 27'h000003e5, 5'd27, 27'h00000054, 32'h00000400,
  1'd1,  5'd11, 27'h0000039e, 5'd29, 27'h00000118, 5'd9, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002a1, 5'd29, 27'h000003a1, 5'd16, 27'h0000004b, 32'h00000400,
  1'd1,  5'd11, 27'h0000024a, 5'd26, 27'h00000340, 5'd27, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000377, 5'd6, 27'h000000cb, 5'd5, 27'h00000137, 32'h00000400,
  1'd1,  5'd20, 27'h00000386, 5'd8, 27'h00000174, 5'd19, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000339, 5'd5, 27'h00000259, 5'd29, 27'h00000169, 32'h00000400,
  1'd1,  5'd24, 27'h000002d7, 5'd20, 27'h000001a5, 5'd5, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003fa, 5'd17, 27'h000002e1, 5'd19, 27'h00000238, 32'h00000400,
  1'd1,  5'd24, 27'h000001cf, 5'd17, 27'h000000c3, 5'd26, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000034f, 5'd27, 27'h00000105, 5'd8, 27'h0000002d, 32'h00000400,
  1'd1,  5'd23, 27'h00000248, 5'd26, 27'h000001bf, 5'd17, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000029d, 5'd26, 27'h000001be, 5'd28, 27'h000002ef, 32'h00000400,
  1'd1,  5'd7, 27'h00000254, 5'd0, 27'h0000036f, 5'd7, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012a, 5'd3, 27'h00000218, 5'd16, 27'h0000018c, 32'h00000400,
  1'd1,  5'd5, 27'h0000018e, 5'd1, 27'h000000a5, 5'd28, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000314, 5'd13, 27'h00000182, 5'd2, 27'h00000022, 32'h00000400,
  1'd1,  5'd5, 27'h00000398, 5'd12, 27'h000003c8, 5'd13, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003fa, 5'd10, 27'h000002dc, 5'd25, 27'h0000034c, 32'h00000400,
  1'd1,  5'd10, 27'h00000097, 5'd23, 27'h000001de, 5'd0, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001e8, 5'd20, 27'h000002fa, 5'd14, 27'h0000009b, 32'h00000400,
  1'd1,  5'd8, 27'h000000d5, 5'd24, 27'h00000158, 5'd22, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000002e, 5'd5, 27'h00000074, 5'd7, 27'h0000024e, 32'h00000400,
  1'd1,  5'd17, 27'h000002b5, 5'd2, 27'h0000020a, 5'd16, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000bd, 5'd0, 27'h00000277, 5'd29, 27'h000003e1, 32'h00000400,
  1'd1,  5'd20, 27'h000000d6, 5'd13, 27'h00000323, 5'd1, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000208, 5'd11, 27'h0000022a, 5'd15, 27'h00000041, 32'h00000400,
  1'd1,  5'd17, 27'h0000031e, 5'd14, 27'h00000054, 5'd22, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000026b, 5'd22, 27'h000003f8, 5'd4, 27'h0000028c, 32'h00000400,
  1'd1,  5'd15, 27'h000002a2, 5'd22, 27'h0000004a, 5'd11, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002fd, 5'd25, 27'h00000263, 5'd21, 27'h00000087, 32'h00000400,
  1'd1,  5'd26, 27'h000000c1, 5'd4, 27'h0000027b, 5'd4, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000031b, 5'd2, 27'h000002cd, 5'd10, 27'h00000373, 32'h00000400,
  1'd1,  5'd26, 27'h00000296, 5'd0, 27'h00000080, 5'd23, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000022e, 5'd12, 27'h000003f5, 5'd4, 27'h00000298, 32'h00000400,
  1'd1,  5'd26, 27'h000001a3, 5'd14, 27'h00000281, 5'd11, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000194, 5'd14, 27'h00000244, 5'd22, 27'h00000162, 32'h00000400,
  1'd1,  5'd30, 27'h000002de, 5'd23, 27'h000000f0, 5'd0, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000b3, 5'd22, 27'h000003cc, 5'd11, 27'h000001c5, 32'h00000400,
  1'd1,  5'd29, 27'h00000103, 5'd20, 27'h000003f4, 5'd25, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b2, 5'd3, 27'h00000245, 5'd2, 27'h0000035d, 32'h00000400,
  1'd1,  5'd8, 27'h0000034c, 5'd1, 27'h0000012d, 5'd13, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000005d, 5'd4, 27'h00000121, 5'd21, 27'h000001c0, 32'h00000400,
  1'd1,  5'd6, 27'h00000352, 5'd14, 27'h00000113, 5'd6, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002ef, 5'd15, 27'h0000005d, 5'd17, 27'h000002da, 32'h00000400,
  1'd1,  5'd8, 27'h00000186, 5'd14, 27'h00000216, 5'd29, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003cc, 5'd22, 27'h00000228, 5'd9, 27'h0000009a, 32'h00000400,
  1'd1,  5'd10, 27'h000000bb, 5'd23, 27'h000002a0, 5'd18, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000039e, 5'd22, 27'h0000014f, 5'd27, 27'h00000251, 32'h00000400,
  1'd1,  5'd17, 27'h00000265, 5'd3, 27'h0000029b, 5'd3, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000027a, 5'd5, 27'h0000004b, 5'd12, 27'h000000e1, 32'h00000400,
  1'd1,  5'd18, 27'h00000059, 5'd4, 27'h00000087, 5'd24, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000031b, 5'd10, 27'h000002a9, 5'd7, 27'h000000f9, 32'h00000400,
  1'd1,  5'd19, 27'h000000c1, 5'd14, 27'h0000039b, 5'd20, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000168, 5'd10, 27'h0000029e, 5'd26, 27'h0000038c, 32'h00000400,
  1'd1,  5'd17, 27'h0000023d, 5'd24, 27'h00000361, 5'd5, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000360, 5'd23, 27'h00000212, 5'd20, 27'h00000258, 32'h00000400,
  1'd1,  5'd17, 27'h00000106, 5'd24, 27'h00000370, 5'd26, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000205, 5'd4, 27'h00000010, 5'd6, 27'h00000224, 32'h00000400,
  1'd1,  5'd26, 27'h00000272, 5'd1, 27'h00000260, 5'd19, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ad, 5'd0, 27'h00000186, 5'd30, 27'h00000001, 32'h00000400,
  1'd1,  5'd28, 27'h00000186, 5'd11, 27'h00000003, 5'd9, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000f2, 5'd11, 27'h00000037, 5'd17, 27'h000002f6, 32'h00000400,
  1'd1,  5'd27, 27'h00000371, 5'd10, 27'h0000018d, 5'd29, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003a3, 5'd24, 27'h00000114, 5'd6, 27'h0000018e, 32'h00000400,
  1'd1,  5'd26, 27'h000002e4, 5'd21, 27'h0000010f, 5'd17, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003bf, 5'd22, 27'h00000107, 5'd28, 27'h00000042, 32'h00000400,
  1'd1,  5'd5, 27'h000001cb, 5'd8, 27'h000001e6, 5'd2, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000289, 5'd9, 27'h00000179, 5'd10, 27'h00000347, 32'h00000400,
  1'd1,  5'd8, 27'h0000018f, 5'd6, 27'h00000329, 5'd23, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ef, 5'd16, 27'h0000031f, 5'd4, 27'h00000141, 32'h00000400,
  1'd1,  5'd6, 27'h00000111, 5'd17, 27'h0000003b, 5'd12, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a0, 5'd16, 27'h00000271, 5'd25, 27'h0000031c, 32'h00000400,
  1'd1,  5'd9, 27'h00000202, 5'd29, 27'h000001cd, 5'd5, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000133, 5'd29, 27'h00000045, 5'd13, 27'h00000358, 32'h00000400,
  1'd1,  5'd8, 27'h00000310, 5'd26, 27'h00000261, 5'd25, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e8, 5'd9, 27'h00000130, 5'd3, 27'h000000f1, 32'h00000400,
  1'd1,  5'd16, 27'h000001cf, 5'd8, 27'h000003f2, 5'd13, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000d0, 5'd9, 27'h0000036e, 5'd25, 27'h0000024d, 32'h00000400,
  1'd1,  5'd18, 27'h0000038c, 5'd15, 27'h000002bb, 5'd1, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000135, 5'd20, 27'h0000010d, 5'd14, 27'h0000027a, 32'h00000400,
  1'd1,  5'd16, 27'h000001ff, 5'd17, 27'h00000001, 5'd21, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000075, 5'd29, 27'h000000d3, 5'd0, 27'h000000e5, 32'h00000400,
  1'd1,  5'd18, 27'h00000168, 5'd28, 27'h0000019e, 5'd13, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000017a, 5'd28, 27'h00000253, 5'd24, 27'h00000097, 32'h00000400,
  1'd1,  5'd26, 27'h000002f8, 5'd8, 27'h00000163, 5'd3, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000022, 5'd8, 27'h00000209, 5'd11, 27'h0000027e, 32'h00000400,
  1'd1,  5'd26, 27'h0000027d, 5'd9, 27'h000001c2, 5'd24, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000007, 5'd17, 27'h00000294, 5'd1, 27'h000003b8, 32'h00000400,
  1'd1,  5'd29, 27'h000000a4, 5'd19, 27'h00000090, 5'd13, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a8, 5'd19, 27'h00000345, 5'd22, 27'h00000236, 32'h00000400,
  1'd1,  5'd26, 27'h00000252, 5'd28, 27'h0000008b, 5'd1, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003d0, 5'd29, 27'h000002c2, 5'd11, 27'h00000049, 32'h00000400,
  1'd1,  5'd28, 27'h000000e8, 5'd26, 27'h00000332, 5'd25, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000010, 5'd9, 27'h000000dc, 5'd5, 27'h00000213, 32'h00000400,
  1'd1,  5'd8, 27'h000003c1, 5'd9, 27'h00000313, 5'd18, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003eb, 5'd7, 27'h0000016f, 5'd29, 27'h000000c4, 32'h00000400,
  1'd1,  5'd6, 27'h00000128, 5'd16, 27'h00000190, 5'd6, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a0, 5'd20, 27'h000001b5, 5'd18, 27'h0000038c, 32'h00000400,
  1'd1,  5'd6, 27'h00000105, 5'd20, 27'h0000005a, 5'd25, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003af, 5'd30, 27'h00000173, 5'd9, 27'h00000340, 32'h00000400,
  1'd1,  5'd8, 27'h00000046, 5'd30, 27'h000001e2, 5'd18, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000220, 5'd28, 27'h00000148, 5'd26, 27'h00000164, 32'h00000400,
  1'd1,  5'd16, 27'h00000018, 5'd5, 27'h000000bb, 5'd7, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f9, 5'd7, 27'h000002da, 5'd19, 27'h00000294, 32'h00000400,
  1'd1,  5'd19, 27'h0000037f, 5'd8, 27'h0000004d, 5'd29, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000096, 5'd19, 27'h000003c6, 5'd5, 27'h00000239, 32'h00000400,
  1'd1,  5'd20, 27'h00000214, 5'd15, 27'h000003ea, 5'd20, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000039a, 5'd20, 27'h000000c2, 5'd30, 27'h000000c2, 32'h00000400,
  1'd1,  5'd19, 27'h000002ea, 5'd30, 27'h00000326, 5'd5, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000b6, 5'd27, 27'h000003f5, 5'd18, 27'h000003ba, 32'h00000400,
  1'd1,  5'd19, 27'h00000381, 5'd30, 27'h0000034e, 5'd30, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000037c, 5'd7, 27'h00000379, 5'd9, 27'h000002e6, 32'h00000400,
  1'd1,  5'd30, 27'h000001ee, 5'd5, 27'h00000231, 5'd16, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000029d, 5'd7, 27'h000002c0, 5'd30, 27'h000000b1, 32'h00000400,
  1'd1,  5'd30, 27'h0000002d, 5'd18, 27'h0000021a, 5'd9, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000030e, 5'd18, 27'h00000089, 5'd17, 27'h0000008f, 32'h00000400,
  1'd1,  5'd30, 27'h000001de, 5'd17, 27'h000002ef, 5'd30, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000096, 5'd26, 27'h000002f1, 5'd5, 27'h0000026a, 32'h00000400,
  1'd1,  5'd28, 27'h00000080, 5'd28, 27'h0000018a, 5'd19, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000146, 5'd30, 27'h000002cb, 5'd26, 27'h00000179, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h00000032, 5'd1, 27'h000001c1, 5'd1, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001ac, 5'd3, 27'h0000000d, 5'd10, 27'h0000018a, 32'h00000400,
  1'd1,  5'd1, 27'h00000325, 5'd2, 27'h0000039a, 5'd22, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003c5, 5'd12, 27'h0000010e, 5'd3, 27'h000003c2, 32'h00000400,
  1'd1,  5'd3, 27'h000000f2, 5'd14, 27'h00000226, 5'd10, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000017a, 5'd12, 27'h00000254, 5'd21, 27'h000002eb, 32'h00000400,
  1'd1,  5'd0, 27'h000002a4, 5'd25, 27'h00000041, 5'd3, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b4, 5'd25, 27'h000000a0, 5'd10, 27'h000002c4, 32'h00000400,
  1'd1,  5'd1, 27'h000001b0, 5'd22, 27'h0000028e, 5'd24, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000c0, 5'd4, 27'h00000258, 5'd0, 27'h00000082, 32'h00000400,
  1'd1,  5'd13, 27'h000003af, 5'd2, 27'h0000012b, 5'd10, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000135, 5'd4, 27'h000003c6, 5'd24, 27'h000001ab, 32'h00000400,
  1'd1,  5'd13, 27'h0000020a, 5'd12, 27'h00000397, 5'd4, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000380, 5'd12, 27'h00000125, 5'd12, 27'h00000399, 32'h00000400,
  1'd1,  5'd12, 27'h00000197, 5'd13, 27'h0000024a, 5'd24, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000028d, 5'd22, 27'h0000024b, 5'd2, 27'h0000037e, 32'h00000400,
  1'd1,  5'd14, 27'h0000021d, 5'd22, 27'h0000037e, 5'd12, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000004a, 5'd23, 27'h000000b3, 5'd21, 27'h00000160, 32'h00000400,
  1'd1,  5'd22, 27'h000001e0, 5'd4, 27'h000002d6, 5'd0, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b8, 5'd4, 27'h0000020c, 5'd10, 27'h00000160, 32'h00000400,
  1'd1,  5'd20, 27'h000003f5, 5'd3, 27'h0000012d, 5'd24, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000342, 5'd13, 27'h000000c5, 5'd1, 27'h0000023f, 32'h00000400,
  1'd1,  5'd22, 27'h000002ba, 5'd12, 27'h000001b2, 5'd10, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000018e, 5'd12, 27'h00000328, 5'd21, 27'h000003d2, 32'h00000400,
  1'd1,  5'd22, 27'h00000239, 5'd25, 27'h000002c9, 5'd0, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002a0, 5'd24, 27'h0000039b, 5'd13, 27'h00000146, 32'h00000400,
  1'd1,  5'd22, 27'h0000032d, 5'd25, 27'h0000033f, 5'd23, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002df, 5'd4, 27'h00000056, 5'd5, 27'h00000365, 32'h00000400,
  1'd1,  5'd3, 27'h0000018d, 5'd5, 27'h0000000d, 5'd20, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000005f, 5'd4, 27'h000003d4, 5'd30, 27'h0000009b, 32'h00000400,
  1'd1,  5'd2, 27'h00000318, 5'd15, 27'h00000001, 5'd8, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a3, 5'd12, 27'h0000003a, 5'd19, 27'h000002bb, 32'h00000400,
  1'd1,  5'd4, 27'h000003de, 5'd11, 27'h00000260, 5'd28, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000010b, 5'd25, 27'h00000012, 5'd9, 27'h000000b0, 32'h00000400,
  1'd1,  5'd0, 27'h000001ff, 5'd22, 27'h000000d4, 5'd18, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a1, 5'd22, 27'h00000193, 5'd30, 27'h00000190, 32'h00000400,
  1'd1,  5'd12, 27'h00000088, 5'd5, 27'h00000073, 5'd6, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000172, 5'd3, 27'h000003e2, 5'd16, 27'h000000a5, 32'h00000400,
  1'd1,  5'd15, 27'h00000111, 5'd1, 27'h0000001a, 5'd29, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a4, 5'd12, 27'h00000042, 5'd6, 27'h000003aa, 32'h00000400,
  1'd1,  5'd10, 27'h000003a1, 5'd13, 27'h0000019e, 5'd16, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000300, 5'd15, 27'h0000007e, 5'd28, 27'h0000026f, 32'h00000400,
  1'd1,  5'd11, 27'h000003f0, 5'd24, 27'h000003c9, 5'd7, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003d6, 5'd22, 27'h00000386, 5'd16, 27'h0000017c, 32'h00000400,
  1'd1,  5'd13, 27'h000000b6, 5'd25, 27'h00000141, 5'd26, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000264, 5'd1, 27'h0000031f, 5'd8, 27'h00000268, 32'h00000400,
  1'd1,  5'd25, 27'h0000022f, 5'd3, 27'h00000337, 5'd17, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ae, 5'd0, 27'h000003ae, 5'd28, 27'h000001ce, 32'h00000400,
  1'd1,  5'd21, 27'h00000272, 5'd10, 27'h0000026a, 5'd6, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000364, 5'd12, 27'h0000034f, 5'd19, 27'h0000007a, 32'h00000400,
  1'd1,  5'd22, 27'h00000096, 5'd12, 27'h0000015a, 5'd30, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000072, 5'd21, 27'h00000126, 5'd5, 27'h000003e2, 32'h00000400,
  1'd1,  5'd25, 27'h0000018b, 5'd23, 27'h00000222, 5'd16, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c6, 5'd25, 27'h000001ae, 5'd27, 27'h00000298, 32'h00000400,
  1'd1,  5'd2, 27'h00000227, 5'd10, 27'h00000130, 5'd0, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000024e, 5'd5, 27'h00000393, 5'd14, 27'h000000ca, 32'h00000400,
  1'd1,  5'd3, 27'h00000142, 5'd9, 27'h00000377, 5'd23, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000086, 5'd16, 27'h000000cf, 5'd2, 27'h000000cb, 32'h00000400,
  1'd1,  5'd4, 27'h00000355, 5'd16, 27'h0000032a, 5'd12, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000015f, 5'd17, 27'h00000306, 5'd20, 27'h00000309, 32'h00000400,
  1'd1,  5'd5, 27'h0000006d, 5'd30, 27'h0000031b, 5'd1, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000013d, 5'd30, 27'h00000119, 5'd11, 27'h000002b6, 32'h00000400,
  1'd1,  5'd3, 27'h00000103, 5'd28, 27'h00000034, 5'd24, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000b2, 5'd7, 27'h000000c4, 5'd1, 27'h000002ca, 32'h00000400,
  1'd1,  5'd14, 27'h00000134, 5'd6, 27'h000001dc, 5'd14, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000031, 5'd5, 27'h00000275, 5'd22, 27'h000002ca, 32'h00000400,
  1'd1,  5'd11, 27'h00000178, 5'd19, 27'h00000099, 5'd0, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002b, 5'd18, 27'h000000f6, 5'd14, 27'h000001be, 32'h00000400,
  1'd1,  5'd12, 27'h0000012f, 5'd18, 27'h00000320, 5'd22, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000039d, 5'd30, 27'h000002e1, 5'd0, 27'h0000010b, 32'h00000400,
  1'd1,  5'd12, 27'h0000019d, 5'd29, 27'h000003e7, 5'd10, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f9, 5'd30, 27'h00000012, 5'd25, 27'h00000072, 32'h00000400,
  1'd1,  5'd23, 27'h000002aa, 5'd8, 27'h000002b8, 5'd3, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002da, 5'd8, 27'h00000238, 5'd12, 27'h00000129, 32'h00000400,
  1'd1,  5'd25, 27'h00000094, 5'd6, 27'h00000040, 5'd20, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000028f, 5'd15, 27'h0000027b, 5'd1, 27'h000000c4, 32'h00000400,
  1'd1,  5'd23, 27'h000000dc, 5'd18, 27'h00000239, 5'd11, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000034e, 5'd16, 27'h000000b3, 5'd22, 27'h000003e1, 32'h00000400,
  1'd1,  5'd24, 27'h000001f0, 5'd29, 27'h00000238, 5'd4, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000bb, 5'd29, 27'h00000046, 5'd13, 27'h000000b9, 32'h00000400,
  1'd1,  5'd23, 27'h0000030a, 5'd25, 27'h00000393, 5'd21, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b7, 5'd6, 27'h00000128, 5'd6, 27'h0000017a, 32'h00000400,
  1'd1,  5'd0, 27'h0000010b, 5'd7, 27'h000001c4, 5'd17, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000284, 5'd8, 27'h00000205, 5'd28, 27'h000003ce, 32'h00000400,
  1'd1,  5'd3, 27'h00000005, 5'd18, 27'h00000294, 5'd8, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000369, 5'd18, 27'h000001f6, 5'd18, 27'h000003e3, 32'h00000400,
  1'd1,  5'd4, 27'h0000012f, 5'd19, 27'h00000042, 5'd25, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000037b, 5'd28, 27'h000003f1, 5'd7, 27'h000002e6, 32'h00000400,
  1'd1,  5'd4, 27'h000000b2, 5'd28, 27'h0000029c, 5'd17, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000f7, 5'd30, 27'h0000025b, 5'd27, 27'h00000300, 32'h00000400,
  1'd1,  5'd14, 27'h00000083, 5'd10, 27'h0000008b, 5'd9, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000273, 5'd9, 27'h00000242, 5'd16, 27'h000001eb, 32'h00000400,
  1'd1,  5'd12, 27'h00000378, 5'd10, 27'h000000f6, 5'd29, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000269, 5'd15, 27'h00000227, 5'd7, 27'h0000019d, 32'h00000400,
  1'd1,  5'd12, 27'h000000f7, 5'd20, 27'h00000023, 5'd17, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e7, 5'd19, 27'h0000016f, 5'd29, 27'h000000b8, 32'h00000400,
  1'd1,  5'd12, 27'h0000034d, 5'd28, 27'h00000349, 5'd6, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000223, 5'd27, 27'h00000330, 5'd17, 27'h000002ec, 32'h00000400,
  1'd1,  5'd13, 27'h00000056, 5'd27, 27'h00000369, 5'd29, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000172, 5'd5, 27'h0000011d, 5'd7, 27'h00000202, 32'h00000400,
  1'd1,  5'd24, 27'h000002b2, 5'd9, 27'h0000030f, 5'd16, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000386, 5'd5, 27'h00000108, 5'd30, 27'h000002f0, 32'h00000400,
  1'd1,  5'd22, 27'h00000395, 5'd19, 27'h000003ac, 5'd7, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000201, 5'd18, 27'h0000004a, 5'd20, 27'h0000023e, 32'h00000400,
  1'd1,  5'd23, 27'h00000366, 5'd20, 27'h0000006d, 5'd30, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006d, 5'd26, 27'h0000035f, 5'd5, 27'h00000299, 32'h00000400,
  1'd1,  5'd25, 27'h0000026c, 5'd30, 27'h00000078, 5'd18, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000396, 5'd27, 27'h00000220, 5'd30, 27'h00000360, 32'h00000400,
  1'd1,  5'd5, 27'h0000036c, 5'd3, 27'h0000001c, 5'd7, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000000c, 5'd4, 27'h0000014c, 5'd16, 27'h0000025c, 32'h00000400,
  1'd1,  5'd8, 27'h000002e1, 5'd2, 27'h00000107, 5'd28, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f1, 5'd14, 27'h0000017f, 5'd1, 27'h0000037b, 32'h00000400,
  1'd1,  5'd9, 27'h000002fc, 5'd12, 27'h0000030f, 5'd13, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000383, 5'd12, 27'h00000163, 5'd22, 27'h000003f4, 32'h00000400,
  1'd1,  5'd6, 27'h000001a6, 5'd21, 27'h0000001c, 5'd1, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000314, 5'd25, 27'h00000025, 5'd10, 27'h000001e0, 32'h00000400,
  1'd1,  5'd8, 27'h000002f5, 5'd23, 27'h00000351, 5'd20, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000341, 5'd3, 27'h0000030a, 5'd9, 27'h000000a9, 32'h00000400,
  1'd1,  5'd17, 27'h00000113, 5'd4, 27'h000001a3, 5'd18, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b5, 5'd3, 27'h000001dd, 5'd27, 27'h000001f0, 32'h00000400,
  1'd1,  5'd17, 27'h0000005d, 5'd13, 27'h00000366, 5'd3, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d4, 5'd14, 27'h0000037d, 5'd14, 27'h00000199, 32'h00000400,
  1'd1,  5'd15, 27'h00000201, 5'd14, 27'h000001ae, 5'd24, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c1, 5'd21, 27'h000003c9, 5'd1, 27'h000003f3, 32'h00000400,
  1'd1,  5'd17, 27'h000002e1, 5'd23, 27'h0000027b, 5'd11, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029d, 5'd24, 27'h000000d9, 5'd21, 27'h00000065, 32'h00000400,
  1'd1,  5'd28, 27'h0000035d, 5'd3, 27'h000001f9, 5'd1, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000023d, 5'd0, 27'h000003a6, 5'd13, 27'h00000215, 32'h00000400,
  1'd1,  5'd28, 27'h000000f1, 5'd1, 27'h000002f7, 5'd24, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d1, 5'd13, 27'h00000351, 5'd1, 27'h00000241, 32'h00000400,
  1'd1,  5'd27, 27'h0000028c, 5'd11, 27'h000002d5, 5'd12, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000309, 5'd10, 27'h0000031c, 5'd23, 27'h0000002c, 32'h00000400,
  1'd1,  5'd26, 27'h000000a1, 5'd21, 27'h000002e8, 5'd2, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000008d, 5'd25, 27'h0000034a, 5'd11, 27'h00000127, 32'h00000400,
  1'd1,  5'd30, 27'h00000199, 5'd23, 27'h000003d1, 5'd23, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000220, 5'd1, 27'h000003ef, 5'd2, 27'h0000003f, 32'h00000400,
  1'd1,  5'd5, 27'h00000304, 5'd0, 27'h00000240, 5'd13, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018b, 5'd3, 27'h0000002e, 5'd21, 27'h00000224, 32'h00000400,
  1'd1,  5'd7, 27'h00000354, 5'd15, 27'h00000059, 5'd5, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000330, 5'd10, 27'h000001c2, 5'd20, 27'h000001b8, 32'h00000400,
  1'd1,  5'd6, 27'h0000033f, 5'd14, 27'h000000a4, 5'd26, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002bd, 5'd24, 27'h0000004b, 5'd8, 27'h0000019c, 32'h00000400,
  1'd1,  5'd7, 27'h00000187, 5'd21, 27'h000003ab, 5'd19, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c7, 5'd21, 27'h000003bc, 5'd30, 27'h000001ed, 32'h00000400,
  1'd1,  5'd19, 27'h000002f4, 5'd4, 27'h00000351, 5'd1, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d5, 5'd3, 27'h0000001a, 5'd11, 27'h00000351, 32'h00000400,
  1'd1,  5'd16, 27'h00000231, 5'd2, 27'h00000114, 5'd23, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000264, 5'd15, 27'h000000fd, 5'd7, 27'h00000331, 32'h00000400,
  1'd1,  5'd19, 27'h000000b4, 5'd14, 27'h0000012a, 5'd16, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003fb, 5'd12, 27'h000002c3, 5'd27, 27'h000003a3, 32'h00000400,
  1'd1,  5'd20, 27'h00000071, 5'd23, 27'h000003d9, 5'd7, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000371, 5'd24, 27'h0000016e, 5'd19, 27'h0000007b, 32'h00000400,
  1'd1,  5'd18, 27'h000000db, 5'd23, 27'h000003ac, 5'd27, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000344, 5'd2, 27'h00000033, 5'd7, 27'h00000187, 32'h00000400,
  1'd1,  5'd29, 27'h00000244, 5'd5, 27'h00000015, 5'd20, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001eb, 5'd0, 27'h000000ec, 5'd29, 27'h000003f9, 32'h00000400,
  1'd1,  5'd30, 27'h00000123, 5'd15, 27'h00000124, 5'd8, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000171, 5'd13, 27'h000003f8, 5'd15, 27'h0000026e, 32'h00000400,
  1'd1,  5'd30, 27'h00000112, 5'd12, 27'h00000329, 5'd29, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003fe, 5'd23, 27'h00000118, 5'd7, 27'h000003bd, 32'h00000400,
  1'd1,  5'd25, 27'h000003ee, 5'd23, 27'h00000067, 5'd16, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f1, 5'd25, 27'h00000352, 5'd29, 27'h0000006f, 32'h00000400,
  1'd1,  5'd5, 27'h00000367, 5'd5, 27'h000003cf, 5'd4, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002b2, 5'd6, 27'h000003f0, 5'd13, 27'h00000032, 32'h00000400,
  1'd1,  5'd7, 27'h000000d7, 5'd8, 27'h00000008, 5'd23, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000373, 5'd19, 27'h00000316, 5'd4, 27'h000003d5, 32'h00000400,
  1'd1,  5'd7, 27'h000000c9, 5'd20, 27'h0000019f, 5'd12, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000028e, 5'd18, 27'h00000386, 5'd21, 27'h00000149, 32'h00000400,
  1'd1,  5'd7, 27'h000001ff, 5'd26, 27'h000003d1, 5'd1, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000260, 5'd26, 27'h00000199, 5'd13, 27'h00000224, 32'h00000400,
  1'd1,  5'd7, 27'h000003dc, 5'd27, 27'h00000087, 5'd22, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d7, 5'd8, 27'h000003f1, 5'd3, 27'h00000342, 32'h00000400,
  1'd1,  5'd20, 27'h000001fe, 5'd8, 27'h0000020e, 5'd15, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c5, 5'd6, 27'h0000021c, 5'd23, 27'h000000b9, 32'h00000400,
  1'd1,  5'd16, 27'h00000087, 5'd16, 27'h0000028b, 5'd3, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000394, 5'd17, 27'h000002af, 5'd12, 27'h000002e2, 32'h00000400,
  1'd1,  5'd15, 27'h000002c8, 5'd19, 27'h00000038, 5'd20, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001e7, 5'd26, 27'h000002c3, 5'd0, 27'h000000de, 32'h00000400,
  1'd1,  5'd19, 27'h000000f2, 5'd28, 27'h00000181, 5'd15, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000202, 5'd27, 27'h0000017a, 5'd22, 27'h000002f8, 32'h00000400,
  1'd1,  5'd28, 27'h000000b4, 5'd7, 27'h0000037c, 5'd3, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002b0, 5'd9, 27'h00000231, 5'd12, 27'h00000256, 32'h00000400,
  1'd1,  5'd29, 27'h000002d1, 5'd9, 27'h00000017, 5'd22, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000022d, 5'd20, 27'h000000c5, 5'd3, 27'h00000155, 32'h00000400,
  1'd1,  5'd29, 27'h00000026, 5'd16, 27'h000000e1, 5'd14, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000322, 5'd19, 27'h00000033, 5'd23, 27'h0000000f, 32'h00000400,
  1'd1,  5'd29, 27'h000002f8, 5'd27, 27'h000003fa, 5'd2, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b7, 5'd29, 27'h000000a1, 5'd14, 27'h000000f1, 32'h00000400,
  1'd1,  5'd27, 27'h0000016a, 5'd28, 27'h000002f2, 5'd21, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000085, 5'd7, 27'h000002e7, 5'd8, 27'h0000010b, 32'h00000400,
  1'd1,  5'd8, 27'h000000a0, 5'd6, 27'h00000125, 5'd17, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000223, 5'd9, 27'h0000015c, 5'd26, 27'h00000221, 32'h00000400,
  1'd1,  5'd7, 27'h00000135, 5'd19, 27'h00000161, 5'd8, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003d5, 5'd20, 27'h00000044, 5'd16, 27'h00000341, 32'h00000400,
  1'd1,  5'd9, 27'h00000106, 5'd18, 27'h00000190, 5'd29, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038d, 5'd27, 27'h000001c9, 5'd8, 27'h00000042, 32'h00000400,
  1'd1,  5'd5, 27'h00000234, 5'd30, 27'h00000196, 5'd19, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033c, 5'd27, 27'h0000001e, 5'd29, 27'h00000038, 32'h00000400,
  1'd1,  5'd17, 27'h000003f4, 5'd8, 27'h0000036e, 5'd7, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000017c, 5'd7, 27'h00000316, 5'd19, 27'h0000000e, 32'h00000400,
  1'd1,  5'd20, 27'h0000015d, 5'd6, 27'h000003e1, 5'd28, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000021e, 5'd19, 27'h000000b6, 5'd9, 27'h0000020e, 32'h00000400,
  1'd1,  5'd18, 27'h00000356, 5'd15, 27'h000003da, 5'd17, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000023a, 5'd18, 27'h000002d9, 5'd26, 27'h00000321, 32'h00000400,
  1'd1,  5'd20, 27'h000001aa, 5'd27, 27'h00000395, 5'd5, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000092, 5'd26, 27'h0000020c, 5'd19, 27'h00000142, 32'h00000400,
  1'd1,  5'd17, 27'h00000007, 5'd29, 27'h00000390, 5'd28, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000183, 5'd5, 27'h00000280, 5'd6, 27'h000000f1, 32'h00000400,
  1'd1,  5'd28, 27'h0000004f, 5'd8, 27'h000000c8, 5'd17, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000164, 5'd5, 27'h000001fb, 5'd29, 27'h0000009d, 32'h00000400,
  1'd1,  5'd29, 27'h00000030, 5'd18, 27'h000003b0, 5'd8, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021c, 5'd20, 27'h000001f8, 5'd16, 27'h00000391, 32'h00000400,
  1'd1,  5'd26, 27'h000003a2, 5'd19, 27'h000001e6, 5'd30, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000077, 5'd27, 27'h0000022e, 5'd6, 27'h0000014f, 32'h00000400,
  1'd1,  5'd29, 27'h0000038e, 5'd30, 27'h000001a2, 5'd18, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000027e, 5'd29, 27'h00000153, 5'd27, 27'h0000016b, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000215, 5'd0, 27'h00000313, 5'd2, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003a6, 5'd4, 27'h00000259, 5'd12, 27'h0000015e, 32'h00000400,
  1'd1,  5'd4, 27'h0000002c, 5'd3, 27'h0000024f, 5'd24, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000125, 5'd11, 27'h000003b4, 5'd1, 27'h000002df, 32'h00000400,
  1'd1,  5'd3, 27'h00000265, 5'd10, 27'h000002f1, 5'd10, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026a, 5'd13, 27'h00000202, 5'd21, 27'h00000292, 32'h00000400,
  1'd1,  5'd1, 27'h000003b0, 5'd22, 27'h00000208, 5'd2, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000254, 5'd23, 27'h00000375, 5'd13, 27'h00000169, 32'h00000400,
  1'd1,  5'd3, 27'h000000fe, 5'd22, 27'h0000038d, 5'd21, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c1, 5'd2, 27'h0000010d, 5'd1, 27'h00000153, 32'h00000400,
  1'd1,  5'd13, 27'h00000296, 5'd1, 27'h0000011b, 5'd12, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000002a, 5'd3, 27'h00000002, 5'd23, 27'h00000028, 32'h00000400,
  1'd1,  5'd14, 27'h00000275, 5'd12, 27'h000001a9, 5'd1, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000183, 5'd14, 27'h000000ce, 5'd11, 27'h0000039d, 32'h00000400,
  1'd1,  5'd13, 27'h0000015c, 5'd12, 27'h0000016d, 5'd20, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c8, 5'd23, 27'h000000d7, 5'd0, 27'h00000374, 32'h00000400,
  1'd1,  5'd12, 27'h00000129, 5'd24, 27'h000001ee, 5'd11, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000026d, 5'd23, 27'h000003fa, 5'd23, 27'h00000110, 32'h00000400,
  1'd1,  5'd21, 27'h000000ff, 5'd0, 27'h00000316, 5'd5, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002cf, 5'd3, 27'h00000126, 5'd13, 27'h000002a9, 32'h00000400,
  1'd1,  5'd20, 27'h00000357, 5'd1, 27'h0000006f, 5'd21, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000008, 5'd15, 27'h0000014e, 5'd1, 27'h00000292, 32'h00000400,
  1'd1,  5'd23, 27'h000001fc, 5'd11, 27'h000000fc, 5'd10, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000226, 5'd14, 27'h00000156, 5'd21, 27'h000002c1, 32'h00000400,
  1'd1,  5'd25, 27'h000001a3, 5'd22, 27'h00000022, 5'd0, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000129, 5'd24, 27'h000002e8, 5'd14, 27'h00000065, 32'h00000400,
  1'd1,  5'd23, 27'h000001c6, 5'd24, 27'h00000010, 5'd23, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000219, 5'd2, 27'h00000243, 5'd7, 27'h0000017e, 32'h00000400,
  1'd1,  5'd0, 27'h000001ae, 5'd3, 27'h00000267, 5'd16, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000232, 5'd0, 27'h0000038b, 5'd27, 27'h00000008, 32'h00000400,
  1'd1,  5'd0, 27'h0000038d, 5'd14, 27'h0000008f, 5'd6, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039a, 5'd15, 27'h000001b9, 5'd17, 27'h000000de, 32'h00000400,
  1'd1,  5'd5, 27'h0000008f, 5'd14, 27'h0000013a, 5'd28, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002c1, 5'd23, 27'h000002a5, 5'd8, 27'h00000368, 32'h00000400,
  1'd1,  5'd2, 27'h000001d3, 5'd24, 27'h000001a9, 5'd17, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000003b, 5'd22, 27'h000001c3, 5'd29, 27'h000002b6, 32'h00000400,
  1'd1,  5'd13, 27'h000001dd, 5'd0, 27'h00000199, 5'd5, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000237, 5'd3, 27'h00000147, 5'd16, 27'h000001d5, 32'h00000400,
  1'd1,  5'd11, 27'h00000289, 5'd1, 27'h0000025a, 5'd26, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000095, 5'd15, 27'h00000129, 5'd9, 27'h00000266, 32'h00000400,
  1'd1,  5'd12, 27'h000002c5, 5'd13, 27'h0000038c, 5'd17, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000280, 5'd10, 27'h000001dd, 5'd27, 27'h0000016f, 32'h00000400,
  1'd1,  5'd13, 27'h00000068, 5'd21, 27'h00000383, 5'd10, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000202, 5'd23, 27'h000003f7, 5'd18, 27'h00000092, 32'h00000400,
  1'd1,  5'd11, 27'h00000162, 5'd24, 27'h0000027a, 5'd30, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000036, 5'd1, 27'h0000031f, 5'd7, 27'h00000092, 32'h00000400,
  1'd1,  5'd20, 27'h0000036c, 5'd4, 27'h00000307, 5'd17, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000001a, 5'd3, 27'h00000388, 5'd27, 27'h0000039b, 32'h00000400,
  1'd1,  5'd21, 27'h0000000a, 5'd10, 27'h00000262, 5'd5, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000014a, 5'd12, 27'h000003c3, 5'd19, 27'h000002c1, 32'h00000400,
  1'd1,  5'd21, 27'h0000023d, 5'd10, 27'h00000236, 5'd30, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000322, 5'd24, 27'h000000cc, 5'd6, 27'h00000094, 32'h00000400,
  1'd1,  5'd21, 27'h000001a7, 5'd25, 27'h0000007d, 5'd19, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000108, 5'd24, 27'h000003d5, 5'd29, 27'h00000139, 32'h00000400,
  1'd1,  5'd4, 27'h000000af, 5'd7, 27'h000002f8, 5'd3, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000189, 5'd7, 27'h00000334, 5'd13, 27'h00000361, 32'h00000400,
  1'd1,  5'd2, 27'h0000021e, 5'd9, 27'h0000035b, 5'd24, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a1, 5'd17, 27'h000002e9, 5'd4, 27'h0000030e, 32'h00000400,
  1'd1,  5'd4, 27'h00000349, 5'd19, 27'h00000383, 5'd10, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002c1, 5'd16, 27'h000000c2, 5'd20, 27'h000002af, 32'h00000400,
  1'd1,  5'd1, 27'h00000221, 5'd30, 27'h00000331, 5'd1, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002eb, 5'd26, 27'h000001c3, 5'd11, 27'h00000302, 32'h00000400,
  1'd1,  5'd5, 27'h00000024, 5'd26, 27'h0000021f, 5'd25, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000d3, 5'd6, 27'h000001dd, 5'd2, 27'h00000019, 32'h00000400,
  1'd1,  5'd12, 27'h0000034d, 5'd9, 27'h000000e0, 5'd14, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000374, 5'd6, 27'h0000007e, 5'd23, 27'h000000e8, 32'h00000400,
  1'd1,  5'd15, 27'h000001c4, 5'd15, 27'h000002c0, 5'd4, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000026, 5'd19, 27'h00000011, 5'd14, 27'h00000157, 32'h00000400,
  1'd1,  5'd12, 27'h00000359, 5'd19, 27'h0000032d, 5'd24, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000229, 5'd28, 27'h000001fd, 5'd0, 27'h000000a8, 32'h00000400,
  1'd1,  5'd12, 27'h00000146, 5'd27, 27'h000003e2, 5'd13, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000243, 5'd27, 27'h0000031d, 5'd21, 27'h00000058, 32'h00000400,
  1'd1,  5'd20, 27'h000003ca, 5'd8, 27'h00000395, 5'd0, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000027c, 5'd7, 27'h000000b3, 5'd10, 27'h00000284, 32'h00000400,
  1'd1,  5'd22, 27'h000001c6, 5'd9, 27'h0000004b, 5'd22, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000141, 5'd20, 27'h00000198, 5'd0, 27'h00000226, 32'h00000400,
  1'd1,  5'd25, 27'h0000006f, 5'd19, 27'h00000131, 5'd15, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000328, 5'd18, 27'h00000132, 5'd21, 27'h0000025c, 32'h00000400,
  1'd1,  5'd25, 27'h000001ce, 5'd29, 27'h000000f9, 5'd0, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000083, 5'd26, 27'h00000134, 5'd14, 27'h0000015f, 32'h00000400,
  1'd1,  5'd25, 27'h00000135, 5'd29, 27'h000001c6, 5'd22, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001fa, 5'd9, 27'h00000310, 5'd9, 27'h0000027d, 32'h00000400,
  1'd1,  5'd0, 27'h00000202, 5'd9, 27'h000003f8, 5'd18, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f2, 5'd5, 27'h000001c8, 5'd28, 27'h000002af, 32'h00000400,
  1'd1,  5'd0, 27'h0000010c, 5'd17, 27'h00000375, 5'd7, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ac, 5'd16, 27'h0000004f, 5'd20, 27'h00000124, 32'h00000400,
  1'd1,  5'd2, 27'h00000355, 5'd15, 27'h000002be, 5'd30, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a8, 5'd27, 27'h00000375, 5'd8, 27'h00000399, 32'h00000400,
  1'd1,  5'd4, 27'h000002f7, 5'd29, 27'h00000070, 5'd17, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b3, 5'd26, 27'h00000162, 5'd29, 27'h000001d2, 32'h00000400,
  1'd1,  5'd10, 27'h00000345, 5'd9, 27'h000002f4, 5'd7, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c4, 5'd5, 27'h000002e0, 5'd20, 27'h000001ff, 32'h00000400,
  1'd1,  5'd12, 27'h000002f6, 5'd6, 27'h000001d4, 5'd26, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001e2, 5'd16, 27'h00000307, 5'd6, 27'h0000007e, 32'h00000400,
  1'd1,  5'd15, 27'h00000180, 5'd15, 27'h00000235, 5'd17, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c4, 5'd17, 27'h00000373, 5'd30, 27'h000003b2, 32'h00000400,
  1'd1,  5'd13, 27'h0000037b, 5'd27, 27'h000003fc, 5'd7, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000009a, 5'd29, 27'h000003ec, 5'd20, 27'h00000203, 32'h00000400,
  1'd1,  5'd13, 27'h00000317, 5'd25, 27'h000003d1, 5'd28, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000e0, 5'd8, 27'h000003b2, 5'd8, 27'h00000294, 32'h00000400,
  1'd1,  5'd24, 27'h00000133, 5'd9, 27'h000000b9, 5'd19, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000dc, 5'd6, 27'h00000135, 5'd30, 27'h0000024e, 32'h00000400,
  1'd1,  5'd24, 27'h000000d1, 5'd16, 27'h00000082, 5'd6, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000069, 5'd19, 27'h0000015c, 5'd18, 27'h0000020c, 32'h00000400,
  1'd1,  5'd21, 27'h0000038e, 5'd15, 27'h00000241, 5'd25, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000002d, 5'd27, 27'h0000000b, 5'd8, 27'h00000321, 32'h00000400,
  1'd1,  5'd21, 27'h00000284, 5'd26, 27'h00000279, 5'd16, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000315, 5'd30, 27'h00000114, 5'd27, 27'h00000241, 32'h00000400,
  1'd1,  5'd7, 27'h0000034e, 5'd4, 27'h000001d9, 5'd5, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d7, 5'd4, 27'h00000083, 5'd17, 27'h0000009f, 32'h00000400,
  1'd1,  5'd8, 27'h0000003e, 5'd3, 27'h0000029c, 5'd30, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000017f, 5'd11, 27'h000003f7, 5'd1, 27'h00000289, 32'h00000400,
  1'd1,  5'd8, 27'h0000021c, 5'd10, 27'h000003f2, 5'd13, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c0, 5'd14, 27'h000003f4, 5'd21, 27'h0000036a, 32'h00000400,
  1'd1,  5'd8, 27'h00000323, 5'd22, 27'h00000112, 5'd4, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ee, 5'd22, 27'h00000214, 5'd11, 27'h0000002b, 32'h00000400,
  1'd1,  5'd10, 27'h00000154, 5'd24, 27'h000003ca, 5'd23, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000021f, 5'd0, 27'h00000326, 5'd6, 27'h000003d8, 32'h00000400,
  1'd1,  5'd16, 27'h0000024d, 5'd1, 27'h000000f8, 5'd17, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003f2, 5'd2, 27'h00000286, 5'd27, 27'h00000216, 32'h00000400,
  1'd1,  5'd16, 27'h0000010c, 5'd12, 27'h00000351, 5'd1, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b2, 5'd10, 27'h00000283, 5'd10, 27'h00000369, 32'h00000400,
  1'd1,  5'd20, 27'h000000e1, 5'd14, 27'h00000319, 5'd22, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000006, 5'd22, 27'h0000035c, 5'd4, 27'h000001f9, 32'h00000400,
  1'd1,  5'd19, 27'h000002dd, 5'd22, 27'h000001d1, 5'd14, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000033a, 5'd25, 27'h000002f6, 5'd24, 27'h0000011f, 32'h00000400,
  1'd1,  5'd28, 27'h00000050, 5'd1, 27'h00000295, 5'd1, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000236, 5'd2, 27'h0000004b, 5'd13, 27'h00000021, 32'h00000400,
  1'd1,  5'd27, 27'h000003f5, 5'd0, 27'h00000270, 5'd24, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000396, 5'd13, 27'h00000258, 5'd2, 27'h00000052, 32'h00000400,
  1'd1,  5'd30, 27'h00000244, 5'd14, 27'h0000010a, 5'd12, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b0, 5'd11, 27'h000002dc, 5'd22, 27'h00000206, 32'h00000400,
  1'd1,  5'd28, 27'h0000015c, 5'd23, 27'h00000369, 5'd3, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000014f, 5'd21, 27'h000003c7, 5'd12, 27'h0000039e, 32'h00000400,
  1'd1,  5'd26, 27'h00000096, 5'd24, 27'h000003d0, 5'd21, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000192, 5'd2, 27'h00000294, 5'd3, 27'h000003a6, 32'h00000400,
  1'd1,  5'd6, 27'h000001e3, 5'd0, 27'h000001ba, 5'd12, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000070, 5'd0, 27'h00000319, 5'd23, 27'h0000004e, 32'h00000400,
  1'd1,  5'd7, 27'h000001b5, 5'd13, 27'h00000237, 5'd9, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000261, 5'd10, 27'h00000291, 5'd20, 27'h00000116, 32'h00000400,
  1'd1,  5'd8, 27'h00000297, 5'd15, 27'h0000018f, 5'd28, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000127, 5'd23, 27'h00000071, 5'd9, 27'h00000235, 32'h00000400,
  1'd1,  5'd8, 27'h000002d4, 5'd20, 27'h0000035c, 5'd19, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001c3, 5'd24, 27'h000001ff, 5'd30, 27'h000002eb, 32'h00000400,
  1'd1,  5'd18, 27'h000002da, 5'd2, 27'h000003ab, 5'd4, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000db, 5'd3, 27'h0000002a, 5'd11, 27'h000002a3, 32'h00000400,
  1'd1,  5'd20, 27'h000000fd, 5'd3, 27'h0000022c, 5'd23, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000007, 5'd14, 27'h00000006, 5'd8, 27'h000001ae, 32'h00000400,
  1'd1,  5'd18, 27'h000002d1, 5'd11, 27'h00000191, 5'd15, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003fe, 5'd14, 27'h00000080, 5'd30, 27'h000002a9, 32'h00000400,
  1'd1,  5'd16, 27'h00000277, 5'd20, 27'h000002dd, 5'd6, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000024c, 5'd22, 27'h0000021a, 5'd19, 27'h00000197, 32'h00000400,
  1'd1,  5'd20, 27'h00000173, 5'd24, 27'h00000249, 5'd28, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003dd, 5'd2, 27'h000002a9, 5'd8, 27'h000003fd, 32'h00000400,
  1'd1,  5'd28, 27'h00000033, 5'd3, 27'h000001dd, 5'd17, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000025f, 5'd0, 27'h000002c7, 5'd26, 27'h000000e6, 32'h00000400,
  1'd1,  5'd26, 27'h0000036e, 5'd11, 27'h00000236, 5'd5, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000051, 5'd14, 27'h0000017d, 5'd17, 27'h000001c6, 32'h00000400,
  1'd1,  5'd29, 27'h00000336, 5'd12, 27'h000002a4, 5'd30, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000251, 5'd25, 27'h00000161, 5'd7, 27'h00000323, 32'h00000400,
  1'd1,  5'd29, 27'h000001a3, 5'd25, 27'h000000b9, 5'd18, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c0, 5'd22, 27'h000001a1, 5'd29, 27'h0000032b, 32'h00000400,
  1'd1,  5'd9, 27'h00000145, 5'd7, 27'h0000019b, 5'd3, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000131, 5'd8, 27'h000002fb, 5'd10, 27'h00000184, 32'h00000400,
  1'd1,  5'd8, 27'h00000102, 5'd8, 27'h000003d4, 5'd20, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003f3, 5'd16, 27'h000001e6, 5'd0, 27'h0000032a, 32'h00000400,
  1'd1,  5'd7, 27'h00000298, 5'd16, 27'h0000012b, 5'd10, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e0, 5'd17, 27'h000001ed, 5'd22, 27'h0000029a, 32'h00000400,
  1'd1,  5'd7, 27'h00000056, 5'd27, 27'h00000323, 5'd1, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c9, 5'd30, 27'h0000024e, 5'd11, 27'h00000027, 32'h00000400,
  1'd1,  5'd6, 27'h00000194, 5'd30, 27'h00000183, 5'd23, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000380, 5'd8, 27'h0000010f, 5'd0, 27'h00000142, 32'h00000400,
  1'd1,  5'd16, 27'h0000009c, 5'd5, 27'h000002b2, 5'd11, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002eb, 5'd8, 27'h000003c3, 5'd23, 27'h000002dd, 32'h00000400,
  1'd1,  5'd15, 27'h00000272, 5'd18, 27'h00000002, 5'd4, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000235, 5'd19, 27'h00000206, 5'd11, 27'h0000005d, 32'h00000400,
  1'd1,  5'd19, 27'h00000016, 5'd20, 27'h0000021a, 5'd25, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000023, 5'd30, 27'h0000008f, 5'd1, 27'h0000017e, 32'h00000400,
  1'd1,  5'd19, 27'h00000201, 5'd26, 27'h00000141, 5'd15, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000244, 5'd27, 27'h000002d6, 5'd21, 27'h0000002a, 32'h00000400,
  1'd1,  5'd28, 27'h000002dd, 5'd6, 27'h0000017e, 5'd4, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000df, 5'd9, 27'h000003a8, 5'd15, 27'h000001ce, 32'h00000400,
  1'd1,  5'd26, 27'h00000187, 5'd7, 27'h000002b1, 5'd23, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000222, 5'd17, 27'h000001e3, 5'd3, 27'h00000324, 32'h00000400,
  1'd1,  5'd28, 27'h000001ab, 5'd18, 27'h0000001b, 5'd12, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000089, 5'd18, 27'h000003f4, 5'd22, 27'h00000153, 32'h00000400,
  1'd1,  5'd26, 27'h000000bd, 5'd28, 27'h000002b9, 5'd1, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000014f, 5'd28, 27'h00000094, 5'd12, 27'h0000036b, 32'h00000400,
  1'd1,  5'd25, 27'h0000035e, 5'd28, 27'h00000320, 5'd24, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000a6, 5'd5, 27'h00000278, 5'd7, 27'h000002a2, 32'h00000400,
  1'd1,  5'd7, 27'h000003a8, 5'd9, 27'h0000001b, 5'd15, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000056, 5'd9, 27'h00000245, 5'd29, 27'h000003b9, 32'h00000400,
  1'd1,  5'd8, 27'h000000f8, 5'd19, 27'h000002d1, 5'd7, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000022b, 5'd19, 27'h0000026a, 5'd16, 27'h00000126, 32'h00000400,
  1'd1,  5'd8, 27'h0000013e, 5'd17, 27'h000001d4, 5'd29, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000f7, 5'd26, 27'h0000028a, 5'd5, 27'h00000306, 32'h00000400,
  1'd1,  5'd5, 27'h000003f3, 5'd28, 27'h00000356, 5'd19, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000004f, 5'd29, 27'h000001bb, 5'd29, 27'h00000019, 32'h00000400,
  1'd1,  5'd19, 27'h00000061, 5'd8, 27'h00000254, 5'd7, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003b4, 5'd5, 27'h000002d3, 5'd16, 27'h000001a4, 32'h00000400,
  1'd1,  5'd16, 27'h0000036e, 5'd9, 27'h000000eb, 5'd28, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f7, 5'd19, 27'h00000302, 5'd7, 27'h00000369, 32'h00000400,
  1'd1,  5'd16, 27'h0000039c, 5'd18, 27'h000000e2, 5'd19, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000234, 5'd15, 27'h00000205, 5'd28, 27'h000002fd, 32'h00000400,
  1'd1,  5'd18, 27'h00000249, 5'd26, 27'h00000034, 5'd8, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002d3, 5'd29, 27'h00000099, 5'd17, 27'h0000004d, 32'h00000400,
  1'd1,  5'd20, 27'h00000286, 5'd30, 27'h000003c0, 5'd28, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000031d, 5'd6, 27'h0000019d, 5'd6, 27'h00000351, 32'h00000400,
  1'd1,  5'd27, 27'h0000000a, 5'd8, 27'h00000050, 5'd16, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038b, 5'd9, 27'h00000150, 5'd30, 27'h000002a9, 32'h00000400,
  1'd1,  5'd30, 27'h00000339, 5'd17, 27'h000003e3, 5'd8, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000006f, 5'd16, 27'h0000005f, 5'd19, 27'h000001fb, 32'h00000400,
  1'd1,  5'd27, 27'h000002a2, 5'd16, 27'h00000252, 5'd28, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034d, 5'd30, 27'h0000038b, 5'd9, 27'h000001b0, 32'h00000400,
  1'd1,  5'd28, 27'h0000012c, 5'd28, 27'h00000059, 5'd18, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003a5, 5'd26, 27'h0000017e, 5'd28, 27'h00000195, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000003c8, 5'd0, 27'h000000af, 5'd3, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000138, 5'd2, 27'h000002b1, 5'd10, 27'h000003a6, 32'h00000400,
  1'd1,  5'd4, 27'h00000220, 5'd3, 27'h00000072, 5'd23, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000272, 5'd12, 27'h000000eb, 5'd2, 27'h0000037e, 32'h00000400,
  1'd1,  5'd4, 27'h00000024, 5'd11, 27'h000000b3, 5'd12, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000b4, 5'd12, 27'h00000363, 5'd25, 27'h0000005c, 32'h00000400,
  1'd1,  5'd3, 27'h000000ef, 5'd24, 27'h00000367, 5'd0, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000341, 5'd23, 27'h00000009, 5'd11, 27'h0000017a, 32'h00000400,
  1'd1,  5'd2, 27'h0000015a, 5'd22, 27'h000000ed, 5'd24, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035c, 5'd4, 27'h000002b2, 5'd0, 27'h00000133, 32'h00000400,
  1'd1,  5'd12, 27'h00000025, 5'd4, 27'h000001e8, 5'd12, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002d2, 5'd0, 27'h000001cb, 5'd22, 27'h00000056, 32'h00000400,
  1'd1,  5'd12, 27'h0000034d, 5'd10, 27'h0000035d, 5'd4, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000181, 5'd13, 27'h00000188, 5'd12, 27'h000002e8, 32'h00000400,
  1'd1,  5'd13, 27'h000003b6, 5'd12, 27'h00000130, 5'd21, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a7, 5'd24, 27'h000001df, 5'd4, 27'h0000028d, 32'h00000400,
  1'd1,  5'd14, 27'h00000050, 5'd24, 27'h000000b6, 5'd14, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000042, 5'd22, 27'h0000005f, 5'd25, 27'h00000268, 32'h00000400,
  1'd1,  5'd23, 27'h00000284, 5'd2, 27'h000003c4, 5'd1, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fb, 5'd2, 27'h000000d5, 5'd12, 27'h000003fa, 32'h00000400,
  1'd1,  5'd25, 27'h00000280, 5'd2, 27'h000002df, 5'd21, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000274, 5'd12, 27'h0000013c, 5'd2, 27'h00000375, 32'h00000400,
  1'd1,  5'd25, 27'h000000e8, 5'd13, 27'h00000075, 5'd11, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000263, 5'd12, 27'h000002a8, 5'd22, 27'h000001e5, 32'h00000400,
  1'd1,  5'd23, 27'h000001c3, 5'd24, 27'h000001fc, 5'd4, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003f4, 5'd23, 27'h00000342, 5'd11, 27'h0000001a, 32'h00000400,
  1'd1,  5'd23, 27'h00000217, 5'd23, 27'h000003eb, 5'd21, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000387, 5'd2, 27'h000001c8, 5'd9, 27'h0000025c, 32'h00000400,
  1'd1,  5'd0, 27'h000000e8, 5'd0, 27'h00000014, 5'd19, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000303, 5'd3, 27'h0000015f, 5'd30, 27'h000000c2, 32'h00000400,
  1'd1,  5'd3, 27'h00000059, 5'd15, 27'h00000010, 5'd6, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000077, 5'd11, 27'h00000166, 5'd19, 27'h000002d7, 32'h00000400,
  1'd1,  5'd4, 27'h0000036f, 5'd12, 27'h00000156, 5'd26, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000021f, 5'd24, 27'h000000fc, 5'd5, 27'h000001bc, 32'h00000400,
  1'd1,  5'd1, 27'h000003a7, 5'd23, 27'h00000154, 5'd18, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000085, 5'd23, 27'h0000028d, 5'd27, 27'h000002f3, 32'h00000400,
  1'd1,  5'd10, 27'h000003a4, 5'd1, 27'h0000009e, 5'd6, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000a7, 5'd0, 27'h000003e4, 5'd19, 27'h000002f2, 32'h00000400,
  1'd1,  5'd11, 27'h00000244, 5'd3, 27'h00000088, 5'd29, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029f, 5'd11, 27'h0000015b, 5'd7, 27'h0000027c, 32'h00000400,
  1'd1,  5'd13, 27'h0000033d, 5'd13, 27'h0000029a, 5'd17, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000165, 5'd13, 27'h00000179, 5'd29, 27'h000000f8, 32'h00000400,
  1'd1,  5'd13, 27'h00000126, 5'd24, 27'h000003e6, 5'd10, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031a, 5'd23, 27'h0000033f, 5'd15, 27'h00000261, 32'h00000400,
  1'd1,  5'd10, 27'h000003df, 5'd22, 27'h0000007f, 5'd29, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032c, 5'd1, 27'h00000130, 5'd7, 27'h00000087, 32'h00000400,
  1'd1,  5'd23, 27'h00000092, 5'd4, 27'h00000259, 5'd15, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c8, 5'd0, 27'h00000261, 5'd27, 27'h00000352, 32'h00000400,
  1'd1,  5'd20, 27'h000003f8, 5'd12, 27'h000003dc, 5'd6, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000201, 5'd10, 27'h000002d6, 5'd15, 27'h000002d8, 32'h00000400,
  1'd1,  5'd23, 27'h00000378, 5'd13, 27'h000000ec, 5'd29, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000190, 5'd23, 27'h00000270, 5'd6, 27'h00000160, 32'h00000400,
  1'd1,  5'd23, 27'h0000033b, 5'd22, 27'h0000034f, 5'd18, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000009, 5'd23, 27'h000003d6, 5'd28, 27'h000003c2, 32'h00000400,
  1'd1,  5'd2, 27'h0000004c, 5'd8, 27'h000001a4, 5'd4, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000018a, 5'd8, 27'h0000038f, 5'd12, 27'h000002b6, 32'h00000400,
  1'd1,  5'd0, 27'h00000104, 5'd7, 27'h000002b9, 5'd24, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f4, 5'd17, 27'h00000282, 5'd1, 27'h00000228, 32'h00000400,
  1'd1,  5'd3, 27'h000002ef, 5'd18, 27'h000003d9, 5'd14, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c7, 5'd18, 27'h0000008e, 5'd22, 27'h000002b0, 32'h00000400,
  1'd1,  5'd2, 27'h000003fc, 5'd30, 27'h0000019a, 5'd3, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c3, 5'd30, 27'h000002b0, 5'd12, 27'h00000325, 32'h00000400,
  1'd1,  5'd4, 27'h0000031a, 5'd30, 27'h00000209, 5'd23, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b9, 5'd5, 27'h00000361, 5'd0, 27'h0000024b, 32'h00000400,
  1'd1,  5'd15, 27'h00000021, 5'd8, 27'h000001a8, 5'd11, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ea, 5'd7, 27'h000003c8, 5'd20, 27'h00000325, 32'h00000400,
  1'd1,  5'd13, 27'h00000303, 5'd19, 27'h000002b9, 5'd1, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e2, 5'd15, 27'h000002fc, 5'd14, 27'h000001a2, 32'h00000400,
  1'd1,  5'd15, 27'h000001cc, 5'd15, 27'h000003a3, 5'd22, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000032e, 5'd29, 27'h000000bb, 5'd2, 27'h000003b9, 32'h00000400,
  1'd1,  5'd10, 27'h000003ae, 5'd30, 27'h000001ee, 5'd11, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c4, 5'd28, 27'h000003f4, 5'd25, 27'h00000285, 32'h00000400,
  1'd1,  5'd21, 27'h00000150, 5'd8, 27'h00000140, 5'd1, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000219, 5'd9, 27'h00000146, 5'd10, 27'h000002e6, 32'h00000400,
  1'd1,  5'd23, 27'h00000373, 5'd8, 27'h00000298, 5'd25, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000000e, 5'd19, 27'h00000388, 5'd2, 27'h000002c1, 32'h00000400,
  1'd1,  5'd22, 27'h00000164, 5'd15, 27'h0000025c, 5'd14, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ce, 5'd19, 27'h00000359, 5'd25, 27'h00000114, 32'h00000400,
  1'd1,  5'd21, 27'h000003c3, 5'd28, 27'h00000299, 5'd1, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000116, 5'd26, 27'h00000156, 5'd10, 27'h0000032e, 32'h00000400,
  1'd1,  5'd25, 27'h00000268, 5'd26, 27'h000001e3, 5'd23, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000021e, 5'd9, 27'h000003cd, 5'd9, 27'h000002e0, 32'h00000400,
  1'd1,  5'd2, 27'h00000079, 5'd6, 27'h00000038, 5'd18, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017a, 5'd9, 27'h00000048, 5'd29, 27'h000003fb, 32'h00000400,
  1'd1,  5'd4, 27'h000001ff, 5'd19, 27'h00000178, 5'd8, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000349, 5'd16, 27'h00000246, 5'd16, 27'h000002f0, 32'h00000400,
  1'd1,  5'd3, 27'h0000004a, 5'd16, 27'h000002c1, 5'd27, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000176, 5'd29, 27'h0000024b, 5'd5, 27'h000001ab, 32'h00000400,
  1'd1,  5'd4, 27'h00000140, 5'd28, 27'h00000283, 5'd15, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d5, 5'd27, 27'h0000023f, 5'd28, 27'h00000069, 32'h00000400,
  1'd1,  5'd13, 27'h00000103, 5'd6, 27'h000002fb, 5'd8, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008f, 5'd7, 27'h000001bd, 5'd15, 27'h000002e2, 32'h00000400,
  1'd1,  5'd14, 27'h00000227, 5'd9, 27'h0000011d, 5'd25, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000005d, 5'd20, 27'h000001e7, 5'd6, 27'h0000008d, 32'h00000400,
  1'd1,  5'd13, 27'h00000282, 5'd19, 27'h0000032e, 5'd17, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013d, 5'd19, 27'h000001fe, 5'd30, 27'h000003e7, 32'h00000400,
  1'd1,  5'd12, 27'h0000011d, 5'd30, 27'h000001fc, 5'd9, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000212, 5'd26, 27'h000001a8, 5'd19, 27'h00000091, 32'h00000400,
  1'd1,  5'd12, 27'h000003fd, 5'd30, 27'h000000ee, 5'd26, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000285, 5'd6, 27'h00000006, 5'd8, 27'h00000060, 32'h00000400,
  1'd1,  5'd22, 27'h0000028b, 5'd5, 27'h000003b6, 5'd20, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000179, 5'd10, 27'h00000008, 5'd26, 27'h00000364, 32'h00000400,
  1'd1,  5'd24, 27'h0000032e, 5'd15, 27'h000002eb, 5'd9, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e6, 5'd20, 27'h000001fe, 5'd19, 27'h000000c3, 32'h00000400,
  1'd1,  5'd22, 27'h00000335, 5'd19, 27'h000000d5, 5'd30, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000035, 5'd27, 27'h00000237, 5'd9, 27'h000001eb, 32'h00000400,
  1'd1,  5'd23, 27'h000000cc, 5'd27, 27'h00000205, 5'd20, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000223, 5'd28, 27'h00000342, 5'd30, 27'h000001b7, 32'h00000400,
  1'd1,  5'd10, 27'h00000036, 5'd1, 27'h00000044, 5'd9, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002b4, 5'd2, 27'h00000178, 5'd18, 27'h000000b2, 32'h00000400,
  1'd1,  5'd7, 27'h0000002f, 5'd0, 27'h0000015d, 5'd29, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000047, 5'd13, 27'h000001eb, 5'd1, 27'h00000291, 32'h00000400,
  1'd1,  5'd6, 27'h00000253, 5'd10, 27'h000001a3, 5'd13, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000034a, 5'd13, 27'h000003f7, 5'd22, 27'h000003cc, 32'h00000400,
  1'd1,  5'd5, 27'h00000146, 5'd23, 27'h000001c0, 5'd3, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000263, 5'd24, 27'h00000139, 5'd13, 27'h00000119, 32'h00000400,
  1'd1,  5'd5, 27'h00000182, 5'd24, 27'h00000141, 5'd22, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000116, 5'd4, 27'h00000100, 5'd7, 27'h000002c1, 32'h00000400,
  1'd1,  5'd16, 27'h000002b6, 5'd3, 27'h00000285, 5'd17, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003e8, 5'd3, 27'h000000d9, 5'd26, 27'h0000008a, 32'h00000400,
  1'd1,  5'd17, 27'h00000000, 5'd10, 27'h00000182, 5'd0, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000015c, 5'd10, 27'h000001be, 5'd13, 27'h00000308, 32'h00000400,
  1'd1,  5'd16, 27'h0000015c, 5'd11, 27'h000000c8, 5'd22, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000187, 5'd24, 27'h0000025f, 5'd0, 27'h00000122, 32'h00000400,
  1'd1,  5'd16, 27'h000003a7, 5'd24, 27'h000000e7, 5'd11, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ef, 5'd24, 27'h000000bb, 5'd21, 27'h0000012f, 32'h00000400,
  1'd1,  5'd30, 27'h0000035a, 5'd5, 27'h0000006c, 5'd0, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000224, 5'd4, 27'h000003ff, 5'd11, 27'h000003b6, 32'h00000400,
  1'd1,  5'd29, 27'h0000004f, 5'd2, 27'h0000003e, 5'd22, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a9, 5'd14, 27'h000002ff, 5'd0, 27'h000001cd, 32'h00000400,
  1'd1,  5'd28, 27'h00000066, 5'd12, 27'h000000fd, 5'd12, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003dd, 5'd13, 27'h00000012, 5'd22, 27'h00000077, 32'h00000400,
  1'd1,  5'd29, 27'h0000029e, 5'd24, 27'h0000011f, 5'd2, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000101, 5'd23, 27'h000003ab, 5'd10, 27'h00000162, 32'h00000400,
  1'd1,  5'd30, 27'h000002e3, 5'd23, 27'h000000c8, 5'd25, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000346, 5'd1, 27'h00000045, 5'd4, 27'h000000b5, 32'h00000400,
  1'd1,  5'd6, 27'h0000038a, 5'd1, 27'h00000074, 5'd11, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c0, 5'd3, 27'h00000118, 5'd22, 27'h00000202, 32'h00000400,
  1'd1,  5'd6, 27'h0000013c, 5'd14, 27'h00000135, 5'd8, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000110, 5'd14, 27'h00000204, 5'd19, 27'h00000289, 32'h00000400,
  1'd1,  5'd6, 27'h0000021f, 5'd10, 27'h00000288, 5'd28, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001bb, 5'd22, 27'h000001e4, 5'd7, 27'h00000205, 32'h00000400,
  1'd1,  5'd10, 27'h0000000e, 5'd21, 27'h00000084, 5'd19, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000124, 5'd20, 27'h0000030f, 5'd26, 27'h0000005e, 32'h00000400,
  1'd1,  5'd16, 27'h000002b1, 5'd1, 27'h000001b4, 5'd0, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002d5, 5'd0, 27'h000000e7, 5'd13, 27'h000000a6, 32'h00000400,
  1'd1,  5'd16, 27'h000000e5, 5'd3, 27'h000000d3, 5'd21, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000023a, 5'd11, 27'h000001c7, 5'd8, 27'h00000389, 32'h00000400,
  1'd1,  5'd17, 27'h000000ad, 5'd14, 27'h000000db, 5'd20, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000084, 5'd14, 27'h000000c4, 5'd26, 27'h00000047, 32'h00000400,
  1'd1,  5'd16, 27'h000003bf, 5'd25, 27'h00000196, 5'd9, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b0, 5'd21, 27'h00000335, 5'd16, 27'h0000002c, 32'h00000400,
  1'd1,  5'd16, 27'h000001ce, 5'd23, 27'h000002b0, 5'd28, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003bc, 5'd1, 27'h000003f7, 5'd7, 27'h000000e9, 32'h00000400,
  1'd1,  5'd30, 27'h0000013c, 5'd1, 27'h000003af, 5'd18, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001b2, 5'd3, 27'h00000041, 5'd30, 27'h000002f3, 32'h00000400,
  1'd1,  5'd30, 27'h000001bb, 5'd14, 27'h000003a3, 5'd7, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000204, 5'd10, 27'h0000035d, 5'd20, 27'h00000040, 32'h00000400,
  1'd1,  5'd30, 27'h00000367, 5'd14, 27'h00000396, 5'd26, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000119, 5'd21, 27'h00000016, 5'd7, 27'h0000014b, 32'h00000400,
  1'd1,  5'd29, 27'h00000322, 5'd23, 27'h00000246, 5'd16, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000145, 5'd21, 27'h000003f3, 5'd26, 27'h0000008f, 32'h00000400,
  1'd1,  5'd9, 27'h0000006f, 5'd9, 27'h00000160, 5'd3, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000318, 5'd10, 27'h0000001b, 5'd13, 27'h00000190, 32'h00000400,
  1'd1,  5'd7, 27'h00000342, 5'd9, 27'h000000e8, 5'd24, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001b9, 5'd18, 27'h0000006b, 5'd3, 27'h00000233, 32'h00000400,
  1'd1,  5'd5, 27'h000001c2, 5'd16, 27'h00000063, 5'd14, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003a6, 5'd17, 27'h000001ea, 5'd21, 27'h00000349, 32'h00000400,
  1'd1,  5'd9, 27'h00000158, 5'd29, 27'h0000000a, 5'd1, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000376, 5'd29, 27'h000000c0, 5'd15, 27'h000000f9, 32'h00000400,
  1'd1,  5'd6, 27'h0000012e, 5'd30, 27'h0000038a, 5'd20, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b8, 5'd10, 27'h0000002f, 5'd1, 27'h0000030a, 32'h00000400,
  1'd1,  5'd16, 27'h00000188, 5'd8, 27'h0000023b, 5'd13, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000027c, 5'd6, 27'h00000206, 5'd22, 27'h000000ac, 32'h00000400,
  1'd1,  5'd17, 27'h00000206, 5'd16, 27'h000003b9, 5'd1, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000256, 5'd15, 27'h000003dd, 5'd12, 27'h00000383, 32'h00000400,
  1'd1,  5'd16, 27'h000002cc, 5'd17, 27'h0000032e, 5'd24, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000188, 5'd26, 27'h0000012f, 5'd1, 27'h0000039d, 32'h00000400,
  1'd1,  5'd18, 27'h000000ca, 5'd25, 27'h00000360, 5'd12, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000045, 5'd26, 27'h0000024a, 5'd25, 27'h000000fb, 32'h00000400,
  1'd1,  5'd30, 27'h00000353, 5'd8, 27'h00000214, 5'd1, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002fe, 5'd10, 27'h00000035, 5'd11, 27'h000001b5, 32'h00000400,
  1'd1,  5'd29, 27'h00000182, 5'd8, 27'h0000016d, 5'd24, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017f, 5'd18, 27'h0000031a, 5'd0, 27'h0000013f, 32'h00000400,
  1'd1,  5'd29, 27'h00000262, 5'd15, 27'h0000039b, 5'd12, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000032d, 5'd20, 27'h00000027, 5'd21, 27'h00000015, 32'h00000400,
  1'd1,  5'd27, 27'h000002f8, 5'd29, 27'h0000021e, 5'd2, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000020d, 5'd26, 27'h0000027b, 5'd12, 27'h00000107, 32'h00000400,
  1'd1,  5'd28, 27'h000002c7, 5'd27, 27'h0000023b, 5'd21, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000159, 5'd5, 27'h00000182, 5'd9, 27'h00000055, 32'h00000400,
  1'd1,  5'd5, 27'h000002bb, 5'd9, 27'h00000284, 5'd18, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033f, 5'd7, 27'h00000301, 5'd27, 27'h000000ac, 32'h00000400,
  1'd1,  5'd9, 27'h0000022e, 5'd18, 27'h000003b8, 5'd9, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000018d, 5'd17, 27'h000003b8, 5'd17, 27'h000000a6, 32'h00000400,
  1'd1,  5'd7, 27'h00000322, 5'd15, 27'h000002c2, 5'd28, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002da, 5'd30, 27'h000000b8, 5'd9, 27'h00000302, 32'h00000400,
  1'd1,  5'd6, 27'h00000042, 5'd26, 27'h00000191, 5'd19, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002cb, 5'd26, 27'h000000a6, 5'd27, 27'h00000259, 32'h00000400,
  1'd1,  5'd16, 27'h0000033d, 5'd10, 27'h00000081, 5'd8, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000033b, 5'd6, 27'h000003b4, 5'd20, 27'h000000fd, 32'h00000400,
  1'd1,  5'd17, 27'h00000207, 5'd5, 27'h0000033b, 5'd26, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000294, 5'd20, 27'h00000280, 5'd5, 27'h00000316, 32'h00000400,
  1'd1,  5'd16, 27'h000002b6, 5'd17, 27'h000003f4, 5'd15, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002fa, 5'd15, 27'h00000327, 5'd28, 27'h000003e9, 32'h00000400,
  1'd1,  5'd20, 27'h00000173, 5'd27, 27'h0000031e, 5'd8, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a7, 5'd29, 27'h000000d2, 5'd16, 27'h00000142, 32'h00000400,
  1'd1,  5'd20, 27'h00000048, 5'd28, 27'h00000367, 5'd29, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000379, 5'd6, 27'h000003e6, 5'd6, 27'h0000027a, 32'h00000400,
  1'd1,  5'd27, 27'h000001a5, 5'd9, 27'h0000002b, 5'd19, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034e, 5'd9, 27'h00000036, 5'd26, 27'h0000030c, 32'h00000400,
  1'd1,  5'd26, 27'h000003df, 5'd17, 27'h000000d1, 5'd10, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c0, 5'd20, 27'h000001a4, 5'd19, 27'h00000192, 32'h00000400,
  1'd1,  5'd26, 27'h000000c5, 5'd17, 27'h00000020, 5'd28, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000072, 5'd28, 27'h000001fd, 5'd8, 27'h00000132, 32'h00000400,
  1'd1,  5'd27, 27'h0000001e, 5'd27, 27'h0000008b, 5'd20, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000139, 5'd30, 27'h000001ea, 5'd28, 27'h000000c5, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000025d, 5'd3, 27'h000000ba, 5'd0, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000039e, 5'd4, 27'h000002f0, 5'd11, 27'h00000061, 32'h00000400,
  1'd1,  5'd2, 27'h00000007, 5'd4, 27'h00000100, 5'd20, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000368, 5'd14, 27'h000000ab, 5'd1, 27'h00000367, 32'h00000400,
  1'd1,  5'd3, 27'h0000029e, 5'd10, 27'h000003b2, 5'd11, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000024e, 5'd11, 27'h000000d3, 5'd21, 27'h0000016d, 32'h00000400,
  1'd1,  5'd1, 27'h0000002f, 5'd23, 27'h000001b3, 5'd1, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012a, 5'd24, 27'h00000036, 5'd12, 27'h00000130, 32'h00000400,
  1'd1,  5'd3, 27'h0000016a, 5'd23, 27'h000003c8, 5'd21, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d9, 5'd4, 27'h000002ce, 5'd1, 27'h00000123, 32'h00000400,
  1'd1,  5'd13, 27'h0000003f, 5'd1, 27'h000000eb, 5'd12, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000132, 5'd2, 27'h000001b7, 5'd24, 27'h000003a1, 32'h00000400,
  1'd1,  5'd11, 27'h000003f5, 5'd14, 27'h000003ef, 5'd0, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000287, 5'd14, 27'h000002c2, 5'd12, 27'h0000033c, 32'h00000400,
  1'd1,  5'd14, 27'h00000158, 5'd11, 27'h000002c9, 5'd25, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000106, 5'd21, 27'h000001e5, 5'd0, 27'h000000b4, 32'h00000400,
  1'd1,  5'd10, 27'h0000031c, 5'd23, 27'h000003b9, 5'd14, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000032, 5'd23, 27'h000001f4, 5'd23, 27'h0000021c, 32'h00000400,
  1'd1,  5'd22, 27'h000000d4, 5'd2, 27'h000002a1, 5'd0, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000172, 5'd4, 27'h00000241, 5'd13, 27'h00000377, 32'h00000400,
  1'd1,  5'd25, 27'h0000033d, 5'd0, 27'h00000032, 5'd23, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000061, 5'd12, 27'h000002e9, 5'd0, 27'h00000260, 32'h00000400,
  1'd1,  5'd23, 27'h00000305, 5'd11, 27'h00000355, 5'd14, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ff, 5'd12, 27'h00000220, 5'd24, 27'h00000286, 32'h00000400,
  1'd1,  5'd22, 27'h00000103, 5'd22, 27'h000001b1, 5'd0, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000285, 5'd20, 27'h000002eb, 5'd14, 27'h0000035f, 32'h00000400,
  1'd1,  5'd25, 27'h00000240, 5'd24, 27'h00000027, 5'd25, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000146, 5'd2, 27'h000000a8, 5'd8, 27'h00000200, 32'h00000400,
  1'd1,  5'd1, 27'h000000d2, 5'd2, 27'h000001f0, 5'd19, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000317, 5'd2, 27'h000003ba, 5'd30, 27'h0000010f, 32'h00000400,
  1'd1,  5'd0, 27'h000003fb, 5'd13, 27'h00000190, 5'd6, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000395, 5'd14, 27'h00000306, 5'd16, 27'h00000383, 32'h00000400,
  1'd1,  5'd2, 27'h000002c9, 5'd10, 27'h000001d9, 5'd26, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ab, 5'd25, 27'h00000305, 5'd5, 27'h000001c4, 32'h00000400,
  1'd1,  5'd1, 27'h0000019a, 5'd21, 27'h00000047, 5'd17, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012e, 5'd21, 27'h000002bb, 5'd26, 27'h00000280, 32'h00000400,
  1'd1,  5'd15, 27'h000000f9, 5'd2, 27'h00000366, 5'd6, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000033f, 5'd4, 27'h00000240, 5'd16, 27'h0000036f, 32'h00000400,
  1'd1,  5'd11, 27'h00000001, 5'd1, 27'h000003f8, 5'd26, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001de, 5'd11, 27'h000002ba, 5'd5, 27'h00000384, 32'h00000400,
  1'd1,  5'd13, 27'h00000303, 5'd13, 27'h0000036a, 5'd19, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001dd, 5'd14, 27'h000001b9, 5'd28, 27'h0000015d, 32'h00000400,
  1'd1,  5'd10, 27'h000001bf, 5'd23, 27'h0000002e, 5'd7, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000a5, 5'd25, 27'h00000010, 5'd19, 27'h00000286, 32'h00000400,
  1'd1,  5'd11, 27'h0000032d, 5'd24, 27'h0000011f, 5'd26, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ac, 5'd1, 27'h000001b1, 5'd7, 27'h00000312, 32'h00000400,
  1'd1,  5'd25, 27'h0000009c, 5'd4, 27'h00000330, 5'd17, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001fc, 5'd2, 27'h000003a3, 5'd26, 27'h0000034d, 32'h00000400,
  1'd1,  5'd22, 27'h0000016c, 5'd13, 27'h000000e0, 5'd5, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000034f, 5'd13, 27'h0000033b, 5'd17, 27'h00000244, 32'h00000400,
  1'd1,  5'd20, 27'h000003fd, 5'd12, 27'h00000367, 5'd26, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000386, 5'd24, 27'h00000286, 5'd5, 27'h000000d4, 32'h00000400,
  1'd1,  5'd22, 27'h00000354, 5'd22, 27'h000002a6, 5'd16, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000011d, 5'd25, 27'h000000b7, 5'd27, 27'h000003c9, 32'h00000400,
  1'd1,  5'd0, 27'h0000003e, 5'd7, 27'h00000356, 5'd2, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003cb, 5'd8, 27'h00000289, 5'd12, 27'h00000353, 32'h00000400,
  1'd1,  5'd0, 27'h000002b8, 5'd9, 27'h0000012b, 5'd21, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b1, 5'd16, 27'h0000024a, 5'd3, 27'h00000158, 32'h00000400,
  1'd1,  5'd1, 27'h000003cc, 5'd17, 27'h000001a9, 5'd11, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000008d, 5'd16, 27'h0000017e, 5'd21, 27'h0000004b, 32'h00000400,
  1'd1,  5'd2, 27'h0000024c, 5'd27, 27'h00000170, 5'd2, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000085, 5'd30, 27'h000000fd, 5'd10, 27'h0000021c, 32'h00000400,
  1'd1,  5'd2, 27'h0000031c, 5'd27, 27'h00000151, 5'd24, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003bf, 5'd9, 27'h00000127, 5'd2, 27'h0000037d, 32'h00000400,
  1'd1,  5'd13, 27'h000003b0, 5'd5, 27'h00000198, 5'd13, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000193, 5'd7, 27'h000000f6, 5'd21, 27'h00000396, 32'h00000400,
  1'd1,  5'd12, 27'h0000010d, 5'd16, 27'h00000064, 5'd3, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000e8, 5'd17, 27'h000003c4, 5'd14, 27'h000000f5, 32'h00000400,
  1'd1,  5'd14, 27'h000003ce, 5'd17, 27'h000001e6, 5'd21, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003d4, 5'd27, 27'h00000138, 5'd1, 27'h000000b6, 32'h00000400,
  1'd1,  5'd12, 27'h000000d2, 5'd30, 27'h00000396, 5'd15, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002ec, 5'd26, 27'h0000005a, 5'd25, 27'h000002f9, 32'h00000400,
  1'd1,  5'd22, 27'h000002a8, 5'd8, 27'h00000233, 5'd4, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000027c, 5'd6, 27'h000000f9, 5'd14, 27'h00000126, 32'h00000400,
  1'd1,  5'd24, 27'h000000e3, 5'd8, 27'h00000194, 5'd22, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000015c, 5'd20, 27'h000000a4, 5'd3, 27'h000002d6, 32'h00000400,
  1'd1,  5'd22, 27'h000000d8, 5'd15, 27'h000002ba, 5'd12, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000004b, 5'd18, 27'h00000159, 5'd22, 27'h00000395, 32'h00000400,
  1'd1,  5'd23, 27'h00000198, 5'd29, 27'h0000015a, 5'd0, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000008e, 5'd27, 27'h0000020e, 5'd14, 27'h00000375, 32'h00000400,
  1'd1,  5'd23, 27'h000000a0, 5'd26, 27'h00000370, 5'd23, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000026c, 5'd5, 27'h000003f3, 5'd5, 27'h00000390, 32'h00000400,
  1'd1,  5'd4, 27'h000002b0, 5'd8, 27'h0000037e, 5'd17, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000254, 5'd6, 27'h00000081, 5'd29, 27'h00000183, 32'h00000400,
  1'd1,  5'd4, 27'h00000260, 5'd20, 27'h0000024b, 5'd6, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000344, 5'd18, 27'h0000026a, 5'd18, 27'h00000053, 32'h00000400,
  1'd1,  5'd3, 27'h000000b8, 5'd19, 27'h00000373, 5'd26, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000339, 5'd29, 27'h0000036a, 5'd8, 27'h00000066, 32'h00000400,
  1'd1,  5'd0, 27'h000003db, 5'd26, 27'h0000033d, 5'd18, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000184, 5'd28, 27'h00000262, 5'd26, 27'h000002c3, 32'h00000400,
  1'd1,  5'd14, 27'h000003d8, 5'd6, 27'h000001ff, 5'd8, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000037, 5'd8, 27'h0000033a, 5'd16, 27'h000003f1, 32'h00000400,
  1'd1,  5'd13, 27'h00000168, 5'd5, 27'h00000368, 5'd26, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000292, 5'd17, 27'h0000038d, 5'd10, 27'h000000a1, 32'h00000400,
  1'd1,  5'd11, 27'h00000080, 5'd17, 27'h0000030e, 5'd17, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000015f, 5'd16, 27'h00000340, 5'd30, 27'h00000321, 32'h00000400,
  1'd1,  5'd13, 27'h000001f9, 5'd29, 27'h00000068, 5'd7, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001cd, 5'd29, 27'h00000399, 5'd17, 27'h00000226, 32'h00000400,
  1'd1,  5'd11, 27'h00000152, 5'd28, 27'h00000211, 5'd27, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002eb, 5'd6, 27'h00000400, 5'd9, 27'h000001b0, 32'h00000400,
  1'd1,  5'd22, 27'h00000390, 5'd8, 27'h00000376, 5'd19, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000af, 5'd6, 27'h000001ad, 5'd30, 27'h00000085, 32'h00000400,
  1'd1,  5'd25, 27'h000001e1, 5'd17, 27'h000001eb, 5'd9, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003e8, 5'd18, 27'h0000020b, 5'd19, 27'h000003b2, 32'h00000400,
  1'd1,  5'd24, 27'h0000001d, 5'd15, 27'h00000225, 5'd30, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000314, 5'd29, 27'h000003a4, 5'd7, 27'h000003d3, 32'h00000400,
  1'd1,  5'd22, 27'h00000218, 5'd28, 27'h00000059, 5'd15, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000188, 5'd29, 27'h000002cf, 5'd28, 27'h0000015b, 32'h00000400,
  1'd1,  5'd9, 27'h0000009b, 5'd0, 27'h00000241, 5'd6, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001f9, 5'd2, 27'h00000243, 5'd17, 27'h00000389, 32'h00000400,
  1'd1,  5'd8, 27'h000001b8, 5'd1, 27'h0000013c, 5'd26, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000010f, 5'd10, 27'h00000346, 5'd4, 27'h000002b2, 32'h00000400,
  1'd1,  5'd5, 27'h0000025d, 5'd11, 27'h000000de, 5'd12, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000194, 5'd15, 27'h00000150, 5'd22, 27'h00000352, 32'h00000400,
  1'd1,  5'd8, 27'h000001b1, 5'd25, 27'h000000da, 5'd4, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000021e, 5'd25, 27'h00000303, 5'd13, 27'h00000107, 32'h00000400,
  1'd1,  5'd10, 27'h00000102, 5'd23, 27'h000002f8, 5'd24, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002cc, 5'd2, 27'h0000012a, 5'd5, 27'h000003a3, 32'h00000400,
  1'd1,  5'd20, 27'h00000053, 5'd5, 27'h00000088, 5'd19, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000161, 5'd3, 27'h000001c9, 5'd27, 27'h0000012e, 32'h00000400,
  1'd1,  5'd17, 27'h000001fd, 5'd11, 27'h000001ba, 5'd2, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000023e, 5'd10, 27'h0000036a, 5'd15, 27'h00000031, 32'h00000400,
  1'd1,  5'd19, 27'h00000175, 5'd11, 27'h000002d8, 5'd22, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b7, 5'd22, 27'h000001a9, 5'd4, 27'h0000014a, 32'h00000400,
  1'd1,  5'd17, 27'h0000007a, 5'd23, 27'h00000191, 5'd10, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031f, 5'd21, 27'h00000228, 5'd24, 27'h00000253, 32'h00000400,
  1'd1,  5'd26, 27'h000000b1, 5'd4, 27'h0000015e, 5'd1, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000034, 5'd0, 27'h0000030a, 5'd12, 27'h00000112, 32'h00000400,
  1'd1,  5'd27, 27'h000002cb, 5'd3, 27'h00000237, 5'd25, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000000d, 5'd13, 27'h00000017, 5'd2, 27'h00000206, 32'h00000400,
  1'd1,  5'd30, 27'h00000103, 5'd12, 27'h000000d9, 5'd12, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c8, 5'd11, 27'h00000078, 5'd23, 27'h00000062, 32'h00000400,
  1'd1,  5'd30, 27'h000001a1, 5'd23, 27'h00000378, 5'd2, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000039b, 5'd21, 27'h00000305, 5'd14, 27'h0000028e, 32'h00000400,
  1'd1,  5'd27, 27'h0000010c, 5'd25, 27'h00000161, 5'd23, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000289, 5'd1, 27'h000000fc, 5'd3, 27'h00000272, 32'h00000400,
  1'd1,  5'd5, 27'h00000191, 5'd3, 27'h00000223, 5'd11, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001e5, 5'd4, 27'h00000102, 5'd21, 27'h00000091, 32'h00000400,
  1'd1,  5'd8, 27'h00000173, 5'd10, 27'h00000227, 5'd7, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000055, 5'd11, 27'h00000019, 5'd17, 27'h0000002d, 32'h00000400,
  1'd1,  5'd5, 27'h00000115, 5'd15, 27'h00000078, 5'd27, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d6, 5'd24, 27'h000000ff, 5'd7, 27'h00000233, 32'h00000400,
  1'd1,  5'd9, 27'h000001e5, 5'd21, 27'h00000399, 5'd16, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000023d, 5'd23, 27'h00000295, 5'd28, 27'h0000022e, 32'h00000400,
  1'd1,  5'd15, 27'h000003dd, 5'd2, 27'h000003c1, 5'd2, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000167, 5'd3, 27'h00000197, 5'd14, 27'h000003d6, 32'h00000400,
  1'd1,  5'd19, 27'h000000b1, 5'd0, 27'h00000328, 5'd24, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000003, 5'd13, 27'h0000003b, 5'd5, 27'h000001c8, 32'h00000400,
  1'd1,  5'd15, 27'h000002d6, 5'd11, 27'h000000b9, 5'd17, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000028c, 5'd12, 27'h00000074, 5'd30, 27'h00000222, 32'h00000400,
  1'd1,  5'd19, 27'h0000004c, 5'd20, 27'h000002c7, 5'd9, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002bc, 5'd21, 27'h000003d2, 5'd20, 27'h000001d2, 32'h00000400,
  1'd1,  5'd20, 27'h00000240, 5'd22, 27'h000003f1, 5'd29, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012e, 5'd2, 27'h0000006e, 5'd6, 27'h000000ec, 32'h00000400,
  1'd1,  5'd30, 27'h00000186, 5'd0, 27'h000003d0, 5'd18, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000159, 5'd4, 27'h000002c0, 5'd30, 27'h000000a3, 32'h00000400,
  1'd1,  5'd27, 27'h00000218, 5'd11, 27'h00000061, 5'd7, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000295, 5'd14, 27'h00000324, 5'd18, 27'h0000032b, 32'h00000400,
  1'd1,  5'd29, 27'h000001cd, 5'd15, 27'h0000006b, 5'd26, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000004a, 5'd21, 27'h000001fc, 5'd9, 27'h000001b8, 32'h00000400,
  1'd1,  5'd29, 27'h0000004a, 5'd21, 27'h000003da, 5'd15, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003fd, 5'd25, 27'h0000018f, 5'd28, 27'h00000378, 32'h00000400,
  1'd1,  5'd7, 27'h000000e0, 5'd8, 27'h00000111, 5'd4, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000221, 5'd7, 27'h000000d3, 5'd14, 27'h000001a9, 32'h00000400,
  1'd1,  5'd8, 27'h00000194, 5'd8, 27'h000000a4, 5'd22, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c3, 5'd15, 27'h00000313, 5'd1, 27'h000002eb, 32'h00000400,
  1'd1,  5'd6, 27'h0000037f, 5'd18, 27'h00000123, 5'd14, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011c, 5'd18, 27'h00000189, 5'd24, 27'h0000039a, 32'h00000400,
  1'd1,  5'd6, 27'h0000029a, 5'd30, 27'h0000036c, 5'd1, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000210, 5'd27, 27'h000000c2, 5'd10, 27'h000003e2, 32'h00000400,
  1'd1,  5'd7, 27'h0000021a, 5'd29, 27'h0000016a, 5'd21, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000302, 5'd10, 27'h000000fa, 5'd0, 27'h0000023e, 32'h00000400,
  1'd1,  5'd15, 27'h000002a1, 5'd9, 27'h00000119, 5'd12, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000388, 5'd8, 27'h00000221, 5'd25, 27'h00000236, 32'h00000400,
  1'd1,  5'd19, 27'h000003fd, 5'd19, 27'h00000347, 5'd4, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000365, 5'd18, 27'h00000052, 5'd14, 27'h000002b0, 32'h00000400,
  1'd1,  5'd17, 27'h00000060, 5'd18, 27'h00000261, 5'd25, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000068, 5'd26, 27'h0000021a, 5'd0, 27'h00000134, 32'h00000400,
  1'd1,  5'd18, 27'h000000ff, 5'd28, 27'h000000fc, 5'd13, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000305, 5'd26, 27'h000000fe, 5'd22, 27'h000001f9, 32'h00000400,
  1'd1,  5'd28, 27'h000003c4, 5'd5, 27'h00000248, 5'd4, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000011d, 5'd10, 27'h00000056, 5'd13, 27'h000003cb, 32'h00000400,
  1'd1,  5'd26, 27'h000000c9, 5'd6, 27'h0000019c, 5'd21, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002fa, 5'd19, 27'h0000027e, 5'd3, 27'h00000351, 32'h00000400,
  1'd1,  5'd27, 27'h000001a1, 5'd17, 27'h00000273, 5'd14, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000225, 5'd18, 27'h000002f5, 5'd25, 27'h000000bd, 32'h00000400,
  1'd1,  5'd29, 27'h00000163, 5'd27, 27'h00000165, 5'd0, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001f1, 5'd25, 27'h000003b6, 5'd11, 27'h000002be, 32'h00000400,
  1'd1,  5'd27, 27'h00000166, 5'd27, 27'h00000306, 5'd20, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000122, 5'd6, 27'h00000097, 5'd6, 27'h00000064, 32'h00000400,
  1'd1,  5'd6, 27'h0000015a, 5'd8, 27'h0000025d, 5'd20, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000234, 5'd7, 27'h0000026c, 5'd25, 27'h000003e4, 32'h00000400,
  1'd1,  5'd10, 27'h0000007b, 5'd17, 27'h0000039b, 5'd8, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000243, 5'd17, 27'h0000038e, 5'd16, 27'h000002ca, 32'h00000400,
  1'd1,  5'd6, 27'h00000226, 5'd16, 27'h000000de, 5'd27, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001dc, 5'd27, 27'h00000218, 5'd8, 27'h00000002, 32'h00000400,
  1'd1,  5'd7, 27'h000000ad, 5'd30, 27'h00000220, 5'd16, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000113, 5'd26, 27'h0000021b, 5'd27, 27'h000003e5, 32'h00000400,
  1'd1,  5'd19, 27'h00000388, 5'd5, 27'h0000023f, 5'd6, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000343, 5'd6, 27'h00000224, 5'd19, 27'h0000021c, 32'h00000400,
  1'd1,  5'd20, 27'h00000076, 5'd6, 27'h0000005c, 5'd30, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000009e, 5'd18, 27'h00000072, 5'd6, 27'h000003eb, 32'h00000400,
  1'd1,  5'd19, 27'h0000009b, 5'd16, 27'h000002cf, 5'd17, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a9, 5'd16, 27'h000001a6, 5'd29, 27'h000003d9, 32'h00000400,
  1'd1,  5'd17, 27'h000003d0, 5'd28, 27'h0000016e, 5'd8, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000008b, 5'd26, 27'h00000361, 5'd18, 27'h000001c5, 32'h00000400,
  1'd1,  5'd15, 27'h000003c5, 5'd29, 27'h000001a7, 5'd27, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000152, 5'd9, 27'h000000ee, 5'd6, 27'h000002e7, 32'h00000400,
  1'd1,  5'd27, 27'h00000221, 5'd9, 27'h00000164, 5'd16, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000040, 5'd7, 27'h000000e2, 5'd27, 27'h000002b0, 32'h00000400,
  1'd1,  5'd28, 27'h00000266, 5'd18, 27'h0000022c, 5'd7, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001cf, 5'd20, 27'h000001ea, 5'd20, 27'h0000029c, 32'h00000400,
  1'd1,  5'd30, 27'h000003cb, 5'd18, 27'h0000001a, 5'd30, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000208, 5'd28, 27'h000003f4, 5'd8, 27'h000000a4, 32'h00000400,
  1'd1,  5'd29, 27'h00000184, 5'd29, 27'h00000214, 5'd15, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000289, 5'd26, 27'h00000277, 5'd28, 27'h00000374, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000003a8, 5'd0, 27'h0000032a, 5'd0, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000023c, 5'd1, 27'h00000106, 5'd12, 27'h000002a8, 32'h00000400,
  1'd1,  5'd2, 27'h00000109, 5'd2, 27'h0000023f, 5'd22, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003a4, 5'd11, 27'h0000025b, 5'd4, 27'h0000028b, 32'h00000400,
  1'd1,  5'd3, 27'h000002e6, 5'd14, 27'h000003e7, 5'd11, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d9, 5'd12, 27'h000002b1, 5'd25, 27'h00000340, 32'h00000400,
  1'd1,  5'd3, 27'h0000007c, 5'd22, 27'h000003e9, 5'd2, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026a, 5'd21, 27'h000002db, 5'd12, 27'h0000014f, 32'h00000400,
  1'd1,  5'd3, 27'h000000e1, 5'd22, 27'h0000014b, 5'd22, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f3, 5'd1, 27'h00000042, 5'd5, 27'h00000044, 32'h00000400,
  1'd1,  5'd14, 27'h0000014a, 5'd0, 27'h00000103, 5'd11, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f0, 5'd1, 27'h000001a5, 5'd21, 27'h00000274, 32'h00000400,
  1'd1,  5'd13, 27'h000000fb, 5'd12, 27'h00000319, 5'd3, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000181, 5'd14, 27'h00000308, 5'd14, 27'h000003ad, 32'h00000400,
  1'd1,  5'd13, 27'h0000036f, 5'd13, 27'h000002dd, 5'd22, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c0, 5'd21, 27'h00000138, 5'd4, 27'h0000015d, 32'h00000400,
  1'd1,  5'd10, 27'h00000170, 5'd25, 27'h000000a6, 5'd11, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000006f, 5'd25, 27'h00000029, 5'd23, 27'h000000aa, 32'h00000400,
  1'd1,  5'd23, 27'h00000347, 5'd0, 27'h000002ab, 5'd2, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000344, 5'd2, 27'h000001c8, 5'd15, 27'h00000158, 32'h00000400,
  1'd1,  5'd21, 27'h00000300, 5'd4, 27'h00000295, 5'd25, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000158, 5'd12, 27'h000001a8, 5'd2, 27'h0000002b, 32'h00000400,
  1'd1,  5'd22, 27'h00000355, 5'd10, 27'h0000028a, 5'd15, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a6, 5'd12, 27'h000000fa, 5'd23, 27'h0000020a, 32'h00000400,
  1'd1,  5'd20, 27'h000003b6, 5'd22, 27'h00000235, 5'd2, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000362, 5'd22, 27'h00000289, 5'd14, 27'h00000059, 32'h00000400,
  1'd1,  5'd23, 27'h000000f4, 5'd25, 27'h00000317, 5'd23, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000261, 5'd4, 27'h0000026c, 5'd8, 27'h00000139, 32'h00000400,
  1'd1,  5'd4, 27'h000000f0, 5'd3, 27'h00000314, 5'd15, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000231, 5'd0, 27'h00000303, 5'd28, 27'h00000380, 32'h00000400,
  1'd1,  5'd3, 27'h0000038b, 5'd11, 27'h000003d5, 5'd7, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d6, 5'd14, 27'h000000d9, 5'd17, 27'h00000352, 32'h00000400,
  1'd1,  5'd4, 27'h0000034c, 5'd15, 27'h0000000c, 5'd29, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b3, 5'd22, 27'h0000024d, 5'd10, 27'h00000016, 32'h00000400,
  1'd1,  5'd4, 27'h000000d6, 5'd25, 27'h00000107, 5'd16, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001cd, 5'd21, 27'h0000033e, 5'd27, 27'h00000002, 32'h00000400,
  1'd1,  5'd12, 27'h000003bb, 5'd2, 27'h00000346, 5'd6, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000172, 5'd3, 27'h00000344, 5'd16, 27'h0000001e, 32'h00000400,
  1'd1,  5'd11, 27'h000002fa, 5'd1, 27'h00000052, 5'd30, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008b, 5'd11, 27'h000000d7, 5'd8, 27'h000001ca, 32'h00000400,
  1'd1,  5'd14, 27'h000003d6, 5'd12, 27'h000003d8, 5'd18, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000396, 5'd12, 27'h00000151, 5'd25, 27'h000003e0, 32'h00000400,
  1'd1,  5'd13, 27'h0000016a, 5'd23, 27'h00000201, 5'd7, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013d, 5'd25, 27'h000001be, 5'd19, 27'h0000024e, 32'h00000400,
  1'd1,  5'd13, 27'h000003f1, 5'd23, 27'h00000356, 5'd28, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001dd, 5'd1, 27'h0000023c, 5'd10, 27'h0000010d, 32'h00000400,
  1'd1,  5'd21, 27'h000003b6, 5'd0, 27'h000002d8, 5'd17, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ff, 5'd0, 27'h00000354, 5'd30, 27'h000003e1, 32'h00000400,
  1'd1,  5'd21, 27'h0000001e, 5'd12, 27'h000001bb, 5'd5, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000295, 5'd14, 27'h0000003b, 5'd18, 27'h00000145, 32'h00000400,
  1'd1,  5'd23, 27'h00000030, 5'd14, 27'h000001db, 5'd28, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ad, 5'd21, 27'h00000311, 5'd10, 27'h000000d8, 32'h00000400,
  1'd1,  5'd24, 27'h00000154, 5'd21, 27'h00000230, 5'd16, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000019b, 5'd23, 27'h000002b6, 5'd27, 27'h00000179, 32'h00000400,
  1'd1,  5'd1, 27'h000001e4, 5'd9, 27'h00000386, 5'd4, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001d9, 5'd5, 27'h00000373, 5'd13, 27'h00000352, 32'h00000400,
  1'd1,  5'd4, 27'h0000017a, 5'd7, 27'h000000b6, 5'd20, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a3, 5'd15, 27'h00000303, 5'd4, 27'h000001f0, 32'h00000400,
  1'd1,  5'd4, 27'h00000189, 5'd18, 27'h00000345, 5'd11, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002b5, 5'd18, 27'h0000036b, 5'd23, 27'h000002a3, 32'h00000400,
  1'd1,  5'd2, 27'h000001f4, 5'd26, 27'h00000376, 5'd5, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000341, 5'd30, 27'h0000005b, 5'd10, 27'h000002d6, 32'h00000400,
  1'd1,  5'd0, 27'h00000219, 5'd30, 27'h00000294, 5'd22, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000374, 5'd5, 27'h000003a5, 5'd3, 27'h00000356, 32'h00000400,
  1'd1,  5'd13, 27'h00000168, 5'd7, 27'h000000fe, 5'd14, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000189, 5'd6, 27'h00000057, 5'd20, 27'h00000369, 32'h00000400,
  1'd1,  5'd13, 27'h00000211, 5'd19, 27'h000001d7, 5'd2, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020f, 5'd18, 27'h000002cf, 5'd13, 27'h000002f2, 32'h00000400,
  1'd1,  5'd10, 27'h000001bc, 5'd18, 27'h000003bc, 5'd22, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000231, 5'd28, 27'h000002bd, 5'd1, 27'h000000fe, 32'h00000400,
  1'd1,  5'd10, 27'h000001bd, 5'd29, 27'h000003f7, 5'd12, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000321, 5'd27, 27'h000001bf, 5'd24, 27'h00000221, 32'h00000400,
  1'd1,  5'd24, 27'h0000039d, 5'd7, 27'h000002cb, 5'd0, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000043, 5'd6, 27'h00000090, 5'd13, 27'h000000d0, 32'h00000400,
  1'd1,  5'd23, 27'h0000023c, 5'd7, 27'h000002d4, 5'd21, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003dc, 5'd19, 27'h0000026b, 5'd4, 27'h000000c4, 32'h00000400,
  1'd1,  5'd23, 27'h0000039b, 5'd17, 27'h0000039a, 5'd10, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000012f, 5'd20, 27'h00000083, 5'd22, 27'h0000031d, 32'h00000400,
  1'd1,  5'd22, 27'h000001bf, 5'd27, 27'h00000143, 5'd0, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002ec, 5'd26, 27'h000000ba, 5'd11, 27'h0000017f, 32'h00000400,
  1'd1,  5'd20, 27'h000003d9, 5'd27, 27'h00000363, 5'd23, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000025, 5'd5, 27'h000000bb, 5'd8, 27'h0000004d, 32'h00000400,
  1'd1,  5'd2, 27'h0000006b, 5'd9, 27'h00000334, 5'd20, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000382, 5'd7, 27'h000003f8, 5'd28, 27'h000002c1, 32'h00000400,
  1'd1,  5'd1, 27'h000003f8, 5'd18, 27'h000003c9, 5'd8, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000027b, 5'd19, 27'h000001d9, 5'd19, 27'h0000006e, 32'h00000400,
  1'd1,  5'd1, 27'h00000134, 5'd17, 27'h000001d0, 5'd30, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003a9, 5'd27, 27'h00000000, 5'd8, 27'h00000243, 32'h00000400,
  1'd1,  5'd3, 27'h000002c1, 5'd29, 27'h000002d4, 5'd18, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000213, 5'd30, 27'h00000236, 5'd26, 27'h000002a6, 32'h00000400,
  1'd1,  5'd11, 27'h00000069, 5'd9, 27'h0000017a, 5'd5, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002e3, 5'd6, 27'h00000205, 5'd15, 27'h000003a2, 32'h00000400,
  1'd1,  5'd11, 27'h000000e1, 5'd6, 27'h000000af, 5'd29, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000072, 5'd20, 27'h000000ee, 5'd8, 27'h00000088, 32'h00000400,
  1'd1,  5'd11, 27'h000000b1, 5'd19, 27'h00000260, 5'd20, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000237, 5'd19, 27'h000001dd, 5'd28, 27'h00000170, 32'h00000400,
  1'd1,  5'd14, 27'h000001d8, 5'd29, 27'h00000250, 5'd8, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000075, 5'd26, 27'h00000091, 5'd19, 27'h000003ed, 32'h00000400,
  1'd1,  5'd12, 27'h0000017d, 5'd28, 27'h000001e3, 5'd26, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000212, 5'd8, 27'h000001b8, 5'd6, 27'h0000035b, 32'h00000400,
  1'd1,  5'd24, 27'h0000001d, 5'd7, 27'h000000d4, 5'd18, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001b2, 5'd8, 27'h0000020d, 5'd28, 27'h00000204, 32'h00000400,
  1'd1,  5'd22, 27'h000002ba, 5'd20, 27'h0000015a, 5'd7, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000268, 5'd16, 27'h00000101, 5'd15, 27'h000003bc, 32'h00000400,
  1'd1,  5'd24, 27'h0000039b, 5'd16, 27'h0000023d, 5'd26, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a7, 5'd27, 27'h0000023a, 5'd6, 27'h00000211, 32'h00000400,
  1'd1,  5'd24, 27'h000002b3, 5'd25, 27'h000003bd, 5'd18, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000279, 5'd28, 27'h000001ca, 5'd27, 27'h000003c4, 32'h00000400,
  1'd1,  5'd6, 27'h000003f4, 5'd0, 27'h0000028e, 5'd8, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000274, 5'd4, 27'h0000014e, 5'd16, 27'h000000d9, 32'h00000400,
  1'd1,  5'd6, 27'h00000150, 5'd0, 27'h00000178, 5'd29, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ce, 5'd11, 27'h0000002a, 5'd4, 27'h000001e7, 32'h00000400,
  1'd1,  5'd9, 27'h000001b7, 5'd10, 27'h00000303, 5'd12, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000114, 5'd12, 27'h00000255, 5'd23, 27'h000003f7, 32'h00000400,
  1'd1,  5'd8, 27'h000000fe, 5'd24, 27'h000002a0, 5'd0, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c0, 5'd24, 27'h00000343, 5'd12, 27'h0000023b, 32'h00000400,
  1'd1,  5'd6, 27'h000002f9, 5'd24, 27'h0000003f, 5'd23, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000033d, 5'd2, 27'h000003db, 5'd8, 27'h000001d5, 32'h00000400,
  1'd1,  5'd19, 27'h00000214, 5'd5, 27'h0000006f, 5'd20, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c9, 5'd0, 27'h00000312, 5'd27, 27'h000003d8, 32'h00000400,
  1'd1,  5'd17, 27'h000002ba, 5'd13, 27'h000002f2, 5'd1, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000218, 5'd12, 27'h00000118, 5'd11, 27'h000000d6, 32'h00000400,
  1'd1,  5'd16, 27'h00000057, 5'd13, 27'h0000004e, 5'd25, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b8, 5'd23, 27'h00000184, 5'd1, 27'h00000387, 32'h00000400,
  1'd1,  5'd18, 27'h00000396, 5'd25, 27'h000000b5, 5'd14, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000240, 5'd25, 27'h00000097, 5'd23, 27'h00000298, 32'h00000400,
  1'd1,  5'd26, 27'h000000ec, 5'd3, 27'h000001f9, 5'd2, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000377, 5'd1, 27'h0000014e, 5'd10, 27'h000001b6, 32'h00000400,
  1'd1,  5'd29, 27'h0000008c, 5'd1, 27'h000002a4, 5'd22, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000370, 5'd13, 27'h0000013d, 5'd0, 27'h00000196, 32'h00000400,
  1'd1,  5'd29, 27'h00000115, 5'd11, 27'h00000314, 5'd13, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000160, 5'd12, 27'h0000021e, 5'd23, 27'h000002fa, 32'h00000400,
  1'd1,  5'd29, 27'h000003b3, 5'd25, 27'h00000125, 5'd0, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000065, 5'd21, 27'h000001ea, 5'd12, 27'h0000001c, 32'h00000400,
  1'd1,  5'd26, 27'h00000047, 5'd20, 27'h0000037d, 5'd22, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000013, 5'd3, 27'h000000f2, 5'd3, 27'h00000014, 32'h00000400,
  1'd1,  5'd9, 27'h0000034a, 5'd0, 27'h0000032a, 5'd15, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034c, 5'd1, 27'h000000c6, 5'd23, 27'h00000356, 32'h00000400,
  1'd1,  5'd9, 27'h0000004a, 5'd13, 27'h00000294, 5'd5, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000131, 5'd12, 27'h0000025e, 5'd18, 27'h0000004d, 32'h00000400,
  1'd1,  5'd6, 27'h000003d8, 5'd14, 27'h00000276, 5'd26, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000df, 5'd24, 27'h00000166, 5'd9, 27'h000000ff, 32'h00000400,
  1'd1,  5'd5, 27'h00000396, 5'd21, 27'h00000133, 5'd19, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000280, 5'd22, 27'h000003bb, 5'd26, 27'h000002e7, 32'h00000400,
  1'd1,  5'd20, 27'h000001ac, 5'd4, 27'h0000000d, 5'd1, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000c7, 5'd3, 27'h000002c1, 5'd11, 27'h000000a4, 32'h00000400,
  1'd1,  5'd18, 27'h000003f5, 5'd4, 27'h000000c2, 5'd22, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000138, 5'd13, 27'h000002be, 5'd7, 27'h00000320, 32'h00000400,
  1'd1,  5'd15, 27'h00000338, 5'd12, 27'h000002d3, 5'd17, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000142, 5'd11, 27'h000003e0, 5'd28, 27'h000003b3, 32'h00000400,
  1'd1,  5'd17, 27'h0000006f, 5'd23, 27'h0000019d, 5'd10, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000019a, 5'd24, 27'h000001bc, 5'd20, 27'h0000027c, 32'h00000400,
  1'd1,  5'd16, 27'h000001df, 5'd22, 27'h00000000, 5'd30, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f8, 5'd0, 27'h00000309, 5'd9, 27'h000002dc, 32'h00000400,
  1'd1,  5'd30, 27'h0000033c, 5'd3, 27'h00000373, 5'd19, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000041, 5'd2, 27'h000002a1, 5'd29, 27'h000002d0, 32'h00000400,
  1'd1,  5'd28, 27'h000001b7, 5'd14, 27'h0000038e, 5'd7, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ff, 5'd12, 27'h0000027b, 5'd20, 27'h00000187, 32'h00000400,
  1'd1,  5'd28, 27'h000000ef, 5'd13, 27'h000002dc, 5'd26, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001cb, 5'd22, 27'h0000033b, 5'd5, 27'h0000017e, 32'h00000400,
  1'd1,  5'd29, 27'h000002e2, 5'd21, 27'h000000ca, 5'd17, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000008e, 5'd25, 27'h0000016f, 5'd30, 27'h000000ef, 32'h00000400,
  1'd1,  5'd9, 27'h0000013f, 5'd7, 27'h00000198, 5'd2, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002de, 5'd8, 27'h0000025c, 5'd10, 27'h0000034c, 32'h00000400,
  1'd1,  5'd8, 27'h00000358, 5'd10, 27'h000000a9, 5'd25, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c2, 5'd16, 27'h000003ad, 5'd2, 27'h0000023b, 32'h00000400,
  1'd1,  5'd7, 27'h000001c5, 5'd15, 27'h000002ec, 5'd13, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003f9, 5'd20, 27'h000001d0, 5'd20, 27'h00000323, 32'h00000400,
  1'd1,  5'd9, 27'h000000f1, 5'd30, 27'h0000037d, 5'd1, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000000e, 5'd28, 27'h0000034f, 5'd12, 27'h000002d3, 32'h00000400,
  1'd1,  5'd7, 27'h000003a0, 5'd28, 27'h000001cd, 5'd25, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000396, 5'd9, 27'h000003cf, 5'd4, 27'h000001f9, 32'h00000400,
  1'd1,  5'd16, 27'h0000035c, 5'd8, 27'h00000107, 5'd14, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ad, 5'd7, 27'h000000d1, 5'd22, 27'h00000179, 32'h00000400,
  1'd1,  5'd15, 27'h000003f6, 5'd16, 27'h0000002f, 5'd5, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000037f, 5'd18, 27'h0000019f, 5'd12, 27'h00000128, 32'h00000400,
  1'd1,  5'd17, 27'h0000021a, 5'd20, 27'h00000127, 5'd21, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001fb, 5'd29, 27'h000000dd, 5'd2, 27'h000000fa, 32'h00000400,
  1'd1,  5'd20, 27'h00000220, 5'd28, 27'h0000027d, 5'd12, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c9, 5'd29, 27'h00000163, 5'd21, 27'h00000368, 32'h00000400,
  1'd1,  5'd30, 27'h00000383, 5'd8, 27'h000001a3, 5'd2, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ed, 5'd6, 27'h0000013a, 5'd10, 27'h000002f3, 32'h00000400,
  1'd1,  5'd28, 27'h0000025e, 5'd9, 27'h00000119, 5'd22, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000024b, 5'd19, 27'h0000021b, 5'd4, 27'h00000210, 32'h00000400,
  1'd1,  5'd29, 27'h000002a5, 5'd17, 27'h00000294, 5'd15, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003f2, 5'd16, 27'h00000167, 5'd20, 27'h00000337, 32'h00000400,
  1'd1,  5'd30, 27'h00000216, 5'd27, 27'h0000014b, 5'd3, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003ec, 5'd29, 27'h0000001c, 5'd11, 27'h000001f2, 32'h00000400,
  1'd1,  5'd28, 27'h000003da, 5'd30, 27'h0000035b, 5'd24, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ba, 5'd6, 27'h00000362, 5'd9, 27'h00000272, 32'h00000400,
  1'd1,  5'd6, 27'h00000056, 5'd10, 27'h00000112, 5'd20, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000290, 5'd5, 27'h000001e6, 5'd27, 27'h000001a2, 32'h00000400,
  1'd1,  5'd8, 27'h000003a7, 5'd19, 27'h0000009a, 5'd7, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ed, 5'd18, 27'h000001ec, 5'd16, 27'h000000ab, 32'h00000400,
  1'd1,  5'd6, 27'h00000100, 5'd17, 27'h00000177, 5'd27, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000051, 5'd30, 27'h0000033b, 5'd5, 27'h000002ad, 32'h00000400,
  1'd1,  5'd6, 27'h0000016f, 5'd26, 27'h000002fd, 5'd18, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007e, 5'd29, 27'h000002ac, 5'd27, 27'h0000008f, 32'h00000400,
  1'd1,  5'd19, 27'h00000312, 5'd7, 27'h00000135, 5'd6, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000198, 5'd10, 27'h00000068, 5'd18, 27'h00000317, 32'h00000400,
  1'd1,  5'd16, 27'h00000116, 5'd8, 27'h00000357, 5'd29, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000027, 5'd18, 27'h0000028b, 5'd8, 27'h0000009f, 32'h00000400,
  1'd1,  5'd18, 27'h0000032f, 5'd17, 27'h000002cc, 5'd17, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002e2, 5'd15, 27'h0000028b, 5'd30, 27'h000000f0, 32'h00000400,
  1'd1,  5'd16, 27'h00000371, 5'd27, 27'h0000026d, 5'd9, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002be, 5'd27, 27'h00000285, 5'd18, 27'h000003cd, 32'h00000400,
  1'd1,  5'd15, 27'h000002ce, 5'd27, 27'h00000189, 5'd27, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000120, 5'd10, 27'h00000106, 5'd7, 27'h000000a0, 32'h00000400,
  1'd1,  5'd25, 27'h00000379, 5'd6, 27'h000002e1, 5'd20, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000024, 5'd7, 27'h000002b7, 5'd26, 27'h00000365, 32'h00000400,
  1'd1,  5'd27, 27'h0000026c, 5'd16, 27'h0000031b, 5'd7, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000002f, 5'd18, 27'h0000005b, 5'd15, 27'h00000354, 32'h00000400,
  1'd1,  5'd26, 27'h000003e3, 5'd20, 27'h000001e4, 5'd27, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000100, 5'd30, 27'h00000175, 5'd7, 27'h000000e5, 32'h00000400,
  1'd1,  5'd28, 27'h000003ce, 5'd29, 27'h000003eb, 5'd19, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002b8, 5'd26, 27'h0000015f, 5'd30, 27'h00000107, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000039b, 5'd2, 27'h0000030f, 5'd4, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000384, 5'd2, 27'h00000218, 5'd10, 27'h000002c2, 32'h00000400,
  1'd1,  5'd4, 27'h00000055, 5'd3, 27'h000002ac, 5'd22, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000037d, 5'd14, 27'h000003be, 5'd0, 27'h000001a8, 32'h00000400,
  1'd1,  5'd0, 27'h000002b8, 5'd12, 27'h00000375, 5'd11, 27'h00000242, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000034, 5'd12, 27'h0000009a, 5'd24, 27'h000001db, 32'h00000400,
  1'd1,  5'd1, 27'h00000298, 5'd24, 27'h00000323, 5'd2, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e9, 5'd25, 27'h00000322, 5'd12, 27'h00000221, 32'h00000400,
  1'd1,  5'd3, 27'h000001fd, 5'd23, 27'h0000002b, 5'd22, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000017, 5'd0, 27'h000003b6, 5'd2, 27'h0000010b, 32'h00000400,
  1'd1,  5'd12, 27'h0000022f, 5'd1, 27'h0000016c, 5'd11, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000005c, 5'd3, 27'h000002de, 5'd23, 27'h00000304, 32'h00000400,
  1'd1,  5'd12, 27'h00000174, 5'd10, 27'h0000039e, 5'd1, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000033b, 5'd13, 27'h00000282, 5'd11, 27'h00000092, 32'h00000400,
  1'd1,  5'd14, 27'h00000239, 5'd13, 27'h0000027d, 5'd20, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003f1, 5'd25, 27'h00000175, 5'd2, 27'h00000075, 32'h00000400,
  1'd1,  5'd12, 27'h00000278, 5'd23, 27'h0000002d, 5'd12, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000d0, 5'd23, 27'h0000027e, 5'd22, 27'h00000307, 32'h00000400,
  1'd1,  5'd21, 27'h00000290, 5'd4, 27'h0000034f, 5'd1, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000010b, 5'd2, 27'h0000018f, 5'd11, 27'h00000303, 32'h00000400,
  1'd1,  5'd22, 27'h000000ad, 5'd4, 27'h00000319, 5'd25, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000006b, 5'd12, 27'h00000216, 5'd3, 27'h0000006a, 32'h00000400,
  1'd1,  5'd23, 27'h0000009c, 5'd13, 27'h000002bc, 5'd11, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000015d, 5'd11, 27'h00000339, 5'd21, 27'h00000154, 32'h00000400,
  1'd1,  5'd21, 27'h000002d9, 5'd25, 27'h00000098, 5'd4, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a2, 5'd23, 27'h000001cd, 5'd11, 27'h000003d4, 32'h00000400,
  1'd1,  5'd23, 27'h000003a3, 5'd23, 27'h00000078, 5'd23, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f2, 5'd0, 27'h0000016e, 5'd5, 27'h0000021b, 32'h00000400,
  1'd1,  5'd2, 27'h000000e0, 5'd2, 27'h00000048, 5'd16, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000200, 5'd3, 27'h0000024f, 5'd30, 27'h000002a2, 32'h00000400,
  1'd1,  5'd0, 27'h00000298, 5'd15, 27'h00000046, 5'd5, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000c4, 5'd12, 27'h00000303, 5'd20, 27'h000001e3, 32'h00000400,
  1'd1,  5'd4, 27'h0000018e, 5'd10, 27'h0000021e, 5'd27, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002d9, 5'd22, 27'h0000013d, 5'd10, 27'h00000033, 32'h00000400,
  1'd1,  5'd2, 27'h00000400, 5'd22, 27'h00000203, 5'd20, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017a, 5'd22, 27'h000001d7, 5'd26, 27'h000003ab, 32'h00000400,
  1'd1,  5'd11, 27'h000002eb, 5'd4, 27'h00000077, 5'd9, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000199, 5'd2, 27'h0000012c, 5'd16, 27'h000002e8, 32'h00000400,
  1'd1,  5'd13, 27'h000000a3, 5'd4, 27'h0000001e, 5'd29, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003b0, 5'd11, 27'h000002eb, 5'd5, 27'h000002e4, 32'h00000400,
  1'd1,  5'd10, 27'h00000192, 5'd12, 27'h0000029b, 5'd19, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000019e, 5'd10, 27'h000003e2, 5'd27, 27'h000001b5, 32'h00000400,
  1'd1,  5'd15, 27'h00000022, 5'd24, 27'h00000160, 5'd7, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000007, 5'd24, 27'h000003a2, 5'd20, 27'h0000014e, 32'h00000400,
  1'd1,  5'd13, 27'h00000152, 5'd24, 27'h00000280, 5'd30, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000335, 5'd1, 27'h00000299, 5'd8, 27'h00000399, 32'h00000400,
  1'd1,  5'd24, 27'h00000046, 5'd3, 27'h000003d9, 5'd20, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000035d, 5'd3, 27'h00000185, 5'd29, 27'h000000e0, 32'h00000400,
  1'd1,  5'd23, 27'h0000036b, 5'd14, 27'h000002fe, 5'd10, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000011, 5'd11, 27'h0000029c, 5'd17, 27'h0000011a, 32'h00000400,
  1'd1,  5'd22, 27'h000002e2, 5'd11, 27'h000003cd, 5'd30, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000036d, 5'd20, 27'h000002e2, 5'd9, 27'h000000d6, 32'h00000400,
  1'd1,  5'd23, 27'h000000bc, 5'd21, 27'h000003a2, 5'd15, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000360, 5'd23, 27'h00000392, 5'd29, 27'h00000243, 32'h00000400,
  1'd1,  5'd0, 27'h0000032b, 5'd8, 27'h00000320, 5'd2, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b9, 5'd8, 27'h00000136, 5'd10, 27'h00000204, 32'h00000400,
  1'd1,  5'd2, 27'h000001db, 5'd6, 27'h000003c3, 5'd22, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026b, 5'd20, 27'h0000017c, 5'd1, 27'h000002d2, 32'h00000400,
  1'd1,  5'd0, 27'h00000196, 5'd15, 27'h00000239, 5'd11, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000178, 5'd20, 27'h0000008f, 5'd20, 27'h00000345, 32'h00000400,
  1'd1,  5'd0, 27'h0000029f, 5'd26, 27'h000000aa, 5'd0, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000011c, 5'd30, 27'h000000de, 5'd11, 27'h000001c2, 32'h00000400,
  1'd1,  5'd0, 27'h00000174, 5'd27, 27'h00000311, 5'd21, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000006a, 5'd7, 27'h00000058, 5'd0, 27'h000003f7, 32'h00000400,
  1'd1,  5'd15, 27'h0000011e, 5'd6, 27'h000003fb, 5'd12, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000032b, 5'd5, 27'h000003dc, 5'd22, 27'h00000079, 32'h00000400,
  1'd1,  5'd14, 27'h00000219, 5'd19, 27'h00000130, 5'd4, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002bc, 5'd16, 27'h00000007, 5'd14, 27'h00000000, 32'h00000400,
  1'd1,  5'd12, 27'h00000171, 5'd16, 27'h000000f8, 5'd24, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000163, 5'd30, 27'h000003fc, 5'd0, 27'h0000036d, 32'h00000400,
  1'd1,  5'd14, 27'h0000019d, 5'd27, 27'h000000db, 5'd12, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000025b, 5'd29, 27'h00000278, 5'd22, 27'h000003bf, 32'h00000400,
  1'd1,  5'd20, 27'h000003cb, 5'd9, 27'h000002b6, 5'd0, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003d5, 5'd6, 27'h0000032c, 5'd13, 27'h00000191, 32'h00000400,
  1'd1,  5'd23, 27'h000002d2, 5'd7, 27'h000003e0, 5'd21, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b3, 5'd17, 27'h0000037e, 5'd3, 27'h00000145, 32'h00000400,
  1'd1,  5'd24, 27'h000001f3, 5'd19, 27'h000001b7, 5'd15, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000281, 5'd19, 27'h0000039e, 5'd24, 27'h000001d5, 32'h00000400,
  1'd1,  5'd24, 27'h00000120, 5'd28, 27'h00000165, 5'd1, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000332, 5'd27, 27'h00000381, 5'd14, 27'h000003c8, 32'h00000400,
  1'd1,  5'd22, 27'h0000013e, 5'd27, 27'h000003eb, 5'd20, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f5, 5'd9, 27'h000002fa, 5'd9, 27'h00000287, 32'h00000400,
  1'd1,  5'd4, 27'h000003d0, 5'd9, 27'h0000027c, 5'd16, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a4, 5'd5, 27'h000002d3, 5'd30, 27'h000003d5, 32'h00000400,
  1'd1,  5'd2, 27'h000001ff, 5'd19, 27'h00000287, 5'd7, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f7, 5'd18, 27'h00000281, 5'd18, 27'h000000ce, 32'h00000400,
  1'd1,  5'd0, 27'h0000025e, 5'd20, 27'h000001b2, 5'd26, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000002c, 5'd29, 27'h00000114, 5'd8, 27'h00000193, 32'h00000400,
  1'd1,  5'd0, 27'h000002de, 5'd27, 27'h00000335, 5'd17, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000018, 5'd30, 27'h000001b8, 5'd26, 27'h00000230, 32'h00000400,
  1'd1,  5'd11, 27'h000000a9, 5'd5, 27'h00000255, 5'd5, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000008f, 5'd5, 27'h00000210, 5'd16, 27'h000001f7, 32'h00000400,
  1'd1,  5'd10, 27'h0000024d, 5'd10, 27'h00000088, 5'd28, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a2, 5'd20, 27'h00000171, 5'd8, 27'h00000093, 32'h00000400,
  1'd1,  5'd11, 27'h00000260, 5'd19, 27'h00000246, 5'd16, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000212, 5'd18, 27'h00000190, 5'd29, 27'h0000015e, 32'h00000400,
  1'd1,  5'd13, 27'h000002cf, 5'd29, 27'h00000074, 5'd8, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000184, 5'd29, 27'h000003ad, 5'd15, 27'h000002e8, 32'h00000400,
  1'd1,  5'd14, 27'h000002e3, 5'd27, 27'h00000375, 5'd29, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000030d, 5'd6, 27'h00000200, 5'd5, 27'h000000e6, 32'h00000400,
  1'd1,  5'd25, 27'h00000229, 5'd8, 27'h00000046, 5'd20, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000029e, 5'd9, 27'h000001fc, 5'd30, 27'h00000020, 32'h00000400,
  1'd1,  5'd23, 27'h0000027e, 5'd17, 27'h00000108, 5'd8, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000029e, 5'd17, 27'h000001f5, 5'd20, 27'h000001d6, 32'h00000400,
  1'd1,  5'd22, 27'h00000370, 5'd18, 27'h00000195, 5'd26, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000e9, 5'd26, 27'h00000358, 5'd9, 27'h000003c6, 32'h00000400,
  1'd1,  5'd23, 27'h000000e2, 5'd30, 27'h0000035f, 5'd16, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000037b, 5'd27, 27'h00000103, 5'd27, 27'h00000345, 32'h00000400,
  1'd1,  5'd6, 27'h00000054, 5'd4, 27'h000003f5, 5'd10, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000010, 5'd4, 27'h000003c5, 5'd15, 27'h00000286, 32'h00000400,
  1'd1,  5'd7, 27'h0000039b, 5'd1, 27'h00000230, 5'd28, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003bf, 5'd10, 27'h000002a4, 5'd1, 27'h0000020f, 32'h00000400,
  1'd1,  5'd6, 27'h00000033, 5'd13, 27'h00000012, 5'd11, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000289, 5'd12, 27'h00000002, 5'd21, 27'h00000162, 32'h00000400,
  1'd1,  5'd7, 27'h000001b3, 5'd20, 27'h0000033c, 5'd0, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000a8, 5'd25, 27'h0000023a, 5'd14, 27'h00000049, 32'h00000400,
  1'd1,  5'd9, 27'h00000329, 5'd23, 27'h00000271, 5'd23, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000253, 5'd1, 27'h0000028a, 5'd6, 27'h00000335, 32'h00000400,
  1'd1,  5'd16, 27'h000002c8, 5'd0, 27'h0000031c, 5'd19, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c6, 5'd2, 27'h0000017b, 5'd30, 27'h00000280, 32'h00000400,
  1'd1,  5'd16, 27'h00000164, 5'd13, 27'h000001c3, 5'd3, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000035a, 5'd10, 27'h00000183, 5'd12, 27'h000000dd, 32'h00000400,
  1'd1,  5'd19, 27'h0000012e, 5'd12, 27'h000002aa, 5'd21, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ab, 5'd22, 27'h000002b9, 5'd4, 27'h000003ba, 32'h00000400,
  1'd1,  5'd20, 27'h00000125, 5'd24, 27'h0000000e, 5'd10, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a4, 5'd24, 27'h00000235, 5'd21, 27'h000001ad, 32'h00000400,
  1'd1,  5'd27, 27'h00000055, 5'd2, 27'h000003a1, 5'd2, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c6, 5'd2, 27'h00000393, 5'd14, 27'h000001bb, 32'h00000400,
  1'd1,  5'd29, 27'h0000036e, 5'd2, 27'h0000037e, 5'd22, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000014a, 5'd14, 27'h000001c7, 5'd2, 27'h00000097, 32'h00000400,
  1'd1,  5'd28, 27'h0000011c, 5'd14, 27'h0000009b, 5'd14, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001c2, 5'd12, 27'h000001c5, 5'd23, 27'h00000319, 32'h00000400,
  1'd1,  5'd30, 27'h00000184, 5'd25, 27'h0000024a, 5'd2, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003b2, 5'd25, 27'h00000242, 5'd12, 27'h0000036a, 32'h00000400,
  1'd1,  5'd27, 27'h00000066, 5'd21, 27'h00000025, 5'd25, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000219, 5'd4, 27'h00000091, 5'd2, 27'h0000007f, 32'h00000400,
  1'd1,  5'd9, 27'h00000300, 5'd3, 27'h00000289, 5'd12, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000013d, 5'd3, 27'h0000010d, 5'd22, 27'h00000333, 32'h00000400,
  1'd1,  5'd8, 27'h000001f3, 5'd12, 27'h00000109, 5'd9, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000379, 5'd14, 27'h0000039b, 5'd16, 27'h00000175, 32'h00000400,
  1'd1,  5'd9, 27'h00000211, 5'd15, 27'h0000019f, 5'd27, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000394, 5'd24, 27'h00000245, 5'd9, 27'h00000130, 32'h00000400,
  1'd1,  5'd8, 27'h0000009a, 5'd22, 27'h00000122, 5'd20, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000198, 5'd25, 27'h00000099, 5'd28, 27'h00000089, 32'h00000400,
  1'd1,  5'd17, 27'h000001d3, 5'd2, 27'h000001a9, 5'd2, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000a7, 5'd5, 27'h0000007e, 5'd11, 27'h000003f9, 32'h00000400,
  1'd1,  5'd20, 27'h00000110, 5'd1, 27'h0000034c, 5'd24, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006b, 5'd13, 27'h000001bb, 5'd9, 27'h0000017e, 32'h00000400,
  1'd1,  5'd19, 27'h000001f3, 5'd14, 27'h0000038b, 5'd20, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000022, 5'd13, 27'h0000028a, 5'd27, 27'h0000015c, 32'h00000400,
  1'd1,  5'd16, 27'h000000a7, 5'd22, 27'h00000028, 5'd9, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000033, 5'd21, 27'h000000da, 5'd17, 27'h00000049, 32'h00000400,
  1'd1,  5'd17, 27'h000001ff, 5'd25, 27'h00000184, 5'd26, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000011f, 5'd2, 27'h00000132, 5'd5, 27'h000001c1, 32'h00000400,
  1'd1,  5'd26, 27'h000002c9, 5'd3, 27'h00000352, 5'd19, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000264, 5'd3, 27'h0000001d, 5'd27, 27'h00000311, 32'h00000400,
  1'd1,  5'd27, 27'h000003ce, 5'd14, 27'h0000003c, 5'd7, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000039d, 5'd11, 27'h00000378, 5'd18, 27'h00000143, 32'h00000400,
  1'd1,  5'd30, 27'h00000075, 5'd12, 27'h00000126, 5'd27, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000232, 5'd23, 27'h000001ea, 5'd5, 27'h0000029d, 32'h00000400,
  1'd1,  5'd28, 27'h00000316, 5'd21, 27'h00000367, 5'd18, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000c8, 5'd24, 27'h0000029a, 5'd30, 27'h00000351, 32'h00000400,
  1'd1,  5'd9, 27'h0000039c, 5'd6, 27'h00000075, 5'd3, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000138, 5'd7, 27'h0000030c, 5'd13, 27'h00000020, 32'h00000400,
  1'd1,  5'd9, 27'h0000038c, 5'd9, 27'h0000016d, 5'd22, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000005, 5'd16, 27'h00000270, 5'd4, 27'h0000031f, 32'h00000400,
  1'd1,  5'd8, 27'h00000240, 5'd17, 27'h000001e7, 5'd15, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038c, 5'd18, 27'h00000285, 5'd24, 27'h0000008b, 32'h00000400,
  1'd1,  5'd5, 27'h00000259, 5'd29, 27'h0000029f, 5'd4, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e3, 5'd28, 27'h00000074, 5'd12, 27'h00000373, 32'h00000400,
  1'd1,  5'd8, 27'h00000256, 5'd27, 27'h00000364, 5'd23, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000263, 5'd6, 27'h000001f4, 5'd4, 27'h00000182, 32'h00000400,
  1'd1,  5'd19, 27'h00000118, 5'd5, 27'h00000361, 5'd14, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a8, 5'd10, 27'h00000151, 5'd23, 27'h00000271, 32'h00000400,
  1'd1,  5'd17, 27'h00000013, 5'd20, 27'h00000269, 5'd1, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000be, 5'd18, 27'h00000135, 5'd12, 27'h00000034, 32'h00000400,
  1'd1,  5'd19, 27'h000002ad, 5'd17, 27'h00000031, 5'd25, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b5, 5'd28, 27'h000000ac, 5'd1, 27'h0000036c, 32'h00000400,
  1'd1,  5'd19, 27'h0000028c, 5'd26, 27'h00000286, 5'd14, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000c6, 5'd26, 27'h0000028a, 5'd23, 27'h000001f8, 32'h00000400,
  1'd1,  5'd28, 27'h00000006, 5'd8, 27'h00000215, 5'd0, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000db, 5'd8, 27'h000000fb, 5'd14, 27'h00000141, 32'h00000400,
  1'd1,  5'd30, 27'h000001c5, 5'd6, 27'h00000111, 5'd25, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b2, 5'd19, 27'h00000371, 5'd4, 27'h00000009, 32'h00000400,
  1'd1,  5'd29, 27'h000003a8, 5'd18, 27'h000001d7, 5'd11, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000144, 5'd18, 27'h0000038c, 5'd24, 27'h00000329, 32'h00000400,
  1'd1,  5'd29, 27'h000003bc, 5'd27, 27'h00000242, 5'd0, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a0, 5'd26, 27'h00000322, 5'd13, 27'h00000199, 32'h00000400,
  1'd1,  5'd26, 27'h000000cc, 5'd30, 27'h00000289, 5'd23, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000271, 5'd7, 27'h0000028a, 5'd9, 27'h000003b5, 32'h00000400,
  1'd1,  5'd5, 27'h000003ca, 5'd5, 27'h000002f0, 5'd19, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000250, 5'd6, 27'h0000021a, 5'd26, 27'h0000017f, 32'h00000400,
  1'd1,  5'd8, 27'h00000091, 5'd19, 27'h00000299, 5'd7, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b7, 5'd15, 27'h0000020c, 5'd18, 27'h000003a2, 32'h00000400,
  1'd1,  5'd7, 27'h00000319, 5'd19, 27'h00000302, 5'd27, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000055, 5'd27, 27'h00000015, 5'd9, 27'h0000020f, 32'h00000400,
  1'd1,  5'd8, 27'h00000167, 5'd29, 27'h000000a3, 5'd17, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e7, 5'd27, 27'h00000345, 5'd26, 27'h000001ca, 32'h00000400,
  1'd1,  5'd20, 27'h0000023e, 5'd7, 27'h0000024c, 5'd8, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b5, 5'd5, 27'h00000284, 5'd18, 27'h00000159, 32'h00000400,
  1'd1,  5'd16, 27'h00000387, 5'd9, 27'h000000ef, 5'd27, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003f9, 5'd15, 27'h00000245, 5'd7, 27'h00000138, 32'h00000400,
  1'd1,  5'd18, 27'h00000114, 5'd20, 27'h000000b7, 5'd17, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000032e, 5'd16, 27'h000002f7, 5'd30, 27'h00000099, 32'h00000400,
  1'd1,  5'd17, 27'h00000387, 5'd28, 27'h000003ed, 5'd8, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000e6, 5'd28, 27'h000002f0, 5'd18, 27'h0000036c, 32'h00000400,
  1'd1,  5'd16, 27'h000003f6, 5'd29, 27'h000002a9, 5'd29, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000320, 5'd8, 27'h00000178, 5'd8, 27'h00000110, 32'h00000400,
  1'd1,  5'd27, 27'h00000199, 5'd7, 27'h00000244, 5'd17, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000014f, 5'd6, 27'h000000de, 5'd28, 27'h00000338, 32'h00000400,
  1'd1,  5'd27, 27'h00000340, 5'd16, 27'h000001d2, 5'd8, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017e, 5'd18, 27'h0000003d, 5'd15, 27'h000002ea, 32'h00000400,
  1'd1,  5'd27, 27'h0000023c, 5'd17, 27'h000002ff, 5'd29, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ef, 5'd29, 27'h0000023f, 5'd10, 27'h000000b0, 32'h00000400,
  1'd1,  5'd26, 27'h000003a9, 5'd30, 27'h00000062, 5'd15, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000064, 5'd26, 27'h0000035a, 5'd26, 27'h0000016f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000042, 5'd1, 27'h0000032b, 5'd0, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000140, 5'd3, 27'h00000272, 5'd14, 27'h00000021, 32'h00000400,
  1'd1,  5'd4, 27'h0000019c, 5'd0, 27'h000001a1, 5'd21, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000018a, 5'd11, 27'h00000183, 5'd1, 27'h0000029d, 32'h00000400,
  1'd1,  5'd3, 27'h0000006d, 5'd10, 27'h000003f0, 5'd12, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000105, 5'd14, 27'h0000012a, 5'd23, 27'h00000106, 32'h00000400,
  1'd1,  5'd3, 27'h00000210, 5'd22, 27'h000003cc, 5'd3, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000001b, 5'd21, 27'h000002a8, 5'd14, 27'h000000e0, 32'h00000400,
  1'd1,  5'd2, 27'h0000015c, 5'd25, 27'h00000277, 5'd24, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000011, 5'd1, 27'h000003b1, 5'd3, 27'h0000000d, 32'h00000400,
  1'd1,  5'd11, 27'h00000005, 5'd1, 27'h00000370, 5'd14, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000134, 5'd0, 27'h000003a3, 5'd25, 27'h00000207, 32'h00000400,
  1'd1,  5'd11, 27'h00000181, 5'd10, 27'h0000022b, 5'd4, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018c, 5'd13, 27'h0000030d, 5'd11, 27'h000000df, 32'h00000400,
  1'd1,  5'd13, 27'h000000bc, 5'd10, 27'h000001b2, 5'd21, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000319, 5'd22, 27'h00000397, 5'd3, 27'h00000025, 32'h00000400,
  1'd1,  5'd14, 27'h000000dd, 5'd21, 27'h00000135, 5'd12, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001b2, 5'd21, 27'h0000036a, 5'd21, 27'h00000140, 32'h00000400,
  1'd1,  5'd23, 27'h000003e6, 5'd4, 27'h000000e3, 5'd4, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000166, 5'd0, 27'h00000066, 5'd11, 27'h00000194, 32'h00000400,
  1'd1,  5'd21, 27'h000001d5, 5'd3, 27'h000001ff, 5'd23, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002ae, 5'd10, 27'h0000018d, 5'd2, 27'h000003f0, 32'h00000400,
  1'd1,  5'd23, 27'h00000193, 5'd13, 27'h0000015e, 5'd14, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000113, 5'd10, 27'h00000177, 5'd23, 27'h000000c2, 32'h00000400,
  1'd1,  5'd22, 27'h0000010f, 5'd22, 27'h000002da, 5'd2, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003db, 5'd20, 27'h0000035a, 5'd10, 27'h00000332, 32'h00000400,
  1'd1,  5'd25, 27'h0000001d, 5'd23, 27'h00000150, 5'd22, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ba, 5'd3, 27'h000002c8, 5'd6, 27'h00000172, 32'h00000400,
  1'd1,  5'd1, 27'h000001fb, 5'd3, 27'h000002d9, 5'd17, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002d4, 5'd0, 27'h0000009c, 5'd27, 27'h000002b3, 32'h00000400,
  1'd1,  5'd1, 27'h000001c4, 5'd10, 27'h000002af, 5'd7, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000027, 5'd13, 27'h000001f5, 5'd17, 27'h00000326, 32'h00000400,
  1'd1,  5'd2, 27'h000002a8, 5'd13, 27'h0000008c, 5'd29, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000059, 5'd23, 27'h00000146, 5'd6, 27'h000001e5, 32'h00000400,
  1'd1,  5'd1, 27'h00000142, 5'd22, 27'h000002f9, 5'd15, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000005f, 5'd21, 27'h00000204, 5'd26, 27'h00000033, 32'h00000400,
  1'd1,  5'd13, 27'h0000038d, 5'd0, 27'h0000003a, 5'd7, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a8, 5'd2, 27'h000000d2, 5'd17, 27'h00000242, 32'h00000400,
  1'd1,  5'd11, 27'h00000046, 5'd4, 27'h000002e6, 5'd28, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000020c, 5'd14, 27'h00000240, 5'd6, 27'h0000016b, 32'h00000400,
  1'd1,  5'd12, 27'h00000142, 5'd11, 27'h00000064, 5'd19, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035a, 5'd11, 27'h00000368, 5'd30, 27'h0000031c, 32'h00000400,
  1'd1,  5'd15, 27'h0000000b, 5'd23, 27'h000002cd, 5'd7, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000004f, 5'd24, 27'h00000070, 5'd18, 27'h00000354, 32'h00000400,
  1'd1,  5'd11, 27'h0000003d, 5'd25, 27'h000000bc, 5'd30, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003fc, 5'd3, 27'h0000004e, 5'd5, 27'h000002c8, 32'h00000400,
  1'd1,  5'd22, 27'h000003b3, 5'd4, 27'h00000044, 5'd18, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001ed, 5'd2, 27'h00000362, 5'd26, 27'h0000031f, 32'h00000400,
  1'd1,  5'd24, 27'h000003b9, 5'd14, 27'h000002e2, 5'd5, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000383, 5'd12, 27'h000000e8, 5'd16, 27'h000001c9, 32'h00000400,
  1'd1,  5'd24, 27'h000003e1, 5'd15, 27'h0000006a, 5'd26, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a7, 5'd21, 27'h00000129, 5'd5, 27'h000003c7, 32'h00000400,
  1'd1,  5'd25, 27'h00000150, 5'd22, 27'h000000e9, 5'd16, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000368, 5'd21, 27'h0000022d, 5'd29, 27'h00000014, 32'h00000400,
  1'd1,  5'd2, 27'h00000235, 5'd9, 27'h00000316, 5'd2, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003af, 5'd6, 27'h0000010c, 5'd13, 27'h000003e4, 32'h00000400,
  1'd1,  5'd0, 27'h0000033d, 5'd8, 27'h000002d2, 5'd24, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b4, 5'd18, 27'h000001a6, 5'd4, 27'h00000346, 32'h00000400,
  1'd1,  5'd4, 27'h000001d6, 5'd17, 27'h00000026, 5'd14, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000199, 5'd19, 27'h000000e5, 5'd24, 27'h0000011d, 32'h00000400,
  1'd1,  5'd2, 27'h00000151, 5'd26, 27'h00000119, 5'd1, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ff, 5'd30, 27'h00000378, 5'd14, 27'h000002c5, 32'h00000400,
  1'd1,  5'd3, 27'h00000205, 5'd27, 27'h00000081, 5'd22, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001d1, 5'd9, 27'h00000172, 5'd4, 27'h000001ad, 32'h00000400,
  1'd1,  5'd10, 27'h000003fb, 5'd10, 27'h00000080, 5'd12, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000185, 5'd7, 27'h00000027, 5'd22, 27'h000003aa, 32'h00000400,
  1'd1,  5'd12, 27'h0000039f, 5'd19, 27'h00000095, 5'd4, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c6, 5'd19, 27'h00000094, 5'd15, 27'h0000004b, 32'h00000400,
  1'd1,  5'd11, 27'h0000013c, 5'd17, 27'h000000d5, 5'd20, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000022e, 5'd30, 27'h00000160, 5'd3, 27'h000002b3, 32'h00000400,
  1'd1,  5'd15, 27'h00000082, 5'd30, 27'h00000379, 5'd10, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000014c, 5'd26, 27'h00000375, 5'd24, 27'h000000fb, 32'h00000400,
  1'd1,  5'd25, 27'h00000105, 5'd5, 27'h000003a8, 5'd1, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000023, 5'd8, 27'h00000117, 5'd12, 27'h00000123, 32'h00000400,
  1'd1,  5'd23, 27'h00000282, 5'd6, 27'h0000016e, 5'd23, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000035f, 5'd19, 27'h0000011a, 5'd1, 27'h00000286, 32'h00000400,
  1'd1,  5'd21, 27'h00000346, 5'd19, 27'h0000017b, 5'd14, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001d9, 5'd19, 27'h00000278, 5'd23, 27'h00000357, 32'h00000400,
  1'd1,  5'd22, 27'h00000006, 5'd30, 27'h000000ad, 5'd1, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000036d, 5'd29, 27'h000000a5, 5'd15, 27'h000000d9, 32'h00000400,
  1'd1,  5'd21, 27'h000000aa, 5'd30, 27'h00000136, 5'd21, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000368, 5'd5, 27'h00000264, 5'd5, 27'h000001b1, 32'h00000400,
  1'd1,  5'd0, 27'h00000152, 5'd9, 27'h000000c3, 5'd18, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000087, 5'd5, 27'h0000011e, 5'd26, 27'h00000322, 32'h00000400,
  1'd1,  5'd3, 27'h00000158, 5'd17, 27'h0000032b, 5'd8, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000091, 5'd17, 27'h000000a4, 5'd15, 27'h00000336, 32'h00000400,
  1'd1,  5'd4, 27'h0000034b, 5'd18, 27'h000000d4, 5'd29, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003e5, 5'd26, 27'h0000029c, 5'd7, 27'h00000283, 32'h00000400,
  1'd1,  5'd0, 27'h000000d4, 5'd28, 27'h00000170, 5'd19, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000126, 5'd29, 27'h000001a0, 5'd28, 27'h000000d6, 32'h00000400,
  1'd1,  5'd13, 27'h00000173, 5'd7, 27'h00000022, 5'd7, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000173, 5'd5, 27'h0000014b, 5'd20, 27'h00000030, 32'h00000400,
  1'd1,  5'd12, 27'h00000303, 5'd6, 27'h000001df, 5'd27, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000281, 5'd17, 27'h000000c4, 5'd8, 27'h00000370, 32'h00000400,
  1'd1,  5'd10, 27'h000003f0, 5'd17, 27'h00000286, 5'd17, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002cf, 5'd17, 27'h00000389, 5'd30, 27'h00000168, 32'h00000400,
  1'd1,  5'd11, 27'h000002db, 5'd28, 27'h000002eb, 5'd7, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000167, 5'd30, 27'h000001b3, 5'd17, 27'h00000160, 32'h00000400,
  1'd1,  5'd10, 27'h000002bc, 5'd28, 27'h00000270, 5'd25, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000039, 5'd6, 27'h0000013a, 5'd6, 27'h0000037c, 32'h00000400,
  1'd1,  5'd25, 27'h000001cb, 5'd8, 27'h0000001d, 5'd19, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000069, 5'd7, 27'h00000189, 5'd30, 27'h000000f8, 32'h00000400,
  1'd1,  5'd25, 27'h00000154, 5'd16, 27'h00000152, 5'd6, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000136, 5'd18, 27'h0000018b, 5'd17, 27'h00000230, 32'h00000400,
  1'd1,  5'd24, 27'h00000263, 5'd20, 27'h0000004f, 5'd26, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000031e, 5'd29, 27'h0000021a, 5'd7, 27'h0000014e, 32'h00000400,
  1'd1,  5'd23, 27'h0000022b, 5'd26, 27'h00000372, 5'd16, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002cc, 5'd26, 27'h0000023d, 5'd30, 27'h00000029, 32'h00000400,
  1'd1,  5'd9, 27'h000003e3, 5'd2, 27'h000000a3, 5'd9, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000016, 5'd3, 27'h000003ea, 5'd20, 27'h00000183, 32'h00000400,
  1'd1,  5'd9, 27'h00000333, 5'd4, 27'h0000018e, 5'd29, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ea, 5'd10, 27'h000001cf, 5'd3, 27'h000002f7, 32'h00000400,
  1'd1,  5'd8, 27'h00000005, 5'd11, 27'h000000c0, 5'd13, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b5, 5'd14, 27'h000001c5, 5'd22, 27'h00000376, 32'h00000400,
  1'd1,  5'd9, 27'h0000032a, 5'd25, 27'h0000009e, 5'd4, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000035f, 5'd21, 27'h000003ff, 5'd12, 27'h0000016a, 32'h00000400,
  1'd1,  5'd7, 27'h000001d6, 5'd23, 27'h0000020d, 5'd21, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f2, 5'd4, 27'h000003b5, 5'd9, 27'h0000015c, 32'h00000400,
  1'd1,  5'd17, 27'h000003d7, 5'd1, 27'h000000f3, 5'd16, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000019e, 5'd4, 27'h0000033e, 5'd26, 27'h00000086, 32'h00000400,
  1'd1,  5'd19, 27'h0000017e, 5'd13, 27'h0000038f, 5'd4, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000160, 5'd12, 27'h000002b3, 5'd13, 27'h0000035c, 32'h00000400,
  1'd1,  5'd15, 27'h000003a3, 5'd12, 27'h000000f7, 5'd21, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000253, 5'd25, 27'h000000e5, 5'd2, 27'h00000153, 32'h00000400,
  1'd1,  5'd19, 27'h00000347, 5'd25, 27'h000000f9, 5'd12, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000013a, 5'd23, 27'h00000014, 5'd24, 27'h00000310, 32'h00000400,
  1'd1,  5'd25, 27'h00000364, 5'd3, 27'h000000e1, 5'd0, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000025, 5'd5, 27'h00000046, 5'd14, 27'h000003b9, 32'h00000400,
  1'd1,  5'd27, 27'h000001d4, 5'd3, 27'h00000052, 5'd23, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000012f, 5'd12, 27'h000001f8, 5'd4, 27'h00000305, 32'h00000400,
  1'd1,  5'd29, 27'h00000110, 5'd14, 27'h000002fe, 5'd10, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f4, 5'd14, 27'h00000361, 5'd25, 27'h000002ab, 32'h00000400,
  1'd1,  5'd28, 27'h00000202, 5'd23, 27'h00000173, 5'd3, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000036a, 5'd21, 27'h00000308, 5'd10, 27'h000003e4, 32'h00000400,
  1'd1,  5'd29, 27'h00000099, 5'd24, 27'h00000272, 5'd23, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000028d, 5'd1, 27'h000000c1, 5'd2, 27'h0000000f, 32'h00000400,
  1'd1,  5'd8, 27'h0000030a, 5'd3, 27'h000003e3, 5'd13, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000022b, 5'd2, 27'h000001f9, 5'd23, 27'h000000b5, 32'h00000400,
  1'd1,  5'd5, 27'h0000012d, 5'd14, 27'h0000028b, 5'd9, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e5, 5'd14, 27'h0000038b, 5'd19, 27'h000000cb, 32'h00000400,
  1'd1,  5'd8, 27'h00000357, 5'd15, 27'h000000ff, 5'd29, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002fa, 5'd21, 27'h0000017c, 5'd5, 27'h000001af, 32'h00000400,
  1'd1,  5'd6, 27'h00000048, 5'd23, 27'h00000188, 5'd19, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000354, 5'd25, 27'h00000235, 5'd30, 27'h0000026c, 32'h00000400,
  1'd1,  5'd19, 27'h0000014b, 5'd3, 27'h000003c2, 5'd0, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000023d, 5'd4, 27'h00000384, 5'd15, 27'h00000171, 32'h00000400,
  1'd1,  5'd18, 27'h0000003f, 5'd2, 27'h0000032a, 5'd23, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f4, 5'd12, 27'h000000d8, 5'd7, 27'h0000038a, 32'h00000400,
  1'd1,  5'd18, 27'h000003a4, 5'd12, 27'h000002cc, 5'd17, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ae, 5'd13, 27'h000001da, 5'd29, 27'h00000083, 32'h00000400,
  1'd1,  5'd17, 27'h00000164, 5'd25, 27'h000001ad, 5'd9, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d7, 5'd22, 27'h000000c1, 5'd19, 27'h00000018, 32'h00000400,
  1'd1,  5'd16, 27'h00000124, 5'd23, 27'h0000029a, 5'd29, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a3, 5'd4, 27'h00000235, 5'd10, 27'h0000012b, 32'h00000400,
  1'd1,  5'd26, 27'h0000003a, 5'd1, 27'h0000028f, 5'd16, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000086, 5'd1, 27'h0000017b, 5'd29, 27'h0000038d, 32'h00000400,
  1'd1,  5'd29, 27'h000003b3, 5'd12, 27'h00000153, 5'd8, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002de, 5'd14, 27'h0000004d, 5'd18, 27'h00000028, 32'h00000400,
  1'd1,  5'd25, 27'h000003ed, 5'd13, 27'h000003d2, 5'd28, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e1, 5'd22, 27'h0000013f, 5'd6, 27'h000003fb, 32'h00000400,
  1'd1,  5'd26, 27'h00000068, 5'd24, 27'h00000126, 5'd17, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000d3, 5'd24, 27'h00000256, 5'd26, 27'h000001a6, 32'h00000400,
  1'd1,  5'd8, 27'h00000167, 5'd9, 27'h000003f2, 5'd1, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000220, 5'd8, 27'h00000381, 5'd10, 27'h0000016c, 32'h00000400,
  1'd1,  5'd8, 27'h0000018c, 5'd9, 27'h00000111, 5'd23, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000224, 5'd18, 27'h0000002e, 5'd2, 27'h0000009e, 32'h00000400,
  1'd1,  5'd6, 27'h000003fb, 5'd20, 27'h000000a4, 5'd10, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000170, 5'd19, 27'h000001a1, 5'd23, 27'h000002cf, 32'h00000400,
  1'd1,  5'd6, 27'h000000aa, 5'd27, 27'h00000383, 5'd1, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c7, 5'd30, 27'h000001b6, 5'd14, 27'h000002c2, 32'h00000400,
  1'd1,  5'd10, 27'h000000a9, 5'd27, 27'h00000240, 5'd24, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e6, 5'd7, 27'h0000006d, 5'd2, 27'h00000040, 32'h00000400,
  1'd1,  5'd18, 27'h00000158, 5'd5, 27'h0000020e, 5'd12, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000008, 5'd6, 27'h000003f1, 5'd24, 27'h0000007a, 32'h00000400,
  1'd1,  5'd19, 27'h00000325, 5'd17, 27'h000003f0, 5'd2, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cd, 5'd16, 27'h0000017a, 5'd14, 27'h00000181, 32'h00000400,
  1'd1,  5'd16, 27'h000003c9, 5'd20, 27'h000000db, 5'd24, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f5, 5'd30, 27'h000002c9, 5'd2, 27'h0000021d, 32'h00000400,
  1'd1,  5'd15, 27'h00000276, 5'd29, 27'h00000239, 5'd15, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cc, 5'd30, 27'h0000022a, 5'd23, 27'h00000249, 32'h00000400,
  1'd1,  5'd29, 27'h00000023, 5'd8, 27'h00000202, 5'd4, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000068, 5'd8, 27'h00000117, 5'd11, 27'h0000007e, 32'h00000400,
  1'd1,  5'd28, 27'h00000261, 5'd9, 27'h000003c9, 5'd24, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000016f, 5'd16, 27'h0000018f, 5'd0, 27'h00000130, 32'h00000400,
  1'd1,  5'd29, 27'h0000006a, 5'd18, 27'h000000d7, 5'd11, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000010f, 5'd20, 27'h00000062, 5'd25, 27'h000002b5, 32'h00000400,
  1'd1,  5'd29, 27'h000003d3, 5'd30, 27'h0000031b, 5'd1, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000e1, 5'd27, 27'h000000f9, 5'd13, 27'h00000393, 32'h00000400,
  1'd1,  5'd30, 27'h0000011d, 5'd30, 27'h000003e4, 5'd24, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000031b, 5'd8, 27'h0000004a, 5'd8, 27'h00000105, 32'h00000400,
  1'd1,  5'd7, 27'h000001c0, 5'd9, 27'h0000009b, 5'd20, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000002b, 5'd8, 27'h000003ba, 5'd26, 27'h000000b7, 32'h00000400,
  1'd1,  5'd5, 27'h00000310, 5'd20, 27'h000000a5, 5'd6, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a1, 5'd16, 27'h000002e7, 5'd18, 27'h000001cd, 32'h00000400,
  1'd1,  5'd8, 27'h000002cd, 5'd17, 27'h00000250, 5'd29, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000029d, 5'd28, 27'h000001e2, 5'd7, 27'h00000084, 32'h00000400,
  1'd1,  5'd5, 27'h000003a5, 5'd29, 27'h000002aa, 5'd18, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cd, 5'd28, 27'h000003c7, 5'd30, 27'h00000018, 32'h00000400,
  1'd1,  5'd16, 27'h0000033a, 5'd6, 27'h000000fe, 5'd8, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002ca, 5'd6, 27'h000002cb, 5'd20, 27'h00000295, 32'h00000400,
  1'd1,  5'd16, 27'h00000248, 5'd5, 27'h0000023f, 5'd29, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000009f, 5'd19, 27'h0000002b, 5'd6, 27'h00000223, 32'h00000400,
  1'd1,  5'd19, 27'h00000298, 5'd18, 27'h00000215, 5'd19, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000020, 5'd20, 27'h00000223, 5'd26, 27'h0000006b, 32'h00000400,
  1'd1,  5'd18, 27'h00000163, 5'd28, 27'h00000308, 5'd9, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ae, 5'd30, 27'h0000009a, 5'd18, 27'h00000148, 32'h00000400,
  1'd1,  5'd19, 27'h000003e3, 5'd26, 27'h0000039c, 5'd30, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d9, 5'd9, 27'h00000079, 5'd10, 27'h000000a4, 32'h00000400,
  1'd1,  5'd27, 27'h0000013c, 5'd7, 27'h00000221, 5'd17, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000008, 5'd10, 27'h00000071, 5'd26, 27'h00000148, 32'h00000400,
  1'd1,  5'd27, 27'h000001bf, 5'd17, 27'h00000107, 5'd9, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b9, 5'd19, 27'h000001a7, 5'd20, 27'h000001df, 32'h00000400,
  1'd1,  5'd28, 27'h00000327, 5'd20, 27'h00000185, 5'd26, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025c, 5'd28, 27'h00000178, 5'd7, 27'h0000039a, 32'h00000400,
  1'd1,  5'd28, 27'h000001ad, 5'd28, 27'h0000002d, 5'd18, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000109, 5'd28, 27'h000003a5, 5'd29, 27'h000000b1, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000387, 5'd2, 27'h000003ca, 5'd1, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f9, 5'd1, 27'h00000358, 5'd11, 27'h0000003b, 32'h00000400,
  1'd1,  5'd4, 27'h000001b5, 5'd3, 27'h0000010a, 5'd25, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e5, 5'd12, 27'h0000037b, 5'd4, 27'h00000111, 32'h00000400,
  1'd1,  5'd1, 27'h000003dc, 5'd11, 27'h000000b9, 5'd10, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000273, 5'd14, 27'h00000382, 5'd25, 27'h0000022c, 32'h00000400,
  1'd1,  5'd1, 27'h000001f6, 5'd22, 27'h000002ed, 5'd4, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b8, 5'd24, 27'h000000d8, 5'd14, 27'h00000069, 32'h00000400,
  1'd1,  5'd0, 27'h00000277, 5'd25, 27'h00000346, 5'd21, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000237, 5'd3, 27'h00000370, 5'd0, 27'h00000092, 32'h00000400,
  1'd1,  5'd13, 27'h00000321, 5'd2, 27'h00000153, 5'd15, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000366, 5'd3, 27'h000001f9, 5'd25, 27'h00000151, 32'h00000400,
  1'd1,  5'd11, 27'h00000212, 5'd13, 27'h000000e4, 5'd3, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000147, 5'd13, 27'h00000248, 5'd10, 27'h00000241, 32'h00000400,
  1'd1,  5'd11, 27'h00000337, 5'd15, 27'h000001a3, 5'd23, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000b3, 5'd20, 27'h0000033f, 5'd1, 27'h00000008, 32'h00000400,
  1'd1,  5'd13, 27'h00000332, 5'd21, 27'h00000122, 5'd13, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000cd, 5'd21, 27'h0000006a, 5'd23, 27'h00000221, 32'h00000400,
  1'd1,  5'd23, 27'h00000011, 5'd1, 27'h000003ae, 5'd4, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002b2, 5'd2, 27'h000000c5, 5'd11, 27'h000003f0, 32'h00000400,
  1'd1,  5'd21, 27'h000000cb, 5'd4, 27'h000003ab, 5'd24, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001db, 5'd13, 27'h000002a7, 5'd4, 27'h0000003d, 32'h00000400,
  1'd1,  5'd21, 27'h00000361, 5'd10, 27'h0000033c, 5'd14, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000127, 5'd14, 27'h00000061, 5'd22, 27'h0000008f, 32'h00000400,
  1'd1,  5'd22, 27'h00000200, 5'd20, 27'h00000389, 5'd3, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000076, 5'd24, 27'h000003c8, 5'd11, 27'h00000121, 32'h00000400,
  1'd1,  5'd23, 27'h000002a0, 5'd23, 27'h0000003f, 5'd24, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000010c, 5'd0, 27'h0000037b, 5'd5, 27'h000003db, 32'h00000400,
  1'd1,  5'd0, 27'h0000023c, 5'd0, 27'h0000018b, 5'd18, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000f7, 5'd4, 27'h000000b7, 5'd28, 27'h000003a9, 32'h00000400,
  1'd1,  5'd1, 27'h00000149, 5'd10, 27'h000003d0, 5'd6, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c2, 5'd11, 27'h000001b0, 5'd16, 27'h00000308, 32'h00000400,
  1'd1,  5'd2, 27'h00000260, 5'd10, 27'h00000182, 5'd28, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000304, 5'd21, 27'h00000096, 5'd6, 27'h00000235, 32'h00000400,
  1'd1,  5'd1, 27'h000002f2, 5'd25, 27'h000002b1, 5'd18, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000357, 5'd20, 27'h0000031e, 5'd27, 27'h00000053, 32'h00000400,
  1'd1,  5'd11, 27'h00000002, 5'd4, 27'h000003eb, 5'd6, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000e8, 5'd2, 27'h0000010e, 5'd16, 27'h00000135, 32'h00000400,
  1'd1,  5'd11, 27'h00000055, 5'd2, 27'h0000028c, 5'd26, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000212, 5'd10, 27'h00000235, 5'd5, 27'h000002f9, 32'h00000400,
  1'd1,  5'd14, 27'h00000045, 5'd12, 27'h00000282, 5'd17, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000310, 5'd14, 27'h000003dc, 5'd28, 27'h000000e2, 32'h00000400,
  1'd1,  5'd10, 27'h00000172, 5'd21, 27'h0000024a, 5'd5, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000267, 5'd23, 27'h00000082, 5'd17, 27'h00000039, 32'h00000400,
  1'd1,  5'd15, 27'h0000015e, 5'd23, 27'h0000002c, 5'd27, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000141, 5'd3, 27'h000002b9, 5'd7, 27'h000000b3, 32'h00000400,
  1'd1,  5'd25, 27'h000000f2, 5'd2, 27'h000000be, 5'd19, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f6, 5'd4, 27'h0000026c, 5'd26, 27'h000001b5, 32'h00000400,
  1'd1,  5'd25, 27'h0000022f, 5'd12, 27'h00000135, 5'd8, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003ba, 5'd10, 27'h000003e7, 5'd17, 27'h000003eb, 32'h00000400,
  1'd1,  5'd21, 27'h0000009a, 5'd13, 27'h000002b2, 5'd28, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000000, 5'd25, 27'h000002d5, 5'd7, 27'h000002b6, 32'h00000400,
  1'd1,  5'd22, 27'h00000316, 5'd23, 27'h00000220, 5'd18, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002c6, 5'd24, 27'h00000400, 5'd30, 27'h00000056, 32'h00000400,
  1'd1,  5'd2, 27'h000001a5, 5'd8, 27'h00000399, 5'd0, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000360, 5'd5, 27'h000002d0, 5'd14, 27'h000002c8, 32'h00000400,
  1'd1,  5'd2, 27'h0000008b, 5'd10, 27'h0000013b, 5'd23, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000208, 5'd17, 27'h00000179, 5'd4, 27'h00000080, 32'h00000400,
  1'd1,  5'd2, 27'h00000299, 5'd18, 27'h00000037, 5'd13, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e4, 5'd17, 27'h0000029f, 5'd22, 27'h000003e9, 32'h00000400,
  1'd1,  5'd2, 27'h000000ef, 5'd30, 27'h000001a1, 5'd2, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000009, 5'd28, 27'h000000df, 5'd11, 27'h0000025c, 32'h00000400,
  1'd1,  5'd0, 27'h00000085, 5'd28, 27'h0000012a, 5'd23, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000015a, 5'd5, 27'h00000226, 5'd5, 27'h000000a1, 32'h00000400,
  1'd1,  5'd12, 27'h00000378, 5'd5, 27'h000003a1, 5'd11, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000357, 5'd8, 27'h000001e6, 5'd24, 27'h000002b1, 32'h00000400,
  1'd1,  5'd15, 27'h0000015d, 5'd16, 27'h000000e5, 5'd2, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001e1, 5'd18, 27'h0000030e, 5'd10, 27'h0000027a, 32'h00000400,
  1'd1,  5'd14, 27'h00000364, 5'd20, 27'h000001d2, 5'd24, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008d, 5'd30, 27'h00000260, 5'd1, 27'h000003fc, 32'h00000400,
  1'd1,  5'd14, 27'h0000026c, 5'd29, 27'h00000246, 5'd14, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034b, 5'd30, 27'h000001ce, 5'd23, 27'h0000024e, 32'h00000400,
  1'd1,  5'd23, 27'h0000020f, 5'd7, 27'h00000238, 5'd0, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fb, 5'd5, 27'h000001fd, 5'd15, 27'h00000034, 32'h00000400,
  1'd1,  5'd23, 27'h00000105, 5'd8, 27'h000003d1, 5'd24, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002cc, 5'd20, 27'h0000014c, 5'd4, 27'h000000ed, 32'h00000400,
  1'd1,  5'd21, 27'h0000001e, 5'd18, 27'h000000fb, 5'd13, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000118, 5'd19, 27'h00000205, 5'd25, 27'h0000002c, 32'h00000400,
  1'd1,  5'd24, 27'h000000a4, 5'd27, 27'h00000198, 5'd3, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000017b, 5'd27, 27'h00000291, 5'd11, 27'h0000008f, 32'h00000400,
  1'd1,  5'd24, 27'h000002d1, 5'd30, 27'h00000127, 5'd21, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000fc, 5'd7, 27'h000002ac, 5'd8, 27'h000000f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000301, 5'd6, 27'h00000141, 5'd16, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000107, 5'd8, 27'h0000010a, 5'd29, 27'h0000019c, 32'h00000400,
  1'd1,  5'd1, 27'h0000032b, 5'd16, 27'h00000275, 5'd10, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000131, 5'd17, 27'h000002a8, 5'd16, 27'h000001e3, 32'h00000400,
  1'd1,  5'd4, 27'h00000189, 5'd15, 27'h000003fa, 5'd29, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000009d, 5'd29, 27'h0000028f, 5'd5, 27'h00000148, 32'h00000400,
  1'd1,  5'd2, 27'h00000181, 5'd25, 27'h000003ba, 5'd17, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000276, 5'd29, 27'h0000027b, 5'd26, 27'h00000358, 32'h00000400,
  1'd1,  5'd13, 27'h00000255, 5'd5, 27'h00000116, 5'd9, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000265, 5'd6, 27'h000002b6, 5'd16, 27'h00000148, 32'h00000400,
  1'd1,  5'd15, 27'h00000110, 5'd9, 27'h00000004, 5'd28, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000009c, 5'd17, 27'h0000031c, 5'd8, 27'h00000210, 32'h00000400,
  1'd1,  5'd11, 27'h0000035d, 5'd16, 27'h00000048, 5'd16, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000af, 5'd15, 27'h0000023f, 5'd27, 27'h00000326, 32'h00000400,
  1'd1,  5'd11, 27'h0000019e, 5'd27, 27'h0000031b, 5'd9, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000036e, 5'd27, 27'h00000028, 5'd16, 27'h00000052, 32'h00000400,
  1'd1,  5'd15, 27'h000001ab, 5'd27, 27'h00000147, 5'd30, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000385, 5'd6, 27'h00000007, 5'd7, 27'h000001a4, 32'h00000400,
  1'd1,  5'd22, 27'h00000084, 5'd5, 27'h00000221, 5'd18, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032e, 5'd5, 27'h000001bc, 5'd27, 27'h000001d5, 32'h00000400,
  1'd1,  5'd25, 27'h000000ff, 5'd16, 27'h00000388, 5'd5, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000073, 5'd17, 27'h00000357, 5'd15, 27'h000003f5, 32'h00000400,
  1'd1,  5'd21, 27'h000000da, 5'd20, 27'h00000180, 5'd30, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000041, 5'd27, 27'h0000038c, 5'd5, 27'h00000140, 32'h00000400,
  1'd1,  5'd24, 27'h000000d2, 5'd27, 27'h00000379, 5'd18, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000015f, 5'd29, 27'h00000273, 5'd29, 27'h0000023e, 32'h00000400,
  1'd1,  5'd9, 27'h00000393, 5'd0, 27'h00000020, 5'd7, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e1, 5'd2, 27'h000002dc, 5'd19, 27'h000002c1, 32'h00000400,
  1'd1,  5'd8, 27'h000003fb, 5'd1, 27'h00000070, 5'd26, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000010d, 5'd13, 27'h000001f6, 5'd4, 27'h000001d8, 32'h00000400,
  1'd1,  5'd9, 27'h000001cf, 5'd10, 27'h00000392, 5'd12, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013e, 5'd13, 27'h000002aa, 5'd25, 27'h000000c2, 32'h00000400,
  1'd1,  5'd6, 27'h00000304, 5'd24, 27'h0000025f, 5'd1, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001dd, 5'd25, 27'h0000012b, 5'd14, 27'h0000029c, 32'h00000400,
  1'd1,  5'd6, 27'h000001fc, 5'd24, 27'h00000059, 5'd23, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002c, 5'd3, 27'h00000125, 5'd9, 27'h00000296, 32'h00000400,
  1'd1,  5'd17, 27'h000003ac, 5'd4, 27'h000002d0, 5'd18, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000081, 5'd1, 27'h0000032b, 5'd30, 27'h000003da, 32'h00000400,
  1'd1,  5'd20, 27'h00000259, 5'd11, 27'h0000030d, 5'd1, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003e4, 5'd15, 27'h000001a0, 5'd14, 27'h0000030c, 32'h00000400,
  1'd1,  5'd16, 27'h00000319, 5'd13, 27'h000002cd, 5'd21, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000019e, 5'd25, 27'h0000015a, 5'd2, 27'h000001e8, 32'h00000400,
  1'd1,  5'd15, 27'h00000263, 5'd23, 27'h00000235, 5'd12, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000016c, 5'd23, 27'h0000010f, 5'd23, 27'h00000039, 32'h00000400,
  1'd1,  5'd28, 27'h000002aa, 5'd3, 27'h000001fd, 5'd2, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e4, 5'd5, 27'h00000090, 5'd10, 27'h000003d1, 32'h00000400,
  1'd1,  5'd29, 27'h00000074, 5'd3, 27'h000003ad, 5'd24, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003aa, 5'd15, 27'h00000109, 5'd5, 27'h00000026, 32'h00000400,
  1'd1,  5'd30, 27'h0000028f, 5'd11, 27'h000003b8, 5'd11, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003cf, 5'd14, 27'h000001c8, 5'd22, 27'h00000304, 32'h00000400,
  1'd1,  5'd30, 27'h0000014e, 5'd22, 27'h00000279, 5'd3, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c0, 5'd21, 27'h000003e3, 5'd12, 27'h000003e8, 32'h00000400,
  1'd1,  5'd30, 27'h0000022c, 5'd24, 27'h000002ea, 5'd23, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003e2, 5'd1, 27'h00000113, 5'd2, 27'h000003ec, 32'h00000400,
  1'd1,  5'd8, 27'h00000365, 5'd2, 27'h0000030c, 5'd13, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002b4, 5'd4, 27'h0000026a, 5'd21, 27'h000001bc, 32'h00000400,
  1'd1,  5'd9, 27'h00000130, 5'd13, 27'h00000207, 5'd7, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000024a, 5'd12, 27'h00000373, 5'd17, 27'h00000210, 32'h00000400,
  1'd1,  5'd6, 27'h000000e7, 5'd12, 27'h000000cc, 5'd26, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002b8, 5'd25, 27'h000002f7, 5'd7, 27'h0000015d, 32'h00000400,
  1'd1,  5'd6, 27'h000001db, 5'd20, 27'h0000030b, 5'd19, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000006f, 5'd21, 27'h0000021f, 5'd25, 27'h000003d8, 32'h00000400,
  1'd1,  5'd15, 27'h000002fe, 5'd2, 27'h00000344, 5'd4, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002bd, 5'd4, 27'h0000017d, 5'd12, 27'h0000018d, 32'h00000400,
  1'd1,  5'd19, 27'h0000037b, 5'd2, 27'h00000131, 5'd23, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000023, 5'd15, 27'h000001d1, 5'd6, 27'h00000287, 32'h00000400,
  1'd1,  5'd16, 27'h00000186, 5'd10, 27'h0000033e, 5'd20, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a9, 5'd13, 27'h0000021b, 5'd30, 27'h00000122, 32'h00000400,
  1'd1,  5'd19, 27'h000001ca, 5'd21, 27'h0000031b, 5'd10, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002a, 5'd24, 27'h0000024d, 5'd20, 27'h000000e5, 32'h00000400,
  1'd1,  5'd20, 27'h00000241, 5'd22, 27'h0000013a, 5'd27, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ab, 5'd1, 27'h00000157, 5'd7, 27'h00000398, 32'h00000400,
  1'd1,  5'd28, 27'h00000364, 5'd0, 27'h000002d5, 5'd17, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000269, 5'd3, 27'h000002f8, 5'd29, 27'h00000065, 32'h00000400,
  1'd1,  5'd27, 27'h0000038b, 5'd12, 27'h000003c6, 5'd8, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000019f, 5'd13, 27'h000003eb, 5'd16, 27'h000003b7, 32'h00000400,
  1'd1,  5'd30, 27'h00000229, 5'd14, 27'h00000332, 5'd28, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c4, 5'd25, 27'h0000016d, 5'd9, 27'h00000095, 32'h00000400,
  1'd1,  5'd26, 27'h00000233, 5'd24, 27'h0000030c, 5'd17, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003bf, 5'd24, 27'h0000009e, 5'd27, 27'h0000010d, 32'h00000400,
  1'd1,  5'd5, 27'h000000ab, 5'd9, 27'h0000028c, 5'd0, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000248, 5'd6, 27'h00000356, 5'd11, 27'h0000001f, 32'h00000400,
  1'd1,  5'd9, 27'h000003f4, 5'd5, 27'h000003b7, 5'd23, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000087, 5'd18, 27'h00000249, 5'd2, 27'h0000035f, 32'h00000400,
  1'd1,  5'd5, 27'h0000010f, 5'd19, 27'h00000356, 5'd14, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002c7, 5'd17, 27'h000002ae, 5'd22, 27'h000003fa, 32'h00000400,
  1'd1,  5'd9, 27'h00000386, 5'd29, 27'h000001dc, 5'd4, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c0, 5'd29, 27'h00000021, 5'd13, 27'h000000d3, 32'h00000400,
  1'd1,  5'd7, 27'h0000035b, 5'd26, 27'h000003f6, 5'd21, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000035, 5'd8, 27'h000001fe, 5'd3, 27'h00000267, 32'h00000400,
  1'd1,  5'd18, 27'h000002a3, 5'd6, 27'h0000026b, 5'd11, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000008c, 5'd7, 27'h000000ae, 5'd22, 27'h00000336, 32'h00000400,
  1'd1,  5'd17, 27'h0000020d, 5'd18, 27'h0000003d, 5'd2, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a7, 5'd20, 27'h0000019a, 5'd12, 27'h0000006a, 32'h00000400,
  1'd1,  5'd18, 27'h000003c7, 5'd17, 27'h000002db, 5'd22, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035e, 5'd27, 27'h0000005e, 5'd0, 27'h000003de, 32'h00000400,
  1'd1,  5'd20, 27'h00000260, 5'd28, 27'h000001dd, 5'd12, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000005d, 5'd30, 27'h0000003a, 5'd22, 27'h00000218, 32'h00000400,
  1'd1,  5'd26, 27'h000000d7, 5'd10, 27'h00000127, 5'd0, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000285, 5'd7, 27'h00000394, 5'd13, 27'h00000300, 32'h00000400,
  1'd1,  5'd29, 27'h000000c7, 5'd7, 27'h0000011d, 5'd22, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e4, 5'd17, 27'h00000068, 5'd2, 27'h00000196, 32'h00000400,
  1'd1,  5'd26, 27'h00000275, 5'd16, 27'h00000114, 5'd15, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f4, 5'd16, 27'h0000036e, 5'd25, 27'h0000021f, 32'h00000400,
  1'd1,  5'd27, 27'h000002d9, 5'd30, 27'h000002c3, 5'd3, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a4, 5'd28, 27'h00000230, 5'd10, 27'h0000023f, 32'h00000400,
  1'd1,  5'd30, 27'h00000136, 5'd29, 27'h0000029b, 5'd20, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000039b, 5'd6, 27'h0000016d, 5'd5, 27'h000001e8, 32'h00000400,
  1'd1,  5'd9, 27'h0000035d, 5'd6, 27'h000000be, 5'd17, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002df, 5'd5, 27'h00000389, 5'd26, 27'h00000210, 32'h00000400,
  1'd1,  5'd7, 27'h00000206, 5'd18, 27'h00000061, 5'd7, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000d8, 5'd16, 27'h000002fd, 5'd15, 27'h000002c6, 32'h00000400,
  1'd1,  5'd7, 27'h000003c3, 5'd19, 27'h000002be, 5'd29, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001bb, 5'd29, 27'h000002e6, 5'd9, 27'h000002bd, 32'h00000400,
  1'd1,  5'd5, 27'h000000fc, 5'd26, 27'h00000183, 5'd17, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000165, 5'd29, 27'h000003e2, 5'd29, 27'h000000ed, 32'h00000400,
  1'd1,  5'd16, 27'h00000237, 5'd10, 27'h00000067, 5'd7, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001f8, 5'd8, 27'h000003ab, 5'd15, 27'h00000232, 32'h00000400,
  1'd1,  5'd17, 27'h00000348, 5'd9, 27'h000002c2, 5'd29, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000282, 5'd17, 27'h00000268, 5'd8, 27'h000000d9, 32'h00000400,
  1'd1,  5'd19, 27'h00000355, 5'd17, 27'h0000001e, 5'd17, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cc, 5'd17, 27'h00000227, 5'd27, 27'h00000065, 32'h00000400,
  1'd1,  5'd19, 27'h0000039a, 5'd26, 27'h0000002b, 5'd6, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000a4, 5'd28, 27'h00000320, 5'd15, 27'h00000377, 32'h00000400,
  1'd1,  5'd17, 27'h0000032f, 5'd30, 27'h00000360, 5'd28, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000bb, 5'd5, 27'h00000171, 5'd5, 27'h0000027f, 32'h00000400,
  1'd1,  5'd28, 27'h00000277, 5'd9, 27'h000003fd, 5'd16, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e8, 5'd6, 27'h00000098, 5'd30, 27'h000003ad, 32'h00000400,
  1'd1,  5'd30, 27'h0000024d, 5'd18, 27'h000001f7, 5'd5, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000002, 5'd19, 27'h00000194, 5'd19, 27'h000001b3, 32'h00000400,
  1'd1,  5'd29, 27'h00000117, 5'd17, 27'h0000000b, 5'd25, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003a1, 5'd28, 27'h000002d9, 5'd6, 27'h000000a4, 32'h00000400,
  1'd1,  5'd27, 27'h0000016d, 5'd30, 27'h000003a0, 5'd18, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000004b, 5'd26, 27'h0000031b, 5'd28, 27'h0000015d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001bc, 5'd4, 27'h00000262, 5'd2, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002d8, 5'd4, 27'h0000037d, 5'd14, 27'h0000035d, 32'h00000400,
  1'd1,  5'd4, 27'h000003e4, 5'd1, 27'h00000043, 5'd23, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000dc, 5'd12, 27'h00000268, 5'd3, 27'h00000049, 32'h00000400,
  1'd1,  5'd4, 27'h00000364, 5'd15, 27'h00000087, 5'd15, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000086, 5'd13, 27'h000003a2, 5'd23, 27'h0000006d, 32'h00000400,
  1'd1,  5'd4, 27'h0000017a, 5'd22, 27'h000003ad, 5'd0, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000218, 5'd22, 27'h0000015c, 5'd14, 27'h000002d6, 32'h00000400,
  1'd1,  5'd3, 27'h00000165, 5'd21, 27'h000000b5, 5'd23, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000171, 5'd2, 27'h0000022a, 5'd3, 27'h00000013, 32'h00000400,
  1'd1,  5'd14, 27'h00000045, 5'd5, 27'h00000012, 5'd10, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d8, 5'd2, 27'h00000363, 5'd24, 27'h000000d0, 32'h00000400,
  1'd1,  5'd15, 27'h0000017c, 5'd13, 27'h0000009e, 5'd4, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000037e, 5'd10, 27'h000001e5, 5'd10, 27'h00000306, 32'h00000400,
  1'd1,  5'd10, 27'h000002b0, 5'd14, 27'h000001e6, 5'd25, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000114, 5'd24, 27'h0000035b, 5'd0, 27'h00000388, 32'h00000400,
  1'd1,  5'd14, 27'h000003a2, 5'd22, 27'h00000019, 5'd10, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000004b, 5'd22, 27'h0000024e, 5'd22, 27'h000002b4, 32'h00000400,
  1'd1,  5'd24, 27'h0000006b, 5'd3, 27'h00000145, 5'd3, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000037a, 5'd3, 27'h000000a3, 5'd14, 27'h000002b3, 32'h00000400,
  1'd1,  5'd24, 27'h000000ae, 5'd4, 27'h00000011, 5'd22, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000005b, 5'd11, 27'h000003a8, 5'd1, 27'h0000017d, 32'h00000400,
  1'd1,  5'd22, 27'h0000026f, 5'd13, 27'h0000027d, 5'd11, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a0, 5'd12, 27'h000000c4, 5'd24, 27'h000000ca, 32'h00000400,
  1'd1,  5'd25, 27'h0000008d, 5'd24, 27'h00000008, 5'd4, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000168, 5'd23, 27'h000001fb, 5'd10, 27'h000001bd, 32'h00000400,
  1'd1,  5'd24, 27'h000002f5, 5'd21, 27'h00000127, 5'd22, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000061, 5'd3, 27'h000002ac, 5'd6, 27'h000002cc, 32'h00000400,
  1'd1,  5'd4, 27'h000002e0, 5'd3, 27'h00000095, 5'd19, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e4, 5'd4, 27'h0000008b, 5'd29, 27'h00000020, 32'h00000400,
  1'd1,  5'd4, 27'h00000341, 5'd13, 27'h00000339, 5'd5, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000361, 5'd12, 27'h000001c1, 5'd18, 27'h000000b8, 32'h00000400,
  1'd1,  5'd1, 27'h000002ca, 5'd10, 27'h000001df, 5'd26, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000009c, 5'd22, 27'h0000004f, 5'd7, 27'h000002fe, 32'h00000400,
  1'd1,  5'd3, 27'h000000fb, 5'd23, 27'h00000378, 5'd16, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000389, 5'd21, 27'h0000005b, 5'd28, 27'h00000227, 32'h00000400,
  1'd1,  5'd13, 27'h00000324, 5'd0, 27'h00000180, 5'd7, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a0, 5'd5, 27'h0000004b, 5'd17, 27'h0000024b, 32'h00000400,
  1'd1,  5'd11, 27'h00000040, 5'd4, 27'h000001d7, 5'd26, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000cc, 5'd10, 27'h000003a7, 5'd9, 27'h00000359, 32'h00000400,
  1'd1,  5'd15, 27'h0000011a, 5'd12, 27'h00000033, 5'd17, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000068, 5'd14, 27'h000002a8, 5'd27, 27'h0000019a, 32'h00000400,
  1'd1,  5'd13, 27'h000000e3, 5'd21, 27'h0000025b, 5'd10, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001fe, 5'd23, 27'h000003ba, 5'd18, 27'h00000316, 32'h00000400,
  1'd1,  5'd13, 27'h0000036a, 5'd25, 27'h00000137, 5'd25, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000373, 5'd2, 27'h0000039d, 5'd7, 27'h00000145, 32'h00000400,
  1'd1,  5'd23, 27'h0000007d, 5'd3, 27'h0000004e, 5'd19, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000233, 5'd4, 27'h0000032c, 5'd29, 27'h000000a2, 32'h00000400,
  1'd1,  5'd25, 27'h0000011d, 5'd14, 27'h00000160, 5'd7, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003be, 5'd12, 27'h000000d5, 5'd16, 27'h000002c2, 32'h00000400,
  1'd1,  5'd24, 27'h000000a9, 5'd12, 27'h0000017b, 5'd29, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000289, 5'd24, 27'h00000251, 5'd8, 27'h000003aa, 32'h00000400,
  1'd1,  5'd25, 27'h0000017d, 5'd24, 27'h00000078, 5'd18, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000261, 5'd23, 27'h00000333, 5'd26, 27'h000001a5, 32'h00000400,
  1'd1,  5'd3, 27'h000000db, 5'd7, 27'h00000049, 5'd3, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000030d, 5'd6, 27'h00000218, 5'd12, 27'h00000315, 32'h00000400,
  1'd1,  5'd0, 27'h000001bf, 5'd5, 27'h00000198, 5'd22, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000054, 5'd16, 27'h0000017a, 5'd3, 27'h00000370, 32'h00000400,
  1'd1,  5'd3, 27'h000001bd, 5'd17, 27'h00000069, 5'd10, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001bc, 5'd18, 27'h000002f3, 5'd24, 27'h000002e4, 32'h00000400,
  1'd1,  5'd2, 27'h00000272, 5'd27, 27'h00000164, 5'd1, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000350, 5'd26, 27'h000002ac, 5'd14, 27'h00000143, 32'h00000400,
  1'd1,  5'd4, 27'h000002da, 5'd27, 27'h00000295, 5'd25, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003db, 5'd6, 27'h000000a4, 5'd2, 27'h00000102, 32'h00000400,
  1'd1,  5'd14, 27'h000002be, 5'd7, 27'h000000a1, 5'd15, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000374, 5'd9, 27'h000000a5, 5'd24, 27'h0000011b, 32'h00000400,
  1'd1,  5'd12, 27'h00000321, 5'd18, 27'h000002a7, 5'd2, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000170, 5'd20, 27'h0000017a, 5'd14, 27'h00000065, 32'h00000400,
  1'd1,  5'd10, 27'h00000337, 5'd18, 27'h0000031d, 5'd24, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000276, 5'd28, 27'h000001b7, 5'd2, 27'h0000026a, 32'h00000400,
  1'd1,  5'd13, 27'h00000380, 5'd30, 27'h00000032, 5'd11, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f0, 5'd30, 27'h0000006c, 5'd21, 27'h000003b8, 32'h00000400,
  1'd1,  5'd25, 27'h0000001e, 5'd7, 27'h00000090, 5'd4, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002cd, 5'd7, 27'h000000e5, 5'd11, 27'h000003ed, 32'h00000400,
  1'd1,  5'd24, 27'h00000250, 5'd9, 27'h000003f8, 5'd24, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000150, 5'd18, 27'h0000019c, 5'd1, 27'h0000021d, 32'h00000400,
  1'd1,  5'd24, 27'h000003eb, 5'd16, 27'h000003d7, 5'd14, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000059, 5'd16, 27'h00000332, 5'd25, 27'h0000011a, 32'h00000400,
  1'd1,  5'd23, 27'h00000308, 5'd29, 27'h00000018, 5'd2, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000336, 5'd27, 27'h0000021d, 5'd12, 27'h00000138, 32'h00000400,
  1'd1,  5'd25, 27'h000000b8, 5'd26, 27'h0000015f, 5'd21, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c1, 5'd8, 27'h0000035b, 5'd9, 27'h00000057, 32'h00000400,
  1'd1,  5'd3, 27'h00000199, 5'd5, 27'h0000039a, 5'd17, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000023f, 5'd5, 27'h000001f6, 5'd28, 27'h00000055, 32'h00000400,
  1'd1,  5'd4, 27'h0000023d, 5'd18, 27'h0000031d, 5'd6, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000378, 5'd19, 27'h0000022c, 5'd19, 27'h0000022d, 32'h00000400,
  1'd1,  5'd4, 27'h0000023b, 5'd16, 27'h00000079, 5'd26, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d4, 5'd27, 27'h000003c2, 5'd5, 27'h0000030a, 32'h00000400,
  1'd1,  5'd1, 27'h000003c9, 5'd28, 27'h00000018, 5'd18, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000023e, 5'd28, 27'h0000019e, 5'd29, 27'h00000335, 32'h00000400,
  1'd1,  5'd14, 27'h000003fc, 5'd9, 27'h00000130, 5'd7, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002c6, 5'd6, 27'h00000288, 5'd20, 27'h000000be, 32'h00000400,
  1'd1,  5'd13, 27'h0000029c, 5'd8, 27'h000002ab, 5'd26, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b0, 5'd18, 27'h00000297, 5'd8, 27'h0000001c, 32'h00000400,
  1'd1,  5'd14, 27'h000003ef, 5'd19, 27'h000000e0, 5'd19, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000199, 5'd19, 27'h000002f1, 5'd29, 27'h000002e1, 32'h00000400,
  1'd1,  5'd15, 27'h000001aa, 5'd26, 27'h00000343, 5'd8, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000293, 5'd29, 27'h000002c4, 5'd18, 27'h00000282, 32'h00000400,
  1'd1,  5'd13, 27'h000000d3, 5'd30, 27'h0000020c, 5'd26, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001e7, 5'd5, 27'h0000029a, 5'd9, 27'h000002ab, 32'h00000400,
  1'd1,  5'd22, 27'h000003cd, 5'd6, 27'h000003f4, 5'd17, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000051, 5'd8, 27'h00000347, 5'd27, 27'h00000002, 32'h00000400,
  1'd1,  5'd22, 27'h00000208, 5'd15, 27'h000003b5, 5'd7, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000032f, 5'd17, 27'h0000037f, 5'd15, 27'h00000343, 32'h00000400,
  1'd1,  5'd22, 27'h000001a5, 5'd20, 27'h0000004a, 5'd30, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000124, 5'd30, 27'h0000002e, 5'd9, 27'h00000044, 32'h00000400,
  1'd1,  5'd22, 27'h000000ff, 5'd28, 27'h000000fd, 5'd19, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000c0, 5'd28, 27'h00000305, 5'd26, 27'h000000f7, 32'h00000400,
  1'd1,  5'd7, 27'h000001f5, 5'd3, 27'h00000000, 5'd9, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000015f, 5'd0, 27'h0000029e, 5'd20, 27'h00000246, 32'h00000400,
  1'd1,  5'd9, 27'h000003e7, 5'd0, 27'h000002cb, 5'd30, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000095, 5'd15, 27'h000001ee, 5'd4, 27'h000001cb, 32'h00000400,
  1'd1,  5'd8, 27'h00000087, 5'd10, 27'h00000353, 5'd14, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002dc, 5'd11, 27'h00000315, 5'd24, 27'h00000143, 32'h00000400,
  1'd1,  5'd7, 27'h00000325, 5'd22, 27'h000001e7, 5'd1, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000c7, 5'd22, 27'h000003c5, 5'd10, 27'h000003f1, 32'h00000400,
  1'd1,  5'd5, 27'h000001b4, 5'd24, 27'h0000023a, 5'd21, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000197, 5'd1, 27'h000000c8, 5'd9, 27'h000000ec, 32'h00000400,
  1'd1,  5'd17, 27'h000001fe, 5'd1, 27'h000000e1, 5'd18, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000024b, 5'd1, 27'h0000002c, 5'd27, 27'h00000006, 32'h00000400,
  1'd1,  5'd20, 27'h0000025e, 5'd12, 27'h00000175, 5'd0, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000025f, 5'd11, 27'h000003ac, 5'd12, 27'h000001de, 32'h00000400,
  1'd1,  5'd20, 27'h00000119, 5'd15, 27'h00000159, 5'd20, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000034b, 5'd24, 27'h0000025d, 5'd0, 27'h000001bb, 32'h00000400,
  1'd1,  5'd20, 27'h0000007f, 5'd23, 27'h000001a7, 5'd13, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f5, 5'd22, 27'h0000015f, 5'd23, 27'h00000183, 32'h00000400,
  1'd1,  5'd26, 27'h00000396, 5'd0, 27'h00000388, 5'd5, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000171, 5'd1, 27'h00000208, 5'd13, 27'h00000337, 32'h00000400,
  1'd1,  5'd26, 27'h00000036, 5'd3, 27'h0000013d, 5'd21, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000372, 5'd13, 27'h0000005e, 5'd0, 27'h00000254, 32'h00000400,
  1'd1,  5'd27, 27'h00000222, 5'd14, 27'h0000003d, 5'd13, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000cf, 5'd12, 27'h00000121, 5'd24, 27'h00000207, 32'h00000400,
  1'd1,  5'd27, 27'h000000da, 5'd21, 27'h0000002a, 5'd5, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000342, 5'd21, 27'h0000017b, 5'd14, 27'h00000180, 32'h00000400,
  1'd1,  5'd27, 27'h0000017d, 5'd23, 27'h000003b1, 5'd22, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000e3, 5'd2, 27'h000003fd, 5'd0, 27'h0000039a, 32'h00000400,
  1'd1,  5'd5, 27'h00000208, 5'd4, 27'h00000306, 5'd10, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000119, 5'd3, 27'h00000151, 5'd22, 27'h000000d5, 32'h00000400,
  1'd1,  5'd6, 27'h00000204, 5'd12, 27'h000002bb, 5'd8, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ed, 5'd10, 27'h00000306, 5'd20, 27'h00000040, 32'h00000400,
  1'd1,  5'd5, 27'h0000039c, 5'd10, 27'h00000247, 5'd25, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002bd, 5'd23, 27'h0000026c, 5'd5, 27'h0000018c, 32'h00000400,
  1'd1,  5'd8, 27'h0000015e, 5'd22, 27'h00000098, 5'd17, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000029, 5'd22, 27'h00000073, 5'd26, 27'h0000024b, 32'h00000400,
  1'd1,  5'd18, 27'h00000190, 5'd0, 27'h000001e3, 5'd2, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002df, 5'd0, 27'h00000108, 5'd12, 27'h00000339, 32'h00000400,
  1'd1,  5'd16, 27'h00000369, 5'd4, 27'h00000290, 5'd24, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000069, 5'd14, 27'h00000247, 5'd7, 27'h000000f9, 32'h00000400,
  1'd1,  5'd18, 27'h0000037c, 5'd13, 27'h00000244, 5'd16, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003ac, 5'd12, 27'h000001b1, 5'd25, 27'h0000039c, 32'h00000400,
  1'd1,  5'd17, 27'h000001e5, 5'd22, 27'h0000019d, 5'd6, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000d0, 5'd21, 27'h0000039e, 5'd19, 27'h0000007e, 32'h00000400,
  1'd1,  5'd18, 27'h0000004f, 5'd25, 27'h000001e7, 5'd30, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003fa, 5'd0, 27'h000001ee, 5'd9, 27'h00000101, 32'h00000400,
  1'd1,  5'd27, 27'h0000028a, 5'd0, 27'h000003e5, 5'd15, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000268, 5'd2, 27'h0000030c, 5'd30, 27'h0000026a, 32'h00000400,
  1'd1,  5'd27, 27'h000003fc, 5'd11, 27'h000001ef, 5'd8, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000038d, 5'd15, 27'h00000059, 5'd19, 27'h00000147, 32'h00000400,
  1'd1,  5'd26, 27'h0000007c, 5'd11, 27'h000000f0, 5'd28, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000028e, 5'd21, 27'h00000223, 5'd9, 27'h0000033c, 32'h00000400,
  1'd1,  5'd29, 27'h00000312, 5'd22, 27'h0000009b, 5'd18, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002ec, 5'd25, 27'h00000061, 5'd29, 27'h00000188, 32'h00000400,
  1'd1,  5'd9, 27'h000003ee, 5'd8, 27'h0000005c, 5'd3, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000112, 5'd5, 27'h000000d7, 5'd15, 27'h000000e8, 32'h00000400,
  1'd1,  5'd9, 27'h000001aa, 5'd6, 27'h0000006a, 5'd24, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000363, 5'd18, 27'h00000390, 5'd3, 27'h000003d5, 32'h00000400,
  1'd1,  5'd5, 27'h00000120, 5'd18, 27'h0000009d, 5'd11, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000119, 5'd19, 27'h000000d6, 5'd24, 27'h000003b6, 32'h00000400,
  1'd1,  5'd9, 27'h000002a7, 5'd28, 27'h000002e4, 5'd3, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000262, 5'd29, 27'h000002cb, 5'd12, 27'h00000208, 32'h00000400,
  1'd1,  5'd8, 27'h0000030f, 5'd28, 27'h00000325, 5'd22, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032a, 5'd9, 27'h00000285, 5'd0, 27'h0000020a, 32'h00000400,
  1'd1,  5'd19, 27'h000000a0, 5'd5, 27'h0000018d, 5'd13, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000014, 5'd6, 27'h0000001b, 5'd24, 27'h000002f0, 32'h00000400,
  1'd1,  5'd20, 27'h000000fd, 5'd18, 27'h0000035f, 5'd0, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ff, 5'd16, 27'h000003f6, 5'd10, 27'h00000392, 32'h00000400,
  1'd1,  5'd20, 27'h00000064, 5'd18, 27'h00000296, 5'd25, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d0, 5'd28, 27'h000003d5, 5'd1, 27'h000002bd, 32'h00000400,
  1'd1,  5'd19, 27'h000000b0, 5'd26, 27'h0000029f, 5'd10, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000242, 5'd28, 27'h0000035b, 5'd25, 27'h00000296, 32'h00000400,
  1'd1,  5'd30, 27'h0000005b, 5'd9, 27'h000001e4, 5'd3, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001e, 5'd7, 27'h00000181, 5'd14, 27'h00000039, 32'h00000400,
  1'd1,  5'd28, 27'h00000290, 5'd8, 27'h00000218, 5'd23, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000020f, 5'd20, 27'h00000215, 5'd4, 27'h0000008c, 32'h00000400,
  1'd1,  5'd28, 27'h00000097, 5'd20, 27'h00000163, 5'd15, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002d1, 5'd19, 27'h000003cc, 5'd23, 27'h000002ab, 32'h00000400,
  1'd1,  5'd30, 27'h00000391, 5'd28, 27'h00000215, 5'd2, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000319, 5'd27, 27'h000001d9, 5'd12, 27'h000002ce, 32'h00000400,
  1'd1,  5'd29, 27'h000003bd, 5'd26, 27'h000000be, 5'd21, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e8, 5'd9, 27'h00000362, 5'd6, 27'h00000125, 32'h00000400,
  1'd1,  5'd6, 27'h000001af, 5'd8, 27'h000000d7, 5'd19, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009e, 5'd6, 27'h00000086, 5'd30, 27'h00000275, 32'h00000400,
  1'd1,  5'd8, 27'h00000088, 5'd18, 27'h00000069, 5'd7, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ea, 5'd18, 27'h00000137, 5'd16, 27'h0000001c, 32'h00000400,
  1'd1,  5'd5, 27'h000000d9, 5'd20, 27'h000001fd, 5'd28, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000f9, 5'd30, 27'h00000095, 5'd8, 27'h000000b0, 32'h00000400,
  1'd1,  5'd6, 27'h00000190, 5'd30, 27'h00000155, 5'd16, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000019e, 5'd30, 27'h00000020, 5'd29, 27'h00000187, 32'h00000400,
  1'd1,  5'd17, 27'h000003a2, 5'd8, 27'h0000030f, 5'd8, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000140, 5'd6, 27'h00000188, 5'd18, 27'h0000003a, 32'h00000400,
  1'd1,  5'd18, 27'h000001f9, 5'd10, 27'h00000010, 5'd26, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a7, 5'd15, 27'h00000253, 5'd5, 27'h0000019c, 32'h00000400,
  1'd1,  5'd18, 27'h000002f7, 5'd15, 27'h000002ce, 5'd18, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000292, 5'd18, 27'h000000df, 5'd28, 27'h000003ae, 32'h00000400,
  1'd1,  5'd19, 27'h000002fe, 5'd30, 27'h0000009e, 5'd6, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001bc, 5'd29, 27'h0000014d, 5'd17, 27'h0000010a, 32'h00000400,
  1'd1,  5'd15, 27'h00000299, 5'd27, 27'h00000115, 5'd26, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002f1, 5'd5, 27'h00000234, 5'd7, 27'h000001cf, 32'h00000400,
  1'd1,  5'd30, 27'h00000248, 5'd7, 27'h00000146, 5'd18, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f7, 5'd9, 27'h00000224, 5'd27, 27'h00000264, 32'h00000400,
  1'd1,  5'd27, 27'h00000071, 5'd16, 27'h00000373, 5'd8, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000011a, 5'd17, 27'h000002be, 5'd17, 27'h0000027e, 32'h00000400,
  1'd1,  5'd28, 27'h000000eb, 5'd20, 27'h0000020c, 5'd29, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000293, 5'd29, 27'h0000018a, 5'd6, 27'h00000169, 32'h00000400,
  1'd1,  5'd29, 27'h00000257, 5'd27, 27'h000001a1, 5'd18, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000036d, 5'd26, 27'h00000305, 5'd30, 27'h00000054, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000003aa, 5'd5, 27'h00000048, 5'd0, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b0, 5'd2, 27'h00000143, 5'd11, 27'h000002ec, 32'h00000400,
  1'd1,  5'd2, 27'h00000133, 5'd1, 27'h000000b9, 5'd21, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000006c, 5'd12, 27'h00000168, 5'd2, 27'h0000002a, 32'h00000400,
  1'd1,  5'd0, 27'h000002e8, 5'd15, 27'h000000a7, 5'd12, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000328, 5'd15, 27'h00000103, 5'd21, 27'h000000bd, 32'h00000400,
  1'd1,  5'd4, 27'h0000013b, 5'd24, 27'h000002d1, 5'd2, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b2, 5'd24, 27'h0000034b, 5'd12, 27'h00000022, 32'h00000400,
  1'd1,  5'd0, 27'h00000248, 5'd21, 27'h00000086, 5'd24, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b5, 5'd2, 27'h000001bf, 5'd3, 27'h00000369, 32'h00000400,
  1'd1,  5'd14, 27'h0000009d, 5'd4, 27'h000003c5, 5'd14, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ff, 5'd1, 27'h000000da, 5'd23, 27'h0000003f, 32'h00000400,
  1'd1,  5'd14, 27'h000001f1, 5'd13, 27'h0000022d, 5'd1, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000194, 5'd15, 27'h00000160, 5'd13, 27'h000001e1, 32'h00000400,
  1'd1,  5'd14, 27'h00000275, 5'd15, 27'h0000000b, 5'd25, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000003e, 5'd25, 27'h00000346, 5'd1, 27'h000003f0, 32'h00000400,
  1'd1,  5'd11, 27'h00000237, 5'd24, 27'h00000126, 5'd11, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003bc, 5'd21, 27'h000002c3, 5'd24, 27'h0000014d, 32'h00000400,
  1'd1,  5'd22, 27'h00000248, 5'd2, 27'h00000212, 5'd3, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000371, 5'd0, 27'h00000221, 5'd14, 27'h000003d8, 32'h00000400,
  1'd1,  5'd22, 27'h000000d1, 5'd0, 27'h0000026d, 5'd21, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000022e, 5'd14, 27'h00000313, 5'd4, 27'h00000301, 32'h00000400,
  1'd1,  5'd24, 27'h00000264, 5'd10, 27'h00000358, 5'd10, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000039b, 5'd10, 27'h000001c4, 5'd24, 27'h0000011d, 32'h00000400,
  1'd1,  5'd24, 27'h000000a7, 5'd25, 27'h000002b6, 5'd1, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fa, 5'd21, 27'h00000200, 5'd14, 27'h00000239, 32'h00000400,
  1'd1,  5'd24, 27'h00000344, 5'd25, 27'h000002e2, 5'd24, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000248, 5'd3, 27'h00000360, 5'd10, 27'h0000005e, 32'h00000400,
  1'd1,  5'd2, 27'h00000242, 5'd3, 27'h0000023b, 5'd18, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c6, 5'd0, 27'h00000181, 5'd29, 27'h00000023, 32'h00000400,
  1'd1,  5'd1, 27'h00000172, 5'd14, 27'h000003c6, 5'd7, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d4, 5'd12, 27'h0000023a, 5'd15, 27'h0000023b, 32'h00000400,
  1'd1,  5'd0, 27'h0000010d, 5'd13, 27'h00000067, 5'd30, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000368, 5'd23, 27'h000000c6, 5'd10, 27'h00000090, 32'h00000400,
  1'd1,  5'd1, 27'h000002a7, 5'd23, 27'h00000179, 5'd16, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fb, 5'd24, 27'h00000037, 5'd30, 27'h000000de, 32'h00000400,
  1'd1,  5'd11, 27'h000003e3, 5'd3, 27'h0000023b, 5'd6, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000019d, 5'd5, 27'h00000014, 5'd15, 27'h00000201, 32'h00000400,
  1'd1,  5'd14, 27'h00000272, 5'd2, 27'h00000287, 5'd28, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001fe, 5'd13, 27'h000000e8, 5'd6, 27'h0000002a, 32'h00000400,
  1'd1,  5'd14, 27'h00000369, 5'd12, 27'h0000014f, 5'd17, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000021b, 5'd13, 27'h00000335, 5'd25, 27'h000003f3, 32'h00000400,
  1'd1,  5'd13, 27'h00000193, 5'd24, 27'h0000002e, 5'd7, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000054, 5'd23, 27'h00000210, 5'd19, 27'h00000091, 32'h00000400,
  1'd1,  5'd11, 27'h00000226, 5'd25, 27'h0000016b, 5'd29, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021e, 5'd1, 27'h0000007c, 5'd9, 27'h000003c2, 32'h00000400,
  1'd1,  5'd25, 27'h0000012e, 5'd0, 27'h0000006b, 5'd19, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d2, 5'd0, 27'h000003bb, 5'd28, 27'h0000021d, 32'h00000400,
  1'd1,  5'd23, 27'h000001c9, 5'd13, 27'h00000094, 5'd8, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002b6, 5'd10, 27'h0000030b, 5'd19, 27'h0000016b, 32'h00000400,
  1'd1,  5'd23, 27'h000000e7, 5'd14, 27'h0000000e, 5'd26, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000027d, 5'd22, 27'h0000006a, 5'd8, 27'h000003e0, 32'h00000400,
  1'd1,  5'd22, 27'h000002aa, 5'd24, 27'h00000173, 5'd18, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000312, 5'd23, 27'h00000292, 5'd28, 27'h00000043, 32'h00000400,
  1'd1,  5'd2, 27'h000001f8, 5'd9, 27'h00000135, 5'd1, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c6, 5'd9, 27'h0000021f, 5'd14, 27'h00000251, 32'h00000400,
  1'd1,  5'd1, 27'h000003cc, 5'd9, 27'h00000235, 5'd23, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000229, 5'd17, 27'h00000105, 5'd4, 27'h000001ed, 32'h00000400,
  1'd1,  5'd1, 27'h00000363, 5'd18, 27'h00000070, 5'd12, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000176, 5'd19, 27'h00000303, 5'd24, 27'h000003e1, 32'h00000400,
  1'd1,  5'd2, 27'h000001d5, 5'd27, 27'h00000257, 5'd0, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000033, 5'd26, 27'h00000074, 5'd13, 27'h00000043, 32'h00000400,
  1'd1,  5'd3, 27'h00000361, 5'd30, 27'h000000f3, 5'd24, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000005f, 5'd9, 27'h000001eb, 5'd3, 27'h000000b6, 32'h00000400,
  1'd1,  5'd11, 27'h0000010a, 5'd8, 27'h00000204, 5'd13, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003df, 5'd5, 27'h00000365, 5'd22, 27'h000003a5, 32'h00000400,
  1'd1,  5'd13, 27'h0000027a, 5'd17, 27'h000001e1, 5'd3, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000139, 5'd20, 27'h0000009f, 5'd15, 27'h00000088, 32'h00000400,
  1'd1,  5'd11, 27'h000001d8, 5'd15, 27'h0000036a, 5'd25, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000052, 5'd28, 27'h000001f4, 5'd4, 27'h000003cc, 32'h00000400,
  1'd1,  5'd14, 27'h00000339, 5'd27, 27'h000003d0, 5'd12, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000287, 5'd27, 27'h00000189, 5'd23, 27'h0000039c, 32'h00000400,
  1'd1,  5'd24, 27'h000002fe, 5'd9, 27'h0000015e, 5'd0, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000179, 5'd6, 27'h0000027e, 5'd12, 27'h000002b5, 32'h00000400,
  1'd1,  5'd24, 27'h000003d4, 5'd7, 27'h000003ab, 5'd23, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001db, 5'd16, 27'h00000199, 5'd4, 27'h00000306, 32'h00000400,
  1'd1,  5'd21, 27'h00000119, 5'd17, 27'h00000061, 5'd10, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000263, 5'd18, 27'h00000302, 5'd23, 27'h0000022d, 32'h00000400,
  1'd1,  5'd24, 27'h00000363, 5'd28, 27'h00000278, 5'd3, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000121, 5'd27, 27'h00000353, 5'd14, 27'h0000034a, 32'h00000400,
  1'd1,  5'd22, 27'h000002b8, 5'd29, 27'h00000240, 5'd21, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000391, 5'd5, 27'h000000b8, 5'd7, 27'h00000309, 32'h00000400,
  1'd1,  5'd1, 27'h00000204, 5'd9, 27'h000001cf, 5'd17, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017f, 5'd8, 27'h00000005, 5'd29, 27'h0000022a, 32'h00000400,
  1'd1,  5'd3, 27'h00000200, 5'd17, 27'h0000006d, 5'd5, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000019, 5'd18, 27'h00000083, 5'd17, 27'h00000267, 32'h00000400,
  1'd1,  5'd3, 27'h000002df, 5'd17, 27'h00000078, 5'd28, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000149, 5'd30, 27'h000003c0, 5'd8, 27'h0000001e, 32'h00000400,
  1'd1,  5'd0, 27'h0000034e, 5'd25, 27'h000003d9, 5'd15, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000026e, 5'd29, 27'h000000ad, 5'd28, 27'h000003af, 32'h00000400,
  1'd1,  5'd11, 27'h0000008a, 5'd7, 27'h00000194, 5'd9, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f8, 5'd8, 27'h00000164, 5'd20, 27'h0000026f, 32'h00000400,
  1'd1,  5'd13, 27'h0000037b, 5'd9, 27'h000002ee, 5'd25, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000369, 5'd16, 27'h00000400, 5'd9, 27'h000001ff, 32'h00000400,
  1'd1,  5'd13, 27'h000001ff, 5'd18, 27'h00000286, 5'd17, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000365, 5'd17, 27'h00000204, 5'd27, 27'h0000004d, 32'h00000400,
  1'd1,  5'd14, 27'h000001f9, 5'd27, 27'h00000380, 5'd7, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000265, 5'd26, 27'h00000333, 5'd17, 27'h000000dd, 32'h00000400,
  1'd1,  5'd10, 27'h000003ea, 5'd28, 27'h0000008b, 5'd28, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002ea, 5'd5, 27'h000000c0, 5'd8, 27'h00000026, 32'h00000400,
  1'd1,  5'd23, 27'h000003b3, 5'd7, 27'h000001bc, 5'd19, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000201, 5'd8, 27'h0000018c, 5'd30, 27'h00000322, 32'h00000400,
  1'd1,  5'd25, 27'h000001ee, 5'd18, 27'h000003b2, 5'd5, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000014a, 5'd16, 27'h0000027c, 5'd19, 27'h0000019b, 32'h00000400,
  1'd1,  5'd21, 27'h000000a7, 5'd17, 27'h000000dc, 5'd26, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000388, 5'd27, 27'h000000c9, 5'd9, 27'h00000232, 32'h00000400,
  1'd1,  5'd25, 27'h00000197, 5'd26, 27'h00000170, 5'd17, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a4, 5'd25, 27'h00000390, 5'd30, 27'h00000196, 32'h00000400,
  1'd1,  5'd10, 27'h00000110, 5'd1, 27'h0000001f, 5'd6, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000013f, 5'd1, 27'h000003f4, 5'd18, 27'h00000138, 32'h00000400,
  1'd1,  5'd7, 27'h000002ad, 5'd3, 27'h000002e9, 5'd27, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001bd, 5'd10, 27'h000003b3, 5'd3, 27'h00000224, 32'h00000400,
  1'd1,  5'd10, 27'h0000000e, 5'd15, 27'h00000128, 5'd15, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000d9, 5'd14, 27'h00000038, 5'd22, 27'h00000119, 32'h00000400,
  1'd1,  5'd7, 27'h00000272, 5'd23, 27'h00000198, 5'd1, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000036d, 5'd24, 27'h000001bc, 5'd15, 27'h0000014a, 32'h00000400,
  1'd1,  5'd6, 27'h000001da, 5'd25, 27'h00000327, 5'd20, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000084, 5'd1, 27'h0000015b, 5'd9, 27'h00000047, 32'h00000400,
  1'd1,  5'd15, 27'h000003c1, 5'd3, 27'h00000199, 5'd18, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000006e, 5'd3, 27'h00000365, 5'd26, 27'h00000224, 32'h00000400,
  1'd1,  5'd15, 27'h000003bb, 5'd14, 27'h0000004b, 5'd2, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039c, 5'd12, 27'h0000030c, 5'd11, 27'h00000079, 32'h00000400,
  1'd1,  5'd16, 27'h000001cd, 5'd12, 27'h0000025f, 5'd22, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000019, 5'd22, 27'h00000302, 5'd0, 27'h00000172, 32'h00000400,
  1'd1,  5'd20, 27'h000001a4, 5'd22, 27'h00000008, 5'd11, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001fb, 5'd22, 27'h00000339, 5'd24, 27'h00000311, 32'h00000400,
  1'd1,  5'd30, 27'h000003f0, 5'd2, 27'h00000032, 5'd0, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002fb, 5'd0, 27'h0000008c, 5'd10, 27'h000001fb, 32'h00000400,
  1'd1,  5'd29, 27'h00000352, 5'd4, 27'h000001f2, 5'd22, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002ee, 5'd14, 27'h00000308, 5'd3, 27'h0000026f, 32'h00000400,
  1'd1,  5'd30, 27'h0000029a, 5'd13, 27'h00000380, 5'd14, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ad, 5'd14, 27'h00000027, 5'd24, 27'h00000374, 32'h00000400,
  1'd1,  5'd30, 27'h0000019d, 5'd20, 27'h0000038a, 5'd0, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ef, 5'd24, 27'h000000ca, 5'd13, 27'h0000005c, 32'h00000400,
  1'd1,  5'd27, 27'h0000006e, 5'd25, 27'h0000001e, 5'd24, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ce, 5'd1, 27'h0000016e, 5'd0, 27'h00000107, 32'h00000400,
  1'd1,  5'd7, 27'h00000263, 5'd3, 27'h0000033f, 5'd14, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000381, 5'd1, 27'h000001e4, 5'd23, 27'h000000a6, 32'h00000400,
  1'd1,  5'd9, 27'h0000012e, 5'd12, 27'h00000174, 5'd9, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000c9, 5'd13, 27'h0000016d, 5'd19, 27'h00000030, 32'h00000400,
  1'd1,  5'd6, 27'h00000260, 5'd12, 27'h000001a6, 5'd26, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002b4, 5'd24, 27'h000001c3, 5'd9, 27'h00000266, 32'h00000400,
  1'd1,  5'd6, 27'h00000057, 5'd23, 27'h000002ff, 5'd17, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000016f, 5'd23, 27'h0000028d, 5'd27, 27'h00000041, 32'h00000400,
  1'd1,  5'd16, 27'h00000369, 5'd4, 27'h000002d3, 5'd3, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000113, 5'd2, 27'h000002d9, 5'd15, 27'h00000178, 32'h00000400,
  1'd1,  5'd20, 27'h00000137, 5'd1, 27'h000001c3, 5'd25, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002fa, 5'd12, 27'h000000c4, 5'd5, 27'h000000be, 32'h00000400,
  1'd1,  5'd19, 27'h00000081, 5'd14, 27'h00000130, 5'd20, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000155, 5'd10, 27'h00000352, 5'd26, 27'h00000009, 32'h00000400,
  1'd1,  5'd17, 27'h0000028e, 5'd21, 27'h000000eb, 5'd7, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000108, 5'd24, 27'h00000100, 5'd17, 27'h0000038e, 32'h00000400,
  1'd1,  5'd16, 27'h00000290, 5'd24, 27'h00000000, 5'd30, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000029f, 5'd4, 27'h00000327, 5'd8, 27'h000000f4, 32'h00000400,
  1'd1,  5'd28, 27'h000003f4, 5'd4, 27'h000003b7, 5'd20, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b9, 5'd1, 27'h00000081, 5'd29, 27'h0000004f, 32'h00000400,
  1'd1,  5'd27, 27'h000000b5, 5'd13, 27'h000003f4, 5'd8, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000008d, 5'd10, 27'h000003c6, 5'd16, 27'h00000209, 32'h00000400,
  1'd1,  5'd26, 27'h000003d4, 5'd11, 27'h000000f1, 5'd28, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000024, 5'd21, 27'h00000108, 5'd5, 27'h000001aa, 32'h00000400,
  1'd1,  5'd26, 27'h000000b0, 5'd24, 27'h00000327, 5'd18, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000026, 5'd22, 27'h00000089, 5'd28, 27'h000000a7, 32'h00000400,
  1'd1,  5'd5, 27'h000002fa, 5'd9, 27'h000003ef, 5'd4, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023d, 5'd9, 27'h00000107, 5'd12, 27'h00000350, 32'h00000400,
  1'd1,  5'd6, 27'h000003ee, 5'd6, 27'h00000029, 5'd25, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003d7, 5'd15, 27'h000003d4, 5'd0, 27'h000001c9, 32'h00000400,
  1'd1,  5'd9, 27'h0000018a, 5'd18, 27'h00000217, 5'd12, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000033, 5'd16, 27'h00000281, 5'd25, 27'h0000031a, 32'h00000400,
  1'd1,  5'd9, 27'h000003ca, 5'd30, 27'h00000041, 5'd2, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003a8, 5'd27, 27'h0000001e, 5'd12, 27'h0000007c, 32'h00000400,
  1'd1,  5'd9, 27'h000002b6, 5'd27, 27'h000002fc, 5'd23, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000226, 5'd5, 27'h00000286, 5'd1, 27'h00000004, 32'h00000400,
  1'd1,  5'd19, 27'h00000142, 5'd6, 27'h0000033c, 5'd12, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000328, 5'd10, 27'h0000010e, 5'd22, 27'h0000004f, 32'h00000400,
  1'd1,  5'd18, 27'h00000375, 5'd18, 27'h00000136, 5'd1, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000104, 5'd16, 27'h00000331, 5'd14, 27'h00000138, 32'h00000400,
  1'd1,  5'd20, 27'h00000151, 5'd16, 27'h00000177, 5'd23, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000085, 5'd28, 27'h00000089, 5'd3, 27'h000000e5, 32'h00000400,
  1'd1,  5'd16, 27'h00000020, 5'd29, 27'h00000296, 5'd11, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000016c, 5'd28, 27'h00000060, 5'd23, 27'h000002b8, 32'h00000400,
  1'd1,  5'd28, 27'h00000082, 5'd6, 27'h00000126, 5'd0, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001bd, 5'd6, 27'h000001f3, 5'd13, 27'h0000026e, 32'h00000400,
  1'd1,  5'd27, 27'h00000180, 5'd6, 27'h00000374, 5'd22, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000213, 5'd20, 27'h000001a6, 5'd3, 27'h00000399, 32'h00000400,
  1'd1,  5'd25, 27'h000003aa, 5'd16, 27'h0000034e, 5'd11, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000029b, 5'd18, 27'h0000002c, 5'd21, 27'h00000207, 32'h00000400,
  1'd1,  5'd27, 27'h00000273, 5'd26, 27'h00000258, 5'd4, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000d2, 5'd30, 27'h0000012c, 5'd11, 27'h000001ac, 32'h00000400,
  1'd1,  5'd26, 27'h000003f8, 5'd26, 27'h00000067, 5'd21, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000e, 5'd9, 27'h0000033b, 5'd9, 27'h000003a0, 32'h00000400,
  1'd1,  5'd8, 27'h0000031e, 5'd9, 27'h00000313, 5'd20, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000323, 5'd9, 27'h00000279, 5'd28, 27'h00000172, 32'h00000400,
  1'd1,  5'd10, 27'h00000119, 5'd19, 27'h00000198, 5'd6, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000e6, 5'd20, 27'h000001f2, 5'd17, 27'h00000022, 32'h00000400,
  1'd1,  5'd6, 27'h000000a2, 5'd18, 27'h0000006e, 5'd28, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000382, 5'd26, 27'h0000031c, 5'd7, 27'h00000216, 32'h00000400,
  1'd1,  5'd5, 27'h000002c9, 5'd30, 27'h000002d9, 5'd19, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000c9, 5'd30, 27'h000000ff, 5'd28, 27'h000002a9, 32'h00000400,
  1'd1,  5'd16, 27'h0000034a, 5'd6, 27'h000003fc, 5'd8, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000091, 5'd9, 27'h000003bb, 5'd15, 27'h0000036a, 32'h00000400,
  1'd1,  5'd15, 27'h00000370, 5'd7, 27'h000000a5, 5'd29, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002c3, 5'd20, 27'h000002a3, 5'd7, 27'h0000034c, 32'h00000400,
  1'd1,  5'd18, 27'h00000397, 5'd20, 27'h00000107, 5'd20, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d7, 5'd18, 27'h0000019a, 5'd29, 27'h0000038f, 32'h00000400,
  1'd1,  5'd18, 27'h000003e6, 5'd29, 27'h0000020a, 5'd7, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001d4, 5'd27, 27'h000003b1, 5'd19, 27'h0000038a, 32'h00000400,
  1'd1,  5'd20, 27'h00000203, 5'd27, 27'h00000391, 5'd25, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001fe, 5'd6, 27'h000003f8, 5'd9, 27'h000003f4, 32'h00000400,
  1'd1,  5'd30, 27'h00000153, 5'd9, 27'h00000144, 5'd19, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007f, 5'd9, 27'h0000034f, 5'd28, 27'h000002d6, 32'h00000400,
  1'd1,  5'd27, 27'h000002c9, 5'd15, 27'h00000307, 5'd9, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007b, 5'd17, 27'h00000396, 5'd20, 27'h000002a4, 32'h00000400,
  1'd1,  5'd28, 27'h00000245, 5'd16, 27'h0000024e, 5'd28, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000170, 5'd26, 27'h00000212, 5'd7, 27'h0000011b, 32'h00000400,
  1'd1,  5'd28, 27'h0000018e, 5'd27, 27'h00000288, 5'd16, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000002e, 5'd27, 27'h000001e6, 5'd26, 27'h000000bb, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000003e7, 5'd3, 27'h00000056, 5'd2, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000086, 5'd1, 27'h00000319, 5'd15, 27'h0000002d, 32'h00000400,
  1'd1,  5'd1, 27'h0000037c, 5'd1, 27'h000001f6, 5'd24, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000fd, 5'd10, 27'h00000292, 5'd4, 27'h000000f2, 32'h00000400,
  1'd1,  5'd0, 27'h00000209, 5'd13, 27'h000002a4, 5'd10, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000047, 5'd10, 27'h000001f0, 5'd20, 27'h000003a0, 32'h00000400,
  1'd1,  5'd1, 27'h0000010d, 5'd21, 27'h0000024d, 5'd3, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000029a, 5'd25, 27'h00000083, 5'd13, 27'h000003b2, 32'h00000400,
  1'd1,  5'd0, 27'h000002e4, 5'd21, 27'h000001ba, 5'd20, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000084, 5'd0, 27'h000001dc, 5'd4, 27'h000003bd, 32'h00000400,
  1'd1,  5'd14, 27'h00000051, 5'd3, 27'h0000039f, 5'd12, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ed, 5'd0, 27'h00000052, 5'd24, 27'h000002e1, 32'h00000400,
  1'd1,  5'd13, 27'h00000103, 5'd14, 27'h000001f1, 5'd5, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038a, 5'd11, 27'h00000241, 5'd10, 27'h000003c0, 32'h00000400,
  1'd1,  5'd14, 27'h0000022c, 5'd10, 27'h000001e0, 5'd24, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000357, 5'd24, 27'h00000348, 5'd2, 27'h00000287, 32'h00000400,
  1'd1,  5'd12, 27'h000001a4, 5'd25, 27'h00000104, 5'd14, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000116, 5'd21, 27'h0000015c, 5'd25, 27'h00000226, 32'h00000400,
  1'd1,  5'd23, 27'h0000034b, 5'd3, 27'h00000046, 5'd4, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000036, 5'd4, 27'h000001b3, 5'd10, 27'h000002b7, 32'h00000400,
  1'd1,  5'd23, 27'h00000257, 5'd1, 27'h00000330, 5'd22, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000037, 5'd11, 27'h000002e9, 5'd0, 27'h000002d7, 32'h00000400,
  1'd1,  5'd21, 27'h0000039a, 5'd12, 27'h000003e1, 5'd11, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000103, 5'd11, 27'h0000010a, 5'd25, 27'h00000247, 32'h00000400,
  1'd1,  5'd21, 27'h00000329, 5'd25, 27'h00000287, 5'd2, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000030c, 5'd22, 27'h00000195, 5'd11, 27'h00000284, 32'h00000400,
  1'd1,  5'd24, 27'h00000028, 5'd25, 27'h000001c2, 5'd20, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000213, 5'd3, 27'h000001c0, 5'd6, 27'h000002d9, 32'h00000400,
  1'd1,  5'd2, 27'h0000021f, 5'd1, 27'h00000031, 5'd18, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000bd, 5'd4, 27'h000003cc, 5'd28, 27'h000002a4, 32'h00000400,
  1'd1,  5'd3, 27'h000001fb, 5'd12, 27'h0000037e, 5'd5, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000ac, 5'd12, 27'h000000d5, 5'd17, 27'h00000271, 32'h00000400,
  1'd1,  5'd0, 27'h000002d9, 5'd11, 27'h000003b6, 5'd28, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000073, 5'd21, 27'h0000026e, 5'd6, 27'h00000042, 32'h00000400,
  1'd1,  5'd5, 27'h000000a6, 5'd23, 27'h00000089, 5'd16, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a7, 5'd23, 27'h00000156, 5'd27, 27'h00000310, 32'h00000400,
  1'd1,  5'd14, 27'h0000019e, 5'd2, 27'h00000147, 5'd5, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000235, 5'd4, 27'h0000019a, 5'd19, 27'h00000080, 32'h00000400,
  1'd1,  5'd13, 27'h00000376, 5'd4, 27'h000000de, 5'd26, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000076, 5'd13, 27'h0000011c, 5'd8, 27'h00000366, 32'h00000400,
  1'd1,  5'd12, 27'h000000d9, 5'd14, 27'h00000192, 5'd20, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000161, 5'd12, 27'h00000302, 5'd27, 27'h0000035b, 32'h00000400,
  1'd1,  5'd12, 27'h000000e1, 5'd24, 27'h00000004, 5'd8, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002a6, 5'd21, 27'h00000376, 5'd17, 27'h00000169, 32'h00000400,
  1'd1,  5'd11, 27'h0000001b, 5'd24, 27'h000001e0, 5'd26, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000387, 5'd1, 27'h000003e1, 5'd10, 27'h0000013a, 32'h00000400,
  1'd1,  5'd22, 27'h0000011f, 5'd2, 27'h00000119, 5'd18, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001cf, 5'd0, 27'h0000004f, 5'd26, 27'h000001e3, 32'h00000400,
  1'd1,  5'd23, 27'h0000035d, 5'd13, 27'h0000002b, 5'd7, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000262, 5'd10, 27'h0000028b, 5'd17, 27'h00000220, 32'h00000400,
  1'd1,  5'd24, 27'h000000d8, 5'd14, 27'h000000bc, 5'd26, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000367, 5'd23, 27'h0000016d, 5'd7, 27'h0000035e, 32'h00000400,
  1'd1,  5'd23, 27'h000000d6, 5'd22, 27'h00000276, 5'd20, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000286, 5'd23, 27'h00000257, 5'd29, 27'h000002c1, 32'h00000400,
  1'd1,  5'd3, 27'h000003c3, 5'd5, 27'h000003c3, 5'd4, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000025, 5'd5, 27'h00000270, 5'd14, 27'h00000211, 32'h00000400,
  1'd1,  5'd3, 27'h0000030a, 5'd8, 27'h000003db, 5'd21, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000320, 5'd19, 27'h0000009d, 5'd1, 27'h00000230, 32'h00000400,
  1'd1,  5'd3, 27'h000001f6, 5'd16, 27'h000003bd, 5'd11, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000032c, 5'd15, 27'h00000266, 5'd22, 27'h000003fc, 32'h00000400,
  1'd1,  5'd3, 27'h00000195, 5'd28, 27'h0000007c, 5'd0, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a8, 5'd29, 27'h000002d1, 5'd11, 27'h000000e1, 32'h00000400,
  1'd1,  5'd3, 27'h00000325, 5'd30, 27'h000001ef, 5'd25, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000083, 5'd6, 27'h0000022d, 5'd0, 27'h00000129, 32'h00000400,
  1'd1,  5'd13, 27'h000003b7, 5'd7, 27'h000002ca, 5'd13, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002d6, 5'd5, 27'h000002be, 5'd21, 27'h00000014, 32'h00000400,
  1'd1,  5'd11, 27'h000001fc, 5'd15, 27'h000002d5, 5'd3, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000125, 5'd20, 27'h0000024b, 5'd10, 27'h0000034a, 32'h00000400,
  1'd1,  5'd10, 27'h0000021d, 5'd18, 27'h0000027c, 5'd22, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008c, 5'd30, 27'h0000010f, 5'd4, 27'h000000b3, 32'h00000400,
  1'd1,  5'd14, 27'h0000027f, 5'd30, 27'h00000390, 5'd14, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000019b, 5'd29, 27'h000000a2, 5'd21, 27'h00000183, 32'h00000400,
  1'd1,  5'd22, 27'h00000057, 5'd8, 27'h00000167, 5'd0, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a6, 5'd8, 27'h000000b8, 5'd14, 27'h00000111, 32'h00000400,
  1'd1,  5'd22, 27'h000001b8, 5'd6, 27'h00000336, 5'd22, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000236, 5'd16, 27'h00000211, 5'd1, 27'h000001cd, 32'h00000400,
  1'd1,  5'd25, 27'h00000232, 5'd19, 27'h00000248, 5'd13, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000019f, 5'd20, 27'h00000286, 5'd24, 27'h000003cb, 32'h00000400,
  1'd1,  5'd23, 27'h000003f6, 5'd27, 27'h000001df, 5'd2, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000024, 5'd30, 27'h0000035b, 5'd14, 27'h00000098, 32'h00000400,
  1'd1,  5'd25, 27'h000000e2, 5'd28, 27'h00000037, 5'd25, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002fe, 5'd10, 27'h000000a9, 5'd5, 27'h0000020e, 32'h00000400,
  1'd1,  5'd0, 27'h000002cb, 5'd7, 27'h00000392, 5'd15, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000065, 5'd8, 27'h000000f9, 5'd29, 27'h000002e2, 32'h00000400,
  1'd1,  5'd2, 27'h00000397, 5'd20, 27'h00000044, 5'd9, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002c3, 5'd18, 27'h00000263, 5'd16, 27'h00000069, 32'h00000400,
  1'd1,  5'd1, 27'h00000251, 5'd17, 27'h000003fc, 5'd30, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f9, 5'd26, 27'h00000322, 5'd6, 27'h0000001f, 32'h00000400,
  1'd1,  5'd2, 27'h0000034f, 5'd26, 27'h000002e8, 5'd16, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e5, 5'd29, 27'h000003a9, 5'd30, 27'h00000077, 32'h00000400,
  1'd1,  5'd13, 27'h0000038c, 5'd9, 27'h00000263, 5'd6, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000003f, 5'd6, 27'h00000012, 5'd19, 27'h000003be, 32'h00000400,
  1'd1,  5'd15, 27'h000001fd, 5'd6, 27'h00000012, 5'd28, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e8, 5'd16, 27'h000000f1, 5'd7, 27'h000001ce, 32'h00000400,
  1'd1,  5'd10, 27'h0000035b, 5'd19, 27'h00000245, 5'd18, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c6, 5'd15, 27'h000003c6, 5'd28, 27'h00000161, 32'h00000400,
  1'd1,  5'd11, 27'h000002a5, 5'd29, 27'h00000339, 5'd9, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a7, 5'd29, 27'h00000136, 5'd18, 27'h0000026e, 32'h00000400,
  1'd1,  5'd14, 27'h00000220, 5'd25, 27'h00000377, 5'd29, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001ea, 5'd8, 27'h000002ad, 5'd6, 27'h00000057, 32'h00000400,
  1'd1,  5'd23, 27'h00000290, 5'd6, 27'h0000015f, 5'd17, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ba, 5'd5, 27'h00000360, 5'd26, 27'h000002a9, 32'h00000400,
  1'd1,  5'd22, 27'h00000102, 5'd16, 27'h000001b8, 5'd9, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000025d, 5'd20, 27'h000000a8, 5'd20, 27'h000000b3, 32'h00000400,
  1'd1,  5'd23, 27'h00000134, 5'd16, 27'h0000005a, 5'd27, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f0, 5'd27, 27'h0000006e, 5'd5, 27'h000002d8, 32'h00000400,
  1'd1,  5'd22, 27'h00000350, 5'd27, 27'h0000019a, 5'd16, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022f, 5'd27, 27'h00000188, 5'd29, 27'h00000174, 32'h00000400,
  1'd1,  5'd8, 27'h00000070, 5'd4, 27'h00000270, 5'd6, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000029, 5'd0, 27'h000002c0, 5'd16, 27'h00000325, 32'h00000400,
  1'd1,  5'd10, 27'h00000143, 5'd3, 27'h000003d3, 5'd27, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a4, 5'd14, 27'h0000007d, 5'd2, 27'h00000261, 32'h00000400,
  1'd1,  5'd6, 27'h00000306, 5'd13, 27'h000001e4, 5'd14, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000080, 5'd14, 27'h0000018a, 5'd22, 27'h000003ef, 32'h00000400,
  1'd1,  5'd5, 27'h00000235, 5'd23, 27'h000001fa, 5'd4, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d4, 5'd21, 27'h000000f8, 5'd14, 27'h000002ec, 32'h00000400,
  1'd1,  5'd7, 27'h00000388, 5'd24, 27'h000002e3, 5'd24, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000028f, 5'd3, 27'h000001ba, 5'd6, 27'h000002e8, 32'h00000400,
  1'd1,  5'd19, 27'h00000162, 5'd0, 27'h0000015f, 5'd17, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035b, 5'd2, 27'h0000025d, 5'd27, 27'h000003e2, 32'h00000400,
  1'd1,  5'd20, 27'h0000000e, 5'd14, 27'h000002d3, 5'd3, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000305, 5'd13, 27'h0000039d, 5'd14, 27'h0000037a, 32'h00000400,
  1'd1,  5'd20, 27'h00000169, 5'd13, 27'h00000345, 5'd21, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000046, 5'd23, 27'h000001f1, 5'd2, 27'h000001c7, 32'h00000400,
  1'd1,  5'd16, 27'h000003a0, 5'd21, 27'h000001e2, 5'd13, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000240, 5'd25, 27'h000002a9, 5'd24, 27'h000002ea, 32'h00000400,
  1'd1,  5'd27, 27'h000001da, 5'd5, 27'h00000019, 5'd0, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000034b, 5'd1, 27'h00000262, 5'd11, 27'h0000032a, 32'h00000400,
  1'd1,  5'd27, 27'h00000179, 5'd2, 27'h000003a6, 5'd21, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000129, 5'd13, 27'h0000019f, 5'd1, 27'h000001bb, 32'h00000400,
  1'd1,  5'd28, 27'h000001eb, 5'd15, 27'h000000c4, 5'd11, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000037c, 5'd11, 27'h00000046, 5'd21, 27'h000002d9, 32'h00000400,
  1'd1,  5'd30, 27'h00000072, 5'd22, 27'h0000021b, 5'd3, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007b, 5'd21, 27'h000000cd, 5'd15, 27'h00000184, 32'h00000400,
  1'd1,  5'd30, 27'h000003dc, 5'd22, 27'h00000045, 5'd22, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ea, 5'd3, 27'h000002d4, 5'd3, 27'h000000fe, 32'h00000400,
  1'd1,  5'd8, 27'h00000228, 5'd3, 27'h00000071, 5'd14, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000fa, 5'd0, 27'h0000017f, 5'd22, 27'h00000254, 32'h00000400,
  1'd1,  5'd6, 27'h0000023d, 5'd12, 27'h000001dc, 5'd7, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000039c, 5'd13, 27'h000000d0, 5'd18, 27'h0000032f, 32'h00000400,
  1'd1,  5'd8, 27'h00000044, 5'd15, 27'h000000d1, 5'd26, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000126, 5'd23, 27'h00000020, 5'd7, 27'h00000021, 32'h00000400,
  1'd1,  5'd6, 27'h000002ef, 5'd23, 27'h000002cc, 5'd18, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000337, 5'd21, 27'h00000142, 5'd26, 27'h00000270, 32'h00000400,
  1'd1,  5'd17, 27'h000003c0, 5'd4, 27'h000002da, 5'd2, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ea, 5'd3, 27'h00000352, 5'd10, 27'h0000026b, 32'h00000400,
  1'd1,  5'd20, 27'h00000027, 5'd0, 27'h00000186, 5'd21, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000074, 5'd12, 27'h000000d1, 5'd10, 27'h000000f4, 32'h00000400,
  1'd1,  5'd16, 27'h000002ac, 5'd12, 27'h00000155, 5'd19, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000055, 5'd12, 27'h00000279, 5'd27, 27'h000001b0, 32'h00000400,
  1'd1,  5'd18, 27'h000003fa, 5'd25, 27'h0000002e, 5'd6, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e7, 5'd23, 27'h0000015a, 5'd15, 27'h00000348, 32'h00000400,
  1'd1,  5'd20, 27'h0000002c, 5'd23, 27'h000003aa, 5'd29, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036a, 5'd0, 27'h0000024d, 5'd10, 27'h00000109, 32'h00000400,
  1'd1,  5'd27, 27'h00000161, 5'd0, 27'h000000cc, 5'd20, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000015e, 5'd4, 27'h000001db, 5'd28, 27'h000003f1, 32'h00000400,
  1'd1,  5'd26, 27'h0000001a, 5'd11, 27'h000001b0, 5'd5, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ed, 5'd13, 27'h0000001e, 5'd19, 27'h000002f9, 32'h00000400,
  1'd1,  5'd30, 27'h00000054, 5'd13, 27'h00000285, 5'd26, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c7, 5'd20, 27'h00000361, 5'd5, 27'h000001a7, 32'h00000400,
  1'd1,  5'd30, 27'h00000285, 5'd21, 27'h0000029e, 5'd17, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000031e, 5'd23, 27'h000000e2, 5'd26, 27'h000001ca, 32'h00000400,
  1'd1,  5'd5, 27'h0000010c, 5'd8, 27'h00000346, 5'd2, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000039d, 5'd6, 27'h0000019d, 5'd12, 27'h0000025d, 32'h00000400,
  1'd1,  5'd5, 27'h00000378, 5'd9, 27'h00000289, 5'd20, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a7, 5'd16, 27'h000003fc, 5'd0, 27'h000003f4, 32'h00000400,
  1'd1,  5'd9, 27'h0000009d, 5'd20, 27'h00000024, 5'd11, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000004, 5'd20, 27'h00000017, 5'd25, 27'h000001ba, 32'h00000400,
  1'd1,  5'd7, 27'h000000e4, 5'd27, 27'h000003fd, 5'd1, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000023, 5'd27, 27'h00000022, 5'd11, 27'h0000001c, 32'h00000400,
  1'd1,  5'd7, 27'h0000007b, 5'd30, 27'h0000031d, 5'd24, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000324, 5'd8, 27'h0000031b, 5'd4, 27'h00000375, 32'h00000400,
  1'd1,  5'd17, 27'h00000019, 5'd6, 27'h0000021c, 5'd13, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d8, 5'd7, 27'h00000084, 5'd24, 27'h0000005b, 32'h00000400,
  1'd1,  5'd17, 27'h00000331, 5'd19, 27'h00000052, 5'd1, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000363, 5'd17, 27'h0000018a, 5'd14, 27'h00000202, 32'h00000400,
  1'd1,  5'd16, 27'h00000105, 5'd17, 27'h00000029, 5'd21, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000034f, 5'd25, 27'h000003a7, 5'd2, 27'h0000031f, 32'h00000400,
  1'd1,  5'd18, 27'h000001b3, 5'd27, 27'h0000000e, 5'd11, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000293, 5'd29, 27'h00000390, 5'd24, 27'h000003a6, 32'h00000400,
  1'd1,  5'd28, 27'h00000045, 5'd8, 27'h00000280, 5'd3, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000283, 5'd9, 27'h00000381, 5'd14, 27'h0000003c, 32'h00000400,
  1'd1,  5'd27, 27'h00000155, 5'd7, 27'h00000187, 5'd23, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000032c, 5'd17, 27'h0000030c, 5'd4, 27'h0000028d, 32'h00000400,
  1'd1,  5'd28, 27'h0000005e, 5'd17, 27'h000001eb, 5'd11, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000010, 5'd19, 27'h000002ef, 5'd21, 27'h00000017, 32'h00000400,
  1'd1,  5'd29, 27'h00000332, 5'd30, 27'h000001ae, 5'd2, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000002c, 5'd26, 27'h00000233, 5'd15, 27'h0000008d, 32'h00000400,
  1'd1,  5'd28, 27'h0000026c, 5'd27, 27'h00000023, 5'd20, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a2, 5'd7, 27'h0000018f, 5'd6, 27'h000003b4, 32'h00000400,
  1'd1,  5'd7, 27'h00000364, 5'd7, 27'h000000e7, 5'd17, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002bf, 5'd7, 27'h0000027c, 5'd30, 27'h0000036f, 32'h00000400,
  1'd1,  5'd8, 27'h000001b8, 5'd16, 27'h00000170, 5'd10, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000010b, 5'd15, 27'h000003b3, 5'd20, 27'h000000bf, 32'h00000400,
  1'd1,  5'd8, 27'h00000180, 5'd17, 27'h000001b1, 5'd30, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d0, 5'd26, 27'h0000028b, 5'd7, 27'h00000257, 32'h00000400,
  1'd1,  5'd7, 27'h00000114, 5'd30, 27'h000001e9, 5'd15, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009c, 5'd29, 27'h00000024, 5'd27, 27'h00000184, 32'h00000400,
  1'd1,  5'd16, 27'h000003c8, 5'd5, 27'h000001da, 5'd5, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000097, 5'd6, 27'h000000aa, 5'd18, 27'h0000009e, 32'h00000400,
  1'd1,  5'd18, 27'h000003f1, 5'd8, 27'h000001d7, 5'd27, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000319, 5'd19, 27'h000002ec, 5'd8, 27'h000001ae, 32'h00000400,
  1'd1,  5'd19, 27'h00000310, 5'd18, 27'h000001a9, 5'd19, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000206, 5'd16, 27'h0000037a, 5'd27, 27'h00000101, 32'h00000400,
  1'd1,  5'd19, 27'h00000022, 5'd26, 27'h00000136, 5'd9, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000312, 5'd27, 27'h000003b9, 5'd15, 27'h00000337, 32'h00000400,
  1'd1,  5'd18, 27'h00000073, 5'd26, 27'h00000268, 5'd26, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000035e, 5'd8, 27'h000000d0, 5'd8, 27'h0000033c, 32'h00000400,
  1'd1,  5'd29, 27'h000002fa, 5'd7, 27'h000003e7, 5'd17, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003ac, 5'd5, 27'h000002b3, 5'd27, 27'h000001ae, 32'h00000400,
  1'd1,  5'd28, 27'h0000036a, 5'd19, 27'h0000002c, 5'd9, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000022b, 5'd16, 27'h00000370, 5'd16, 27'h000003f7, 32'h00000400,
  1'd1,  5'd26, 27'h000000b9, 5'd18, 27'h0000021d, 5'd28, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000a9, 5'd25, 27'h000003bc, 5'd6, 27'h000003e5, 32'h00000400,
  1'd1,  5'd26, 27'h00000028, 5'd26, 27'h00000075, 5'd17, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000357, 5'd26, 27'h00000173, 5'd26, 27'h00000116, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000146, 5'd4, 27'h00000348, 5'd3, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000326, 5'd0, 27'h00000073, 5'd11, 27'h000001f8, 32'h00000400,
  1'd1,  5'd3, 27'h000001c7, 5'd0, 27'h00000260, 5'd22, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000220, 5'd14, 27'h00000189, 5'd0, 27'h00000109, 32'h00000400,
  1'd1,  5'd2, 27'h000001c3, 5'd11, 27'h00000246, 5'd12, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000216, 5'd13, 27'h0000007b, 5'd22, 27'h0000030a, 32'h00000400,
  1'd1,  5'd1, 27'h000001f8, 5'd23, 27'h000000d7, 5'd2, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000023d, 5'd23, 27'h000001e8, 5'd13, 27'h0000020d, 32'h00000400,
  1'd1,  5'd3, 27'h0000029f, 5'd24, 27'h000003d3, 5'd23, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f7, 5'd2, 27'h0000001f, 5'd2, 27'h00000292, 32'h00000400,
  1'd1,  5'd10, 27'h000002fc, 5'd3, 27'h0000008b, 5'd12, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003aa, 5'd1, 27'h00000048, 5'd23, 27'h000003c7, 32'h00000400,
  1'd1,  5'd11, 27'h000002d7, 5'd13, 27'h00000017, 5'd1, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011f, 5'd13, 27'h000001f9, 5'd11, 27'h000002cf, 32'h00000400,
  1'd1,  5'd10, 27'h000003b5, 5'd12, 27'h000003a1, 5'd24, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035e, 5'd20, 27'h0000039c, 5'd4, 27'h0000013b, 32'h00000400,
  1'd1,  5'd15, 27'h000000c3, 5'd24, 27'h00000186, 5'd12, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000243, 5'd25, 27'h00000174, 5'd20, 27'h00000323, 32'h00000400,
  1'd1,  5'd25, 27'h000002cb, 5'd0, 27'h000003c4, 5'd4, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000036e, 5'd4, 27'h000000df, 5'd13, 27'h00000256, 32'h00000400,
  1'd1,  5'd21, 27'h000002dc, 5'd3, 27'h000000fa, 5'd22, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003e7, 5'd10, 27'h00000342, 5'd3, 27'h0000027e, 32'h00000400,
  1'd1,  5'd23, 27'h00000151, 5'd11, 27'h000000ec, 5'd11, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000025d, 5'd13, 27'h000000df, 5'd22, 27'h000003bd, 32'h00000400,
  1'd1,  5'd25, 27'h00000302, 5'd24, 27'h00000032, 5'd1, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000062, 5'd22, 27'h000002b9, 5'd12, 27'h000001bf, 32'h00000400,
  1'd1,  5'd21, 27'h0000027c, 5'd23, 27'h000002d5, 5'd25, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000fc, 5'd3, 27'h000001a2, 5'd9, 27'h00000323, 32'h00000400,
  1'd1,  5'd3, 27'h00000210, 5'd5, 27'h00000023, 5'd18, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000325, 5'd2, 27'h000003f3, 5'd27, 27'h0000031d, 32'h00000400,
  1'd1,  5'd3, 27'h000002cc, 5'd12, 27'h0000024f, 5'd9, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000012f, 5'd12, 27'h000000f4, 5'd15, 27'h00000284, 32'h00000400,
  1'd1,  5'd4, 27'h00000092, 5'd13, 27'h000001f0, 5'd26, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000323, 5'd25, 27'h000001d9, 5'd8, 27'h00000256, 32'h00000400,
  1'd1,  5'd1, 27'h000001f0, 5'd21, 27'h000001fd, 5'd16, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000047, 5'd21, 27'h000003fe, 5'd26, 27'h00000050, 32'h00000400,
  1'd1,  5'd14, 27'h000000b7, 5'd3, 27'h000000ee, 5'd8, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f5, 5'd2, 27'h0000034c, 5'd18, 27'h0000003e, 32'h00000400,
  1'd1,  5'd10, 27'h0000015c, 5'd1, 27'h0000007f, 5'd26, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000007d, 5'd11, 27'h00000183, 5'd6, 27'h00000341, 32'h00000400,
  1'd1,  5'd13, 27'h0000031e, 5'd13, 27'h00000241, 5'd17, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000134, 5'd12, 27'h0000007c, 5'd28, 27'h00000315, 32'h00000400,
  1'd1,  5'd12, 27'h00000039, 5'd24, 27'h00000144, 5'd7, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000387, 5'd23, 27'h00000236, 5'd15, 27'h00000379, 32'h00000400,
  1'd1,  5'd10, 27'h000001c3, 5'd22, 27'h00000221, 5'd29, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000158, 5'd2, 27'h000000e2, 5'd9, 27'h000000ec, 32'h00000400,
  1'd1,  5'd22, 27'h00000372, 5'd3, 27'h000000b7, 5'd18, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000036d, 5'd3, 27'h00000335, 5'd26, 27'h00000071, 32'h00000400,
  1'd1,  5'd24, 27'h0000035c, 5'd11, 27'h000002b6, 5'd7, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000147, 5'd13, 27'h00000073, 5'd20, 27'h00000159, 32'h00000400,
  1'd1,  5'd23, 27'h00000374, 5'd13, 27'h00000228, 5'd27, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d5, 5'd25, 27'h000002d0, 5'd7, 27'h000000df, 32'h00000400,
  1'd1,  5'd21, 27'h000001af, 5'd24, 27'h000002d4, 5'd19, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e4, 5'd22, 27'h00000364, 5'd28, 27'h000001d7, 32'h00000400,
  1'd1,  5'd1, 27'h00000267, 5'd5, 27'h000000c0, 5'd2, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000015, 5'd5, 27'h000000ea, 5'd13, 27'h00000349, 32'h00000400,
  1'd1,  5'd1, 27'h0000020f, 5'd6, 27'h0000019d, 5'd21, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000297, 5'd16, 27'h00000306, 5'd0, 27'h0000021c, 32'h00000400,
  1'd1,  5'd0, 27'h000001e7, 5'd18, 27'h0000024c, 5'd13, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000059, 5'd19, 27'h00000294, 5'd21, 27'h00000070, 32'h00000400,
  1'd1,  5'd3, 27'h0000036f, 5'd28, 27'h00000056, 5'd4, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000008f, 5'd29, 27'h0000024c, 5'd14, 27'h000003a2, 32'h00000400,
  1'd1,  5'd4, 27'h000003e7, 5'd29, 27'h000003df, 5'd21, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031f, 5'd6, 27'h00000252, 5'd1, 27'h00000121, 32'h00000400,
  1'd1,  5'd10, 27'h000002cd, 5'd5, 27'h000001c6, 5'd10, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000245, 5'd10, 27'h00000122, 5'd23, 27'h000002a9, 32'h00000400,
  1'd1,  5'd15, 27'h00000043, 5'd16, 27'h00000203, 5'd1, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b6, 5'd18, 27'h00000368, 5'd11, 27'h000003de, 32'h00000400,
  1'd1,  5'd12, 27'h000002f5, 5'd16, 27'h000001be, 5'd24, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000010e, 5'd30, 27'h00000010, 5'd3, 27'h000003a2, 32'h00000400,
  1'd1,  5'd11, 27'h0000013f, 5'd26, 27'h00000252, 5'd13, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001b4, 5'd29, 27'h00000359, 5'd24, 27'h00000257, 32'h00000400,
  1'd1,  5'd21, 27'h000000fd, 5'd9, 27'h0000024b, 5'd3, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000179, 5'd10, 27'h000000be, 5'd10, 27'h000001aa, 32'h00000400,
  1'd1,  5'd22, 27'h0000007b, 5'd9, 27'h000002b5, 5'd25, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032a, 5'd15, 27'h000003a0, 5'd2, 27'h00000033, 32'h00000400,
  1'd1,  5'd21, 27'h00000374, 5'd15, 27'h00000201, 5'd14, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000052, 5'd16, 27'h00000084, 5'd22, 27'h0000032d, 32'h00000400,
  1'd1,  5'd24, 27'h000003d9, 5'd30, 27'h00000345, 5'd3, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003eb, 5'd28, 27'h00000197, 5'd12, 27'h000002c7, 32'h00000400,
  1'd1,  5'd24, 27'h000002aa, 5'd29, 27'h00000184, 5'd22, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000026b, 5'd8, 27'h0000034c, 5'd9, 27'h0000035b, 32'h00000400,
  1'd1,  5'd4, 27'h000003ef, 5'd7, 27'h000000bc, 5'd17, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000365, 5'd9, 27'h00000291, 5'd29, 27'h00000031, 32'h00000400,
  1'd1,  5'd3, 27'h000000a3, 5'd15, 27'h00000284, 5'd5, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000af, 5'd16, 27'h000001c9, 5'd18, 27'h00000023, 32'h00000400,
  1'd1,  5'd1, 27'h000003e1, 5'd17, 27'h00000378, 5'd28, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000033c, 5'd29, 27'h00000013, 5'd6, 27'h000003b9, 32'h00000400,
  1'd1,  5'd0, 27'h000000a5, 5'd26, 27'h000001b1, 5'd18, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032c, 5'd26, 27'h000000e6, 5'd28, 27'h00000290, 32'h00000400,
  1'd1,  5'd10, 27'h00000163, 5'd9, 27'h000002ef, 5'd6, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000123, 5'd6, 27'h00000025, 5'd17, 27'h000002fb, 32'h00000400,
  1'd1,  5'd11, 27'h0000008d, 5'd6, 27'h000002f9, 5'd30, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fa, 5'd19, 27'h000003ba, 5'd6, 27'h00000138, 32'h00000400,
  1'd1,  5'd12, 27'h00000075, 5'd16, 27'h000001ce, 5'd17, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003bb, 5'd16, 27'h0000038c, 5'd28, 27'h00000023, 32'h00000400,
  1'd1,  5'd11, 27'h00000343, 5'd30, 27'h00000261, 5'd6, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c3, 5'd30, 27'h0000038a, 5'd20, 27'h000001db, 32'h00000400,
  1'd1,  5'd14, 27'h00000136, 5'd28, 27'h000002ea, 5'd27, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ba, 5'd5, 27'h000000cb, 5'd8, 27'h0000003c, 32'h00000400,
  1'd1,  5'd25, 27'h0000016d, 5'd7, 27'h0000021e, 5'd18, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000231, 5'd7, 27'h00000073, 5'd28, 27'h0000014f, 32'h00000400,
  1'd1,  5'd22, 27'h00000330, 5'd17, 27'h000000bd, 5'd7, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fb, 5'd17, 27'h0000032e, 5'd18, 27'h00000376, 32'h00000400,
  1'd1,  5'd22, 27'h00000287, 5'd18, 27'h0000039c, 5'd30, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000136, 5'd27, 27'h0000025f, 5'd8, 27'h000002f3, 32'h00000400,
  1'd1,  5'd21, 27'h00000170, 5'd27, 27'h000003f9, 5'd18, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c9, 5'd25, 27'h000003dc, 5'd29, 27'h00000276, 32'h00000400,
  1'd1,  5'd5, 27'h00000252, 5'd4, 27'h00000296, 5'd5, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002ea, 5'd0, 27'h00000260, 5'd18, 27'h0000027c, 32'h00000400,
  1'd1,  5'd10, 27'h000000e2, 5'd1, 27'h0000007f, 5'd30, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e5, 5'd15, 27'h000001cc, 5'd3, 27'h0000028e, 32'h00000400,
  1'd1,  5'd6, 27'h00000312, 5'd12, 27'h00000368, 5'd11, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e2, 5'd13, 27'h0000024f, 5'd23, 27'h000003c5, 32'h00000400,
  1'd1,  5'd8, 27'h000002db, 5'd22, 27'h000003e1, 5'd3, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000f9, 5'd21, 27'h00000362, 5'd12, 27'h000000e1, 32'h00000400,
  1'd1,  5'd8, 27'h00000120, 5'd24, 27'h000000a8, 5'd22, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000036, 5'd3, 27'h000002c0, 5'd6, 27'h00000372, 32'h00000400,
  1'd1,  5'd17, 27'h00000153, 5'd4, 27'h000003ab, 5'd18, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ff, 5'd1, 27'h00000186, 5'd27, 27'h0000015f, 32'h00000400,
  1'd1,  5'd16, 27'h00000233, 5'd12, 27'h000000d0, 5'd0, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000398, 5'd12, 27'h00000059, 5'd14, 27'h00000352, 32'h00000400,
  1'd1,  5'd20, 27'h00000007, 5'd15, 27'h000001a1, 5'd21, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000093, 5'd22, 27'h00000296, 5'd4, 27'h00000180, 32'h00000400,
  1'd1,  5'd19, 27'h000002d3, 5'd23, 27'h000002fe, 5'd11, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002e8, 5'd24, 27'h0000005a, 5'd20, 27'h000002f6, 32'h00000400,
  1'd1,  5'd28, 27'h000003e7, 5'd0, 27'h0000010e, 5'd0, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ed, 5'd0, 27'h000003de, 5'd14, 27'h0000015a, 32'h00000400,
  1'd1,  5'd28, 27'h00000268, 5'd2, 27'h00000096, 5'd22, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b3, 5'd14, 27'h00000304, 5'd4, 27'h00000000, 32'h00000400,
  1'd1,  5'd30, 27'h0000019a, 5'd15, 27'h000001bd, 5'd12, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000231, 5'd12, 27'h00000370, 5'd22, 27'h00000372, 32'h00000400,
  1'd1,  5'd25, 27'h000003d1, 5'd23, 27'h000003ba, 5'd1, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f2, 5'd21, 27'h00000067, 5'd13, 27'h000003c7, 32'h00000400,
  1'd1,  5'd28, 27'h000002d0, 5'd20, 27'h0000034e, 5'd23, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000f7, 5'd3, 27'h00000281, 5'd1, 27'h000003a0, 32'h00000400,
  1'd1,  5'd7, 27'h000003a2, 5'd0, 27'h00000060, 5'd10, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000010b, 5'd1, 27'h0000015e, 5'd22, 27'h0000014d, 32'h00000400,
  1'd1,  5'd8, 27'h000000e3, 5'd11, 27'h00000173, 5'd5, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000cc, 5'd12, 27'h000002e6, 5'd18, 27'h000000e3, 32'h00000400,
  1'd1,  5'd5, 27'h000002f5, 5'd11, 27'h000000fd, 5'd27, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d0, 5'd21, 27'h0000035a, 5'd5, 27'h0000021d, 32'h00000400,
  1'd1,  5'd6, 27'h000000ba, 5'd24, 27'h000000a4, 5'd20, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000365, 5'd24, 27'h0000027e, 5'd29, 27'h000001ec, 32'h00000400,
  1'd1,  5'd19, 27'h00000039, 5'd2, 27'h000001be, 5'd1, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000094, 5'd1, 27'h000001b2, 5'd14, 27'h000001f6, 32'h00000400,
  1'd1,  5'd16, 27'h00000275, 5'd3, 27'h00000158, 5'd21, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001c4, 5'd10, 27'h00000374, 5'd9, 27'h000002bf, 32'h00000400,
  1'd1,  5'd20, 27'h00000223, 5'd11, 27'h000000ff, 5'd17, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000217, 5'd12, 27'h00000354, 5'd29, 27'h000003ba, 32'h00000400,
  1'd1,  5'd19, 27'h000002f8, 5'd23, 27'h00000329, 5'd9, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000096, 5'd25, 27'h000002cc, 5'd18, 27'h00000059, 32'h00000400,
  1'd1,  5'd17, 27'h00000322, 5'd22, 27'h00000369, 5'd27, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000035a, 5'd2, 27'h00000246, 5'd7, 27'h00000062, 32'h00000400,
  1'd1,  5'd28, 27'h000003a7, 5'd0, 27'h00000298, 5'd17, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000024c, 5'd2, 27'h00000186, 5'd30, 27'h00000087, 32'h00000400,
  1'd1,  5'd28, 27'h0000021c, 5'd13, 27'h0000035e, 5'd9, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000304, 5'd11, 27'h00000277, 5'd18, 27'h000000e7, 32'h00000400,
  1'd1,  5'd27, 27'h0000007d, 5'd10, 27'h0000027f, 5'd30, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000172, 5'd20, 27'h0000030b, 5'd5, 27'h000001d6, 32'h00000400,
  1'd1,  5'd26, 27'h000002a1, 5'd23, 27'h00000380, 5'd15, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000009a, 5'd25, 27'h00000206, 5'd28, 27'h0000002b, 32'h00000400,
  1'd1,  5'd5, 27'h00000147, 5'd5, 27'h00000392, 5'd3, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000189, 5'd9, 27'h00000282, 5'd10, 27'h000001d6, 32'h00000400,
  1'd1,  5'd6, 27'h0000009e, 5'd5, 27'h0000037c, 5'd22, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a5, 5'd18, 27'h00000064, 5'd1, 27'h000000b3, 32'h00000400,
  1'd1,  5'd8, 27'h0000009f, 5'd16, 27'h000001de, 5'd14, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003bc, 5'd20, 27'h000000b3, 5'd22, 27'h0000035a, 32'h00000400,
  1'd1,  5'd8, 27'h00000273, 5'd26, 27'h000003ac, 5'd4, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000366, 5'd30, 27'h000003c7, 5'd14, 27'h000003c5, 32'h00000400,
  1'd1,  5'd7, 27'h00000353, 5'd28, 27'h0000008d, 5'd23, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003a0, 5'd6, 27'h0000022b, 5'd5, 27'h00000039, 32'h00000400,
  1'd1,  5'd18, 27'h0000013c, 5'd6, 27'h000000b8, 5'd13, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ff, 5'd9, 27'h000002e5, 5'd25, 27'h00000251, 32'h00000400,
  1'd1,  5'd18, 27'h0000004a, 5'd19, 27'h000002c8, 5'd1, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000001b, 5'd19, 27'h00000318, 5'd13, 27'h000001c7, 32'h00000400,
  1'd1,  5'd20, 27'h0000022d, 5'd15, 27'h0000032b, 5'd25, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001dd, 5'd29, 27'h0000028b, 5'd2, 27'h0000001d, 32'h00000400,
  1'd1,  5'd16, 27'h00000262, 5'd28, 27'h000002d3, 5'd14, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000005d, 5'd30, 27'h00000141, 5'd24, 27'h0000007b, 32'h00000400,
  1'd1,  5'd29, 27'h000000c7, 5'd6, 27'h000002f4, 5'd2, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000c7, 5'd7, 27'h00000009, 5'd15, 27'h0000006f, 32'h00000400,
  1'd1,  5'd28, 27'h0000017e, 5'd7, 27'h00000346, 5'd24, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000015b, 5'd15, 27'h00000291, 5'd3, 27'h00000373, 32'h00000400,
  1'd1,  5'd28, 27'h00000209, 5'd20, 27'h000001a7, 5'd14, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001ac, 5'd19, 27'h000001c3, 5'd23, 27'h000003e9, 32'h00000400,
  1'd1,  5'd30, 27'h0000038e, 5'd29, 27'h000000a5, 5'd3, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000027d, 5'd30, 27'h0000036f, 5'd14, 27'h00000356, 32'h00000400,
  1'd1,  5'd29, 27'h00000239, 5'd28, 27'h000003a2, 5'd25, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000110, 5'd7, 27'h0000017a, 5'd6, 27'h0000005a, 32'h00000400,
  1'd1,  5'd9, 27'h0000003c, 5'd9, 27'h00000398, 5'd16, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000b3, 5'd6, 27'h0000031c, 5'd26, 27'h000003a0, 32'h00000400,
  1'd1,  5'd6, 27'h0000023c, 5'd19, 27'h000000ca, 5'd5, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000052, 5'd18, 27'h00000118, 5'd20, 27'h0000010d, 32'h00000400,
  1'd1,  5'd5, 27'h00000382, 5'd18, 27'h00000129, 5'd27, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000231, 5'd28, 27'h000003fc, 5'd8, 27'h000001e1, 32'h00000400,
  1'd1,  5'd8, 27'h00000245, 5'd25, 27'h000003a6, 5'd19, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c6, 5'd29, 27'h00000028, 5'd29, 27'h000001af, 32'h00000400,
  1'd1,  5'd17, 27'h000001f5, 5'd9, 27'h000000bc, 5'd6, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000036d, 5'd6, 27'h00000302, 5'd17, 27'h0000023f, 32'h00000400,
  1'd1,  5'd17, 27'h00000329, 5'd7, 27'h000001e2, 5'd29, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000002e, 5'd18, 27'h0000009f, 5'd7, 27'h00000354, 32'h00000400,
  1'd1,  5'd17, 27'h00000088, 5'd20, 27'h00000073, 5'd18, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000027a, 5'd18, 27'h000000a4, 5'd27, 27'h0000002d, 32'h00000400,
  1'd1,  5'd16, 27'h00000212, 5'd29, 27'h000001ee, 5'd5, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000017a, 5'd28, 27'h00000246, 5'd17, 27'h0000008c, 32'h00000400,
  1'd1,  5'd17, 27'h0000019c, 5'd30, 27'h000001dc, 5'd30, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000008a, 5'd7, 27'h000002ba, 5'd9, 27'h00000298, 32'h00000400,
  1'd1,  5'd30, 27'h000002e2, 5'd8, 27'h0000006f, 5'd19, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000018b, 5'd7, 27'h000003be, 5'd27, 27'h000002c5, 32'h00000400,
  1'd1,  5'd30, 27'h0000007a, 5'd15, 27'h00000280, 5'd6, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036d, 5'd15, 27'h000003fe, 5'd17, 27'h00000241, 32'h00000400,
  1'd1,  5'd30, 27'h000002aa, 5'd17, 27'h00000129, 5'd30, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000167, 5'd28, 27'h00000019, 5'd9, 27'h00000348, 32'h00000400,
  1'd1,  5'd29, 27'h000001d0, 5'd28, 27'h00000316, 5'd17, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012d, 5'd29, 27'h00000198, 5'd29, 27'h00000006, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000002de, 5'd1, 27'h000000c0, 5'd2, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000004d, 5'd5, 27'h00000038, 5'd11, 27'h00000215, 32'h00000400,
  1'd1,  5'd4, 27'h000000be, 5'd1, 27'h00000248, 5'd24, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000222, 5'd14, 27'h0000032f, 5'd3, 27'h000000ba, 32'h00000400,
  1'd1,  5'd0, 27'h00000131, 5'd14, 27'h000003be, 5'd11, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000110, 5'd13, 27'h0000016a, 5'd25, 27'h000001b2, 32'h00000400,
  1'd1,  5'd2, 27'h00000212, 5'd24, 27'h000001cf, 5'd1, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000384, 5'd23, 27'h000001ec, 5'd13, 27'h00000105, 32'h00000400,
  1'd1,  5'd0, 27'h000000fd, 5'd24, 27'h000003bf, 5'd24, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000025d, 5'd0, 27'h00000256, 5'd0, 27'h00000006, 32'h00000400,
  1'd1,  5'd13, 27'h0000024a, 5'd2, 27'h00000302, 5'd15, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003af, 5'd2, 27'h00000237, 5'd23, 27'h00000160, 32'h00000400,
  1'd1,  5'd13, 27'h000002c7, 5'd14, 27'h00000330, 5'd0, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000178, 5'd12, 27'h000002c4, 5'd14, 27'h00000010, 32'h00000400,
  1'd1,  5'd14, 27'h00000170, 5'd11, 27'h000001b1, 5'd25, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000047, 5'd21, 27'h000002c6, 5'd3, 27'h00000084, 32'h00000400,
  1'd1,  5'd14, 27'h0000003e, 5'd23, 27'h000002ae, 5'd14, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000373, 5'd25, 27'h00000231, 5'd24, 27'h000001dc, 32'h00000400,
  1'd1,  5'd23, 27'h00000218, 5'd3, 27'h000003ba, 5'd2, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000132, 5'd1, 27'h0000010c, 5'd13, 27'h00000197, 32'h00000400,
  1'd1,  5'd20, 27'h000003f2, 5'd3, 27'h00000003, 5'd21, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002dd, 5'd14, 27'h00000110, 5'd3, 27'h0000007e, 32'h00000400,
  1'd1,  5'd23, 27'h00000208, 5'd11, 27'h00000221, 5'd11, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002cd, 5'd14, 27'h000002e5, 5'd23, 27'h00000203, 32'h00000400,
  1'd1,  5'd23, 27'h0000032e, 5'd22, 27'h00000015, 5'd4, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000300, 5'd24, 27'h00000388, 5'd12, 27'h0000031b, 32'h00000400,
  1'd1,  5'd25, 27'h00000159, 5'd22, 27'h00000259, 5'd22, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000062, 5'd4, 27'h000002ae, 5'd7, 27'h000003d7, 32'h00000400,
  1'd1,  5'd3, 27'h000001da, 5'd4, 27'h00000153, 5'd15, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002dc, 5'd2, 27'h00000127, 5'd29, 27'h00000177, 32'h00000400,
  1'd1,  5'd0, 27'h00000139, 5'd13, 27'h000001d8, 5'd9, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000db, 5'd14, 27'h0000021d, 5'd18, 27'h000002e2, 32'h00000400,
  1'd1,  5'd4, 27'h00000044, 5'd11, 27'h000002e8, 5'd30, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d3, 5'd24, 27'h0000012c, 5'd5, 27'h000001ab, 32'h00000400,
  1'd1,  5'd0, 27'h0000021a, 5'd20, 27'h00000367, 5'd19, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000009c, 5'd24, 27'h000003ba, 5'd28, 27'h00000193, 32'h00000400,
  1'd1,  5'd14, 27'h000002b7, 5'd2, 27'h00000079, 5'd9, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f5, 5'd3, 27'h000001ff, 5'd18, 27'h00000127, 32'h00000400,
  1'd1,  5'd10, 27'h00000374, 5'd5, 27'h00000081, 5'd29, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c6, 5'd13, 27'h00000260, 5'd9, 27'h0000008e, 32'h00000400,
  1'd1,  5'd11, 27'h00000110, 5'd15, 27'h000000c9, 5'd17, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000399, 5'd11, 27'h0000004a, 5'd26, 27'h00000327, 32'h00000400,
  1'd1,  5'd11, 27'h0000001e, 5'd25, 27'h0000006c, 5'd7, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000256, 5'd20, 27'h0000038b, 5'd19, 27'h000002e0, 32'h00000400,
  1'd1,  5'd14, 27'h000000a3, 5'd24, 27'h000003f6, 5'd29, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c4, 5'd2, 27'h000003b0, 5'd7, 27'h00000115, 32'h00000400,
  1'd1,  5'd25, 27'h000002ba, 5'd2, 27'h000001da, 5'd16, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019d, 5'd1, 27'h0000016a, 5'd28, 27'h0000023e, 32'h00000400,
  1'd1,  5'd24, 27'h0000019a, 5'd11, 27'h000000d9, 5'd9, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000213, 5'd12, 27'h0000005c, 5'd19, 27'h0000022b, 32'h00000400,
  1'd1,  5'd23, 27'h000002a5, 5'd13, 27'h000002df, 5'd29, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003da, 5'd21, 27'h0000016e, 5'd5, 27'h000002f2, 32'h00000400,
  1'd1,  5'd25, 27'h00000173, 5'd24, 27'h00000098, 5'd16, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000158, 5'd24, 27'h0000024f, 5'd27, 27'h00000163, 32'h00000400,
  1'd1,  5'd0, 27'h00000253, 5'd9, 27'h000002b6, 5'd2, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022d, 5'd6, 27'h00000233, 5'd14, 27'h00000297, 32'h00000400,
  1'd1,  5'd1, 27'h0000020f, 5'd6, 27'h000003b3, 5'd24, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000000d, 5'd20, 27'h000001c3, 5'd4, 27'h000000ff, 32'h00000400,
  1'd1,  5'd4, 27'h00000334, 5'd16, 27'h000002e6, 5'd15, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003ab, 5'd19, 27'h00000333, 5'd21, 27'h0000008e, 32'h00000400,
  1'd1,  5'd1, 27'h00000350, 5'd29, 27'h000001e9, 5'd1, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a8, 5'd28, 27'h00000156, 5'd14, 27'h000000aa, 32'h00000400,
  1'd1,  5'd2, 27'h00000242, 5'd26, 27'h000001d6, 5'd24, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002c9, 5'd8, 27'h00000367, 5'd4, 27'h00000311, 32'h00000400,
  1'd1,  5'd10, 27'h000003e9, 5'd9, 27'h0000039f, 5'd13, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c1, 5'd7, 27'h00000390, 5'd22, 27'h000003fa, 32'h00000400,
  1'd1,  5'd12, 27'h000003e1, 5'd17, 27'h000001b7, 5'd0, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000218, 5'd18, 27'h000001ca, 5'd12, 27'h000003f1, 32'h00000400,
  1'd1,  5'd10, 27'h00000238, 5'd16, 27'h000001a5, 5'd23, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000325, 5'd30, 27'h000001cd, 5'd2, 27'h00000368, 32'h00000400,
  1'd1,  5'd15, 27'h000001b9, 5'd30, 27'h00000113, 5'd11, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000169, 5'd26, 27'h000000ef, 5'd22, 27'h00000104, 32'h00000400,
  1'd1,  5'd21, 27'h00000211, 5'd9, 27'h00000314, 5'd4, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000f3, 5'd5, 27'h00000184, 5'd12, 27'h0000022f, 32'h00000400,
  1'd1,  5'd22, 27'h000003d6, 5'd6, 27'h000003b3, 5'd22, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000398, 5'd17, 27'h0000007a, 5'd4, 27'h000003ee, 32'h00000400,
  1'd1,  5'd24, 27'h000002ca, 5'd19, 27'h000003f6, 5'd13, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002b8, 5'd15, 27'h0000029b, 5'd24, 27'h00000286, 32'h00000400,
  1'd1,  5'd21, 27'h000003ab, 5'd29, 27'h0000014f, 5'd1, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000033c, 5'd27, 27'h0000003d, 5'd12, 27'h000003e1, 32'h00000400,
  1'd1,  5'd22, 27'h00000172, 5'd30, 27'h00000241, 5'd23, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027a, 5'd7, 27'h000000d8, 5'd9, 27'h000000a2, 32'h00000400,
  1'd1,  5'd0, 27'h0000034c, 5'd9, 27'h000001b6, 5'd17, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000009b, 5'd7, 27'h000001b7, 5'd29, 27'h0000013a, 32'h00000400,
  1'd1,  5'd3, 27'h000002f5, 5'd18, 27'h0000031d, 5'd6, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000023e, 5'd20, 27'h000001f7, 5'd18, 27'h00000219, 32'h00000400,
  1'd1,  5'd3, 27'h0000017f, 5'd16, 27'h00000266, 5'd29, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000206, 5'd29, 27'h00000257, 5'd6, 27'h000003d9, 32'h00000400,
  1'd1,  5'd3, 27'h000003af, 5'd26, 27'h000002da, 5'd17, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000020d, 5'd29, 27'h00000194, 5'd27, 27'h00000209, 32'h00000400,
  1'd1,  5'd11, 27'h000001e5, 5'd6, 27'h000003f1, 5'd9, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000275, 5'd9, 27'h0000017c, 5'd18, 27'h000002f6, 32'h00000400,
  1'd1,  5'd14, 27'h0000008e, 5'd7, 27'h0000032e, 5'd30, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001bb, 5'd17, 27'h000002f9, 5'd6, 27'h00000088, 32'h00000400,
  1'd1,  5'd10, 27'h00000249, 5'd18, 27'h00000307, 5'd17, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000400, 5'd16, 27'h00000386, 5'd26, 27'h00000046, 32'h00000400,
  1'd1,  5'd10, 27'h000002f7, 5'd26, 27'h0000005b, 5'd7, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e7, 5'd29, 27'h000000ac, 5'd19, 27'h00000037, 32'h00000400,
  1'd1,  5'd14, 27'h000000ea, 5'd28, 27'h000003e2, 5'd28, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b5, 5'd7, 27'h00000271, 5'd6, 27'h000000dc, 32'h00000400,
  1'd1,  5'd25, 27'h0000018c, 5'd6, 27'h000000e4, 5'd15, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002ce, 5'd8, 27'h00000224, 5'd30, 27'h00000187, 32'h00000400,
  1'd1,  5'd21, 27'h000003a3, 5'd16, 27'h000001b8, 5'd6, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b2, 5'd15, 27'h000002ea, 5'd20, 27'h00000143, 32'h00000400,
  1'd1,  5'd24, 27'h000000bc, 5'd19, 27'h000003b2, 5'd27, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000399, 5'd27, 27'h00000136, 5'd8, 27'h00000121, 32'h00000400,
  1'd1,  5'd23, 27'h000003cb, 5'd27, 27'h00000381, 5'd19, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002a2, 5'd26, 27'h0000029b, 5'd26, 27'h00000281, 32'h00000400,
  1'd1,  5'd6, 27'h0000001e, 5'd4, 27'h0000019c, 5'd8, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e8, 5'd3, 27'h00000223, 5'd16, 27'h000000f7, 32'h00000400,
  1'd1,  5'd7, 27'h00000205, 5'd0, 27'h000000cc, 5'd30, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e0, 5'd12, 27'h000003dd, 5'd4, 27'h00000150, 32'h00000400,
  1'd1,  5'd9, 27'h000002fe, 5'd12, 27'h000001a1, 5'd11, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a0, 5'd13, 27'h000002b8, 5'd24, 27'h000000a3, 32'h00000400,
  1'd1,  5'd8, 27'h00000223, 5'd24, 27'h000002fd, 5'd0, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d1, 5'd24, 27'h00000045, 5'd14, 27'h00000088, 32'h00000400,
  1'd1,  5'd9, 27'h000002f5, 5'd20, 27'h00000330, 5'd24, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000198, 5'd1, 27'h000000fd, 5'd7, 27'h000000ed, 32'h00000400,
  1'd1,  5'd17, 27'h00000236, 5'd5, 27'h00000094, 5'd19, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029f, 5'd0, 27'h000000de, 5'd28, 27'h00000237, 32'h00000400,
  1'd1,  5'd20, 27'h00000165, 5'd12, 27'h000003a8, 5'd4, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003ea, 5'd15, 27'h000001f7, 5'd15, 27'h00000104, 32'h00000400,
  1'd1,  5'd16, 27'h000002b3, 5'd15, 27'h000001dc, 5'd25, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000017, 5'd22, 27'h00000144, 5'd2, 27'h00000202, 32'h00000400,
  1'd1,  5'd17, 27'h00000019, 5'd23, 27'h00000353, 5'd13, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000b5, 5'd21, 27'h000003d8, 5'd24, 27'h00000243, 32'h00000400,
  1'd1,  5'd28, 27'h000000f3, 5'd4, 27'h00000325, 5'd5, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ac, 5'd4, 27'h000002d1, 5'd11, 27'h0000019c, 32'h00000400,
  1'd1,  5'd30, 27'h00000183, 5'd0, 27'h00000005, 5'd23, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f3, 5'd11, 27'h000000d4, 5'd4, 27'h000001b5, 32'h00000400,
  1'd1,  5'd29, 27'h0000032f, 5'd14, 27'h000002b5, 5'd10, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000155, 5'd12, 27'h00000105, 5'd23, 27'h00000089, 32'h00000400,
  1'd1,  5'd27, 27'h000002e3, 5'd23, 27'h00000018, 5'd2, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ee, 5'd25, 27'h000000c2, 5'd13, 27'h000000f6, 32'h00000400,
  1'd1,  5'd30, 27'h0000004e, 5'd23, 27'h000003bf, 5'd21, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000292, 5'd3, 27'h00000211, 5'd1, 27'h00000217, 32'h00000400,
  1'd1,  5'd10, 27'h00000033, 5'd3, 27'h0000003b, 5'd14, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002fe, 5'd0, 27'h000000ce, 5'd23, 27'h00000014, 32'h00000400,
  1'd1,  5'd8, 27'h000002ce, 5'd13, 27'h000003ed, 5'd8, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e5, 5'd12, 27'h00000134, 5'd19, 27'h000000c1, 32'h00000400,
  1'd1,  5'd10, 27'h00000148, 5'd12, 27'h000002ff, 5'd28, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000268, 5'd20, 27'h0000032a, 5'd8, 27'h00000071, 32'h00000400,
  1'd1,  5'd7, 27'h0000027d, 5'd24, 27'h00000346, 5'd18, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000156, 5'd25, 27'h000001c3, 5'd30, 27'h00000272, 32'h00000400,
  1'd1,  5'd17, 27'h000001d8, 5'd3, 27'h00000377, 5'd4, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000034b, 5'd2, 27'h00000240, 5'd11, 27'h000003b3, 32'h00000400,
  1'd1,  5'd17, 27'h000002b0, 5'd2, 27'h00000151, 5'd22, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000278, 5'd12, 27'h0000001c, 5'd8, 27'h0000004b, 32'h00000400,
  1'd1,  5'd18, 27'h000002ff, 5'd12, 27'h00000386, 5'd20, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000027f, 5'd11, 27'h000000e5, 5'd27, 27'h00000058, 32'h00000400,
  1'd1,  5'd16, 27'h000001ff, 5'd24, 27'h000001e6, 5'd6, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000f0, 5'd25, 27'h000000e1, 5'd20, 27'h00000131, 32'h00000400,
  1'd1,  5'd15, 27'h00000294, 5'd22, 27'h0000019a, 5'd29, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000033e, 5'd1, 27'h0000011d, 5'd8, 27'h000003c0, 32'h00000400,
  1'd1,  5'd27, 27'h00000391, 5'd1, 27'h000000bc, 5'd16, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a3, 5'd3, 27'h00000069, 5'd30, 27'h000000e2, 32'h00000400,
  1'd1,  5'd27, 27'h000002a1, 5'd13, 27'h00000269, 5'd9, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002ea, 5'd13, 27'h00000061, 5'd19, 27'h0000024f, 32'h00000400,
  1'd1,  5'd29, 27'h000001a1, 5'd13, 27'h000003bd, 5'd30, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e7, 5'd25, 27'h00000267, 5'd7, 27'h000000c1, 32'h00000400,
  1'd1,  5'd29, 27'h0000011c, 5'd25, 27'h000001d8, 5'd16, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001dd, 5'd22, 27'h00000347, 5'd27, 27'h0000008b, 32'h00000400,
  1'd1,  5'd8, 27'h00000017, 5'd8, 27'h000002ae, 5'd4, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000279, 5'd10, 27'h0000002b, 5'd11, 27'h00000041, 32'h00000400,
  1'd1,  5'd7, 27'h000000ff, 5'd7, 27'h0000030e, 5'd22, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000018, 5'd18, 27'h000000b3, 5'd3, 27'h00000185, 32'h00000400,
  1'd1,  5'd8, 27'h000001e7, 5'd17, 27'h00000009, 5'd13, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038e, 5'd15, 27'h000003ba, 5'd24, 27'h000002ac, 32'h00000400,
  1'd1,  5'd5, 27'h000003ec, 5'd27, 27'h000000a4, 5'd3, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000095, 5'd30, 27'h000003ac, 5'd15, 27'h00000082, 32'h00000400,
  1'd1,  5'd8, 27'h00000248, 5'd26, 27'h00000180, 5'd22, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000de, 5'd6, 27'h00000172, 5'd4, 27'h00000017, 32'h00000400,
  1'd1,  5'd18, 27'h0000004d, 5'd5, 27'h000002cc, 5'd13, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d0, 5'd5, 27'h000003d6, 5'd24, 27'h000002e3, 32'h00000400,
  1'd1,  5'd16, 27'h000003e4, 5'd17, 27'h00000083, 5'd2, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000a8, 5'd16, 27'h0000018f, 5'd13, 27'h00000303, 32'h00000400,
  1'd1,  5'd16, 27'h000001aa, 5'd19, 27'h000001f2, 5'd21, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000276, 5'd27, 27'h00000004, 5'd2, 27'h00000180, 32'h00000400,
  1'd1,  5'd19, 27'h00000071, 5'd28, 27'h00000313, 5'd13, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ae, 5'd30, 27'h000003c0, 5'd24, 27'h000000b1, 32'h00000400,
  1'd1,  5'd26, 27'h00000266, 5'd8, 27'h00000361, 5'd2, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000101, 5'd5, 27'h0000010e, 5'd11, 27'h0000001a, 32'h00000400,
  1'd1,  5'd28, 27'h000003f8, 5'd9, 27'h000001a0, 5'd21, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000320, 5'd15, 27'h0000021c, 5'd1, 27'h00000372, 32'h00000400,
  1'd1,  5'd27, 27'h000000f1, 5'd16, 27'h0000025d, 5'd11, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000e1, 5'd17, 27'h00000004, 5'd23, 27'h00000056, 32'h00000400,
  1'd1,  5'd26, 27'h00000263, 5'd30, 27'h0000025e, 5'd2, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000048, 5'd26, 27'h00000353, 5'd10, 27'h0000018b, 32'h00000400,
  1'd1,  5'd29, 27'h00000311, 5'd26, 27'h00000040, 5'd20, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000018b, 5'd9, 27'h000003fc, 5'd5, 27'h0000023c, 32'h00000400,
  1'd1,  5'd7, 27'h00000398, 5'd6, 27'h00000340, 5'd16, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e5, 5'd6, 27'h000002b5, 5'd30, 27'h00000109, 32'h00000400,
  1'd1,  5'd8, 27'h000000c2, 5'd18, 27'h000000a8, 5'd6, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e3, 5'd17, 27'h00000035, 5'd16, 27'h00000317, 32'h00000400,
  1'd1,  5'd7, 27'h000001fe, 5'd17, 27'h00000281, 5'd26, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002a9, 5'd28, 27'h00000381, 5'd7, 27'h00000125, 32'h00000400,
  1'd1,  5'd8, 27'h0000011b, 5'd27, 27'h000001d5, 5'd17, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000198, 5'd28, 27'h0000000f, 5'd28, 27'h00000138, 32'h00000400,
  1'd1,  5'd15, 27'h000002c8, 5'd8, 27'h00000073, 5'd8, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001f2, 5'd9, 27'h000001ff, 5'd18, 27'h0000005c, 32'h00000400,
  1'd1,  5'd16, 27'h00000152, 5'd9, 27'h0000001c, 5'd27, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002e1, 5'd16, 27'h00000304, 5'd10, 27'h000000d1, 32'h00000400,
  1'd1,  5'd19, 27'h0000028d, 5'd17, 27'h000002b3, 5'd16, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d6, 5'd16, 27'h00000072, 5'd28, 27'h00000322, 32'h00000400,
  1'd1,  5'd15, 27'h00000360, 5'd27, 27'h0000016d, 5'd10, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000149, 5'd28, 27'h000002f2, 5'd15, 27'h0000039c, 32'h00000400,
  1'd1,  5'd19, 27'h000003c8, 5'd30, 27'h000002fc, 5'd26, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000009d, 5'd8, 27'h00000332, 5'd8, 27'h000003a2, 32'h00000400,
  1'd1,  5'd29, 27'h0000036c, 5'd8, 27'h000003a8, 5'd17, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000078, 5'd7, 27'h00000375, 5'd27, 27'h0000039c, 32'h00000400,
  1'd1,  5'd30, 27'h00000272, 5'd17, 27'h000002e6, 5'd6, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001aa, 5'd16, 27'h000002ae, 5'd19, 27'h000001bc, 32'h00000400,
  1'd1,  5'd29, 27'h000002a5, 5'd16, 27'h0000025a, 5'd29, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ec, 5'd29, 27'h0000002c, 5'd6, 27'h0000014d, 32'h00000400,
  1'd1,  5'd26, 27'h000002a3, 5'd29, 27'h0000025e, 5'd18, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b3, 5'd26, 27'h000001db, 5'd30, 27'h00000007, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000084, 5'd3, 27'h00000258, 5'd0, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000390, 5'd2, 27'h000003c8, 5'd10, 27'h0000015e, 32'h00000400,
  1'd1,  5'd2, 27'h00000158, 5'd0, 27'h00000324, 5'd21, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000399, 5'd10, 27'h00000232, 5'd4, 27'h00000349, 32'h00000400,
  1'd1,  5'd1, 27'h0000023c, 5'd14, 27'h0000013b, 5'd14, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000012, 5'd14, 27'h000001bd, 5'd23, 27'h00000133, 32'h00000400,
  1'd1,  5'd0, 27'h000000cf, 5'd24, 27'h000002bf, 5'd1, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000017e, 5'd23, 27'h00000018, 5'd11, 27'h0000011d, 32'h00000400,
  1'd1,  5'd1, 27'h000001b2, 5'd25, 27'h0000000e, 5'd25, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000324, 5'd3, 27'h000002aa, 5'd3, 27'h00000355, 32'h00000400,
  1'd1,  5'd14, 27'h00000077, 5'd2, 27'h00000169, 5'd10, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f0, 5'd1, 27'h00000226, 5'd22, 27'h0000010a, 32'h00000400,
  1'd1,  5'd14, 27'h000001da, 5'd14, 27'h000003e6, 5'd4, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000018d, 5'd11, 27'h0000013f, 5'd14, 27'h000003d2, 32'h00000400,
  1'd1,  5'd13, 27'h00000199, 5'd11, 27'h00000154, 5'd21, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002c8, 5'd23, 27'h00000165, 5'd2, 27'h0000035f, 32'h00000400,
  1'd1,  5'd15, 27'h0000000e, 5'd23, 27'h000000ef, 5'd12, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d1, 5'd20, 27'h000003b2, 5'd24, 27'h000000ae, 32'h00000400,
  1'd1,  5'd22, 27'h0000016c, 5'd2, 27'h000002f9, 5'd4, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000020b, 5'd3, 27'h000001d0, 5'd13, 27'h000003da, 32'h00000400,
  1'd1,  5'd21, 27'h000000af, 5'd1, 27'h00000324, 5'd23, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000294, 5'd11, 27'h000000b2, 5'd0, 27'h000001eb, 32'h00000400,
  1'd1,  5'd23, 27'h000002c3, 5'd11, 27'h00000189, 5'd14, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001fb, 5'd11, 27'h000000db, 5'd20, 27'h000003fd, 32'h00000400,
  1'd1,  5'd24, 27'h00000152, 5'd25, 27'h000000de, 5'd5, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b3, 5'd23, 27'h0000038d, 5'd13, 27'h00000052, 32'h00000400,
  1'd1,  5'd24, 27'h00000078, 5'd21, 27'h0000021a, 5'd24, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000136, 5'd0, 27'h0000034f, 5'd7, 27'h000002cb, 32'h00000400,
  1'd1,  5'd1, 27'h00000385, 5'd5, 27'h00000087, 5'd16, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000132, 5'd4, 27'h00000161, 5'd30, 27'h000000fd, 32'h00000400,
  1'd1,  5'd1, 27'h000001dc, 5'd13, 27'h00000319, 5'd8, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000057, 5'd10, 27'h00000390, 5'd17, 27'h000002d5, 32'h00000400,
  1'd1,  5'd0, 27'h000002cd, 5'd11, 27'h000000eb, 5'd28, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000350, 5'd23, 27'h000003e3, 5'd9, 27'h00000098, 32'h00000400,
  1'd1,  5'd4, 27'h00000317, 5'd23, 27'h00000251, 5'd18, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d3, 5'd25, 27'h00000213, 5'd26, 27'h0000036d, 32'h00000400,
  1'd1,  5'd12, 27'h0000010e, 5'd0, 27'h00000106, 5'd8, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000004c, 5'd4, 27'h000000cd, 5'd18, 27'h00000184, 32'h00000400,
  1'd1,  5'd15, 27'h0000014f, 5'd2, 27'h0000015a, 5'd30, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002b2, 5'd11, 27'h000003d0, 5'd6, 27'h000000ec, 32'h00000400,
  1'd1,  5'd14, 27'h000003af, 5'd13, 27'h0000038c, 5'd19, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000386, 5'd10, 27'h0000018e, 5'd29, 27'h0000032d, 32'h00000400,
  1'd1,  5'd15, 27'h000000ef, 5'd24, 27'h000002a7, 5'd8, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a9, 5'd24, 27'h000002b4, 5'd16, 27'h0000034a, 32'h00000400,
  1'd1,  5'd13, 27'h000001a5, 5'd23, 27'h00000286, 5'd30, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000373, 5'd4, 27'h0000021d, 5'd6, 27'h00000325, 32'h00000400,
  1'd1,  5'd20, 27'h000002d4, 5'd3, 27'h00000057, 5'd19, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000315, 5'd3, 27'h000001ad, 5'd30, 27'h000001b8, 32'h00000400,
  1'd1,  5'd24, 27'h0000039c, 5'd11, 27'h000002a8, 5'd9, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a0, 5'd14, 27'h0000023e, 5'd19, 27'h00000072, 32'h00000400,
  1'd1,  5'd25, 27'h00000014, 5'd12, 27'h000003a5, 5'd28, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000269, 5'd22, 27'h00000152, 5'd7, 27'h00000067, 32'h00000400,
  1'd1,  5'd23, 27'h00000161, 5'd23, 27'h00000056, 5'd19, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038e, 5'd22, 27'h0000024f, 5'd29, 27'h000002de, 32'h00000400,
  1'd1,  5'd2, 27'h000000ba, 5'd5, 27'h000001fb, 5'd4, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000259, 5'd5, 27'h000001d6, 5'd13, 27'h00000052, 32'h00000400,
  1'd1,  5'd4, 27'h00000110, 5'd9, 27'h00000335, 5'd22, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000250, 5'd19, 27'h000000b5, 5'd2, 27'h00000241, 32'h00000400,
  1'd1,  5'd2, 27'h00000171, 5'd20, 27'h0000021d, 5'd14, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000171, 5'd19, 27'h00000224, 5'd22, 27'h00000371, 32'h00000400,
  1'd1,  5'd3, 27'h00000024, 5'd28, 27'h00000327, 5'd3, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000086, 5'd30, 27'h00000073, 5'd15, 27'h00000127, 32'h00000400,
  1'd1,  5'd1, 27'h00000246, 5'd28, 27'h000001fc, 5'd22, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000281, 5'd8, 27'h00000216, 5'd0, 27'h000003f6, 32'h00000400,
  1'd1,  5'd14, 27'h0000004b, 5'd9, 27'h000000f4, 5'd10, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003dc, 5'd5, 27'h000002c0, 5'd23, 27'h00000221, 32'h00000400,
  1'd1,  5'd15, 27'h000000cf, 5'd19, 27'h0000030c, 5'd4, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000341, 5'd18, 27'h0000035a, 5'd12, 27'h0000020f, 32'h00000400,
  1'd1,  5'd12, 27'h00000089, 5'd16, 27'h000001da, 5'd22, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a4, 5'd26, 27'h0000032a, 5'd3, 27'h000002c5, 32'h00000400,
  1'd1,  5'd10, 27'h000003a7, 5'd26, 27'h000002f4, 5'd11, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000019f, 5'd27, 27'h000000bd, 5'd24, 27'h00000047, 32'h00000400,
  1'd1,  5'd25, 27'h0000004b, 5'd8, 27'h000002a2, 5'd1, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000011b, 5'd7, 27'h00000398, 5'd12, 27'h00000286, 32'h00000400,
  1'd1,  5'd22, 27'h00000120, 5'd9, 27'h0000002c, 5'd22, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038a, 5'd16, 27'h000003d3, 5'd0, 27'h000002db, 32'h00000400,
  1'd1,  5'd21, 27'h00000199, 5'd16, 27'h000001ba, 5'd13, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000000c, 5'd20, 27'h000000fe, 5'd25, 27'h0000030c, 32'h00000400,
  1'd1,  5'd22, 27'h000002e1, 5'd28, 27'h000002f6, 5'd4, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000003b, 5'd30, 27'h0000006c, 5'd12, 27'h000002b1, 32'h00000400,
  1'd1,  5'd24, 27'h00000106, 5'd29, 27'h0000020f, 5'd22, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000c7, 5'd9, 27'h00000369, 5'd6, 27'h000002f2, 32'h00000400,
  1'd1,  5'd0, 27'h00000219, 5'd7, 27'h0000011d, 5'd19, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020f, 5'd7, 27'h0000002e, 5'd29, 27'h00000186, 32'h00000400,
  1'd1,  5'd0, 27'h00000357, 5'd15, 27'h000002cd, 5'd6, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000357, 5'd19, 27'h00000274, 5'd17, 27'h00000249, 32'h00000400,
  1'd1,  5'd4, 27'h00000086, 5'd17, 27'h00000170, 5'd29, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000015b, 5'd27, 27'h000001e4, 5'd7, 27'h00000132, 32'h00000400,
  1'd1,  5'd5, 27'h00000013, 5'd27, 27'h00000152, 5'd17, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000223, 5'd26, 27'h0000023b, 5'd28, 27'h0000002c, 32'h00000400,
  1'd1,  5'd13, 27'h000000cd, 5'd8, 27'h00000044, 5'd8, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000382, 5'd9, 27'h000003ba, 5'd17, 27'h00000212, 32'h00000400,
  1'd1,  5'd13, 27'h000002a9, 5'd7, 27'h00000086, 5'd29, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021b, 5'd16, 27'h00000331, 5'd6, 27'h00000031, 32'h00000400,
  1'd1,  5'd10, 27'h000002c7, 5'd16, 27'h0000008a, 5'd16, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002ce, 5'd20, 27'h00000215, 5'd30, 27'h000003a2, 32'h00000400,
  1'd1,  5'd14, 27'h00000127, 5'd26, 27'h00000121, 5'd6, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c6, 5'd30, 27'h00000060, 5'd18, 27'h000001d1, 32'h00000400,
  1'd1,  5'd12, 27'h000001c9, 5'd30, 27'h000000e9, 5'd30, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fa, 5'd8, 27'h00000275, 5'd9, 27'h000001ea, 32'h00000400,
  1'd1,  5'd22, 27'h0000013e, 5'd9, 27'h00000032, 5'd15, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000020f, 5'd5, 27'h0000039f, 5'd28, 27'h000001f0, 32'h00000400,
  1'd1,  5'd20, 27'h00000315, 5'd17, 27'h00000250, 5'd9, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000066, 5'd19, 27'h00000129, 5'd18, 27'h000002ec, 32'h00000400,
  1'd1,  5'd22, 27'h000000a2, 5'd18, 27'h00000123, 5'd26, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000c5, 5'd26, 27'h000000ed, 5'd10, 27'h0000005c, 32'h00000400,
  1'd1,  5'd23, 27'h000003b4, 5'd26, 27'h00000133, 5'd15, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000050, 5'd26, 27'h000000cf, 5'd26, 27'h00000279, 32'h00000400,
  1'd1,  5'd6, 27'h00000170, 5'd3, 27'h00000272, 5'd6, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000a6, 5'd1, 27'h00000149, 5'd16, 27'h0000018c, 32'h00000400,
  1'd1,  5'd8, 27'h000002b1, 5'd1, 27'h000001fa, 5'd30, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011a, 5'd13, 27'h00000191, 5'd0, 27'h0000036d, 32'h00000400,
  1'd1,  5'd8, 27'h00000330, 5'd15, 27'h000001d2, 5'd10, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a1, 5'd14, 27'h00000133, 5'd21, 27'h0000029d, 32'h00000400,
  1'd1,  5'd5, 27'h000000cf, 5'd21, 27'h00000107, 5'd2, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000192, 5'd23, 27'h00000119, 5'd14, 27'h00000387, 32'h00000400,
  1'd1,  5'd9, 27'h00000046, 5'd25, 27'h000002d5, 5'd20, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000302, 5'd4, 27'h00000088, 5'd7, 27'h0000037f, 32'h00000400,
  1'd1,  5'd17, 27'h00000341, 5'd0, 27'h00000290, 5'd18, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000269, 5'd4, 27'h0000016d, 5'd27, 27'h0000019e, 32'h00000400,
  1'd1,  5'd18, 27'h000000c1, 5'd11, 27'h00000223, 5'd3, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000363, 5'd13, 27'h00000046, 5'd10, 27'h000002d3, 32'h00000400,
  1'd1,  5'd16, 27'h0000038a, 5'd11, 27'h00000321, 5'd23, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000214, 5'd21, 27'h000001f7, 5'd4, 27'h000001e2, 32'h00000400,
  1'd1,  5'd17, 27'h00000295, 5'd22, 27'h00000286, 5'd14, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000003a, 5'd25, 27'h00000146, 5'd24, 27'h00000309, 32'h00000400,
  1'd1,  5'd30, 27'h00000205, 5'd4, 27'h000000ee, 5'd1, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a9, 5'd4, 27'h0000031a, 5'd14, 27'h0000030e, 32'h00000400,
  1'd1,  5'd30, 27'h000003a7, 5'd4, 27'h0000033b, 5'd25, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000016, 5'd11, 27'h00000087, 5'd5, 27'h00000071, 32'h00000400,
  1'd1,  5'd28, 27'h00000227, 5'd10, 27'h00000391, 5'd13, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003aa, 5'd12, 27'h0000001c, 5'd21, 27'h00000232, 32'h00000400,
  1'd1,  5'd26, 27'h0000019a, 5'd23, 27'h000000ed, 5'd4, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b8, 5'd22, 27'h000001b4, 5'd14, 27'h000000d9, 32'h00000400,
  1'd1,  5'd29, 27'h000002f3, 5'd21, 27'h000002b1, 5'd22, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031f, 5'd0, 27'h000003d0, 5'd0, 27'h000000cd, 32'h00000400,
  1'd1,  5'd5, 27'h00000281, 5'd3, 27'h00000388, 5'd12, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000025b, 5'd2, 27'h0000005b, 5'd24, 27'h00000040, 32'h00000400,
  1'd1,  5'd7, 27'h00000265, 5'd15, 27'h00000081, 5'd8, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000226, 5'd12, 27'h000000ac, 5'd17, 27'h0000020f, 32'h00000400,
  1'd1,  5'd8, 27'h00000091, 5'd12, 27'h000002d9, 5'd28, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003be, 5'd23, 27'h00000336, 5'd5, 27'h00000265, 32'h00000400,
  1'd1,  5'd8, 27'h00000222, 5'd25, 27'h00000317, 5'd16, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000338, 5'd22, 27'h0000013c, 5'd29, 27'h000000f4, 32'h00000400,
  1'd1,  5'd19, 27'h0000031f, 5'd5, 27'h00000003, 5'd4, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003ce, 5'd1, 27'h0000001d, 5'd13, 27'h0000015a, 32'h00000400,
  1'd1,  5'd15, 27'h000003a7, 5'd2, 27'h00000208, 5'd21, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000367, 5'd11, 27'h000002fa, 5'd6, 27'h000000c5, 32'h00000400,
  1'd1,  5'd20, 27'h00000017, 5'd13, 27'h00000169, 5'd17, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000285, 5'd12, 27'h00000092, 5'd28, 27'h000002c2, 32'h00000400,
  1'd1,  5'd17, 27'h000001a5, 5'd23, 27'h00000004, 5'd6, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002ca, 5'd24, 27'h0000013c, 5'd17, 27'h0000034e, 32'h00000400,
  1'd1,  5'd18, 27'h000002c9, 5'd24, 27'h000000bb, 5'd29, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003d8, 5'd4, 27'h000000a7, 5'd9, 27'h000001ea, 32'h00000400,
  1'd1,  5'd29, 27'h00000136, 5'd0, 27'h000001dd, 5'd15, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000330, 5'd0, 27'h000000c2, 5'd30, 27'h000000c9, 32'h00000400,
  1'd1,  5'd27, 27'h0000035d, 5'd10, 27'h000001df, 5'd10, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b0, 5'd11, 27'h000002f8, 5'd16, 27'h00000192, 32'h00000400,
  1'd1,  5'd30, 27'h000002fd, 5'd15, 27'h0000016d, 5'd30, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000098, 5'd20, 27'h00000321, 5'd8, 27'h0000035d, 32'h00000400,
  1'd1,  5'd28, 27'h000001ce, 5'd25, 27'h0000004e, 5'd19, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003fe, 5'd22, 27'h000001fd, 5'd26, 27'h000002bc, 32'h00000400,
  1'd1,  5'd7, 27'h00000371, 5'd9, 27'h0000035b, 5'd2, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000030f, 5'd5, 27'h0000020b, 5'd13, 27'h00000017, 32'h00000400,
  1'd1,  5'd7, 27'h0000024c, 5'd6, 27'h00000061, 5'd23, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000126, 5'd19, 27'h0000021a, 5'd3, 27'h000002de, 32'h00000400,
  1'd1,  5'd10, 27'h0000002a, 5'd19, 27'h000003ea, 5'd11, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b3, 5'd19, 27'h0000037f, 5'd25, 27'h000002a8, 32'h00000400,
  1'd1,  5'd6, 27'h000000cc, 5'd29, 27'h0000038a, 5'd2, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000100, 5'd30, 27'h000000e4, 5'd12, 27'h000002bc, 32'h00000400,
  1'd1,  5'd8, 27'h0000010a, 5'd30, 27'h00000159, 5'd25, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000033d, 5'd5, 27'h00000384, 5'd1, 27'h000000d2, 32'h00000400,
  1'd1,  5'd15, 27'h00000326, 5'd6, 27'h0000008a, 5'd11, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000171, 5'd8, 27'h000000b9, 5'd24, 27'h00000245, 32'h00000400,
  1'd1,  5'd20, 27'h000001ad, 5'd19, 27'h0000023f, 5'd1, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d0, 5'd17, 27'h000001c9, 5'd13, 27'h000002bb, 32'h00000400,
  1'd1,  5'd20, 27'h000000a1, 5'd19, 27'h00000194, 5'd23, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f6, 5'd26, 27'h00000381, 5'd1, 27'h000000e2, 32'h00000400,
  1'd1,  5'd19, 27'h000001cb, 5'd28, 27'h00000211, 5'd11, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000172, 5'd27, 27'h000000d5, 5'd22, 27'h00000388, 32'h00000400,
  1'd1,  5'd26, 27'h0000007b, 5'd6, 27'h000003a0, 5'd3, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000384, 5'd5, 27'h00000280, 5'd13, 27'h0000029a, 32'h00000400,
  1'd1,  5'd29, 27'h000003e5, 5'd6, 27'h00000329, 5'd22, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e6, 5'd19, 27'h000001eb, 5'd3, 27'h000000c5, 32'h00000400,
  1'd1,  5'd29, 27'h00000169, 5'd15, 27'h0000036f, 5'd14, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000033c, 5'd20, 27'h00000134, 5'd25, 27'h00000326, 32'h00000400,
  1'd1,  5'd29, 27'h000002d8, 5'd28, 27'h00000015, 5'd4, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ce, 5'd29, 27'h0000026f, 5'd13, 27'h0000017b, 32'h00000400,
  1'd1,  5'd26, 27'h0000010a, 5'd28, 27'h00000059, 5'd25, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000027, 5'd7, 27'h00000046, 5'd7, 27'h000001fe, 32'h00000400,
  1'd1,  5'd9, 27'h000000c2, 5'd8, 27'h0000032b, 5'd18, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000382, 5'd9, 27'h00000311, 5'd26, 27'h000001f7, 32'h00000400,
  1'd1,  5'd6, 27'h00000130, 5'd19, 27'h000001d8, 5'd8, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002bc, 5'd15, 27'h0000034b, 5'd19, 27'h00000092, 32'h00000400,
  1'd1,  5'd10, 27'h00000111, 5'd16, 27'h00000131, 5'd30, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b2, 5'd26, 27'h000001e5, 5'd9, 27'h00000017, 32'h00000400,
  1'd1,  5'd6, 27'h0000037d, 5'd27, 27'h00000025, 5'd16, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000d3, 5'd28, 27'h000001e5, 5'd28, 27'h00000310, 32'h00000400,
  1'd1,  5'd16, 27'h0000006e, 5'd9, 27'h000001eb, 5'd9, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002cd, 5'd9, 27'h0000027a, 5'd20, 27'h00000082, 32'h00000400,
  1'd1,  5'd18, 27'h000000ae, 5'd7, 27'h0000014f, 5'd26, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000094, 5'd18, 27'h000003bb, 5'd6, 27'h00000273, 32'h00000400,
  1'd1,  5'd17, 27'h000000c7, 5'd17, 27'h00000370, 5'd16, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f4, 5'd16, 27'h000002ea, 5'd27, 27'h00000082, 32'h00000400,
  1'd1,  5'd17, 27'h00000265, 5'd26, 27'h000003d6, 5'd5, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ef, 5'd25, 27'h000003ae, 5'd20, 27'h0000018f, 32'h00000400,
  1'd1,  5'd17, 27'h000003c9, 5'd27, 27'h0000032a, 5'd29, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003d8, 5'd7, 27'h00000095, 5'd8, 27'h0000003e, 32'h00000400,
  1'd1,  5'd30, 27'h0000036b, 5'd9, 27'h000002fe, 5'd16, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000010f, 5'd6, 27'h000000b2, 5'd26, 27'h00000280, 32'h00000400,
  1'd1,  5'd30, 27'h0000027c, 5'd17, 27'h000003b0, 5'd8, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000313, 5'd19, 27'h000002cf, 5'd20, 27'h0000004d, 32'h00000400,
  1'd1,  5'd26, 27'h00000062, 5'd17, 27'h000001fb, 5'd26, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000005d, 5'd29, 27'h00000081, 5'd9, 27'h00000154, 32'h00000400,
  1'd1,  5'd29, 27'h000001e7, 5'd29, 27'h00000217, 5'd16, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000009d, 5'd29, 27'h000002d8, 5'd29, 27'h0000039f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000002b8, 5'd1, 27'h00000117, 5'd4, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002d9, 5'd2, 27'h0000016f, 5'd12, 27'h000002ff, 32'h00000400,
  1'd1,  5'd3, 27'h000000b9, 5'd2, 27'h00000180, 5'd25, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000001e, 5'd14, 27'h00000135, 5'd2, 27'h00000274, 32'h00000400,
  1'd1,  5'd3, 27'h0000007f, 5'd11, 27'h00000013, 5'd10, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000009e, 5'd14, 27'h000003de, 5'd21, 27'h0000009e, 32'h00000400,
  1'd1,  5'd2, 27'h000000fe, 5'd24, 27'h000003e1, 5'd4, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002cc, 5'd23, 27'h0000015c, 5'd12, 27'h0000039e, 32'h00000400,
  1'd1,  5'd4, 27'h0000027a, 5'd21, 27'h000001b6, 5'd20, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003dd, 5'd4, 27'h00000150, 5'd5, 27'h000000a9, 32'h00000400,
  1'd1,  5'd14, 27'h00000028, 5'd0, 27'h0000008d, 5'd11, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031a, 5'd4, 27'h000002c3, 5'd21, 27'h00000303, 32'h00000400,
  1'd1,  5'd14, 27'h000002d5, 5'd14, 27'h00000392, 5'd5, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c1, 5'd14, 27'h00000107, 5'd13, 27'h00000142, 32'h00000400,
  1'd1,  5'd11, 27'h0000023c, 5'd11, 27'h00000276, 5'd22, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000031, 5'd25, 27'h0000033a, 5'd1, 27'h000003d8, 32'h00000400,
  1'd1,  5'd12, 27'h00000027, 5'd22, 27'h00000030, 5'd11, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000167, 5'd21, 27'h00000037, 5'd22, 27'h00000126, 32'h00000400,
  1'd1,  5'd25, 27'h00000232, 5'd1, 27'h00000272, 5'd0, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000103, 5'd2, 27'h0000028f, 5'd10, 27'h00000196, 32'h00000400,
  1'd1,  5'd23, 27'h00000304, 5'd3, 27'h0000039e, 5'd23, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000378, 5'd10, 27'h0000036e, 5'd2, 27'h000003ab, 32'h00000400,
  1'd1,  5'd25, 27'h00000010, 5'd11, 27'h000001d2, 5'd10, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000dd, 5'd13, 27'h00000244, 5'd24, 27'h000000b5, 32'h00000400,
  1'd1,  5'd25, 27'h00000301, 5'd22, 27'h000002a4, 5'd3, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000332, 5'd24, 27'h000000c2, 5'd13, 27'h00000047, 32'h00000400,
  1'd1,  5'd21, 27'h00000125, 5'd24, 27'h0000013d, 5'd21, 27'h00000242, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000240, 5'd3, 27'h000001ba, 5'd9, 27'h0000038e, 32'h00000400,
  1'd1,  5'd3, 27'h00000011, 5'd1, 27'h0000014f, 5'd18, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003ce, 5'd2, 27'h00000089, 5'd26, 27'h0000037a, 32'h00000400,
  1'd1,  5'd5, 27'h00000055, 5'd11, 27'h00000153, 5'd7, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000351, 5'd13, 27'h0000025c, 5'd15, 27'h00000222, 32'h00000400,
  1'd1,  5'd4, 27'h00000207, 5'd13, 27'h00000049, 5'd29, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b0, 5'd22, 27'h00000395, 5'd9, 27'h00000394, 32'h00000400,
  1'd1,  5'd2, 27'h00000009, 5'd22, 27'h0000021c, 5'd17, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000022e, 5'd21, 27'h000000fc, 5'd30, 27'h00000283, 32'h00000400,
  1'd1,  5'd15, 27'h000001a0, 5'd4, 27'h000000fb, 5'd5, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000332, 5'd4, 27'h00000116, 5'd19, 27'h00000022, 32'h00000400,
  1'd1,  5'd12, 27'h00000245, 5'd2, 27'h0000010d, 5'd28, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f1, 5'd14, 27'h00000129, 5'd5, 27'h0000017a, 32'h00000400,
  1'd1,  5'd13, 27'h000001bb, 5'd12, 27'h000000d9, 5'd18, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001f2, 5'd14, 27'h000003b1, 5'd27, 27'h000001bd, 32'h00000400,
  1'd1,  5'd13, 27'h00000259, 5'd23, 27'h0000005c, 5'd6, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000341, 5'd23, 27'h00000352, 5'd16, 27'h0000033a, 32'h00000400,
  1'd1,  5'd13, 27'h000002da, 5'd23, 27'h0000038e, 5'd28, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000257, 5'd0, 27'h00000056, 5'd8, 27'h000000dd, 32'h00000400,
  1'd1,  5'd22, 27'h00000083, 5'd5, 27'h0000001f, 5'd17, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000366, 5'd3, 27'h000003ab, 5'd29, 27'h00000350, 32'h00000400,
  1'd1,  5'd22, 27'h000002c8, 5'd14, 27'h00000100, 5'd9, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d9, 5'd14, 27'h000001df, 5'd17, 27'h00000046, 32'h00000400,
  1'd1,  5'd21, 27'h00000309, 5'd11, 27'h000000c3, 5'd29, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000027d, 5'd24, 27'h00000163, 5'd8, 27'h0000009f, 32'h00000400,
  1'd1,  5'd22, 27'h000001c7, 5'd21, 27'h0000022c, 5'd18, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000026, 5'd23, 27'h000000c3, 5'd27, 27'h00000065, 32'h00000400,
  1'd1,  5'd4, 27'h0000034d, 5'd5, 27'h000002c4, 5'd4, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000206, 5'd9, 27'h000002fa, 5'd14, 27'h00000304, 32'h00000400,
  1'd1,  5'd4, 27'h000000ec, 5'd7, 27'h00000055, 5'd22, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000038e, 5'd19, 27'h0000034a, 5'd2, 27'h00000271, 32'h00000400,
  1'd1,  5'd3, 27'h000002a1, 5'd16, 27'h00000328, 5'd10, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000030c, 5'd16, 27'h00000203, 5'd21, 27'h000000c0, 32'h00000400,
  1'd1,  5'd3, 27'h000000e9, 5'd30, 27'h0000027f, 5'd4, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ba, 5'd29, 27'h0000030d, 5'd12, 27'h0000002d, 32'h00000400,
  1'd1,  5'd4, 27'h0000039e, 5'd27, 27'h00000305, 5'd25, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003de, 5'd5, 27'h000002d5, 5'd2, 27'h000001db, 32'h00000400,
  1'd1,  5'd10, 27'h0000028d, 5'd9, 27'h00000267, 5'd12, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000059, 5'd7, 27'h0000031c, 5'd21, 27'h00000299, 32'h00000400,
  1'd1,  5'd14, 27'h0000014f, 5'd18, 27'h00000269, 5'd2, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c5, 5'd18, 27'h000001ef, 5'd11, 27'h00000107, 32'h00000400,
  1'd1,  5'd11, 27'h00000003, 5'd17, 27'h000003c0, 5'd22, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003bc, 5'd26, 27'h000003eb, 5'd1, 27'h000000bb, 32'h00000400,
  1'd1,  5'd13, 27'h00000053, 5'd30, 27'h00000099, 5'd13, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000249, 5'd28, 27'h0000027d, 5'd21, 27'h00000391, 32'h00000400,
  1'd1,  5'd22, 27'h00000325, 5'd9, 27'h0000030c, 5'd3, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002cc, 5'd9, 27'h000003ef, 5'd14, 27'h000000ef, 32'h00000400,
  1'd1,  5'd20, 27'h000003ec, 5'd9, 27'h00000184, 5'd22, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000247, 5'd16, 27'h00000259, 5'd4, 27'h00000230, 32'h00000400,
  1'd1,  5'd21, 27'h0000023e, 5'd16, 27'h00000107, 5'd15, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000003d, 5'd17, 27'h00000337, 5'd23, 27'h00000106, 32'h00000400,
  1'd1,  5'd23, 27'h0000021c, 5'd30, 27'h00000265, 5'd4, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000232, 5'd29, 27'h000001fe, 5'd12, 27'h000000b2, 32'h00000400,
  1'd1,  5'd24, 27'h0000021f, 5'd26, 27'h0000022d, 5'd25, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000f5, 5'd9, 27'h000002be, 5'd5, 27'h00000184, 32'h00000400,
  1'd1,  5'd3, 27'h000003af, 5'd9, 27'h000002e0, 5'd15, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000016, 5'd6, 27'h000000b7, 5'd26, 27'h00000130, 32'h00000400,
  1'd1,  5'd2, 27'h000002ee, 5'd16, 27'h00000124, 5'd8, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000085, 5'd17, 27'h00000394, 5'd19, 27'h00000269, 32'h00000400,
  1'd1,  5'd3, 27'h000001c4, 5'd19, 27'h00000119, 5'd30, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000064, 5'd28, 27'h00000040, 5'd5, 27'h000003bb, 32'h00000400,
  1'd1,  5'd3, 27'h00000304, 5'd29, 27'h000001cf, 5'd16, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000013, 5'd28, 27'h000001a5, 5'd30, 27'h000003bb, 32'h00000400,
  1'd1,  5'd14, 27'h000003a9, 5'd7, 27'h00000058, 5'd8, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000006f, 5'd9, 27'h00000026, 5'd16, 27'h00000193, 32'h00000400,
  1'd1,  5'd12, 27'h00000382, 5'd8, 27'h000002a6, 5'd26, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000371, 5'd17, 27'h000001c7, 5'd6, 27'h00000342, 32'h00000400,
  1'd1,  5'd14, 27'h00000091, 5'd18, 27'h000000cc, 5'd18, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000035d, 5'd19, 27'h000000f8, 5'd27, 27'h000001b7, 32'h00000400,
  1'd1,  5'd12, 27'h00000271, 5'd26, 27'h000003e3, 5'd8, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000166, 5'd26, 27'h000003df, 5'd16, 27'h00000039, 32'h00000400,
  1'd1,  5'd15, 27'h000001f8, 5'd26, 27'h0000022a, 5'd29, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000021, 5'd9, 27'h00000317, 5'd10, 27'h00000088, 32'h00000400,
  1'd1,  5'd24, 27'h000003e1, 5'd5, 27'h000003fb, 5'd17, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d0, 5'd5, 27'h00000380, 5'd26, 27'h0000009d, 32'h00000400,
  1'd1,  5'd25, 27'h00000216, 5'd16, 27'h0000026a, 5'd9, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000008b, 5'd19, 27'h000003d2, 5'd15, 27'h000003e3, 32'h00000400,
  1'd1,  5'd24, 27'h00000346, 5'd18, 27'h0000033f, 5'd30, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003b3, 5'd27, 27'h00000371, 5'd5, 27'h00000362, 32'h00000400,
  1'd1,  5'd22, 27'h00000249, 5'd26, 27'h00000172, 5'd17, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001db, 5'd29, 27'h0000039f, 5'd26, 27'h00000391, 32'h00000400,
  1'd1,  5'd8, 27'h00000075, 5'd4, 27'h000001b8, 5'd8, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000007d, 5'd4, 27'h0000004d, 5'd17, 27'h00000033, 32'h00000400,
  1'd1,  5'd9, 27'h000003b7, 5'd3, 27'h000001dd, 5'd29, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000269, 5'd14, 27'h000000e0, 5'd0, 27'h00000243, 32'h00000400,
  1'd1,  5'd7, 27'h00000033, 5'd11, 27'h00000289, 5'd13, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002e3, 5'd13, 27'h00000016, 5'd21, 27'h000002e2, 32'h00000400,
  1'd1,  5'd10, 27'h00000136, 5'd25, 27'h0000005e, 5'd1, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000017e, 5'd20, 27'h000002ba, 5'd12, 27'h00000302, 32'h00000400,
  1'd1,  5'd9, 27'h000002ba, 5'd22, 27'h000003ae, 5'd22, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021f, 5'd2, 27'h00000095, 5'd6, 27'h0000027a, 32'h00000400,
  1'd1,  5'd17, 27'h00000212, 5'd3, 27'h00000087, 5'd17, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000385, 5'd4, 27'h000001fd, 5'd27, 27'h00000387, 32'h00000400,
  1'd1,  5'd20, 27'h000000c9, 5'd13, 27'h00000107, 5'd0, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000221, 5'd11, 27'h0000032f, 5'd13, 27'h000003eb, 32'h00000400,
  1'd1,  5'd17, 27'h000002bc, 5'd11, 27'h00000380, 5'd21, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000152, 5'd22, 27'h0000003d, 5'd4, 27'h000000be, 32'h00000400,
  1'd1,  5'd18, 27'h00000133, 5'd25, 27'h000002f2, 5'd15, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d6, 5'd23, 27'h000002f1, 5'd21, 27'h00000395, 32'h00000400,
  1'd1,  5'd29, 27'h000003ea, 5'd1, 27'h0000032e, 5'd1, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000312, 5'd2, 27'h000002ab, 5'd14, 27'h00000227, 32'h00000400,
  1'd1,  5'd27, 27'h000001e6, 5'd2, 27'h0000036c, 5'd21, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000020c, 5'd12, 27'h00000285, 5'd2, 27'h00000085, 32'h00000400,
  1'd1,  5'd28, 27'h000001db, 5'd11, 27'h0000018b, 5'd14, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002ab, 5'd11, 27'h0000029f, 5'd24, 27'h00000334, 32'h00000400,
  1'd1,  5'd28, 27'h0000012d, 5'd21, 27'h00000334, 5'd3, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000215, 5'd23, 27'h0000004a, 5'd11, 27'h00000191, 32'h00000400,
  1'd1,  5'd26, 27'h00000381, 5'd24, 27'h0000007e, 5'd22, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000a6, 5'd0, 27'h00000278, 5'd3, 27'h00000391, 32'h00000400,
  1'd1,  5'd7, 27'h0000014f, 5'd4, 27'h000002ce, 5'd10, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000053, 5'd2, 27'h000000e8, 5'd24, 27'h0000002b, 32'h00000400,
  1'd1,  5'd6, 27'h000001bb, 5'd11, 27'h00000035, 5'd8, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f6, 5'd11, 27'h000003cc, 5'd20, 27'h0000023d, 32'h00000400,
  1'd1,  5'd6, 27'h000003f4, 5'd14, 27'h0000028c, 5'd28, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000333, 5'd21, 27'h000001f6, 5'd6, 27'h000000af, 32'h00000400,
  1'd1,  5'd7, 27'h000002d9, 5'd22, 27'h000001bc, 5'd17, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000ff, 5'd21, 27'h00000112, 5'd26, 27'h000003be, 32'h00000400,
  1'd1,  5'd17, 27'h00000180, 5'd4, 27'h000001b6, 5'd0, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000035f, 5'd2, 27'h000002cd, 5'd10, 27'h000003ac, 32'h00000400,
  1'd1,  5'd16, 27'h00000020, 5'd2, 27'h0000015a, 5'd22, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cc, 5'd11, 27'h00000165, 5'd5, 27'h000003e1, 32'h00000400,
  1'd1,  5'd16, 27'h00000043, 5'd13, 27'h00000220, 5'd20, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000fa, 5'd11, 27'h0000015d, 5'd26, 27'h00000306, 32'h00000400,
  1'd1,  5'd16, 27'h0000012e, 5'd22, 27'h00000293, 5'd9, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001e, 5'd21, 27'h0000013f, 5'd16, 27'h0000016c, 32'h00000400,
  1'd1,  5'd17, 27'h000003a1, 5'd24, 27'h0000022f, 5'd26, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b2, 5'd1, 27'h000002f5, 5'd5, 27'h00000339, 32'h00000400,
  1'd1,  5'd28, 27'h000003d1, 5'd1, 27'h0000017a, 5'd20, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000fc, 5'd1, 27'h0000016c, 5'd30, 27'h000002c3, 32'h00000400,
  1'd1,  5'd27, 27'h0000023f, 5'd12, 27'h00000012, 5'd6, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000024e, 5'd13, 27'h00000198, 5'd16, 27'h00000052, 32'h00000400,
  1'd1,  5'd29, 27'h00000391, 5'd11, 27'h000002eb, 5'd28, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e9, 5'd20, 27'h000003a9, 5'd9, 27'h000002b0, 32'h00000400,
  1'd1,  5'd26, 27'h000001f2, 5'd22, 27'h00000259, 5'd15, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000213, 5'd22, 27'h000003cf, 5'd27, 27'h00000046, 32'h00000400,
  1'd1,  5'd10, 27'h00000027, 5'd5, 27'h000002c8, 5'd1, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f1, 5'd7, 27'h000003e2, 5'd12, 27'h000001c1, 32'h00000400,
  1'd1,  5'd10, 27'h00000049, 5'd10, 27'h000000b4, 5'd25, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002b9, 5'd19, 27'h0000013f, 5'd4, 27'h000003e9, 32'h00000400,
  1'd1,  5'd7, 27'h00000395, 5'd15, 27'h00000232, 5'd15, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000115, 5'd18, 27'h000000d1, 5'd22, 27'h00000354, 32'h00000400,
  1'd1,  5'd6, 27'h000003dc, 5'd27, 27'h0000038d, 5'd5, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000029, 5'd26, 27'h000000df, 5'd14, 27'h0000007a, 32'h00000400,
  1'd1,  5'd8, 27'h000002a4, 5'd28, 27'h000000c9, 5'd21, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000052, 5'd6, 27'h00000106, 5'd1, 27'h00000077, 32'h00000400,
  1'd1,  5'd18, 27'h00000152, 5'd7, 27'h000001a8, 5'd15, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000050, 5'd9, 27'h000002d2, 5'd21, 27'h000002c5, 32'h00000400,
  1'd1,  5'd18, 27'h0000022c, 5'd15, 27'h000003d6, 5'd2, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d2, 5'd16, 27'h000002e8, 5'd11, 27'h00000216, 32'h00000400,
  1'd1,  5'd17, 27'h000001fa, 5'd17, 27'h00000175, 5'd21, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000017c, 5'd26, 27'h000001d8, 5'd2, 27'h0000030c, 32'h00000400,
  1'd1,  5'd20, 27'h0000008a, 5'd27, 27'h000002c1, 5'd15, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000024d, 5'd27, 27'h00000133, 5'd24, 27'h00000094, 32'h00000400,
  1'd1,  5'd30, 27'h000000d4, 5'd9, 27'h0000023f, 5'd4, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000013b, 5'd7, 27'h000001ad, 5'd12, 27'h000003ce, 32'h00000400,
  1'd1,  5'd28, 27'h000000fa, 5'd5, 27'h00000117, 5'd23, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b5, 5'd18, 27'h00000188, 5'd1, 27'h000002dd, 32'h00000400,
  1'd1,  5'd26, 27'h000002f6, 5'd19, 27'h000000b3, 5'd13, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000229, 5'd17, 27'h00000368, 5'd22, 27'h00000325, 32'h00000400,
  1'd1,  5'd28, 27'h00000007, 5'd30, 27'h00000358, 5'd0, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000010d, 5'd25, 27'h0000038d, 5'd12, 27'h00000382, 32'h00000400,
  1'd1,  5'd27, 27'h000000a6, 5'd29, 27'h0000008a, 5'd21, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000020e, 5'd5, 27'h00000299, 5'd5, 27'h000003dc, 32'h00000400,
  1'd1,  5'd5, 27'h0000031b, 5'd6, 27'h000002f5, 5'd18, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d8, 5'd7, 27'h000003a2, 5'd26, 27'h00000318, 32'h00000400,
  1'd1,  5'd8, 27'h0000033a, 5'd18, 27'h00000047, 5'd8, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021e, 5'd16, 27'h00000088, 5'd19, 27'h00000296, 32'h00000400,
  1'd1,  5'd5, 27'h0000023d, 5'd15, 27'h0000036e, 5'd28, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000003b, 5'd30, 27'h0000025b, 5'd9, 27'h00000027, 32'h00000400,
  1'd1,  5'd5, 27'h00000233, 5'd28, 27'h000002fa, 5'd15, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000039c, 5'd26, 27'h00000265, 5'd28, 27'h000000b5, 32'h00000400,
  1'd1,  5'd19, 27'h0000001f, 5'd6, 27'h0000026d, 5'd8, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000101, 5'd5, 27'h000002a2, 5'd20, 27'h00000066, 32'h00000400,
  1'd1,  5'd18, 27'h000000ea, 5'd5, 27'h000002bd, 5'd30, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a1, 5'd18, 27'h000002b2, 5'd7, 27'h00000328, 32'h00000400,
  1'd1,  5'd16, 27'h00000003, 5'd17, 27'h0000001c, 5'd16, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d5, 5'd18, 27'h00000166, 5'd30, 27'h0000012e, 32'h00000400,
  1'd1,  5'd18, 27'h00000309, 5'd26, 27'h0000007d, 5'd6, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001cd, 5'd28, 27'h000002a3, 5'd16, 27'h000003a5, 32'h00000400,
  1'd1,  5'd16, 27'h00000396, 5'd29, 27'h00000043, 5'd30, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000004d, 5'd6, 27'h00000339, 5'd7, 27'h00000340, 32'h00000400,
  1'd1,  5'd29, 27'h000003d8, 5'd6, 27'h0000033e, 5'd16, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000038d, 5'd7, 27'h000001f0, 5'd28, 27'h000001f8, 32'h00000400,
  1'd1,  5'd28, 27'h000001a6, 5'd15, 27'h0000037d, 5'd9, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002ba, 5'd18, 27'h00000067, 5'd18, 27'h0000017a, 32'h00000400,
  1'd1,  5'd30, 27'h000002c4, 5'd17, 27'h0000028f, 5'd29, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e8, 5'd27, 27'h000001da, 5'd7, 27'h000002a0, 32'h00000400,
  1'd1,  5'd30, 27'h000002cc, 5'd27, 27'h00000172, 5'd17, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003da, 5'd30, 27'h000002ba, 5'd28, 27'h000000ca, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001e9, 5'd0, 27'h00000199, 5'd1, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000e3, 5'd2, 27'h000001dc, 5'd12, 27'h0000004a, 32'h00000400,
  1'd1,  5'd0, 27'h00000033, 5'd0, 27'h00000311, 5'd25, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000001b, 5'd14, 27'h0000011a, 5'd2, 27'h0000014e, 32'h00000400,
  1'd1,  5'd3, 27'h00000244, 5'd13, 27'h00000166, 5'd12, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000004b, 5'd10, 27'h00000369, 5'd21, 27'h00000026, 32'h00000400,
  1'd1,  5'd1, 27'h0000017e, 5'd22, 27'h00000001, 5'd1, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000035, 5'd24, 27'h000002dd, 5'd14, 27'h0000028f, 32'h00000400,
  1'd1,  5'd1, 27'h000001b9, 5'd24, 27'h000000a2, 5'd23, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003b7, 5'd0, 27'h00000131, 5'd0, 27'h000002bd, 32'h00000400,
  1'd1,  5'd12, 27'h00000070, 5'd4, 27'h00000362, 5'd13, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e3, 5'd1, 27'h000003ea, 5'd24, 27'h000002d3, 32'h00000400,
  1'd1,  5'd13, 27'h0000022f, 5'd10, 27'h000001bb, 5'd3, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003a5, 5'd11, 27'h000001ef, 5'd12, 27'h00000207, 32'h00000400,
  1'd1,  5'd11, 27'h000001d1, 5'd11, 27'h000002f4, 5'd24, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000024c, 5'd22, 27'h0000039b, 5'd2, 27'h000003e8, 32'h00000400,
  1'd1,  5'd13, 27'h00000073, 5'd23, 27'h0000028e, 5'd13, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000039c, 5'd23, 27'h00000174, 5'd24, 27'h0000011d, 32'h00000400,
  1'd1,  5'd22, 27'h000002ae, 5'd0, 27'h00000187, 5'd0, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002b8, 5'd3, 27'h00000182, 5'd12, 27'h000000c9, 32'h00000400,
  1'd1,  5'd23, 27'h0000014b, 5'd1, 27'h000000b9, 5'd24, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000003e, 5'd12, 27'h00000350, 5'd3, 27'h000001ed, 32'h00000400,
  1'd1,  5'd22, 27'h000003f3, 5'd10, 27'h00000308, 5'd14, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000027d, 5'd13, 27'h000000c1, 5'd24, 27'h000003a0, 32'h00000400,
  1'd1,  5'd23, 27'h00000205, 5'd23, 27'h000000e4, 5'd4, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000217, 5'd24, 27'h00000359, 5'd14, 27'h00000240, 32'h00000400,
  1'd1,  5'd24, 27'h00000008, 5'd21, 27'h00000320, 5'd23, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000c9, 5'd3, 27'h00000254, 5'd5, 27'h00000321, 32'h00000400,
  1'd1,  5'd3, 27'h00000335, 5'd1, 27'h0000005b, 5'd17, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000046, 5'd0, 27'h00000199, 5'd28, 27'h0000038a, 32'h00000400,
  1'd1,  5'd3, 27'h000003bb, 5'd12, 27'h00000184, 5'd6, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000292, 5'd11, 27'h0000023b, 5'd15, 27'h00000338, 32'h00000400,
  1'd1,  5'd0, 27'h00000299, 5'd10, 27'h0000024e, 5'd28, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000036d, 5'd22, 27'h000001af, 5'd9, 27'h00000071, 32'h00000400,
  1'd1,  5'd1, 27'h00000082, 5'd22, 27'h00000355, 5'd20, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001be, 5'd23, 27'h000001fb, 5'd27, 27'h00000234, 32'h00000400,
  1'd1,  5'd13, 27'h000000bd, 5'd1, 27'h0000013c, 5'd9, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000017c, 5'd4, 27'h0000034e, 5'd19, 27'h000001b0, 32'h00000400,
  1'd1,  5'd12, 27'h00000077, 5'd4, 27'h00000353, 5'd29, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000338, 5'd14, 27'h000000e9, 5'd9, 27'h00000147, 32'h00000400,
  1'd1,  5'd12, 27'h000002b0, 5'd12, 27'h0000011f, 5'd18, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c0, 5'd12, 27'h0000035e, 5'd28, 27'h00000311, 32'h00000400,
  1'd1,  5'd12, 27'h000002db, 5'd22, 27'h00000299, 5'd8, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001c2, 5'd23, 27'h000001d8, 5'd16, 27'h000002b1, 32'h00000400,
  1'd1,  5'd12, 27'h000003ec, 5'd21, 27'h000002c1, 5'd28, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e5, 5'd1, 27'h000002d1, 5'd9, 27'h000001a7, 32'h00000400,
  1'd1,  5'd24, 27'h000001f2, 5'd2, 27'h00000260, 5'd19, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001db, 5'd1, 27'h000000f7, 5'd26, 27'h000003c4, 32'h00000400,
  1'd1,  5'd21, 27'h00000287, 5'd10, 27'h00000180, 5'd7, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000002, 5'd14, 27'h000003df, 5'd19, 27'h00000008, 32'h00000400,
  1'd1,  5'd23, 27'h000003bc, 5'd11, 27'h000000a5, 5'd28, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031e, 5'd21, 27'h000001e3, 5'd6, 27'h00000393, 32'h00000400,
  1'd1,  5'd22, 27'h00000058, 5'd22, 27'h00000300, 5'd19, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000006a, 5'd25, 27'h00000020, 5'd28, 27'h00000120, 32'h00000400,
  1'd1,  5'd0, 27'h00000341, 5'd9, 27'h000003d8, 5'd2, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a3, 5'd5, 27'h000001d2, 5'd11, 27'h00000279, 32'h00000400,
  1'd1,  5'd4, 27'h0000029e, 5'd9, 27'h00000180, 5'd25, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002e6, 5'd18, 27'h000001b2, 5'd0, 27'h00000032, 32'h00000400,
  1'd1,  5'd2, 27'h0000025c, 5'd18, 27'h000000f7, 5'd15, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000022, 5'd16, 27'h000002e9, 5'd22, 27'h00000130, 32'h00000400,
  1'd1,  5'd4, 27'h000002f5, 5'd29, 27'h0000003e, 5'd0, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c7, 5'd27, 27'h00000305, 5'd10, 27'h00000198, 32'h00000400,
  1'd1,  5'd0, 27'h0000011e, 5'd27, 27'h00000289, 5'd21, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b6, 5'd8, 27'h00000247, 5'd3, 27'h0000006b, 32'h00000400,
  1'd1,  5'd13, 27'h00000113, 5'd7, 27'h00000385, 5'd14, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000192, 5'd5, 27'h00000295, 5'd25, 27'h000000ce, 32'h00000400,
  1'd1,  5'd13, 27'h00000291, 5'd18, 27'h0000011f, 5'd0, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000204, 5'd19, 27'h00000230, 5'd13, 27'h0000006c, 32'h00000400,
  1'd1,  5'd12, 27'h000003f1, 5'd20, 27'h000001ab, 5'd23, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000226, 5'd26, 27'h00000123, 5'd0, 27'h0000017f, 32'h00000400,
  1'd1,  5'd11, 27'h00000026, 5'd26, 27'h00000198, 5'd14, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000350, 5'd29, 27'h000001e0, 5'd24, 27'h0000014b, 32'h00000400,
  1'd1,  5'd22, 27'h000002f8, 5'd7, 27'h0000023e, 5'd1, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000011c, 5'd10, 27'h00000026, 5'd13, 27'h0000027a, 32'h00000400,
  1'd1,  5'd21, 27'h00000216, 5'd5, 27'h000000c2, 5'd20, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038b, 5'd15, 27'h0000029f, 5'd4, 27'h000002eb, 32'h00000400,
  1'd1,  5'd23, 27'h00000066, 5'd17, 27'h0000005e, 5'd11, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000363, 5'd19, 27'h00000040, 5'd20, 27'h00000381, 32'h00000400,
  1'd1,  5'd23, 27'h00000136, 5'd30, 27'h000001c1, 5'd3, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000213, 5'd29, 27'h00000110, 5'd12, 27'h00000068, 32'h00000400,
  1'd1,  5'd25, 27'h000000b5, 5'd29, 27'h00000240, 5'd24, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000018e, 5'd7, 27'h000003bf, 5'd5, 27'h00000278, 32'h00000400,
  1'd1,  5'd3, 27'h000001db, 5'd8, 27'h000001e6, 5'd18, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017c, 5'd6, 27'h00000190, 5'd26, 27'h000003dc, 32'h00000400,
  1'd1,  5'd0, 27'h0000021d, 5'd20, 27'h000001e8, 5'd9, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000008e, 5'd16, 27'h00000193, 5'd19, 27'h000003ab, 32'h00000400,
  1'd1,  5'd0, 27'h0000014a, 5'd17, 27'h000000d2, 5'd25, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000362, 5'd30, 27'h000000b7, 5'd7, 27'h000002af, 32'h00000400,
  1'd1,  5'd4, 27'h00000043, 5'd30, 27'h000000b0, 5'd16, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000138, 5'd30, 27'h0000012a, 5'd27, 27'h0000010e, 32'h00000400,
  1'd1,  5'd10, 27'h00000347, 5'd7, 27'h00000260, 5'd9, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f1, 5'd9, 27'h00000186, 5'd19, 27'h000001c0, 32'h00000400,
  1'd1,  5'd14, 27'h0000015f, 5'd9, 27'h00000046, 5'd29, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000a2, 5'd18, 27'h00000378, 5'd6, 27'h000000a6, 32'h00000400,
  1'd1,  5'd15, 27'h00000114, 5'd16, 27'h00000354, 5'd19, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000164, 5'd20, 27'h00000127, 5'd27, 27'h00000138, 32'h00000400,
  1'd1,  5'd10, 27'h00000372, 5'd27, 27'h0000024f, 5'd6, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017b, 5'd30, 27'h0000019a, 5'd19, 27'h00000193, 32'h00000400,
  1'd1,  5'd15, 27'h000001ff, 5'd29, 27'h00000063, 5'd30, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002f5, 5'd8, 27'h000002b9, 5'd9, 27'h000002fd, 32'h00000400,
  1'd1,  5'd24, 27'h0000014a, 5'd6, 27'h0000001e, 5'd18, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a9, 5'd8, 27'h000003f1, 5'd27, 27'h000003dd, 32'h00000400,
  1'd1,  5'd24, 27'h00000034, 5'd17, 27'h000001d6, 5'd7, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002a7, 5'd19, 27'h000003fc, 5'd15, 27'h000003c2, 32'h00000400,
  1'd1,  5'd21, 27'h000000ef, 5'd16, 27'h00000065, 5'd30, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000037, 5'd27, 27'h000000bf, 5'd8, 27'h00000288, 32'h00000400,
  1'd1,  5'd23, 27'h00000343, 5'd29, 27'h000003e8, 5'd17, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000129, 5'd26, 27'h00000001, 5'd28, 27'h0000020c, 32'h00000400,
  1'd1,  5'd10, 27'h00000097, 5'd1, 27'h000003a1, 5'd7, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000af, 5'd0, 27'h0000000b, 5'd17, 27'h00000045, 32'h00000400,
  1'd1,  5'd6, 27'h0000033d, 5'd2, 27'h000003bc, 5'd30, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000016, 5'd14, 27'h0000020b, 5'd1, 27'h00000243, 32'h00000400,
  1'd1,  5'd7, 27'h000002e2, 5'd11, 27'h00000165, 5'd15, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ec, 5'd15, 27'h0000007d, 5'd24, 27'h0000014f, 32'h00000400,
  1'd1,  5'd6, 27'h00000264, 5'd24, 27'h000002e7, 5'd2, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000354, 5'd21, 27'h00000365, 5'd14, 27'h00000228, 32'h00000400,
  1'd1,  5'd7, 27'h00000392, 5'd23, 27'h000000af, 5'd22, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000294, 5'd2, 27'h000001b2, 5'd5, 27'h0000013c, 32'h00000400,
  1'd1,  5'd17, 27'h000002dd, 5'd1, 27'h00000007, 5'd19, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000117, 5'd0, 27'h000000e2, 5'd27, 27'h0000020b, 32'h00000400,
  1'd1,  5'd19, 27'h0000005e, 5'd12, 27'h00000346, 5'd0, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f5, 5'd15, 27'h0000012e, 5'd11, 27'h000001d7, 32'h00000400,
  1'd1,  5'd19, 27'h0000007b, 5'd12, 27'h0000039b, 5'd22, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000218, 5'd21, 27'h00000329, 5'd0, 27'h00000172, 32'h00000400,
  1'd1,  5'd16, 27'h0000001b, 5'd22, 27'h000003d5, 5'd15, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a3, 5'd24, 27'h000003f0, 5'd22, 27'h00000348, 32'h00000400,
  1'd1,  5'd29, 27'h000001be, 5'd0, 27'h000002f4, 5'd3, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000304, 5'd4, 27'h000003e4, 5'd14, 27'h0000019c, 32'h00000400,
  1'd1,  5'd28, 27'h00000168, 5'd4, 27'h00000005, 5'd22, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000138, 5'd11, 27'h000002db, 5'd4, 27'h00000301, 32'h00000400,
  1'd1,  5'd26, 27'h000001b7, 5'd11, 27'h000000a6, 5'd13, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000023, 5'd10, 27'h0000035b, 5'd23, 27'h0000011e, 32'h00000400,
  1'd1,  5'd27, 27'h0000005d, 5'd25, 27'h0000024f, 5'd3, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000395, 5'd23, 27'h00000005, 5'd12, 27'h000000c1, 32'h00000400,
  1'd1,  5'd27, 27'h00000391, 5'd21, 27'h00000205, 5'd21, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e9, 5'd0, 27'h00000112, 5'd3, 27'h00000212, 32'h00000400,
  1'd1,  5'd9, 27'h0000009c, 5'd3, 27'h00000096, 5'd15, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000155, 5'd4, 27'h000003a2, 5'd22, 27'h000003cf, 32'h00000400,
  1'd1,  5'd7, 27'h0000030a, 5'd15, 27'h00000150, 5'd5, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003d3, 5'd12, 27'h00000005, 5'd16, 27'h00000077, 32'h00000400,
  1'd1,  5'd6, 27'h000003e9, 5'd14, 27'h0000030f, 5'd29, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000030f, 5'd20, 27'h000003a1, 5'd6, 27'h000000ca, 32'h00000400,
  1'd1,  5'd9, 27'h000003d4, 5'd25, 27'h0000011a, 5'd17, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000119, 5'd24, 27'h00000227, 5'd26, 27'h00000022, 32'h00000400,
  1'd1,  5'd20, 27'h000001c8, 5'd1, 27'h00000060, 5'd2, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000100, 5'd4, 27'h000001e0, 5'd11, 27'h000000cc, 32'h00000400,
  1'd1,  5'd20, 27'h0000014a, 5'd0, 27'h0000025a, 5'd23, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001d0, 5'd14, 27'h000003ad, 5'd10, 27'h000000ac, 32'h00000400,
  1'd1,  5'd16, 27'h00000390, 5'd11, 27'h000003a5, 5'd19, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000092, 5'd11, 27'h0000005f, 5'd26, 27'h000002a2, 32'h00000400,
  1'd1,  5'd18, 27'h000002f4, 5'd21, 27'h00000311, 5'd9, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000013c, 5'd21, 27'h00000367, 5'd18, 27'h000001af, 32'h00000400,
  1'd1,  5'd17, 27'h00000039, 5'd23, 27'h0000038c, 5'd30, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a3, 5'd0, 27'h000000bc, 5'd5, 27'h00000153, 32'h00000400,
  1'd1,  5'd28, 27'h00000152, 5'd1, 27'h0000006b, 5'd20, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ed, 5'd2, 27'h00000379, 5'd26, 27'h000000ac, 32'h00000400,
  1'd1,  5'd26, 27'h0000023d, 5'd11, 27'h0000034e, 5'd7, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d3, 5'd13, 27'h000000d4, 5'd18, 27'h000000b0, 32'h00000400,
  1'd1,  5'd27, 27'h00000271, 5'd11, 27'h0000026d, 5'd28, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000018, 5'd24, 27'h00000126, 5'd7, 27'h000001ba, 32'h00000400,
  1'd1,  5'd28, 27'h0000024b, 5'd23, 27'h0000003d, 5'd16, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000264, 5'd25, 27'h0000006b, 5'd27, 27'h00000115, 32'h00000400,
  1'd1,  5'd7, 27'h000001f3, 5'd10, 27'h00000066, 5'd1, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002f6, 5'd7, 27'h000003c0, 5'd14, 27'h00000393, 32'h00000400,
  1'd1,  5'd6, 27'h00000114, 5'd7, 27'h000001a1, 5'd22, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000275, 5'd17, 27'h00000148, 5'd2, 27'h0000030f, 32'h00000400,
  1'd1,  5'd6, 27'h00000208, 5'd20, 27'h000000ec, 5'd11, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000017d, 5'd15, 27'h00000306, 5'd24, 27'h00000330, 32'h00000400,
  1'd1,  5'd5, 27'h000001e5, 5'd25, 27'h0000037f, 5'd2, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ed, 5'd29, 27'h0000031c, 5'd12, 27'h000003e4, 32'h00000400,
  1'd1,  5'd7, 27'h00000105, 5'd25, 27'h000003ee, 5'd20, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000054, 5'd7, 27'h000002e2, 5'd1, 27'h000002e4, 32'h00000400,
  1'd1,  5'd20, 27'h000000d2, 5'd7, 27'h00000127, 5'd13, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002f3, 5'd5, 27'h000003f2, 5'd21, 27'h000001bb, 32'h00000400,
  1'd1,  5'd17, 27'h00000232, 5'd18, 27'h0000024e, 5'd3, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000016d, 5'd16, 27'h00000192, 5'd11, 27'h00000167, 32'h00000400,
  1'd1,  5'd18, 27'h0000026c, 5'd17, 27'h00000252, 5'd23, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002c0, 5'd25, 27'h0000035b, 5'd4, 27'h00000204, 32'h00000400,
  1'd1,  5'd15, 27'h00000212, 5'd28, 27'h00000229, 5'd13, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ea, 5'd29, 27'h00000358, 5'd23, 27'h000003ea, 32'h00000400,
  1'd1,  5'd26, 27'h00000068, 5'd8, 27'h000001a1, 5'd4, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000309, 5'd8, 27'h00000054, 5'd11, 27'h000000ea, 32'h00000400,
  1'd1,  5'd28, 27'h00000260, 5'd7, 27'h0000012f, 5'd24, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000001a, 5'd20, 27'h0000016d, 5'd1, 27'h0000022e, 32'h00000400,
  1'd1,  5'd29, 27'h0000032b, 5'd17, 27'h000003f1, 5'd15, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000326, 5'd19, 27'h000003c3, 5'd23, 27'h000000ac, 32'h00000400,
  1'd1,  5'd30, 27'h000000b0, 5'd26, 27'h0000007a, 5'd0, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000002b, 5'd26, 27'h00000268, 5'd13, 27'h00000048, 32'h00000400,
  1'd1,  5'd30, 27'h000001bc, 5'd28, 27'h00000061, 5'd23, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d5, 5'd8, 27'h0000018b, 5'd9, 27'h0000005c, 32'h00000400,
  1'd1,  5'd7, 27'h00000032, 5'd10, 27'h00000034, 5'd18, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000038, 5'd9, 27'h00000039, 5'd30, 27'h000002df, 32'h00000400,
  1'd1,  5'd9, 27'h00000377, 5'd16, 27'h000000de, 5'd6, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000395, 5'd17, 27'h00000219, 5'd18, 27'h00000159, 32'h00000400,
  1'd1,  5'd6, 27'h000003c8, 5'd18, 27'h000003bd, 5'd29, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a2, 5'd27, 27'h000002dc, 5'd5, 27'h00000352, 32'h00000400,
  1'd1,  5'd6, 27'h0000019b, 5'd27, 27'h00000069, 5'd17, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ce, 5'd29, 27'h000002cb, 5'd29, 27'h0000039e, 32'h00000400,
  1'd1,  5'd18, 27'h00000050, 5'd6, 27'h000001c2, 5'd5, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000380, 5'd8, 27'h000000ba, 5'd16, 27'h00000159, 32'h00000400,
  1'd1,  5'd19, 27'h00000346, 5'd6, 27'h0000014d, 5'd27, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000007a, 5'd17, 27'h000003ba, 5'd7, 27'h00000113, 32'h00000400,
  1'd1,  5'd16, 27'h0000024a, 5'd16, 27'h00000392, 5'd16, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000065, 5'd17, 27'h000000bb, 5'd30, 27'h000002e2, 32'h00000400,
  1'd1,  5'd17, 27'h0000011d, 5'd28, 27'h0000021d, 5'd6, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000246, 5'd27, 27'h0000029d, 5'd17, 27'h00000140, 32'h00000400,
  1'd1,  5'd19, 27'h000001c1, 5'd28, 27'h000002da, 5'd28, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000028f, 5'd5, 27'h000002df, 5'd6, 27'h00000150, 32'h00000400,
  1'd1,  5'd30, 27'h000003f0, 5'd6, 27'h0000038e, 5'd18, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000027a, 5'd5, 27'h000000c8, 5'd29, 27'h00000001, 32'h00000400,
  1'd1,  5'd26, 27'h0000027f, 5'd18, 27'h000003f3, 5'd6, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024a, 5'd16, 27'h0000002f, 5'd17, 27'h00000287, 32'h00000400,
  1'd1,  5'd27, 27'h0000029d, 5'd19, 27'h00000368, 5'd27, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c5, 5'd27, 27'h0000006c, 5'd5, 27'h000002ad, 32'h00000400,
  1'd1,  5'd27, 27'h00000157, 5'd26, 27'h000001c7, 5'd15, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000357, 5'd29, 27'h00000273, 5'd29, 27'h00000230, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003f9, 5'd1, 27'h000000ab, 5'd3, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000134, 5'd3, 27'h0000031f, 5'd11, 27'h00000233, 32'h00000400,
  1'd1,  5'd0, 27'h0000018f, 5'd2, 27'h000002b7, 5'd23, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000320, 5'd13, 27'h000003a6, 5'd0, 27'h00000342, 32'h00000400,
  1'd1,  5'd2, 27'h000003b7, 5'd12, 27'h0000036f, 5'd13, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ee, 5'd12, 27'h000001bf, 5'd24, 27'h00000110, 32'h00000400,
  1'd1,  5'd4, 27'h0000011d, 5'd21, 27'h000002ae, 5'd1, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000fa, 5'd24, 27'h000001e9, 5'd14, 27'h000003fe, 32'h00000400,
  1'd1,  5'd2, 27'h00000313, 5'd23, 27'h00000266, 5'd24, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f2, 5'd5, 27'h0000006a, 5'd0, 27'h00000391, 32'h00000400,
  1'd1,  5'd11, 27'h000000bc, 5'd2, 27'h0000020c, 5'd13, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000015, 5'd3, 27'h000003cd, 5'd25, 27'h000002d6, 32'h00000400,
  1'd1,  5'd11, 27'h000002ff, 5'd10, 27'h000002aa, 5'd1, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000062, 5'd11, 27'h000000df, 5'd10, 27'h00000350, 32'h00000400,
  1'd1,  5'd11, 27'h00000228, 5'd11, 27'h0000037c, 5'd23, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000342, 5'd21, 27'h00000006, 5'd2, 27'h00000010, 32'h00000400,
  1'd1,  5'd13, 27'h00000105, 5'd24, 27'h00000009, 5'd13, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029b, 5'd23, 27'h0000024d, 5'd22, 27'h000003bf, 32'h00000400,
  1'd1,  5'd22, 27'h000002ca, 5'd3, 27'h0000011c, 5'd1, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003fa, 5'd3, 27'h000003eb, 5'd13, 27'h000001ab, 32'h00000400,
  1'd1,  5'd24, 27'h00000098, 5'd4, 27'h00000377, 5'd22, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003b8, 5'd15, 27'h0000004e, 5'd3, 27'h00000267, 32'h00000400,
  1'd1,  5'd20, 27'h00000336, 5'd14, 27'h00000133, 5'd14, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000036a, 5'd11, 27'h0000022a, 5'd22, 27'h000001b9, 32'h00000400,
  1'd1,  5'd22, 27'h0000029c, 5'd25, 27'h0000032d, 5'd2, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000002c, 5'd22, 27'h000000bd, 5'd11, 27'h000002e3, 32'h00000400,
  1'd1,  5'd22, 27'h00000259, 5'd22, 27'h0000011e, 5'd23, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a2, 5'd3, 27'h000003e5, 5'd7, 27'h00000391, 32'h00000400,
  1'd1,  5'd4, 27'h00000129, 5'd3, 27'h00000283, 5'd18, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a6, 5'd2, 27'h000003df, 5'd25, 27'h000003fa, 32'h00000400,
  1'd1,  5'd1, 27'h00000242, 5'd15, 27'h000001b4, 5'd6, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000035a, 5'd14, 27'h000001dd, 5'd19, 27'h000002dd, 32'h00000400,
  1'd1,  5'd4, 27'h00000270, 5'd11, 27'h00000097, 5'd27, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000018f, 5'd23, 27'h00000311, 5'd5, 27'h000002c4, 32'h00000400,
  1'd1,  5'd1, 27'h000001d9, 5'd24, 27'h00000258, 5'd18, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000280, 5'd24, 27'h000002bd, 5'd29, 27'h0000021f, 32'h00000400,
  1'd1,  5'd14, 27'h000000f7, 5'd4, 27'h000000b6, 5'd5, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000011, 5'd3, 27'h0000004c, 5'd16, 27'h000002e9, 32'h00000400,
  1'd1,  5'd11, 27'h000000e0, 5'd4, 27'h000002dd, 5'd25, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000016c, 5'd11, 27'h000002bb, 5'd9, 27'h000003bf, 32'h00000400,
  1'd1,  5'd14, 27'h000001cd, 5'd13, 27'h00000144, 5'd17, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fb, 5'd14, 27'h0000011e, 5'd29, 27'h00000051, 32'h00000400,
  1'd1,  5'd13, 27'h000003fa, 5'd25, 27'h000000a0, 5'd7, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001da, 5'd24, 27'h000001cd, 5'd16, 27'h0000003f, 32'h00000400,
  1'd1,  5'd12, 27'h00000075, 5'd24, 27'h000001f6, 5'd28, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d2, 5'd1, 27'h000000e0, 5'd7, 27'h0000000a, 32'h00000400,
  1'd1,  5'd24, 27'h000000ac, 5'd4, 27'h000001be, 5'd19, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000161, 5'd1, 27'h00000313, 5'd28, 27'h0000036c, 32'h00000400,
  1'd1,  5'd25, 27'h000001bd, 5'd14, 27'h0000016f, 5'd6, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001f3, 5'd12, 27'h00000106, 5'd16, 27'h000001a0, 32'h00000400,
  1'd1,  5'd25, 27'h00000336, 5'd15, 27'h000001f3, 5'd29, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000001b, 5'd25, 27'h00000132, 5'd9, 27'h0000001f, 32'h00000400,
  1'd1,  5'd24, 27'h00000107, 5'd23, 27'h00000310, 5'd18, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000303, 5'd23, 27'h000002ae, 5'd29, 27'h00000038, 32'h00000400,
  1'd1,  5'd3, 27'h00000384, 5'd8, 27'h00000117, 5'd2, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e8, 5'd8, 27'h000002d3, 5'd14, 27'h000001ab, 32'h00000400,
  1'd1,  5'd4, 27'h00000231, 5'd6, 27'h0000018d, 5'd25, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000018, 5'd18, 27'h00000042, 5'd1, 27'h000003a6, 32'h00000400,
  1'd1,  5'd0, 27'h0000015c, 5'd17, 27'h00000162, 5'd14, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000230, 5'd19, 27'h00000185, 5'd22, 27'h000001ac, 32'h00000400,
  1'd1,  5'd3, 27'h00000129, 5'd29, 27'h000001e6, 5'd1, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000122, 5'd30, 27'h00000311, 5'd15, 27'h00000121, 32'h00000400,
  1'd1,  5'd3, 27'h0000022e, 5'd30, 27'h000001a8, 5'd25, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000084, 5'd9, 27'h000002f7, 5'd3, 27'h00000322, 32'h00000400,
  1'd1,  5'd11, 27'h000002aa, 5'd6, 27'h0000017a, 5'd10, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000268, 5'd5, 27'h000003c8, 5'd22, 27'h000002cc, 32'h00000400,
  1'd1,  5'd14, 27'h000003da, 5'd17, 27'h00000242, 5'd2, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000008a, 5'd19, 27'h00000079, 5'd15, 27'h000001d7, 32'h00000400,
  1'd1,  5'd15, 27'h000001d8, 5'd20, 27'h0000000e, 5'd25, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000094, 5'd28, 27'h00000222, 5'd4, 27'h0000029b, 32'h00000400,
  1'd1,  5'd12, 27'h0000005a, 5'd27, 27'h000001e8, 5'd11, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000182, 5'd30, 27'h00000282, 5'd23, 27'h000001d4, 32'h00000400,
  1'd1,  5'd22, 27'h00000122, 5'd8, 27'h0000017b, 5'd0, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000046, 5'd8, 27'h0000003a, 5'd11, 27'h000003c2, 32'h00000400,
  1'd1,  5'd21, 27'h0000025b, 5'd7, 27'h0000020c, 5'd21, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002da, 5'd19, 27'h0000025e, 5'd1, 27'h000001b6, 32'h00000400,
  1'd1,  5'd21, 27'h000001cc, 5'd19, 27'h00000359, 5'd13, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001e4, 5'd19, 27'h00000103, 5'd23, 27'h00000075, 32'h00000400,
  1'd1,  5'd24, 27'h000003d8, 5'd29, 27'h0000004c, 5'd3, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000138, 5'd27, 27'h000003bb, 5'd11, 27'h00000212, 32'h00000400,
  1'd1,  5'd24, 27'h000003b2, 5'd28, 27'h00000188, 5'd21, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000024d, 5'd9, 27'h00000266, 5'd6, 27'h00000064, 32'h00000400,
  1'd1,  5'd0, 27'h00000347, 5'd6, 27'h0000013e, 5'd16, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000357, 5'd5, 27'h0000036f, 5'd27, 27'h00000054, 32'h00000400,
  1'd1,  5'd1, 27'h00000157, 5'd15, 27'h000003ef, 5'd8, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000003d, 5'd16, 27'h0000035f, 5'd20, 27'h00000217, 32'h00000400,
  1'd1,  5'd1, 27'h00000297, 5'd20, 27'h0000005d, 5'd28, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000195, 5'd29, 27'h00000257, 5'd10, 27'h0000003b, 32'h00000400,
  1'd1,  5'd1, 27'h000002a7, 5'd27, 27'h000001ee, 5'd18, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000144, 5'd30, 27'h000001bf, 5'd26, 27'h00000312, 32'h00000400,
  1'd1,  5'd12, 27'h00000200, 5'd6, 27'h00000367, 5'd7, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000139, 5'd8, 27'h00000291, 5'd17, 27'h000002f9, 32'h00000400,
  1'd1,  5'd14, 27'h0000022e, 5'd7, 27'h000003a6, 5'd30, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000012d, 5'd18, 27'h00000345, 5'd8, 27'h000003bf, 32'h00000400,
  1'd1,  5'd15, 27'h0000007d, 5'd19, 27'h0000030a, 5'd20, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000039c, 5'd17, 27'h000002c4, 5'd30, 27'h000001b3, 32'h00000400,
  1'd1,  5'd15, 27'h0000019d, 5'd29, 27'h00000342, 5'd6, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000029a, 5'd29, 27'h00000374, 5'd17, 27'h000002da, 32'h00000400,
  1'd1,  5'd13, 27'h00000008, 5'd28, 27'h00000095, 5'd28, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b8, 5'd6, 27'h0000019b, 5'd9, 27'h0000039b, 32'h00000400,
  1'd1,  5'd21, 27'h0000019a, 5'd5, 27'h000000bf, 5'd16, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003e5, 5'd9, 27'h00000306, 5'd28, 27'h00000061, 32'h00000400,
  1'd1,  5'd23, 27'h0000012a, 5'd16, 27'h000001fc, 5'd8, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000172, 5'd16, 27'h00000060, 5'd20, 27'h000000a4, 32'h00000400,
  1'd1,  5'd23, 27'h000003eb, 5'd16, 27'h000000f3, 5'd29, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000179, 5'd28, 27'h00000192, 5'd6, 27'h0000037e, 32'h00000400,
  1'd1,  5'd21, 27'h000000ca, 5'd29, 27'h0000035c, 5'd17, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002e7, 5'd28, 27'h000002f0, 5'd27, 27'h000000b8, 32'h00000400,
  1'd1,  5'd7, 27'h000002c4, 5'd1, 27'h000003fe, 5'd9, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000021c, 5'd3, 27'h000003b5, 5'd20, 27'h00000226, 32'h00000400,
  1'd1,  5'd10, 27'h000000a0, 5'd3, 27'h00000382, 5'd30, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a9, 5'd11, 27'h0000019a, 5'd2, 27'h000001eb, 32'h00000400,
  1'd1,  5'd9, 27'h000002f4, 5'd11, 27'h0000007e, 5'd15, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000229, 5'd12, 27'h00000140, 5'd24, 27'h000001a6, 32'h00000400,
  1'd1,  5'd9, 27'h00000188, 5'd23, 27'h0000018d, 5'd1, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000382, 5'd21, 27'h0000013b, 5'd11, 27'h0000033a, 32'h00000400,
  1'd1,  5'd9, 27'h000001e2, 5'd25, 27'h00000167, 5'd21, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000017, 5'd4, 27'h0000005d, 5'd6, 27'h000000c7, 32'h00000400,
  1'd1,  5'd18, 27'h000001be, 5'd1, 27'h000003dd, 5'd18, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ac, 5'd2, 27'h000003ac, 5'd26, 27'h0000031f, 32'h00000400,
  1'd1,  5'd18, 27'h0000000a, 5'd10, 27'h000001fe, 5'd3, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000034c, 5'd10, 27'h00000272, 5'd14, 27'h00000200, 32'h00000400,
  1'd1,  5'd19, 27'h0000038a, 5'd12, 27'h00000383, 5'd22, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000162, 5'd24, 27'h000001ec, 5'd3, 27'h00000173, 32'h00000400,
  1'd1,  5'd19, 27'h00000399, 5'd22, 27'h000001c3, 5'd13, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000004f, 5'd22, 27'h000002e8, 5'd23, 27'h000001f2, 32'h00000400,
  1'd1,  5'd30, 27'h000003f4, 5'd4, 27'h000001c7, 5'd0, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003d1, 5'd3, 27'h00000005, 5'd10, 27'h00000202, 32'h00000400,
  1'd1,  5'd27, 27'h000002c3, 5'd1, 27'h00000349, 5'd22, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000269, 5'd14, 27'h0000034e, 5'd4, 27'h00000100, 32'h00000400,
  1'd1,  5'd29, 27'h000003c7, 5'd12, 27'h0000038e, 5'd10, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000040, 5'd14, 27'h00000336, 5'd25, 27'h000002c8, 32'h00000400,
  1'd1,  5'd28, 27'h0000003c, 5'd21, 27'h0000000a, 5'd0, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c7, 5'd21, 27'h00000092, 5'd10, 27'h00000371, 32'h00000400,
  1'd1,  5'd29, 27'h00000253, 5'd21, 27'h0000018f, 5'd21, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000022f, 5'd0, 27'h000002bf, 5'd2, 27'h0000008c, 32'h00000400,
  1'd1,  5'd8, 27'h0000026f, 5'd2, 27'h00000308, 5'd12, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031b, 5'd2, 27'h0000002b, 5'd21, 27'h000002ee, 32'h00000400,
  1'd1,  5'd10, 27'h0000001a, 5'd15, 27'h000000dd, 5'd8, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f9, 5'd12, 27'h00000388, 5'd17, 27'h0000010b, 32'h00000400,
  1'd1,  5'd5, 27'h0000017b, 5'd14, 27'h00000306, 5'd29, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d5, 5'd24, 27'h000002d7, 5'd5, 27'h000000f5, 32'h00000400,
  1'd1,  5'd5, 27'h00000331, 5'd22, 27'h00000106, 5'd19, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000280, 5'd23, 27'h000001ba, 5'd26, 27'h000003ef, 32'h00000400,
  1'd1,  5'd19, 27'h000001d9, 5'd0, 27'h000001ba, 5'd0, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000018c, 5'd1, 27'h000002c2, 5'd11, 27'h00000215, 32'h00000400,
  1'd1,  5'd20, 27'h0000014d, 5'd0, 27'h0000030c, 5'd21, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e4, 5'd12, 27'h00000051, 5'd6, 27'h000000cc, 32'h00000400,
  1'd1,  5'd18, 27'h0000032a, 5'd13, 27'h0000028e, 5'd17, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000284, 5'd14, 27'h000001c3, 5'd26, 27'h000001a0, 32'h00000400,
  1'd1,  5'd18, 27'h00000223, 5'd25, 27'h0000018e, 5'd6, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003f3, 5'd22, 27'h000003e0, 5'd18, 27'h000003e1, 32'h00000400,
  1'd1,  5'd19, 27'h0000027a, 5'd25, 27'h000001f9, 5'd29, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000054, 5'd3, 27'h00000311, 5'd9, 27'h00000305, 32'h00000400,
  1'd1,  5'd29, 27'h0000029a, 5'd5, 27'h0000006b, 5'd16, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000383, 5'd0, 27'h00000163, 5'd27, 27'h00000057, 32'h00000400,
  1'd1,  5'd26, 27'h000003f8, 5'd15, 27'h00000150, 5'd7, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000193, 5'd11, 27'h000003eb, 5'd20, 27'h00000081, 32'h00000400,
  1'd1,  5'd30, 27'h00000353, 5'd10, 27'h000003c5, 5'd28, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000015a, 5'd24, 27'h000003b0, 5'd9, 27'h000001e2, 32'h00000400,
  1'd1,  5'd28, 27'h00000399, 5'd25, 27'h00000049, 5'd18, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001df, 5'd24, 27'h000003d1, 5'd26, 27'h00000000, 32'h00000400,
  1'd1,  5'd8, 27'h00000062, 5'd7, 27'h000003cf, 5'd1, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000078, 5'd6, 27'h00000115, 5'd14, 27'h000003ea, 32'h00000400,
  1'd1,  5'd5, 27'h00000270, 5'd6, 27'h0000030f, 5'd22, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e5, 5'd17, 27'h00000233, 5'd1, 27'h000001df, 32'h00000400,
  1'd1,  5'd8, 27'h0000006b, 5'd20, 27'h00000111, 5'd12, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002d4, 5'd15, 27'h000002c0, 5'd24, 27'h000003de, 32'h00000400,
  1'd1,  5'd9, 27'h000001fe, 5'd29, 27'h000000da, 5'd2, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000012d, 5'd27, 27'h0000000d, 5'd15, 27'h00000135, 32'h00000400,
  1'd1,  5'd8, 27'h00000348, 5'd26, 27'h000003d6, 5'd21, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000036c, 5'd7, 27'h00000376, 5'd2, 27'h0000007c, 32'h00000400,
  1'd1,  5'd20, 27'h00000079, 5'd10, 27'h0000005e, 5'd12, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003fe, 5'd9, 27'h000002b6, 5'd22, 27'h000001c3, 32'h00000400,
  1'd1,  5'd16, 27'h00000306, 5'd16, 27'h00000200, 5'd0, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d6, 5'd16, 27'h000001c8, 5'd14, 27'h000002ff, 32'h00000400,
  1'd1,  5'd18, 27'h00000048, 5'd17, 27'h0000019f, 5'd20, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000a6, 5'd27, 27'h00000050, 5'd1, 27'h000000f8, 32'h00000400,
  1'd1,  5'd18, 27'h000000af, 5'd28, 27'h0000028c, 5'd11, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016e, 5'd27, 27'h00000089, 5'd23, 27'h0000032e, 32'h00000400,
  1'd1,  5'd29, 27'h00000304, 5'd7, 27'h00000056, 5'd4, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b5, 5'd7, 27'h00000072, 5'd12, 27'h000000be, 32'h00000400,
  1'd1,  5'd30, 27'h00000044, 5'd5, 27'h000000fe, 5'd25, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000009, 5'd19, 27'h00000324, 5'd0, 27'h00000385, 32'h00000400,
  1'd1,  5'd29, 27'h0000024c, 5'd20, 27'h00000247, 5'd10, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000008c, 5'd19, 27'h00000117, 5'd23, 27'h000001c4, 32'h00000400,
  1'd1,  5'd29, 27'h00000229, 5'd28, 27'h00000191, 5'd0, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000020c, 5'd30, 27'h0000038b, 5'd10, 27'h00000259, 32'h00000400,
  1'd1,  5'd26, 27'h000003c6, 5'd26, 27'h000002fc, 5'd21, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000010a, 5'd6, 27'h0000011a, 5'd9, 27'h0000008f, 32'h00000400,
  1'd1,  5'd8, 27'h00000134, 5'd8, 27'h000002d6, 5'd18, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c2, 5'd7, 27'h000000d9, 5'd29, 27'h000003c0, 32'h00000400,
  1'd1,  5'd8, 27'h000001fd, 5'd18, 27'h000003fc, 5'd7, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001f7, 5'd18, 27'h00000073, 5'd18, 27'h00000217, 32'h00000400,
  1'd1,  5'd6, 27'h0000028c, 5'd19, 27'h000003f2, 5'd29, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a0, 5'd27, 27'h00000097, 5'd5, 27'h00000351, 32'h00000400,
  1'd1,  5'd7, 27'h000000c5, 5'd30, 27'h000001ce, 5'd17, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e8, 5'd27, 27'h000003d4, 5'd30, 27'h0000006e, 32'h00000400,
  1'd1,  5'd18, 27'h00000018, 5'd9, 27'h00000209, 5'd9, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002b1, 5'd5, 27'h00000126, 5'd15, 27'h00000376, 32'h00000400,
  1'd1,  5'd17, 27'h00000022, 5'd8, 27'h00000280, 5'd25, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000061, 5'd17, 27'h00000363, 5'd6, 27'h000003d8, 32'h00000400,
  1'd1,  5'd19, 27'h000000f0, 5'd17, 27'h0000030e, 5'd19, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000177, 5'd16, 27'h00000010, 5'd30, 27'h00000006, 32'h00000400,
  1'd1,  5'd19, 27'h00000138, 5'd30, 27'h00000207, 5'd5, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000026d, 5'd27, 27'h000001ba, 5'd18, 27'h000000b1, 32'h00000400,
  1'd1,  5'd19, 27'h00000258, 5'd29, 27'h000001cb, 5'd28, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000365, 5'd8, 27'h000000d2, 5'd6, 27'h00000011, 32'h00000400,
  1'd1,  5'd27, 27'h00000076, 5'd8, 27'h0000027f, 5'd18, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003ef, 5'd8, 27'h000001e6, 5'd26, 27'h000000b4, 32'h00000400,
  1'd1,  5'd27, 27'h00000196, 5'd18, 27'h0000009c, 5'd8, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000038f, 5'd18, 27'h000000a5, 5'd19, 27'h00000361, 32'h00000400,
  1'd1,  5'd29, 27'h00000224, 5'd16, 27'h000002c1, 5'd29, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000287, 5'd25, 27'h000003e6, 5'd6, 27'h000002a2, 32'h00000400,
  1'd1,  5'd27, 27'h0000032c, 5'd30, 27'h00000147, 5'd16, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000a8, 5'd27, 27'h000002a0, 5'd29, 27'h000003ae, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000201, 5'd0, 27'h0000035b, 5'd2, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000af, 5'd0, 27'h000000bb, 5'd14, 27'h000003e9, 32'h00000400,
  1'd1,  5'd2, 27'h00000276, 5'd0, 27'h0000019d, 5'd24, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000325, 5'd15, 27'h00000119, 5'd4, 27'h00000298, 32'h00000400,
  1'd1,  5'd0, 27'h00000063, 5'd10, 27'h00000334, 5'd12, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000323, 5'd13, 27'h000002b9, 5'd22, 27'h0000021b, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd25, 27'h000000b4, 5'd0, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000018d, 5'd24, 27'h00000102, 5'd10, 27'h0000039e, 32'h00000400,
  1'd1,  5'd0, 27'h00000321, 5'd24, 27'h000001b0, 5'd25, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002cc, 5'd1, 27'h000000bf, 5'd2, 27'h00000324, 32'h00000400,
  1'd1,  5'd14, 27'h000001bf, 5'd3, 27'h00000157, 5'd12, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001e0, 5'd3, 27'h00000140, 5'd21, 27'h0000010f, 32'h00000400,
  1'd1,  5'd10, 27'h000003a0, 5'd12, 27'h0000011a, 5'd1, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000142, 5'd13, 27'h0000029d, 5'd14, 27'h000002a6, 32'h00000400,
  1'd1,  5'd15, 27'h000001bc, 5'd12, 27'h00000140, 5'd24, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000396, 5'd24, 27'h0000018e, 5'd0, 27'h00000394, 32'h00000400,
  1'd1,  5'd11, 27'h00000084, 5'd24, 27'h00000299, 5'd11, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000030b, 5'd24, 27'h000002c8, 5'd20, 27'h000003f4, 32'h00000400,
  1'd1,  5'd21, 27'h000001ac, 5'd3, 27'h000003a0, 5'd1, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002d1, 5'd4, 27'h0000019f, 5'd14, 27'h00000001, 32'h00000400,
  1'd1,  5'd23, 27'h000003a1, 5'd3, 27'h00000082, 5'd24, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000030, 5'd11, 27'h00000067, 5'd4, 27'h00000331, 32'h00000400,
  1'd1,  5'd23, 27'h000001e3, 5'd12, 27'h00000204, 5'd15, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002f5, 5'd12, 27'h00000027, 5'd22, 27'h0000034e, 32'h00000400,
  1'd1,  5'd20, 27'h00000366, 5'd24, 27'h00000352, 5'd3, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000276, 5'd22, 27'h0000004a, 5'd14, 27'h000001fd, 32'h00000400,
  1'd1,  5'd21, 27'h0000005b, 5'd20, 27'h000003a6, 5'd22, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001c0, 5'd2, 27'h000000d6, 5'd10, 27'h000000f7, 32'h00000400,
  1'd1,  5'd1, 27'h000002af, 5'd2, 27'h0000005a, 5'd17, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b9, 5'd0, 27'h00000174, 5'd29, 27'h000001b3, 32'h00000400,
  1'd1,  5'd4, 27'h000003b8, 5'd11, 27'h0000033e, 5'd8, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000001, 5'd15, 27'h000000aa, 5'd18, 27'h0000015d, 32'h00000400,
  1'd1,  5'd2, 27'h000001e6, 5'd10, 27'h00000273, 5'd29, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000367, 5'd23, 27'h00000394, 5'd5, 27'h000000e1, 32'h00000400,
  1'd1,  5'd3, 27'h000001b4, 5'd23, 27'h00000359, 5'd20, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000035, 5'd25, 27'h00000230, 5'd26, 27'h00000355, 32'h00000400,
  1'd1,  5'd13, 27'h00000356, 5'd2, 27'h000002f5, 5'd5, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000340, 5'd3, 27'h0000030b, 5'd19, 27'h00000169, 32'h00000400,
  1'd1,  5'd12, 27'h0000020b, 5'd0, 27'h00000218, 5'd29, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ff, 5'd10, 27'h0000026d, 5'd5, 27'h0000011f, 32'h00000400,
  1'd1,  5'd10, 27'h0000021d, 5'd13, 27'h00000266, 5'd19, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b0, 5'd13, 27'h000000d3, 5'd29, 27'h0000007c, 32'h00000400,
  1'd1,  5'd14, 27'h00000054, 5'd23, 27'h000003fc, 5'd5, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000199, 5'd21, 27'h000003cc, 5'd20, 27'h00000012, 32'h00000400,
  1'd1,  5'd10, 27'h0000036e, 5'd24, 27'h000002e7, 5'd26, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002fe, 5'd3, 27'h000003d3, 5'd7, 27'h00000052, 32'h00000400,
  1'd1,  5'd24, 27'h0000034b, 5'd1, 27'h0000014e, 5'd18, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000039, 5'd4, 27'h00000345, 5'd28, 27'h000003e7, 32'h00000400,
  1'd1,  5'd21, 27'h0000021b, 5'd13, 27'h00000124, 5'd8, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000302, 5'd14, 27'h000002be, 5'd18, 27'h000001bb, 32'h00000400,
  1'd1,  5'd22, 27'h000002b9, 5'd11, 27'h00000262, 5'd27, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a0, 5'd23, 27'h00000152, 5'd5, 27'h00000295, 32'h00000400,
  1'd1,  5'd21, 27'h000000f6, 5'd22, 27'h00000031, 5'd16, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003cd, 5'd21, 27'h000001a1, 5'd30, 27'h00000300, 32'h00000400,
  1'd1,  5'd1, 27'h000000cb, 5'd7, 27'h000000af, 5'd1, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000089, 5'd8, 27'h0000024f, 5'd10, 27'h000001c9, 32'h00000400,
  1'd1,  5'd0, 27'h00000271, 5'd8, 27'h00000277, 5'd22, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002be, 5'd18, 27'h000001b4, 5'd2, 27'h00000222, 32'h00000400,
  1'd1,  5'd1, 27'h00000329, 5'd19, 27'h00000195, 5'd10, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000028e, 5'd18, 27'h000001c9, 5'd25, 27'h000002e2, 32'h00000400,
  1'd1,  5'd2, 27'h00000233, 5'd27, 27'h00000222, 5'd5, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000140, 5'd29, 27'h00000192, 5'd12, 27'h000002e3, 32'h00000400,
  1'd1,  5'd0, 27'h000002cb, 5'd27, 27'h000003d4, 5'd25, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000240, 5'd6, 27'h0000027b, 5'd3, 27'h0000025d, 32'h00000400,
  1'd1,  5'd13, 27'h00000288, 5'd6, 27'h00000078, 5'd11, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000b2, 5'd6, 27'h00000265, 5'd21, 27'h00000174, 32'h00000400,
  1'd1,  5'd11, 27'h0000003a, 5'd17, 27'h0000037a, 5'd2, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000377, 5'd18, 27'h00000382, 5'd12, 27'h0000021c, 32'h00000400,
  1'd1,  5'd11, 27'h00000026, 5'd16, 27'h00000027, 5'd24, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000092, 5'd30, 27'h00000368, 5'd0, 27'h000002ab, 32'h00000400,
  1'd1,  5'd14, 27'h00000360, 5'd26, 27'h000003df, 5'd11, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000247, 5'd27, 27'h0000010c, 5'd21, 27'h00000227, 32'h00000400,
  1'd1,  5'd25, 27'h00000200, 5'd9, 27'h0000014a, 5'd1, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000024e, 5'd7, 27'h000002b8, 5'd13, 27'h000003cd, 32'h00000400,
  1'd1,  5'd22, 27'h0000032b, 5'd6, 27'h0000010c, 5'd24, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000207, 5'd18, 27'h0000035c, 5'd0, 27'h000003ef, 32'h00000400,
  1'd1,  5'd23, 27'h000000cb, 5'd17, 27'h000001c1, 5'd11, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000190, 5'd17, 27'h0000021d, 5'd22, 27'h000000d2, 32'h00000400,
  1'd1,  5'd25, 27'h00000167, 5'd27, 27'h00000238, 5'd1, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e2, 5'd29, 27'h00000203, 5'd11, 27'h0000028e, 32'h00000400,
  1'd1,  5'd24, 27'h000003f1, 5'd28, 27'h00000186, 5'd24, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002c3, 5'd6, 27'h000003f2, 5'd7, 27'h000002a0, 32'h00000400,
  1'd1,  5'd3, 27'h00000319, 5'd7, 27'h00000368, 5'd17, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000212, 5'd5, 27'h0000030d, 5'd29, 27'h00000032, 32'h00000400,
  1'd1,  5'd3, 27'h0000002c, 5'd17, 27'h0000013b, 5'd7, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000284, 5'd17, 27'h000001e7, 5'd20, 27'h00000083, 32'h00000400,
  1'd1,  5'd2, 27'h000000ce, 5'd18, 27'h00000269, 5'd28, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000043, 5'd27, 27'h00000337, 5'd6, 27'h0000010b, 32'h00000400,
  1'd1,  5'd4, 27'h000000f2, 5'd30, 27'h000001ab, 5'd19, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000202, 5'd28, 27'h00000273, 5'd27, 27'h000003fd, 32'h00000400,
  1'd1,  5'd11, 27'h0000015b, 5'd5, 27'h00000180, 5'd9, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001c5, 5'd5, 27'h00000267, 5'd16, 27'h0000029d, 32'h00000400,
  1'd1,  5'd14, 27'h00000235, 5'd9, 27'h00000275, 5'd30, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003bc, 5'd15, 27'h000002ae, 5'd8, 27'h000003aa, 32'h00000400,
  1'd1,  5'd12, 27'h00000077, 5'd17, 27'h00000102, 5'd18, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029a, 5'd17, 27'h00000105, 5'd30, 27'h00000047, 32'h00000400,
  1'd1,  5'd13, 27'h0000008f, 5'd28, 27'h00000075, 5'd8, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000081, 5'd27, 27'h00000125, 5'd15, 27'h00000262, 32'h00000400,
  1'd1,  5'd10, 27'h000002f9, 5'd28, 27'h000003b2, 5'd26, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000ec, 5'd7, 27'h00000312, 5'd8, 27'h00000128, 32'h00000400,
  1'd1,  5'd20, 27'h000002ec, 5'd7, 27'h000002e1, 5'd16, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ba, 5'd9, 27'h000000c1, 5'd28, 27'h00000081, 32'h00000400,
  1'd1,  5'd22, 27'h00000167, 5'd18, 27'h000001e5, 5'd7, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000032a, 5'd17, 27'h000003e4, 5'd19, 27'h0000038b, 32'h00000400,
  1'd1,  5'd20, 27'h00000396, 5'd17, 27'h00000349, 5'd28, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000bd, 5'd30, 27'h000000a9, 5'd5, 27'h000003a9, 32'h00000400,
  1'd1,  5'd22, 27'h00000338, 5'd30, 27'h000000ad, 5'd19, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000002c, 5'd26, 27'h000001ec, 5'd30, 27'h000003a1, 32'h00000400,
  1'd1,  5'd5, 27'h000000cd, 5'd1, 27'h0000004d, 5'd9, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000221, 5'd0, 27'h000000bc, 5'd16, 27'h00000122, 32'h00000400,
  1'd1,  5'd6, 27'h00000013, 5'd1, 27'h000000a4, 5'd30, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000047, 5'd14, 27'h000000fd, 5'd3, 27'h000000bb, 32'h00000400,
  1'd1,  5'd5, 27'h00000348, 5'd12, 27'h000000d6, 5'd12, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000022c, 5'd14, 27'h000001c1, 5'd23, 27'h00000167, 32'h00000400,
  1'd1,  5'd5, 27'h000000f0, 5'd22, 27'h000003a3, 5'd3, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000f1, 5'd21, 27'h000003d6, 5'd11, 27'h00000174, 32'h00000400,
  1'd1,  5'd10, 27'h00000050, 5'd25, 27'h0000028e, 5'd20, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000003b, 5'd2, 27'h000000df, 5'd7, 27'h0000023b, 32'h00000400,
  1'd1,  5'd19, 27'h000003d3, 5'd1, 27'h000002e5, 5'd20, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000137, 5'd4, 27'h000000e2, 5'd29, 27'h0000006f, 32'h00000400,
  1'd1,  5'd17, 27'h0000013b, 5'd12, 27'h00000255, 5'd4, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e3, 5'd14, 27'h000000c3, 5'd13, 27'h00000286, 32'h00000400,
  1'd1,  5'd17, 27'h0000019c, 5'd11, 27'h00000382, 5'd24, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e5, 5'd25, 27'h00000124, 5'd0, 27'h00000116, 32'h00000400,
  1'd1,  5'd15, 27'h00000278, 5'd25, 27'h000001aa, 5'd14, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000004f, 5'd21, 27'h0000030f, 5'd25, 27'h000001fc, 32'h00000400,
  1'd1,  5'd27, 27'h00000196, 5'd4, 27'h0000029a, 5'd0, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000384, 5'd1, 27'h0000034a, 5'd15, 27'h000000fc, 32'h00000400,
  1'd1,  5'd27, 27'h00000279, 5'd1, 27'h0000021d, 5'd25, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001bf, 5'd13, 27'h00000128, 5'd1, 27'h000001f2, 32'h00000400,
  1'd1,  5'd29, 27'h00000267, 5'd10, 27'h000001ca, 5'd11, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000055, 5'd14, 27'h00000224, 5'd24, 27'h0000005f, 32'h00000400,
  1'd1,  5'd27, 27'h000000eb, 5'd21, 27'h0000023b, 5'd3, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000169, 5'd21, 27'h00000026, 5'd11, 27'h0000036c, 32'h00000400,
  1'd1,  5'd26, 27'h000003f5, 5'd24, 27'h000003f6, 5'd20, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c3, 5'd4, 27'h00000236, 5'd1, 27'h0000035d, 32'h00000400,
  1'd1,  5'd6, 27'h000003a4, 5'd0, 27'h00000307, 5'd15, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000377, 5'd1, 27'h0000005d, 5'd24, 27'h00000167, 32'h00000400,
  1'd1,  5'd9, 27'h000001b7, 5'd12, 27'h0000035a, 5'd5, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ee, 5'd15, 27'h000000ed, 5'd16, 27'h000002ad, 32'h00000400,
  1'd1,  5'd9, 27'h000000ca, 5'd12, 27'h00000103, 5'd28, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d8, 5'd22, 27'h00000331, 5'd9, 27'h0000019c, 32'h00000400,
  1'd1,  5'd9, 27'h000001ed, 5'd23, 27'h00000308, 5'd19, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e5, 5'd21, 27'h00000154, 5'd29, 27'h000003d0, 32'h00000400,
  1'd1,  5'd15, 27'h00000342, 5'd1, 27'h00000221, 5'd4, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000012d, 5'd5, 27'h00000021, 5'd13, 27'h000003f9, 32'h00000400,
  1'd1,  5'd19, 27'h00000212, 5'd3, 27'h00000302, 5'd24, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d0, 5'd13, 27'h000001df, 5'd9, 27'h0000031f, 32'h00000400,
  1'd1,  5'd15, 27'h000002f0, 5'd10, 27'h000003be, 5'd17, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003bb, 5'd12, 27'h000001a9, 5'd28, 27'h0000012e, 32'h00000400,
  1'd1,  5'd16, 27'h00000310, 5'd24, 27'h000000ed, 5'd10, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001fe, 5'd23, 27'h0000022d, 5'd19, 27'h0000000b, 32'h00000400,
  1'd1,  5'd16, 27'h000002c9, 5'd24, 27'h0000016f, 5'd26, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b9, 5'd4, 27'h00000385, 5'd7, 27'h00000328, 32'h00000400,
  1'd1,  5'd29, 27'h000002b8, 5'd4, 27'h0000024a, 5'd16, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000094, 5'd2, 27'h00000024, 5'd27, 27'h00000207, 32'h00000400,
  1'd1,  5'd27, 27'h0000011b, 5'd11, 27'h000001b0, 5'd8, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000312, 5'd13, 27'h0000021c, 5'd16, 27'h000003f2, 32'h00000400,
  1'd1,  5'd27, 27'h00000124, 5'd11, 27'h000003c1, 5'd26, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ae, 5'd22, 27'h000002ad, 5'd6, 27'h000000b5, 32'h00000400,
  1'd1,  5'd30, 27'h000003c0, 5'd24, 27'h0000014e, 5'd18, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000013d, 5'd25, 27'h00000316, 5'd27, 27'h00000024, 32'h00000400,
  1'd1,  5'd9, 27'h000000b5, 5'd7, 27'h000001b6, 5'd2, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034e, 5'd9, 27'h00000202, 5'd15, 27'h00000104, 32'h00000400,
  1'd1,  5'd5, 27'h0000021b, 5'd9, 27'h00000363, 5'd24, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000351, 5'd19, 27'h00000244, 5'd0, 27'h000000d0, 32'h00000400,
  1'd1,  5'd6, 27'h00000203, 5'd16, 27'h000003fc, 5'd13, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000015e, 5'd19, 27'h0000029b, 5'd22, 27'h000002b3, 32'h00000400,
  1'd1,  5'd5, 27'h00000314, 5'd28, 27'h0000012f, 5'd4, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011a, 5'd26, 27'h0000035a, 5'd14, 27'h000002dd, 32'h00000400,
  1'd1,  5'd8, 27'h00000256, 5'd26, 27'h000001ee, 5'd24, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000130, 5'd6, 27'h000001e0, 5'd0, 27'h0000029e, 32'h00000400,
  1'd1,  5'd18, 27'h00000188, 5'd8, 27'h00000015, 5'd12, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001b0, 5'd8, 27'h000002ba, 5'd21, 27'h000003e1, 32'h00000400,
  1'd1,  5'd19, 27'h000001cc, 5'd19, 27'h00000379, 5'd0, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000298, 5'd19, 27'h0000009c, 5'd11, 27'h0000012b, 32'h00000400,
  1'd1,  5'd19, 27'h0000022c, 5'd15, 27'h0000026f, 5'd21, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000028c, 5'd29, 27'h0000018e, 5'd0, 27'h00000300, 32'h00000400,
  1'd1,  5'd16, 27'h00000006, 5'd27, 27'h000003b3, 5'd12, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000272, 5'd28, 27'h000002eb, 5'd22, 27'h00000191, 32'h00000400,
  1'd1,  5'd29, 27'h00000172, 5'd5, 27'h000002b6, 5'd3, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e1, 5'd9, 27'h00000243, 5'd13, 27'h0000018f, 32'h00000400,
  1'd1,  5'd28, 27'h000001cb, 5'd6, 27'h000000c8, 5'd25, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000026b, 5'd16, 27'h000001a9, 5'd4, 27'h000003a6, 32'h00000400,
  1'd1,  5'd27, 27'h000002eb, 5'd20, 27'h0000005b, 5'd13, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003fc, 5'd17, 27'h000003e6, 5'd23, 27'h000000a5, 32'h00000400,
  1'd1,  5'd29, 27'h0000003f, 5'd27, 27'h00000130, 5'd3, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001c8, 5'd30, 27'h00000376, 5'd15, 27'h00000162, 32'h00000400,
  1'd1,  5'd28, 27'h00000230, 5'd28, 27'h00000374, 5'd23, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000001a, 5'd6, 27'h000001cd, 5'd9, 27'h0000028f, 32'h00000400,
  1'd1,  5'd5, 27'h00000100, 5'd6, 27'h000003bc, 5'd19, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000014b, 5'd10, 27'h00000015, 5'd27, 27'h000003a2, 32'h00000400,
  1'd1,  5'd9, 27'h0000020b, 5'd20, 27'h000002a0, 5'd6, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002e9, 5'd17, 27'h000000f8, 5'd15, 27'h0000034e, 32'h00000400,
  1'd1,  5'd6, 27'h00000066, 5'd15, 27'h000003a1, 5'd30, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d3, 5'd26, 27'h000002f5, 5'd8, 27'h00000382, 32'h00000400,
  1'd1,  5'd6, 27'h00000390, 5'd30, 27'h00000084, 5'd16, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ae, 5'd29, 27'h00000054, 5'd28, 27'h0000036b, 32'h00000400,
  1'd1,  5'd20, 27'h000002a9, 5'd7, 27'h000003bf, 5'd6, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000292, 5'd6, 27'h00000374, 5'd18, 27'h000000d7, 32'h00000400,
  1'd1,  5'd18, 27'h00000181, 5'd7, 27'h000002b0, 5'd26, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000005a, 5'd19, 27'h00000234, 5'd6, 27'h00000309, 32'h00000400,
  1'd1,  5'd18, 27'h000003d1, 5'd15, 27'h00000242, 5'd19, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002e3, 5'd17, 27'h000000f9, 5'd28, 27'h00000016, 32'h00000400,
  1'd1,  5'd19, 27'h000001b0, 5'd28, 27'h000000b9, 5'd5, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000026a, 5'd29, 27'h0000012f, 5'd18, 27'h000001f4, 32'h00000400,
  1'd1,  5'd16, 27'h00000103, 5'd29, 27'h00000025, 5'd29, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019c, 5'd7, 27'h00000065, 5'd8, 27'h000001ad, 32'h00000400,
  1'd1,  5'd27, 27'h00000355, 5'd8, 27'h00000309, 5'd19, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002cb, 5'd6, 27'h000000f6, 5'd28, 27'h0000019b, 32'h00000400,
  1'd1,  5'd27, 27'h000003ae, 5'd18, 27'h00000229, 5'd7, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000005, 5'd18, 27'h000000e3, 5'd20, 27'h00000157, 32'h00000400,
  1'd1,  5'd30, 27'h0000013d, 5'd15, 27'h00000232, 5'd29, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000362, 5'd29, 27'h00000029, 5'd6, 27'h000001a8, 32'h00000400,
  1'd1,  5'd27, 27'h0000005d, 5'd28, 27'h000001a5, 5'd16, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002bd, 5'd30, 27'h000000c5, 5'd29, 27'h00000048, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000109, 5'd0, 27'h000001b2, 5'd4, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000157, 5'd2, 27'h0000021b, 5'd14, 27'h0000009c, 32'h00000400,
  1'd1,  5'd4, 27'h0000027d, 5'd0, 27'h000003b2, 5'd23, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000338, 5'd12, 27'h0000002f, 5'd3, 27'h000000c6, 32'h00000400,
  1'd1,  5'd2, 27'h00000300, 5'd13, 27'h0000016b, 5'd10, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002dd, 5'd12, 27'h00000014, 5'd22, 27'h000003a1, 32'h00000400,
  1'd1,  5'd1, 27'h000000b5, 5'd21, 27'h000003d2, 5'd4, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000136, 5'd22, 27'h000002c9, 5'd10, 27'h00000386, 32'h00000400,
  1'd1,  5'd3, 27'h00000125, 5'd25, 27'h00000276, 5'd21, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035a, 5'd1, 27'h00000173, 5'd1, 27'h00000249, 32'h00000400,
  1'd1,  5'd10, 27'h0000015d, 5'd0, 27'h000001a1, 5'd13, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000001c, 5'd2, 27'h00000368, 5'd24, 27'h00000232, 32'h00000400,
  1'd1,  5'd14, 27'h0000031c, 5'd13, 27'h0000030a, 5'd1, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000272, 5'd12, 27'h00000270, 5'd10, 27'h000002c7, 32'h00000400,
  1'd1,  5'd14, 27'h00000390, 5'd12, 27'h000002b3, 5'd25, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000001a, 5'd23, 27'h000000b1, 5'd1, 27'h0000008d, 32'h00000400,
  1'd1,  5'd11, 27'h0000034e, 5'd23, 27'h00000267, 5'd10, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038f, 5'd24, 27'h000002bb, 5'd25, 27'h000002b4, 32'h00000400,
  1'd1,  5'd22, 27'h0000014c, 5'd1, 27'h0000031b, 5'd0, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000030a, 5'd2, 27'h00000307, 5'd11, 27'h000002ec, 32'h00000400,
  1'd1,  5'd25, 27'h000002f4, 5'd0, 27'h00000174, 5'd22, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b3, 5'd11, 27'h00000113, 5'd2, 27'h000000d6, 32'h00000400,
  1'd1,  5'd22, 27'h000000a2, 5'd13, 27'h000000bb, 5'd11, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b1, 5'd13, 27'h00000195, 5'd24, 27'h0000015c, 32'h00000400,
  1'd1,  5'd22, 27'h000001e9, 5'd23, 27'h0000015f, 5'd3, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000a8, 5'd24, 27'h000002ad, 5'd14, 27'h0000000e, 32'h00000400,
  1'd1,  5'd22, 27'h000001a6, 5'd22, 27'h00000336, 5'd25, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000010c, 5'd3, 27'h0000011d, 5'd8, 27'h000001b6, 32'h00000400,
  1'd1,  5'd3, 27'h0000034c, 5'd1, 27'h000000bf, 5'd20, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000138, 5'd2, 27'h00000352, 5'd27, 27'h00000294, 32'h00000400,
  1'd1,  5'd0, 27'h00000168, 5'd12, 27'h00000227, 5'd9, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000208, 5'd11, 27'h00000120, 5'd19, 27'h00000237, 32'h00000400,
  1'd1,  5'd2, 27'h00000294, 5'd10, 27'h000001e9, 5'd27, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000c9, 5'd20, 27'h000003ce, 5'd9, 27'h00000079, 32'h00000400,
  1'd1,  5'd0, 27'h00000355, 5'd24, 27'h000003c6, 5'd18, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000003e, 5'd23, 27'h000000bb, 5'd30, 27'h00000013, 32'h00000400,
  1'd1,  5'd11, 27'h000002d8, 5'd2, 27'h000000e1, 5'd5, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000037d, 5'd4, 27'h00000103, 5'd19, 27'h00000146, 32'h00000400,
  1'd1,  5'd12, 27'h000001a8, 5'd2, 27'h00000212, 5'd30, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000012b, 5'd15, 27'h00000195, 5'd8, 27'h000003b4, 32'h00000400,
  1'd1,  5'd11, 27'h00000340, 5'd14, 27'h00000340, 5'd16, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ae, 5'd14, 27'h000000eb, 5'd29, 27'h00000233, 32'h00000400,
  1'd1,  5'd10, 27'h000001a1, 5'd25, 27'h0000026b, 5'd8, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000030d, 5'd24, 27'h00000327, 5'd19, 27'h00000253, 32'h00000400,
  1'd1,  5'd14, 27'h00000121, 5'd24, 27'h00000235, 5'd26, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b6, 5'd1, 27'h00000076, 5'd8, 27'h000000ac, 32'h00000400,
  1'd1,  5'd25, 27'h000002ef, 5'd1, 27'h000003a6, 5'd15, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000041, 5'd4, 27'h000000a3, 5'd25, 27'h000003f2, 32'h00000400,
  1'd1,  5'd21, 27'h00000353, 5'd15, 27'h00000183, 5'd7, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000081, 5'd14, 27'h00000038, 5'd18, 27'h000001c1, 32'h00000400,
  1'd1,  5'd23, 27'h0000018d, 5'd13, 27'h0000037c, 5'd28, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000108, 5'd25, 27'h00000070, 5'd10, 27'h00000055, 32'h00000400,
  1'd1,  5'd22, 27'h000000f7, 5'd24, 27'h000003ae, 5'd16, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000031e, 5'd21, 27'h000001db, 5'd30, 27'h00000241, 32'h00000400,
  1'd1,  5'd2, 27'h000002fc, 5'd7, 27'h00000038, 5'd2, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000047, 5'd7, 27'h000001f2, 5'd10, 27'h000002a6, 32'h00000400,
  1'd1,  5'd4, 27'h0000037e, 5'd8, 27'h000001ca, 5'd23, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000f7, 5'd15, 27'h000002d3, 5'd3, 27'h00000319, 32'h00000400,
  1'd1,  5'd1, 27'h00000340, 5'd19, 27'h000002d7, 5'd14, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000144, 5'd16, 27'h00000076, 5'd24, 27'h00000098, 32'h00000400,
  1'd1,  5'd3, 27'h00000080, 5'd30, 27'h000003b5, 5'd5, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000216, 5'd28, 27'h00000322, 5'd15, 27'h000001f7, 32'h00000400,
  1'd1,  5'd2, 27'h000002c9, 5'd26, 27'h00000309, 5'd25, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000cd, 5'd7, 27'h00000057, 5'd0, 27'h000001ba, 32'h00000400,
  1'd1,  5'd15, 27'h000001cf, 5'd6, 27'h000000d3, 5'd10, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a5, 5'd9, 27'h00000314, 5'd23, 27'h00000183, 32'h00000400,
  1'd1,  5'd10, 27'h000003b3, 5'd17, 27'h00000003, 5'd3, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000320, 5'd16, 27'h00000282, 5'd14, 27'h000000a3, 32'h00000400,
  1'd1,  5'd13, 27'h000001fb, 5'd17, 27'h00000076, 5'd22, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001ed, 5'd28, 27'h000000e7, 5'd2, 27'h000002dd, 32'h00000400,
  1'd1,  5'd12, 27'h00000073, 5'd29, 27'h0000024c, 5'd15, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001b3, 5'd30, 27'h0000014d, 5'd25, 27'h000000bc, 32'h00000400,
  1'd1,  5'd22, 27'h000002ee, 5'd5, 27'h000002b9, 5'd1, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000287, 5'd5, 27'h0000036c, 5'd12, 27'h00000319, 32'h00000400,
  1'd1,  5'd22, 27'h00000295, 5'd6, 27'h000003c9, 5'd24, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002c0, 5'd18, 27'h00000159, 5'd2, 27'h00000117, 32'h00000400,
  1'd1,  5'd22, 27'h000001eb, 5'd15, 27'h0000033a, 5'd13, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000005d, 5'd18, 27'h00000053, 5'd21, 27'h00000170, 32'h00000400,
  1'd1,  5'd22, 27'h000002c3, 5'd28, 27'h00000030, 5'd2, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000212, 5'd29, 27'h00000069, 5'd14, 27'h0000023e, 32'h00000400,
  1'd1,  5'd25, 27'h00000096, 5'd29, 27'h00000354, 5'd21, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000037b, 5'd7, 27'h0000035c, 5'd6, 27'h00000303, 32'h00000400,
  1'd1,  5'd4, 27'h000000bc, 5'd5, 27'h0000020f, 5'd17, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000083, 5'd8, 27'h0000027e, 5'd27, 27'h00000181, 32'h00000400,
  1'd1,  5'd4, 27'h00000009, 5'd17, 27'h00000025, 5'd7, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002d0, 5'd18, 27'h000000bd, 5'd18, 27'h000003e6, 32'h00000400,
  1'd1,  5'd2, 27'h000000ae, 5'd18, 27'h00000314, 5'd28, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028c, 5'd28, 27'h000001be, 5'd9, 27'h00000054, 32'h00000400,
  1'd1,  5'd3, 27'h000001ea, 5'd27, 27'h0000021f, 5'd18, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a8, 5'd26, 27'h000003b5, 5'd27, 27'h0000034c, 32'h00000400,
  1'd1,  5'd12, 27'h000002e4, 5'd8, 27'h000002e5, 5'd8, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ee, 5'd8, 27'h000002f0, 5'd20, 27'h000000e1, 32'h00000400,
  1'd1,  5'd13, 27'h0000023b, 5'd7, 27'h000003f1, 5'd27, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000036c, 5'd16, 27'h0000024b, 5'd6, 27'h0000033c, 32'h00000400,
  1'd1,  5'd11, 27'h0000022e, 5'd16, 27'h000003fe, 5'd18, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f7, 5'd20, 27'h000000c5, 5'd26, 27'h00000023, 32'h00000400,
  1'd1,  5'd11, 27'h000001d2, 5'd27, 27'h0000007f, 5'd8, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d4, 5'd29, 27'h00000022, 5'd15, 27'h00000372, 32'h00000400,
  1'd1,  5'd11, 27'h000003f2, 5'd29, 27'h000002f3, 5'd27, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000021, 5'd8, 27'h000000aa, 5'd7, 27'h0000001b, 32'h00000400,
  1'd1,  5'd25, 27'h00000151, 5'd7, 27'h0000025c, 5'd17, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001f5, 5'd7, 27'h0000035d, 5'd27, 27'h000001f4, 32'h00000400,
  1'd1,  5'd21, 27'h000001a7, 5'd16, 27'h00000103, 5'd5, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000039d, 5'd18, 27'h0000008a, 5'd15, 27'h00000264, 32'h00000400,
  1'd1,  5'd23, 27'h00000306, 5'd20, 27'h000000bd, 5'd28, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000031f, 5'd28, 27'h000001dc, 5'd7, 27'h00000032, 32'h00000400,
  1'd1,  5'd22, 27'h000000b6, 5'd27, 27'h00000046, 5'd20, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ea, 5'd29, 27'h000001ad, 5'd30, 27'h00000377, 32'h00000400,
  1'd1,  5'd9, 27'h000002a7, 5'd5, 27'h00000099, 5'd6, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000375, 5'd4, 27'h000001ac, 5'd17, 27'h000003e6, 32'h00000400,
  1'd1,  5'd5, 27'h000003c8, 5'd3, 27'h000002e1, 5'd26, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ac, 5'd12, 27'h000000c5, 5'd1, 27'h00000306, 32'h00000400,
  1'd1,  5'd5, 27'h00000390, 5'd14, 27'h000003c0, 5'd11, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ef, 5'd12, 27'h000003b1, 5'd23, 27'h0000018a, 32'h00000400,
  1'd1,  5'd6, 27'h00000377, 5'd23, 27'h00000146, 5'd2, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003aa, 5'd25, 27'h000000a2, 5'd14, 27'h00000212, 32'h00000400,
  1'd1,  5'd10, 27'h0000004b, 5'd24, 27'h00000365, 5'd22, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000017, 5'd0, 27'h00000133, 5'd7, 27'h00000046, 32'h00000400,
  1'd1,  5'd17, 27'h00000232, 5'd1, 27'h00000197, 5'd19, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000217, 5'd2, 27'h0000009e, 5'd26, 27'h000002b7, 32'h00000400,
  1'd1,  5'd16, 27'h000002f8, 5'd12, 27'h00000102, 5'd1, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000146, 5'd15, 27'h00000073, 5'd12, 27'h00000383, 32'h00000400,
  1'd1,  5'd19, 27'h00000264, 5'd14, 27'h000003b2, 5'd23, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000046, 5'd23, 27'h0000029b, 5'd0, 27'h000000c7, 32'h00000400,
  1'd1,  5'd20, 27'h00000109, 5'd21, 27'h00000136, 5'd11, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000022, 5'd23, 27'h000000e1, 5'd20, 27'h0000035b, 32'h00000400,
  1'd1,  5'd28, 27'h00000241, 5'd2, 27'h00000140, 5'd1, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000130, 5'd0, 27'h000003d9, 5'd10, 27'h00000251, 32'h00000400,
  1'd1,  5'd29, 27'h0000028f, 5'd4, 27'h0000012c, 5'd23, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003d0, 5'd13, 27'h00000217, 5'd1, 27'h000002c2, 32'h00000400,
  1'd1,  5'd27, 27'h0000007d, 5'd13, 27'h0000025f, 5'd14, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c6, 5'd10, 27'h00000312, 5'd23, 27'h00000126, 32'h00000400,
  1'd1,  5'd26, 27'h00000361, 5'd22, 27'h000001aa, 5'd1, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000278, 5'd25, 27'h000001f7, 5'd11, 27'h00000175, 32'h00000400,
  1'd1,  5'd26, 27'h000000ac, 5'd22, 27'h000002a7, 5'd21, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000007, 5'd3, 27'h00000367, 5'd1, 27'h000002b4, 32'h00000400,
  1'd1,  5'd9, 27'h00000085, 5'd4, 27'h0000039f, 5'd14, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000045, 5'd4, 27'h000002ab, 5'd22, 27'h00000108, 32'h00000400,
  1'd1,  5'd5, 27'h00000123, 5'd12, 27'h00000094, 5'd9, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000200, 5'd11, 27'h000002ab, 5'd18, 27'h0000007f, 32'h00000400,
  1'd1,  5'd8, 27'h00000166, 5'd13, 27'h000000fa, 5'd30, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002a2, 5'd24, 27'h00000301, 5'd6, 27'h0000007c, 32'h00000400,
  1'd1,  5'd9, 27'h000003ed, 5'd22, 27'h000000c4, 5'd18, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f8, 5'd23, 27'h00000277, 5'd30, 27'h00000097, 32'h00000400,
  1'd1,  5'd17, 27'h00000380, 5'd3, 27'h00000054, 5'd0, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e6, 5'd2, 27'h0000022e, 5'd10, 27'h0000033a, 32'h00000400,
  1'd1,  5'd16, 27'h0000026c, 5'd3, 27'h0000031c, 5'd23, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000024f, 5'd13, 27'h00000378, 5'd6, 27'h00000209, 32'h00000400,
  1'd1,  5'd19, 27'h000000bc, 5'd10, 27'h00000384, 5'd16, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000153, 5'd13, 27'h00000107, 5'd26, 27'h00000036, 32'h00000400,
  1'd1,  5'd19, 27'h000003e4, 5'd21, 27'h00000072, 5'd9, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029b, 5'd22, 27'h00000007, 5'd20, 27'h00000153, 32'h00000400,
  1'd1,  5'd18, 27'h000003a8, 5'd20, 27'h000003ba, 5'd27, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000018a, 5'd2, 27'h00000081, 5'd6, 27'h000001ac, 32'h00000400,
  1'd1,  5'd26, 27'h00000041, 5'd0, 27'h0000031b, 5'd17, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003da, 5'd4, 27'h000003e2, 5'd28, 27'h00000364, 32'h00000400,
  1'd1,  5'd29, 27'h00000201, 5'd13, 27'h0000000a, 5'd8, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000038d, 5'd11, 27'h000002aa, 5'd15, 27'h0000034a, 32'h00000400,
  1'd1,  5'd29, 27'h0000023b, 5'd14, 27'h0000025f, 5'd28, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000012d, 5'd22, 27'h00000397, 5'd6, 27'h00000314, 32'h00000400,
  1'd1,  5'd30, 27'h000002ef, 5'd21, 27'h0000007d, 5'd18, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000bf, 5'd23, 27'h00000290, 5'd26, 27'h000001a9, 32'h00000400,
  1'd1,  5'd8, 27'h000003bc, 5'd5, 27'h0000017e, 5'd2, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a6, 5'd8, 27'h00000222, 5'd14, 27'h0000000b, 32'h00000400,
  1'd1,  5'd9, 27'h00000004, 5'd9, 27'h000000b7, 5'd23, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000248, 5'd17, 27'h00000211, 5'd3, 27'h000003ac, 32'h00000400,
  1'd1,  5'd10, 27'h00000076, 5'd18, 27'h00000374, 5'd11, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034e, 5'd18, 27'h000000b5, 5'd22, 27'h000002ea, 32'h00000400,
  1'd1,  5'd6, 27'h000001cd, 5'd29, 27'h00000200, 5'd3, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000343, 5'd27, 27'h000000d7, 5'd12, 27'h0000033f, 32'h00000400,
  1'd1,  5'd9, 27'h0000020d, 5'd27, 27'h000002da, 5'd22, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000017, 5'd7, 27'h0000038d, 5'd1, 27'h00000189, 32'h00000400,
  1'd1,  5'd16, 27'h000000f0, 5'd5, 27'h000000d8, 5'd11, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000068, 5'd5, 27'h000000b9, 5'd24, 27'h00000393, 32'h00000400,
  1'd1,  5'd17, 27'h00000199, 5'd16, 27'h000002d4, 5'd4, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000390, 5'd15, 27'h000003c1, 5'd13, 27'h000000de, 32'h00000400,
  1'd1,  5'd20, 27'h00000121, 5'd18, 27'h000001f4, 5'd22, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d6, 5'd28, 27'h0000013f, 5'd0, 27'h0000027a, 32'h00000400,
  1'd1,  5'd15, 27'h0000024f, 5'd26, 27'h00000331, 5'd15, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000347, 5'd27, 27'h0000027f, 5'd25, 27'h00000114, 32'h00000400,
  1'd1,  5'd26, 27'h000003fe, 5'd7, 27'h0000038f, 5'd3, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000008c, 5'd5, 27'h000001f6, 5'd11, 27'h0000007a, 32'h00000400,
  1'd1,  5'd30, 27'h000000a6, 5'd8, 27'h000000fc, 5'd21, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000035d, 5'd20, 27'h00000057, 5'd3, 27'h00000163, 32'h00000400,
  1'd1,  5'd27, 27'h00000246, 5'd18, 27'h000001e5, 5'd14, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000030a, 5'd18, 27'h0000026f, 5'd22, 27'h0000004d, 32'h00000400,
  1'd1,  5'd27, 27'h00000059, 5'd28, 27'h000000bf, 5'd3, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000f, 5'd26, 27'h000000f8, 5'd10, 27'h00000215, 32'h00000400,
  1'd1,  5'd30, 27'h0000023b, 5'd27, 27'h00000318, 5'd22, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000018a, 5'd10, 27'h00000150, 5'd8, 27'h000002b3, 32'h00000400,
  1'd1,  5'd5, 27'h000003cc, 5'd6, 27'h00000322, 5'd16, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000035b, 5'd6, 27'h000001d3, 5'd29, 27'h0000004e, 32'h00000400,
  1'd1,  5'd9, 27'h00000355, 5'd18, 27'h00000303, 5'd8, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000031d, 5'd16, 27'h000000d1, 5'd16, 27'h00000299, 32'h00000400,
  1'd1,  5'd7, 27'h0000022b, 5'd18, 27'h0000002b, 5'd27, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000364, 5'd30, 27'h000003c1, 5'd7, 27'h000001eb, 32'h00000400,
  1'd1,  5'd5, 27'h0000038c, 5'd29, 27'h000002f3, 5'd17, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032f, 5'd26, 27'h00000207, 5'd29, 27'h000003ba, 32'h00000400,
  1'd1,  5'd15, 27'h0000022f, 5'd9, 27'h00000218, 5'd6, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000234, 5'd6, 27'h00000153, 5'd19, 27'h0000024a, 32'h00000400,
  1'd1,  5'd16, 27'h00000176, 5'd10, 27'h000000f4, 5'd27, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002eb, 5'd18, 27'h00000332, 5'd7, 27'h00000365, 32'h00000400,
  1'd1,  5'd18, 27'h00000085, 5'd18, 27'h000001dd, 5'd20, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001a3, 5'd15, 27'h000002bb, 5'd27, 27'h000002b5, 32'h00000400,
  1'd1,  5'd20, 27'h00000252, 5'd30, 27'h00000041, 5'd7, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ee, 5'd27, 27'h000003fa, 5'd18, 27'h000002d6, 32'h00000400,
  1'd1,  5'd18, 27'h0000015b, 5'd28, 27'h000000ef, 5'd26, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003be, 5'd6, 27'h000003de, 5'd8, 27'h0000000c, 32'h00000400,
  1'd1,  5'd30, 27'h0000034a, 5'd6, 27'h000001ec, 5'd16, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000106, 5'd9, 27'h00000020, 5'd28, 27'h000003b5, 32'h00000400,
  1'd1,  5'd28, 27'h00000389, 5'd20, 27'h00000200, 5'd8, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000032c, 5'd19, 27'h000000b9, 5'd15, 27'h000002ec, 32'h00000400,
  1'd1,  5'd28, 27'h000001cb, 5'd18, 27'h000003e4, 5'd29, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000029d, 5'd28, 27'h00000006, 5'd8, 27'h00000153, 32'h00000400,
  1'd1,  5'd26, 27'h000000d8, 5'd27, 27'h000002ff, 5'd19, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000197, 5'd30, 27'h00000154, 5'd30, 27'h00000320, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000002ff, 5'd2, 27'h00000124, 5'd1, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000331, 5'd3, 27'h00000017, 5'd14, 27'h000001fe, 32'h00000400,
  1'd1,  5'd1, 27'h000000ba, 5'd0, 27'h00000001, 5'd22, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d0, 5'd11, 27'h000002ef, 5'd5, 27'h000000a4, 32'h00000400,
  1'd1,  5'd4, 27'h00000211, 5'd12, 27'h00000264, 5'd12, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ef, 5'd14, 27'h0000029f, 5'd23, 27'h000003cb, 32'h00000400,
  1'd1,  5'd4, 27'h000001ee, 5'd21, 27'h00000203, 5'd0, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003e3, 5'd21, 27'h000002c5, 5'd13, 27'h00000158, 32'h00000400,
  1'd1,  5'd0, 27'h000003e8, 5'd25, 27'h000000fb, 5'd22, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000217, 5'd1, 27'h00000080, 5'd3, 27'h000003dd, 32'h00000400,
  1'd1,  5'd12, 27'h000003af, 5'd3, 27'h000002ed, 5'd14, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000274, 5'd0, 27'h0000012e, 5'd20, 27'h000002b0, 32'h00000400,
  1'd1,  5'd11, 27'h00000272, 5'd14, 27'h00000139, 5'd2, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d9, 5'd12, 27'h0000015c, 5'd13, 27'h000001ed, 32'h00000400,
  1'd1,  5'd14, 27'h00000336, 5'd10, 27'h00000218, 5'd23, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035a, 5'd21, 27'h00000372, 5'd0, 27'h00000008, 32'h00000400,
  1'd1,  5'd13, 27'h00000244, 5'd23, 27'h0000012e, 5'd13, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000060, 5'd25, 27'h0000012a, 5'd25, 27'h0000000c, 32'h00000400,
  1'd1,  5'd20, 27'h00000346, 5'd2, 27'h00000115, 5'd3, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001a3, 5'd2, 27'h00000307, 5'd14, 27'h0000020c, 32'h00000400,
  1'd1,  5'd21, 27'h00000226, 5'd5, 27'h00000050, 5'd22, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000153, 5'd13, 27'h000000c3, 5'd0, 27'h0000034a, 32'h00000400,
  1'd1,  5'd22, 27'h000000e5, 5'd10, 27'h0000036e, 5'd11, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000001a, 5'd13, 27'h00000329, 5'd24, 27'h00000178, 32'h00000400,
  1'd1,  5'd22, 27'h0000004c, 5'd23, 27'h00000061, 5'd2, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000210, 5'd23, 27'h000002cd, 5'd14, 27'h00000316, 32'h00000400,
  1'd1,  5'd22, 27'h0000006c, 5'd25, 27'h000000a1, 5'd25, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002fe, 5'd3, 27'h0000001d, 5'd9, 27'h000001ad, 32'h00000400,
  1'd1,  5'd1, 27'h000002c4, 5'd1, 27'h000003d1, 5'd16, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d9, 5'd3, 27'h000002d3, 5'd26, 27'h0000018d, 32'h00000400,
  1'd1,  5'd1, 27'h0000021b, 5'd15, 27'h0000000c, 5'd6, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002b9, 5'd13, 27'h0000002a, 5'd17, 27'h0000006b, 32'h00000400,
  1'd1,  5'd3, 27'h0000002d, 5'd12, 27'h000003a5, 5'd29, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000008d, 5'd23, 27'h00000213, 5'd8, 27'h000002dc, 32'h00000400,
  1'd1,  5'd4, 27'h000003eb, 5'd24, 27'h00000166, 5'd16, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000393, 5'd21, 27'h000002de, 5'd29, 27'h00000020, 32'h00000400,
  1'd1,  5'd13, 27'h0000029a, 5'd5, 27'h000000aa, 5'd7, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000038f, 5'd1, 27'h0000005a, 5'd17, 27'h00000314, 32'h00000400,
  1'd1,  5'd11, 27'h00000214, 5'd1, 27'h0000005f, 5'd27, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000148, 5'd13, 27'h00000315, 5'd9, 27'h00000101, 32'h00000400,
  1'd1,  5'd11, 27'h00000278, 5'd15, 27'h00000140, 5'd17, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000006d, 5'd12, 27'h0000036c, 5'd26, 27'h000001ef, 32'h00000400,
  1'd1,  5'd11, 27'h00000364, 5'd24, 27'h0000014a, 5'd6, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000123, 5'd21, 27'h00000112, 5'd19, 27'h000002a3, 32'h00000400,
  1'd1,  5'd11, 27'h000003c3, 5'd25, 27'h0000015a, 5'd27, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000013a, 5'd1, 27'h000001b1, 5'd8, 27'h0000034c, 32'h00000400,
  1'd1,  5'd22, 27'h000003ec, 5'd2, 27'h00000151, 5'd16, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000392, 5'd5, 27'h00000061, 5'd30, 27'h000002fd, 32'h00000400,
  1'd1,  5'd25, 27'h00000088, 5'd12, 27'h00000165, 5'd7, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003c2, 5'd11, 27'h0000002e, 5'd19, 27'h000003b6, 32'h00000400,
  1'd1,  5'd22, 27'h000003a7, 5'd13, 27'h000003bb, 5'd27, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000200, 5'd25, 27'h000000da, 5'd7, 27'h00000202, 32'h00000400,
  1'd1,  5'd25, 27'h00000070, 5'd25, 27'h00000240, 5'd18, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000016e, 5'd25, 27'h0000017b, 5'd26, 27'h00000226, 32'h00000400,
  1'd1,  5'd1, 27'h00000306, 5'd8, 27'h00000320, 5'd2, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000008a, 5'd7, 27'h00000264, 5'd13, 27'h000000fa, 32'h00000400,
  1'd1,  5'd2, 27'h000001dd, 5'd8, 27'h00000037, 5'd21, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000191, 5'd16, 27'h00000258, 5'd0, 27'h000002e6, 32'h00000400,
  1'd1,  5'd3, 27'h00000261, 5'd16, 27'h000003eb, 5'd13, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000145, 5'd16, 27'h000000ba, 5'd25, 27'h00000172, 32'h00000400,
  1'd1,  5'd1, 27'h00000085, 5'd30, 27'h00000281, 5'd2, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000371, 5'd28, 27'h00000162, 5'd11, 27'h000000f4, 32'h00000400,
  1'd1,  5'd0, 27'h000002f1, 5'd30, 27'h0000035e, 5'd24, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001f0, 5'd8, 27'h0000025a, 5'd0, 27'h0000029b, 32'h00000400,
  1'd1,  5'd11, 27'h00000247, 5'd7, 27'h00000171, 5'd15, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000391, 5'd8, 27'h0000022b, 5'd25, 27'h000002e8, 32'h00000400,
  1'd1,  5'd14, 27'h00000386, 5'd20, 27'h0000018e, 5'd0, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000011, 5'd19, 27'h0000028d, 5'd11, 27'h000000db, 32'h00000400,
  1'd1,  5'd10, 27'h00000369, 5'd17, 27'h000001dc, 5'd22, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000320, 5'd29, 27'h000000ac, 5'd3, 27'h00000176, 32'h00000400,
  1'd1,  5'd10, 27'h000002ec, 5'd27, 27'h0000009a, 5'd14, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000345, 5'd30, 27'h000000a5, 5'd21, 27'h000002b1, 32'h00000400,
  1'd1,  5'd21, 27'h0000019e, 5'd8, 27'h00000338, 5'd0, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002a5, 5'd6, 27'h0000022f, 5'd10, 27'h000001f5, 32'h00000400,
  1'd1,  5'd22, 27'h0000035e, 5'd9, 27'h000002c3, 5'd23, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032e, 5'd18, 27'h000003d3, 5'd2, 27'h0000031d, 32'h00000400,
  1'd1,  5'd24, 27'h0000002c, 5'd19, 27'h00000162, 5'd15, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000011a, 5'd20, 27'h000000b3, 5'd22, 27'h0000032b, 32'h00000400,
  1'd1,  5'd23, 27'h000003d1, 5'd26, 27'h000001a2, 5'd4, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000081, 5'd28, 27'h000002fe, 5'd13, 27'h000001f4, 32'h00000400,
  1'd1,  5'd21, 27'h000003a3, 5'd29, 27'h00000301, 5'd23, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000c2, 5'd6, 27'h00000023, 5'd7, 27'h0000025f, 32'h00000400,
  1'd1,  5'd3, 27'h0000023b, 5'd6, 27'h000001ac, 5'd16, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003cc, 5'd10, 27'h000000b4, 5'd28, 27'h000002f9, 32'h00000400,
  1'd1,  5'd2, 27'h0000019e, 5'd15, 27'h0000027b, 5'd8, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c0, 5'd17, 27'h000002ad, 5'd16, 27'h00000400, 32'h00000400,
  1'd1,  5'd5, 27'h0000007c, 5'd18, 27'h0000028f, 5'd27, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000260, 5'd29, 27'h00000376, 5'd5, 27'h00000341, 32'h00000400,
  1'd1,  5'd1, 27'h00000108, 5'd25, 27'h000003a4, 5'd17, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000d8, 5'd30, 27'h000000cf, 5'd30, 27'h00000038, 32'h00000400,
  1'd1,  5'd13, 27'h00000084, 5'd5, 27'h00000341, 5'd7, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f2, 5'd6, 27'h00000000, 5'd15, 27'h000003b5, 32'h00000400,
  1'd1,  5'd12, 27'h0000030f, 5'd7, 27'h00000299, 5'd28, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000030a, 5'd16, 27'h000002c2, 5'd10, 27'h00000015, 32'h00000400,
  1'd1,  5'd11, 27'h0000031d, 5'd18, 27'h000002d0, 5'd19, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000203, 5'd16, 27'h000000d9, 5'd26, 27'h000002c3, 32'h00000400,
  1'd1,  5'd14, 27'h00000069, 5'd30, 27'h00000159, 5'd5, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000320, 5'd29, 27'h000002e7, 5'd18, 27'h0000029b, 32'h00000400,
  1'd1,  5'd12, 27'h00000162, 5'd30, 27'h0000038b, 5'd27, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000028d, 5'd5, 27'h00000298, 5'd10, 27'h0000005a, 32'h00000400,
  1'd1,  5'd24, 27'h000002e2, 5'd7, 27'h000000a1, 5'd15, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000070, 5'd10, 27'h000000e0, 5'd30, 27'h000002d1, 32'h00000400,
  1'd1,  5'd21, 27'h00000213, 5'd16, 27'h000000f6, 5'd8, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003bb, 5'd16, 27'h0000021c, 5'd15, 27'h000003a4, 32'h00000400,
  1'd1,  5'd23, 27'h000002a0, 5'd16, 27'h0000021a, 5'd27, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000340, 5'd28, 27'h000000d5, 5'd9, 27'h0000004e, 32'h00000400,
  1'd1,  5'd22, 27'h0000026d, 5'd29, 27'h00000294, 5'd16, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001ad, 5'd29, 27'h000001c3, 5'd29, 27'h000003ac, 32'h00000400,
  1'd1,  5'd10, 27'h0000001b, 5'd1, 27'h000001df, 5'd5, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000153, 5'd0, 27'h00000024, 5'd19, 27'h0000011b, 32'h00000400,
  1'd1,  5'd9, 27'h0000019f, 5'd1, 27'h00000087, 5'd27, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000309, 5'd10, 27'h00000375, 5'd1, 27'h00000109, 32'h00000400,
  1'd1,  5'd9, 27'h000003e7, 5'd12, 27'h00000190, 5'd10, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000269, 5'd10, 27'h000001f2, 5'd20, 27'h00000367, 32'h00000400,
  1'd1,  5'd8, 27'h000003ed, 5'd21, 27'h0000023e, 5'd3, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c5, 5'd20, 27'h0000031b, 5'd12, 27'h00000384, 32'h00000400,
  1'd1,  5'd9, 27'h0000016e, 5'd21, 27'h000000c6, 5'd25, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d9, 5'd3, 27'h000002d8, 5'd5, 27'h0000033c, 32'h00000400,
  1'd1,  5'd16, 27'h000002f3, 5'd2, 27'h0000008a, 5'd18, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d8, 5'd2, 27'h00000096, 5'd26, 27'h0000020e, 32'h00000400,
  1'd1,  5'd19, 27'h0000010f, 5'd11, 27'h0000018b, 5'd4, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000389, 5'd13, 27'h0000003e, 5'd14, 27'h000000b3, 32'h00000400,
  1'd1,  5'd20, 27'h00000048, 5'd13, 27'h00000212, 5'd22, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000004b, 5'd23, 27'h0000000e, 5'd2, 27'h0000000a, 32'h00000400,
  1'd1,  5'd19, 27'h000000c0, 5'd22, 27'h000002ce, 5'd11, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000226, 5'd25, 27'h00000270, 5'd22, 27'h00000356, 32'h00000400,
  1'd1,  5'd28, 27'h00000151, 5'd4, 27'h0000000f, 5'd0, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000334, 5'd3, 27'h0000036f, 5'd12, 27'h0000008d, 32'h00000400,
  1'd1,  5'd26, 27'h000003b0, 5'd3, 27'h00000158, 5'd21, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000397, 5'd13, 27'h00000115, 5'd4, 27'h00000239, 32'h00000400,
  1'd1,  5'd28, 27'h00000213, 5'd12, 27'h0000011b, 5'd12, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ea, 5'd12, 27'h000000b3, 5'd24, 27'h000003ed, 32'h00000400,
  1'd1,  5'd29, 27'h000002dc, 5'd25, 27'h0000011c, 5'd1, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ee, 5'd23, 27'h0000025a, 5'd15, 27'h00000192, 32'h00000400,
  1'd1,  5'd28, 27'h00000242, 5'd22, 27'h00000242, 5'd21, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000222, 5'd2, 27'h000003c8, 5'd4, 27'h00000341, 32'h00000400,
  1'd1,  5'd7, 27'h00000109, 5'd1, 27'h0000016d, 5'd12, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000396, 5'd3, 27'h000002a0, 5'd25, 27'h00000303, 32'h00000400,
  1'd1,  5'd10, 27'h000000a3, 5'd13, 27'h0000024e, 5'd5, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e6, 5'd10, 27'h00000238, 5'd20, 27'h000000bc, 32'h00000400,
  1'd1,  5'd10, 27'h000000cb, 5'd12, 27'h000003bb, 5'd28, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001f3, 5'd25, 27'h00000227, 5'd8, 27'h00000083, 32'h00000400,
  1'd1,  5'd7, 27'h0000023e, 5'd24, 27'h00000081, 5'd16, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000373, 5'd23, 27'h00000266, 5'd30, 27'h00000260, 32'h00000400,
  1'd1,  5'd16, 27'h000002c4, 5'd2, 27'h00000157, 5'd3, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000028, 5'd4, 27'h000000c3, 5'd11, 27'h0000005d, 32'h00000400,
  1'd1,  5'd17, 27'h00000277, 5'd0, 27'h0000029c, 5'd20, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000017a, 5'd12, 27'h00000301, 5'd8, 27'h000001db, 32'h00000400,
  1'd1,  5'd20, 27'h000000e6, 5'd13, 27'h000000c1, 5'd19, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000351, 5'd11, 27'h0000015c, 5'd26, 27'h000003e5, 32'h00000400,
  1'd1,  5'd16, 27'h0000020e, 5'd25, 27'h00000186, 5'd5, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ee, 5'd22, 27'h0000024c, 5'd18, 27'h000002a0, 32'h00000400,
  1'd1,  5'd19, 27'h0000006d, 5'd23, 27'h0000029a, 5'd26, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000321, 5'd0, 27'h000001a0, 5'd8, 27'h00000011, 32'h00000400,
  1'd1,  5'd29, 27'h00000198, 5'd3, 27'h00000303, 5'd16, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a3, 5'd3, 27'h0000036e, 5'd30, 27'h000002bf, 32'h00000400,
  1'd1,  5'd27, 27'h000000b2, 5'd14, 27'h00000001, 5'd8, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000274, 5'd11, 27'h00000086, 5'd20, 27'h00000094, 32'h00000400,
  1'd1,  5'd30, 27'h00000277, 5'd10, 27'h0000030c, 5'd27, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000249, 5'd25, 27'h000001b0, 5'd8, 27'h000002bb, 32'h00000400,
  1'd1,  5'd26, 27'h000002d2, 5'd21, 27'h000000dc, 5'd18, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000038d, 5'd25, 27'h00000193, 5'd29, 27'h0000026b, 32'h00000400,
  1'd1,  5'd7, 27'h00000131, 5'd9, 27'h000002f2, 5'd3, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000119, 5'd8, 27'h000000f7, 5'd13, 27'h00000352, 32'h00000400,
  1'd1,  5'd6, 27'h00000017, 5'd7, 27'h00000152, 5'd20, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000301, 5'd17, 27'h00000347, 5'd2, 27'h000003ed, 32'h00000400,
  1'd1,  5'd7, 27'h000002e1, 5'd20, 27'h00000273, 5'd15, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000006d, 5'd19, 27'h00000358, 5'd21, 27'h00000052, 32'h00000400,
  1'd1,  5'd5, 27'h00000280, 5'd26, 27'h0000019c, 5'd0, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000150, 5'd28, 27'h00000011, 5'd14, 27'h00000045, 32'h00000400,
  1'd1,  5'd5, 27'h0000034f, 5'd26, 27'h0000021d, 5'd20, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000105, 5'd6, 27'h00000310, 5'd3, 27'h000003a2, 32'h00000400,
  1'd1,  5'd19, 27'h000003e3, 5'd6, 27'h00000368, 5'd13, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000037, 5'd7, 27'h000002ed, 5'd22, 27'h00000140, 32'h00000400,
  1'd1,  5'd20, 27'h000001d9, 5'd20, 27'h0000026b, 5'd3, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000028b, 5'd19, 27'h000000fd, 5'd14, 27'h000000be, 32'h00000400,
  1'd1,  5'd20, 27'h00000001, 5'd16, 27'h00000048, 5'd23, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000020, 5'd29, 27'h00000218, 5'd1, 27'h00000181, 32'h00000400,
  1'd1,  5'd18, 27'h00000333, 5'd30, 27'h000002af, 5'd11, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000051, 5'd28, 27'h0000022a, 5'd24, 27'h0000002c, 32'h00000400,
  1'd1,  5'd30, 27'h0000034f, 5'd5, 27'h000000c7, 5'd1, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000051, 5'd7, 27'h000003a6, 5'd12, 27'h000001b8, 32'h00000400,
  1'd1,  5'd26, 27'h00000047, 5'd8, 27'h0000028c, 5'd23, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003fb, 5'd20, 27'h00000132, 5'd3, 27'h000003e0, 32'h00000400,
  1'd1,  5'd29, 27'h000003ea, 5'd20, 27'h00000229, 5'd11, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000037c, 5'd19, 27'h0000025d, 5'd21, 27'h000002b4, 32'h00000400,
  1'd1,  5'd26, 27'h0000014d, 5'd29, 27'h000002fd, 5'd3, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000014c, 5'd28, 27'h00000224, 5'd14, 27'h00000214, 32'h00000400,
  1'd1,  5'd30, 27'h0000007a, 5'd26, 27'h000000f7, 5'd24, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000212, 5'd7, 27'h00000274, 5'd10, 27'h000000ee, 32'h00000400,
  1'd1,  5'd9, 27'h00000037, 5'd7, 27'h000002dc, 5'd17, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f3, 5'd9, 27'h0000017d, 5'd26, 27'h000003a2, 32'h00000400,
  1'd1,  5'd8, 27'h000001b8, 5'd15, 27'h0000032d, 5'd8, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000298, 5'd17, 27'h0000007e, 5'd16, 27'h0000004f, 32'h00000400,
  1'd1,  5'd9, 27'h000003d7, 5'd18, 27'h0000026f, 5'd26, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000134, 5'd28, 27'h0000028e, 5'd5, 27'h000003de, 32'h00000400,
  1'd1,  5'd5, 27'h0000011d, 5'd29, 27'h0000009c, 5'd19, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000114, 5'd27, 27'h00000335, 5'd26, 27'h000000ab, 32'h00000400,
  1'd1,  5'd18, 27'h000002f9, 5'd8, 27'h000000fc, 5'd9, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000287, 5'd7, 27'h00000339, 5'd16, 27'h0000002e, 32'h00000400,
  1'd1,  5'd15, 27'h00000286, 5'd8, 27'h00000288, 5'd26, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000024d, 5'd15, 27'h0000025b, 5'd5, 27'h000002ac, 32'h00000400,
  1'd1,  5'd20, 27'h00000243, 5'd19, 27'h00000071, 5'd20, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000a8, 5'd18, 27'h00000131, 5'd26, 27'h000001b3, 32'h00000400,
  1'd1,  5'd17, 27'h00000056, 5'd27, 27'h000002a9, 5'd7, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000299, 5'd26, 27'h00000081, 5'd16, 27'h00000116, 32'h00000400,
  1'd1,  5'd16, 27'h00000002, 5'd28, 27'h0000030d, 5'd26, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c8, 5'd6, 27'h000000c4, 5'd6, 27'h0000032f, 32'h00000400,
  1'd1,  5'd29, 27'h00000116, 5'd8, 27'h000002a2, 5'd18, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000186, 5'd8, 27'h00000135, 5'd28, 27'h00000202, 32'h00000400,
  1'd1,  5'd29, 27'h00000354, 5'd16, 27'h000000af, 5'd8, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000187, 5'd20, 27'h0000024c, 5'd17, 27'h0000009e, 32'h00000400,
  1'd1,  5'd27, 27'h00000208, 5'd20, 27'h0000023b, 5'd26, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000001c, 5'd29, 27'h000002a9, 5'd5, 27'h0000013a, 32'h00000400,
  1'd1,  5'd28, 27'h0000030c, 5'd30, 27'h000001a6, 5'd18, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e9, 5'd29, 27'h00000272, 5'd28, 27'h00000198, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000112, 5'd3, 27'h000001f3, 5'd0, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000160, 5'd0, 27'h00000095, 5'd11, 27'h000003d4, 32'h00000400,
  1'd1,  5'd2, 27'h00000152, 5'd0, 27'h00000217, 5'd20, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003ff, 5'd13, 27'h00000396, 5'd3, 27'h00000179, 32'h00000400,
  1'd1,  5'd1, 27'h0000022f, 5'd12, 27'h0000002c, 5'd13, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000007e, 5'd10, 27'h00000223, 5'd22, 27'h000000de, 32'h00000400,
  1'd1,  5'd3, 27'h0000010a, 5'd24, 27'h00000231, 5'd4, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000006c, 5'd23, 27'h000003fc, 5'd11, 27'h00000278, 32'h00000400,
  1'd1,  5'd2, 27'h000002a0, 5'd24, 27'h0000002d, 5'd23, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003bd, 5'd2, 27'h000001eb, 5'd1, 27'h0000037e, 32'h00000400,
  1'd1,  5'd12, 27'h000001a1, 5'd3, 27'h000002f2, 5'd13, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000d9, 5'd4, 27'h000003c5, 5'd22, 27'h0000024f, 32'h00000400,
  1'd1,  5'd11, 27'h0000034b, 5'd14, 27'h00000127, 5'd1, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000158, 5'd10, 27'h00000177, 5'd10, 27'h0000018b, 32'h00000400,
  1'd1,  5'd11, 27'h00000106, 5'd11, 27'h000002b1, 5'd25, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fc, 5'd23, 27'h000003fb, 5'd3, 27'h000001a8, 32'h00000400,
  1'd1,  5'd10, 27'h0000024b, 5'd22, 27'h0000016f, 5'd11, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a8, 5'd22, 27'h000002af, 5'd21, 27'h00000245, 32'h00000400,
  1'd1,  5'd25, 27'h0000017d, 5'd3, 27'h000003b2, 5'd1, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000393, 5'd4, 27'h00000031, 5'd13, 27'h0000013c, 32'h00000400,
  1'd1,  5'd23, 27'h0000024d, 5'd3, 27'h0000003b, 5'd22, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000293, 5'd15, 27'h00000120, 5'd3, 27'h0000012b, 32'h00000400,
  1'd1,  5'd24, 27'h00000210, 5'd14, 27'h000003fd, 5'd14, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002ff, 5'd13, 27'h0000039b, 5'd22, 27'h00000387, 32'h00000400,
  1'd1,  5'd24, 27'h000001ff, 5'd25, 27'h000000f0, 5'd2, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000212, 5'd23, 27'h0000029a, 5'd12, 27'h000002d3, 32'h00000400,
  1'd1,  5'd21, 27'h0000004b, 5'd22, 27'h000000ab, 5'd21, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000392, 5'd3, 27'h00000279, 5'd8, 27'h00000345, 32'h00000400,
  1'd1,  5'd4, 27'h00000040, 5'd3, 27'h00000324, 5'd16, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e6, 5'd1, 27'h0000013d, 5'd28, 27'h00000169, 32'h00000400,
  1'd1,  5'd0, 27'h000001df, 5'd12, 27'h0000039a, 5'd8, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003e4, 5'd12, 27'h00000293, 5'd20, 27'h000000fa, 32'h00000400,
  1'd1,  5'd1, 27'h0000002c, 5'd11, 27'h000000ad, 5'd26, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a8, 5'd22, 27'h00000066, 5'd8, 27'h00000364, 32'h00000400,
  1'd1,  5'd0, 27'h00000241, 5'd20, 27'h000003ab, 5'd17, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000074, 5'd24, 27'h00000040, 5'd29, 27'h000002e2, 32'h00000400,
  1'd1,  5'd11, 27'h000001f3, 5'd0, 27'h00000269, 5'd6, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003c5, 5'd1, 27'h0000001c, 5'd17, 27'h000000db, 32'h00000400,
  1'd1,  5'd11, 27'h000003dc, 5'd0, 27'h00000168, 5'd27, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000e6, 5'd11, 27'h00000359, 5'd8, 27'h00000390, 32'h00000400,
  1'd1,  5'd13, 27'h00000311, 5'd11, 27'h00000014, 5'd18, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000021c, 5'd10, 27'h000003e2, 5'd29, 27'h00000179, 32'h00000400,
  1'd1,  5'd10, 27'h000003b6, 5'd23, 27'h0000019a, 5'd9, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000021c, 5'd25, 27'h00000213, 5'd17, 27'h00000279, 32'h00000400,
  1'd1,  5'd13, 27'h000003fe, 5'd20, 27'h000002b3, 5'd30, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e1, 5'd0, 27'h00000184, 5'd8, 27'h00000053, 32'h00000400,
  1'd1,  5'd25, 27'h00000345, 5'd5, 27'h0000000c, 5'd20, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000032a, 5'd0, 27'h00000116, 5'd29, 27'h0000003d, 32'h00000400,
  1'd1,  5'd24, 27'h000000a6, 5'd12, 27'h00000270, 5'd5, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002aa, 5'd13, 27'h00000177, 5'd20, 27'h00000267, 32'h00000400,
  1'd1,  5'd25, 27'h0000008b, 5'd13, 27'h000002d7, 5'd26, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000022c, 5'd20, 27'h000002fb, 5'd6, 27'h00000174, 32'h00000400,
  1'd1,  5'd24, 27'h00000125, 5'd22, 27'h00000104, 5'd20, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b3, 5'd23, 27'h000001c8, 5'd30, 27'h000000bd, 32'h00000400,
  1'd1,  5'd4, 27'h000000ee, 5'd6, 27'h000002df, 5'd0, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000036a, 5'd8, 27'h000000e5, 5'd12, 27'h000003e8, 32'h00000400,
  1'd1,  5'd3, 27'h00000195, 5'd9, 27'h000003aa, 5'd21, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f3, 5'd19, 27'h00000086, 5'd0, 27'h000002bd, 32'h00000400,
  1'd1,  5'd1, 27'h0000036e, 5'd15, 27'h00000218, 5'd10, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003ae, 5'd16, 27'h00000014, 5'd24, 27'h0000036f, 32'h00000400,
  1'd1,  5'd4, 27'h00000368, 5'd26, 27'h00000297, 5'd0, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000082, 5'd26, 27'h000001a7, 5'd12, 27'h000000c9, 32'h00000400,
  1'd1,  5'd2, 27'h000003eb, 5'd30, 27'h00000110, 5'd23, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001b2, 5'd7, 27'h0000014a, 5'd1, 27'h0000009a, 32'h00000400,
  1'd1,  5'd11, 27'h0000028c, 5'd5, 27'h0000015d, 5'd14, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a2, 5'd9, 27'h0000039a, 5'd21, 27'h00000210, 32'h00000400,
  1'd1,  5'd11, 27'h0000032a, 5'd18, 27'h00000125, 5'd2, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000099, 5'd19, 27'h000001ef, 5'd14, 27'h000001d9, 32'h00000400,
  1'd1,  5'd12, 27'h00000051, 5'd18, 27'h000002ca, 5'd20, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000309, 5'd27, 27'h00000116, 5'd4, 27'h000001bd, 32'h00000400,
  1'd1,  5'd13, 27'h000000da, 5'd30, 27'h00000288, 5'd14, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000378, 5'd26, 27'h00000220, 5'd21, 27'h0000036f, 32'h00000400,
  1'd1,  5'd21, 27'h0000003b, 5'd5, 27'h00000354, 5'd1, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000018a, 5'd8, 27'h00000142, 5'd11, 27'h000003f7, 32'h00000400,
  1'd1,  5'd21, 27'h00000305, 5'd9, 27'h0000037d, 5'd20, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000199, 5'd16, 27'h00000352, 5'd3, 27'h0000024a, 32'h00000400,
  1'd1,  5'd21, 27'h00000232, 5'd17, 27'h00000200, 5'd11, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000014c, 5'd20, 27'h00000065, 5'd24, 27'h00000270, 32'h00000400,
  1'd1,  5'd21, 27'h00000222, 5'd26, 27'h0000026e, 5'd4, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003c8, 5'd27, 27'h0000011a, 5'd15, 27'h000001cb, 32'h00000400,
  1'd1,  5'd22, 27'h0000005e, 5'd28, 27'h00000172, 5'd24, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000f4, 5'd10, 27'h00000065, 5'd8, 27'h0000003f, 32'h00000400,
  1'd1,  5'd4, 27'h000001f5, 5'd5, 27'h0000023a, 5'd19, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001f9, 5'd9, 27'h000000e1, 5'd30, 27'h00000326, 32'h00000400,
  1'd1,  5'd3, 27'h000001f0, 5'd18, 27'h0000031d, 5'd10, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000198, 5'd19, 27'h000001f0, 5'd16, 27'h000001fd, 32'h00000400,
  1'd1,  5'd2, 27'h00000240, 5'd17, 27'h00000249, 5'd26, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000193, 5'd26, 27'h00000077, 5'd7, 27'h0000024f, 32'h00000400,
  1'd1,  5'd4, 27'h00000170, 5'd26, 27'h00000325, 5'd16, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001b8, 5'd28, 27'h00000312, 5'd26, 27'h0000017d, 32'h00000400,
  1'd1,  5'd13, 27'h00000245, 5'd7, 27'h000001c6, 5'd6, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000e9, 5'd5, 27'h000000ef, 5'd16, 27'h00000305, 32'h00000400,
  1'd1,  5'd10, 27'h00000187, 5'd7, 27'h000002d8, 5'd26, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b8, 5'd20, 27'h0000007d, 5'd9, 27'h000001bb, 32'h00000400,
  1'd1,  5'd12, 27'h00000400, 5'd19, 27'h000003cc, 5'd20, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000198, 5'd19, 27'h000003a2, 5'd30, 27'h00000024, 32'h00000400,
  1'd1,  5'd11, 27'h00000276, 5'd27, 27'h0000002b, 5'd7, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f5, 5'd28, 27'h000000ee, 5'd17, 27'h0000003d, 32'h00000400,
  1'd1,  5'd15, 27'h000001bb, 5'd28, 27'h00000312, 5'd25, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002b8, 5'd8, 27'h00000139, 5'd8, 27'h000002ec, 32'h00000400,
  1'd1,  5'd24, 27'h000002d2, 5'd6, 27'h00000334, 5'd15, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000320, 5'd9, 27'h00000305, 5'd27, 27'h000003aa, 32'h00000400,
  1'd1,  5'd21, 27'h0000020a, 5'd15, 27'h00000213, 5'd8, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000014, 5'd18, 27'h00000314, 5'd15, 27'h00000229, 32'h00000400,
  1'd1,  5'd21, 27'h00000258, 5'd19, 27'h00000045, 5'd29, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000259, 5'd27, 27'h00000211, 5'd6, 27'h000000d3, 32'h00000400,
  1'd1,  5'd22, 27'h00000011, 5'd28, 27'h000002e4, 5'd19, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d7, 5'd27, 27'h00000029, 5'd26, 27'h00000190, 32'h00000400,
  1'd1,  5'd7, 27'h0000000d, 5'd2, 27'h0000035d, 5'd7, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000123, 5'd0, 27'h0000024b, 5'd17, 27'h0000008c, 32'h00000400,
  1'd1,  5'd9, 27'h00000296, 5'd1, 27'h000002d1, 5'd27, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000016c, 5'd11, 27'h00000051, 5'd2, 27'h00000037, 32'h00000400,
  1'd1,  5'd6, 27'h000001ef, 5'd14, 27'h000003b9, 5'd14, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000026f, 5'd10, 27'h0000020e, 5'd24, 27'h00000220, 32'h00000400,
  1'd1,  5'd7, 27'h00000289, 5'd23, 27'h0000035d, 5'd3, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000199, 5'd23, 27'h000000c1, 5'd10, 27'h000002a1, 32'h00000400,
  1'd1,  5'd10, 27'h0000004a, 5'd21, 27'h00000002, 5'd21, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000138, 5'd4, 27'h0000020c, 5'd9, 27'h000000bd, 32'h00000400,
  1'd1,  5'd18, 27'h000000ba, 5'd1, 27'h00000242, 5'd19, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002f6, 5'd2, 27'h00000331, 5'd28, 27'h0000039c, 32'h00000400,
  1'd1,  5'd19, 27'h000003f9, 5'd13, 27'h000000b4, 5'd4, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b1, 5'd12, 27'h0000008f, 5'd11, 27'h0000027e, 32'h00000400,
  1'd1,  5'd16, 27'h000002f5, 5'd13, 27'h00000234, 5'd22, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000233, 5'd24, 27'h0000015a, 5'd1, 27'h0000003f, 32'h00000400,
  1'd1,  5'd17, 27'h0000023a, 5'd25, 27'h000002ec, 5'd14, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000037, 5'd24, 27'h0000015b, 5'd21, 27'h000002ab, 32'h00000400,
  1'd1,  5'd29, 27'h0000000e, 5'd3, 27'h00000136, 5'd4, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000010, 5'd2, 27'h00000330, 5'd11, 27'h000001f8, 32'h00000400,
  1'd1,  5'd26, 27'h00000121, 5'd4, 27'h0000020e, 5'd20, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000193, 5'd13, 27'h000003f1, 5'd0, 27'h000003df, 32'h00000400,
  1'd1,  5'd26, 27'h000000d6, 5'd14, 27'h000000eb, 5'd12, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000338, 5'd11, 27'h00000204, 5'd25, 27'h000002b8, 32'h00000400,
  1'd1,  5'd30, 27'h000001be, 5'd21, 27'h0000023b, 5'd5, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b1, 5'd25, 27'h000002ca, 5'd14, 27'h0000029e, 32'h00000400,
  1'd1,  5'd27, 27'h000003dd, 5'd21, 27'h00000035, 5'd23, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000256, 5'd0, 27'h000000d1, 5'd0, 27'h000003e1, 32'h00000400,
  1'd1,  5'd9, 27'h0000000e, 5'd4, 27'h00000001, 5'd11, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000303, 5'd1, 27'h0000039b, 5'd21, 27'h000003b7, 32'h00000400,
  1'd1,  5'd9, 27'h000001b5, 5'd11, 27'h000002b4, 5'd5, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000010, 5'd12, 27'h00000284, 5'd16, 27'h000000f3, 32'h00000400,
  1'd1,  5'd7, 27'h00000075, 5'd10, 27'h0000019e, 5'd30, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000004d, 5'd24, 27'h00000206, 5'd9, 27'h000000f2, 32'h00000400,
  1'd1,  5'd9, 27'h000001c0, 5'd24, 27'h0000002d, 5'd18, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001db, 5'd20, 27'h000003f2, 5'd29, 27'h0000011c, 32'h00000400,
  1'd1,  5'd16, 27'h00000216, 5'd4, 27'h00000378, 5'd0, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000173, 5'd2, 27'h000003a9, 5'd11, 27'h00000063, 32'h00000400,
  1'd1,  5'd19, 27'h00000254, 5'd2, 27'h00000196, 5'd24, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f1, 5'd11, 27'h00000042, 5'd8, 27'h00000391, 32'h00000400,
  1'd1,  5'd16, 27'h0000016c, 5'd13, 27'h00000171, 5'd18, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000025, 5'd11, 27'h0000012e, 5'd30, 27'h0000022e, 32'h00000400,
  1'd1,  5'd20, 27'h0000024c, 5'd22, 27'h0000006d, 5'd9, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000007a, 5'd21, 27'h000002ed, 5'd20, 27'h0000008b, 32'h00000400,
  1'd1,  5'd20, 27'h000000ef, 5'd23, 27'h0000028a, 5'd29, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003fe, 5'd1, 27'h0000011c, 5'd8, 27'h00000286, 32'h00000400,
  1'd1,  5'd27, 27'h0000022d, 5'd3, 27'h00000187, 5'd17, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000356, 5'd2, 27'h000003a8, 5'd28, 27'h000003c9, 32'h00000400,
  1'd1,  5'd27, 27'h00000189, 5'd13, 27'h0000014c, 5'd6, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000215, 5'd15, 27'h00000009, 5'd16, 27'h000003df, 32'h00000400,
  1'd1,  5'd30, 27'h0000023d, 5'd12, 27'h00000364, 5'd27, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000032, 5'd23, 27'h000001c5, 5'd7, 27'h00000236, 32'h00000400,
  1'd1,  5'd26, 27'h000000a2, 5'd25, 27'h00000162, 5'd15, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000d5, 5'd24, 27'h00000261, 5'd29, 27'h000001a7, 32'h00000400,
  1'd1,  5'd9, 27'h000003db, 5'd7, 27'h00000015, 5'd2, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000325, 5'd10, 27'h00000096, 5'd12, 27'h000003d1, 32'h00000400,
  1'd1,  5'd5, 27'h00000327, 5'd8, 27'h00000206, 5'd23, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000157, 5'd16, 27'h00000217, 5'd4, 27'h000003ce, 32'h00000400,
  1'd1,  5'd9, 27'h000000e0, 5'd15, 27'h00000388, 5'd15, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000331, 5'd16, 27'h0000008c, 5'd22, 27'h000002f4, 32'h00000400,
  1'd1,  5'd6, 27'h000001f8, 5'd30, 27'h000000c1, 5'd3, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000044, 5'd26, 27'h00000151, 5'd11, 27'h000002f8, 32'h00000400,
  1'd1,  5'd6, 27'h000003c6, 5'd26, 27'h0000026f, 5'd22, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002e8, 5'd5, 27'h00000199, 5'd0, 27'h000002ea, 32'h00000400,
  1'd1,  5'd20, 27'h00000094, 5'd7, 27'h0000008b, 5'd14, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000238, 5'd8, 27'h000000ca, 5'd22, 27'h00000166, 32'h00000400,
  1'd1,  5'd17, 27'h00000151, 5'd17, 27'h0000029b, 5'd2, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000265, 5'd18, 27'h00000142, 5'd14, 27'h00000290, 32'h00000400,
  1'd1,  5'd17, 27'h0000011e, 5'd18, 27'h00000005, 5'd24, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019b, 5'd27, 27'h0000001d, 5'd3, 27'h000001fd, 32'h00000400,
  1'd1,  5'd16, 27'h000003a0, 5'd30, 27'h00000149, 5'd15, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000074, 5'd27, 27'h00000382, 5'd24, 27'h00000325, 32'h00000400,
  1'd1,  5'd29, 27'h000003f2, 5'd10, 27'h0000001e, 5'd3, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003aa, 5'd6, 27'h00000257, 5'd14, 27'h000000e6, 32'h00000400,
  1'd1,  5'd25, 27'h00000378, 5'd8, 27'h00000012, 5'd22, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000109, 5'd17, 27'h00000222, 5'd3, 27'h000003eb, 32'h00000400,
  1'd1,  5'd28, 27'h000002c4, 5'd18, 27'h0000030a, 5'd13, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021f, 5'd19, 27'h000001a0, 5'd24, 27'h00000353, 32'h00000400,
  1'd1,  5'd28, 27'h00000015, 5'd30, 27'h000000f1, 5'd1, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023a, 5'd27, 27'h00000373, 5'd14, 27'h000001f6, 32'h00000400,
  1'd1,  5'd28, 27'h000000ed, 5'd27, 27'h00000208, 5'd21, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c8, 5'd5, 27'h000001b2, 5'd5, 27'h00000123, 32'h00000400,
  1'd1,  5'd9, 27'h0000025f, 5'd8, 27'h000003ef, 5'd18, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021e, 5'd5, 27'h00000106, 5'd26, 27'h000002c1, 32'h00000400,
  1'd1,  5'd8, 27'h00000378, 5'd16, 27'h00000049, 5'd8, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000037, 5'd17, 27'h00000391, 5'd15, 27'h00000256, 32'h00000400,
  1'd1,  5'd7, 27'h00000262, 5'd17, 27'h00000231, 5'd27, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000226, 5'd28, 27'h0000024b, 5'd9, 27'h000002a5, 32'h00000400,
  1'd1,  5'd7, 27'h000000ca, 5'd25, 27'h000003ce, 5'd19, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ab, 5'd27, 27'h00000239, 5'd26, 27'h0000010c, 32'h00000400,
  1'd1,  5'd18, 27'h000000b2, 5'd10, 27'h0000000c, 5'd8, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000017, 5'd6, 27'h000001c4, 5'd18, 27'h000003a4, 32'h00000400,
  1'd1,  5'd16, 27'h00000265, 5'd5, 27'h00000276, 5'd29, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000008e, 5'd17, 27'h000002df, 5'd8, 27'h0000024a, 32'h00000400,
  1'd1,  5'd18, 27'h00000361, 5'd18, 27'h000002b4, 5'd16, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000347, 5'd17, 27'h000001de, 5'd29, 27'h0000006f, 32'h00000400,
  1'd1,  5'd20, 27'h0000022c, 5'd26, 27'h00000131, 5'd6, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000010c, 5'd26, 27'h000001ad, 5'd16, 27'h00000172, 32'h00000400,
  1'd1,  5'd17, 27'h00000191, 5'd26, 27'h00000398, 5'd30, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001fc, 5'd8, 27'h00000097, 5'd9, 27'h00000290, 32'h00000400,
  1'd1,  5'd26, 27'h000003d4, 5'd8, 27'h000003aa, 5'd16, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000036c, 5'd9, 27'h000000ae, 5'd29, 27'h000002c8, 32'h00000400,
  1'd1,  5'd25, 27'h00000377, 5'd17, 27'h000003e3, 5'd8, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000341, 5'd17, 27'h0000019b, 5'd19, 27'h00000361, 32'h00000400,
  1'd1,  5'd27, 27'h000000eb, 5'd16, 27'h000003e7, 5'd26, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f5, 5'd27, 27'h00000037, 5'd6, 27'h0000035d, 32'h00000400,
  1'd1,  5'd30, 27'h000003be, 5'd29, 27'h00000397, 5'd17, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d4, 5'd28, 27'h000003c6, 5'd25, 27'h000003af, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h00000075, 5'd0, 27'h000002ce, 5'd4, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000104, 5'd0, 27'h00000103, 5'd13, 27'h00000075, 32'h00000400,
  1'd1,  5'd4, 27'h0000017a, 5'd1, 27'h0000018f, 5'd22, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000189, 5'd12, 27'h000000a3, 5'd1, 27'h000000c6, 32'h00000400,
  1'd1,  5'd3, 27'h00000379, 5'd11, 27'h0000021f, 5'd11, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000254, 5'd12, 27'h000003dc, 5'd20, 27'h00000362, 32'h00000400,
  1'd1,  5'd4, 27'h000002bb, 5'd25, 27'h00000225, 5'd3, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000129, 5'd21, 27'h00000354, 5'd15, 27'h00000068, 32'h00000400,
  1'd1,  5'd0, 27'h000002e5, 5'd20, 27'h000003c4, 5'd20, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000001c, 5'd5, 27'h0000001b, 5'd4, 27'h00000326, 32'h00000400,
  1'd1,  5'd10, 27'h000003af, 5'd5, 27'h00000024, 5'd11, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000015b, 5'd0, 27'h000001ef, 5'd23, 27'h0000037c, 32'h00000400,
  1'd1,  5'd11, 27'h000002f5, 5'd11, 27'h00000242, 5'd1, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000392, 5'd14, 27'h0000029b, 5'd11, 27'h0000011d, 32'h00000400,
  1'd1,  5'd12, 27'h00000356, 5'd12, 27'h0000035c, 5'd22, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ab, 5'd23, 27'h000002cc, 5'd3, 27'h000000f3, 32'h00000400,
  1'd1,  5'd11, 27'h0000025c, 5'd23, 27'h0000022f, 5'd12, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000005a, 5'd21, 27'h00000146, 5'd21, 27'h000000df, 32'h00000400,
  1'd1,  5'd24, 27'h000000b4, 5'd5, 27'h0000006b, 5'd2, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000304, 5'd1, 27'h000003f4, 5'd10, 27'h00000240, 32'h00000400,
  1'd1,  5'd21, 27'h000000c6, 5'd1, 27'h00000151, 5'd25, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000000c, 5'd10, 27'h00000333, 5'd1, 27'h00000064, 32'h00000400,
  1'd1,  5'd21, 27'h00000111, 5'd13, 27'h000002a6, 5'd10, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b6, 5'd13, 27'h00000371, 5'd21, 27'h000003ea, 32'h00000400,
  1'd1,  5'd25, 27'h000002ae, 5'd21, 27'h0000013b, 5'd4, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b5, 5'd25, 27'h000002fa, 5'd12, 27'h000003b7, 32'h00000400,
  1'd1,  5'd24, 27'h0000021d, 5'd23, 27'h00000378, 5'd22, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000317, 5'd0, 27'h000001fe, 5'd7, 27'h00000071, 32'h00000400,
  1'd1,  5'd4, 27'h00000082, 5'd1, 27'h000000c4, 5'd16, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000006f, 5'd3, 27'h000000ea, 5'd28, 27'h00000291, 32'h00000400,
  1'd1,  5'd3, 27'h000000ab, 5'd13, 27'h000000e9, 5'd6, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000007a, 5'd14, 27'h000000f0, 5'd15, 27'h00000366, 32'h00000400,
  1'd1,  5'd0, 27'h000000fe, 5'd10, 27'h0000027e, 5'd28, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002b9, 5'd21, 27'h0000035a, 5'd7, 27'h00000127, 32'h00000400,
  1'd1,  5'd4, 27'h00000085, 5'd23, 27'h000001e6, 5'd18, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000065, 5'd24, 27'h0000020b, 5'd29, 27'h0000035e, 32'h00000400,
  1'd1,  5'd11, 27'h00000294, 5'd3, 27'h000000c0, 5'd8, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001fe, 5'd3, 27'h000000f1, 5'd17, 27'h000002d4, 32'h00000400,
  1'd1,  5'd15, 27'h0000013e, 5'd4, 27'h00000254, 5'd28, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001a6, 5'd11, 27'h00000292, 5'd7, 27'h000002f0, 32'h00000400,
  1'd1,  5'd14, 27'h000001ec, 5'd12, 27'h00000167, 5'd19, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029b, 5'd15, 27'h0000002a, 5'd30, 27'h0000035f, 32'h00000400,
  1'd1,  5'd13, 27'h00000005, 5'd23, 27'h000003ba, 5'd6, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000022d, 5'd23, 27'h000000b6, 5'd15, 27'h00000275, 32'h00000400,
  1'd1,  5'd13, 27'h000001ff, 5'd25, 27'h00000106, 5'd29, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000180, 5'd2, 27'h0000012a, 5'd6, 27'h000001ad, 32'h00000400,
  1'd1,  5'd24, 27'h00000250, 5'd1, 27'h000002f9, 5'd16, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001de, 5'd0, 27'h0000034e, 5'd29, 27'h0000023a, 32'h00000400,
  1'd1,  5'd21, 27'h000001f1, 5'd11, 27'h00000213, 5'd6, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003bd, 5'd12, 27'h0000016b, 5'd17, 27'h000000f4, 32'h00000400,
  1'd1,  5'd22, 27'h000000cd, 5'd15, 27'h0000007f, 5'd30, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000067, 5'd22, 27'h00000060, 5'd5, 27'h00000376, 32'h00000400,
  1'd1,  5'd20, 27'h00000340, 5'd22, 27'h0000036b, 5'd20, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000c6, 5'd24, 27'h00000009, 5'd29, 27'h00000298, 32'h00000400,
  1'd1,  5'd1, 27'h000003f3, 5'd9, 27'h00000103, 5'd4, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000002b, 5'd9, 27'h000002f1, 5'd13, 27'h000003fe, 32'h00000400,
  1'd1,  5'd4, 27'h00000265, 5'd8, 27'h000002df, 5'd20, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000af, 5'd18, 27'h000003aa, 5'd1, 27'h00000254, 32'h00000400,
  1'd1,  5'd3, 27'h00000065, 5'd19, 27'h00000087, 5'd11, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002ea, 5'd20, 27'h00000034, 5'd22, 27'h00000134, 32'h00000400,
  1'd1,  5'd0, 27'h0000001d, 5'd26, 27'h00000296, 5'd4, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ec, 5'd30, 27'h00000083, 5'd12, 27'h00000054, 32'h00000400,
  1'd1,  5'd3, 27'h00000196, 5'd27, 27'h00000364, 5'd21, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000027a, 5'd5, 27'h000001bc, 5'd4, 27'h00000264, 32'h00000400,
  1'd1,  5'd12, 27'h00000000, 5'd5, 27'h000001f4, 5'd14, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000073, 5'd8, 27'h00000058, 5'd23, 27'h000001d7, 32'h00000400,
  1'd1,  5'd14, 27'h000000cc, 5'd20, 27'h000001d5, 5'd2, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000262, 5'd18, 27'h00000397, 5'd14, 27'h00000100, 32'h00000400,
  1'd1,  5'd10, 27'h00000266, 5'd16, 27'h00000087, 5'd21, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d8, 5'd26, 27'h00000291, 5'd1, 27'h0000006f, 32'h00000400,
  1'd1,  5'd12, 27'h000002fa, 5'd30, 27'h000001ed, 5'd10, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001de, 5'd28, 27'h000001be, 5'd21, 27'h0000012a, 32'h00000400,
  1'd1,  5'd24, 27'h000001c3, 5'd5, 27'h0000023b, 5'd3, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ff, 5'd6, 27'h000000f1, 5'd14, 27'h00000332, 32'h00000400,
  1'd1,  5'd25, 27'h0000017e, 5'd6, 27'h000002bb, 5'd23, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000131, 5'd19, 27'h000002e6, 5'd1, 27'h00000354, 32'h00000400,
  1'd1,  5'd22, 27'h00000278, 5'd16, 27'h000000c9, 5'd13, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001c, 5'd15, 27'h00000330, 5'd22, 27'h0000030e, 32'h00000400,
  1'd1,  5'd21, 27'h00000133, 5'd30, 27'h00000231, 5'd0, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f9, 5'd28, 27'h0000038e, 5'd14, 27'h0000018b, 32'h00000400,
  1'd1,  5'd20, 27'h00000341, 5'd28, 27'h0000001b, 5'd21, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000048, 5'd5, 27'h000000bd, 5'd7, 27'h0000006f, 32'h00000400,
  1'd1,  5'd2, 27'h000000a5, 5'd10, 27'h000000ef, 5'd20, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000112, 5'd9, 27'h000003a4, 5'd26, 27'h0000013c, 32'h00000400,
  1'd1,  5'd3, 27'h0000026e, 5'd20, 27'h00000063, 5'd6, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000c6, 5'd17, 27'h00000291, 5'd19, 27'h000001aa, 32'h00000400,
  1'd1,  5'd1, 27'h00000262, 5'd15, 27'h00000217, 5'd30, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000364, 5'd28, 27'h00000218, 5'd6, 27'h00000282, 32'h00000400,
  1'd1,  5'd2, 27'h0000030e, 5'd30, 27'h000002fc, 5'd18, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038a, 5'd29, 27'h000003e4, 5'd29, 27'h000002cc, 32'h00000400,
  1'd1,  5'd12, 27'h0000039e, 5'd8, 27'h00000392, 5'd7, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000000a, 5'd6, 27'h00000272, 5'd18, 27'h00000145, 32'h00000400,
  1'd1,  5'd11, 27'h00000088, 5'd5, 27'h00000175, 5'd29, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000365, 5'd18, 27'h000001e4, 5'd5, 27'h000003d0, 32'h00000400,
  1'd1,  5'd14, 27'h0000013d, 5'd16, 27'h00000308, 5'd17, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003bc, 5'd16, 27'h000002c0, 5'd29, 27'h0000036c, 32'h00000400,
  1'd1,  5'd11, 27'h00000381, 5'd28, 27'h0000009e, 5'd9, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000267, 5'd26, 27'h00000195, 5'd17, 27'h000001d2, 32'h00000400,
  1'd1,  5'd14, 27'h00000263, 5'd27, 27'h000003e6, 5'd26, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000d4, 5'd5, 27'h000001ca, 5'd5, 27'h00000307, 32'h00000400,
  1'd1,  5'd21, 27'h00000108, 5'd9, 27'h0000023b, 5'd15, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000dd, 5'd5, 27'h0000023f, 5'd29, 27'h0000033b, 32'h00000400,
  1'd1,  5'd23, 27'h00000336, 5'd20, 27'h00000177, 5'd7, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b7, 5'd16, 27'h0000015f, 5'd18, 27'h00000226, 32'h00000400,
  1'd1,  5'd25, 27'h000001a4, 5'd17, 27'h00000220, 5'd28, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000258, 5'd30, 27'h000002b5, 5'd5, 27'h000002c9, 32'h00000400,
  1'd1,  5'd25, 27'h00000318, 5'd30, 27'h0000026f, 5'd19, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a3, 5'd29, 27'h000000c4, 5'd28, 27'h000000b0, 32'h00000400,
  1'd1,  5'd7, 27'h000002ae, 5'd2, 27'h00000287, 5'd6, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000cf, 5'd3, 27'h00000052, 5'd19, 27'h000003e3, 32'h00000400,
  1'd1,  5'd6, 27'h00000293, 5'd0, 27'h0000002f, 5'd28, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000328, 5'd12, 27'h0000015a, 5'd4, 27'h00000198, 32'h00000400,
  1'd1,  5'd5, 27'h0000039e, 5'd10, 27'h00000344, 5'd12, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c2, 5'd11, 27'h000001b7, 5'd24, 27'h000000d4, 32'h00000400,
  1'd1,  5'd6, 27'h000001ac, 5'd22, 27'h000000be, 5'd0, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000273, 5'd23, 27'h000002fa, 5'd14, 27'h000003c3, 32'h00000400,
  1'd1,  5'd6, 27'h00000045, 5'd24, 27'h000003be, 5'd22, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001c9, 5'd3, 27'h0000000b, 5'd6, 27'h000001e8, 32'h00000400,
  1'd1,  5'd17, 27'h0000038e, 5'd1, 27'h00000208, 5'd16, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000046, 5'd2, 27'h00000154, 5'd29, 27'h00000082, 32'h00000400,
  1'd1,  5'd19, 27'h00000208, 5'd11, 27'h0000020e, 5'd0, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000046, 5'd10, 27'h0000030c, 5'd11, 27'h00000201, 32'h00000400,
  1'd1,  5'd16, 27'h00000354, 5'd15, 27'h0000018f, 5'd25, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000341, 5'd22, 27'h0000034b, 5'd4, 27'h000000d9, 32'h00000400,
  1'd1,  5'd17, 27'h000002b4, 5'd25, 27'h000001f5, 5'd15, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002be, 5'd20, 27'h000003db, 5'd22, 27'h000000bf, 32'h00000400,
  1'd1,  5'd27, 27'h0000006f, 5'd3, 27'h00000187, 5'd2, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000ce, 5'd1, 27'h00000026, 5'd11, 27'h000000eb, 32'h00000400,
  1'd1,  5'd28, 27'h000001c2, 5'd2, 27'h00000160, 5'd23, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a8, 5'd11, 27'h00000251, 5'd3, 27'h00000337, 32'h00000400,
  1'd1,  5'd26, 27'h0000014b, 5'd14, 27'h0000037f, 5'd10, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000dc, 5'd14, 27'h0000003c, 5'd22, 27'h0000007a, 32'h00000400,
  1'd1,  5'd28, 27'h000003c3, 5'd23, 27'h000000de, 5'd1, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000176, 5'd24, 27'h0000039a, 5'd13, 27'h000001a7, 32'h00000400,
  1'd1,  5'd30, 27'h0000014e, 5'd24, 27'h0000014f, 5'd24, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000a4, 5'd1, 27'h000000cb, 5'd0, 27'h00000069, 32'h00000400,
  1'd1,  5'd8, 27'h00000336, 5'd1, 27'h000000fb, 5'd13, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ec, 5'd0, 27'h000002e8, 5'd22, 27'h000000a1, 32'h00000400,
  1'd1,  5'd8, 27'h000001de, 5'd12, 27'h000000e5, 5'd7, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ea, 5'd11, 27'h00000041, 5'd16, 27'h0000018b, 32'h00000400,
  1'd1,  5'd8, 27'h0000016b, 5'd14, 27'h000002ee, 5'd30, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000313, 5'd21, 27'h000001f7, 5'd6, 27'h00000100, 32'h00000400,
  1'd1,  5'd9, 27'h000003a9, 5'd21, 27'h00000019, 5'd20, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000019b, 5'd24, 27'h0000026a, 5'd26, 27'h00000073, 32'h00000400,
  1'd1,  5'd19, 27'h00000231, 5'd0, 27'h000000fa, 5'd4, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001fe, 5'd4, 27'h000001a6, 5'd13, 27'h000000ac, 32'h00000400,
  1'd1,  5'd17, 27'h000000d5, 5'd4, 27'h000001d3, 5'd24, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d9, 5'd14, 27'h00000293, 5'd7, 27'h0000023c, 32'h00000400,
  1'd1,  5'd18, 27'h000002e0, 5'd14, 27'h00000009, 5'd19, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000031d, 5'd11, 27'h0000017b, 5'd30, 27'h000000f9, 32'h00000400,
  1'd1,  5'd16, 27'h00000162, 5'd23, 27'h000003ad, 5'd6, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029b, 5'd21, 27'h000000b5, 5'd17, 27'h000002f1, 32'h00000400,
  1'd1,  5'd15, 27'h00000319, 5'd21, 27'h000000f4, 5'd27, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012e, 5'd3, 27'h00000204, 5'd7, 27'h00000197, 32'h00000400,
  1'd1,  5'd28, 27'h00000282, 5'd2, 27'h000001e9, 5'd16, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ed, 5'd2, 27'h000002f3, 5'd27, 27'h0000024a, 32'h00000400,
  1'd1,  5'd28, 27'h000000bb, 5'd14, 27'h000003c3, 5'd9, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000376, 5'd10, 27'h0000037a, 5'd16, 27'h0000013c, 32'h00000400,
  1'd1,  5'd29, 27'h000000cb, 5'd15, 27'h000001dd, 5'd30, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000026b, 5'd22, 27'h0000039d, 5'd5, 27'h000000c4, 32'h00000400,
  1'd1,  5'd30, 27'h000001c1, 5'd25, 27'h00000275, 5'd16, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000372, 5'd23, 27'h0000002a, 5'd28, 27'h00000029, 32'h00000400,
  1'd1,  5'd9, 27'h00000049, 5'd5, 27'h00000154, 5'd0, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000193, 5'd6, 27'h00000230, 5'd10, 27'h000003eb, 32'h00000400,
  1'd1,  5'd5, 27'h0000011a, 5'd5, 27'h00000366, 5'd22, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a1, 5'd16, 27'h00000369, 5'd1, 27'h00000351, 32'h00000400,
  1'd1,  5'd7, 27'h00000029, 5'd18, 27'h000000ef, 5'd14, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000329, 5'd15, 27'h00000231, 5'd25, 27'h00000228, 32'h00000400,
  1'd1,  5'd9, 27'h0000001c, 5'd27, 27'h000003a8, 5'd1, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000323, 5'd26, 27'h00000168, 5'd15, 27'h00000165, 32'h00000400,
  1'd1,  5'd6, 27'h000003dc, 5'd28, 27'h000001d7, 5'd24, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000152, 5'd5, 27'h000003ea, 5'd0, 27'h0000017d, 32'h00000400,
  1'd1,  5'd18, 27'h00000127, 5'd9, 27'h0000003d, 5'd14, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000039c, 5'd8, 27'h00000304, 5'd23, 27'h000001d6, 32'h00000400,
  1'd1,  5'd16, 27'h0000005a, 5'd19, 27'h0000009c, 5'd0, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003ed, 5'd17, 27'h000003f0, 5'd11, 27'h0000031a, 32'h00000400,
  1'd1,  5'd19, 27'h0000003f, 5'd20, 27'h0000027b, 5'd25, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002e6, 5'd26, 27'h000000ba, 5'd4, 27'h00000316, 32'h00000400,
  1'd1,  5'd18, 27'h000002c4, 5'd27, 27'h0000010c, 5'd12, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ec, 5'd28, 27'h0000038a, 5'd21, 27'h0000013f, 32'h00000400,
  1'd1,  5'd30, 27'h00000035, 5'd8, 27'h00000210, 5'd2, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000378, 5'd10, 27'h00000074, 5'd12, 27'h0000028d, 32'h00000400,
  1'd1,  5'd30, 27'h00000143, 5'd7, 27'h000001b6, 5'd22, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f3, 5'd16, 27'h00000026, 5'd2, 27'h00000300, 32'h00000400,
  1'd1,  5'd28, 27'h000003bf, 5'd16, 27'h00000248, 5'd12, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001f7, 5'd20, 27'h000001cb, 5'd21, 27'h0000034b, 32'h00000400,
  1'd1,  5'd29, 27'h0000026b, 5'd28, 27'h0000010d, 5'd2, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000361, 5'd26, 27'h00000033, 5'd13, 27'h0000038d, 32'h00000400,
  1'd1,  5'd26, 27'h0000006b, 5'd27, 27'h00000356, 5'd24, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001fc, 5'd9, 27'h0000034a, 5'd6, 27'h0000016a, 32'h00000400,
  1'd1,  5'd7, 27'h000001bc, 5'd6, 27'h00000318, 5'd20, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000225, 5'd5, 27'h00000374, 5'd30, 27'h00000393, 32'h00000400,
  1'd1,  5'd5, 27'h0000010b, 5'd16, 27'h0000011d, 5'd5, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000011f, 5'd15, 27'h00000206, 5'd18, 27'h0000024e, 32'h00000400,
  1'd1,  5'd6, 27'h000002c3, 5'd20, 27'h000000dc, 5'd30, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e6, 5'd27, 27'h0000016d, 5'd8, 27'h00000227, 32'h00000400,
  1'd1,  5'd7, 27'h0000006c, 5'd27, 27'h00000348, 5'd18, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002fc, 5'd30, 27'h00000228, 5'd27, 27'h000001b8, 32'h00000400,
  1'd1,  5'd20, 27'h00000091, 5'd8, 27'h000002f5, 5'd6, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000276, 5'd6, 27'h000002f2, 5'd18, 27'h0000023d, 32'h00000400,
  1'd1,  5'd18, 27'h000002b7, 5'd7, 27'h000002af, 5'd29, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000005, 5'd19, 27'h000002d4, 5'd7, 27'h000001a0, 32'h00000400,
  1'd1,  5'd19, 27'h00000167, 5'd19, 27'h000002c9, 5'd20, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003ef, 5'd17, 27'h0000007f, 5'd29, 27'h00000057, 32'h00000400,
  1'd1,  5'd17, 27'h0000038f, 5'd27, 27'h000003b7, 5'd5, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000189, 5'd26, 27'h000001be, 5'd20, 27'h00000144, 32'h00000400,
  1'd1,  5'd19, 27'h00000252, 5'd28, 27'h00000105, 5'd30, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000028f, 5'd8, 27'h00000164, 5'd6, 27'h000002e4, 32'h00000400,
  1'd1,  5'd30, 27'h00000204, 5'd6, 27'h000003c6, 5'd18, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000120, 5'd8, 27'h000000d6, 5'd28, 27'h000002a9, 32'h00000400,
  1'd1,  5'd30, 27'h0000039a, 5'd17, 27'h000000b1, 5'd7, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001a7, 5'd15, 27'h000002d4, 5'd17, 27'h00000362, 32'h00000400,
  1'd1,  5'd28, 27'h000001c0, 5'd19, 27'h00000340, 5'd27, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000000c, 5'd28, 27'h00000046, 5'd8, 27'h00000285, 32'h00000400,
  1'd1,  5'd26, 27'h000000c2, 5'd26, 27'h00000025, 5'd16, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000287, 5'd30, 27'h000001c5, 5'd30, 27'h000003d2, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000002c6, 5'd1, 27'h00000169, 5'd1, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000338, 5'd3, 27'h0000004a, 5'd15, 27'h00000122, 32'h00000400,
  1'd1,  5'd3, 27'h000000cf, 5'd4, 27'h00000353, 5'd21, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000193, 5'd13, 27'h000002b9, 5'd0, 27'h0000031c, 32'h00000400,
  1'd1,  5'd3, 27'h0000034b, 5'd13, 27'h000002fc, 5'd13, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a8, 5'd11, 27'h00000116, 5'd23, 27'h00000152, 32'h00000400,
  1'd1,  5'd0, 27'h00000179, 5'd23, 27'h000001ac, 5'd4, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003dc, 5'd23, 27'h000003c4, 5'd11, 27'h000001e0, 32'h00000400,
  1'd1,  5'd2, 27'h000002e7, 5'd22, 27'h0000029f, 5'd21, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000109, 5'd4, 27'h000001b4, 5'd3, 27'h00000331, 32'h00000400,
  1'd1,  5'd14, 27'h0000022a, 5'd3, 27'h00000160, 5'd12, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000121, 5'd2, 27'h00000085, 5'd22, 27'h00000096, 32'h00000400,
  1'd1,  5'd11, 27'h000002da, 5'd11, 27'h00000279, 5'd1, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000069, 5'd14, 27'h000001fc, 5'd15, 27'h00000065, 32'h00000400,
  1'd1,  5'd13, 27'h000003d3, 5'd12, 27'h00000016, 5'd21, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029f, 5'd23, 27'h000003f7, 5'd1, 27'h000000bb, 32'h00000400,
  1'd1,  5'd12, 27'h0000029d, 5'd23, 27'h0000014f, 5'd13, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000060, 5'd22, 27'h000002bf, 5'd23, 27'h00000125, 32'h00000400,
  1'd1,  5'd24, 27'h00000372, 5'd2, 27'h00000260, 5'd1, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000288, 5'd1, 27'h0000027d, 5'd10, 27'h00000354, 32'h00000400,
  1'd1,  5'd20, 27'h00000377, 5'd4, 27'h000001a6, 5'd20, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000000f, 5'd10, 27'h000001f7, 5'd1, 27'h00000028, 32'h00000400,
  1'd1,  5'd21, 27'h00000190, 5'd12, 27'h00000021, 5'd10, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a2, 5'd10, 27'h0000030d, 5'd25, 27'h000002af, 32'h00000400,
  1'd1,  5'd24, 27'h000001fc, 5'd22, 27'h0000010f, 5'd3, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000f4, 5'd20, 27'h0000037b, 5'd12, 27'h00000140, 32'h00000400,
  1'd1,  5'd23, 27'h00000021, 5'd25, 27'h0000020b, 5'd24, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000029e, 5'd2, 27'h000000cd, 5'd7, 27'h00000333, 32'h00000400,
  1'd1,  5'd0, 27'h000000ef, 5'd1, 27'h000002a2, 5'd16, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002ce, 5'd5, 27'h0000004c, 5'd29, 27'h00000101, 32'h00000400,
  1'd1,  5'd1, 27'h000000e1, 5'd14, 27'h0000020b, 5'd8, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002ae, 5'd13, 27'h000002ec, 5'd16, 27'h0000034a, 32'h00000400,
  1'd1,  5'd0, 27'h000001e9, 5'd12, 27'h0000039d, 5'd28, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b9, 5'd21, 27'h0000017b, 5'd7, 27'h00000020, 32'h00000400,
  1'd1,  5'd1, 27'h000001b5, 5'd24, 27'h0000021a, 5'd18, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000114, 5'd24, 27'h0000039d, 5'd30, 27'h00000098, 32'h00000400,
  1'd1,  5'd13, 27'h000002d1, 5'd0, 27'h000003a7, 5'd10, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ce, 5'd2, 27'h00000328, 5'd20, 27'h0000024a, 32'h00000400,
  1'd1,  5'd14, 27'h0000035f, 5'd0, 27'h000000b1, 5'd30, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000242, 5'd13, 27'h00000224, 5'd9, 27'h000003a9, 32'h00000400,
  1'd1,  5'd13, 27'h00000357, 5'd15, 27'h0000000d, 5'd19, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000276, 5'd12, 27'h000003e2, 5'd30, 27'h00000330, 32'h00000400,
  1'd1,  5'd10, 27'h000002f0, 5'd23, 27'h00000183, 5'd9, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000004e, 5'd24, 27'h0000010e, 5'd20, 27'h00000107, 32'h00000400,
  1'd1,  5'd11, 27'h00000250, 5'd22, 27'h000003ad, 5'd27, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c9, 5'd2, 27'h00000234, 5'd7, 27'h00000258, 32'h00000400,
  1'd1,  5'd22, 27'h00000382, 5'd1, 27'h00000223, 5'd18, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000015f, 5'd1, 27'h0000031d, 5'd26, 27'h00000233, 32'h00000400,
  1'd1,  5'd23, 27'h00000100, 5'd12, 27'h0000006b, 5'd5, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000092, 5'd12, 27'h0000024b, 5'd20, 27'h0000015d, 32'h00000400,
  1'd1,  5'd23, 27'h000003ac, 5'd13, 27'h0000018b, 5'd26, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000005, 5'd21, 27'h00000317, 5'd6, 27'h000002ab, 32'h00000400,
  1'd1,  5'd22, 27'h0000011f, 5'd23, 27'h00000091, 5'd18, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000005c, 5'd20, 27'h000002fd, 5'd27, 27'h00000120, 32'h00000400,
  1'd1,  5'd1, 27'h00000368, 5'd9, 27'h000002af, 5'd1, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000091, 5'd8, 27'h000003ab, 5'd13, 27'h000000e4, 32'h00000400,
  1'd1,  5'd3, 27'h000002cc, 5'd9, 27'h0000031b, 5'd23, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ee, 5'd18, 27'h00000094, 5'd2, 27'h00000259, 32'h00000400,
  1'd1,  5'd0, 27'h00000168, 5'd18, 27'h000003d7, 5'd11, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000067, 5'd20, 27'h00000270, 5'd21, 27'h000001a1, 32'h00000400,
  1'd1,  5'd1, 27'h0000031b, 5'd26, 27'h000002c8, 5'd1, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000206, 5'd28, 27'h000002c4, 5'd13, 27'h00000206, 32'h00000400,
  1'd1,  5'd0, 27'h000002b5, 5'd26, 27'h00000152, 5'd22, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001de, 5'd7, 27'h000001ea, 5'd3, 27'h00000169, 32'h00000400,
  1'd1,  5'd13, 27'h00000050, 5'd8, 27'h000003b4, 5'd12, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000118, 5'd9, 27'h00000368, 5'd22, 27'h00000304, 32'h00000400,
  1'd1,  5'd14, 27'h000002e0, 5'd16, 27'h00000188, 5'd0, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001b9, 5'd16, 27'h0000026e, 5'd11, 27'h0000020e, 32'h00000400,
  1'd1,  5'd10, 27'h000002dc, 5'd17, 27'h000003c3, 5'd22, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000072, 5'd26, 27'h000001ce, 5'd0, 27'h000000b9, 32'h00000400,
  1'd1,  5'd11, 27'h00000204, 5'd27, 27'h000001e5, 5'd13, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000019, 5'd27, 27'h0000039c, 5'd24, 27'h00000087, 32'h00000400,
  1'd1,  5'd22, 27'h0000031a, 5'd10, 27'h000000cb, 5'd1, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000287, 5'd7, 27'h00000333, 5'd10, 27'h000003f6, 32'h00000400,
  1'd1,  5'd21, 27'h000000ef, 5'd5, 27'h0000039a, 5'd24, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a7, 5'd15, 27'h000003ee, 5'd4, 27'h000002e9, 32'h00000400,
  1'd1,  5'd23, 27'h000003bd, 5'd17, 27'h000003e3, 5'd13, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003f9, 5'd18, 27'h00000235, 5'd23, 27'h000001ae, 32'h00000400,
  1'd1,  5'd20, 27'h000003db, 5'd27, 27'h0000005b, 5'd1, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034c, 5'd28, 27'h00000217, 5'd10, 27'h0000018f, 32'h00000400,
  1'd1,  5'd21, 27'h000003a3, 5'd27, 27'h00000353, 5'd23, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000346, 5'd7, 27'h000003f0, 5'd5, 27'h000002b1, 32'h00000400,
  1'd1,  5'd4, 27'h00000144, 5'd9, 27'h00000273, 5'd19, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000137, 5'd7, 27'h0000022a, 5'd26, 27'h00000144, 32'h00000400,
  1'd1,  5'd3, 27'h00000159, 5'd20, 27'h00000205, 5'd9, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000033, 5'd20, 27'h000000de, 5'd15, 27'h000003c7, 32'h00000400,
  1'd1,  5'd1, 27'h0000012a, 5'd16, 27'h00000281, 5'd30, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002df, 5'd27, 27'h0000020c, 5'd9, 27'h000001b4, 32'h00000400,
  1'd1,  5'd1, 27'h00000212, 5'd27, 27'h0000018a, 5'd20, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e4, 5'd30, 27'h00000327, 5'd28, 27'h00000145, 32'h00000400,
  1'd1,  5'd13, 27'h00000278, 5'd8, 27'h00000133, 5'd7, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000299, 5'd9, 27'h0000017f, 5'd19, 27'h00000168, 32'h00000400,
  1'd1,  5'd11, 27'h00000337, 5'd8, 27'h00000198, 5'd29, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029d, 5'd15, 27'h00000232, 5'd7, 27'h0000033b, 32'h00000400,
  1'd1,  5'd14, 27'h000001f2, 5'd19, 27'h00000194, 5'd20, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000b7, 5'd18, 27'h000002cd, 5'd26, 27'h00000120, 32'h00000400,
  1'd1,  5'd11, 27'h00000004, 5'd27, 27'h00000208, 5'd6, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c2, 5'd27, 27'h00000148, 5'd17, 27'h00000046, 32'h00000400,
  1'd1,  5'd12, 27'h0000034c, 5'd29, 27'h000002ed, 5'd30, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e6, 5'd9, 27'h000003e6, 5'd6, 27'h000002d2, 32'h00000400,
  1'd1,  5'd25, 27'h00000296, 5'd5, 27'h000002a6, 5'd18, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000017b, 5'd9, 27'h00000314, 5'd28, 27'h0000014f, 32'h00000400,
  1'd1,  5'd25, 27'h00000150, 5'd19, 27'h0000005b, 5'd5, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000129, 5'd16, 27'h00000336, 5'd18, 27'h00000270, 32'h00000400,
  1'd1,  5'd21, 27'h00000118, 5'd20, 27'h000001e8, 5'd29, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000060, 5'd27, 27'h000001e5, 5'd5, 27'h000002cd, 32'h00000400,
  1'd1,  5'd22, 27'h00000156, 5'd29, 27'h000003bc, 5'd20, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000019d, 5'd26, 27'h00000377, 5'd27, 27'h000002e9, 32'h00000400,
  1'd1,  5'd6, 27'h0000012d, 5'd2, 27'h00000018, 5'd5, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000023f, 5'd4, 27'h000000c8, 5'd19, 27'h00000284, 32'h00000400,
  1'd1,  5'd9, 27'h0000023f, 5'd2, 27'h000003ff, 5'd26, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000011c, 5'd14, 27'h00000219, 5'd4, 27'h000002de, 32'h00000400,
  1'd1,  5'd5, 27'h000001f2, 5'd11, 27'h00000262, 5'd10, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000360, 5'd12, 27'h00000280, 5'd22, 27'h0000021c, 32'h00000400,
  1'd1,  5'd5, 27'h000000ae, 5'd22, 27'h000000e3, 5'd2, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000283, 5'd20, 27'h000002d0, 5'd12, 27'h000001eb, 32'h00000400,
  1'd1,  5'd8, 27'h0000028e, 5'd20, 27'h000002b8, 5'd24, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000107, 5'd1, 27'h0000011e, 5'd6, 27'h000000d9, 32'h00000400,
  1'd1,  5'd19, 27'h000002c6, 5'd0, 27'h000002a6, 5'd17, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002c0, 5'd4, 27'h00000212, 5'd28, 27'h00000131, 32'h00000400,
  1'd1,  5'd20, 27'h00000056, 5'd13, 27'h000002b5, 5'd3, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000012b, 5'd11, 27'h000003ce, 5'd13, 27'h000003fb, 32'h00000400,
  1'd1,  5'd19, 27'h00000105, 5'd11, 27'h000002a7, 5'd25, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000017c, 5'd22, 27'h0000028c, 5'd4, 27'h000001c8, 32'h00000400,
  1'd1,  5'd17, 27'h000002aa, 5'd22, 27'h0000000b, 5'd13, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ef, 5'd20, 27'h000002e1, 5'd22, 27'h000000f2, 32'h00000400,
  1'd1,  5'd29, 27'h0000010c, 5'd1, 27'h00000101, 5'd2, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000d, 5'd0, 27'h00000103, 5'd10, 27'h00000323, 32'h00000400,
  1'd1,  5'd26, 27'h000003ee, 5'd2, 27'h00000336, 5'd24, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002bb, 5'd14, 27'h0000003f, 5'd4, 27'h00000095, 32'h00000400,
  1'd1,  5'd29, 27'h000000c6, 5'd14, 27'h0000015f, 5'd11, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000246, 5'd13, 27'h000002fc, 5'd24, 27'h000000cf, 32'h00000400,
  1'd1,  5'd29, 27'h00000244, 5'd20, 27'h000003f8, 5'd2, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b1, 5'd21, 27'h000002ee, 5'd13, 27'h0000022e, 32'h00000400,
  1'd1,  5'd27, 27'h00000173, 5'd21, 27'h000001b5, 5'd22, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002cf, 5'd3, 27'h000003cb, 5'd0, 27'h00000247, 32'h00000400,
  1'd1,  5'd5, 27'h000002fa, 5'd1, 27'h00000112, 5'd12, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d6, 5'd3, 27'h000000c6, 5'd22, 27'h0000015c, 32'h00000400,
  1'd1,  5'd8, 27'h00000341, 5'd13, 27'h0000003b, 5'd6, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000289, 5'd12, 27'h0000029e, 5'd19, 27'h00000391, 32'h00000400,
  1'd1,  5'd5, 27'h00000313, 5'd15, 27'h00000075, 5'd27, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000025, 5'd25, 27'h00000099, 5'd9, 27'h00000067, 32'h00000400,
  1'd1,  5'd8, 27'h000002f5, 5'd25, 27'h00000183, 5'd17, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000c2, 5'd22, 27'h0000026f, 5'd26, 27'h000001d0, 32'h00000400,
  1'd1,  5'd19, 27'h00000070, 5'd4, 27'h00000039, 5'd0, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000184, 5'd0, 27'h00000387, 5'd15, 27'h0000002e, 32'h00000400,
  1'd1,  5'd15, 27'h000002a2, 5'd4, 27'h000002e8, 5'd25, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000016, 5'd11, 27'h000000d3, 5'd5, 27'h000000cc, 32'h00000400,
  1'd1,  5'd18, 27'h0000035e, 5'd15, 27'h000000e5, 5'd19, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000027d, 5'd11, 27'h00000124, 5'd26, 27'h000003a8, 32'h00000400,
  1'd1,  5'd15, 27'h00000354, 5'd23, 27'h000002ea, 5'd7, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a4, 5'd21, 27'h000003b0, 5'd20, 27'h0000017f, 32'h00000400,
  1'd1,  5'd19, 27'h00000369, 5'd25, 27'h0000034a, 5'd29, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000275, 5'd4, 27'h0000006f, 5'd9, 27'h0000027a, 32'h00000400,
  1'd1,  5'd27, 27'h00000200, 5'd1, 27'h00000282, 5'd18, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002ca, 5'd4, 27'h00000197, 5'd28, 27'h000002cf, 32'h00000400,
  1'd1,  5'd29, 27'h00000366, 5'd14, 27'h00000121, 5'd6, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f5, 5'd15, 27'h0000004d, 5'd15, 27'h000002ab, 32'h00000400,
  1'd1,  5'd26, 27'h00000000, 5'd12, 27'h00000080, 5'd28, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e9, 5'd25, 27'h000002f2, 5'd7, 27'h00000055, 32'h00000400,
  1'd1,  5'd30, 27'h00000391, 5'd21, 27'h00000341, 5'd20, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000018a, 5'd22, 27'h000003c4, 5'd30, 27'h000003d5, 32'h00000400,
  1'd1,  5'd7, 27'h00000033, 5'd9, 27'h000003a7, 5'd4, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003fc, 5'd9, 27'h00000029, 5'd13, 27'h0000021d, 32'h00000400,
  1'd1,  5'd6, 27'h000001bb, 5'd5, 27'h000000ef, 5'd23, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000235, 5'd15, 27'h0000032f, 5'd4, 27'h000002b7, 32'h00000400,
  1'd1,  5'd9, 27'h0000027d, 5'd17, 27'h0000003b, 5'd14, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003b4, 5'd20, 27'h00000044, 5'd22, 27'h000001e0, 32'h00000400,
  1'd1,  5'd8, 27'h00000149, 5'd28, 27'h00000284, 5'd0, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000015, 5'd29, 27'h00000076, 5'd10, 27'h00000318, 32'h00000400,
  1'd1,  5'd6, 27'h00000059, 5'd29, 27'h000001c4, 5'd24, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000130, 5'd8, 27'h00000305, 5'd1, 27'h00000019, 32'h00000400,
  1'd1,  5'd18, 27'h0000009b, 5'd8, 27'h0000011f, 5'd14, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000307, 5'd5, 27'h00000242, 5'd23, 27'h000002e9, 32'h00000400,
  1'd1,  5'd15, 27'h00000236, 5'd16, 27'h00000273, 5'd3, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003a0, 5'd20, 27'h000000af, 5'd10, 27'h000003e2, 32'h00000400,
  1'd1,  5'd20, 27'h000001ca, 5'd15, 27'h00000299, 5'd22, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e9, 5'd29, 27'h000001cb, 5'd2, 27'h000001dd, 32'h00000400,
  1'd1,  5'd18, 27'h00000030, 5'd29, 27'h000003bd, 5'd14, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000121, 5'd29, 27'h0000001d, 5'd20, 27'h000002ff, 32'h00000400,
  1'd1,  5'd25, 27'h00000372, 5'd9, 27'h000001b2, 5'd3, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021d, 5'd8, 27'h00000296, 5'd13, 27'h00000372, 32'h00000400,
  1'd1,  5'd29, 27'h0000034c, 5'd7, 27'h0000022c, 5'd21, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000377, 5'd16, 27'h000001d5, 5'd3, 27'h000000d2, 32'h00000400,
  1'd1,  5'd27, 27'h000000c4, 5'd15, 27'h00000240, 5'd12, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000139, 5'd16, 27'h000001b4, 5'd20, 27'h00000338, 32'h00000400,
  1'd1,  5'd30, 27'h00000081, 5'd28, 27'h00000218, 5'd4, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ad, 5'd28, 27'h0000036a, 5'd12, 27'h00000240, 32'h00000400,
  1'd1,  5'd26, 27'h000000e3, 5'd27, 27'h0000024f, 5'd23, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000215, 5'd5, 27'h00000114, 5'd5, 27'h000002af, 32'h00000400,
  1'd1,  5'd6, 27'h00000265, 5'd7, 27'h000001a3, 5'd19, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000002b, 5'd6, 27'h000002d5, 5'd30, 27'h000003fe, 32'h00000400,
  1'd1,  5'd8, 27'h000000ee, 5'd19, 27'h000001dd, 5'd5, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000334, 5'd16, 27'h000000e7, 5'd18, 27'h000000df, 32'h00000400,
  1'd1,  5'd6, 27'h00000075, 5'd18, 27'h000003dd, 5'd30, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002ba, 5'd29, 27'h00000369, 5'd7, 27'h000002a9, 32'h00000400,
  1'd1,  5'd5, 27'h00000267, 5'd29, 27'h0000020b, 5'd16, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000007b, 5'd30, 27'h0000035b, 5'd26, 27'h0000037a, 32'h00000400,
  1'd1,  5'd16, 27'h00000307, 5'd8, 27'h000000be, 5'd7, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000011d, 5'd6, 27'h0000034e, 5'd17, 27'h000003f1, 32'h00000400,
  1'd1,  5'd18, 27'h000003df, 5'd8, 27'h000003b2, 5'd28, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000038e, 5'd15, 27'h000002f4, 5'd9, 27'h000002c5, 32'h00000400,
  1'd1,  5'd16, 27'h00000164, 5'd16, 27'h00000281, 5'd17, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000013, 5'd17, 27'h000003f5, 5'd28, 27'h000000d5, 32'h00000400,
  1'd1,  5'd16, 27'h000000e4, 5'd29, 27'h00000239, 5'd6, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000228, 5'd29, 27'h0000025c, 5'd15, 27'h000002cf, 32'h00000400,
  1'd1,  5'd18, 27'h00000265, 5'd27, 27'h00000397, 5'd27, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000241, 5'd7, 27'h000001f3, 5'd9, 27'h000003af, 32'h00000400,
  1'd1,  5'd27, 27'h0000013d, 5'd6, 27'h00000165, 5'd20, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000275, 5'd6, 27'h000001de, 5'd26, 27'h00000264, 32'h00000400,
  1'd1,  5'd26, 27'h00000339, 5'd15, 27'h0000035b, 5'd6, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000032a, 5'd15, 27'h0000031f, 5'd16, 27'h000000e2, 32'h00000400,
  1'd1,  5'd27, 27'h0000024b, 5'd16, 27'h000002bd, 5'd28, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001cb, 5'd30, 27'h00000396, 5'd7, 27'h0000022a, 32'h00000400,
  1'd1,  5'd29, 27'h00000028, 5'd26, 27'h0000038d, 5'd19, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d1, 5'd26, 27'h000002b9, 5'd27, 27'h00000098, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h00000078, 5'd2, 27'h000003a0, 5'd0, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d5, 5'd3, 27'h00000263, 5'd12, 27'h00000359, 32'h00000400,
  1'd1,  5'd1, 27'h000000ef, 5'd2, 27'h0000000c, 5'd21, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000205, 5'd11, 27'h0000006e, 5'd0, 27'h0000028a, 32'h00000400,
  1'd1,  5'd1, 27'h000000ac, 5'd12, 27'h000000ff, 5'd11, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000cb, 5'd10, 27'h000001cc, 5'd24, 27'h00000260, 32'h00000400,
  1'd1,  5'd3, 27'h00000252, 5'd20, 27'h000002b0, 5'd4, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000312, 5'd24, 27'h000003df, 5'd12, 27'h0000012e, 32'h00000400,
  1'd1,  5'd2, 27'h0000038b, 5'd21, 27'h0000022b, 5'd25, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003a7, 5'd4, 27'h00000359, 5'd3, 27'h0000035d, 32'h00000400,
  1'd1,  5'd13, 27'h00000390, 5'd1, 27'h0000014f, 5'd14, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000050, 5'd0, 27'h000001d0, 5'd21, 27'h000002c1, 32'h00000400,
  1'd1,  5'd13, 27'h000001cd, 5'd12, 27'h000002d1, 5'd2, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002ce, 5'd12, 27'h000001d1, 5'd11, 27'h000000cc, 32'h00000400,
  1'd1,  5'd14, 27'h0000025b, 5'd13, 27'h000001ad, 5'd20, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000012d, 5'd20, 27'h00000309, 5'd1, 27'h00000303, 32'h00000400,
  1'd1,  5'd11, 27'h000003e7, 5'd25, 27'h0000031b, 5'd12, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000003b, 5'd21, 27'h00000013, 5'd23, 27'h00000157, 32'h00000400,
  1'd1,  5'd25, 27'h0000028e, 5'd4, 27'h00000051, 5'd2, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000230, 5'd3, 27'h00000386, 5'd11, 27'h00000050, 32'h00000400,
  1'd1,  5'd24, 27'h00000375, 5'd0, 27'h000001f3, 5'd21, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f0, 5'd11, 27'h000001ce, 5'd4, 27'h000003c9, 32'h00000400,
  1'd1,  5'd22, 27'h000003ea, 5'd10, 27'h0000029a, 5'd15, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000285, 5'd14, 27'h00000012, 5'd23, 27'h000000dc, 32'h00000400,
  1'd1,  5'd21, 27'h00000018, 5'd21, 27'h000001f1, 5'd4, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a6, 5'd23, 27'h00000325, 5'd13, 27'h000001cc, 32'h00000400,
  1'd1,  5'd21, 27'h0000012e, 5'd22, 27'h00000195, 5'd22, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000000a, 5'd0, 27'h00000238, 5'd8, 27'h000000ad, 32'h00000400,
  1'd1,  5'd3, 27'h0000011a, 5'd0, 27'h000000e4, 5'd18, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000022, 5'd0, 27'h0000008c, 5'd26, 27'h0000021f, 32'h00000400,
  1'd1,  5'd2, 27'h0000014d, 5'd13, 27'h00000201, 5'd5, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a6, 5'd12, 27'h000002e4, 5'd17, 27'h00000162, 32'h00000400,
  1'd1,  5'd0, 27'h000002f7, 5'd15, 27'h0000007b, 5'd28, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000af, 5'd23, 27'h000003d2, 5'd9, 27'h000003f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000021, 5'd25, 27'h0000023a, 5'd16, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000023e, 5'd23, 27'h00000330, 5'd26, 27'h0000023c, 32'h00000400,
  1'd1,  5'd14, 27'h00000268, 5'd4, 27'h000000d0, 5'd5, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000317, 5'd0, 27'h0000008d, 5'd16, 27'h000001cb, 32'h00000400,
  1'd1,  5'd14, 27'h0000016f, 5'd0, 27'h00000064, 5'd28, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000098, 5'd13, 27'h0000029c, 5'd5, 27'h00000246, 32'h00000400,
  1'd1,  5'd13, 27'h00000345, 5'd10, 27'h000002b0, 5'd18, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e1, 5'd12, 27'h000003ea, 5'd26, 27'h000000ff, 32'h00000400,
  1'd1,  5'd10, 27'h000003ce, 5'd21, 27'h00000155, 5'd9, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000005c, 5'd22, 27'h00000336, 5'd20, 27'h000000c9, 32'h00000400,
  1'd1,  5'd14, 27'h000001c4, 5'd24, 27'h00000332, 5'd26, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000160, 5'd4, 27'h00000111, 5'd10, 27'h0000012e, 32'h00000400,
  1'd1,  5'd23, 27'h00000239, 5'd0, 27'h00000324, 5'd17, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000256, 5'd1, 27'h00000276, 5'd28, 27'h0000027b, 32'h00000400,
  1'd1,  5'd21, 27'h00000349, 5'd11, 27'h000002d7, 5'd9, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ba, 5'd13, 27'h00000066, 5'd17, 27'h00000075, 32'h00000400,
  1'd1,  5'd21, 27'h0000031d, 5'd14, 27'h000003dc, 5'd26, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000337, 5'd20, 27'h000003f0, 5'd7, 27'h00000134, 32'h00000400,
  1'd1,  5'd22, 27'h00000026, 5'd24, 27'h000003ae, 5'd20, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d3, 5'd24, 27'h00000245, 5'd26, 27'h000003e8, 32'h00000400,
  1'd1,  5'd0, 27'h0000008b, 5'd9, 27'h0000029e, 5'd1, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000011a, 5'd9, 27'h00000383, 5'd11, 27'h00000271, 32'h00000400,
  1'd1,  5'd0, 27'h000000c7, 5'd8, 27'h00000047, 5'd25, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000011, 5'd18, 27'h000000d9, 5'd0, 27'h00000026, 32'h00000400,
  1'd1,  5'd4, 27'h00000359, 5'd19, 27'h00000391, 5'd10, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000388, 5'd17, 27'h000000c5, 5'd23, 27'h0000021d, 32'h00000400,
  1'd1,  5'd3, 27'h00000323, 5'd29, 27'h000001ce, 5'd2, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000a6, 5'd30, 27'h00000160, 5'd14, 27'h000002a9, 32'h00000400,
  1'd1,  5'd2, 27'h0000010b, 5'd28, 27'h0000005a, 5'd23, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034b, 5'd5, 27'h000001a3, 5'd4, 27'h0000003c, 32'h00000400,
  1'd1,  5'd12, 27'h0000003a, 5'd5, 27'h00000229, 5'd15, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000047, 5'd7, 27'h00000046, 5'd23, 27'h000002a8, 32'h00000400,
  1'd1,  5'd13, 27'h00000092, 5'd20, 27'h0000009a, 5'd4, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003ea, 5'd18, 27'h0000037d, 5'd14, 27'h00000017, 32'h00000400,
  1'd1,  5'd11, 27'h000003f7, 5'd18, 27'h000003fc, 5'd25, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000153, 5'd27, 27'h0000022f, 5'd4, 27'h000002e7, 32'h00000400,
  1'd1,  5'd13, 27'h00000070, 5'd30, 27'h000003b6, 5'd12, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000002a, 5'd30, 27'h000002bf, 5'd24, 27'h0000007f, 32'h00000400,
  1'd1,  5'd22, 27'h000002e7, 5'd8, 27'h000001f3, 5'd2, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000068, 5'd5, 27'h000002d0, 5'd12, 27'h00000288, 32'h00000400,
  1'd1,  5'd23, 27'h000000aa, 5'd7, 27'h000000f7, 5'd22, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bd, 5'd19, 27'h000002c5, 5'd1, 27'h000002f7, 32'h00000400,
  1'd1,  5'd21, 27'h0000009b, 5'd17, 27'h0000037b, 5'd12, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000168, 5'd16, 27'h000000bf, 5'd22, 27'h000000f1, 32'h00000400,
  1'd1,  5'd22, 27'h000002a3, 5'd26, 27'h000001d9, 5'd3, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b2, 5'd29, 27'h00000009, 5'd11, 27'h00000239, 32'h00000400,
  1'd1,  5'd25, 27'h000000c4, 5'd26, 27'h000001ad, 5'd24, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000033a, 5'd10, 27'h000000a8, 5'd9, 27'h00000172, 32'h00000400,
  1'd1,  5'd1, 27'h000001e0, 5'd5, 27'h000001cd, 5'd18, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000357, 5'd6, 27'h0000039d, 5'd29, 27'h00000368, 32'h00000400,
  1'd1,  5'd1, 27'h0000016f, 5'd20, 27'h00000026, 5'd8, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001eb, 5'd15, 27'h0000033b, 5'd17, 27'h0000007b, 32'h00000400,
  1'd1,  5'd3, 27'h00000364, 5'd19, 27'h000000e1, 5'd29, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000027e, 5'd29, 27'h00000031, 5'd7, 27'h000001c7, 32'h00000400,
  1'd1,  5'd3, 27'h00000386, 5'd30, 27'h00000053, 5'd19, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c4, 5'd29, 27'h000000b0, 5'd26, 27'h00000022, 32'h00000400,
  1'd1,  5'd12, 27'h000001a3, 5'd6, 27'h00000210, 5'd5, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000013f, 5'd7, 27'h000001b0, 5'd19, 27'h00000260, 32'h00000400,
  1'd1,  5'd12, 27'h0000026d, 5'd5, 27'h0000025d, 5'd26, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000301, 5'd19, 27'h0000000b, 5'd9, 27'h00000077, 32'h00000400,
  1'd1,  5'd11, 27'h0000002a, 5'd16, 27'h00000181, 5'd20, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000219, 5'd18, 27'h00000254, 5'd26, 27'h000000c1, 32'h00000400,
  1'd1,  5'd12, 27'h00000252, 5'd27, 27'h000001d1, 5'd5, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000151, 5'd26, 27'h00000244, 5'd16, 27'h00000189, 32'h00000400,
  1'd1,  5'd11, 27'h0000001b, 5'd26, 27'h00000144, 5'd29, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000385, 5'd5, 27'h00000252, 5'd6, 27'h00000260, 32'h00000400,
  1'd1,  5'd24, 27'h00000269, 5'd9, 27'h0000037c, 5'd17, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000c9, 5'd5, 27'h000001a9, 5'd27, 27'h00000210, 32'h00000400,
  1'd1,  5'd21, 27'h00000075, 5'd18, 27'h00000251, 5'd6, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000022c, 5'd15, 27'h000002a7, 5'd18, 27'h00000158, 32'h00000400,
  1'd1,  5'd20, 27'h0000038e, 5'd18, 27'h0000002f, 5'd29, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000189, 5'd30, 27'h000000fb, 5'd5, 27'h00000122, 32'h00000400,
  1'd1,  5'd25, 27'h000001be, 5'd26, 27'h0000030a, 5'd18, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000139, 5'd29, 27'h000001c0, 5'd30, 27'h000001f3, 32'h00000400,
  1'd1,  5'd8, 27'h0000020a, 5'd1, 27'h000002d3, 5'd8, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000144, 5'd2, 27'h000000bf, 5'd20, 27'h00000177, 32'h00000400,
  1'd1,  5'd8, 27'h00000035, 5'd4, 27'h00000166, 5'd26, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000051, 5'd13, 27'h0000020a, 5'd4, 27'h000003ca, 32'h00000400,
  1'd1,  5'd6, 27'h000002e3, 5'd12, 27'h000001ee, 5'd12, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000256, 5'd12, 27'h00000351, 5'd25, 27'h00000151, 32'h00000400,
  1'd1,  5'd7, 27'h000000ce, 5'd20, 27'h0000035c, 5'd4, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a2, 5'd23, 27'h000000c2, 5'd15, 27'h0000012c, 32'h00000400,
  1'd1,  5'd7, 27'h00000199, 5'd23, 27'h00000062, 5'd21, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a4, 5'd2, 27'h000000ca, 5'd5, 27'h000003a9, 32'h00000400,
  1'd1,  5'd15, 27'h00000271, 5'd3, 27'h0000026c, 5'd15, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000156, 5'd1, 27'h000003aa, 5'd30, 27'h0000002d, 32'h00000400,
  1'd1,  5'd18, 27'h000002d1, 5'd10, 27'h000002e4, 5'd3, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000079, 5'd15, 27'h0000011d, 5'd12, 27'h00000190, 32'h00000400,
  1'd1,  5'd18, 27'h00000348, 5'd11, 27'h00000361, 5'd24, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000061, 5'd22, 27'h000000cd, 5'd0, 27'h00000322, 32'h00000400,
  1'd1,  5'd18, 27'h0000021d, 5'd22, 27'h000000d5, 5'd11, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000324, 5'd22, 27'h00000280, 5'd25, 27'h000000e2, 32'h00000400,
  1'd1,  5'd28, 27'h000001e2, 5'd0, 27'h000000a3, 5'd3, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b7, 5'd4, 27'h000001b2, 5'd15, 27'h000000a3, 32'h00000400,
  1'd1,  5'd26, 27'h000003e2, 5'd0, 27'h00000059, 5'd24, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000316, 5'd15, 27'h0000003b, 5'd1, 27'h0000016f, 32'h00000400,
  1'd1,  5'd25, 27'h000003fc, 5'd14, 27'h000001dd, 5'd14, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d0, 5'd13, 27'h0000018e, 5'd20, 27'h000003b3, 32'h00000400,
  1'd1,  5'd29, 27'h000001b9, 5'd25, 27'h00000043, 5'd0, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000112, 5'd24, 27'h00000270, 5'd13, 27'h00000324, 32'h00000400,
  1'd1,  5'd29, 27'h00000119, 5'd23, 27'h00000170, 5'd24, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000026d, 5'd4, 27'h000000c4, 5'd2, 27'h000003de, 32'h00000400,
  1'd1,  5'd7, 27'h000001b8, 5'd4, 27'h00000378, 5'd12, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a5, 5'd5, 27'h0000000d, 5'd20, 27'h00000349, 32'h00000400,
  1'd1,  5'd6, 27'h0000026a, 5'd14, 27'h00000379, 5'd8, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000060, 5'd13, 27'h00000270, 5'd19, 27'h0000034e, 32'h00000400,
  1'd1,  5'd7, 27'h00000125, 5'd15, 27'h0000019f, 5'd28, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000030f, 5'd23, 27'h00000177, 5'd7, 27'h000001de, 32'h00000400,
  1'd1,  5'd9, 27'h000003f2, 5'd22, 27'h00000387, 5'd15, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000216, 5'd25, 27'h000001b2, 5'd29, 27'h00000223, 32'h00000400,
  1'd1,  5'd20, 27'h0000014c, 5'd4, 27'h000002ec, 5'd4, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e4, 5'd0, 27'h00000317, 5'd12, 27'h0000025f, 32'h00000400,
  1'd1,  5'd17, 27'h000003fd, 5'd3, 27'h0000034f, 5'd24, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ec, 5'd11, 27'h0000017b, 5'd9, 27'h000003e6, 32'h00000400,
  1'd1,  5'd18, 27'h000002fb, 5'd13, 27'h000002ce, 5'd16, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000276, 5'd15, 27'h000000a1, 5'd30, 27'h000003b0, 32'h00000400,
  1'd1,  5'd17, 27'h0000024a, 5'd24, 27'h000002bb, 5'd6, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000292, 5'd23, 27'h000002f6, 5'd17, 27'h00000207, 32'h00000400,
  1'd1,  5'd18, 27'h000002cb, 5'd24, 27'h0000010b, 5'd27, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e0, 5'd1, 27'h00000072, 5'd6, 27'h000003d7, 32'h00000400,
  1'd1,  5'd26, 27'h0000020b, 5'd4, 27'h000003c8, 5'd16, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000030, 5'd4, 27'h0000021a, 5'd30, 27'h000002b1, 32'h00000400,
  1'd1,  5'd29, 27'h00000330, 5'd10, 27'h000001ad, 5'd8, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001b7, 5'd13, 27'h0000010f, 5'd17, 27'h000000fb, 32'h00000400,
  1'd1,  5'd28, 27'h000002c1, 5'd14, 27'h0000002d, 5'd30, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002e4, 5'd24, 27'h00000235, 5'd7, 27'h00000383, 32'h00000400,
  1'd1,  5'd29, 27'h0000026c, 5'd21, 27'h000002ef, 5'd19, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000001c, 5'd23, 27'h0000029c, 5'd27, 27'h00000175, 32'h00000400,
  1'd1,  5'd5, 27'h0000025b, 5'd9, 27'h00000252, 5'd4, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000360, 5'd6, 27'h00000087, 5'd13, 27'h000002be, 32'h00000400,
  1'd1,  5'd8, 27'h0000034d, 5'd5, 27'h00000132, 5'd22, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000009c, 5'd18, 27'h00000056, 5'd3, 27'h000002fb, 32'h00000400,
  1'd1,  5'd8, 27'h0000028e, 5'd20, 27'h000000a2, 5'd11, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ee, 5'd16, 27'h000000b0, 5'd25, 27'h0000012a, 32'h00000400,
  1'd1,  5'd8, 27'h00000362, 5'd28, 27'h000002e4, 5'd3, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000d4, 5'd30, 27'h00000121, 5'd11, 27'h00000071, 32'h00000400,
  1'd1,  5'd5, 27'h00000211, 5'd27, 27'h00000334, 5'd23, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000026, 5'd10, 27'h00000094, 5'd4, 27'h000003e7, 32'h00000400,
  1'd1,  5'd18, 27'h00000146, 5'd9, 27'h000002f2, 5'd12, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000328, 5'd6, 27'h0000006b, 5'd21, 27'h000001b7, 32'h00000400,
  1'd1,  5'd15, 27'h00000227, 5'd20, 27'h00000106, 5'd3, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000168, 5'd17, 27'h00000254, 5'd15, 27'h0000003a, 32'h00000400,
  1'd1,  5'd17, 27'h00000327, 5'd16, 27'h000003b9, 5'd22, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000008a, 5'd29, 27'h000003fb, 5'd4, 27'h00000170, 32'h00000400,
  1'd1,  5'd16, 27'h00000372, 5'd30, 27'h000003e9, 5'd11, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002cf, 5'd28, 27'h0000027f, 5'd22, 27'h000000b0, 32'h00000400,
  1'd1,  5'd28, 27'h00000124, 5'd6, 27'h00000233, 5'd2, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000011d, 5'd10, 27'h00000096, 5'd11, 27'h0000014b, 32'h00000400,
  1'd1,  5'd29, 27'h0000032d, 5'd6, 27'h000002dc, 5'd24, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a2, 5'd18, 27'h0000032b, 5'd0, 27'h00000020, 32'h00000400,
  1'd1,  5'd26, 27'h000000c2, 5'd20, 27'h0000022c, 5'd13, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000026c, 5'd20, 27'h00000266, 5'd20, 27'h000003e0, 32'h00000400,
  1'd1,  5'd29, 27'h000001b2, 5'd27, 27'h0000010a, 5'd1, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000103, 5'd30, 27'h00000346, 5'd12, 27'h00000302, 32'h00000400,
  1'd1,  5'd30, 27'h00000282, 5'd26, 27'h000000c3, 5'd23, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c5, 5'd9, 27'h0000035c, 5'd7, 27'h00000023, 32'h00000400,
  1'd1,  5'd9, 27'h00000054, 5'd9, 27'h000002d0, 5'd17, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f6, 5'd10, 27'h00000135, 5'd26, 27'h00000023, 32'h00000400,
  1'd1,  5'd5, 27'h000001c8, 5'd19, 27'h0000028c, 5'd9, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000364, 5'd18, 27'h00000344, 5'd17, 27'h000003da, 32'h00000400,
  1'd1,  5'd10, 27'h00000042, 5'd19, 27'h00000077, 5'd28, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001c3, 5'd29, 27'h0000003c, 5'd5, 27'h00000130, 32'h00000400,
  1'd1,  5'd6, 27'h0000006f, 5'd28, 27'h0000021a, 5'd15, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a8, 5'd26, 27'h00000065, 5'd29, 27'h00000346, 32'h00000400,
  1'd1,  5'd16, 27'h000002c5, 5'd6, 27'h00000346, 5'd8, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039b, 5'd9, 27'h00000182, 5'd19, 27'h000000ca, 32'h00000400,
  1'd1,  5'd17, 27'h00000173, 5'd10, 27'h00000037, 5'd27, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000308, 5'd16, 27'h00000299, 5'd9, 27'h00000396, 32'h00000400,
  1'd1,  5'd15, 27'h00000208, 5'd17, 27'h0000018d, 5'd18, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000077, 5'd19, 27'h000001f9, 5'd27, 27'h000000a5, 32'h00000400,
  1'd1,  5'd19, 27'h00000260, 5'd28, 27'h000001ad, 5'd5, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000e9, 5'd28, 27'h0000012f, 5'd18, 27'h00000380, 32'h00000400,
  1'd1,  5'd16, 27'h0000011f, 5'd26, 27'h00000262, 5'd28, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012f, 5'd5, 27'h00000336, 5'd9, 27'h000001af, 32'h00000400,
  1'd1,  5'd26, 27'h00000380, 5'd9, 27'h00000218, 5'd18, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000277, 5'd7, 27'h00000278, 5'd28, 27'h0000038a, 32'h00000400,
  1'd1,  5'd25, 27'h00000392, 5'd18, 27'h000001e1, 5'd6, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001f, 5'd19, 27'h0000034f, 5'd20, 27'h00000059, 32'h00000400,
  1'd1,  5'd28, 27'h00000384, 5'd17, 27'h00000301, 5'd27, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000009b, 5'd27, 27'h000003f6, 5'd6, 27'h000002dd, 32'h00000400,
  1'd1,  5'd26, 27'h0000022c, 5'd28, 27'h00000018, 5'd16, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003b2, 5'd27, 27'h00000347, 5'd27, 27'h000001fd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000002bf, 5'd0, 27'h000000d9, 5'd3, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000029e, 5'd1, 27'h00000195, 5'd11, 27'h0000024d, 32'h00000400,
  1'd1,  5'd2, 27'h00000184, 5'd2, 27'h00000053, 5'd23, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000157, 5'd14, 27'h000003df, 5'd3, 27'h0000000c, 32'h00000400,
  1'd1,  5'd0, 27'h000001aa, 5'd14, 27'h000003d6, 5'd14, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000282, 5'd11, 27'h00000083, 5'd21, 27'h0000036a, 32'h00000400,
  1'd1,  5'd3, 27'h00000171, 5'd21, 27'h0000007f, 5'd3, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000013d, 5'd23, 27'h00000019, 5'd13, 27'h000003a3, 32'h00000400,
  1'd1,  5'd2, 27'h000002b8, 5'd24, 27'h00000021, 5'd22, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000016d, 5'd4, 27'h0000016a, 5'd3, 27'h000001ee, 32'h00000400,
  1'd1,  5'd15, 27'h000001a3, 5'd1, 27'h00000084, 5'd15, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000142, 5'd0, 27'h000003b7, 5'd25, 27'h000002ed, 32'h00000400,
  1'd1,  5'd15, 27'h0000009e, 5'd10, 27'h000002de, 5'd2, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001bb, 5'd12, 27'h0000033c, 5'd10, 27'h0000029f, 32'h00000400,
  1'd1,  5'd11, 27'h000001c0, 5'd11, 27'h00000075, 5'd22, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f3, 5'd24, 27'h0000026c, 5'd1, 27'h000003a6, 32'h00000400,
  1'd1,  5'd13, 27'h000000be, 5'd21, 27'h0000020a, 5'd14, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000147, 5'd24, 27'h00000218, 5'd22, 27'h0000031d, 32'h00000400,
  1'd1,  5'd24, 27'h00000098, 5'd2, 27'h00000358, 5'd0, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001a0, 5'd0, 27'h000001da, 5'd14, 27'h000000e4, 32'h00000400,
  1'd1,  5'd21, 27'h000002c6, 5'd1, 27'h0000038b, 5'd22, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000076, 5'd12, 27'h000001dd, 5'd3, 27'h000003fe, 32'h00000400,
  1'd1,  5'd21, 27'h000002b5, 5'd13, 27'h0000036d, 5'd13, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003c4, 5'd15, 27'h00000125, 5'd24, 27'h0000020f, 32'h00000400,
  1'd1,  5'd24, 27'h000003cb, 5'd22, 27'h00000197, 5'd3, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e4, 5'd21, 27'h0000020b, 5'd14, 27'h00000146, 32'h00000400,
  1'd1,  5'd20, 27'h000003fb, 5'd25, 27'h000001a5, 5'd22, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001af, 5'd1, 27'h000003e2, 5'd7, 27'h000000f5, 32'h00000400,
  1'd1,  5'd1, 27'h000001da, 5'd4, 27'h00000271, 5'd15, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c5, 5'd4, 27'h00000063, 5'd29, 27'h000001c4, 32'h00000400,
  1'd1,  5'd1, 27'h00000233, 5'd15, 27'h000000ed, 5'd6, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002dd, 5'd10, 27'h00000216, 5'd18, 27'h0000005b, 32'h00000400,
  1'd1,  5'd0, 27'h00000278, 5'd15, 27'h000001fe, 5'd29, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000a8, 5'd24, 27'h000000c6, 5'd5, 27'h000001dd, 32'h00000400,
  1'd1,  5'd1, 27'h00000177, 5'd21, 27'h000001da, 5'd20, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000235, 5'd25, 27'h00000187, 5'd29, 27'h00000268, 32'h00000400,
  1'd1,  5'd11, 27'h00000328, 5'd0, 27'h00000095, 5'd7, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003aa, 5'd2, 27'h000000f0, 5'd16, 27'h000001cd, 32'h00000400,
  1'd1,  5'd14, 27'h00000287, 5'd1, 27'h0000016a, 5'd28, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000186, 5'd11, 27'h000002a7, 5'd6, 27'h000000cd, 32'h00000400,
  1'd1,  5'd13, 27'h0000027b, 5'd11, 27'h00000338, 5'd20, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000113, 5'd10, 27'h0000029a, 5'd25, 27'h000003ad, 32'h00000400,
  1'd1,  5'd14, 27'h00000351, 5'd20, 27'h000003b2, 5'd5, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000277, 5'd22, 27'h00000399, 5'd20, 27'h0000013d, 32'h00000400,
  1'd1,  5'd15, 27'h0000019a, 5'd24, 27'h0000001d, 5'd29, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ac, 5'd2, 27'h000000aa, 5'd6, 27'h000002f9, 32'h00000400,
  1'd1,  5'd21, 27'h00000106, 5'd0, 27'h0000004b, 5'd18, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000309, 5'd2, 27'h000001ab, 5'd30, 27'h0000001e, 32'h00000400,
  1'd1,  5'd25, 27'h000002a5, 5'd11, 27'h000003f2, 5'd5, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000032, 5'd13, 27'h0000031d, 5'd16, 27'h00000207, 32'h00000400,
  1'd1,  5'd20, 27'h00000390, 5'd10, 27'h00000341, 5'd28, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003b3, 5'd23, 27'h000000c4, 5'd5, 27'h00000152, 32'h00000400,
  1'd1,  5'd24, 27'h000003a7, 5'd24, 27'h00000236, 5'd19, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002c7, 5'd21, 27'h00000267, 5'd28, 27'h000003e3, 32'h00000400,
  1'd1,  5'd1, 27'h000002d6, 5'd5, 27'h000003e8, 5'd2, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000066, 5'd9, 27'h000000f6, 5'd11, 27'h0000004d, 32'h00000400,
  1'd1,  5'd4, 27'h000002d3, 5'd6, 27'h00000358, 5'd25, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d3, 5'd15, 27'h00000283, 5'd0, 27'h0000034f, 32'h00000400,
  1'd1,  5'd2, 27'h00000041, 5'd17, 27'h0000019c, 5'd15, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000031f, 5'd17, 27'h00000359, 5'd22, 27'h00000328, 32'h00000400,
  1'd1,  5'd1, 27'h000000cf, 5'd30, 27'h00000113, 5'd3, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000004e, 5'd28, 27'h00000172, 5'd15, 27'h0000016e, 32'h00000400,
  1'd1,  5'd2, 27'h0000007f, 5'd27, 27'h0000001d, 5'd20, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001b0, 5'd5, 27'h000003d0, 5'd5, 27'h0000005e, 32'h00000400,
  1'd1,  5'd15, 27'h00000020, 5'd7, 27'h00000051, 5'd11, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000249, 5'd5, 27'h000003ab, 5'd25, 27'h000002b1, 32'h00000400,
  1'd1,  5'd13, 27'h000003ff, 5'd20, 27'h00000203, 5'd2, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000332, 5'd18, 27'h000002aa, 5'd11, 27'h00000157, 32'h00000400,
  1'd1,  5'd12, 27'h00000223, 5'd17, 27'h000002fe, 5'd25, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000310, 5'd26, 27'h000002e4, 5'd0, 27'h0000023a, 32'h00000400,
  1'd1,  5'd10, 27'h000003d4, 5'd30, 27'h00000330, 5'd10, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000119, 5'd29, 27'h0000008b, 5'd21, 27'h00000280, 32'h00000400,
  1'd1,  5'd25, 27'h00000346, 5'd10, 27'h000000b7, 5'd3, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000ad, 5'd5, 27'h00000293, 5'd14, 27'h000003e6, 32'h00000400,
  1'd1,  5'd21, 27'h000000d4, 5'd6, 27'h00000006, 5'd21, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000212, 5'd16, 27'h00000027, 5'd4, 27'h000003ea, 32'h00000400,
  1'd1,  5'd24, 27'h000003d2, 5'd16, 27'h000003ed, 5'd13, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000083, 5'd19, 27'h000002d2, 5'd21, 27'h00000205, 32'h00000400,
  1'd1,  5'd21, 27'h0000035c, 5'd27, 27'h00000117, 5'd3, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000e2, 5'd29, 27'h000003e8, 5'd13, 27'h0000021b, 32'h00000400,
  1'd1,  5'd24, 27'h000002d1, 5'd28, 27'h0000007a, 5'd20, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000274, 5'd10, 27'h00000018, 5'd7, 27'h00000047, 32'h00000400,
  1'd1,  5'd5, 27'h00000003, 5'd9, 27'h0000030d, 5'd18, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000022e, 5'd9, 27'h0000004b, 5'd27, 27'h00000231, 32'h00000400,
  1'd1,  5'd2, 27'h00000399, 5'd17, 27'h000003a3, 5'd8, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d9, 5'd19, 27'h0000022b, 5'd15, 27'h0000026d, 32'h00000400,
  1'd1,  5'd4, 27'h00000311, 5'd18, 27'h00000018, 5'd27, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003ce, 5'd30, 27'h000001e3, 5'd5, 27'h0000030e, 32'h00000400,
  1'd1,  5'd1, 27'h000002e5, 5'd30, 27'h0000039c, 5'd19, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000021a, 5'd30, 27'h0000007f, 5'd27, 27'h0000013e, 32'h00000400,
  1'd1,  5'd10, 27'h00000189, 5'd8, 27'h00000176, 5'd9, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e3, 5'd8, 27'h00000342, 5'd19, 27'h00000140, 32'h00000400,
  1'd1,  5'd13, 27'h00000036, 5'd6, 27'h000001f3, 5'd28, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000365, 5'd20, 27'h000000a7, 5'd8, 27'h000001ca, 32'h00000400,
  1'd1,  5'd12, 27'h000001b6, 5'd16, 27'h000000e4, 5'd16, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000de, 5'd15, 27'h000002d7, 5'd26, 27'h0000001d, 32'h00000400,
  1'd1,  5'd13, 27'h00000258, 5'd26, 27'h00000235, 5'd9, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000001e, 5'd29, 27'h00000064, 5'd16, 27'h000002ca, 32'h00000400,
  1'd1,  5'd10, 27'h0000039c, 5'd29, 27'h000002bd, 5'd27, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002a7, 5'd9, 27'h00000313, 5'd9, 27'h00000313, 32'h00000400,
  1'd1,  5'd20, 27'h000002d8, 5'd6, 27'h00000365, 5'd17, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002bb, 5'd10, 27'h0000011c, 5'd26, 27'h00000236, 32'h00000400,
  1'd1,  5'd25, 27'h000000fb, 5'd20, 27'h00000181, 5'd7, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000153, 5'd18, 27'h00000143, 5'd15, 27'h000003bb, 32'h00000400,
  1'd1,  5'd24, 27'h00000134, 5'd18, 27'h00000284, 5'd26, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000146, 5'd27, 27'h000001b4, 5'd9, 27'h00000332, 32'h00000400,
  1'd1,  5'd23, 27'h000000bb, 5'd26, 27'h00000166, 5'd17, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003a2, 5'd28, 27'h000002df, 5'd26, 27'h000002cd, 32'h00000400,
  1'd1,  5'd8, 27'h00000066, 5'd0, 27'h000002ec, 5'd6, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000254, 5'd2, 27'h00000395, 5'd19, 27'h000003e5, 32'h00000400,
  1'd1,  5'd9, 27'h0000023f, 5'd1, 27'h00000159, 5'd28, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000261, 5'd10, 27'h00000377, 5'd2, 27'h0000018b, 32'h00000400,
  1'd1,  5'd6, 27'h0000004b, 5'd14, 27'h0000023f, 5'd11, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000015d, 5'd11, 27'h00000003, 5'd24, 27'h000000e3, 32'h00000400,
  1'd1,  5'd8, 27'h0000014f, 5'd21, 27'h00000113, 5'd1, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000356, 5'd20, 27'h000003b4, 5'd11, 27'h0000012b, 32'h00000400,
  1'd1,  5'd7, 27'h000003ea, 5'd24, 27'h0000035c, 5'd22, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003f9, 5'd0, 27'h00000050, 5'd8, 27'h000000e5, 32'h00000400,
  1'd1,  5'd18, 27'h00000310, 5'd4, 27'h00000245, 5'd17, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b2, 5'd0, 27'h0000003c, 5'd26, 27'h00000055, 32'h00000400,
  1'd1,  5'd16, 27'h000001e5, 5'd12, 27'h0000001a, 5'd1, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000343, 5'd11, 27'h00000140, 5'd14, 27'h0000000f, 32'h00000400,
  1'd1,  5'd18, 27'h0000028c, 5'd14, 27'h00000092, 5'd24, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003f3, 5'd21, 27'h00000118, 5'd0, 27'h000002ae, 32'h00000400,
  1'd1,  5'd17, 27'h00000367, 5'd20, 27'h00000322, 5'd10, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003e7, 5'd25, 27'h000001b9, 5'd21, 27'h0000028c, 32'h00000400,
  1'd1,  5'd27, 27'h00000220, 5'd2, 27'h00000015, 5'd0, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000392, 5'd0, 27'h000003c4, 5'd11, 27'h000001c0, 32'h00000400,
  1'd1,  5'd28, 27'h000000bc, 5'd4, 27'h00000255, 5'd24, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000164, 5'd13, 27'h00000177, 5'd3, 27'h0000005c, 32'h00000400,
  1'd1,  5'd28, 27'h0000003b, 5'd11, 27'h00000217, 5'd11, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000013f, 5'd13, 27'h000000b4, 5'd21, 27'h0000000f, 32'h00000400,
  1'd1,  5'd27, 27'h0000006b, 5'd22, 27'h00000200, 5'd3, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002fb, 5'd21, 27'h00000223, 5'd10, 27'h00000374, 32'h00000400,
  1'd1,  5'd26, 27'h000002c1, 5'd23, 27'h000003c0, 5'd21, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000077, 5'd1, 27'h00000249, 5'd0, 27'h000001db, 32'h00000400,
  1'd1,  5'd7, 27'h0000023f, 5'd1, 27'h00000355, 5'd10, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001bc, 5'd3, 27'h0000029b, 5'd21, 27'h0000039e, 32'h00000400,
  1'd1,  5'd5, 27'h000000d0, 5'd12, 27'h00000352, 5'd8, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000bc, 5'd10, 27'h000001a1, 5'd16, 27'h0000005e, 32'h00000400,
  1'd1,  5'd9, 27'h0000033e, 5'd10, 27'h000001d1, 5'd27, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ae, 5'd22, 27'h0000023a, 5'd7, 27'h00000051, 32'h00000400,
  1'd1,  5'd6, 27'h0000003d, 5'd24, 27'h0000016f, 5'd20, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ad, 5'd21, 27'h000001b7, 5'd27, 27'h000000c8, 32'h00000400,
  1'd1,  5'd20, 27'h000000bf, 5'd5, 27'h00000023, 5'd2, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000283, 5'd4, 27'h00000062, 5'd11, 27'h000003b8, 32'h00000400,
  1'd1,  5'd18, 27'h00000132, 5'd1, 27'h00000203, 5'd24, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000c0, 5'd11, 27'h0000033e, 5'd9, 27'h000001c8, 32'h00000400,
  1'd1,  5'd19, 27'h0000005c, 5'd14, 27'h000002e3, 5'd15, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001cb, 5'd14, 27'h000002e4, 5'd29, 27'h00000155, 32'h00000400,
  1'd1,  5'd16, 27'h00000285, 5'd22, 27'h0000035c, 5'd5, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002fd, 5'd22, 27'h00000313, 5'd19, 27'h000000e3, 32'h00000400,
  1'd1,  5'd19, 27'h000003d0, 5'd21, 27'h00000020, 5'd29, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000020f, 5'd4, 27'h000002ae, 5'd9, 27'h000002fb, 32'h00000400,
  1'd1,  5'd29, 27'h00000032, 5'd4, 27'h00000040, 5'd17, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a0, 5'd1, 27'h00000260, 5'd26, 27'h00000358, 32'h00000400,
  1'd1,  5'd26, 27'h00000394, 5'd14, 27'h000002ec, 5'd6, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000128, 5'd15, 27'h0000002f, 5'd18, 27'h00000231, 32'h00000400,
  1'd1,  5'd28, 27'h000003aa, 5'd12, 27'h00000343, 5'd28, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e3, 5'd23, 27'h00000207, 5'd7, 27'h0000025b, 32'h00000400,
  1'd1,  5'd29, 27'h000003d3, 5'd21, 27'h00000011, 5'd17, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006a, 5'd22, 27'h00000089, 5'd27, 27'h000002ea, 32'h00000400,
  1'd1,  5'd5, 27'h00000320, 5'd6, 27'h00000365, 5'd0, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002b9, 5'd8, 27'h000001be, 5'd12, 27'h000002ec, 32'h00000400,
  1'd1,  5'd8, 27'h000003e3, 5'd6, 27'h0000002d, 5'd22, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002fe, 5'd19, 27'h0000022c, 5'd1, 27'h000003d9, 32'h00000400,
  1'd1,  5'd6, 27'h00000182, 5'd20, 27'h00000127, 5'd12, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000026d, 5'd18, 27'h00000329, 5'd24, 27'h0000006d, 32'h00000400,
  1'd1,  5'd9, 27'h00000113, 5'd30, 27'h00000340, 5'd1, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000092, 5'd28, 27'h000001be, 5'd11, 27'h00000340, 32'h00000400,
  1'd1,  5'd7, 27'h00000308, 5'd29, 27'h000001d6, 5'd23, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000021f, 5'd6, 27'h000002b0, 5'd1, 27'h000003cd, 32'h00000400,
  1'd1,  5'd19, 27'h000001c0, 5'd8, 27'h00000125, 5'd12, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000019d, 5'd9, 27'h0000023c, 5'd23, 27'h000002f3, 32'h00000400,
  1'd1,  5'd17, 27'h00000232, 5'd18, 27'h0000032d, 5'd4, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000081, 5'd15, 27'h000002ed, 5'd14, 27'h0000035e, 32'h00000400,
  1'd1,  5'd18, 27'h00000113, 5'd20, 27'h0000013f, 5'd25, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000250, 5'd30, 27'h00000345, 5'd2, 27'h00000007, 32'h00000400,
  1'd1,  5'd18, 27'h0000022a, 5'd28, 27'h000003f6, 5'd11, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f9, 5'd26, 27'h000002c6, 5'd24, 27'h00000168, 32'h00000400,
  1'd1,  5'd29, 27'h0000030a, 5'd9, 27'h000003fd, 5'd2, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000fe, 5'd8, 27'h000002e8, 5'd14, 27'h00000292, 32'h00000400,
  1'd1,  5'd26, 27'h0000036f, 5'd9, 27'h000002db, 5'd23, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000224, 5'd19, 27'h00000242, 5'd4, 27'h00000067, 32'h00000400,
  1'd1,  5'd26, 27'h000001d7, 5'd16, 27'h00000013, 5'd10, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012f, 5'd15, 27'h00000313, 5'd24, 27'h0000019e, 32'h00000400,
  1'd1,  5'd28, 27'h00000241, 5'd28, 27'h00000207, 5'd1, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000175, 5'd28, 27'h00000291, 5'd12, 27'h0000009e, 32'h00000400,
  1'd1,  5'd27, 27'h0000024e, 5'd28, 27'h0000028e, 5'd21, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000367, 5'd9, 27'h000003a0, 5'd10, 27'h00000082, 32'h00000400,
  1'd1,  5'd5, 27'h0000031e, 5'd5, 27'h0000026f, 5'd16, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000025f, 5'd5, 27'h00000184, 5'd30, 27'h00000316, 32'h00000400,
  1'd1,  5'd6, 27'h000002a7, 5'd17, 27'h0000011a, 5'd5, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000056, 5'd18, 27'h000000f5, 5'd19, 27'h00000201, 32'h00000400,
  1'd1,  5'd7, 27'h00000157, 5'd20, 27'h0000026e, 5'd27, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001f0, 5'd27, 27'h00000240, 5'd5, 27'h000000d5, 32'h00000400,
  1'd1,  5'd5, 27'h000000d5, 5'd26, 27'h0000032b, 5'd19, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000242, 5'd29, 27'h0000034f, 5'd27, 27'h000002b0, 32'h00000400,
  1'd1,  5'd16, 27'h00000317, 5'd9, 27'h0000009d, 5'd6, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000167, 5'd8, 27'h0000029b, 5'd18, 27'h0000019f, 32'h00000400,
  1'd1,  5'd20, 27'h00000161, 5'd7, 27'h00000101, 5'd30, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000261, 5'd19, 27'h000001d5, 5'd8, 27'h0000001d, 32'h00000400,
  1'd1,  5'd19, 27'h000001a5, 5'd18, 27'h00000066, 5'd16, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000032c, 5'd19, 27'h000002d4, 5'd29, 27'h00000065, 32'h00000400,
  1'd1,  5'd19, 27'h000002f5, 5'd28, 27'h0000037a, 5'd7, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000261, 5'd28, 27'h000001ed, 5'd17, 27'h0000006c, 32'h00000400,
  1'd1,  5'd16, 27'h0000001e, 5'd28, 27'h000001d0, 5'd27, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000025c, 5'd8, 27'h000002d6, 5'd6, 27'h000000e7, 32'h00000400,
  1'd1,  5'd26, 27'h00000052, 5'd7, 27'h000001af, 5'd17, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000229, 5'd5, 27'h00000311, 5'd26, 27'h00000043, 32'h00000400,
  1'd1,  5'd30, 27'h00000159, 5'd16, 27'h0000024d, 5'd5, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000019c, 5'd18, 27'h000003d1, 5'd20, 27'h0000029b, 32'h00000400,
  1'd1,  5'd28, 27'h000002b2, 5'd16, 27'h00000281, 5'd27, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c7, 5'd27, 27'h00000311, 5'd6, 27'h0000014b, 32'h00000400,
  1'd1,  5'd30, 27'h00000033, 5'd30, 27'h000001a0, 5'd19, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000108, 5'd26, 27'h00000193, 5'd27, 27'h0000021d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000128, 5'd3, 27'h000003f5, 5'd3, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000029c, 5'd1, 27'h0000018a, 5'd11, 27'h000002b2, 32'h00000400,
  1'd1,  5'd2, 27'h0000010a, 5'd0, 27'h0000037f, 5'd21, 27'h00000257, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000211, 5'd11, 27'h00000264, 5'd2, 27'h000000e8, 32'h00000400,
  1'd1,  5'd0, 27'h00000253, 5'd14, 27'h0000013a, 5'd12, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000081, 5'd12, 27'h0000038e, 5'd24, 27'h00000231, 32'h00000400,
  1'd1,  5'd0, 27'h0000026b, 5'd21, 27'h00000172, 5'd4, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e8, 5'd22, 27'h00000118, 5'd13, 27'h00000303, 32'h00000400,
  1'd1,  5'd2, 27'h0000027c, 5'd23, 27'h000002ff, 5'd23, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000206, 5'd4, 27'h0000000e, 5'd2, 27'h00000078, 32'h00000400,
  1'd1,  5'd12, 27'h00000343, 5'd1, 27'h000001d7, 5'd14, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000241, 5'd0, 27'h00000274, 5'd24, 27'h0000013e, 32'h00000400,
  1'd1,  5'd13, 27'h0000008f, 5'd13, 27'h0000016a, 5'd1, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000006c, 5'd11, 27'h00000068, 5'd14, 27'h00000299, 32'h00000400,
  1'd1,  5'd12, 27'h0000033e, 5'd14, 27'h00000187, 5'd24, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000135, 5'd25, 27'h000000cb, 5'd2, 27'h000002b0, 32'h00000400,
  1'd1,  5'd11, 27'h000001eb, 5'd23, 27'h0000030e, 5'd12, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000001d, 5'd24, 27'h000001cd, 5'd23, 27'h00000256, 32'h00000400,
  1'd1,  5'd21, 27'h00000258, 5'd0, 27'h0000021b, 5'd4, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002f4, 5'd2, 27'h00000379, 5'd13, 27'h00000221, 32'h00000400,
  1'd1,  5'd24, 27'h00000001, 5'd3, 27'h00000061, 5'd20, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000017a, 5'd12, 27'h00000266, 5'd1, 27'h00000180, 32'h00000400,
  1'd1,  5'd22, 27'h000001b4, 5'd15, 27'h00000077, 5'd11, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001dd, 5'd12, 27'h0000008f, 5'd23, 27'h00000184, 32'h00000400,
  1'd1,  5'd21, 27'h000000da, 5'd21, 27'h00000346, 5'd3, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000096, 5'd25, 27'h000000d1, 5'd12, 27'h00000196, 32'h00000400,
  1'd1,  5'd21, 27'h00000377, 5'd22, 27'h00000226, 5'd24, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b2, 5'd0, 27'h00000165, 5'd8, 27'h000002c6, 32'h00000400,
  1'd1,  5'd4, 27'h00000358, 5'd3, 27'h000000af, 5'd17, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000e4, 5'd4, 27'h00000140, 5'd30, 27'h00000263, 32'h00000400,
  1'd1,  5'd4, 27'h0000024d, 5'd11, 27'h00000100, 5'd6, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001da, 5'd12, 27'h00000186, 5'd19, 27'h00000387, 32'h00000400,
  1'd1,  5'd3, 27'h000002cc, 5'd12, 27'h00000349, 5'd28, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000092, 5'd24, 27'h00000132, 5'd6, 27'h000000a8, 32'h00000400,
  1'd1,  5'd2, 27'h000001cc, 5'd21, 27'h0000005e, 5'd15, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a4, 5'd20, 27'h00000374, 5'd30, 27'h00000326, 32'h00000400,
  1'd1,  5'd11, 27'h0000016f, 5'd2, 27'h00000027, 5'd8, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000174, 5'd2, 27'h00000309, 5'd16, 27'h00000359, 32'h00000400,
  1'd1,  5'd14, 27'h000000ee, 5'd2, 27'h0000028f, 5'd28, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000010b, 5'd14, 27'h0000018a, 5'd6, 27'h000000c6, 32'h00000400,
  1'd1,  5'd10, 27'h000003d8, 5'd15, 27'h0000003a, 5'd19, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000063, 5'd12, 27'h0000025a, 5'd27, 27'h0000030f, 32'h00000400,
  1'd1,  5'd12, 27'h000001d4, 5'd21, 27'h00000267, 5'd9, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000028b, 5'd24, 27'h000001a5, 5'd15, 27'h000003c3, 32'h00000400,
  1'd1,  5'd10, 27'h000001dc, 5'd25, 27'h00000178, 5'd29, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002a0, 5'd2, 27'h000002ee, 5'd10, 27'h00000107, 32'h00000400,
  1'd1,  5'd23, 27'h00000339, 5'd4, 27'h00000185, 5'd18, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000030f, 5'd3, 27'h00000210, 5'd29, 27'h000003d4, 32'h00000400,
  1'd1,  5'd25, 27'h000002f1, 5'd12, 27'h000002c7, 5'd7, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000062, 5'd14, 27'h000003ee, 5'd20, 27'h00000281, 32'h00000400,
  1'd1,  5'd23, 27'h000002a6, 5'd12, 27'h00000385, 5'd29, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000035a, 5'd23, 27'h000001c4, 5'd9, 27'h000000bf, 32'h00000400,
  1'd1,  5'd20, 27'h000002d0, 5'd23, 27'h00000113, 5'd20, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000110, 5'd22, 27'h0000026c, 5'd28, 27'h000000b3, 32'h00000400,
  1'd1,  5'd0, 27'h000002ad, 5'd6, 27'h00000131, 5'd4, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000023, 5'd5, 27'h00000366, 5'd13, 27'h0000035c, 32'h00000400,
  1'd1,  5'd2, 27'h00000300, 5'd7, 27'h0000027f, 5'd23, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000314, 5'd16, 27'h000003a1, 5'd4, 27'h0000003f, 32'h00000400,
  1'd1,  5'd5, 27'h00000027, 5'd17, 27'h00000338, 5'd13, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000f0, 5'd20, 27'h0000020f, 5'd23, 27'h00000272, 32'h00000400,
  1'd1,  5'd3, 27'h0000030d, 5'd30, 27'h0000025c, 5'd4, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f1, 5'd29, 27'h000000b7, 5'd14, 27'h00000321, 32'h00000400,
  1'd1,  5'd4, 27'h00000128, 5'd27, 27'h00000243, 5'd25, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001d0, 5'd7, 27'h0000030b, 5'd3, 27'h0000039a, 32'h00000400,
  1'd1,  5'd12, 27'h0000015e, 5'd7, 27'h0000018a, 5'd12, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000015b, 5'd5, 27'h000002fd, 5'd21, 27'h00000331, 32'h00000400,
  1'd1,  5'd10, 27'h00000357, 5'd20, 27'h00000144, 5'd0, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002a1, 5'd17, 27'h0000021f, 5'd13, 27'h000000e2, 32'h00000400,
  1'd1,  5'd12, 27'h000000ae, 5'd17, 27'h00000097, 5'd22, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000022b, 5'd26, 27'h0000023c, 5'd1, 27'h00000091, 32'h00000400,
  1'd1,  5'd12, 27'h00000223, 5'd29, 27'h000002df, 5'd14, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f5, 5'd26, 27'h0000035f, 5'd21, 27'h000003f6, 32'h00000400,
  1'd1,  5'd23, 27'h0000023d, 5'd7, 27'h00000374, 5'd2, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000183, 5'd6, 27'h000003b4, 5'd11, 27'h000001a5, 32'h00000400,
  1'd1,  5'd24, 27'h000000ff, 5'd6, 27'h0000018a, 5'd21, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034d, 5'd16, 27'h000000ee, 5'd4, 27'h000003ef, 32'h00000400,
  1'd1,  5'd23, 27'h0000020c, 5'd19, 27'h00000204, 5'd10, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000031, 5'd16, 27'h000001fe, 5'd22, 27'h000003e4, 32'h00000400,
  1'd1,  5'd23, 27'h000003d4, 5'd25, 27'h000003ba, 5'd3, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f1, 5'd27, 27'h000001b7, 5'd10, 27'h00000227, 32'h00000400,
  1'd1,  5'd20, 27'h000003b8, 5'd26, 27'h00000115, 5'd24, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000011e, 5'd6, 27'h00000125, 5'd5, 27'h000002fb, 32'h00000400,
  1'd1,  5'd2, 27'h00000068, 5'd8, 27'h0000006a, 5'd18, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000006c, 5'd7, 27'h00000259, 5'd28, 27'h000002e6, 32'h00000400,
  1'd1,  5'd4, 27'h0000002b, 5'd16, 27'h00000371, 5'd9, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000062, 5'd15, 27'h00000228, 5'd20, 27'h000000a9, 32'h00000400,
  1'd1,  5'd2, 27'h000000ba, 5'd18, 27'h0000035b, 5'd26, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000385, 5'd29, 27'h00000268, 5'd7, 27'h000000e4, 32'h00000400,
  1'd1,  5'd3, 27'h000001bf, 5'd27, 27'h000001f7, 5'd15, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000f9, 5'd29, 27'h000000b7, 5'd30, 27'h0000029e, 32'h00000400,
  1'd1,  5'd14, 27'h0000014c, 5'd6, 27'h0000011e, 5'd7, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000027, 5'd9, 27'h0000030b, 5'd17, 27'h000002f7, 32'h00000400,
  1'd1,  5'd14, 27'h000002b5, 5'd9, 27'h0000035a, 5'd30, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000277, 5'd18, 27'h000000fe, 5'd7, 27'h000002ed, 32'h00000400,
  1'd1,  5'd14, 27'h00000170, 5'd20, 27'h00000212, 5'd17, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a1, 5'd18, 27'h00000376, 5'd27, 27'h000002f1, 32'h00000400,
  1'd1,  5'd14, 27'h00000312, 5'd26, 27'h000001c1, 5'd7, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000012f, 5'd26, 27'h000003b9, 5'd16, 27'h00000332, 32'h00000400,
  1'd1,  5'd12, 27'h0000017c, 5'd30, 27'h00000045, 5'd27, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000118, 5'd8, 27'h000002f0, 5'd7, 27'h000002e2, 32'h00000400,
  1'd1,  5'd23, 27'h00000172, 5'd5, 27'h00000388, 5'd17, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000350, 5'd7, 27'h00000278, 5'd29, 27'h000001e9, 32'h00000400,
  1'd1,  5'd23, 27'h0000007d, 5'd17, 27'h0000012a, 5'd8, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002aa, 5'd20, 27'h000000dd, 5'd19, 27'h00000248, 32'h00000400,
  1'd1,  5'd23, 27'h000000d1, 5'd17, 27'h00000025, 5'd27, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000006b, 5'd26, 27'h00000377, 5'd5, 27'h000001d3, 32'h00000400,
  1'd1,  5'd22, 27'h00000275, 5'd30, 27'h00000270, 5'd18, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002fa, 5'd27, 27'h000001c3, 5'd28, 27'h000000bc, 32'h00000400,
  1'd1,  5'd5, 27'h00000309, 5'd3, 27'h00000007, 5'd5, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002ee, 5'd0, 27'h000001d5, 5'd18, 27'h00000294, 32'h00000400,
  1'd1,  5'd6, 27'h0000018d, 5'd4, 27'h000000cd, 5'd26, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e5, 5'd14, 27'h000000e1, 5'd4, 27'h00000176, 32'h00000400,
  1'd1,  5'd9, 27'h00000186, 5'd10, 27'h00000372, 5'd12, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e1, 5'd10, 27'h0000027c, 5'd23, 27'h0000035f, 32'h00000400,
  1'd1,  5'd7, 27'h000003fa, 5'd22, 27'h00000268, 5'd4, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a0, 5'd21, 27'h00000218, 5'd14, 27'h0000019e, 32'h00000400,
  1'd1,  5'd5, 27'h0000012d, 5'd22, 27'h000001dc, 5'd25, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001db, 5'd1, 27'h0000010e, 5'd8, 27'h00000372, 32'h00000400,
  1'd1,  5'd17, 27'h00000235, 5'd4, 27'h000002f4, 5'd18, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000109, 5'd4, 27'h0000017e, 5'd26, 27'h0000014a, 32'h00000400,
  1'd1,  5'd18, 27'h000001a7, 5'd10, 27'h000003ee, 5'd2, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006f, 5'd13, 27'h000001ee, 5'd14, 27'h000003f4, 32'h00000400,
  1'd1,  5'd16, 27'h0000038c, 5'd15, 27'h000000f4, 5'd22, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000c8, 5'd24, 27'h0000012b, 5'd2, 27'h000000e4, 32'h00000400,
  1'd1,  5'd20, 27'h0000026a, 5'd22, 27'h00000199, 5'd15, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000015d, 5'd21, 27'h00000071, 5'd24, 27'h00000064, 32'h00000400,
  1'd1,  5'd26, 27'h00000007, 5'd4, 27'h000003c5, 5'd3, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000085, 5'd4, 27'h00000306, 5'd12, 27'h000002b2, 32'h00000400,
  1'd1,  5'd30, 27'h000002bd, 5'd2, 27'h0000001e, 5'd22, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000002, 5'd12, 27'h00000154, 5'd3, 27'h0000031a, 32'h00000400,
  1'd1,  5'd28, 27'h00000104, 5'd13, 27'h000002fa, 5'd15, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000016b, 5'd14, 27'h000000d0, 5'd22, 27'h00000329, 32'h00000400,
  1'd1,  5'd30, 27'h000000af, 5'd24, 27'h00000076, 5'd1, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000242, 5'd25, 27'h000000fb, 5'd13, 27'h000002ea, 32'h00000400,
  1'd1,  5'd29, 27'h000002bf, 5'd23, 27'h000001fe, 5'd22, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d4, 5'd0, 27'h00000022, 5'd1, 27'h000002f2, 32'h00000400,
  1'd1,  5'd6, 27'h00000187, 5'd0, 27'h00000306, 5'd13, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000019c, 5'd3, 27'h00000001, 5'd22, 27'h000003b2, 32'h00000400,
  1'd1,  5'd9, 27'h0000004b, 5'd10, 27'h000001ea, 5'd6, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000093, 5'd14, 27'h00000120, 5'd19, 27'h000001cc, 32'h00000400,
  1'd1,  5'd8, 27'h000002e4, 5'd11, 27'h000000fd, 5'd30, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e2, 5'd23, 27'h00000272, 5'd6, 27'h00000149, 32'h00000400,
  1'd1,  5'd10, 27'h00000151, 5'd25, 27'h00000256, 5'd17, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e6, 5'd25, 27'h0000024f, 5'd26, 27'h00000206, 32'h00000400,
  1'd1,  5'd20, 27'h00000217, 5'd1, 27'h00000242, 5'd1, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000118, 5'd0, 27'h000003c8, 5'd12, 27'h00000081, 32'h00000400,
  1'd1,  5'd16, 27'h000003f5, 5'd2, 27'h000002f0, 5'd24, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000321, 5'd13, 27'h00000185, 5'd10, 27'h0000010c, 32'h00000400,
  1'd1,  5'd18, 27'h000001fa, 5'd11, 27'h00000201, 5'd20, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000016f, 5'd11, 27'h00000275, 5'd28, 27'h000001c2, 32'h00000400,
  1'd1,  5'd19, 27'h00000239, 5'd22, 27'h00000292, 5'd9, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000dc, 5'd22, 27'h00000314, 5'd15, 27'h0000034e, 32'h00000400,
  1'd1,  5'd16, 27'h0000001e, 5'd21, 27'h0000016a, 5'd30, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000390, 5'd4, 27'h0000016b, 5'd5, 27'h000002e7, 32'h00000400,
  1'd1,  5'd28, 27'h000002b9, 5'd4, 27'h000001c3, 5'd15, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000236, 5'd1, 27'h000000a6, 5'd27, 27'h00000150, 32'h00000400,
  1'd1,  5'd29, 27'h00000186, 5'd12, 27'h000000ec, 5'd9, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003cd, 5'd14, 27'h00000157, 5'd19, 27'h0000010f, 32'h00000400,
  1'd1,  5'd30, 27'h00000100, 5'd14, 27'h00000144, 5'd28, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000134, 5'd22, 27'h000000a4, 5'd8, 27'h0000006f, 32'h00000400,
  1'd1,  5'd26, 27'h00000097, 5'd25, 27'h000001b0, 5'd16, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c2, 5'd21, 27'h00000109, 5'd27, 27'h000003ee, 32'h00000400,
  1'd1,  5'd7, 27'h00000308, 5'd8, 27'h0000033e, 5'd4, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000357, 5'd6, 27'h0000022f, 5'd12, 27'h0000018d, 32'h00000400,
  1'd1,  5'd5, 27'h00000349, 5'd5, 27'h000001b4, 5'd23, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000266, 5'd16, 27'h00000141, 5'd3, 27'h000000c7, 32'h00000400,
  1'd1,  5'd10, 27'h0000005d, 5'd17, 27'h00000041, 5'd14, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000010c, 5'd18, 27'h000003e3, 5'd25, 27'h0000006a, 32'h00000400,
  1'd1,  5'd6, 27'h000001db, 5'd29, 27'h00000044, 5'd4, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e6, 5'd29, 27'h000002af, 5'd12, 27'h0000003f, 32'h00000400,
  1'd1,  5'd5, 27'h000003da, 5'd26, 27'h0000019e, 5'd21, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000110, 5'd5, 27'h00000227, 5'd1, 27'h000000bf, 32'h00000400,
  1'd1,  5'd20, 27'h00000020, 5'd7, 27'h000000eb, 5'd12, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000136, 5'd5, 27'h00000150, 5'd21, 27'h000000c6, 32'h00000400,
  1'd1,  5'd15, 27'h0000035b, 5'd19, 27'h00000274, 5'd2, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000022d, 5'd20, 27'h000001c1, 5'd14, 27'h000002c8, 32'h00000400,
  1'd1,  5'd16, 27'h000003b1, 5'd20, 27'h000000b8, 5'd21, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000321, 5'd30, 27'h00000330, 5'd2, 27'h00000093, 32'h00000400,
  1'd1,  5'd16, 27'h000000c3, 5'd30, 27'h00000390, 5'd10, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000318, 5'd28, 27'h00000175, 5'd21, 27'h000003cb, 32'h00000400,
  1'd1,  5'd26, 27'h00000138, 5'd5, 27'h000000f8, 5'd3, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000b0, 5'd6, 27'h000002e0, 5'd11, 27'h0000029d, 32'h00000400,
  1'd1,  5'd25, 27'h00000385, 5'd6, 27'h00000239, 5'd23, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003bb, 5'd16, 27'h000000d8, 5'd0, 27'h0000003a, 32'h00000400,
  1'd1,  5'd26, 27'h000002bd, 5'd19, 27'h000000bd, 5'd15, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000264, 5'd18, 27'h00000381, 5'd25, 27'h00000156, 32'h00000400,
  1'd1,  5'd27, 27'h00000221, 5'd26, 27'h0000001c, 5'd1, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001da, 5'd27, 27'h000001a6, 5'd12, 27'h0000008d, 32'h00000400,
  1'd1,  5'd29, 27'h0000014b, 5'd27, 27'h000000d3, 5'd25, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000185, 5'd9, 27'h00000134, 5'd5, 27'h000003a9, 32'h00000400,
  1'd1,  5'd8, 27'h00000118, 5'd6, 27'h0000013b, 5'd18, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000249, 5'd8, 27'h0000006c, 5'd27, 27'h000000f5, 32'h00000400,
  1'd1,  5'd6, 27'h00000322, 5'd20, 27'h000000d0, 5'd6, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000001f, 5'd17, 27'h00000290, 5'd17, 27'h000003bd, 32'h00000400,
  1'd1,  5'd8, 27'h000003b6, 5'd17, 27'h000003a0, 5'd29, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000000f, 5'd25, 27'h000003b5, 5'd9, 27'h00000272, 32'h00000400,
  1'd1,  5'd8, 27'h00000053, 5'd26, 27'h0000012a, 5'd16, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002d6, 5'd30, 27'h0000010f, 5'd30, 27'h0000023c, 32'h00000400,
  1'd1,  5'd17, 27'h000002ea, 5'd5, 27'h00000254, 5'd5, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000271, 5'd9, 27'h0000031a, 5'd18, 27'h000003f5, 32'h00000400,
  1'd1,  5'd16, 27'h00000125, 5'd5, 27'h000002f0, 5'd28, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000009d, 5'd20, 27'h0000028c, 5'd6, 27'h000001cf, 32'h00000400,
  1'd1,  5'd20, 27'h00000209, 5'd20, 27'h0000025f, 5'd15, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000d4, 5'd17, 27'h00000157, 5'd30, 27'h000002da, 32'h00000400,
  1'd1,  5'd15, 27'h000003a8, 5'd28, 27'h000001d5, 5'd5, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000036a, 5'd28, 27'h000002e4, 5'd19, 27'h00000379, 32'h00000400,
  1'd1,  5'd17, 27'h00000351, 5'd29, 27'h000003e3, 5'd28, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d0, 5'd5, 27'h0000038e, 5'd9, 27'h00000218, 32'h00000400,
  1'd1,  5'd25, 27'h000003c9, 5'd9, 27'h0000037c, 5'd16, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000010a, 5'd9, 27'h00000288, 5'd29, 27'h00000064, 32'h00000400,
  1'd1,  5'd30, 27'h00000319, 5'd19, 27'h00000260, 5'd8, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000180, 5'd17, 27'h00000261, 5'd17, 27'h000001ac, 32'h00000400,
  1'd1,  5'd27, 27'h00000297, 5'd16, 27'h000002cb, 5'd29, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ed, 5'd29, 27'h00000334, 5'd8, 27'h00000115, 32'h00000400,
  1'd1,  5'd29, 27'h00000021, 5'd29, 27'h00000340, 5'd17, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000354, 5'd27, 27'h00000358, 5'd29, 27'h000002f5, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000000ef, 5'd1, 27'h00000328, 5'd1, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000330, 5'd4, 27'h000003eb, 5'd11, 27'h000001a6, 32'h00000400,
  1'd1,  5'd1, 27'h000000b9, 5'd3, 27'h000003d4, 5'd23, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000dc, 5'd14, 27'h00000208, 5'd2, 27'h00000113, 32'h00000400,
  1'd1,  5'd0, 27'h00000028, 5'd12, 27'h00000177, 5'd15, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000047, 5'd10, 27'h000001c4, 5'd22, 27'h000002d9, 32'h00000400,
  1'd1,  5'd4, 27'h00000029, 5'd22, 27'h00000290, 5'd0, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023a, 5'd25, 27'h0000022d, 5'd14, 27'h00000041, 32'h00000400,
  1'd1,  5'd4, 27'h000002a7, 5'd23, 27'h00000302, 5'd25, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021f, 5'd3, 27'h000002ec, 5'd0, 27'h0000010b, 32'h00000400,
  1'd1,  5'd11, 27'h000002f4, 5'd3, 27'h00000078, 5'd13, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000021e, 5'd3, 27'h0000028e, 5'd22, 27'h0000006c, 32'h00000400,
  1'd1,  5'd12, 27'h00000183, 5'd14, 27'h000002dd, 5'd5, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d2, 5'd14, 27'h0000012b, 5'd14, 27'h00000241, 32'h00000400,
  1'd1,  5'd14, 27'h00000268, 5'd10, 27'h0000028c, 5'd22, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000002c, 5'd23, 27'h0000021b, 5'd0, 27'h000000fd, 32'h00000400,
  1'd1,  5'd11, 27'h000001c7, 5'd24, 27'h0000012c, 5'd13, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000054, 5'd21, 27'h00000075, 5'd25, 27'h000000ac, 32'h00000400,
  1'd1,  5'd23, 27'h0000018d, 5'd4, 27'h000002e0, 5'd2, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001f7, 5'd1, 27'h00000372, 5'd14, 27'h0000037c, 32'h00000400,
  1'd1,  5'd21, 27'h00000129, 5'd1, 27'h00000054, 5'd25, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a1, 5'd10, 27'h00000192, 5'd4, 27'h00000394, 32'h00000400,
  1'd1,  5'd22, 27'h000003a6, 5'd12, 27'h0000028c, 5'd12, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002ff, 5'd11, 27'h0000010e, 5'd20, 27'h0000030c, 32'h00000400,
  1'd1,  5'd24, 27'h00000077, 5'd25, 27'h00000064, 5'd4, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000042, 5'd25, 27'h000002f0, 5'd12, 27'h00000194, 32'h00000400,
  1'd1,  5'd25, 27'h000001a6, 5'd23, 27'h000000a5, 5'd25, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028b, 5'd3, 27'h000001c7, 5'd7, 27'h00000005, 32'h00000400,
  1'd1,  5'd2, 27'h00000005, 5'd2, 27'h000002b7, 5'd18, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003be, 5'd2, 27'h00000212, 5'd26, 27'h0000014c, 32'h00000400,
  1'd1,  5'd1, 27'h0000018b, 5'd14, 27'h000000c7, 5'd5, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000201, 5'd13, 27'h0000028d, 5'd18, 27'h000002dc, 32'h00000400,
  1'd1,  5'd3, 27'h00000084, 5'd11, 27'h0000012c, 5'd29, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d4, 5'd23, 27'h00000339, 5'd9, 27'h000003b5, 32'h00000400,
  1'd1,  5'd3, 27'h00000104, 5'd22, 27'h0000015a, 5'd16, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001dc, 5'd24, 27'h00000365, 5'd27, 27'h000002f4, 32'h00000400,
  1'd1,  5'd12, 27'h0000031c, 5'd2, 27'h0000032c, 5'd5, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d9, 5'd2, 27'h000000d7, 5'd16, 27'h00000221, 32'h00000400,
  1'd1,  5'd14, 27'h00000016, 5'd0, 27'h00000114, 5'd30, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000351, 5'd14, 27'h00000314, 5'd9, 27'h000001c4, 32'h00000400,
  1'd1,  5'd13, 27'h0000034e, 5'd12, 27'h0000019a, 5'd19, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034f, 5'd11, 27'h000002f8, 5'd28, 27'h00000157, 32'h00000400,
  1'd1,  5'd10, 27'h00000330, 5'd25, 27'h000001a5, 5'd10, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000029, 5'd23, 27'h000002ea, 5'd19, 27'h0000025d, 32'h00000400,
  1'd1,  5'd10, 27'h00000391, 5'd22, 27'h000000ad, 5'd29, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000088, 5'd4, 27'h00000103, 5'd6, 27'h000003c9, 32'h00000400,
  1'd1,  5'd24, 27'h00000021, 5'd2, 27'h0000039a, 5'd19, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000029c, 5'd0, 27'h00000359, 5'd28, 27'h00000113, 32'h00000400,
  1'd1,  5'd25, 27'h000000f4, 5'd14, 27'h000001ca, 5'd8, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003cd, 5'd14, 27'h00000318, 5'd17, 27'h0000020f, 32'h00000400,
  1'd1,  5'd24, 27'h00000204, 5'd10, 27'h000002f8, 5'd26, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a2, 5'd23, 27'h00000252, 5'd5, 27'h000002e2, 32'h00000400,
  1'd1,  5'd25, 27'h0000002f, 5'd24, 27'h000001b2, 5'd19, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000227, 5'd23, 27'h0000014e, 5'd30, 27'h000003f2, 32'h00000400,
  1'd1,  5'd0, 27'h0000035c, 5'd6, 27'h000003a4, 5'd1, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000118, 5'd8, 27'h0000008f, 5'd12, 27'h000002c1, 32'h00000400,
  1'd1,  5'd2, 27'h000001e5, 5'd7, 27'h00000078, 5'd21, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000096, 5'd20, 27'h000000e2, 5'd4, 27'h000003e3, 32'h00000400,
  1'd1,  5'd4, 27'h000001de, 5'd16, 27'h000001c4, 5'd14, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000116, 5'd17, 27'h00000029, 5'd23, 27'h00000097, 32'h00000400,
  1'd1,  5'd2, 27'h00000234, 5'd27, 27'h0000038c, 5'd4, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000138, 5'd26, 27'h00000002, 5'd11, 27'h00000269, 32'h00000400,
  1'd1,  5'd4, 27'h00000312, 5'd27, 27'h000000fc, 5'd21, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000033d, 5'd5, 27'h00000327, 5'd1, 27'h000003e8, 32'h00000400,
  1'd1,  5'd10, 27'h00000229, 5'd9, 27'h000000c0, 5'd10, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e9, 5'd7, 27'h0000032f, 5'd22, 27'h000000a1, 32'h00000400,
  1'd1,  5'd12, 27'h00000379, 5'd19, 27'h00000307, 5'd4, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000022, 5'd16, 27'h00000119, 5'd12, 27'h000000ff, 32'h00000400,
  1'd1,  5'd14, 27'h00000387, 5'd19, 27'h000000f3, 5'd21, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003cd, 5'd26, 27'h0000035f, 5'd2, 27'h0000013c, 32'h00000400,
  1'd1,  5'd11, 27'h000003ed, 5'd26, 27'h000001ec, 5'd15, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029e, 5'd27, 27'h0000023a, 5'd25, 27'h0000024a, 32'h00000400,
  1'd1,  5'd22, 27'h000001ac, 5'd9, 27'h000003cd, 5'd2, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fa, 5'd8, 27'h000003b8, 5'd14, 27'h00000337, 32'h00000400,
  1'd1,  5'd21, 27'h0000015d, 5'd8, 27'h000000d0, 5'd22, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003c2, 5'd20, 27'h000001c4, 5'd3, 27'h00000171, 32'h00000400,
  1'd1,  5'd25, 27'h00000140, 5'd19, 27'h00000020, 5'd10, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000015d, 5'd16, 27'h000001ce, 5'd23, 27'h000002e4, 32'h00000400,
  1'd1,  5'd22, 27'h0000005c, 5'd30, 27'h0000015d, 5'd5, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000278, 5'd30, 27'h0000004f, 5'd14, 27'h00000047, 32'h00000400,
  1'd1,  5'd23, 27'h0000001b, 5'd26, 27'h00000256, 5'd20, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c9, 5'd5, 27'h00000290, 5'd6, 27'h000003a2, 32'h00000400,
  1'd1,  5'd0, 27'h000003d3, 5'd5, 27'h00000143, 5'd16, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f0, 5'd10, 27'h00000058, 5'd26, 27'h00000116, 32'h00000400,
  1'd1,  5'd2, 27'h000001e5, 5'd15, 27'h000003bd, 5'd7, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000a7, 5'd17, 27'h000000c8, 5'd19, 27'h000000d1, 32'h00000400,
  1'd1,  5'd0, 27'h000003fc, 5'd17, 27'h00000330, 5'd29, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000017e, 5'd28, 27'h000001c1, 5'd6, 27'h000001fc, 32'h00000400,
  1'd1,  5'd2, 27'h000003b7, 5'd30, 27'h00000102, 5'd15, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000194, 5'd27, 27'h00000213, 5'd30, 27'h00000111, 32'h00000400,
  1'd1,  5'd12, 27'h000000a3, 5'd6, 27'h000003d3, 5'd8, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000319, 5'd9, 27'h00000224, 5'd16, 27'h000000d6, 32'h00000400,
  1'd1,  5'd15, 27'h000001c7, 5'd6, 27'h0000018d, 5'd28, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000dd, 5'd17, 27'h00000355, 5'd9, 27'h00000162, 32'h00000400,
  1'd1,  5'd12, 27'h0000008a, 5'd19, 27'h000002a0, 5'd19, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000026a, 5'd15, 27'h00000346, 5'd28, 27'h0000006f, 32'h00000400,
  1'd1,  5'd13, 27'h00000282, 5'd30, 27'h000002a2, 5'd6, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000194, 5'd27, 27'h000002d7, 5'd16, 27'h0000015d, 32'h00000400,
  1'd1,  5'd10, 27'h0000033a, 5'd30, 27'h0000027d, 5'd26, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000373, 5'd5, 27'h00000256, 5'd6, 27'h000001e2, 32'h00000400,
  1'd1,  5'd22, 27'h000002eb, 5'd5, 27'h000003c6, 5'd16, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000c5, 5'd8, 27'h00000222, 5'd28, 27'h000003bc, 32'h00000400,
  1'd1,  5'd24, 27'h000001e6, 5'd20, 27'h00000065, 5'd9, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000000e, 5'd18, 27'h00000144, 5'd19, 27'h000003b2, 32'h00000400,
  1'd1,  5'd22, 27'h0000039d, 5'd16, 27'h000000b7, 5'd26, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ec, 5'd29, 27'h00000254, 5'd5, 27'h000002c7, 32'h00000400,
  1'd1,  5'd21, 27'h000001d1, 5'd26, 27'h000002d7, 5'd17, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001cb, 5'd28, 27'h000003fb, 5'd30, 27'h00000365, 32'h00000400,
  1'd1,  5'd7, 27'h00000009, 5'd0, 27'h000000f1, 5'd8, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ab, 5'd5, 27'h00000008, 5'd15, 27'h00000225, 32'h00000400,
  1'd1,  5'd10, 27'h00000150, 5'd4, 27'h000002ba, 5'd28, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000309, 5'd13, 27'h00000210, 5'd4, 27'h000002cb, 32'h00000400,
  1'd1,  5'd9, 27'h00000090, 5'd15, 27'h000001b4, 5'd15, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000036e, 5'd12, 27'h000001ff, 5'd24, 27'h00000167, 32'h00000400,
  1'd1,  5'd8, 27'h0000018b, 5'd23, 27'h00000359, 5'd0, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000020f, 5'd23, 27'h000002bb, 5'd12, 27'h00000350, 32'h00000400,
  1'd1,  5'd7, 27'h00000275, 5'd22, 27'h0000036a, 5'd24, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000034c, 5'd1, 27'h0000019a, 5'd9, 27'h0000013d, 32'h00000400,
  1'd1,  5'd15, 27'h000002b3, 5'd2, 27'h00000050, 5'd18, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000188, 5'd4, 27'h000003ae, 5'd30, 27'h00000353, 32'h00000400,
  1'd1,  5'd18, 27'h0000019c, 5'd14, 27'h000001d6, 5'd1, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002c7, 5'd11, 27'h00000378, 5'd15, 27'h000001c8, 32'h00000400,
  1'd1,  5'd15, 27'h0000037d, 5'd14, 27'h00000148, 5'd21, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001a8, 5'd25, 27'h000001a1, 5'd0, 27'h00000123, 32'h00000400,
  1'd1,  5'd19, 27'h000002a0, 5'd23, 27'h0000035b, 5'd11, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000399, 5'd20, 27'h000003cf, 5'd24, 27'h000003b1, 32'h00000400,
  1'd1,  5'd26, 27'h0000007c, 5'd4, 27'h00000168, 5'd2, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f5, 5'd1, 27'h0000005a, 5'd10, 27'h000002d7, 32'h00000400,
  1'd1,  5'd27, 27'h00000001, 5'd0, 27'h000002ae, 5'd23, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b2, 5'd10, 27'h00000252, 5'd4, 27'h00000310, 32'h00000400,
  1'd1,  5'd28, 27'h000002b8, 5'd12, 27'h00000217, 5'd15, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000be, 5'd10, 27'h00000181, 5'd22, 27'h00000159, 32'h00000400,
  1'd1,  5'd30, 27'h00000309, 5'd20, 27'h00000309, 5'd1, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000044, 5'd22, 27'h0000027b, 5'd14, 27'h000000a1, 32'h00000400,
  1'd1,  5'd27, 27'h000002d2, 5'd25, 27'h000000eb, 5'd21, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000261, 5'd1, 27'h0000013f, 5'd1, 27'h0000029d, 32'h00000400,
  1'd1,  5'd10, 27'h00000045, 5'd0, 27'h00000049, 5'd12, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000381, 5'd1, 27'h00000202, 5'd22, 27'h00000285, 32'h00000400,
  1'd1,  5'd9, 27'h0000010a, 5'd13, 27'h00000259, 5'd6, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000056, 5'd10, 27'h0000027c, 5'd20, 27'h000000c8, 32'h00000400,
  1'd1,  5'd6, 27'h00000188, 5'd10, 27'h0000022a, 5'd27, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000022, 5'd23, 27'h0000021d, 5'd9, 27'h000002a9, 32'h00000400,
  1'd1,  5'd6, 27'h000001ce, 5'd21, 27'h00000145, 5'd20, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000074, 5'd23, 27'h00000219, 5'd27, 27'h000000f9, 32'h00000400,
  1'd1,  5'd16, 27'h00000024, 5'd0, 27'h000000d2, 5'd0, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000c3, 5'd3, 27'h0000027e, 5'd10, 27'h000002de, 32'h00000400,
  1'd1,  5'd19, 27'h000003bb, 5'd4, 27'h000001c9, 5'd21, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000036d, 5'd14, 27'h000001b2, 5'd8, 27'h00000311, 32'h00000400,
  1'd1,  5'd16, 27'h00000183, 5'd12, 27'h000001fe, 5'd16, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000286, 5'd10, 27'h0000024f, 5'd28, 27'h000002e6, 32'h00000400,
  1'd1,  5'd15, 27'h00000388, 5'd24, 27'h0000038e, 5'd5, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000005e, 5'd21, 27'h00000101, 5'd19, 27'h00000354, 32'h00000400,
  1'd1,  5'd20, 27'h000000e0, 5'd25, 27'h00000131, 5'd26, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f9, 5'd0, 27'h0000016b, 5'd6, 27'h00000138, 32'h00000400,
  1'd1,  5'd28, 27'h0000006d, 5'd4, 27'h0000024b, 5'd18, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000004a, 5'd4, 27'h0000020f, 5'd27, 27'h0000011c, 32'h00000400,
  1'd1,  5'd26, 27'h00000331, 5'd10, 27'h00000386, 5'd6, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d8, 5'd12, 27'h00000072, 5'd17, 27'h000003a1, 32'h00000400,
  1'd1,  5'd28, 27'h000002d2, 5'd14, 27'h00000297, 5'd26, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000014e, 5'd21, 27'h00000145, 5'd6, 27'h00000076, 32'h00000400,
  1'd1,  5'd30, 27'h000002ee, 5'd22, 27'h00000351, 5'd19, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000167, 5'd20, 27'h000002d8, 5'd27, 27'h0000015f, 32'h00000400,
  1'd1,  5'd7, 27'h00000145, 5'd6, 27'h000001fc, 5'd1, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003c5, 5'd7, 27'h000002b6, 5'd13, 27'h000000be, 32'h00000400,
  1'd1,  5'd7, 27'h00000388, 5'd5, 27'h00000324, 5'd22, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000158, 5'd18, 27'h000001b8, 5'd1, 27'h0000038a, 32'h00000400,
  1'd1,  5'd5, 27'h0000012f, 5'd17, 27'h00000365, 5'd15, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000bd, 5'd16, 27'h0000005b, 5'd25, 27'h0000029c, 32'h00000400,
  1'd1,  5'd9, 27'h000001b2, 5'd26, 27'h000001b0, 5'd1, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003d4, 5'd30, 27'h00000325, 5'd11, 27'h00000136, 32'h00000400,
  1'd1,  5'd7, 27'h0000023d, 5'd28, 27'h0000012e, 5'd23, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003bc, 5'd7, 27'h00000025, 5'd3, 27'h0000008d, 32'h00000400,
  1'd1,  5'd18, 27'h0000038c, 5'd5, 27'h000000ef, 5'd10, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000027, 5'd5, 27'h000003f2, 5'd23, 27'h0000036d, 32'h00000400,
  1'd1,  5'd18, 27'h00000004, 5'd17, 27'h00000130, 5'd2, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000393, 5'd16, 27'h00000367, 5'd12, 27'h0000006d, 32'h00000400,
  1'd1,  5'd16, 27'h000002b1, 5'd19, 27'h00000013, 5'd25, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002cb, 5'd29, 27'h0000033c, 5'd2, 27'h00000381, 32'h00000400,
  1'd1,  5'd20, 27'h00000038, 5'd28, 27'h000000ef, 5'd11, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002d4, 5'd28, 27'h00000292, 5'd21, 27'h000000f1, 32'h00000400,
  1'd1,  5'd28, 27'h0000039e, 5'd9, 27'h0000034d, 5'd4, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000246, 5'd5, 27'h0000010c, 5'd11, 27'h00000210, 32'h00000400,
  1'd1,  5'd28, 27'h0000020c, 5'd8, 27'h0000012e, 5'd23, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000187, 5'd19, 27'h00000240, 5'd0, 27'h00000282, 32'h00000400,
  1'd1,  5'd29, 27'h000000e7, 5'd18, 27'h000003b1, 5'd14, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000058, 5'd15, 27'h00000337, 5'd22, 27'h000003af, 32'h00000400,
  1'd1,  5'd28, 27'h00000165, 5'd26, 27'h00000244, 5'd3, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000022f, 5'd29, 27'h00000180, 5'd11, 27'h000003a2, 32'h00000400,
  1'd1,  5'd25, 27'h000003ec, 5'd26, 27'h0000034a, 5'd25, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000170, 5'd7, 27'h000003ce, 5'd10, 27'h00000037, 32'h00000400,
  1'd1,  5'd6, 27'h00000027, 5'd6, 27'h000003ad, 5'd17, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000162, 5'd8, 27'h00000174, 5'd27, 27'h0000025f, 32'h00000400,
  1'd1,  5'd5, 27'h000002c9, 5'd16, 27'h000001e0, 5'd6, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002db, 5'd15, 27'h000002ca, 5'd17, 27'h00000392, 32'h00000400,
  1'd1,  5'd7, 27'h00000177, 5'd15, 27'h00000386, 5'd27, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000036, 5'd30, 27'h00000373, 5'd6, 27'h000002bc, 32'h00000400,
  1'd1,  5'd8, 27'h000000c5, 5'd28, 27'h0000037a, 5'd16, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000046, 5'd28, 27'h000001cb, 5'd26, 27'h000003fe, 32'h00000400,
  1'd1,  5'd19, 27'h000001d1, 5'd9, 27'h0000002c, 5'd5, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000148, 5'd7, 27'h000001b7, 5'd19, 27'h000003aa, 32'h00000400,
  1'd1,  5'd17, 27'h000001be, 5'd10, 27'h0000010b, 5'd29, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000028c, 5'd20, 27'h000000f7, 5'd9, 27'h00000377, 32'h00000400,
  1'd1,  5'd17, 27'h00000048, 5'd20, 27'h00000072, 5'd19, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000112, 5'd20, 27'h00000230, 5'd27, 27'h000002b9, 32'h00000400,
  1'd1,  5'd18, 27'h0000026a, 5'd27, 27'h00000360, 5'd8, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003bd, 5'd30, 27'h00000298, 5'd19, 27'h00000110, 32'h00000400,
  1'd1,  5'd18, 27'h000002b7, 5'd28, 27'h00000360, 5'd27, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000188, 5'd7, 27'h000001ed, 5'd10, 27'h000000ec, 32'h00000400,
  1'd1,  5'd27, 27'h000002b1, 5'd8, 27'h0000034e, 5'd17, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a3, 5'd7, 27'h000002d5, 5'd30, 27'h000002f0, 32'h00000400,
  1'd1,  5'd30, 27'h0000018e, 5'd15, 27'h00000367, 5'd8, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000031d, 5'd17, 27'h000000c1, 5'd18, 27'h000000a3, 32'h00000400,
  1'd1,  5'd25, 27'h000003c0, 5'd18, 27'h00000110, 5'd27, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e1, 5'd29, 27'h000002cb, 5'd8, 27'h00000396, 32'h00000400,
  1'd1,  5'd27, 27'h000000ea, 5'd29, 27'h00000175, 5'd20, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000247, 5'd29, 27'h00000099, 5'd27, 27'h000003ed, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003cd, 5'd1, 27'h0000006d, 5'd1, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b3, 5'd3, 27'h0000006a, 5'd11, 27'h00000163, 32'h00000400,
  1'd1,  5'd3, 27'h000000e0, 5'd2, 27'h00000343, 5'd21, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001fc, 5'd11, 27'h000003c7, 5'd1, 27'h0000001d, 32'h00000400,
  1'd1,  5'd3, 27'h00000382, 5'd12, 27'h00000346, 5'd14, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000d6, 5'd10, 27'h000003ba, 5'd21, 27'h000001e2, 32'h00000400,
  1'd1,  5'd1, 27'h00000172, 5'd22, 27'h000003b1, 5'd0, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002dc, 5'd24, 27'h0000005d, 5'd14, 27'h000002df, 32'h00000400,
  1'd1,  5'd2, 27'h0000021a, 5'd24, 27'h000000d2, 5'd22, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000304, 5'd1, 27'h0000020a, 5'd1, 27'h0000035d, 32'h00000400,
  1'd1,  5'd10, 27'h000002c6, 5'd2, 27'h000003c4, 5'd13, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035d, 5'd2, 27'h000002e6, 5'd24, 27'h000002b3, 32'h00000400,
  1'd1,  5'd15, 27'h0000016c, 5'd14, 27'h000002e6, 5'd0, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000357, 5'd12, 27'h00000055, 5'd14, 27'h000003a5, 32'h00000400,
  1'd1,  5'd11, 27'h0000000e, 5'd13, 27'h000003bc, 5'd21, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000110, 5'd21, 27'h000003b2, 5'd1, 27'h000002ae, 32'h00000400,
  1'd1,  5'd10, 27'h000002bb, 5'd21, 27'h00000039, 5'd13, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000117, 5'd23, 27'h000003f2, 5'd24, 27'h000003d5, 32'h00000400,
  1'd1,  5'd20, 27'h000002e3, 5'd5, 27'h00000029, 5'd1, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000182, 5'd1, 27'h00000345, 5'd14, 27'h000000ae, 32'h00000400,
  1'd1,  5'd24, 27'h000002e6, 5'd4, 27'h000001f4, 5'd23, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ec, 5'd12, 27'h0000006c, 5'd1, 27'h00000060, 32'h00000400,
  1'd1,  5'd22, 27'h00000231, 5'd11, 27'h0000029c, 5'd11, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000330, 5'd14, 27'h00000375, 5'd25, 27'h000000ce, 32'h00000400,
  1'd1,  5'd23, 27'h0000005f, 5'd22, 27'h00000103, 5'd3, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034d, 5'd21, 27'h000002ad, 5'd11, 27'h0000033d, 32'h00000400,
  1'd1,  5'd25, 27'h000001c6, 5'd23, 27'h00000375, 5'd22, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000044, 5'd2, 27'h000002fe, 5'd7, 27'h0000004c, 32'h00000400,
  1'd1,  5'd1, 27'h000003a8, 5'd0, 27'h0000039f, 5'd18, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000179, 5'd1, 27'h0000006c, 5'd27, 27'h000000de, 32'h00000400,
  1'd1,  5'd1, 27'h000002b8, 5'd14, 27'h00000254, 5'd5, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000dc, 5'd13, 27'h0000013d, 5'd17, 27'h000002a4, 32'h00000400,
  1'd1,  5'd2, 27'h0000027c, 5'd13, 27'h000002fb, 5'd29, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000207, 5'd21, 27'h0000013d, 5'd7, 27'h000001ea, 32'h00000400,
  1'd1,  5'd4, 27'h000003f1, 5'd23, 27'h000000ff, 5'd16, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000018, 5'd25, 27'h000002b9, 5'd28, 27'h00000177, 32'h00000400,
  1'd1,  5'd15, 27'h000000b7, 5'd0, 27'h00000000, 5'd5, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000224, 5'd2, 27'h0000024f, 5'd20, 27'h00000166, 32'h00000400,
  1'd1,  5'd10, 27'h00000216, 5'd4, 27'h00000393, 5'd30, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001d9, 5'd14, 27'h00000009, 5'd5, 27'h000001a1, 32'h00000400,
  1'd1,  5'd13, 27'h00000066, 5'd12, 27'h000000f2, 5'd19, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002fb, 5'd14, 27'h000000b1, 5'd26, 27'h000002f2, 32'h00000400,
  1'd1,  5'd11, 27'h000001e3, 5'd25, 27'h00000144, 5'd6, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f3, 5'd25, 27'h0000019c, 5'd18, 27'h000002ad, 32'h00000400,
  1'd1,  5'd15, 27'h00000116, 5'd21, 27'h00000108, 5'd26, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000197, 5'd2, 27'h000002b8, 5'd6, 27'h000000c5, 32'h00000400,
  1'd1,  5'd22, 27'h0000000b, 5'd0, 27'h000002dd, 5'd15, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003cb, 5'd0, 27'h0000011c, 5'd28, 27'h00000004, 32'h00000400,
  1'd1,  5'd25, 27'h000002f4, 5'd14, 27'h00000116, 5'd8, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000291, 5'd13, 27'h0000028a, 5'd19, 27'h00000283, 32'h00000400,
  1'd1,  5'd23, 27'h000002a6, 5'd11, 27'h000003c4, 5'd27, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000295, 5'd21, 27'h00000077, 5'd9, 27'h000003df, 32'h00000400,
  1'd1,  5'd21, 27'h0000009a, 5'd22, 27'h00000260, 5'd19, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000142, 5'd23, 27'h0000027a, 5'd28, 27'h000002aa, 32'h00000400,
  1'd1,  5'd0, 27'h000001d9, 5'd8, 27'h000000c8, 5'd3, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000cd, 5'd9, 27'h000003be, 5'd13, 27'h00000393, 32'h00000400,
  1'd1,  5'd3, 27'h000000c8, 5'd5, 27'h000000cf, 5'd24, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000072, 5'd16, 27'h0000036b, 5'd4, 27'h00000179, 32'h00000400,
  1'd1,  5'd1, 27'h000000b0, 5'd20, 27'h0000020b, 5'd10, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001d9, 5'd20, 27'h000001ac, 5'd25, 27'h000001a6, 32'h00000400,
  1'd1,  5'd2, 27'h00000096, 5'd29, 27'h00000381, 5'd3, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000220, 5'd29, 27'h00000010, 5'd14, 27'h000000d0, 32'h00000400,
  1'd1,  5'd0, 27'h000002b7, 5'd29, 27'h00000275, 5'd25, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000019a, 5'd7, 27'h0000008d, 5'd2, 27'h000001f1, 32'h00000400,
  1'd1,  5'd14, 27'h00000305, 5'd7, 27'h0000033c, 5'd11, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000046, 5'd9, 27'h000000fb, 5'd23, 27'h00000226, 32'h00000400,
  1'd1,  5'd14, 27'h000000d9, 5'd20, 27'h0000009e, 5'd2, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001e2, 5'd17, 27'h000003c4, 5'd15, 27'h00000094, 32'h00000400,
  1'd1,  5'd10, 27'h00000181, 5'd16, 27'h000002fc, 5'd24, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000341, 5'd29, 27'h0000006a, 5'd3, 27'h00000265, 32'h00000400,
  1'd1,  5'd12, 27'h000002c7, 5'd26, 27'h000002fe, 5'd15, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000040, 5'd30, 27'h00000116, 5'd23, 27'h0000015c, 32'h00000400,
  1'd1,  5'd24, 27'h000001ef, 5'd5, 27'h00000252, 5'd2, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000bd, 5'd8, 27'h000001d8, 5'd14, 27'h000002aa, 32'h00000400,
  1'd1,  5'd21, 27'h00000241, 5'd6, 27'h00000282, 5'd21, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001e5, 5'd16, 27'h00000288, 5'd1, 27'h000002a4, 32'h00000400,
  1'd1,  5'd24, 27'h00000081, 5'd19, 27'h00000371, 5'd12, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000016, 5'd17, 27'h0000005f, 5'd24, 27'h000000af, 32'h00000400,
  1'd1,  5'd25, 27'h0000034e, 5'd28, 27'h0000034f, 5'd1, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000019e, 5'd26, 27'h00000057, 5'd12, 27'h00000325, 32'h00000400,
  1'd1,  5'd24, 27'h00000158, 5'd29, 27'h00000309, 5'd22, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c8, 5'd6, 27'h000001cd, 5'd9, 27'h00000286, 32'h00000400,
  1'd1,  5'd0, 27'h00000037, 5'd7, 27'h000001f4, 5'd15, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000001a, 5'd5, 27'h00000208, 5'd29, 27'h000003a7, 32'h00000400,
  1'd1,  5'd4, 27'h000003a9, 5'd20, 27'h0000020e, 5'd7, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000e6, 5'd17, 27'h00000025, 5'd15, 27'h000003a3, 32'h00000400,
  1'd1,  5'd0, 27'h00000348, 5'd16, 27'h00000113, 5'd28, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000010c, 5'd26, 27'h000002c7, 5'd7, 27'h000002fd, 32'h00000400,
  1'd1,  5'd0, 27'h00000007, 5'd28, 27'h000003c8, 5'd16, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000011, 5'd28, 27'h00000038, 5'd26, 27'h00000326, 32'h00000400,
  1'd1,  5'd14, 27'h0000002c, 5'd5, 27'h000001f6, 5'd8, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001cc, 5'd5, 27'h000001bc, 5'd15, 27'h000002f4, 32'h00000400,
  1'd1,  5'd15, 27'h0000008c, 5'd8, 27'h000000b5, 5'd26, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000005d, 5'd17, 27'h0000019d, 5'd9, 27'h000002ea, 32'h00000400,
  1'd1,  5'd15, 27'h00000109, 5'd16, 27'h0000036a, 5'd15, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008b, 5'd20, 27'h00000192, 5'd28, 27'h0000004d, 32'h00000400,
  1'd1,  5'd15, 27'h00000158, 5'd30, 27'h00000375, 5'd7, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000146, 5'd29, 27'h00000338, 5'd17, 27'h0000035a, 32'h00000400,
  1'd1,  5'd13, 27'h000000ca, 5'd27, 27'h000000f6, 5'd30, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000147, 5'd10, 27'h00000119, 5'd8, 27'h0000035d, 32'h00000400,
  1'd1,  5'd24, 27'h000002f0, 5'd5, 27'h00000120, 5'd17, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000369, 5'd8, 27'h000003a2, 5'd28, 27'h0000024f, 32'h00000400,
  1'd1,  5'd22, 27'h00000079, 5'd19, 27'h000000b4, 5'd6, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003c6, 5'd18, 27'h000001d5, 5'd16, 27'h00000279, 32'h00000400,
  1'd1,  5'd21, 27'h00000101, 5'd16, 27'h000002de, 5'd29, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000146, 5'd26, 27'h000000ca, 5'd9, 27'h00000053, 32'h00000400,
  1'd1,  5'd23, 27'h0000029d, 5'd30, 27'h0000023d, 5'd17, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ba, 5'd28, 27'h00000231, 5'd28, 27'h000003d9, 32'h00000400,
  1'd1,  5'd8, 27'h000003eb, 5'd4, 27'h000002ba, 5'd8, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000230, 5'd0, 27'h000000e3, 5'd18, 27'h0000010a, 32'h00000400,
  1'd1,  5'd7, 27'h00000032, 5'd3, 27'h00000172, 5'd28, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001c1, 5'd13, 27'h000003f5, 5'd5, 27'h0000004b, 32'h00000400,
  1'd1,  5'd8, 27'h0000024c, 5'd14, 27'h00000296, 5'd14, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000029e, 5'd12, 27'h000000d9, 5'd25, 27'h00000215, 32'h00000400,
  1'd1,  5'd9, 27'h0000029a, 5'd25, 27'h000001f8, 5'd4, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000164, 5'd21, 27'h0000014f, 5'd13, 27'h00000165, 32'h00000400,
  1'd1,  5'd6, 27'h00000339, 5'd22, 27'h0000016e, 5'd24, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003ec, 5'd0, 27'h000003ef, 5'd9, 27'h00000215, 32'h00000400,
  1'd1,  5'd17, 27'h000001fd, 5'd4, 27'h00000130, 5'd19, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032a, 5'd2, 27'h00000274, 5'd26, 27'h00000299, 32'h00000400,
  1'd1,  5'd19, 27'h000001bf, 5'd15, 27'h000001a8, 5'd1, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001dd, 5'd13, 27'h0000022d, 5'd10, 27'h00000381, 32'h00000400,
  1'd1,  5'd18, 27'h00000189, 5'd13, 27'h00000123, 5'd20, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000048, 5'd24, 27'h0000017c, 5'd2, 27'h0000026d, 32'h00000400,
  1'd1,  5'd18, 27'h00000077, 5'd23, 27'h000002e9, 5'd11, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000074, 5'd24, 27'h00000276, 5'd25, 27'h0000002b, 32'h00000400,
  1'd1,  5'd30, 27'h0000030a, 5'd3, 27'h00000139, 5'd5, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000052, 5'd2, 27'h0000007c, 5'd13, 27'h000000ac, 32'h00000400,
  1'd1,  5'd29, 27'h000003f0, 5'd1, 27'h0000038e, 5'd24, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000375, 5'd15, 27'h0000007f, 5'd1, 27'h00000005, 32'h00000400,
  1'd1,  5'd30, 27'h0000018d, 5'd12, 27'h000002ba, 5'd14, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000203, 5'd12, 27'h00000041, 5'd24, 27'h0000018a, 32'h00000400,
  1'd1,  5'd30, 27'h000003e3, 5'd21, 27'h0000003d, 5'd1, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000375, 5'd21, 27'h00000330, 5'd14, 27'h00000197, 32'h00000400,
  1'd1,  5'd30, 27'h0000029d, 5'd25, 27'h000001c4, 5'd22, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000026d, 5'd4, 27'h000000ee, 5'd1, 27'h000000bb, 32'h00000400,
  1'd1,  5'd10, 27'h0000002a, 5'd4, 27'h00000274, 5'd15, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000030d, 5'd1, 27'h0000022a, 5'd23, 27'h000000a2, 32'h00000400,
  1'd1,  5'd5, 27'h00000332, 5'd14, 27'h00000252, 5'd5, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000113, 5'd10, 27'h000002c9, 5'd16, 27'h00000096, 32'h00000400,
  1'd1,  5'd7, 27'h0000020c, 5'd14, 27'h00000000, 5'd28, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d7, 5'd24, 27'h0000030d, 5'd6, 27'h0000022b, 32'h00000400,
  1'd1,  5'd8, 27'h0000027f, 5'd25, 27'h000002d5, 5'd20, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ac, 5'd21, 27'h00000336, 5'd28, 27'h00000168, 32'h00000400,
  1'd1,  5'd18, 27'h0000000d, 5'd4, 27'h0000038f, 5'd0, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001bf, 5'd0, 27'h00000273, 5'd11, 27'h000002af, 32'h00000400,
  1'd1,  5'd18, 27'h00000364, 5'd1, 27'h0000038a, 5'd23, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000035c, 5'd10, 27'h00000321, 5'd10, 27'h000000cb, 32'h00000400,
  1'd1,  5'd16, 27'h0000033a, 5'd13, 27'h000001bc, 5'd19, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000030d, 5'd14, 27'h0000023f, 5'd27, 27'h00000191, 32'h00000400,
  1'd1,  5'd20, 27'h00000208, 5'd25, 27'h000002fd, 5'd8, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000351, 5'd23, 27'h000000d3, 5'd17, 27'h00000028, 32'h00000400,
  1'd1,  5'd17, 27'h000000b1, 5'd25, 27'h000002ca, 5'd27, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000175, 5'd4, 27'h000000d4, 5'd9, 27'h000003d8, 32'h00000400,
  1'd1,  5'd30, 27'h000002fb, 5'd0, 27'h00000084, 5'd18, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000054, 5'd2, 27'h000000d2, 5'd29, 27'h000003c1, 32'h00000400,
  1'd1,  5'd26, 27'h00000300, 5'd11, 27'h0000035e, 5'd9, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000146, 5'd11, 27'h00000313, 5'd17, 27'h000000b9, 32'h00000400,
  1'd1,  5'd29, 27'h00000155, 5'd10, 27'h000002a9, 5'd29, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c5, 5'd21, 27'h0000017b, 5'd6, 27'h00000235, 32'h00000400,
  1'd1,  5'd27, 27'h000002f7, 5'd25, 27'h00000218, 5'd19, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024c, 5'd25, 27'h00000216, 5'd29, 27'h00000287, 32'h00000400,
  1'd1,  5'd8, 27'h000003eb, 5'd8, 27'h00000295, 5'd4, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000013f, 5'd7, 27'h00000115, 5'd12, 27'h000003c5, 32'h00000400,
  1'd1,  5'd10, 27'h000000ed, 5'd8, 27'h0000012d, 5'd24, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000e6, 5'd16, 27'h0000024b, 5'd0, 27'h000002e6, 32'h00000400,
  1'd1,  5'd6, 27'h00000211, 5'd18, 27'h0000033e, 5'd14, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000089, 5'd15, 27'h0000034b, 5'd25, 27'h0000032e, 32'h00000400,
  1'd1,  5'd7, 27'h00000314, 5'd27, 27'h000002fd, 5'd2, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b9, 5'd26, 27'h00000010, 5'd10, 27'h0000030e, 32'h00000400,
  1'd1,  5'd8, 27'h000001c1, 5'd28, 27'h000002c8, 5'd21, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000345, 5'd8, 27'h000000d9, 5'd2, 27'h0000021a, 32'h00000400,
  1'd1,  5'd18, 27'h000003d0, 5'd6, 27'h0000034e, 5'd12, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000c5, 5'd9, 27'h00000102, 5'd25, 27'h00000253, 32'h00000400,
  1'd1,  5'd16, 27'h0000020b, 5'd19, 27'h0000014f, 5'd4, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000205, 5'd17, 27'h00000019, 5'd13, 27'h0000038f, 32'h00000400,
  1'd1,  5'd18, 27'h00000182, 5'd18, 27'h0000033b, 5'd24, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001c, 5'd30, 27'h0000038c, 5'd3, 27'h000002c9, 32'h00000400,
  1'd1,  5'd15, 27'h00000331, 5'd29, 27'h00000039, 5'd15, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000297, 5'd27, 27'h000000b5, 5'd21, 27'h000002c1, 32'h00000400,
  1'd1,  5'd28, 27'h000000cd, 5'd7, 27'h0000013d, 5'd2, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003c6, 5'd9, 27'h000002aa, 5'd11, 27'h000001ba, 32'h00000400,
  1'd1,  5'd28, 27'h000002f2, 5'd8, 27'h000003b4, 5'd20, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000023, 5'd17, 27'h00000232, 5'd1, 27'h000000f3, 32'h00000400,
  1'd1,  5'd27, 27'h0000014c, 5'd17, 27'h0000025a, 5'd11, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001b7, 5'd15, 27'h0000024e, 5'd21, 27'h00000191, 32'h00000400,
  1'd1,  5'd26, 27'h000000cb, 5'd30, 27'h000003bc, 5'd4, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001f0, 5'd29, 27'h00000330, 5'd12, 27'h0000018c, 32'h00000400,
  1'd1,  5'd27, 27'h00000003, 5'd27, 27'h000003e0, 5'd24, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001d7, 5'd8, 27'h00000219, 5'd9, 27'h00000197, 32'h00000400,
  1'd1,  5'd6, 27'h000000e2, 5'd6, 27'h000001a1, 5'd17, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003bc, 5'd8, 27'h0000001f, 5'd27, 27'h000001ce, 32'h00000400,
  1'd1,  5'd8, 27'h000000e5, 5'd17, 27'h0000000c, 5'd9, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002fe, 5'd19, 27'h0000033d, 5'd18, 27'h00000218, 32'h00000400,
  1'd1,  5'd10, 27'h000000bd, 5'd16, 27'h00000291, 5'd29, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000018b, 5'd28, 27'h0000031b, 5'd9, 27'h00000158, 32'h00000400,
  1'd1,  5'd8, 27'h000003ef, 5'd27, 27'h000000e9, 5'd18, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e3, 5'd28, 27'h000000c0, 5'd27, 27'h0000010b, 32'h00000400,
  1'd1,  5'd18, 27'h000002ce, 5'd6, 27'h000000e0, 5'd5, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029f, 5'd7, 27'h00000223, 5'd18, 27'h00000341, 32'h00000400,
  1'd1,  5'd18, 27'h0000022f, 5'd8, 27'h000001e9, 5'd26, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000349, 5'd16, 27'h000001ec, 5'd6, 27'h00000166, 32'h00000400,
  1'd1,  5'd17, 27'h000001f8, 5'd17, 27'h00000379, 5'd19, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000379, 5'd20, 27'h0000026d, 5'd28, 27'h0000003c, 32'h00000400,
  1'd1,  5'd18, 27'h0000006d, 5'd29, 27'h000003e4, 5'd9, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f9, 5'd28, 27'h000002b2, 5'd19, 27'h000000b4, 32'h00000400,
  1'd1,  5'd16, 27'h000002fb, 5'd30, 27'h00000179, 5'd27, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000096, 5'd8, 27'h000003f1, 5'd6, 27'h0000008e, 32'h00000400,
  1'd1,  5'd27, 27'h00000047, 5'd5, 27'h00000121, 5'd20, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ef, 5'd6, 27'h0000034f, 5'd30, 27'h00000181, 32'h00000400,
  1'd1,  5'd27, 27'h000002d4, 5'd15, 27'h0000038c, 5'd10, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000332, 5'd19, 27'h00000226, 5'd19, 27'h0000027a, 32'h00000400,
  1'd1,  5'd30, 27'h000003db, 5'd19, 27'h000001b9, 5'd28, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000015a, 5'd29, 27'h000003a1, 5'd7, 27'h0000017b, 32'h00000400,
  1'd1,  5'd27, 27'h00000207, 5'd30, 27'h000002b0, 5'd19, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000155, 5'd26, 27'h00000186, 5'd26, 27'h0000037d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000017d, 5'd1, 27'h000000b8, 5'd1, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e1, 5'd1, 27'h000001a3, 5'd13, 27'h0000001d, 32'h00000400,
  1'd1,  5'd1, 27'h000000d4, 5'd0, 27'h00000032, 5'd21, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000062, 5'd13, 27'h000002d6, 5'd3, 27'h000003d5, 32'h00000400,
  1'd1,  5'd0, 27'h00000229, 5'd14, 27'h00000335, 5'd12, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000009a, 5'd11, 27'h000002e3, 5'd23, 27'h0000035d, 32'h00000400,
  1'd1,  5'd2, 27'h0000028c, 5'd21, 27'h000000bd, 5'd4, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000070, 5'd25, 27'h0000033c, 5'd13, 27'h000002bc, 32'h00000400,
  1'd1,  5'd0, 27'h000003dc, 5'd22, 27'h00000050, 5'd21, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000075, 5'd1, 27'h000003ac, 5'd5, 27'h0000003c, 32'h00000400,
  1'd1,  5'd13, 27'h00000004, 5'd4, 27'h00000359, 5'd15, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000218, 5'd0, 27'h0000009d, 5'd22, 27'h000002d3, 32'h00000400,
  1'd1,  5'd10, 27'h000001ae, 5'd14, 27'h00000199, 5'd4, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000204, 5'd14, 27'h000002f2, 5'd13, 27'h00000393, 32'h00000400,
  1'd1,  5'd10, 27'h0000026d, 5'd13, 27'h00000151, 5'd21, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000165, 5'd24, 27'h00000336, 5'd5, 27'h00000090, 32'h00000400,
  1'd1,  5'd11, 27'h00000340, 5'd24, 27'h00000276, 5'd10, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001fd, 5'd25, 27'h0000011c, 5'd25, 27'h000002d7, 32'h00000400,
  1'd1,  5'd23, 27'h000001f3, 5'd4, 27'h00000333, 5'd4, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000018c, 5'd3, 27'h000000f1, 5'd12, 27'h00000368, 32'h00000400,
  1'd1,  5'd20, 27'h000002ab, 5'd3, 27'h000002ad, 5'd21, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000025e, 5'd11, 27'h000003a4, 5'd1, 27'h000000b4, 32'h00000400,
  1'd1,  5'd24, 27'h000000c0, 5'd12, 27'h0000005b, 5'd14, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000375, 5'd14, 27'h0000021a, 5'd20, 27'h00000340, 32'h00000400,
  1'd1,  5'd24, 27'h00000034, 5'd24, 27'h000002f4, 5'd4, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000018e, 5'd23, 27'h000003a1, 5'd10, 27'h0000021c, 32'h00000400,
  1'd1,  5'd21, 27'h00000051, 5'd22, 27'h00000048, 5'd21, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f4, 5'd1, 27'h000000f9, 5'd8, 27'h00000057, 32'h00000400,
  1'd1,  5'd3, 27'h00000146, 5'd1, 27'h000001ea, 5'd18, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000034b, 5'd4, 27'h00000145, 5'd29, 27'h00000085, 32'h00000400,
  1'd1,  5'd3, 27'h000001d0, 5'd13, 27'h00000023, 5'd5, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000291, 5'd15, 27'h00000135, 5'd20, 27'h0000028b, 32'h00000400,
  1'd1,  5'd4, 27'h00000309, 5'd10, 27'h0000025c, 5'd30, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000038e, 5'd21, 27'h000003ec, 5'd9, 27'h0000027f, 32'h00000400,
  1'd1,  5'd0, 27'h000003bc, 5'd23, 27'h000001ac, 5'd17, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000045, 5'd22, 27'h000001d0, 5'd30, 27'h000002fe, 32'h00000400,
  1'd1,  5'd13, 27'h00000056, 5'd4, 27'h0000035d, 5'd5, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f6, 5'd1, 27'h000002ff, 5'd16, 27'h000001dd, 32'h00000400,
  1'd1,  5'd11, 27'h000002a7, 5'd3, 27'h000000a1, 5'd29, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002a3, 5'd13, 27'h00000032, 5'd7, 27'h0000036b, 32'h00000400,
  1'd1,  5'd15, 27'h000001ea, 5'd10, 27'h000003be, 5'd19, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002dc, 5'd15, 27'h000001f1, 5'd30, 27'h000001d6, 32'h00000400,
  1'd1,  5'd14, 27'h00000306, 5'd21, 27'h000003d8, 5'd5, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000127, 5'd25, 27'h000001e1, 5'd16, 27'h000002bb, 32'h00000400,
  1'd1,  5'd14, 27'h000003ab, 5'd22, 27'h0000037b, 5'd27, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000166, 5'd3, 27'h000003cd, 5'd9, 27'h0000031d, 32'h00000400,
  1'd1,  5'd24, 27'h00000206, 5'd4, 27'h0000039f, 5'd18, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002c1, 5'd3, 27'h0000038a, 5'd25, 27'h0000036b, 32'h00000400,
  1'd1,  5'd21, 27'h000003f8, 5'd14, 27'h0000022f, 5'd6, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000128, 5'd11, 27'h000000a8, 5'd19, 27'h0000013d, 32'h00000400,
  1'd1,  5'd25, 27'h000002b3, 5'd11, 27'h0000015d, 5'd28, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000033a, 5'd22, 27'h000000da, 5'd5, 27'h00000361, 32'h00000400,
  1'd1,  5'd24, 27'h000000c3, 5'd23, 27'h00000380, 5'd16, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000003f, 5'd22, 27'h000000b3, 5'd30, 27'h0000015b, 32'h00000400,
  1'd1,  5'd0, 27'h00000392, 5'd10, 27'h000000bc, 5'd1, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000066, 5'd5, 27'h0000016c, 5'd15, 27'h00000134, 32'h00000400,
  1'd1,  5'd0, 27'h0000016b, 5'd6, 27'h00000097, 5'd21, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f4, 5'd19, 27'h000002e9, 5'd3, 27'h00000063, 32'h00000400,
  1'd1,  5'd1, 27'h0000032b, 5'd19, 27'h0000013d, 5'd12, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003cd, 5'd16, 27'h0000033f, 5'd25, 27'h0000034e, 32'h00000400,
  1'd1,  5'd0, 27'h00000216, 5'd29, 27'h00000365, 5'd3, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000012b, 5'd28, 27'h00000328, 5'd13, 27'h0000020d, 32'h00000400,
  1'd1,  5'd2, 27'h0000012f, 5'd26, 27'h000002ac, 5'd20, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029c, 5'd6, 27'h00000137, 5'd3, 27'h0000032f, 32'h00000400,
  1'd1,  5'd11, 27'h00000196, 5'd6, 27'h00000312, 5'd11, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002e3, 5'd10, 27'h00000147, 5'd23, 27'h00000341, 32'h00000400,
  1'd1,  5'd10, 27'h00000314, 5'd19, 27'h00000264, 5'd2, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025d, 5'd16, 27'h00000399, 5'd12, 27'h000001c2, 32'h00000400,
  1'd1,  5'd11, 27'h00000086, 5'd18, 27'h00000218, 5'd23, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000025e, 5'd28, 27'h0000019a, 5'd4, 27'h00000342, 32'h00000400,
  1'd1,  5'd15, 27'h000001da, 5'd30, 27'h000003af, 5'd10, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000032f, 5'd29, 27'h000002f5, 5'd24, 27'h000001cd, 32'h00000400,
  1'd1,  5'd23, 27'h000002bb, 5'd9, 27'h000001f3, 5'd4, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000375, 5'd10, 27'h00000073, 5'd13, 27'h0000016e, 32'h00000400,
  1'd1,  5'd24, 27'h00000127, 5'd6, 27'h000001e1, 5'd25, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000292, 5'd19, 27'h000003e6, 5'd4, 27'h0000002a, 32'h00000400,
  1'd1,  5'd22, 27'h000002d0, 5'd17, 27'h000001df, 5'd15, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000020f, 5'd15, 27'h000003d6, 5'd21, 27'h000000d6, 32'h00000400,
  1'd1,  5'd23, 27'h000003a3, 5'd27, 27'h00000006, 5'd4, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000018c, 5'd26, 27'h00000091, 5'd10, 27'h000001bf, 32'h00000400,
  1'd1,  5'd22, 27'h00000032, 5'd27, 27'h000000bf, 5'd24, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000385, 5'd5, 27'h00000155, 5'd9, 27'h00000157, 32'h00000400,
  1'd1,  5'd1, 27'h000001d6, 5'd9, 27'h000002e5, 5'd18, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000035a, 5'd7, 27'h00000023, 5'd29, 27'h00000305, 32'h00000400,
  1'd1,  5'd0, 27'h00000025, 5'd16, 27'h000003de, 5'd9, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000052, 5'd19, 27'h000003e1, 5'd18, 27'h000001b9, 32'h00000400,
  1'd1,  5'd2, 27'h000000a3, 5'd17, 27'h00000320, 5'd29, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002e2, 5'd28, 27'h00000108, 5'd6, 27'h000003cf, 32'h00000400,
  1'd1,  5'd0, 27'h00000110, 5'd28, 27'h000002d6, 5'd19, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000212, 5'd26, 27'h00000088, 5'd30, 27'h0000002c, 32'h00000400,
  1'd1,  5'd14, 27'h000001d4, 5'd6, 27'h00000273, 5'd8, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000341, 5'd9, 27'h0000022f, 5'd17, 27'h000001d2, 32'h00000400,
  1'd1,  5'd13, 27'h00000309, 5'd7, 27'h00000059, 5'd28, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000054, 5'd19, 27'h000003b7, 5'd9, 27'h000002a5, 32'h00000400,
  1'd1,  5'd14, 27'h00000185, 5'd19, 27'h0000004f, 5'd15, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021b, 5'd17, 27'h0000013f, 5'd29, 27'h0000019a, 32'h00000400,
  1'd1,  5'd11, 27'h00000062, 5'd30, 27'h00000349, 5'd6, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001be, 5'd30, 27'h00000359, 5'd18, 27'h000003ad, 32'h00000400,
  1'd1,  5'd13, 27'h00000052, 5'd30, 27'h0000034a, 5'd26, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000186, 5'd5, 27'h0000022d, 5'd9, 27'h00000176, 32'h00000400,
  1'd1,  5'd21, 27'h00000395, 5'd7, 27'h0000026b, 5'd20, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000115, 5'd9, 27'h00000188, 5'd30, 27'h0000019f, 32'h00000400,
  1'd1,  5'd21, 27'h00000310, 5'd16, 27'h000000b3, 5'd6, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d1, 5'd18, 27'h0000000b, 5'd20, 27'h0000029e, 32'h00000400,
  1'd1,  5'd23, 27'h00000358, 5'd18, 27'h000002cf, 5'd29, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ff, 5'd30, 27'h00000138, 5'd6, 27'h00000349, 32'h00000400,
  1'd1,  5'd25, 27'h000000c1, 5'd26, 27'h00000066, 5'd19, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000327, 5'd30, 27'h00000380, 5'd27, 27'h0000039e, 32'h00000400,
  1'd1,  5'd6, 27'h0000034f, 5'd2, 27'h0000022d, 5'd7, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000031f, 5'd2, 27'h000000b3, 5'd16, 27'h00000197, 32'h00000400,
  1'd1,  5'd5, 27'h000001d4, 5'd0, 27'h0000015f, 5'd28, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e7, 5'd15, 27'h000000c1, 5'd0, 27'h000003e3, 32'h00000400,
  1'd1,  5'd7, 27'h000002b1, 5'd13, 27'h00000211, 5'd11, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020b, 5'd10, 27'h00000211, 5'd21, 27'h00000134, 32'h00000400,
  1'd1,  5'd8, 27'h0000016e, 5'd20, 27'h000002ca, 5'd2, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000213, 5'd24, 27'h000000a2, 5'd10, 27'h000002ef, 32'h00000400,
  1'd1,  5'd8, 27'h000001a1, 5'd25, 27'h00000203, 5'd22, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000024a, 5'd0, 27'h0000023d, 5'd10, 27'h00000052, 32'h00000400,
  1'd1,  5'd17, 27'h00000067, 5'd3, 27'h0000002f, 5'd19, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000032b, 5'd0, 27'h00000361, 5'd29, 27'h000003f3, 32'h00000400,
  1'd1,  5'd16, 27'h00000089, 5'd13, 27'h0000010c, 5'd2, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000361, 5'd13, 27'h00000382, 5'd14, 27'h000001ee, 32'h00000400,
  1'd1,  5'd19, 27'h000000bf, 5'd13, 27'h000000fc, 5'd23, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ad, 5'd21, 27'h00000231, 5'd4, 27'h00000215, 32'h00000400,
  1'd1,  5'd16, 27'h000000e1, 5'd25, 27'h00000255, 5'd11, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001bc, 5'd21, 27'h0000013a, 5'd22, 27'h00000342, 32'h00000400,
  1'd1,  5'd27, 27'h000003cb, 5'd1, 27'h000001d4, 5'd1, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002e9, 5'd2, 27'h0000031f, 5'd10, 27'h000002c8, 32'h00000400,
  1'd1,  5'd29, 27'h000001a5, 5'd3, 27'h0000018f, 5'd23, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001ad, 5'd14, 27'h0000027c, 5'd1, 27'h0000029c, 32'h00000400,
  1'd1,  5'd27, 27'h00000165, 5'd13, 27'h0000038d, 5'd14, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000005e, 5'd14, 27'h00000376, 5'd21, 27'h000003c8, 32'h00000400,
  1'd1,  5'd29, 27'h00000055, 5'd24, 27'h00000060, 5'd4, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000001, 5'd22, 27'h0000031d, 5'd14, 27'h000003e4, 32'h00000400,
  1'd1,  5'd26, 27'h000000b3, 5'd25, 27'h0000023a, 5'd23, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000015d, 5'd0, 27'h000003a2, 5'd1, 27'h00000290, 32'h00000400,
  1'd1,  5'd6, 27'h0000004d, 5'd1, 27'h00000315, 5'd10, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000075, 5'd4, 27'h00000141, 5'd22, 27'h000001a7, 32'h00000400,
  1'd1,  5'd9, 27'h00000152, 5'd12, 27'h0000005c, 5'd9, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000143, 5'd13, 27'h00000064, 5'd17, 27'h000001f0, 32'h00000400,
  1'd1,  5'd7, 27'h000001ed, 5'd15, 27'h0000000e, 5'd30, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000014d, 5'd25, 27'h00000268, 5'd8, 27'h000001ae, 32'h00000400,
  1'd1,  5'd5, 27'h0000019a, 5'd23, 27'h00000042, 5'd16, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000310, 5'd24, 27'h00000166, 5'd26, 27'h0000030d, 32'h00000400,
  1'd1,  5'd15, 27'h00000283, 5'd2, 27'h000001ce, 5'd4, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000320, 5'd1, 27'h000002c1, 5'd12, 27'h00000196, 32'h00000400,
  1'd1,  5'd18, 27'h0000020a, 5'd1, 27'h00000340, 5'd22, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000030e, 5'd14, 27'h00000390, 5'd7, 27'h0000029e, 32'h00000400,
  1'd1,  5'd20, 27'h000001cb, 5'd15, 27'h000001d4, 5'd15, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000014a, 5'd14, 27'h00000189, 5'd30, 27'h0000008a, 32'h00000400,
  1'd1,  5'd16, 27'h00000373, 5'd20, 27'h000002fa, 5'd8, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000153, 5'd25, 27'h00000170, 5'd19, 27'h00000064, 32'h00000400,
  1'd1,  5'd17, 27'h00000299, 5'd24, 27'h00000118, 5'd28, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f3, 5'd2, 27'h0000036e, 5'd9, 27'h00000344, 32'h00000400,
  1'd1,  5'd27, 27'h00000274, 5'd0, 27'h00000185, 5'd19, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000398, 5'd3, 27'h00000227, 5'd27, 27'h000001af, 32'h00000400,
  1'd1,  5'd30, 27'h0000030a, 5'd13, 27'h000001cc, 5'd6, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b4, 5'd11, 27'h0000038b, 5'd15, 27'h00000333, 32'h00000400,
  1'd1,  5'd26, 27'h00000215, 5'd11, 27'h000003c2, 5'd27, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000030b, 5'd21, 27'h000000ab, 5'd5, 27'h000002c6, 32'h00000400,
  1'd1,  5'd30, 27'h00000165, 5'd23, 27'h000001fb, 5'd15, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000026f, 5'd23, 27'h0000027a, 5'd25, 27'h0000037f, 32'h00000400,
  1'd1,  5'd5, 27'h000000bd, 5'd6, 27'h000002df, 5'd1, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000027e, 5'd6, 27'h00000227, 5'd10, 27'h00000350, 32'h00000400,
  1'd1,  5'd7, 27'h000003f0, 5'd9, 27'h00000315, 5'd24, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ba, 5'd17, 27'h00000015, 5'd2, 27'h00000142, 32'h00000400,
  1'd1,  5'd6, 27'h0000038e, 5'd19, 27'h000000d6, 5'd12, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000157, 5'd15, 27'h000003b8, 5'd24, 27'h00000156, 32'h00000400,
  1'd1,  5'd8, 27'h0000036a, 5'd26, 27'h00000057, 5'd2, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000091, 5'd27, 27'h000003ba, 5'd15, 27'h00000004, 32'h00000400,
  1'd1,  5'd8, 27'h0000024c, 5'd30, 27'h00000198, 5'd22, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000004f, 5'd7, 27'h00000115, 5'd1, 27'h000002e6, 32'h00000400,
  1'd1,  5'd17, 27'h0000018a, 5'd6, 27'h0000014b, 5'd14, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ee, 5'd9, 27'h000002af, 5'd22, 27'h00000232, 32'h00000400,
  1'd1,  5'd18, 27'h000003f4, 5'd15, 27'h0000030e, 5'd4, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000042, 5'd19, 27'h0000015f, 5'd12, 27'h00000132, 32'h00000400,
  1'd1,  5'd17, 27'h0000035f, 5'd18, 27'h000001f6, 5'd23, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ed, 5'd29, 27'h00000376, 5'd0, 27'h0000006d, 32'h00000400,
  1'd1,  5'd19, 27'h0000006c, 5'd27, 27'h0000012f, 5'd15, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000010c, 5'd29, 27'h000000c2, 5'd23, 27'h000000b2, 32'h00000400,
  1'd1,  5'd25, 27'h00000386, 5'd6, 27'h00000124, 5'd0, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000038e, 5'd7, 27'h000002f6, 5'd15, 27'h00000131, 32'h00000400,
  1'd1,  5'd28, 27'h000001ca, 5'd6, 27'h000000b0, 5'd24, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000390, 5'd17, 27'h00000335, 5'd3, 27'h00000081, 32'h00000400,
  1'd1,  5'd26, 27'h000003ab, 5'd19, 27'h00000122, 5'd14, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ab, 5'd18, 27'h0000000b, 5'd21, 27'h000002fd, 32'h00000400,
  1'd1,  5'd27, 27'h000003b2, 5'd26, 27'h000003bd, 5'd3, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000006b, 5'd28, 27'h00000233, 5'd11, 27'h000002ab, 32'h00000400,
  1'd1,  5'd30, 27'h00000053, 5'd28, 27'h00000206, 5'd20, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001ef, 5'd8, 27'h00000353, 5'd10, 27'h0000001c, 32'h00000400,
  1'd1,  5'd8, 27'h0000035a, 5'd5, 27'h000000c3, 5'd19, 27'h000002a9, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000032b, 5'd8, 27'h00000195, 5'd25, 27'h000003f8, 32'h00000400,
  1'd1,  5'd8, 27'h0000012d, 5'd19, 27'h00000170, 5'd8, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000022, 5'd20, 27'h000001d1, 5'd16, 27'h00000339, 32'h00000400,
  1'd1,  5'd9, 27'h00000237, 5'd17, 27'h000000ec, 5'd29, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000011b, 5'd28, 27'h000000ca, 5'd9, 27'h000000d5, 32'h00000400,
  1'd1,  5'd5, 27'h00000116, 5'd26, 27'h000003fe, 5'd18, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000033d, 5'd29, 27'h000000fa, 5'd29, 27'h000002b5, 32'h00000400,
  1'd1,  5'd16, 27'h000002fb, 5'd9, 27'h000001fd, 5'd6, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c8, 5'd10, 27'h00000022, 5'd20, 27'h00000278, 32'h00000400,
  1'd1,  5'd17, 27'h0000014a, 5'd7, 27'h000000c8, 5'd27, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001d8, 5'd17, 27'h000003b0, 5'd7, 27'h00000178, 32'h00000400,
  1'd1,  5'd18, 27'h00000198, 5'd16, 27'h000002ff, 5'd15, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000294, 5'd16, 27'h0000007e, 5'd26, 27'h00000277, 32'h00000400,
  1'd1,  5'd18, 27'h00000327, 5'd26, 27'h0000009f, 5'd6, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003dd, 5'd29, 27'h000003a1, 5'd15, 27'h0000036e, 32'h00000400,
  1'd1,  5'd16, 27'h000002e7, 5'd30, 27'h0000018e, 5'd27, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000015, 5'd5, 27'h000003f3, 5'd6, 27'h0000033f, 32'h00000400,
  1'd1,  5'd30, 27'h000003db, 5'd9, 27'h00000365, 5'd19, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000018d, 5'd8, 27'h000001ce, 5'd27, 27'h0000009a, 32'h00000400,
  1'd1,  5'd30, 27'h000000df, 5'd18, 27'h00000075, 5'd7, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001cf, 5'd20, 27'h000000da, 5'd18, 27'h000003b0, 32'h00000400,
  1'd1,  5'd27, 27'h00000018, 5'd17, 27'h000000d2, 5'd27, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003b9, 5'd28, 27'h0000025a, 5'd6, 27'h000002d9, 32'h00000400,
  1'd1,  5'd29, 27'h0000027c, 5'd29, 27'h00000315, 5'd17, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c6, 5'd28, 27'h00000013, 5'd29, 27'h000002dd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000125, 5'd0, 27'h00000066, 5'd4, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e7, 5'd4, 27'h00000251, 5'd12, 27'h00000102, 32'h00000400,
  1'd1,  5'd4, 27'h000001c5, 5'd4, 27'h000001ba, 5'd25, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000129, 5'd12, 27'h000001f9, 5'd1, 27'h00000193, 32'h00000400,
  1'd1,  5'd2, 27'h0000006c, 5'd14, 27'h0000015d, 5'd13, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000015, 5'd13, 27'h000003f6, 5'd21, 27'h000003b6, 32'h00000400,
  1'd1,  5'd0, 27'h000000ee, 5'd24, 27'h00000361, 5'd0, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000335, 5'd24, 27'h00000095, 5'd14, 27'h000002e7, 32'h00000400,
  1'd1,  5'd0, 27'h00000025, 5'd24, 27'h0000033c, 5'd24, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c9, 5'd3, 27'h00000108, 5'd3, 27'h000001cb, 32'h00000400,
  1'd1,  5'd12, 27'h00000120, 5'd2, 27'h000000df, 5'd11, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001a3, 5'd0, 27'h00000337, 5'd22, 27'h000003aa, 32'h00000400,
  1'd1,  5'd11, 27'h0000033d, 5'd15, 27'h000000f6, 5'd3, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000234, 5'd12, 27'h00000114, 5'd13, 27'h0000012e, 32'h00000400,
  1'd1,  5'd11, 27'h0000034f, 5'd14, 27'h000000af, 5'd21, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013d, 5'd20, 27'h000002bb, 5'd2, 27'h00000139, 32'h00000400,
  1'd1,  5'd11, 27'h00000225, 5'd25, 27'h000000c7, 5'd10, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000094, 5'd23, 27'h0000039c, 5'd22, 27'h0000006f, 32'h00000400,
  1'd1,  5'd21, 27'h000003d3, 5'd0, 27'h000000ab, 5'd0, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002de, 5'd1, 27'h000002f5, 5'd12, 27'h00000250, 32'h00000400,
  1'd1,  5'd21, 27'h00000066, 5'd0, 27'h000003f4, 5'd24, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000052, 5'd13, 27'h000002b0, 5'd3, 27'h00000076, 32'h00000400,
  1'd1,  5'd20, 27'h000002ca, 5'd12, 27'h000003c4, 5'd14, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000020f, 5'd10, 27'h00000192, 5'd23, 27'h000001bb, 32'h00000400,
  1'd1,  5'd24, 27'h000003cd, 5'd24, 27'h0000025b, 5'd1, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000092, 5'd22, 27'h0000019c, 5'd14, 27'h00000266, 32'h00000400,
  1'd1,  5'd25, 27'h000000b9, 5'd24, 27'h000001e5, 5'd23, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000171, 5'd4, 27'h0000034a, 5'd8, 27'h0000035b, 32'h00000400,
  1'd1,  5'd3, 27'h00000018, 5'd1, 27'h000003a7, 5'd20, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002e2, 5'd3, 27'h00000132, 5'd27, 27'h00000064, 32'h00000400,
  1'd1,  5'd0, 27'h0000018a, 5'd10, 27'h000002b3, 5'd6, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000030d, 5'd15, 27'h0000017f, 5'd19, 27'h000003cf, 32'h00000400,
  1'd1,  5'd3, 27'h00000100, 5'd13, 27'h000003c6, 5'd29, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000011f, 5'd24, 27'h000002b1, 5'd8, 27'h000003a1, 32'h00000400,
  1'd1,  5'd1, 27'h000000ee, 5'd24, 27'h00000350, 5'd17, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000129, 5'd24, 27'h00000097, 5'd30, 27'h0000018b, 32'h00000400,
  1'd1,  5'd13, 27'h0000022b, 5'd1, 27'h000003fc, 5'd8, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000026e, 5'd0, 27'h00000296, 5'd17, 27'h000002c9, 32'h00000400,
  1'd1,  5'd12, 27'h000001e8, 5'd0, 27'h00000340, 5'd28, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035b, 5'd13, 27'h0000039e, 5'd8, 27'h0000008e, 32'h00000400,
  1'd1,  5'd11, 27'h000001c8, 5'd10, 27'h000003bc, 5'd16, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000105, 5'd12, 27'h000002d5, 5'd27, 27'h000002ae, 32'h00000400,
  1'd1,  5'd13, 27'h0000030a, 5'd21, 27'h00000389, 5'd5, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000019c, 5'd21, 27'h0000036d, 5'd16, 27'h000002d0, 32'h00000400,
  1'd1,  5'd14, 27'h00000143, 5'd25, 27'h0000007f, 5'd27, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a8, 5'd4, 27'h00000152, 5'd9, 27'h000003af, 32'h00000400,
  1'd1,  5'd21, 27'h000001c9, 5'd2, 27'h0000024b, 5'd18, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ce, 5'd3, 27'h0000016d, 5'd29, 27'h000002e9, 32'h00000400,
  1'd1,  5'd25, 27'h00000229, 5'd11, 27'h000003dc, 5'd7, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000324, 5'd13, 27'h000003d5, 5'd18, 27'h000000fd, 32'h00000400,
  1'd1,  5'd25, 27'h0000011b, 5'd11, 27'h0000027f, 5'd30, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000018e, 5'd24, 27'h00000080, 5'd9, 27'h000001f5, 32'h00000400,
  1'd1,  5'd24, 27'h000002cc, 5'd21, 27'h000002b2, 5'd19, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a5, 5'd23, 27'h0000028d, 5'd27, 27'h00000280, 32'h00000400,
  1'd1,  5'd1, 27'h00000299, 5'd8, 27'h00000143, 5'd1, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ba, 5'd9, 27'h000002b2, 5'd15, 27'h0000012c, 32'h00000400,
  1'd1,  5'd1, 27'h000001b1, 5'd7, 27'h00000123, 5'd21, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000009e, 5'd19, 27'h000000b1, 5'd0, 27'h00000249, 32'h00000400,
  1'd1,  5'd2, 27'h00000298, 5'd17, 27'h000002c2, 5'd12, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000019f, 5'd19, 27'h000002d5, 5'd24, 27'h0000004a, 32'h00000400,
  1'd1,  5'd3, 27'h00000266, 5'd30, 27'h0000016c, 5'd0, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000000a, 5'd26, 27'h000002ba, 5'd10, 27'h00000168, 32'h00000400,
  1'd1,  5'd5, 27'h00000033, 5'd29, 27'h00000078, 5'd22, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029e, 5'd7, 27'h00000014, 5'd4, 27'h0000001e, 32'h00000400,
  1'd1,  5'd10, 27'h0000036b, 5'd5, 27'h00000297, 5'd10, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e6, 5'd8, 27'h00000230, 5'd25, 27'h0000022c, 32'h00000400,
  1'd1,  5'd10, 27'h000003e5, 5'd15, 27'h000002e8, 5'd2, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000032b, 5'd17, 27'h00000186, 5'd12, 27'h00000298, 32'h00000400,
  1'd1,  5'd14, 27'h00000331, 5'd20, 27'h0000023f, 5'd23, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000022b, 5'd26, 27'h000001c5, 5'd0, 27'h00000047, 32'h00000400,
  1'd1,  5'd12, 27'h000003bb, 5'd28, 27'h000002e4, 5'd11, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c2, 5'd30, 27'h00000243, 5'd21, 27'h00000395, 32'h00000400,
  1'd1,  5'd24, 27'h00000080, 5'd7, 27'h00000085, 5'd0, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000029a, 5'd8, 27'h00000019, 5'd10, 27'h00000377, 32'h00000400,
  1'd1,  5'd23, 27'h000003da, 5'd7, 27'h00000162, 5'd24, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000fb, 5'd17, 27'h000001f7, 5'd3, 27'h000003cd, 32'h00000400,
  1'd1,  5'd23, 27'h000003dd, 5'd18, 27'h000003fb, 5'd10, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000219, 5'd19, 27'h0000023b, 5'd21, 27'h000003e2, 32'h00000400,
  1'd1,  5'd24, 27'h0000013e, 5'd29, 27'h00000156, 5'd2, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000bb, 5'd29, 27'h00000150, 5'd13, 27'h00000033, 32'h00000400,
  1'd1,  5'd24, 27'h0000016b, 5'd28, 27'h0000000c, 5'd22, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000144, 5'd6, 27'h00000164, 5'd6, 27'h0000037f, 32'h00000400,
  1'd1,  5'd1, 27'h000000c4, 5'd8, 27'h000003b7, 5'd17, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000376, 5'd5, 27'h00000361, 5'd27, 27'h0000022c, 32'h00000400,
  1'd1,  5'd3, 27'h00000218, 5'd15, 27'h00000210, 5'd6, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000144, 5'd17, 27'h00000398, 5'd16, 27'h000000f5, 32'h00000400,
  1'd1,  5'd4, 27'h00000011, 5'd17, 27'h00000331, 5'd29, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000286, 5'd29, 27'h000001b1, 5'd5, 27'h00000333, 32'h00000400,
  1'd1,  5'd4, 27'h0000031e, 5'd28, 27'h00000201, 5'd17, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000007e, 5'd29, 27'h00000132, 5'd26, 27'h0000009c, 32'h00000400,
  1'd1,  5'd14, 27'h0000005d, 5'd5, 27'h000000e7, 5'd5, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000015b, 5'd6, 27'h000000ff, 5'd19, 27'h00000312, 32'h00000400,
  1'd1,  5'd12, 27'h00000019, 5'd5, 27'h00000330, 5'd28, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000245, 5'd17, 27'h0000007d, 5'd6, 27'h00000350, 32'h00000400,
  1'd1,  5'd13, 27'h0000019d, 5'd20, 27'h00000075, 5'd17, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000017b, 5'd18, 27'h000002a5, 5'd26, 27'h000001be, 32'h00000400,
  1'd1,  5'd10, 27'h000003d7, 5'd27, 27'h000000ca, 5'd9, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000003e, 5'd29, 27'h00000366, 5'd16, 27'h00000266, 32'h00000400,
  1'd1,  5'd15, 27'h000000ec, 5'd28, 27'h000000ca, 5'd26, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000018f, 5'd7, 27'h0000035f, 5'd6, 27'h000003ad, 32'h00000400,
  1'd1,  5'd20, 27'h0000038f, 5'd5, 27'h0000024c, 5'd15, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000024e, 5'd6, 27'h00000152, 5'd27, 27'h000003c4, 32'h00000400,
  1'd1,  5'd23, 27'h00000254, 5'd17, 27'h0000038c, 5'd7, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000364, 5'd17, 27'h00000072, 5'd20, 27'h00000069, 32'h00000400,
  1'd1,  5'd21, 27'h00000296, 5'd19, 27'h0000012c, 5'd29, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000030f, 5'd26, 27'h000003b5, 5'd10, 27'h000000a6, 32'h00000400,
  1'd1,  5'd21, 27'h00000318, 5'd27, 27'h000003cb, 5'd17, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000304, 5'd30, 27'h000000c6, 5'd30, 27'h00000342, 32'h00000400,
  1'd1,  5'd8, 27'h00000298, 5'd0, 27'h000000fe, 5'd7, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000031a, 5'd4, 27'h00000387, 5'd19, 27'h00000350, 32'h00000400,
  1'd1,  5'd5, 27'h00000228, 5'd2, 27'h0000012d, 5'd28, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000395, 5'd13, 27'h000003f0, 5'd4, 27'h000003cb, 32'h00000400,
  1'd1,  5'd6, 27'h000002bc, 5'd11, 27'h00000109, 5'd11, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f7, 5'd12, 27'h0000013e, 5'd24, 27'h00000200, 32'h00000400,
  1'd1,  5'd5, 27'h00000362, 5'd24, 27'h000003ec, 5'd3, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000016c, 5'd25, 27'h00000315, 5'd11, 27'h0000037a, 32'h00000400,
  1'd1,  5'd9, 27'h0000008c, 5'd20, 27'h00000386, 5'd24, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000133, 5'd3, 27'h0000036a, 5'd9, 27'h00000122, 32'h00000400,
  1'd1,  5'd20, 27'h0000010e, 5'd4, 27'h00000148, 5'd19, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000032c, 5'd2, 27'h00000169, 5'd29, 27'h00000172, 32'h00000400,
  1'd1,  5'd19, 27'h000001bb, 5'd11, 27'h000000d0, 5'd2, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009c, 5'd14, 27'h00000198, 5'd10, 27'h00000194, 32'h00000400,
  1'd1,  5'd16, 27'h00000355, 5'd13, 27'h000001fe, 5'd24, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000013e, 5'd24, 27'h0000025d, 5'd2, 27'h0000015d, 32'h00000400,
  1'd1,  5'd16, 27'h000003a2, 5'd22, 27'h00000111, 5'd14, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ac, 5'd25, 27'h0000028e, 5'd24, 27'h000000f6, 32'h00000400,
  1'd1,  5'd29, 27'h0000006a, 5'd2, 27'h000002b0, 5'd2, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000043, 5'd4, 27'h00000048, 5'd11, 27'h00000099, 32'h00000400,
  1'd1,  5'd27, 27'h00000297, 5'd4, 27'h000002a0, 5'd25, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006f, 5'd10, 27'h00000177, 5'd3, 27'h00000336, 32'h00000400,
  1'd1,  5'd29, 27'h000003a1, 5'd15, 27'h00000194, 5'd11, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003b8, 5'd11, 27'h00000277, 5'd23, 27'h0000003d, 32'h00000400,
  1'd1,  5'd30, 27'h00000398, 5'd23, 27'h000001f8, 5'd1, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c0, 5'd23, 27'h00000079, 5'd14, 27'h000001bd, 32'h00000400,
  1'd1,  5'd26, 27'h00000079, 5'd22, 27'h000001b1, 5'd22, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000009e, 5'd0, 27'h00000208, 5'd1, 27'h0000000f, 32'h00000400,
  1'd1,  5'd5, 27'h000002f8, 5'd3, 27'h0000016d, 5'd12, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000319, 5'd4, 27'h0000008f, 5'd24, 27'h000002c0, 32'h00000400,
  1'd1,  5'd9, 27'h0000021b, 5'd11, 27'h00000279, 5'd8, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000182, 5'd14, 27'h0000022d, 5'd15, 27'h00000227, 32'h00000400,
  1'd1,  5'd7, 27'h00000356, 5'd12, 27'h00000246, 5'd28, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000025c, 5'd22, 27'h0000012c, 5'd10, 27'h00000010, 32'h00000400,
  1'd1,  5'd8, 27'h00000101, 5'd22, 27'h000002cd, 5'd16, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000247, 5'd24, 27'h00000141, 5'd28, 27'h0000025d, 32'h00000400,
  1'd1,  5'd18, 27'h000000d6, 5'd2, 27'h000001dc, 5'd4, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003cb, 5'd0, 27'h00000122, 5'd11, 27'h00000226, 32'h00000400,
  1'd1,  5'd17, 27'h0000038a, 5'd4, 27'h000001dc, 5'd23, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000101, 5'd13, 27'h000000c0, 5'd6, 27'h00000082, 32'h00000400,
  1'd1,  5'd19, 27'h000000d3, 5'd11, 27'h00000212, 5'd17, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000dc, 5'd14, 27'h000000de, 5'd27, 27'h000000a0, 32'h00000400,
  1'd1,  5'd17, 27'h000001f3, 5'd23, 27'h0000016c, 5'd7, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000020a, 5'd25, 27'h0000003c, 5'd17, 27'h000003ac, 32'h00000400,
  1'd1,  5'd18, 27'h0000028c, 5'd22, 27'h0000003b, 5'd26, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a0, 5'd4, 27'h0000010e, 5'd6, 27'h00000272, 32'h00000400,
  1'd1,  5'd30, 27'h00000287, 5'd2, 27'h000003a3, 5'd18, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000023f, 5'd1, 27'h00000115, 5'd28, 27'h000003f9, 32'h00000400,
  1'd1,  5'd26, 27'h0000029e, 5'd11, 27'h000002a1, 5'd7, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ac, 5'd10, 27'h000002ab, 5'd15, 27'h0000023c, 32'h00000400,
  1'd1,  5'd28, 27'h0000024c, 5'd14, 27'h0000038d, 5'd26, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002eb, 5'd21, 27'h0000013c, 5'd6, 27'h000002f6, 32'h00000400,
  1'd1,  5'd28, 27'h00000132, 5'd22, 27'h00000163, 5'd16, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000076, 5'd23, 27'h00000317, 5'd26, 27'h000002d7, 32'h00000400,
  1'd1,  5'd8, 27'h00000376, 5'd6, 27'h000000d6, 5'd0, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003b4, 5'd7, 27'h00000338, 5'd14, 27'h00000354, 32'h00000400,
  1'd1,  5'd8, 27'h000001e9, 5'd6, 27'h00000090, 5'd25, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000037, 5'd18, 27'h0000031e, 5'd2, 27'h00000014, 32'h00000400,
  1'd1,  5'd9, 27'h000000c4, 5'd17, 27'h000000d6, 5'd15, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000027e, 5'd19, 27'h00000080, 5'd25, 27'h0000011f, 32'h00000400,
  1'd1,  5'd9, 27'h0000038c, 5'd27, 27'h0000006e, 5'd3, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000379, 5'd26, 27'h000001bc, 5'd11, 27'h000003dd, 32'h00000400,
  1'd1,  5'd8, 27'h0000023c, 5'd29, 27'h000002bf, 5'd23, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000384, 5'd8, 27'h000001f0, 5'd3, 27'h000002df, 32'h00000400,
  1'd1,  5'd20, 27'h0000022c, 5'd7, 27'h00000231, 5'd13, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000372, 5'd8, 27'h0000031c, 5'd22, 27'h00000016, 32'h00000400,
  1'd1,  5'd17, 27'h00000319, 5'd18, 27'h000001d6, 5'd2, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030b, 5'd16, 27'h0000031b, 5'd11, 27'h00000233, 32'h00000400,
  1'd1,  5'd19, 27'h00000366, 5'd16, 27'h0000016d, 5'd25, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000030, 5'd27, 27'h0000012c, 5'd1, 27'h000002b1, 32'h00000400,
  1'd1,  5'd20, 27'h0000019c, 5'd30, 27'h00000046, 5'd13, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000221, 5'd29, 27'h000000d3, 5'd21, 27'h0000007c, 32'h00000400,
  1'd1,  5'd26, 27'h00000189, 5'd6, 27'h000003ee, 5'd2, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b8, 5'd7, 27'h0000020a, 5'd10, 27'h0000032c, 32'h00000400,
  1'd1,  5'd29, 27'h000003f9, 5'd7, 27'h0000004f, 5'd20, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003cf, 5'd19, 27'h0000037f, 5'd3, 27'h000000cd, 32'h00000400,
  1'd1,  5'd29, 27'h0000001f, 5'd16, 27'h0000024a, 5'd12, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001e8, 5'd19, 27'h00000218, 5'd24, 27'h00000230, 32'h00000400,
  1'd1,  5'd28, 27'h00000337, 5'd28, 27'h00000170, 5'd1, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000023c, 5'd30, 27'h0000038f, 5'd14, 27'h0000019f, 32'h00000400,
  1'd1,  5'd27, 27'h000000d9, 5'd25, 27'h0000036f, 5'd23, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000249, 5'd8, 27'h0000037f, 5'd6, 27'h000003d8, 32'h00000400,
  1'd1,  5'd9, 27'h000002fd, 5'd7, 27'h000000e4, 5'd18, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000010e, 5'd9, 27'h000003ce, 5'd28, 27'h0000023b, 32'h00000400,
  1'd1,  5'd9, 27'h00000274, 5'd19, 27'h000001c3, 5'd5, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000184, 5'd16, 27'h0000013e, 5'd19, 27'h000003be, 32'h00000400,
  1'd1,  5'd8, 27'h000002cf, 5'd19, 27'h00000036, 5'd30, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001d1, 5'd29, 27'h00000135, 5'd7, 27'h0000025c, 32'h00000400,
  1'd1,  5'd6, 27'h0000016e, 5'd28, 27'h0000014d, 5'd17, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000024a, 5'd27, 27'h0000007b, 5'd27, 27'h00000348, 32'h00000400,
  1'd1,  5'd16, 27'h0000025f, 5'd5, 27'h00000291, 5'd7, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000021f, 5'd6, 27'h000003ac, 5'd20, 27'h0000012d, 32'h00000400,
  1'd1,  5'd17, 27'h0000002b, 5'd9, 27'h00000355, 5'd26, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000127, 5'd19, 27'h000003c3, 5'd5, 27'h000003bf, 32'h00000400,
  1'd1,  5'd19, 27'h000001a7, 5'd19, 27'h000000bb, 5'd15, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000141, 5'd16, 27'h000000a3, 5'd26, 27'h000002e8, 32'h00000400,
  1'd1,  5'd16, 27'h000003d8, 5'd30, 27'h000000e3, 5'd9, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002bf, 5'd30, 27'h000001e5, 5'd19, 27'h00000068, 32'h00000400,
  1'd1,  5'd16, 27'h000003d6, 5'd30, 27'h0000005a, 5'd26, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000013f, 5'd6, 27'h00000175, 5'd8, 27'h000000a2, 32'h00000400,
  1'd1,  5'd29, 27'h00000303, 5'd6, 27'h000002f8, 5'd16, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000273, 5'd6, 27'h000003e6, 5'd27, 27'h0000031c, 32'h00000400,
  1'd1,  5'd29, 27'h000001b6, 5'd17, 27'h00000324, 5'd9, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000342, 5'd17, 27'h0000021d, 5'd17, 27'h00000352, 32'h00000400,
  1'd1,  5'd26, 27'h00000018, 5'd16, 27'h00000312, 5'd28, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000303, 5'd30, 27'h000000fc, 5'd6, 27'h000001c0, 32'h00000400,
  1'd1,  5'd28, 27'h00000016, 5'd28, 27'h000000c0, 5'd17, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000025e, 5'd26, 27'h0000022e, 5'd26, 27'h0000031b, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h00000013, 5'd0, 27'h00000126, 5'd1, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000c5, 5'd4, 27'h000002a9, 5'd10, 27'h00000193, 32'h00000400,
  1'd1,  5'd0, 27'h00000003, 5'd5, 27'h00000079, 5'd21, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000031f, 5'd13, 27'h00000058, 5'd0, 27'h000003f3, 32'h00000400,
  1'd1,  5'd3, 27'h000001fc, 5'd12, 27'h000001ad, 5'd15, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000268, 5'd14, 27'h000000bb, 5'd22, 27'h00000391, 32'h00000400,
  1'd1,  5'd1, 27'h000003c5, 5'd24, 27'h00000174, 5'd4, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000152, 5'd23, 27'h000001a7, 5'd12, 27'h0000019a, 32'h00000400,
  1'd1,  5'd2, 27'h000001cc, 5'd22, 27'h00000343, 5'd24, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a2, 5'd0, 27'h00000176, 5'd1, 27'h0000034c, 32'h00000400,
  1'd1,  5'd12, 27'h00000399, 5'd0, 27'h00000248, 5'd12, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000397, 5'd3, 27'h000001da, 5'd23, 27'h00000339, 32'h00000400,
  1'd1,  5'd13, 27'h000003be, 5'd15, 27'h00000114, 5'd2, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a0, 5'd13, 27'h00000262, 5'd15, 27'h00000120, 32'h00000400,
  1'd1,  5'd14, 27'h0000007b, 5'd14, 27'h000002bc, 5'd24, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e6, 5'd20, 27'h000002f2, 5'd0, 27'h00000218, 32'h00000400,
  1'd1,  5'd11, 27'h00000203, 5'd21, 27'h0000005e, 5'd10, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000fb, 5'd22, 27'h00000394, 5'd24, 27'h0000017d, 32'h00000400,
  1'd1,  5'd21, 27'h0000028a, 5'd4, 27'h00000286, 5'd2, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f8, 5'd0, 27'h00000258, 5'd11, 27'h0000038b, 32'h00000400,
  1'd1,  5'd23, 27'h00000220, 5'd3, 27'h000002aa, 5'd21, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000a0, 5'd15, 27'h0000006d, 5'd3, 27'h0000012a, 32'h00000400,
  1'd1,  5'd23, 27'h000000fb, 5'd11, 27'h00000357, 5'd11, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038f, 5'd10, 27'h0000028d, 5'd23, 27'h0000015d, 32'h00000400,
  1'd1,  5'd20, 27'h000003f5, 5'd25, 27'h00000019, 5'd4, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000008b, 5'd22, 27'h00000357, 5'd12, 27'h000003f4, 32'h00000400,
  1'd1,  5'd25, 27'h00000190, 5'd25, 27'h0000030e, 5'd23, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000007d, 5'd3, 27'h0000038e, 5'd7, 27'h000002bb, 32'h00000400,
  1'd1,  5'd2, 27'h00000348, 5'd4, 27'h00000008, 5'd18, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000233, 5'd0, 27'h000001b3, 5'd29, 27'h0000006d, 32'h00000400,
  1'd1,  5'd2, 27'h000001fc, 5'd14, 27'h000003e1, 5'd5, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000386, 5'd12, 27'h00000356, 5'd16, 27'h0000010c, 32'h00000400,
  1'd1,  5'd0, 27'h0000015e, 5'd11, 27'h000003b2, 5'd30, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e8, 5'd24, 27'h00000391, 5'd8, 27'h00000298, 32'h00000400,
  1'd1,  5'd1, 27'h0000018f, 5'd23, 27'h000000d0, 5'd19, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000037, 5'd22, 27'h000000c2, 5'd29, 27'h00000051, 32'h00000400,
  1'd1,  5'd12, 27'h00000029, 5'd1, 27'h000001a5, 5'd5, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c2, 5'd1, 27'h0000016e, 5'd15, 27'h000003b5, 32'h00000400,
  1'd1,  5'd13, 27'h0000001e, 5'd5, 27'h000000a0, 5'd28, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001ef, 5'd13, 27'h00000082, 5'd9, 27'h000002d2, 32'h00000400,
  1'd1,  5'd14, 27'h000001c2, 5'd14, 27'h000001d3, 5'd15, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000034, 5'd11, 27'h000002f9, 5'd25, 27'h000003a3, 32'h00000400,
  1'd1,  5'd10, 27'h00000280, 5'd23, 27'h000002f1, 5'd6, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000161, 5'd24, 27'h0000037f, 5'd17, 27'h000002b3, 32'h00000400,
  1'd1,  5'd13, 27'h0000013c, 5'd21, 27'h00000020, 5'd30, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c3, 5'd2, 27'h000001c7, 5'd10, 27'h00000084, 32'h00000400,
  1'd1,  5'd21, 27'h0000008b, 5'd4, 27'h0000010e, 5'd19, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000027, 5'd4, 27'h00000248, 5'd29, 27'h000003bd, 32'h00000400,
  1'd1,  5'd24, 27'h00000103, 5'd12, 27'h000003af, 5'd5, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000086, 5'd15, 27'h0000018f, 5'd19, 27'h000001c3, 32'h00000400,
  1'd1,  5'd24, 27'h000000ed, 5'd12, 27'h00000259, 5'd28, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000249, 5'd21, 27'h00000269, 5'd5, 27'h000002c2, 32'h00000400,
  1'd1,  5'd22, 27'h00000107, 5'd23, 27'h000003ad, 5'd16, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000235, 5'd22, 27'h000000ae, 5'd28, 27'h000001df, 32'h00000400,
  1'd1,  5'd0, 27'h000002a5, 5'd6, 27'h00000041, 5'd1, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003e2, 5'd6, 27'h000000ac, 5'd14, 27'h0000014d, 32'h00000400,
  1'd1,  5'd4, 27'h00000300, 5'd7, 27'h00000062, 5'd21, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e3, 5'd16, 27'h0000012e, 5'd1, 27'h0000029e, 32'h00000400,
  1'd1,  5'd1, 27'h000002b9, 5'd15, 27'h000002c7, 5'd13, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002e8, 5'd16, 27'h00000096, 5'd24, 27'h000001ef, 32'h00000400,
  1'd1,  5'd3, 27'h000002ae, 5'd29, 27'h000001a2, 5'd3, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000c0, 5'd26, 27'h000000c3, 5'd15, 27'h000000d3, 32'h00000400,
  1'd1,  5'd2, 27'h000001a0, 5'd27, 27'h0000011f, 5'd22, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000063, 5'd5, 27'h00000299, 5'd4, 27'h000000b6, 32'h00000400,
  1'd1,  5'd15, 27'h0000002a, 5'd9, 27'h000002c8, 5'd14, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000e3, 5'd10, 27'h00000109, 5'd21, 27'h0000006a, 32'h00000400,
  1'd1,  5'd13, 27'h0000023c, 5'd15, 27'h00000349, 5'd2, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ad, 5'd15, 27'h000003b8, 5'd14, 27'h00000111, 32'h00000400,
  1'd1,  5'd12, 27'h00000197, 5'd15, 27'h000003fb, 5'd24, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000da, 5'd26, 27'h00000008, 5'd4, 27'h00000105, 32'h00000400,
  1'd1,  5'd15, 27'h0000010b, 5'd28, 27'h000001ed, 5'd10, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d1, 5'd30, 27'h0000019c, 5'd21, 27'h0000008f, 32'h00000400,
  1'd1,  5'd25, 27'h0000011f, 5'd7, 27'h0000024f, 5'd5, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e4, 5'd6, 27'h0000017e, 5'd13, 27'h0000021a, 32'h00000400,
  1'd1,  5'd23, 27'h00000008, 5'd10, 27'h00000105, 5'd22, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c9, 5'd18, 27'h000003f4, 5'd2, 27'h000001ea, 32'h00000400,
  1'd1,  5'd22, 27'h00000069, 5'd15, 27'h0000031f, 5'd15, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000307, 5'd19, 27'h00000389, 5'd22, 27'h00000074, 32'h00000400,
  1'd1,  5'd21, 27'h00000055, 5'd29, 27'h0000023b, 5'd4, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000038, 5'd30, 27'h00000179, 5'd14, 27'h00000033, 32'h00000400,
  1'd1,  5'd20, 27'h00000392, 5'd28, 27'h00000039, 5'd24, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000356, 5'd7, 27'h0000000d, 5'd8, 27'h00000174, 32'h00000400,
  1'd1,  5'd1, 27'h000002ca, 5'd5, 27'h000002a0, 5'd17, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000245, 5'd5, 27'h00000270, 5'd26, 27'h00000314, 32'h00000400,
  1'd1,  5'd2, 27'h000003e5, 5'd19, 27'h00000012, 5'd7, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012c, 5'd16, 27'h00000203, 5'd20, 27'h00000108, 32'h00000400,
  1'd1,  5'd4, 27'h000003bb, 5'd19, 27'h00000097, 5'd28, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000021b, 5'd28, 27'h0000033f, 5'd6, 27'h00000111, 32'h00000400,
  1'd1,  5'd2, 27'h00000391, 5'd27, 27'h000003bc, 5'd16, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c3, 5'd27, 27'h00000316, 5'd27, 27'h0000009e, 32'h00000400,
  1'd1,  5'd10, 27'h00000305, 5'd9, 27'h00000067, 5'd9, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000050, 5'd8, 27'h00000160, 5'd19, 27'h000002e8, 32'h00000400,
  1'd1,  5'd12, 27'h000002bc, 5'd8, 27'h00000164, 5'd30, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000258, 5'd17, 27'h00000358, 5'd6, 27'h000002fe, 32'h00000400,
  1'd1,  5'd13, 27'h000002b0, 5'd18, 27'h00000303, 5'd20, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000351, 5'd17, 27'h00000042, 5'd30, 27'h0000018a, 32'h00000400,
  1'd1,  5'd14, 27'h000000ca, 5'd29, 27'h0000011c, 5'd5, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000372, 5'd27, 27'h00000100, 5'd15, 27'h000002d9, 32'h00000400,
  1'd1,  5'd14, 27'h0000001a, 5'd30, 27'h000001d1, 5'd26, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000023f, 5'd6, 27'h00000389, 5'd7, 27'h000002fa, 32'h00000400,
  1'd1,  5'd24, 27'h000001c9, 5'd9, 27'h00000371, 5'd18, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000017, 5'd7, 27'h00000030, 5'd27, 27'h00000380, 32'h00000400,
  1'd1,  5'd21, 27'h000003b1, 5'd20, 27'h00000173, 5'd7, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000142, 5'd19, 27'h00000284, 5'd16, 27'h00000305, 32'h00000400,
  1'd1,  5'd21, 27'h00000054, 5'd18, 27'h00000353, 5'd30, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001c9, 5'd26, 27'h0000027c, 5'd6, 27'h000000ff, 32'h00000400,
  1'd1,  5'd21, 27'h00000076, 5'd27, 27'h0000005c, 5'd17, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000035c, 5'd30, 27'h0000011c, 5'd28, 27'h000003f1, 32'h00000400,
  1'd1,  5'd6, 27'h000003f6, 5'd0, 27'h000003db, 5'd6, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c5, 5'd1, 27'h000001b9, 5'd16, 27'h00000057, 32'h00000400,
  1'd1,  5'd10, 27'h00000008, 5'd1, 27'h00000189, 5'd27, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000173, 5'd12, 27'h0000019b, 5'd2, 27'h00000253, 32'h00000400,
  1'd1,  5'd7, 27'h000002b7, 5'd15, 27'h000001ae, 5'd10, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ab, 5'd12, 27'h00000235, 5'd24, 27'h00000070, 32'h00000400,
  1'd1,  5'd8, 27'h000000e9, 5'd21, 27'h0000035d, 5'd1, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000008b, 5'd23, 27'h00000192, 5'd10, 27'h0000032b, 32'h00000400,
  1'd1,  5'd9, 27'h000001e4, 5'd24, 27'h000003af, 5'd25, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000f7, 5'd1, 27'h000002eb, 5'd7, 27'h000000cf, 32'h00000400,
  1'd1,  5'd17, 27'h00000373, 5'd2, 27'h000001c6, 5'd16, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006c, 5'd4, 27'h0000038c, 5'd28, 27'h00000272, 32'h00000400,
  1'd1,  5'd16, 27'h0000039c, 5'd13, 27'h0000036f, 5'd0, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000213, 5'd13, 27'h0000036a, 5'd13, 27'h00000083, 32'h00000400,
  1'd1,  5'd19, 27'h0000002e, 5'd12, 27'h00000238, 5'd23, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000dd, 5'd21, 27'h000001bb, 5'd1, 27'h0000037a, 32'h00000400,
  1'd1,  5'd20, 27'h000001fc, 5'd22, 27'h00000196, 5'd13, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000037d, 5'd22, 27'h0000012e, 5'd21, 27'h000000fc, 32'h00000400,
  1'd1,  5'd28, 27'h0000015c, 5'd2, 27'h0000022b, 5'd4, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000a4, 5'd5, 27'h00000008, 5'd13, 27'h000001b4, 32'h00000400,
  1'd1,  5'd29, 27'h00000217, 5'd2, 27'h00000101, 5'd21, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c6, 5'd14, 27'h000003a7, 5'd1, 27'h000001f0, 32'h00000400,
  1'd1,  5'd27, 27'h000000b7, 5'd11, 27'h00000246, 5'd14, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023b, 5'd15, 27'h00000031, 5'd23, 27'h000001b6, 32'h00000400,
  1'd1,  5'd28, 27'h00000293, 5'd21, 27'h000002d9, 5'd4, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000017a, 5'd22, 27'h0000032c, 5'd11, 27'h00000229, 32'h00000400,
  1'd1,  5'd27, 27'h00000075, 5'd21, 27'h0000016c, 5'd23, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021e, 5'd2, 27'h0000035a, 5'd3, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h00000017, 5'd3, 27'h000001b6, 5'd13, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000c2, 5'd3, 27'h00000112, 5'd25, 27'h00000313, 32'h00000400,
  1'd1,  5'd9, 27'h0000010e, 5'd13, 27'h000000e0, 5'd7, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e8, 5'd12, 27'h000001d8, 5'd16, 27'h00000271, 32'h00000400,
  1'd1,  5'd9, 27'h000003e0, 5'd10, 27'h000003c9, 5'd28, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005b, 5'd25, 27'h00000031, 5'd9, 27'h00000279, 32'h00000400,
  1'd1,  5'd9, 27'h000000bd, 5'd25, 27'h00000009, 5'd16, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002cc, 5'd24, 27'h00000355, 5'd29, 27'h00000298, 32'h00000400,
  1'd1,  5'd20, 27'h000001c1, 5'd3, 27'h00000359, 5'd2, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000234, 5'd0, 27'h0000039a, 5'd15, 27'h00000156, 32'h00000400,
  1'd1,  5'd16, 27'h000002f0, 5'd1, 27'h00000227, 5'd22, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000288, 5'd15, 27'h000001e9, 5'd10, 27'h0000002d, 32'h00000400,
  1'd1,  5'd16, 27'h000000af, 5'd12, 27'h0000030c, 5'd18, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a3, 5'd11, 27'h00000168, 5'd28, 27'h000003f0, 32'h00000400,
  1'd1,  5'd18, 27'h000001de, 5'd23, 27'h0000029a, 5'd5, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035c, 5'd22, 27'h00000197, 5'd20, 27'h00000186, 32'h00000400,
  1'd1,  5'd17, 27'h0000003d, 5'd25, 27'h00000098, 5'd30, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000017d, 5'd1, 27'h00000112, 5'd8, 27'h0000005d, 32'h00000400,
  1'd1,  5'd29, 27'h0000018e, 5'd3, 27'h00000202, 5'd18, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000193, 5'd2, 27'h0000002b, 5'd28, 27'h000002f2, 32'h00000400,
  1'd1,  5'd29, 27'h000000b1, 5'd14, 27'h00000392, 5'd7, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000378, 5'd15, 27'h000000da, 5'd20, 27'h0000024a, 32'h00000400,
  1'd1,  5'd27, 27'h000000df, 5'd13, 27'h00000050, 5'd29, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000308, 5'd24, 27'h000001cb, 5'd6, 27'h000001b1, 32'h00000400,
  1'd1,  5'd30, 27'h00000000, 5'd24, 27'h000001cd, 5'd19, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000123, 5'd22, 27'h00000067, 5'd27, 27'h00000381, 32'h00000400,
  1'd1,  5'd9, 27'h00000164, 5'd8, 27'h000003f1, 5'd3, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000221, 5'd5, 27'h00000210, 5'd11, 27'h000001af, 32'h00000400,
  1'd1,  5'd7, 27'h0000038d, 5'd7, 27'h00000280, 5'd24, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032b, 5'd16, 27'h00000191, 5'd2, 27'h0000009d, 32'h00000400,
  1'd1,  5'd9, 27'h0000019c, 5'd16, 27'h00000394, 5'd13, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000001, 5'd20, 27'h00000090, 5'd24, 27'h00000248, 32'h00000400,
  1'd1,  5'd6, 27'h0000011b, 5'd27, 27'h000003f6, 5'd4, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e0, 5'd28, 27'h000003af, 5'd11, 27'h00000024, 32'h00000400,
  1'd1,  5'd6, 27'h000003c5, 5'd28, 27'h00000025, 5'd21, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000292, 5'd5, 27'h000000cc, 5'd2, 27'h0000007d, 32'h00000400,
  1'd1,  5'd15, 27'h0000037e, 5'd9, 27'h000001fa, 5'd11, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000f8, 5'd9, 27'h0000015d, 5'd23, 27'h00000389, 32'h00000400,
  1'd1,  5'd20, 27'h00000125, 5'd18, 27'h000001e6, 5'd2, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d5, 5'd20, 27'h0000000b, 5'd10, 27'h000002b0, 32'h00000400,
  1'd1,  5'd19, 27'h00000235, 5'd19, 27'h000003d3, 5'd23, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d0, 5'd27, 27'h00000141, 5'd2, 27'h000000b9, 32'h00000400,
  1'd1,  5'd17, 27'h000001fd, 5'd30, 27'h000001b1, 5'd13, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000251, 5'd29, 27'h0000032a, 5'd22, 27'h0000028e, 32'h00000400,
  1'd1,  5'd30, 27'h00000228, 5'd6, 27'h000003dc, 5'd0, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000350, 5'd8, 27'h00000150, 5'd14, 27'h000000ff, 32'h00000400,
  1'd1,  5'd28, 27'h0000014f, 5'd5, 27'h000001ed, 5'd21, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b6, 5'd20, 27'h00000181, 5'd1, 27'h000003cc, 32'h00000400,
  1'd1,  5'd30, 27'h000001ab, 5'd20, 27'h0000004c, 5'd12, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000322, 5'd18, 27'h0000002f, 5'd24, 27'h0000018b, 32'h00000400,
  1'd1,  5'd26, 27'h000000ee, 5'd27, 27'h00000082, 5'd2, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000022c, 5'd27, 27'h000003f0, 5'd11, 27'h000003f2, 32'h00000400,
  1'd1,  5'd29, 27'h00000272, 5'd28, 27'h0000038d, 5'd23, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000028c, 5'd7, 27'h00000157, 5'd9, 27'h00000334, 32'h00000400,
  1'd1,  5'd7, 27'h000001d9, 5'd9, 27'h0000018c, 5'd18, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000185, 5'd8, 27'h00000264, 5'd27, 27'h0000027b, 32'h00000400,
  1'd1,  5'd5, 27'h00000318, 5'd20, 27'h00000069, 5'd7, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e1, 5'd19, 27'h000002ad, 5'd15, 27'h00000310, 32'h00000400,
  1'd1,  5'd9, 27'h000001f8, 5'd19, 27'h00000398, 5'd26, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000360, 5'd30, 27'h00000039, 5'd5, 27'h000000c4, 32'h00000400,
  1'd1,  5'd7, 27'h00000222, 5'd26, 27'h000000ed, 5'd18, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f2, 5'd27, 27'h000000ec, 5'd29, 27'h000000b2, 32'h00000400,
  1'd1,  5'd18, 27'h0000016d, 5'd10, 27'h0000004e, 5'd8, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000249, 5'd9, 27'h0000032a, 5'd17, 27'h0000002a, 32'h00000400,
  1'd1,  5'd18, 27'h0000038b, 5'd6, 27'h000003f6, 5'd29, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000029c, 5'd18, 27'h000000e8, 5'd6, 27'h00000134, 32'h00000400,
  1'd1,  5'd19, 27'h00000351, 5'd15, 27'h00000330, 5'd18, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b8, 5'd20, 27'h00000019, 5'd28, 27'h000001b5, 32'h00000400,
  1'd1,  5'd17, 27'h0000014d, 5'd26, 27'h0000021d, 5'd6, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000127, 5'd28, 27'h000003d8, 5'd18, 27'h00000343, 32'h00000400,
  1'd1,  5'd15, 27'h00000375, 5'd26, 27'h00000146, 5'd27, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000079, 5'd9, 27'h0000012f, 5'd5, 27'h00000326, 32'h00000400,
  1'd1,  5'd26, 27'h0000025e, 5'd7, 27'h0000023a, 5'd18, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001fd, 5'd9, 27'h0000020a, 5'd26, 27'h00000256, 32'h00000400,
  1'd1,  5'd28, 27'h00000005, 5'd16, 27'h00000205, 5'd10, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000357, 5'd18, 27'h00000120, 5'd16, 27'h000003b2, 32'h00000400,
  1'd1,  5'd29, 27'h000000a7, 5'd17, 27'h0000005e, 5'd27, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a6, 5'd29, 27'h00000099, 5'd6, 27'h000003ca, 32'h00000400,
  1'd1,  5'd29, 27'h000000ff, 5'd29, 27'h000002a6, 5'd17, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000005c, 5'd26, 27'h000002c3, 5'd30, 27'h00000352, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000002a4, 5'd4, 27'h000001a6, 5'd2, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000099, 5'd2, 27'h000003b7, 5'd15, 27'h00000071, 32'h00000400,
  1'd1,  5'd2, 27'h00000263, 5'd2, 27'h0000024b, 5'd23, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000f9, 5'd12, 27'h00000152, 5'd1, 27'h00000271, 32'h00000400,
  1'd1,  5'd2, 27'h000002a2, 5'd12, 27'h00000109, 5'd11, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000314, 5'd14, 27'h0000000c, 5'd21, 27'h000001a7, 32'h00000400,
  1'd1,  5'd4, 27'h00000037, 5'd21, 27'h000001bd, 5'd2, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000254, 5'd24, 27'h00000312, 5'd14, 27'h000003ca, 32'h00000400,
  1'd1,  5'd3, 27'h0000007a, 5'd21, 27'h00000222, 5'd23, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000039b, 5'd1, 27'h000000a3, 5'd2, 27'h000002ce, 32'h00000400,
  1'd1,  5'd13, 27'h0000033d, 5'd0, 27'h00000133, 5'd14, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003cd, 5'd1, 27'h0000003b, 5'd21, 27'h00000158, 32'h00000400,
  1'd1,  5'd12, 27'h00000279, 5'd13, 27'h000002b5, 5'd2, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000266, 5'd13, 27'h000000b6, 5'd14, 27'h000000a6, 32'h00000400,
  1'd1,  5'd14, 27'h0000029f, 5'd11, 27'h00000088, 5'd20, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d7, 5'd24, 27'h000003ae, 5'd2, 27'h0000005a, 32'h00000400,
  1'd1,  5'd13, 27'h0000037a, 5'd23, 27'h00000173, 5'd13, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e1, 5'd24, 27'h000001e2, 5'd24, 27'h00000320, 32'h00000400,
  1'd1,  5'd25, 27'h00000327, 5'd3, 27'h000001c8, 5'd2, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b7, 5'd1, 27'h000003ac, 5'd13, 27'h0000029f, 32'h00000400,
  1'd1,  5'd21, 27'h00000304, 5'd2, 27'h000001c9, 5'd24, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000032e, 5'd10, 27'h0000036e, 5'd5, 27'h0000007b, 32'h00000400,
  1'd1,  5'd25, 27'h00000262, 5'd13, 27'h00000127, 5'd10, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000126, 5'd10, 27'h000001e3, 5'd23, 27'h00000136, 32'h00000400,
  1'd1,  5'd24, 27'h0000028e, 5'd24, 27'h0000010f, 5'd3, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000019f, 5'd24, 27'h000001b6, 5'd15, 27'h00000022, 32'h00000400,
  1'd1,  5'd22, 27'h00000157, 5'd22, 27'h000002df, 5'd21, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001ef, 5'd1, 27'h000002af, 5'd8, 27'h000000a0, 32'h00000400,
  1'd1,  5'd1, 27'h00000070, 5'd2, 27'h0000014c, 5'd18, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000391, 5'd4, 27'h000002e4, 5'd29, 27'h00000261, 32'h00000400,
  1'd1,  5'd2, 27'h000002ee, 5'd11, 27'h000000ae, 5'd7, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002e1, 5'd13, 27'h0000034e, 5'd16, 27'h00000118, 32'h00000400,
  1'd1,  5'd3, 27'h000003c8, 5'd12, 27'h0000007b, 5'd29, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014c, 5'd24, 27'h000001fe, 5'd8, 27'h0000003c, 32'h00000400,
  1'd1,  5'd3, 27'h000001dc, 5'd22, 27'h00000203, 5'd17, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001b4, 5'd20, 27'h00000386, 5'd30, 27'h00000097, 32'h00000400,
  1'd1,  5'd14, 27'h000000c3, 5'd1, 27'h00000184, 5'd8, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000063, 5'd2, 27'h0000002b, 5'd16, 27'h00000355, 32'h00000400,
  1'd1,  5'd12, 27'h000001ae, 5'd4, 27'h00000265, 5'd29, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000171, 5'd13, 27'h00000300, 5'd5, 27'h000003a8, 32'h00000400,
  1'd1,  5'd15, 27'h0000005f, 5'd14, 27'h00000329, 5'd16, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000299, 5'd11, 27'h00000058, 5'd30, 27'h0000020c, 32'h00000400,
  1'd1,  5'd12, 27'h0000005f, 5'd22, 27'h00000020, 5'd5, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ed, 5'd24, 27'h00000321, 5'd17, 27'h0000004c, 32'h00000400,
  1'd1,  5'd15, 27'h000001ca, 5'd25, 27'h0000030f, 5'd30, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000374, 5'd4, 27'h000002e1, 5'd8, 27'h000000a4, 32'h00000400,
  1'd1,  5'd24, 27'h000000fc, 5'd1, 27'h0000001d, 5'd15, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000060, 5'd1, 27'h00000029, 5'd27, 27'h000000ed, 32'h00000400,
  1'd1,  5'd23, 27'h000002a1, 5'd10, 27'h0000039b, 5'd8, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e4, 5'd12, 27'h000002c2, 5'd17, 27'h0000014f, 32'h00000400,
  1'd1,  5'd24, 27'h00000214, 5'd13, 27'h0000017d, 5'd30, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001a1, 5'd22, 27'h00000266, 5'd7, 27'h000000d7, 32'h00000400,
  1'd1,  5'd23, 27'h0000035d, 5'd20, 27'h000003e9, 5'd18, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022f, 5'd23, 27'h000003a4, 5'd29, 27'h00000080, 32'h00000400,
  1'd1,  5'd4, 27'h0000021b, 5'd7, 27'h0000037f, 5'd4, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000004d, 5'd10, 27'h00000109, 5'd15, 27'h0000011f, 32'h00000400,
  1'd1,  5'd4, 27'h00000250, 5'd8, 27'h0000020b, 5'd22, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000010f, 5'd15, 27'h00000354, 5'd3, 27'h000000c2, 32'h00000400,
  1'd1,  5'd0, 27'h000002f6, 5'd17, 27'h00000140, 5'd13, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000018b, 5'd19, 27'h00000307, 5'd25, 27'h0000001b, 32'h00000400,
  1'd1,  5'd3, 27'h000001a4, 5'd28, 27'h00000197, 5'd2, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000c6, 5'd29, 27'h000001eb, 5'd10, 27'h000003ab, 32'h00000400,
  1'd1,  5'd3, 27'h000001be, 5'd30, 27'h00000162, 5'd20, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000120, 5'd7, 27'h000001ad, 5'd3, 27'h000001b7, 32'h00000400,
  1'd1,  5'd11, 27'h000002ee, 5'd7, 27'h000000a0, 5'd12, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000289, 5'd5, 27'h0000029b, 5'd25, 27'h00000007, 32'h00000400,
  1'd1,  5'd10, 27'h000002c6, 5'd17, 27'h0000038a, 5'd2, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000393, 5'd20, 27'h000001b4, 5'd11, 27'h00000196, 32'h00000400,
  1'd1,  5'd11, 27'h000002c5, 5'd18, 27'h00000250, 5'd22, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001af, 5'd28, 27'h00000235, 5'd2, 27'h000003b8, 32'h00000400,
  1'd1,  5'd12, 27'h000003b3, 5'd30, 27'h00000058, 5'd12, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000186, 5'd27, 27'h0000032c, 5'd22, 27'h00000322, 32'h00000400,
  1'd1,  5'd22, 27'h000002fe, 5'd9, 27'h0000013c, 5'd3, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000013c, 5'd8, 27'h0000004f, 5'd11, 27'h000003aa, 32'h00000400,
  1'd1,  5'd22, 27'h0000011f, 5'd5, 27'h000003ec, 5'd23, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000068, 5'd20, 27'h0000023c, 5'd2, 27'h00000203, 32'h00000400,
  1'd1,  5'd23, 27'h000001cf, 5'd15, 27'h00000375, 5'd13, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000000c, 5'd15, 27'h000003cb, 5'd25, 27'h00000057, 32'h00000400,
  1'd1,  5'd21, 27'h00000370, 5'd27, 27'h000003d3, 5'd2, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001c5, 5'd27, 27'h000000ea, 5'd13, 27'h000001d2, 32'h00000400,
  1'd1,  5'd20, 27'h0000033b, 5'd29, 27'h00000122, 5'd22, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039b, 5'd8, 27'h0000001d, 5'd6, 27'h000003fc, 32'h00000400,
  1'd1,  5'd1, 27'h0000038d, 5'd7, 27'h0000018d, 5'd16, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000378, 5'd7, 27'h000001bf, 5'd27, 27'h00000383, 32'h00000400,
  1'd1,  5'd3, 27'h00000199, 5'd20, 27'h00000254, 5'd9, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001dc, 5'd18, 27'h00000204, 5'd19, 27'h000000df, 32'h00000400,
  1'd1,  5'd4, 27'h00000360, 5'd17, 27'h000002d8, 5'd26, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000167, 5'd27, 27'h00000118, 5'd7, 27'h00000305, 32'h00000400,
  1'd1,  5'd4, 27'h000001ab, 5'd25, 27'h0000035b, 5'd16, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000095, 5'd29, 27'h00000172, 5'd30, 27'h000000f0, 32'h00000400,
  1'd1,  5'd10, 27'h000003cb, 5'd6, 27'h00000291, 5'd7, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f5, 5'd7, 27'h00000389, 5'd18, 27'h00000282, 32'h00000400,
  1'd1,  5'd14, 27'h000003e8, 5'd9, 27'h00000332, 5'd27, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000001, 5'd20, 27'h0000008e, 5'd8, 27'h000002f7, 32'h00000400,
  1'd1,  5'd11, 27'h0000023b, 5'd17, 27'h00000147, 5'd19, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000fe, 5'd20, 27'h00000154, 5'd30, 27'h0000026b, 32'h00000400,
  1'd1,  5'd14, 27'h000000a3, 5'd27, 27'h00000166, 5'd8, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000031e, 5'd27, 27'h0000031e, 5'd16, 27'h0000022c, 32'h00000400,
  1'd1,  5'd11, 27'h00000127, 5'd29, 27'h000000ad, 5'd30, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002bb, 5'd7, 27'h00000307, 5'd7, 27'h00000382, 32'h00000400,
  1'd1,  5'd21, 27'h00000284, 5'd8, 27'h0000023f, 5'd19, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ee, 5'd7, 27'h0000014a, 5'd27, 27'h000000d6, 32'h00000400,
  1'd1,  5'd23, 27'h000003cf, 5'd18, 27'h000001c7, 5'd5, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000186, 5'd18, 27'h00000002, 5'd15, 27'h00000207, 32'h00000400,
  1'd1,  5'd24, 27'h000002b0, 5'd15, 27'h00000230, 5'd26, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000099, 5'd30, 27'h00000226, 5'd9, 27'h000003f6, 32'h00000400,
  1'd1,  5'd21, 27'h000000a5, 5'd30, 27'h00000065, 5'd18, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a9, 5'd30, 27'h00000317, 5'd28, 27'h00000311, 32'h00000400,
  1'd1,  5'd5, 27'h00000182, 5'd0, 27'h00000217, 5'd5, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000d, 5'd2, 27'h00000336, 5'd19, 27'h0000003b, 32'h00000400,
  1'd1,  5'd7, 27'h000000bf, 5'd2, 27'h000000ac, 5'd30, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000030d, 5'd10, 27'h000003de, 5'd1, 27'h0000038f, 32'h00000400,
  1'd1,  5'd9, 27'h000002c7, 5'd12, 27'h000002e9, 5'd13, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003b3, 5'd14, 27'h000000d4, 5'd22, 27'h0000025d, 32'h00000400,
  1'd1,  5'd7, 27'h00000329, 5'd24, 27'h0000020f, 5'd5, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000322, 5'd20, 27'h00000334, 5'd13, 27'h00000006, 32'h00000400,
  1'd1,  5'd6, 27'h00000326, 5'd22, 27'h00000153, 5'd23, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000373, 5'd1, 27'h000000eb, 5'd6, 27'h00000086, 32'h00000400,
  1'd1,  5'd19, 27'h00000335, 5'd2, 27'h00000355, 5'd19, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000191, 5'd0, 27'h000001a5, 5'd28, 27'h00000202, 32'h00000400,
  1'd1,  5'd17, 27'h000002c2, 5'd13, 27'h0000004a, 5'd4, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002fb, 5'd13, 27'h000001e6, 5'd10, 27'h0000034f, 32'h00000400,
  1'd1,  5'd17, 27'h000003b0, 5'd15, 27'h0000005a, 5'd22, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002c9, 5'd23, 27'h000001a0, 5'd4, 27'h00000083, 32'h00000400,
  1'd1,  5'd17, 27'h000003c9, 5'd25, 27'h0000018d, 5'd13, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000029f, 5'd24, 27'h00000162, 5'd24, 27'h000003d9, 32'h00000400,
  1'd1,  5'd30, 27'h0000027a, 5'd5, 27'h0000007b, 5'd2, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a8, 5'd0, 27'h00000149, 5'd10, 27'h000003d9, 32'h00000400,
  1'd1,  5'd27, 27'h0000018a, 5'd2, 27'h000003e8, 5'd21, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003a2, 5'd11, 27'h0000012b, 5'd3, 27'h00000236, 32'h00000400,
  1'd1,  5'd28, 27'h000001a8, 5'd11, 27'h00000081, 5'd13, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000312, 5'd12, 27'h000001d8, 5'd24, 27'h000002e4, 32'h00000400,
  1'd1,  5'd26, 27'h000003a4, 5'd22, 27'h00000025, 5'd1, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019e, 5'd23, 27'h00000297, 5'd14, 27'h0000025b, 32'h00000400,
  1'd1,  5'd25, 27'h00000394, 5'd25, 27'h00000292, 5'd22, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000031b, 5'd3, 27'h00000201, 5'd1, 27'h00000291, 32'h00000400,
  1'd1,  5'd9, 27'h0000036c, 5'd1, 27'h000001b7, 5'd10, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018f, 5'd2, 27'h000001a6, 5'd21, 27'h00000108, 32'h00000400,
  1'd1,  5'd9, 27'h00000101, 5'd11, 27'h000003a8, 5'd7, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000139, 5'd10, 27'h00000351, 5'd16, 27'h00000061, 32'h00000400,
  1'd1,  5'd5, 27'h00000100, 5'd14, 27'h000003e0, 5'd29, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023f, 5'd23, 27'h00000056, 5'd7, 27'h00000224, 32'h00000400,
  1'd1,  5'd6, 27'h000001b7, 5'd22, 27'h00000208, 5'd19, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ba, 5'd23, 27'h0000013b, 5'd29, 27'h000001a2, 32'h00000400,
  1'd1,  5'd16, 27'h00000284, 5'd4, 27'h000002a6, 5'd4, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000026f, 5'd2, 27'h00000051, 5'd13, 27'h0000030b, 32'h00000400,
  1'd1,  5'd20, 27'h000000bf, 5'd2, 27'h000002de, 5'd24, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b4, 5'd14, 27'h000001f9, 5'd9, 27'h00000235, 32'h00000400,
  1'd1,  5'd15, 27'h0000028f, 5'd10, 27'h000002bf, 5'd15, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000225, 5'd15, 27'h000000d9, 5'd29, 27'h0000038d, 32'h00000400,
  1'd1,  5'd17, 27'h000001a2, 5'd23, 27'h0000039e, 5'd7, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000028d, 5'd25, 27'h000002c4, 5'd16, 27'h00000248, 32'h00000400,
  1'd1,  5'd16, 27'h00000057, 5'd21, 27'h000003a4, 5'd30, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000011b, 5'd3, 27'h000002ee, 5'd6, 27'h00000082, 32'h00000400,
  1'd1,  5'd30, 27'h0000035d, 5'd5, 27'h00000031, 5'd18, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000fe, 5'd2, 27'h0000021d, 5'd27, 27'h00000007, 32'h00000400,
  1'd1,  5'd28, 27'h000000b3, 5'd11, 27'h0000031d, 5'd7, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b9, 5'd13, 27'h000003d8, 5'd17, 27'h0000022f, 32'h00000400,
  1'd1,  5'd29, 27'h000002fe, 5'd14, 27'h000001b2, 5'd26, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000d1, 5'd22, 27'h000001ba, 5'd7, 27'h00000399, 32'h00000400,
  1'd1,  5'd26, 27'h00000308, 5'd24, 27'h0000018f, 5'd18, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000266, 5'd25, 27'h00000018, 5'd28, 27'h000003f3, 32'h00000400,
  1'd1,  5'd9, 27'h000000b2, 5'd8, 27'h0000023a, 5'd3, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000018f, 5'd10, 27'h00000077, 5'd14, 27'h00000278, 32'h00000400,
  1'd1,  5'd8, 27'h00000013, 5'd6, 27'h000001c3, 5'd23, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000213, 5'd17, 27'h00000217, 5'd2, 27'h00000317, 32'h00000400,
  1'd1,  5'd7, 27'h0000007a, 5'd18, 27'h0000036c, 5'd12, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fc, 5'd17, 27'h000000b9, 5'd22, 27'h000001d7, 32'h00000400,
  1'd1,  5'd9, 27'h00000353, 5'd29, 27'h000001a3, 5'd0, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000075, 5'd30, 27'h0000003f, 5'd12, 27'h0000010d, 32'h00000400,
  1'd1,  5'd9, 27'h00000242, 5'd29, 27'h000001f4, 5'd21, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000034f, 5'd7, 27'h0000008e, 5'd1, 27'h000000c3, 32'h00000400,
  1'd1,  5'd17, 27'h0000017f, 5'd7, 27'h00000268, 5'd11, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000087, 5'd7, 27'h000003ca, 5'd24, 27'h000003fb, 32'h00000400,
  1'd1,  5'd20, 27'h00000045, 5'd17, 27'h00000340, 5'd2, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ff, 5'd15, 27'h00000256, 5'd13, 27'h000003d9, 32'h00000400,
  1'd1,  5'd16, 27'h0000038f, 5'd19, 27'h000003f7, 5'd21, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002aa, 5'd27, 27'h0000035c, 5'd0, 27'h0000004e, 32'h00000400,
  1'd1,  5'd17, 27'h00000129, 5'd29, 27'h00000084, 5'd11, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000e2, 5'd29, 27'h00000296, 5'd24, 27'h0000023f, 32'h00000400,
  1'd1,  5'd28, 27'h00000062, 5'd9, 27'h00000204, 5'd2, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000014, 5'd7, 27'h0000000b, 5'd13, 27'h0000037f, 32'h00000400,
  1'd1,  5'd27, 27'h0000002e, 5'd10, 27'h00000053, 5'd21, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e9, 5'd19, 27'h000002e7, 5'd0, 27'h00000126, 32'h00000400,
  1'd1,  5'd27, 27'h000003dc, 5'd18, 27'h00000222, 5'd15, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000055, 5'd19, 27'h0000008e, 5'd21, 27'h00000194, 32'h00000400,
  1'd1,  5'd29, 27'h000000ef, 5'd26, 27'h00000315, 5'd1, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000078, 5'd29, 27'h000002cb, 5'd14, 27'h000001c8, 32'h00000400,
  1'd1,  5'd30, 27'h00000032, 5'd29, 27'h00000248, 5'd23, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000145, 5'd7, 27'h0000021c, 5'd6, 27'h00000319, 32'h00000400,
  1'd1,  5'd10, 27'h000000a9, 5'd7, 27'h00000214, 5'd17, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000001c, 5'd7, 27'h000000ed, 5'd30, 27'h0000028a, 32'h00000400,
  1'd1,  5'd10, 27'h00000155, 5'd19, 27'h0000012e, 5'd6, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000162, 5'd17, 27'h00000181, 5'd16, 27'h00000126, 32'h00000400,
  1'd1,  5'd7, 27'h00000079, 5'd19, 27'h00000020, 5'd30, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000072, 5'd29, 27'h000002bf, 5'd5, 27'h00000257, 32'h00000400,
  1'd1,  5'd10, 27'h000000f7, 5'd26, 27'h00000125, 5'd20, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000008c, 5'd30, 27'h000000b2, 5'd27, 27'h0000031e, 32'h00000400,
  1'd1,  5'd19, 27'h000000af, 5'd6, 27'h00000300, 5'd6, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f1, 5'd5, 27'h000000e5, 5'd20, 27'h0000005e, 32'h00000400,
  1'd1,  5'd17, 27'h00000080, 5'd7, 27'h00000107, 5'd26, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ae, 5'd18, 27'h00000131, 5'd7, 27'h00000067, 32'h00000400,
  1'd1,  5'd17, 27'h00000339, 5'd16, 27'h0000039e, 5'd20, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000022b, 5'd19, 27'h000003fc, 5'd27, 27'h0000000d, 32'h00000400,
  1'd1,  5'd17, 27'h0000038e, 5'd28, 27'h000003b6, 5'd7, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001e9, 5'd30, 27'h00000112, 5'd18, 27'h000003e6, 32'h00000400,
  1'd1,  5'd18, 27'h00000080, 5'd26, 27'h00000090, 5'd30, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003cd, 5'd5, 27'h0000029a, 5'd8, 27'h0000019d, 32'h00000400,
  1'd1,  5'd30, 27'h000003fd, 5'd7, 27'h0000004a, 5'd20, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000013d, 5'd5, 27'h000000e7, 5'd30, 27'h000003e8, 32'h00000400,
  1'd1,  5'd29, 27'h0000023c, 5'd17, 27'h00000244, 5'd5, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b1, 5'd19, 27'h0000038c, 5'd19, 27'h000002c9, 32'h00000400,
  1'd1,  5'd30, 27'h000000f6, 5'd16, 27'h0000000e, 5'd26, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003db, 5'd26, 27'h000000ec, 5'd6, 27'h000001ec, 32'h00000400,
  1'd1,  5'd26, 27'h000002bd, 5'd30, 27'h0000023c, 5'd18, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000004a, 5'd27, 27'h00000383, 5'd28, 27'h000000f6, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000000b6, 5'd4, 27'h00000177, 5'd0, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d1, 5'd1, 27'h0000026a, 5'd12, 27'h000003ae, 32'h00000400,
  1'd1,  5'd0, 27'h0000026a, 5'd1, 27'h00000336, 5'd22, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000039f, 5'd14, 27'h00000147, 5'd0, 27'h0000027e, 32'h00000400,
  1'd1,  5'd4, 27'h0000006e, 5'd10, 27'h00000278, 5'd14, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000cf, 5'd12, 27'h0000037a, 5'd21, 27'h0000008b, 32'h00000400,
  1'd1,  5'd1, 27'h000000b0, 5'd24, 27'h0000027c, 5'd3, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ce, 5'd21, 27'h00000268, 5'd13, 27'h000003b3, 32'h00000400,
  1'd1,  5'd3, 27'h0000028c, 5'd24, 27'h00000163, 5'd23, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003ba, 5'd1, 27'h000003dd, 5'd4, 27'h0000032f, 32'h00000400,
  1'd1,  5'd15, 27'h0000013b, 5'd4, 27'h00000078, 5'd12, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000144, 5'd2, 27'h0000003b, 5'd25, 27'h0000027b, 32'h00000400,
  1'd1,  5'd13, 27'h0000037b, 5'd11, 27'h0000005e, 5'd0, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000289, 5'd10, 27'h0000018c, 5'd10, 27'h000003a1, 32'h00000400,
  1'd1,  5'd15, 27'h0000019a, 5'd10, 27'h00000279, 5'd24, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000033d, 5'd24, 27'h000002d6, 5'd1, 27'h000003cf, 32'h00000400,
  1'd1,  5'd11, 27'h00000294, 5'd22, 27'h00000313, 5'd14, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000003f, 5'd21, 27'h000000d1, 5'd24, 27'h0000005a, 32'h00000400,
  1'd1,  5'd24, 27'h00000095, 5'd4, 27'h000003a6, 5'd2, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d3, 5'd3, 27'h000002a8, 5'd11, 27'h0000018d, 32'h00000400,
  1'd1,  5'd25, 27'h00000098, 5'd0, 27'h0000025d, 5'd21, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d9, 5'd10, 27'h000003e0, 5'd3, 27'h00000114, 32'h00000400,
  1'd1,  5'd22, 27'h0000004b, 5'd12, 27'h00000063, 5'd13, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001bb, 5'd12, 27'h000000a8, 5'd24, 27'h00000193, 32'h00000400,
  1'd1,  5'd24, 27'h0000009a, 5'd21, 27'h00000113, 5'd2, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f9, 5'd24, 27'h00000078, 5'd15, 27'h000001f8, 32'h00000400,
  1'd1,  5'd22, 27'h000000eb, 5'd21, 27'h000001c3, 5'd23, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000070, 5'd3, 27'h000002ad, 5'd8, 27'h00000241, 32'h00000400,
  1'd1,  5'd3, 27'h00000158, 5'd1, 27'h000001ff, 5'd19, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000091, 5'd3, 27'h0000034b, 5'd27, 27'h00000175, 32'h00000400,
  1'd1,  5'd4, 27'h00000261, 5'd13, 27'h0000000d, 5'd9, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000229, 5'd15, 27'h000000d6, 5'd19, 27'h000003f4, 32'h00000400,
  1'd1,  5'd4, 27'h00000355, 5'd13, 27'h0000027a, 5'd30, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000007a, 5'd22, 27'h000002ad, 5'd5, 27'h00000115, 32'h00000400,
  1'd1,  5'd3, 27'h0000020b, 5'd21, 27'h0000034c, 5'd20, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000020b, 5'd23, 27'h0000004f, 5'd29, 27'h00000098, 32'h00000400,
  1'd1,  5'd14, 27'h000000b5, 5'd3, 27'h000002f5, 5'd6, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000038f, 5'd0, 27'h00000328, 5'd20, 27'h000000d2, 32'h00000400,
  1'd1,  5'd13, 27'h0000030e, 5'd4, 27'h0000031a, 5'd27, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000a2, 5'd13, 27'h00000229, 5'd5, 27'h00000323, 32'h00000400,
  1'd1,  5'd13, 27'h0000021d, 5'd11, 27'h0000000a, 5'd18, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f1, 5'd15, 27'h000001ce, 5'd27, 27'h0000039a, 32'h00000400,
  1'd1,  5'd14, 27'h00000051, 5'd24, 27'h0000016b, 5'd7, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000c6, 5'd23, 27'h00000113, 5'd18, 27'h000002dd, 32'h00000400,
  1'd1,  5'd10, 27'h0000032f, 5'd22, 27'h0000022d, 5'd26, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000296, 5'd4, 27'h000003fb, 5'd9, 27'h000000c2, 32'h00000400,
  1'd1,  5'd23, 27'h000003a7, 5'd0, 27'h0000006f, 5'd15, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001df, 5'd3, 27'h00000281, 5'd30, 27'h0000004a, 32'h00000400,
  1'd1,  5'd24, 27'h0000012f, 5'd12, 27'h000000dc, 5'd6, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000000c, 5'd11, 27'h000001c1, 5'd19, 27'h0000022a, 32'h00000400,
  1'd1,  5'd22, 27'h0000018c, 5'd14, 27'h00000117, 5'd28, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002de, 5'd21, 27'h00000143, 5'd10, 27'h00000069, 32'h00000400,
  1'd1,  5'd23, 27'h00000184, 5'd22, 27'h00000162, 5'd15, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002fe, 5'd22, 27'h0000019e, 5'd30, 27'h0000016b, 32'h00000400,
  1'd1,  5'd2, 27'h0000002b, 5'd9, 27'h000002fc, 5'd3, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000008a, 5'd9, 27'h00000209, 5'd11, 27'h00000318, 32'h00000400,
  1'd1,  5'd5, 27'h00000080, 5'd8, 27'h00000280, 5'd25, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000324, 5'd19, 27'h000003ae, 5'd3, 27'h0000038a, 32'h00000400,
  1'd1,  5'd3, 27'h00000107, 5'd17, 27'h0000021a, 5'd11, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000144, 5'd16, 27'h000001cd, 5'd24, 27'h00000180, 32'h00000400,
  1'd1,  5'd0, 27'h000003e2, 5'd28, 27'h00000240, 5'd3, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000024e, 5'd30, 27'h00000185, 5'd10, 27'h000002e3, 32'h00000400,
  1'd1,  5'd4, 27'h00000224, 5'd30, 27'h000003b3, 5'd23, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000082, 5'd6, 27'h00000010, 5'd3, 27'h0000000b, 32'h00000400,
  1'd1,  5'd11, 27'h0000005e, 5'd5, 27'h000002bd, 5'd13, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000228, 5'd9, 27'h0000001c, 5'd21, 27'h00000127, 32'h00000400,
  1'd1,  5'd11, 27'h0000021d, 5'd17, 27'h0000011d, 5'd4, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000024d, 5'd19, 27'h000001ac, 5'd14, 27'h00000354, 32'h00000400,
  1'd1,  5'd14, 27'h000001d0, 5'd17, 27'h00000084, 5'd22, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f8, 5'd29, 27'h000003ab, 5'd0, 27'h000002d1, 32'h00000400,
  1'd1,  5'd14, 27'h00000068, 5'd29, 27'h00000230, 5'd13, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029f, 5'd30, 27'h0000001d, 5'd21, 27'h00000187, 32'h00000400,
  1'd1,  5'd24, 27'h00000150, 5'd6, 27'h00000110, 5'd1, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000f2, 5'd6, 27'h000000cc, 5'd13, 27'h00000027, 32'h00000400,
  1'd1,  5'd24, 27'h000002f5, 5'd7, 27'h000002eb, 5'd23, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002fc, 5'd16, 27'h00000379, 5'd4, 27'h000002f0, 32'h00000400,
  1'd1,  5'd23, 27'h000001e6, 5'd16, 27'h000000b3, 5'd13, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000023, 5'd20, 27'h00000220, 5'd23, 27'h000001fd, 32'h00000400,
  1'd1,  5'd23, 27'h000001e3, 5'd28, 27'h0000028a, 5'd4, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000fb, 5'd28, 27'h000001f2, 5'd11, 27'h000003b4, 32'h00000400,
  1'd1,  5'd21, 27'h00000288, 5'd28, 27'h000001a5, 5'd22, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000345, 5'd8, 27'h000001e3, 5'd5, 27'h0000013a, 32'h00000400,
  1'd1,  5'd4, 27'h000001b3, 5'd8, 27'h00000034, 5'd17, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000311, 5'd8, 27'h00000166, 5'd29, 27'h0000007d, 32'h00000400,
  1'd1,  5'd0, 27'h0000007d, 5'd20, 27'h000001de, 5'd8, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000004a, 5'd20, 27'h00000178, 5'd18, 27'h000002d7, 32'h00000400,
  1'd1,  5'd1, 27'h000001db, 5'd16, 27'h00000276, 5'd26, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a9, 5'd28, 27'h000001e6, 5'd9, 27'h0000001f, 32'h00000400,
  1'd1,  5'd4, 27'h0000035b, 5'd27, 27'h00000181, 5'd17, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000156, 5'd30, 27'h000002e6, 5'd27, 27'h0000029e, 32'h00000400,
  1'd1,  5'd12, 27'h000002fc, 5'd10, 27'h000000e9, 5'd9, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003ea, 5'd10, 27'h0000002c, 5'd17, 27'h000002ef, 32'h00000400,
  1'd1,  5'd10, 27'h000002dd, 5'd7, 27'h0000014e, 5'd30, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000a3, 5'd16, 27'h0000022c, 5'd6, 27'h00000207, 32'h00000400,
  1'd1,  5'd13, 27'h0000024c, 5'd18, 27'h00000396, 5'd16, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ee, 5'd18, 27'h000001e8, 5'd30, 27'h000003cb, 32'h00000400,
  1'd1,  5'd11, 27'h000001fc, 5'd28, 27'h00000237, 5'd5, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000002e, 5'd26, 27'h0000037a, 5'd16, 27'h00000368, 32'h00000400,
  1'd1,  5'd13, 27'h000002b5, 5'd29, 27'h0000020d, 5'd30, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000143, 5'd7, 27'h0000035f, 5'd7, 27'h00000382, 32'h00000400,
  1'd1,  5'd24, 27'h00000214, 5'd8, 27'h000003e5, 5'd18, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000029e, 5'd7, 27'h00000193, 5'd29, 27'h0000016e, 32'h00000400,
  1'd1,  5'd22, 27'h0000037d, 5'd20, 27'h000001d9, 5'd5, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000033d, 5'd17, 27'h00000328, 5'd16, 27'h00000061, 32'h00000400,
  1'd1,  5'd23, 27'h000002f4, 5'd16, 27'h0000007b, 5'd29, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000242, 5'd29, 27'h000000d0, 5'd8, 27'h000003f2, 32'h00000400,
  1'd1,  5'd24, 27'h000002a4, 5'd30, 27'h000002ae, 5'd20, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ae, 5'd29, 27'h000001f8, 5'd29, 27'h00000154, 32'h00000400,
  1'd1,  5'd6, 27'h0000026b, 5'd0, 27'h000002ee, 5'd10, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001bd, 5'd4, 27'h000003fa, 5'd15, 27'h00000321, 32'h00000400,
  1'd1,  5'd5, 27'h00000166, 5'd3, 27'h00000036, 5'd30, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000032f, 5'd13, 27'h000000cd, 5'd3, 27'h00000169, 32'h00000400,
  1'd1,  5'd6, 27'h0000017a, 5'd13, 27'h00000006, 5'd14, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000126, 5'd14, 27'h0000003e, 5'd25, 27'h0000019a, 32'h00000400,
  1'd1,  5'd7, 27'h00000026, 5'd22, 27'h000000db, 5'd2, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003a, 5'd21, 27'h0000019d, 5'd14, 27'h000002ca, 32'h00000400,
  1'd1,  5'd8, 27'h0000027d, 5'd24, 27'h000002f6, 5'd24, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000016e, 5'd5, 27'h00000091, 5'd8, 27'h000003bd, 32'h00000400,
  1'd1,  5'd18, 27'h00000273, 5'd2, 27'h00000033, 5'd15, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000036f, 5'd3, 27'h000001e1, 5'd30, 27'h00000181, 32'h00000400,
  1'd1,  5'd15, 27'h00000385, 5'd12, 27'h000001d7, 5'd0, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c7, 5'd11, 27'h00000053, 5'd12, 27'h0000039f, 32'h00000400,
  1'd1,  5'd20, 27'h000000fe, 5'd14, 27'h0000027f, 5'd22, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029d, 5'd24, 27'h000001f6, 5'd4, 27'h0000011b, 32'h00000400,
  1'd1,  5'd20, 27'h00000075, 5'd23, 27'h0000009c, 5'd10, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000009b, 5'd24, 27'h0000021b, 5'd23, 27'h00000356, 32'h00000400,
  1'd1,  5'd29, 27'h000002f1, 5'd1, 27'h0000011c, 5'd1, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e5, 5'd0, 27'h00000073, 5'd11, 27'h0000002e, 32'h00000400,
  1'd1,  5'd29, 27'h000001e1, 5'd0, 27'h0000014c, 5'd21, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000050, 5'd13, 27'h0000020f, 5'd2, 27'h00000394, 32'h00000400,
  1'd1,  5'd29, 27'h00000067, 5'd11, 27'h0000006b, 5'd14, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000bf, 5'd14, 27'h00000302, 5'd25, 27'h00000114, 32'h00000400,
  1'd1,  5'd29, 27'h000002fe, 5'd21, 27'h0000028d, 5'd3, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000032, 5'd22, 27'h00000034, 5'd11, 27'h000003c7, 32'h00000400,
  1'd1,  5'd29, 27'h00000102, 5'd23, 27'h000000d9, 5'd25, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001c0, 5'd2, 27'h000002da, 5'd2, 27'h00000305, 32'h00000400,
  1'd1,  5'd7, 27'h0000036a, 5'd4, 27'h0000025c, 5'd10, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000012, 5'd2, 27'h000002db, 5'd25, 27'h00000242, 32'h00000400,
  1'd1,  5'd5, 27'h00000254, 5'd10, 27'h0000039f, 5'd7, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000348, 5'd12, 27'h00000396, 5'd19, 27'h00000315, 32'h00000400,
  1'd1,  5'd8, 27'h00000094, 5'd11, 27'h0000025a, 5'd26, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c8, 5'd25, 27'h0000026c, 5'd5, 27'h0000031a, 32'h00000400,
  1'd1,  5'd7, 27'h000002b9, 5'd21, 27'h0000014d, 5'd18, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000195, 5'd23, 27'h00000212, 5'd28, 27'h000001e1, 32'h00000400,
  1'd1,  5'd18, 27'h00000256, 5'd3, 27'h0000017b, 5'd4, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000076, 5'd1, 27'h000000b8, 5'd11, 27'h00000190, 32'h00000400,
  1'd1,  5'd15, 27'h00000385, 5'd0, 27'h000001f3, 5'd25, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002f2, 5'd11, 27'h00000338, 5'd5, 27'h00000378, 32'h00000400,
  1'd1,  5'd18, 27'h00000054, 5'd10, 27'h00000315, 5'd19, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002cd, 5'd11, 27'h0000024b, 5'd29, 27'h000001e1, 32'h00000400,
  1'd1,  5'd18, 27'h000000f7, 5'd22, 27'h00000028, 5'd5, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000397, 5'd20, 27'h000002d6, 5'd17, 27'h000001c8, 32'h00000400,
  1'd1,  5'd20, 27'h000001f7, 5'd23, 27'h00000171, 5'd26, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f6, 5'd0, 27'h0000004f, 5'd6, 27'h000002f9, 32'h00000400,
  1'd1,  5'd26, 27'h0000019f, 5'd4, 27'h0000017e, 5'd20, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000329, 5'd1, 27'h00000090, 5'd27, 27'h000000d8, 32'h00000400,
  1'd1,  5'd27, 27'h00000237, 5'd12, 27'h0000038e, 5'd8, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d5, 5'd13, 27'h00000317, 5'd17, 27'h0000023e, 32'h00000400,
  1'd1,  5'd29, 27'h000001d6, 5'd14, 27'h00000291, 5'd26, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000019a, 5'd23, 27'h00000218, 5'd7, 27'h0000039e, 32'h00000400,
  1'd1,  5'd30, 27'h0000027d, 5'd21, 27'h000001a0, 5'd16, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000100, 5'd24, 27'h00000000, 5'd27, 27'h000000d0, 32'h00000400,
  1'd1,  5'd6, 27'h00000103, 5'd10, 27'h0000003a, 5'd4, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000e7, 5'd10, 27'h00000028, 5'd12, 27'h0000023d, 32'h00000400,
  1'd1,  5'd5, 27'h00000295, 5'd6, 27'h000000b2, 5'd21, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a3, 5'd19, 27'h00000141, 5'd0, 27'h00000115, 32'h00000400,
  1'd1,  5'd5, 27'h000003c6, 5'd17, 27'h00000130, 5'd10, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002b8, 5'd16, 27'h000003bf, 5'd22, 27'h00000062, 32'h00000400,
  1'd1,  5'd5, 27'h00000304, 5'd27, 27'h00000201, 5'd4, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000010d, 5'd30, 27'h00000214, 5'd12, 27'h000001bd, 32'h00000400,
  1'd1,  5'd9, 27'h0000002b, 5'd30, 27'h0000021e, 5'd21, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039b, 5'd6, 27'h00000145, 5'd0, 27'h0000015d, 32'h00000400,
  1'd1,  5'd18, 27'h000002e6, 5'd9, 27'h00000289, 5'd12, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000281, 5'd7, 27'h00000347, 5'd21, 27'h00000077, 32'h00000400,
  1'd1,  5'd18, 27'h00000169, 5'd17, 27'h00000316, 5'd2, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000081, 5'd17, 27'h000001ea, 5'd10, 27'h00000196, 32'h00000400,
  1'd1,  5'd17, 27'h00000346, 5'd15, 27'h000002da, 5'd22, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000018, 5'd29, 27'h0000028b, 5'd2, 27'h0000003d, 32'h00000400,
  1'd1,  5'd18, 27'h000001ed, 5'd29, 27'h000001cb, 5'd12, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000029c, 5'd29, 27'h000003ef, 5'd24, 27'h00000008, 32'h00000400,
  1'd1,  5'd26, 27'h00000017, 5'd5, 27'h0000029a, 5'd0, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000257, 5'd7, 27'h00000275, 5'd10, 27'h0000017c, 32'h00000400,
  1'd1,  5'd29, 27'h000002d3, 5'd8, 27'h0000016d, 5'd21, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000031, 5'd19, 27'h00000310, 5'd1, 27'h000003d8, 32'h00000400,
  1'd1,  5'd28, 27'h00000235, 5'd20, 27'h0000028b, 5'd13, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000087, 5'd19, 27'h00000222, 5'd21, 27'h0000004a, 32'h00000400,
  1'd1,  5'd29, 27'h00000246, 5'd27, 27'h0000001d, 5'd1, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000049, 5'd30, 27'h00000244, 5'd14, 27'h00000057, 32'h00000400,
  1'd1,  5'd27, 27'h0000004c, 5'd28, 27'h0000026c, 5'd22, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002b7, 5'd7, 27'h00000333, 5'd8, 27'h0000035b, 32'h00000400,
  1'd1,  5'd8, 27'h000002e6, 5'd7, 27'h000000f5, 5'd16, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000012a, 5'd5, 27'h000003f6, 5'd27, 27'h0000026e, 32'h00000400,
  1'd1,  5'd8, 27'h0000024c, 5'd20, 27'h00000172, 5'd6, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000112, 5'd20, 27'h000000b1, 5'd19, 27'h0000029e, 32'h00000400,
  1'd1,  5'd7, 27'h000002b6, 5'd16, 27'h00000091, 5'd28, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013d, 5'd30, 27'h0000011d, 5'd5, 27'h0000024f, 32'h00000400,
  1'd1,  5'd8, 27'h000001ff, 5'd30, 27'h00000215, 5'd17, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000084, 5'd27, 27'h00000282, 5'd27, 27'h00000321, 32'h00000400,
  1'd1,  5'd19, 27'h000000fc, 5'd7, 27'h00000227, 5'd7, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003e7, 5'd6, 27'h00000042, 5'd18, 27'h00000102, 32'h00000400,
  1'd1,  5'd18, 27'h000000e2, 5'd5, 27'h00000280, 5'd27, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000015e, 5'd18, 27'h000001fd, 5'd6, 27'h0000004a, 32'h00000400,
  1'd1,  5'd16, 27'h000003ea, 5'd18, 27'h00000086, 5'd18, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006d, 5'd19, 27'h000002a7, 5'd27, 27'h000002a4, 32'h00000400,
  1'd1,  5'd18, 27'h00000199, 5'd26, 27'h000000a7, 5'd9, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000325, 5'd28, 27'h00000131, 5'd15, 27'h00000341, 32'h00000400,
  1'd1,  5'd17, 27'h000003dc, 5'd26, 27'h0000025e, 5'd27, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000172, 5'd6, 27'h00000366, 5'd9, 27'h000000b2, 32'h00000400,
  1'd1,  5'd29, 27'h000001e1, 5'd8, 27'h000001da, 5'd16, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000029e, 5'd6, 27'h000003e7, 5'd27, 27'h0000013f, 32'h00000400,
  1'd1,  5'd30, 27'h00000078, 5'd16, 27'h000000aa, 5'd8, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000388, 5'd17, 27'h0000013e, 5'd19, 27'h0000037d, 32'h00000400,
  1'd1,  5'd27, 27'h0000015b, 5'd20, 27'h00000172, 5'd28, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b9, 5'd29, 27'h0000016d, 5'd6, 27'h000000e1, 32'h00000400,
  1'd1,  5'd30, 27'h00000219, 5'd29, 27'h00000247, 5'd18, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a7, 5'd28, 27'h000001b6, 5'd26, 27'h000001fc, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000117, 5'd2, 27'h000002f5, 5'd2, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000224, 5'd1, 27'h00000149, 5'd12, 27'h00000198, 32'h00000400,
  1'd1,  5'd4, 27'h0000012b, 5'd2, 27'h00000313, 5'd22, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002fc, 5'd14, 27'h00000385, 5'd1, 27'h00000057, 32'h00000400,
  1'd1,  5'd1, 27'h00000345, 5'd15, 27'h00000168, 5'd13, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000c9, 5'd11, 27'h00000323, 5'd25, 27'h00000115, 32'h00000400,
  1'd1,  5'd2, 27'h000000db, 5'd25, 27'h00000154, 5'd3, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000003f, 5'd21, 27'h00000136, 5'd10, 27'h000002bb, 32'h00000400,
  1'd1,  5'd4, 27'h00000296, 5'd22, 27'h0000014c, 5'd23, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000078, 5'd4, 27'h000002e6, 5'd1, 27'h00000202, 32'h00000400,
  1'd1,  5'd15, 27'h00000031, 5'd1, 27'h00000331, 5'd15, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000009d, 5'd1, 27'h00000071, 5'd23, 27'h000003ee, 32'h00000400,
  1'd1,  5'd13, 27'h000003ff, 5'd13, 27'h000003bf, 5'd1, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000169, 5'd12, 27'h0000004b, 5'd14, 27'h000001c8, 32'h00000400,
  1'd1,  5'd11, 27'h000002ec, 5'd12, 27'h00000195, 5'd22, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000365, 5'd21, 27'h000001c7, 5'd0, 27'h00000050, 32'h00000400,
  1'd1,  5'd11, 27'h000000a5, 5'd22, 27'h00000047, 5'd13, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000055, 5'd21, 27'h00000214, 5'd21, 27'h0000018a, 32'h00000400,
  1'd1,  5'd22, 27'h000003fb, 5'd0, 27'h000001b2, 5'd0, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000f3, 5'd4, 27'h0000004d, 5'd15, 27'h0000009b, 32'h00000400,
  1'd1,  5'd22, 27'h000003bc, 5'd0, 27'h00000241, 5'd20, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e1, 5'd11, 27'h000002d9, 5'd1, 27'h00000003, 32'h00000400,
  1'd1,  5'd22, 27'h00000213, 5'd13, 27'h00000387, 5'd13, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002c0, 5'd12, 27'h000000ad, 5'd25, 27'h00000113, 32'h00000400,
  1'd1,  5'd25, 27'h00000156, 5'd25, 27'h00000320, 5'd0, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000179, 5'd25, 27'h00000271, 5'd12, 27'h00000347, 32'h00000400,
  1'd1,  5'd25, 27'h00000177, 5'd23, 27'h00000048, 5'd21, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000f9, 5'd4, 27'h000003ef, 5'd7, 27'h0000011e, 32'h00000400,
  1'd1,  5'd0, 27'h0000020f, 5'd0, 27'h00000053, 5'd15, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a6, 5'd2, 27'h00000250, 5'd25, 27'h000003a1, 32'h00000400,
  1'd1,  5'd1, 27'h000002d6, 5'd14, 27'h000002c5, 5'd10, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000287, 5'd13, 27'h0000003c, 5'd20, 27'h000000c7, 32'h00000400,
  1'd1,  5'd4, 27'h00000335, 5'd14, 27'h00000127, 5'd25, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000043, 5'd24, 27'h00000182, 5'd9, 27'h0000035b, 32'h00000400,
  1'd1,  5'd2, 27'h00000135, 5'd20, 27'h000002f1, 5'd18, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000349, 5'd24, 27'h000002fd, 5'd27, 27'h000003fa, 32'h00000400,
  1'd1,  5'd13, 27'h0000024e, 5'd0, 27'h000001a0, 5'd7, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003b, 5'd3, 27'h000002d5, 5'd18, 27'h0000006b, 32'h00000400,
  1'd1,  5'd12, 27'h000003a4, 5'd3, 27'h000000c6, 5'd26, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000d7, 5'd13, 27'h0000021f, 5'd6, 27'h00000073, 32'h00000400,
  1'd1,  5'd13, 27'h0000028c, 5'd14, 27'h00000329, 5'd16, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000011f, 5'd12, 27'h000001d9, 5'd30, 27'h00000395, 32'h00000400,
  1'd1,  5'd10, 27'h0000019b, 5'd23, 27'h0000039e, 5'd6, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c5, 5'd21, 27'h0000001f, 5'd19, 27'h000000f9, 32'h00000400,
  1'd1,  5'd13, 27'h000001c7, 5'd22, 27'h000002c1, 5'd27, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000039b, 5'd4, 27'h00000211, 5'd6, 27'h000001b3, 32'h00000400,
  1'd1,  5'd20, 27'h000003d4, 5'd2, 27'h0000004f, 5'd17, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000380, 5'd3, 27'h0000002f, 5'd30, 27'h00000242, 32'h00000400,
  1'd1,  5'd24, 27'h000000ff, 5'd13, 27'h00000058, 5'd5, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e9, 5'd15, 27'h00000098, 5'd17, 27'h0000001c, 32'h00000400,
  1'd1,  5'd24, 27'h0000002f, 5'd14, 27'h00000241, 5'd28, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001bd, 5'd24, 27'h00000070, 5'd6, 27'h00000222, 32'h00000400,
  1'd1,  5'd25, 27'h0000033b, 5'd24, 27'h0000038e, 5'd18, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c9, 5'd22, 27'h000002ed, 5'd30, 27'h00000249, 32'h00000400,
  1'd1,  5'd0, 27'h00000262, 5'd6, 27'h00000327, 5'd5, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b8, 5'd9, 27'h0000012d, 5'd12, 27'h00000283, 32'h00000400,
  1'd1,  5'd2, 27'h0000032f, 5'd9, 27'h0000014f, 5'd23, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000205, 5'd15, 27'h0000027e, 5'd5, 27'h00000047, 32'h00000400,
  1'd1,  5'd1, 27'h000002b4, 5'd16, 27'h00000181, 5'd14, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000279, 5'd18, 27'h00000276, 5'd24, 27'h0000035f, 32'h00000400,
  1'd1,  5'd0, 27'h000003ed, 5'd30, 27'h00000225, 5'd2, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001df, 5'd27, 27'h00000028, 5'd12, 27'h000003e7, 32'h00000400,
  1'd1,  5'd3, 27'h00000032, 5'd27, 27'h00000077, 5'd23, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000198, 5'd7, 27'h0000006b, 5'd4, 27'h00000189, 32'h00000400,
  1'd1,  5'd14, 27'h00000335, 5'd8, 27'h0000038e, 5'd15, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f2, 5'd5, 27'h000002ae, 5'd21, 27'h00000223, 32'h00000400,
  1'd1,  5'd14, 27'h000001d3, 5'd20, 27'h00000056, 5'd4, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000039c, 5'd15, 27'h000002b9, 5'd13, 27'h00000077, 32'h00000400,
  1'd1,  5'd12, 27'h00000308, 5'd16, 27'h00000386, 5'd25, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000eb, 5'd27, 27'h000000ec, 5'd4, 27'h00000314, 32'h00000400,
  1'd1,  5'd14, 27'h0000000d, 5'd26, 27'h0000010d, 5'd11, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002a8, 5'd29, 27'h00000400, 5'd25, 27'h00000042, 32'h00000400,
  1'd1,  5'd23, 27'h00000201, 5'd9, 27'h00000392, 5'd3, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001e2, 5'd6, 27'h000003a9, 5'd12, 27'h000002f8, 32'h00000400,
  1'd1,  5'd21, 27'h0000017c, 5'd8, 27'h0000025b, 5'd22, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000008b, 5'd20, 27'h00000242, 5'd3, 27'h000002e7, 32'h00000400,
  1'd1,  5'd25, 27'h00000058, 5'd20, 27'h00000264, 5'd13, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000367, 5'd16, 27'h0000025d, 5'd21, 27'h000003f2, 32'h00000400,
  1'd1,  5'd22, 27'h000002c3, 5'd29, 27'h00000238, 5'd1, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ce, 5'd25, 27'h000003a7, 5'd12, 27'h00000054, 32'h00000400,
  1'd1,  5'd21, 27'h00000000, 5'd28, 27'h0000017f, 5'd24, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000170, 5'd5, 27'h000002c6, 5'd10, 27'h00000044, 32'h00000400,
  1'd1,  5'd0, 27'h000000c3, 5'd8, 27'h000001dc, 5'd17, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f2, 5'd6, 27'h00000195, 5'd30, 27'h0000010e, 32'h00000400,
  1'd1,  5'd2, 27'h0000019a, 5'd17, 27'h0000016a, 5'd9, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000009b, 5'd16, 27'h000003fd, 5'd18, 27'h00000348, 32'h00000400,
  1'd1,  5'd2, 27'h00000012, 5'd19, 27'h00000289, 5'd27, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000034a, 5'd29, 27'h0000031e, 5'd5, 27'h00000370, 32'h00000400,
  1'd1,  5'd1, 27'h000000b6, 5'd28, 27'h00000204, 5'd16, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000d1, 5'd26, 27'h00000113, 5'd29, 27'h00000288, 32'h00000400,
  1'd1,  5'd15, 27'h00000015, 5'd6, 27'h00000104, 5'd8, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000032a, 5'd9, 27'h00000115, 5'd18, 27'h000002b4, 32'h00000400,
  1'd1,  5'd14, 27'h000001c0, 5'd6, 27'h000003a6, 5'd29, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000034b, 5'd15, 27'h000002b1, 5'd7, 27'h00000078, 32'h00000400,
  1'd1,  5'd10, 27'h00000392, 5'd20, 27'h0000000d, 5'd19, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000031e, 5'd19, 27'h0000018e, 5'd27, 27'h00000111, 32'h00000400,
  1'd1,  5'd11, 27'h00000195, 5'd29, 27'h00000254, 5'd8, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002fd, 5'd28, 27'h0000000d, 5'd15, 27'h000002fd, 32'h00000400,
  1'd1,  5'd13, 27'h00000200, 5'd28, 27'h000001a6, 5'd30, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000027a, 5'd5, 27'h00000238, 5'd7, 27'h00000270, 32'h00000400,
  1'd1,  5'd22, 27'h00000347, 5'd9, 27'h000000fd, 5'd17, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000016f, 5'd9, 27'h00000310, 5'd26, 27'h00000079, 32'h00000400,
  1'd1,  5'd24, 27'h000003f2, 5'd19, 27'h00000222, 5'd8, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fa, 5'd16, 27'h000002b8, 5'd15, 27'h000003a5, 32'h00000400,
  1'd1,  5'd24, 27'h0000018f, 5'd20, 27'h000000a6, 5'd29, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000fd, 5'd30, 27'h000000f7, 5'd8, 27'h000001b6, 32'h00000400,
  1'd1,  5'd24, 27'h000000cf, 5'd27, 27'h00000387, 5'd19, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000030, 5'd30, 27'h00000117, 5'd27, 27'h0000015a, 32'h00000400,
  1'd1,  5'd5, 27'h000003b8, 5'd2, 27'h000002fc, 5'd6, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000035e, 5'd0, 27'h00000021, 5'd16, 27'h0000019d, 32'h00000400,
  1'd1,  5'd6, 27'h00000344, 5'd4, 27'h00000168, 5'd29, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ad, 5'd15, 27'h0000002b, 5'd0, 27'h00000267, 32'h00000400,
  1'd1,  5'd5, 27'h000003cb, 5'd11, 27'h000003b2, 5'd11, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000331, 5'd11, 27'h000000c4, 5'd25, 27'h0000019b, 32'h00000400,
  1'd1,  5'd5, 27'h00000294, 5'd25, 27'h00000172, 5'd2, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000196, 5'd23, 27'h000000f0, 5'd13, 27'h00000338, 32'h00000400,
  1'd1,  5'd5, 27'h0000026c, 5'd22, 27'h0000019d, 5'd25, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000179, 5'd1, 27'h0000020d, 5'd5, 27'h000002cd, 32'h00000400,
  1'd1,  5'd15, 27'h000002af, 5'd2, 27'h00000094, 5'd19, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d6, 5'd4, 27'h0000012e, 5'd29, 27'h000001ee, 32'h00000400,
  1'd1,  5'd16, 27'h00000333, 5'd10, 27'h000002f0, 5'd2, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c0, 5'd12, 27'h000000e1, 5'd14, 27'h0000010a, 32'h00000400,
  1'd1,  5'd17, 27'h000000e4, 5'd11, 27'h00000020, 5'd21, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000236, 5'd21, 27'h000003c1, 5'd4, 27'h0000036b, 32'h00000400,
  1'd1,  5'd16, 27'h000003e9, 5'd21, 27'h000002cd, 5'd11, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e5, 5'd24, 27'h00000080, 5'd25, 27'h000000ff, 32'h00000400,
  1'd1,  5'd29, 27'h0000014e, 5'd2, 27'h000001c8, 5'd3, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000266, 5'd1, 27'h000002e7, 5'd12, 27'h000003dc, 32'h00000400,
  1'd1,  5'd28, 27'h0000009a, 5'd3, 27'h000002b2, 5'd23, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000011, 5'd12, 27'h00000139, 5'd4, 27'h00000124, 32'h00000400,
  1'd1,  5'd27, 27'h000000e7, 5'd11, 27'h00000075, 5'd12, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000010c, 5'd13, 27'h00000022, 5'd23, 27'h00000023, 32'h00000400,
  1'd1,  5'd26, 27'h00000363, 5'd23, 27'h000001ca, 5'd3, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000015a, 5'd23, 27'h00000090, 5'd12, 27'h000002b1, 32'h00000400,
  1'd1,  5'd29, 27'h0000031d, 5'd22, 27'h000003f2, 5'd21, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000036e, 5'd1, 27'h000003c0, 5'd0, 27'h00000334, 32'h00000400,
  1'd1,  5'd10, 27'h00000009, 5'd0, 27'h0000039e, 5'd13, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000005d, 5'd2, 27'h00000034, 5'd25, 27'h000000bf, 32'h00000400,
  1'd1,  5'd7, 27'h000003fb, 5'd10, 27'h0000024a, 5'd9, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d7, 5'd10, 27'h00000201, 5'd17, 27'h0000032b, 32'h00000400,
  1'd1,  5'd6, 27'h000002b7, 5'd12, 27'h00000118, 5'd26, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000178, 5'd22, 27'h000002d2, 5'd10, 27'h00000053, 32'h00000400,
  1'd1,  5'd7, 27'h00000246, 5'd23, 27'h000001f4, 5'd16, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000317, 5'd23, 27'h000000e4, 5'd27, 27'h0000011f, 32'h00000400,
  1'd1,  5'd16, 27'h0000018a, 5'd3, 27'h00000283, 5'd0, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000001a, 5'd0, 27'h00000043, 5'd14, 27'h00000027, 32'h00000400,
  1'd1,  5'd15, 27'h000002b1, 5'd3, 27'h00000310, 5'd21, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000237, 5'd12, 27'h000003c8, 5'd9, 27'h0000019f, 32'h00000400,
  1'd1,  5'd18, 27'h0000025a, 5'd13, 27'h0000030f, 5'd17, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002ed, 5'd11, 27'h0000028c, 5'd28, 27'h000002df, 32'h00000400,
  1'd1,  5'd17, 27'h000002ac, 5'd21, 27'h0000028e, 5'd8, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000054, 5'd23, 27'h000003d6, 5'd16, 27'h0000022f, 32'h00000400,
  1'd1,  5'd17, 27'h000001ec, 5'd22, 27'h00000169, 5'd29, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000035f, 5'd4, 27'h000003d8, 5'd5, 27'h000002d7, 32'h00000400,
  1'd1,  5'd26, 27'h00000080, 5'd1, 27'h0000025f, 5'd17, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000009a, 5'd1, 27'h00000306, 5'd30, 27'h000001bd, 32'h00000400,
  1'd1,  5'd26, 27'h00000269, 5'd14, 27'h000003ea, 5'd5, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b2, 5'd11, 27'h000002cb, 5'd18, 27'h00000217, 32'h00000400,
  1'd1,  5'd28, 27'h0000032b, 5'd14, 27'h000001b3, 5'd27, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000100, 5'd25, 27'h0000006f, 5'd8, 27'h0000022d, 32'h00000400,
  1'd1,  5'd29, 27'h00000008, 5'd22, 27'h000003ba, 5'd17, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000178, 5'd20, 27'h0000038f, 5'd30, 27'h000001a2, 32'h00000400,
  1'd1,  5'd7, 27'h000001dd, 5'd6, 27'h00000288, 5'd2, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000039e, 5'd8, 27'h0000033c, 5'd11, 27'h00000208, 32'h00000400,
  1'd1,  5'd8, 27'h00000271, 5'd5, 27'h00000155, 5'd21, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023b, 5'd17, 27'h00000343, 5'd2, 27'h00000306, 32'h00000400,
  1'd1,  5'd6, 27'h0000034d, 5'd17, 27'h0000036d, 5'd10, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002b3, 5'd16, 27'h00000055, 5'd24, 27'h0000038f, 32'h00000400,
  1'd1,  5'd7, 27'h000000d0, 5'd27, 27'h000001c0, 5'd1, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ee, 5'd28, 27'h0000010f, 5'd11, 27'h0000017b, 32'h00000400,
  1'd1,  5'd7, 27'h0000032e, 5'd27, 27'h00000249, 5'd23, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000227, 5'd9, 27'h0000012b, 5'd2, 27'h00000359, 32'h00000400,
  1'd1,  5'd20, 27'h00000250, 5'd7, 27'h0000001f, 5'd13, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000022f, 5'd6, 27'h000003b5, 5'd25, 27'h0000020e, 32'h00000400,
  1'd1,  5'd17, 27'h0000008e, 5'd16, 27'h00000288, 5'd4, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000213, 5'd17, 27'h0000034d, 5'd12, 27'h00000125, 32'h00000400,
  1'd1,  5'd20, 27'h00000290, 5'd16, 27'h00000191, 5'd24, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000db, 5'd27, 27'h00000372, 5'd1, 27'h0000030d, 32'h00000400,
  1'd1,  5'd15, 27'h00000205, 5'd30, 27'h00000035, 5'd13, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000019, 5'd29, 27'h0000033b, 5'd24, 27'h0000010e, 32'h00000400,
  1'd1,  5'd28, 27'h00000324, 5'd6, 27'h000000b0, 5'd1, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000010c, 5'd10, 27'h0000003a, 5'd12, 27'h000002df, 32'h00000400,
  1'd1,  5'd29, 27'h000003f0, 5'd10, 27'h00000005, 5'd24, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003af, 5'd18, 27'h000002e8, 5'd3, 27'h000003d4, 32'h00000400,
  1'd1,  5'd28, 27'h0000001c, 5'd15, 27'h00000210, 5'd11, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002fa, 5'd20, 27'h0000004d, 5'd23, 27'h00000322, 32'h00000400,
  1'd1,  5'd29, 27'h00000089, 5'd28, 27'h0000038c, 5'd4, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000010b, 5'd28, 27'h000002dd, 5'd13, 27'h000001b4, 32'h00000400,
  1'd1,  5'd30, 27'h00000316, 5'd29, 27'h0000022a, 5'd21, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000029a, 5'd10, 27'h000000f5, 5'd5, 27'h00000206, 32'h00000400,
  1'd1,  5'd5, 27'h00000169, 5'd9, 27'h000000c7, 5'd19, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000141, 5'd6, 27'h00000347, 5'd28, 27'h00000050, 32'h00000400,
  1'd1,  5'd8, 27'h000000d4, 5'd17, 27'h000002e3, 5'd5, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000133, 5'd17, 27'h000003d7, 5'd18, 27'h0000005a, 32'h00000400,
  1'd1,  5'd9, 27'h000002f5, 5'd17, 27'h0000030a, 5'd30, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002f0, 5'd29, 27'h00000333, 5'd9, 27'h00000050, 32'h00000400,
  1'd1,  5'd8, 27'h00000350, 5'd28, 27'h00000190, 5'd16, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000027, 5'd26, 27'h0000022b, 5'd25, 27'h00000397, 32'h00000400,
  1'd1,  5'd15, 27'h000003da, 5'd5, 27'h000003a9, 5'd8, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a5, 5'd6, 27'h00000174, 5'd16, 27'h000003da, 32'h00000400,
  1'd1,  5'd20, 27'h0000016c, 5'd10, 27'h000000c6, 5'd27, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002da, 5'd16, 27'h000003de, 5'd5, 27'h000003b7, 32'h00000400,
  1'd1,  5'd19, 27'h000000f8, 5'd15, 27'h000003c3, 5'd17, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000269, 5'd16, 27'h0000038d, 5'd30, 27'h000003e4, 32'h00000400,
  1'd1,  5'd19, 27'h0000038f, 5'd29, 27'h0000001c, 5'd9, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000174, 5'd29, 27'h00000271, 5'd17, 27'h0000029b, 32'h00000400,
  1'd1,  5'd20, 27'h0000008c, 5'd26, 27'h00000150, 5'd27, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000035a, 5'd9, 27'h000000ff, 5'd6, 27'h000003f7, 32'h00000400,
  1'd1,  5'd27, 27'h000000de, 5'd6, 27'h0000011a, 5'd20, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000229, 5'd5, 27'h000000ff, 5'd28, 27'h0000004e, 32'h00000400,
  1'd1,  5'd27, 27'h000000c1, 5'd16, 27'h00000380, 5'd7, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f2, 5'd17, 27'h00000116, 5'd16, 27'h000000f9, 32'h00000400,
  1'd1,  5'd27, 27'h000000e9, 5'd16, 27'h00000052, 5'd29, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000026d, 5'd27, 27'h00000075, 5'd8, 27'h000001f9, 32'h00000400,
  1'd1,  5'd27, 27'h0000026d, 5'd28, 27'h000003f8, 5'd16, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019f, 5'd26, 27'h00000342, 5'd25, 27'h0000037c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000265, 5'd3, 27'h000001a0, 5'd4, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a6, 5'd4, 27'h0000024f, 5'd11, 27'h000003da, 32'h00000400,
  1'd1,  5'd4, 27'h00000217, 5'd4, 27'h000001e4, 5'd23, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003cf, 5'd10, 27'h0000030d, 5'd5, 27'h00000023, 32'h00000400,
  1'd1,  5'd0, 27'h0000016b, 5'd11, 27'h000002f4, 5'd15, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000106, 5'd12, 27'h00000170, 5'd22, 27'h00000142, 32'h00000400,
  1'd1,  5'd0, 27'h0000019d, 5'd21, 27'h000002df, 5'd4, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002f9, 5'd21, 27'h000002f0, 5'd13, 27'h00000271, 32'h00000400,
  1'd1,  5'd2, 27'h00000334, 5'd21, 27'h00000245, 5'd21, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001ec, 5'd2, 27'h00000217, 5'd4, 27'h000000a8, 32'h00000400,
  1'd1,  5'd11, 27'h00000053, 5'd1, 27'h000002ab, 5'd15, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000247, 5'd4, 27'h000002c7, 5'd24, 27'h00000128, 32'h00000400,
  1'd1,  5'd13, 27'h00000141, 5'd12, 27'h0000005c, 5'd3, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e6, 5'd11, 27'h00000060, 5'd11, 27'h00000160, 32'h00000400,
  1'd1,  5'd11, 27'h000003cf, 5'd11, 27'h000000d5, 5'd22, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000145, 5'd25, 27'h000001d4, 5'd2, 27'h000002a6, 32'h00000400,
  1'd1,  5'd12, 27'h00000353, 5'd24, 27'h00000125, 5'd10, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000286, 5'd21, 27'h00000024, 5'd25, 27'h00000010, 32'h00000400,
  1'd1,  5'd21, 27'h00000300, 5'd4, 27'h000003fd, 5'd4, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002cc, 5'd3, 27'h000002aa, 5'd14, 27'h00000178, 32'h00000400,
  1'd1,  5'd22, 27'h00000374, 5'd1, 27'h000002d8, 5'd22, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f8, 5'd12, 27'h000002f7, 5'd5, 27'h00000006, 32'h00000400,
  1'd1,  5'd25, 27'h000002bb, 5'd14, 27'h00000308, 5'd14, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000223, 5'd13, 27'h000002a7, 5'd21, 27'h000002b3, 32'h00000400,
  1'd1,  5'd22, 27'h000000d2, 5'd24, 27'h00000027, 5'd1, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000023a, 5'd21, 27'h000002cf, 5'd12, 27'h000000fb, 32'h00000400,
  1'd1,  5'd24, 27'h000000cc, 5'd25, 27'h000000c3, 5'd21, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ad, 5'd2, 27'h0000005e, 5'd5, 27'h00000252, 32'h00000400,
  1'd1,  5'd4, 27'h0000016d, 5'd5, 27'h00000031, 5'd19, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000007, 5'd4, 27'h0000038c, 5'd30, 27'h00000239, 32'h00000400,
  1'd1,  5'd0, 27'h000003fc, 5'd13, 27'h000002ce, 5'd7, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d0, 5'd14, 27'h00000385, 5'd17, 27'h000003a1, 32'h00000400,
  1'd1,  5'd0, 27'h000003ab, 5'd15, 27'h000001b5, 5'd30, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000062, 5'd24, 27'h0000003e, 5'd7, 27'h00000193, 32'h00000400,
  1'd1,  5'd1, 27'h000002b1, 5'd23, 27'h0000020d, 5'd15, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017e, 5'd22, 27'h0000037d, 5'd27, 27'h00000069, 32'h00000400,
  1'd1,  5'd11, 27'h00000086, 5'd4, 27'h00000392, 5'd9, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001fd, 5'd1, 27'h00000286, 5'd20, 27'h000001ba, 32'h00000400,
  1'd1,  5'd12, 27'h000002e0, 5'd2, 27'h0000021a, 5'd30, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001ed, 5'd14, 27'h000001ec, 5'd7, 27'h000001a6, 32'h00000400,
  1'd1,  5'd12, 27'h00000300, 5'd15, 27'h000001a1, 5'd18, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000232, 5'd14, 27'h00000080, 5'd28, 27'h0000020e, 32'h00000400,
  1'd1,  5'd14, 27'h0000013e, 5'd21, 27'h000003a0, 5'd8, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000056, 5'd24, 27'h00000081, 5'd19, 27'h00000065, 32'h00000400,
  1'd1,  5'd12, 27'h00000217, 5'd21, 27'h00000058, 5'd29, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000232, 5'd4, 27'h000003fb, 5'd6, 27'h0000020c, 32'h00000400,
  1'd1,  5'd22, 27'h00000212, 5'd1, 27'h000003bd, 5'd18, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000030d, 5'd1, 27'h000003ab, 5'd29, 27'h0000036c, 32'h00000400,
  1'd1,  5'd21, 27'h000001eb, 5'd13, 27'h0000036d, 5'd8, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000145, 5'd11, 27'h000000f0, 5'd20, 27'h0000001b, 32'h00000400,
  1'd1,  5'd21, 27'h000001f7, 5'd14, 27'h0000036c, 5'd26, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001a1, 5'd25, 27'h00000055, 5'd6, 27'h0000025a, 32'h00000400,
  1'd1,  5'd24, 27'h000001b6, 5'd21, 27'h000002b8, 5'd15, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001bf, 5'd23, 27'h00000279, 5'd28, 27'h00000312, 32'h00000400,
  1'd1,  5'd0, 27'h00000060, 5'd5, 27'h0000024a, 5'd4, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000309, 5'd10, 27'h0000002c, 5'd12, 27'h00000044, 32'h00000400,
  1'd1,  5'd3, 27'h000003a8, 5'd6, 27'h00000095, 5'd22, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000de, 5'd19, 27'h00000260, 5'd2, 27'h0000009d, 32'h00000400,
  1'd1,  5'd4, 27'h000002e1, 5'd17, 27'h00000341, 5'd12, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000007a, 5'd20, 27'h00000212, 5'd21, 27'h00000012, 32'h00000400,
  1'd1,  5'd2, 27'h000001b2, 5'd30, 27'h000002a4, 5'd2, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000018b, 5'd27, 27'h00000050, 5'd10, 27'h0000020c, 32'h00000400,
  1'd1,  5'd4, 27'h0000006b, 5'd27, 27'h000001df, 5'd23, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000116, 5'd9, 27'h00000058, 5'd1, 27'h0000026f, 32'h00000400,
  1'd1,  5'd15, 27'h000001b7, 5'd9, 27'h000002c8, 5'd14, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ed, 5'd9, 27'h000002ca, 5'd21, 27'h0000023f, 32'h00000400,
  1'd1,  5'd11, 27'h0000032b, 5'd17, 27'h000002e4, 5'd2, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000e8, 5'd19, 27'h00000396, 5'd13, 27'h00000213, 32'h00000400,
  1'd1,  5'd11, 27'h000003e6, 5'd17, 27'h000000eb, 5'd23, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f8, 5'd27, 27'h000002e9, 5'd1, 27'h0000037a, 32'h00000400,
  1'd1,  5'd15, 27'h00000004, 5'd26, 27'h0000026d, 5'd12, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e9, 5'd30, 27'h00000068, 5'd23, 27'h0000003b, 32'h00000400,
  1'd1,  5'd23, 27'h000000fc, 5'd6, 27'h000000ba, 5'd2, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001b0, 5'd7, 27'h00000147, 5'd13, 27'h00000349, 32'h00000400,
  1'd1,  5'd23, 27'h00000213, 5'd8, 27'h000001da, 5'd21, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ed, 5'd19, 27'h00000334, 5'd1, 27'h00000265, 32'h00000400,
  1'd1,  5'd22, 27'h0000009d, 5'd19, 27'h000003c3, 5'd11, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000015, 5'd16, 27'h00000116, 5'd23, 27'h000002e9, 32'h00000400,
  1'd1,  5'd25, 27'h0000023d, 5'd29, 27'h00000355, 5'd4, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b5, 5'd28, 27'h0000012c, 5'd12, 27'h00000264, 32'h00000400,
  1'd1,  5'd25, 27'h0000002c, 5'd26, 27'h00000376, 5'd24, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000009b, 5'd7, 27'h00000215, 5'd5, 27'h00000314, 32'h00000400,
  1'd1,  5'd2, 27'h00000345, 5'd8, 27'h000000c8, 5'd18, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002b0, 5'd6, 27'h00000145, 5'd27, 27'h000000bd, 32'h00000400,
  1'd1,  5'd0, 27'h000003c4, 5'd17, 27'h000002c3, 5'd6, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e4, 5'd18, 27'h000002d1, 5'd16, 27'h000001a1, 32'h00000400,
  1'd1,  5'd0, 27'h00000286, 5'd20, 27'h00000254, 5'd27, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fb, 5'd28, 27'h00000371, 5'd6, 27'h00000110, 32'h00000400,
  1'd1,  5'd3, 27'h00000114, 5'd27, 27'h00000160, 5'd16, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b0, 5'd27, 27'h0000019a, 5'd26, 27'h00000183, 32'h00000400,
  1'd1,  5'd15, 27'h00000167, 5'd5, 27'h000003ff, 5'd5, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002a8, 5'd6, 27'h000001ed, 5'd19, 27'h00000139, 32'h00000400,
  1'd1,  5'd13, 27'h00000280, 5'd6, 27'h0000029e, 5'd30, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000fb, 5'd19, 27'h00000158, 5'd8, 27'h0000024d, 32'h00000400,
  1'd1,  5'd14, 27'h0000002d, 5'd16, 27'h0000002c, 5'd20, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d2, 5'd18, 27'h000000db, 5'd30, 27'h0000030c, 32'h00000400,
  1'd1,  5'd13, 27'h00000138, 5'd29, 27'h00000304, 5'd5, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a1, 5'd27, 27'h000001c7, 5'd16, 27'h000000f8, 32'h00000400,
  1'd1,  5'd11, 27'h000001ed, 5'd30, 27'h00000227, 5'd29, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d6, 5'd8, 27'h0000020f, 5'd10, 27'h000000d2, 32'h00000400,
  1'd1,  5'd23, 27'h00000155, 5'd10, 27'h000000eb, 5'd18, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000015f, 5'd9, 27'h000002e2, 5'd27, 27'h00000349, 32'h00000400,
  1'd1,  5'd24, 27'h00000205, 5'd17, 27'h000000df, 5'd6, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000328, 5'd20, 27'h0000029a, 5'd18, 27'h00000268, 32'h00000400,
  1'd1,  5'd21, 27'h0000033f, 5'd18, 27'h00000019, 5'd29, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000036f, 5'd30, 27'h0000012f, 5'd7, 27'h00000314, 32'h00000400,
  1'd1,  5'd24, 27'h00000202, 5'd27, 27'h000002e1, 5'd20, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000351, 5'd30, 27'h00000135, 5'd27, 27'h00000355, 32'h00000400,
  1'd1,  5'd6, 27'h000002b6, 5'd3, 27'h000000a5, 5'd9, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001b9, 5'd0, 27'h000002b5, 5'd20, 27'h00000270, 32'h00000400,
  1'd1,  5'd5, 27'h000002c4, 5'd3, 27'h000000c6, 5'd28, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ed, 5'd10, 27'h0000026f, 5'd4, 27'h00000081, 32'h00000400,
  1'd1,  5'd7, 27'h000002a0, 5'd10, 27'h00000272, 5'd11, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000077, 5'd11, 27'h000002bb, 5'd20, 27'h000003c3, 32'h00000400,
  1'd1,  5'd5, 27'h00000265, 5'd20, 27'h00000365, 5'd4, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000c2, 5'd24, 27'h000001e6, 5'd10, 27'h000002f8, 32'h00000400,
  1'd1,  5'd7, 27'h0000038c, 5'd24, 27'h00000077, 5'd21, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000103, 5'd2, 27'h0000033b, 5'd9, 27'h00000007, 32'h00000400,
  1'd1,  5'd19, 27'h0000021b, 5'd3, 27'h000000e2, 5'd20, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000330, 5'd0, 27'h000003e4, 5'd28, 27'h000003ad, 32'h00000400,
  1'd1,  5'd18, 27'h00000098, 5'd15, 27'h000001c4, 5'd3, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001cf, 5'd12, 27'h000000cc, 5'd10, 27'h000001b5, 32'h00000400,
  1'd1,  5'd19, 27'h0000007e, 5'd14, 27'h00000153, 5'd23, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002a2, 5'd24, 27'h0000000b, 5'd3, 27'h000003a8, 32'h00000400,
  1'd1,  5'd16, 27'h00000272, 5'd24, 27'h000001cf, 5'd12, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000031b, 5'd25, 27'h00000261, 5'd25, 27'h000002bf, 32'h00000400,
  1'd1,  5'd28, 27'h000003dc, 5'd0, 27'h0000008c, 5'd2, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000394, 5'd0, 27'h00000046, 5'd12, 27'h000001da, 32'h00000400,
  1'd1,  5'd29, 27'h0000000b, 5'd3, 27'h00000265, 5'd22, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b3, 5'd10, 27'h00000263, 5'd4, 27'h00000298, 32'h00000400,
  1'd1,  5'd29, 27'h00000240, 5'd14, 27'h00000285, 5'd15, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000027a, 5'd13, 27'h0000009d, 5'd23, 27'h000001e4, 32'h00000400,
  1'd1,  5'd27, 27'h0000017d, 5'd21, 27'h000000a3, 5'd3, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000021b, 5'd22, 27'h00000052, 5'd15, 27'h000000d6, 32'h00000400,
  1'd1,  5'd28, 27'h00000388, 5'd21, 27'h000000c7, 5'd21, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000127, 5'd3, 27'h00000313, 5'd0, 27'h00000287, 32'h00000400,
  1'd1,  5'd6, 27'h000002ef, 5'd4, 27'h0000021e, 5'd14, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000171, 5'd0, 27'h000003d8, 5'd25, 27'h00000122, 32'h00000400,
  1'd1,  5'd5, 27'h000003cc, 5'd11, 27'h000001e3, 5'd6, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000087, 5'd10, 27'h000001aa, 5'd16, 27'h000003b1, 32'h00000400,
  1'd1,  5'd6, 27'h000001ea, 5'd14, 27'h000003b6, 5'd28, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000369, 5'd23, 27'h00000012, 5'd5, 27'h000000ef, 32'h00000400,
  1'd1,  5'd8, 27'h00000020, 5'd23, 27'h00000285, 5'd19, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000170, 5'd22, 27'h00000320, 5'd30, 27'h00000343, 32'h00000400,
  1'd1,  5'd17, 27'h0000029d, 5'd2, 27'h00000273, 5'd0, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000358, 5'd0, 27'h00000111, 5'd15, 27'h00000177, 32'h00000400,
  1'd1,  5'd16, 27'h00000275, 5'd4, 27'h000002ee, 5'd24, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ea, 5'd12, 27'h0000009b, 5'd7, 27'h00000023, 32'h00000400,
  1'd1,  5'd18, 27'h00000133, 5'd14, 27'h00000038, 5'd16, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000109, 5'd13, 27'h00000021, 5'd28, 27'h00000377, 32'h00000400,
  1'd1,  5'd16, 27'h000001ea, 5'd24, 27'h0000038a, 5'd10, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003fc, 5'd24, 27'h00000343, 5'd18, 27'h00000159, 32'h00000400,
  1'd1,  5'd20, 27'h0000009f, 5'd23, 27'h0000027d, 5'd29, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000033d, 5'd0, 27'h0000023a, 5'd7, 27'h0000001d, 32'h00000400,
  1'd1,  5'd30, 27'h00000045, 5'd1, 27'h000000d1, 5'd17, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a5, 5'd3, 27'h00000275, 5'd27, 27'h000002fa, 32'h00000400,
  1'd1,  5'd29, 27'h0000034a, 5'd13, 27'h000001c4, 5'd8, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001a2, 5'd15, 27'h0000009f, 5'd18, 27'h000002bc, 32'h00000400,
  1'd1,  5'd27, 27'h00000078, 5'd12, 27'h0000020e, 5'd29, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000331, 5'd25, 27'h00000078, 5'd7, 27'h000002a5, 32'h00000400,
  1'd1,  5'd30, 27'h000002fc, 5'd21, 27'h00000113, 5'd17, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000213, 5'd22, 27'h000002e9, 5'd28, 27'h00000161, 32'h00000400,
  1'd1,  5'd6, 27'h000002de, 5'd7, 27'h000002fd, 5'd1, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000034b, 5'd6, 27'h000001e5, 5'd11, 27'h0000000d, 32'h00000400,
  1'd1,  5'd8, 27'h000003fd, 5'd5, 27'h000000c0, 5'd21, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003de, 5'd17, 27'h000000f4, 5'd4, 27'h00000276, 32'h00000400,
  1'd1,  5'd8, 27'h00000007, 5'd17, 27'h00000224, 5'd13, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002db, 5'd15, 27'h000003f7, 5'd23, 27'h000002eb, 32'h00000400,
  1'd1,  5'd7, 27'h00000066, 5'd28, 27'h000003cd, 5'd0, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003aa, 5'd27, 27'h00000025, 5'd14, 27'h00000310, 32'h00000400,
  1'd1,  5'd8, 27'h000001bb, 5'd30, 27'h00000364, 5'd22, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001dd, 5'd5, 27'h0000015b, 5'd1, 27'h0000025e, 32'h00000400,
  1'd1,  5'd16, 27'h0000023f, 5'd5, 27'h00000390, 5'd10, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e5, 5'd6, 27'h000001e2, 5'd20, 27'h00000355, 32'h00000400,
  1'd1,  5'd19, 27'h00000048, 5'd16, 27'h000000b1, 5'd2, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000029b, 5'd16, 27'h000002e6, 5'd13, 27'h00000056, 32'h00000400,
  1'd1,  5'd18, 27'h0000029f, 5'd16, 27'h00000306, 5'd21, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039e, 5'd30, 27'h0000011b, 5'd3, 27'h00000279, 32'h00000400,
  1'd1,  5'd17, 27'h000002b2, 5'd26, 27'h000003f6, 5'd10, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000032, 5'd27, 27'h000003c4, 5'd22, 27'h000000a9, 32'h00000400,
  1'd1,  5'd27, 27'h0000027b, 5'd7, 27'h000003b2, 5'd4, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a8, 5'd7, 27'h00000002, 5'd15, 27'h00000124, 32'h00000400,
  1'd1,  5'd30, 27'h00000328, 5'd9, 27'h00000062, 5'd23, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000058, 5'd18, 27'h000001a0, 5'd0, 27'h000000fa, 32'h00000400,
  1'd1,  5'd30, 27'h0000026b, 5'd20, 27'h00000127, 5'd15, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000280, 5'd17, 27'h0000026b, 5'd22, 27'h00000119, 32'h00000400,
  1'd1,  5'd26, 27'h00000360, 5'd26, 27'h000003eb, 5'd2, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000044, 5'd27, 27'h00000352, 5'd12, 27'h0000018d, 32'h00000400,
  1'd1,  5'd27, 27'h00000371, 5'd28, 27'h00000223, 5'd22, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000040, 5'd5, 27'h000003e6, 5'd7, 27'h0000003c, 32'h00000400,
  1'd1,  5'd6, 27'h0000003e, 5'd9, 27'h00000304, 5'd19, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001e2, 5'd7, 27'h0000026d, 5'd26, 27'h00000045, 32'h00000400,
  1'd1,  5'd6, 27'h0000036c, 5'd18, 27'h00000163, 5'd8, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005e, 5'd17, 27'h00000178, 5'd16, 27'h0000039a, 32'h00000400,
  1'd1,  5'd5, 27'h000001b4, 5'd19, 27'h00000344, 5'd29, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d8, 5'd27, 27'h0000015a, 5'd9, 27'h00000071, 32'h00000400,
  1'd1,  5'd7, 27'h00000227, 5'd30, 27'h00000285, 5'd16, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000125, 5'd30, 27'h00000313, 5'd28, 27'h00000142, 32'h00000400,
  1'd1,  5'd18, 27'h00000289, 5'd8, 27'h000001b7, 5'd8, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000265, 5'd7, 27'h000001ce, 5'd16, 27'h00000197, 32'h00000400,
  1'd1,  5'd16, 27'h000003e2, 5'd9, 27'h000003df, 5'd26, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000258, 5'd17, 27'h000001e8, 5'd6, 27'h000001b7, 32'h00000400,
  1'd1,  5'd15, 27'h00000384, 5'd17, 27'h000000ad, 5'd20, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000027c, 5'd18, 27'h0000018e, 5'd26, 27'h0000008b, 32'h00000400,
  1'd1,  5'd16, 27'h00000175, 5'd26, 27'h00000010, 5'd10, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000228, 5'd30, 27'h00000069, 5'd18, 27'h00000213, 32'h00000400,
  1'd1,  5'd17, 27'h000003ad, 5'd29, 27'h00000313, 5'd27, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000008b, 5'd9, 27'h00000213, 5'd5, 27'h000002fa, 32'h00000400,
  1'd1,  5'd26, 27'h00000279, 5'd8, 27'h00000329, 5'd20, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ad, 5'd8, 27'h000003b9, 5'd29, 27'h00000326, 32'h00000400,
  1'd1,  5'd26, 27'h000002fd, 5'd19, 27'h00000387, 5'd8, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d5, 5'd15, 27'h0000025b, 5'd17, 27'h0000012a, 32'h00000400,
  1'd1,  5'd27, 27'h0000019f, 5'd17, 27'h000000af, 5'd27, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000018f, 5'd29, 27'h000002bf, 5'd8, 27'h00000153, 32'h00000400,
  1'd1,  5'd29, 27'h00000125, 5'd29, 27'h0000015d, 5'd15, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000110, 5'd27, 27'h00000241, 5'd29, 27'h0000016f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000243, 5'd2, 27'h0000006a, 5'd1, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014c, 5'd2, 27'h000003ad, 5'd14, 27'h000003e9, 32'h00000400,
  1'd1,  5'd2, 27'h000002d6, 5'd4, 27'h000003d5, 5'd22, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000016e, 5'd12, 27'h0000025a, 5'd3, 27'h0000037d, 32'h00000400,
  1'd1,  5'd0, 27'h0000019b, 5'd11, 27'h000000c1, 5'd12, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001f1, 5'd12, 27'h00000389, 5'd24, 27'h0000015f, 32'h00000400,
  1'd1,  5'd1, 27'h0000028c, 5'd21, 27'h00000001, 5'd2, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ae, 5'd24, 27'h00000162, 5'd15, 27'h000001aa, 32'h00000400,
  1'd1,  5'd4, 27'h00000105, 5'd21, 27'h0000014a, 5'd23, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000035, 5'd3, 27'h00000392, 5'd2, 27'h0000012a, 32'h00000400,
  1'd1,  5'd11, 27'h000000ae, 5'd2, 27'h0000030f, 5'd12, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001da, 5'd3, 27'h0000037c, 5'd24, 27'h000003de, 32'h00000400,
  1'd1,  5'd15, 27'h00000017, 5'd11, 27'h00000171, 5'd4, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002c, 5'd10, 27'h00000201, 5'd13, 27'h000003ba, 32'h00000400,
  1'd1,  5'd11, 27'h000002ee, 5'd12, 27'h00000149, 5'd25, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000368, 5'd21, 27'h00000274, 5'd0, 27'h0000002d, 32'h00000400,
  1'd1,  5'd11, 27'h000002f6, 5'd21, 27'h00000292, 5'd14, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000022b, 5'd22, 27'h00000032, 5'd21, 27'h000000cc, 32'h00000400,
  1'd1,  5'd22, 27'h000003c8, 5'd2, 27'h0000025a, 5'd0, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b0, 5'd0, 27'h00000365, 5'd14, 27'h00000395, 32'h00000400,
  1'd1,  5'd23, 27'h000000cf, 5'd0, 27'h000000bf, 5'd23, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000114, 5'd12, 27'h0000014d, 5'd3, 27'h00000315, 32'h00000400,
  1'd1,  5'd21, 27'h000001ed, 5'd14, 27'h0000003d, 5'd11, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000154, 5'd10, 27'h00000367, 5'd23, 27'h000001b0, 32'h00000400,
  1'd1,  5'd24, 27'h00000260, 5'd23, 27'h00000264, 5'd2, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000360, 5'd22, 27'h0000017a, 5'd10, 27'h000002b4, 32'h00000400,
  1'd1,  5'd22, 27'h0000002d, 5'd22, 27'h0000011d, 5'd22, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000030b, 5'd2, 27'h000002de, 5'd6, 27'h0000030c, 32'h00000400,
  1'd1,  5'd2, 27'h0000014a, 5'd0, 27'h00000069, 5'd17, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000aa, 5'd1, 27'h000001c7, 5'd30, 27'h000001bf, 32'h00000400,
  1'd1,  5'd2, 27'h0000002e, 5'd10, 27'h000001d9, 5'd10, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002f0, 5'd10, 27'h0000027e, 5'd19, 27'h00000141, 32'h00000400,
  1'd1,  5'd1, 27'h00000198, 5'd14, 27'h00000104, 5'd28, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000315, 5'd25, 27'h00000086, 5'd8, 27'h00000349, 32'h00000400,
  1'd1,  5'd0, 27'h00000253, 5'd21, 27'h00000303, 5'd18, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d7, 5'd23, 27'h00000249, 5'd29, 27'h0000025a, 32'h00000400,
  1'd1,  5'd13, 27'h000000ed, 5'd0, 27'h00000153, 5'd9, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000132, 5'd0, 27'h00000096, 5'd16, 27'h00000179, 32'h00000400,
  1'd1,  5'd11, 27'h00000117, 5'd0, 27'h0000033d, 5'd29, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f0, 5'd13, 27'h00000172, 5'd7, 27'h000000e7, 32'h00000400,
  1'd1,  5'd14, 27'h00000195, 5'd13, 27'h00000065, 5'd15, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000eb, 5'd15, 27'h000000f0, 5'd26, 27'h00000316, 32'h00000400,
  1'd1,  5'd10, 27'h000002a3, 5'd22, 27'h00000055, 5'd6, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f5, 5'd25, 27'h00000263, 5'd16, 27'h000002dd, 32'h00000400,
  1'd1,  5'd14, 27'h00000158, 5'd25, 27'h00000337, 5'd25, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e0, 5'd2, 27'h000000dd, 5'd5, 27'h00000287, 32'h00000400,
  1'd1,  5'd22, 27'h000001d9, 5'd2, 27'h00000389, 5'd17, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003b9, 5'd1, 27'h000003e9, 5'd28, 27'h00000036, 32'h00000400,
  1'd1,  5'd21, 27'h00000354, 5'd10, 27'h00000333, 5'd6, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a5, 5'd13, 27'h00000215, 5'd20, 27'h00000046, 32'h00000400,
  1'd1,  5'd23, 27'h0000007a, 5'd13, 27'h000000a4, 5'd29, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ba, 5'd21, 27'h00000290, 5'd9, 27'h0000015b, 32'h00000400,
  1'd1,  5'd23, 27'h000000af, 5'd24, 27'h00000127, 5'd16, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000250, 5'd23, 27'h0000003a, 5'd28, 27'h000001b7, 32'h00000400,
  1'd1,  5'd1, 27'h000003f0, 5'd5, 27'h000002b5, 5'd2, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a7, 5'd7, 27'h000000bc, 5'd15, 27'h000000d3, 32'h00000400,
  1'd1,  5'd2, 27'h00000050, 5'd8, 27'h00000250, 5'd21, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000023, 5'd16, 27'h000000a8, 5'd1, 27'h0000018d, 32'h00000400,
  1'd1,  5'd3, 27'h0000006e, 5'd18, 27'h00000182, 5'd13, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b8, 5'd17, 27'h000001d1, 5'd22, 27'h0000028d, 32'h00000400,
  1'd1,  5'd0, 27'h0000011d, 5'd26, 27'h00000234, 5'd0, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000009a, 5'd27, 27'h000000bd, 5'd13, 27'h00000126, 32'h00000400,
  1'd1,  5'd5, 27'h00000013, 5'd27, 27'h00000283, 5'd21, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000d0, 5'd6, 27'h00000008, 5'd0, 27'h0000026c, 32'h00000400,
  1'd1,  5'd14, 27'h00000355, 5'd8, 27'h0000028d, 5'd14, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003e1, 5'd10, 27'h000000ab, 5'd25, 27'h0000012a, 32'h00000400,
  1'd1,  5'd13, 27'h000003f9, 5'd17, 27'h00000381, 5'd3, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002c6, 5'd17, 27'h000001fd, 5'd10, 27'h00000330, 32'h00000400,
  1'd1,  5'd12, 27'h0000026e, 5'd16, 27'h0000007e, 5'd23, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013b, 5'd30, 27'h000002ca, 5'd0, 27'h000002e6, 32'h00000400,
  1'd1,  5'd10, 27'h00000243, 5'd26, 27'h000000a9, 5'd12, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ad, 5'd26, 27'h00000296, 5'd25, 27'h00000162, 32'h00000400,
  1'd1,  5'd23, 27'h000003cf, 5'd10, 27'h0000008f, 5'd3, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a9, 5'd10, 27'h00000127, 5'd14, 27'h0000026a, 32'h00000400,
  1'd1,  5'd22, 27'h000002d0, 5'd10, 27'h00000083, 5'd24, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000345, 5'd15, 27'h000002f3, 5'd1, 27'h0000013d, 32'h00000400,
  1'd1,  5'd23, 27'h000002ed, 5'd16, 27'h000003d3, 5'd12, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031d, 5'd19, 27'h00000144, 5'd25, 27'h00000234, 32'h00000400,
  1'd1,  5'd21, 27'h0000020b, 5'd27, 27'h00000282, 5'd2, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001bd, 5'd30, 27'h00000212, 5'd11, 27'h00000226, 32'h00000400,
  1'd1,  5'd24, 27'h00000210, 5'd26, 27'h00000028, 5'd20, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000008a, 5'd8, 27'h00000386, 5'd9, 27'h000003b4, 32'h00000400,
  1'd1,  5'd1, 27'h0000007e, 5'd10, 27'h00000012, 5'd20, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000103, 5'd9, 27'h000001b5, 5'd30, 27'h00000282, 32'h00000400,
  1'd1,  5'd2, 27'h000003f5, 5'd19, 27'h000002bb, 5'd7, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c3, 5'd18, 27'h000002f1, 5'd16, 27'h0000024b, 32'h00000400,
  1'd1,  5'd2, 27'h000001e3, 5'd16, 27'h0000019b, 5'd29, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000019a, 5'd29, 27'h0000022c, 5'd7, 27'h00000236, 32'h00000400,
  1'd1,  5'd1, 27'h00000365, 5'd30, 27'h0000020c, 5'd17, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003d5, 5'd26, 27'h000001a2, 5'd27, 27'h000000fb, 32'h00000400,
  1'd1,  5'd14, 27'h00000397, 5'd7, 27'h00000277, 5'd7, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000152, 5'd8, 27'h00000223, 5'd20, 27'h000001d7, 32'h00000400,
  1'd1,  5'd11, 27'h00000278, 5'd9, 27'h0000024a, 5'd28, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000d7, 5'd17, 27'h0000039f, 5'd9, 27'h00000075, 32'h00000400,
  1'd1,  5'd11, 27'h0000035e, 5'd19, 27'h0000025b, 5'd18, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000108, 5'd17, 27'h0000024c, 5'd30, 27'h00000228, 32'h00000400,
  1'd1,  5'd12, 27'h00000396, 5'd26, 27'h00000297, 5'd6, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000190, 5'd29, 27'h0000012a, 5'd16, 27'h00000257, 32'h00000400,
  1'd1,  5'd12, 27'h000003e3, 5'd27, 27'h000001d6, 5'd28, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000031f, 5'd10, 27'h0000004f, 5'd9, 27'h0000001b, 32'h00000400,
  1'd1,  5'd24, 27'h00000020, 5'd5, 27'h0000029a, 5'd16, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d4, 5'd5, 27'h000000c4, 5'd27, 27'h000002cb, 32'h00000400,
  1'd1,  5'd24, 27'h00000377, 5'd15, 27'h0000024b, 5'd6, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000010f, 5'd18, 27'h0000008c, 5'd20, 27'h00000091, 32'h00000400,
  1'd1,  5'd24, 27'h00000141, 5'd19, 27'h0000027b, 5'd30, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000134, 5'd28, 27'h000002d1, 5'd6, 27'h000002a1, 32'h00000400,
  1'd1,  5'd20, 27'h00000342, 5'd26, 27'h000000af, 5'd16, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002eb, 5'd29, 27'h00000039, 5'd27, 27'h0000008b, 32'h00000400,
  1'd1,  5'd9, 27'h000001a9, 5'd2, 27'h0000018b, 5'd8, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000356, 5'd3, 27'h000000e0, 5'd16, 27'h0000028f, 32'h00000400,
  1'd1,  5'd5, 27'h000003a6, 5'd2, 27'h000003d1, 5'd26, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000008d, 5'd11, 27'h000001c1, 5'd1, 27'h00000370, 32'h00000400,
  1'd1,  5'd7, 27'h00000050, 5'd13, 27'h000003aa, 5'd12, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000033d, 5'd12, 27'h000001bb, 5'd22, 27'h00000031, 32'h00000400,
  1'd1,  5'd7, 27'h00000136, 5'd23, 27'h000001e8, 5'd1, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000263, 5'd23, 27'h0000010d, 5'd10, 27'h000001be, 32'h00000400,
  1'd1,  5'd7, 27'h00000063, 5'd22, 27'h000002b0, 5'd22, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a7, 5'd0, 27'h00000346, 5'd7, 27'h00000162, 32'h00000400,
  1'd1,  5'd17, 27'h0000022f, 5'd2, 27'h000000d3, 5'd19, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000029d, 5'd3, 27'h00000088, 5'd25, 27'h00000379, 32'h00000400,
  1'd1,  5'd20, 27'h00000152, 5'd14, 27'h00000141, 5'd4, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ef, 5'd14, 27'h0000031e, 5'd13, 27'h000001d2, 32'h00000400,
  1'd1,  5'd16, 27'h000001e1, 5'd11, 27'h000003c9, 5'd25, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000323, 5'd22, 27'h0000008f, 5'd1, 27'h0000027c, 32'h00000400,
  1'd1,  5'd17, 27'h000003f4, 5'd22, 27'h00000381, 5'd12, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000fb, 5'd25, 27'h00000060, 5'd21, 27'h0000026d, 32'h00000400,
  1'd1,  5'd29, 27'h00000331, 5'd3, 27'h000000f7, 5'd2, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000190, 5'd3, 27'h0000016f, 5'd14, 27'h000001c1, 32'h00000400,
  1'd1,  5'd30, 27'h000000d9, 5'd0, 27'h000002ac, 5'd25, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b5, 5'd12, 27'h000003fd, 5'd2, 27'h00000128, 32'h00000400,
  1'd1,  5'd25, 27'h000003b2, 5'd10, 27'h00000341, 5'd13, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b0, 5'd15, 27'h000000b8, 5'd23, 27'h00000304, 32'h00000400,
  1'd1,  5'd29, 27'h0000029a, 5'd22, 27'h000000c4, 5'd3, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000be, 5'd21, 27'h000003d2, 5'd11, 27'h000000c3, 32'h00000400,
  1'd1,  5'd29, 27'h000002f3, 5'd21, 27'h00000117, 5'd25, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038c, 5'd0, 27'h00000391, 5'd2, 27'h00000071, 32'h00000400,
  1'd1,  5'd7, 27'h0000026f, 5'd4, 27'h000001fe, 5'd12, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000214, 5'd0, 27'h00000385, 5'd24, 27'h000000b9, 32'h00000400,
  1'd1,  5'd5, 27'h0000022c, 5'd12, 27'h00000293, 5'd7, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000d5, 5'd14, 27'h0000011b, 5'd18, 27'h000003f6, 32'h00000400,
  1'd1,  5'd7, 27'h000002dd, 5'd13, 27'h00000046, 5'd29, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000210, 5'd24, 27'h000003c3, 5'd6, 27'h000001aa, 32'h00000400,
  1'd1,  5'd5, 27'h0000039d, 5'd24, 27'h0000019f, 5'd16, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000363, 5'd21, 27'h00000158, 5'd26, 27'h000001fd, 32'h00000400,
  1'd1,  5'd17, 27'h0000032b, 5'd1, 27'h00000140, 5'd0, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000169, 5'd1, 27'h00000350, 5'd11, 27'h00000371, 32'h00000400,
  1'd1,  5'd19, 27'h00000135, 5'd3, 27'h000002d9, 5'd23, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000008b, 5'd13, 27'h000000f2, 5'd7, 27'h000001b1, 32'h00000400,
  1'd1,  5'd17, 27'h00000083, 5'd11, 27'h0000039d, 5'd16, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000079, 5'd14, 27'h00000192, 5'd27, 27'h00000185, 32'h00000400,
  1'd1,  5'd18, 27'h0000026f, 5'd25, 27'h000002cd, 5'd8, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000399, 5'd24, 27'h00000310, 5'd17, 27'h00000266, 32'h00000400,
  1'd1,  5'd17, 27'h000001f4, 5'd23, 27'h0000024d, 5'd29, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d4, 5'd3, 27'h00000193, 5'd9, 27'h00000199, 32'h00000400,
  1'd1,  5'd27, 27'h0000032f, 5'd0, 27'h000002b7, 5'd18, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000347, 5'd0, 27'h0000016e, 5'd29, 27'h000000f3, 32'h00000400,
  1'd1,  5'd28, 27'h00000336, 5'd12, 27'h000002a2, 5'd7, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000276, 5'd12, 27'h000000c0, 5'd16, 27'h000000b6, 32'h00000400,
  1'd1,  5'd29, 27'h00000069, 5'd14, 27'h00000295, 5'd30, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000b3, 5'd23, 27'h0000021b, 5'd6, 27'h00000168, 32'h00000400,
  1'd1,  5'd25, 27'h000003ef, 5'd22, 27'h0000034f, 5'd17, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000396, 5'd22, 27'h0000010c, 5'd29, 27'h0000029d, 32'h00000400,
  1'd1,  5'd7, 27'h0000033a, 5'd5, 27'h000001d4, 5'd3, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000227, 5'd8, 27'h000003f1, 5'd11, 27'h0000038a, 32'h00000400,
  1'd1,  5'd7, 27'h0000022a, 5'd10, 27'h00000133, 5'd23, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a2, 5'd16, 27'h0000006a, 5'd4, 27'h000001cc, 32'h00000400,
  1'd1,  5'd7, 27'h00000364, 5'd19, 27'h000002a5, 5'd13, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000035, 5'd16, 27'h0000011b, 5'd23, 27'h000000d7, 32'h00000400,
  1'd1,  5'd9, 27'h00000131, 5'd30, 27'h000001aa, 5'd3, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000175, 5'd29, 27'h0000011c, 5'd11, 27'h0000019c, 32'h00000400,
  1'd1,  5'd7, 27'h000001ea, 5'd29, 27'h000001db, 5'd22, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ba, 5'd7, 27'h00000309, 5'd1, 27'h0000036f, 32'h00000400,
  1'd1,  5'd20, 27'h0000020c, 5'd9, 27'h000003f7, 5'd13, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000220, 5'd7, 27'h00000270, 5'd22, 27'h000003bf, 32'h00000400,
  1'd1,  5'd18, 27'h000002e9, 5'd16, 27'h000003b8, 5'd0, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000245, 5'd18, 27'h00000273, 5'd11, 27'h00000357, 32'h00000400,
  1'd1,  5'd16, 27'h00000223, 5'd19, 27'h00000143, 5'd23, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003d6, 5'd28, 27'h000002f1, 5'd3, 27'h00000351, 32'h00000400,
  1'd1,  5'd20, 27'h0000010a, 5'd28, 27'h0000003e, 5'd10, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000227, 5'd26, 27'h000002b2, 5'd25, 27'h00000236, 32'h00000400,
  1'd1,  5'd28, 27'h000001fc, 5'd9, 27'h00000325, 5'd2, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000277, 5'd6, 27'h00000240, 5'd13, 27'h000000b8, 32'h00000400,
  1'd1,  5'd29, 27'h000002c4, 5'd8, 27'h000002fc, 5'd23, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ba, 5'd19, 27'h00000206, 5'd2, 27'h000000b7, 32'h00000400,
  1'd1,  5'd26, 27'h000002ba, 5'd18, 27'h0000026b, 5'd12, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000383, 5'd18, 27'h00000038, 5'd21, 27'h000002c7, 32'h00000400,
  1'd1,  5'd28, 27'h00000254, 5'd29, 27'h0000006f, 5'd0, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000375, 5'd27, 27'h0000016d, 5'd11, 27'h000002f7, 32'h00000400,
  1'd1,  5'd30, 27'h0000004d, 5'd30, 27'h00000338, 5'd20, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000151, 5'd7, 27'h00000103, 5'd9, 27'h00000355, 32'h00000400,
  1'd1,  5'd9, 27'h00000065, 5'd7, 27'h00000223, 5'd18, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000377, 5'd7, 27'h00000130, 5'd26, 27'h00000120, 32'h00000400,
  1'd1,  5'd9, 27'h00000308, 5'd15, 27'h00000325, 5'd9, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000027b, 5'd16, 27'h00000279, 5'd17, 27'h0000002c, 32'h00000400,
  1'd1,  5'd6, 27'h000000ab, 5'd17, 27'h00000329, 5'd26, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000008f, 5'd27, 27'h000000f3, 5'd10, 27'h000000c0, 32'h00000400,
  1'd1,  5'd5, 27'h000001de, 5'd27, 27'h000002c2, 5'd17, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000015d, 5'd28, 27'h00000243, 5'd30, 27'h00000201, 32'h00000400,
  1'd1,  5'd19, 27'h0000018b, 5'd5, 27'h0000033f, 5'd5, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000030f, 5'd9, 27'h0000035d, 5'd18, 27'h0000035f, 32'h00000400,
  1'd1,  5'd16, 27'h000002ee, 5'd7, 27'h0000003e, 5'd26, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000091, 5'd18, 27'h000000e1, 5'd7, 27'h000003a8, 32'h00000400,
  1'd1,  5'd16, 27'h000002c2, 5'd17, 27'h00000318, 5'd19, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001fe, 5'd17, 27'h0000008b, 5'd29, 27'h0000002c, 32'h00000400,
  1'd1,  5'd17, 27'h00000186, 5'd27, 27'h0000034a, 5'd6, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000070, 5'd29, 27'h000003d1, 5'd20, 27'h00000086, 32'h00000400,
  1'd1,  5'd20, 27'h00000221, 5'd30, 27'h000000fe, 5'd26, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003c9, 5'd5, 27'h00000119, 5'd7, 27'h000001af, 32'h00000400,
  1'd1,  5'd30, 27'h000001ca, 5'd7, 27'h000002b2, 5'd19, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021a, 5'd9, 27'h000000b8, 5'd29, 27'h0000009f, 32'h00000400,
  1'd1,  5'd27, 27'h0000017d, 5'd18, 27'h000002ee, 5'd5, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000066, 5'd16, 27'h0000018d, 5'd18, 27'h00000321, 32'h00000400,
  1'd1,  5'd28, 27'h000003f8, 5'd15, 27'h000003e0, 5'd26, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000031a, 5'd29, 27'h00000108, 5'd6, 27'h000000f5, 32'h00000400,
  1'd1,  5'd26, 27'h000003e5, 5'd30, 27'h000003bd, 5'd16, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000000d, 5'd27, 27'h00000393, 5'd26, 27'h000003b2, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000032f, 5'd2, 27'h000000d8, 5'd1, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000014, 5'd1, 27'h0000025b, 5'd14, 27'h000000e8, 32'h00000400,
  1'd1,  5'd3, 27'h000002ef, 5'd2, 27'h00000299, 5'd22, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f6, 5'd11, 27'h00000168, 5'd4, 27'h00000220, 32'h00000400,
  1'd1,  5'd2, 27'h0000016e, 5'd14, 27'h00000200, 5'd14, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001bb, 5'd14, 27'h000002b9, 5'd20, 27'h000003d2, 32'h00000400,
  1'd1,  5'd4, 27'h000001d3, 5'd25, 27'h00000007, 5'd3, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000152, 5'd22, 27'h00000095, 5'd13, 27'h000000f9, 32'h00000400,
  1'd1,  5'd4, 27'h000002aa, 5'd25, 27'h00000005, 5'd21, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000023, 5'd1, 27'h000002b9, 5'd1, 27'h0000010a, 32'h00000400,
  1'd1,  5'd12, 27'h0000014b, 5'd0, 27'h00000219, 5'd13, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e6, 5'd3, 27'h00000221, 5'd22, 27'h000002cf, 32'h00000400,
  1'd1,  5'd14, 27'h000002e6, 5'd14, 27'h00000293, 5'd0, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000061, 5'd11, 27'h0000038f, 5'd14, 27'h00000165, 32'h00000400,
  1'd1,  5'd11, 27'h00000125, 5'd14, 27'h0000035f, 5'd21, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000030f, 5'd21, 27'h00000228, 5'd3, 27'h000001f8, 32'h00000400,
  1'd1,  5'd13, 27'h0000033a, 5'd23, 27'h0000016e, 5'd11, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003eb, 5'd24, 27'h00000061, 5'd23, 27'h000000d2, 32'h00000400,
  1'd1,  5'd22, 27'h00000341, 5'd2, 27'h000002f8, 5'd0, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000345, 5'd2, 27'h00000172, 5'd11, 27'h000002c9, 32'h00000400,
  1'd1,  5'd23, 27'h00000114, 5'd3, 27'h0000019c, 5'd25, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001fc, 5'd14, 27'h00000250, 5'd4, 27'h0000020b, 32'h00000400,
  1'd1,  5'd20, 27'h000002f5, 5'd10, 27'h00000209, 5'd13, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000034, 5'd11, 27'h000000ad, 5'd24, 27'h00000121, 32'h00000400,
  1'd1,  5'd24, 27'h000002dd, 5'd24, 27'h0000032b, 5'd1, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000304, 5'd23, 27'h00000038, 5'd12, 27'h00000326, 32'h00000400,
  1'd1,  5'd22, 27'h0000016d, 5'd25, 27'h000000b6, 5'd21, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000008e, 5'd4, 27'h0000005b, 5'd6, 27'h0000021b, 32'h00000400,
  1'd1,  5'd4, 27'h00000288, 5'd1, 27'h000001e4, 5'd17, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000384, 5'd1, 27'h000002df, 5'd27, 27'h00000279, 32'h00000400,
  1'd1,  5'd3, 27'h00000231, 5'd14, 27'h00000089, 5'd6, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000c6, 5'd12, 27'h00000107, 5'd20, 27'h0000024c, 32'h00000400,
  1'd1,  5'd1, 27'h000001b4, 5'd11, 27'h00000227, 5'd28, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000024b, 5'd22, 27'h000003ea, 5'd7, 27'h000002de, 32'h00000400,
  1'd1,  5'd1, 27'h000003b7, 5'd21, 27'h000000b7, 5'd18, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000005, 5'd20, 27'h000002ad, 5'd28, 27'h000001c1, 32'h00000400,
  1'd1,  5'd14, 27'h00000281, 5'd4, 27'h00000211, 5'd9, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000318, 5'd2, 27'h00000337, 5'd17, 27'h0000013b, 32'h00000400,
  1'd1,  5'd12, 27'h0000003c, 5'd0, 27'h000000c7, 5'd28, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000038b, 5'd14, 27'h000001ad, 5'd8, 27'h00000272, 32'h00000400,
  1'd1,  5'd11, 27'h000002d1, 5'd15, 27'h00000066, 5'd17, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000386, 5'd13, 27'h000000dc, 5'd28, 27'h0000001f, 32'h00000400,
  1'd1,  5'd13, 27'h0000030a, 5'd25, 27'h0000000d, 5'd8, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002bb, 5'd25, 27'h000002aa, 5'd19, 27'h000002a3, 32'h00000400,
  1'd1,  5'd12, 27'h00000114, 5'd22, 27'h00000246, 5'd26, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002b0, 5'd1, 27'h00000316, 5'd5, 27'h000001f6, 32'h00000400,
  1'd1,  5'd24, 27'h00000359, 5'd1, 27'h000002d5, 5'd17, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002cc, 5'd1, 27'h000003da, 5'd26, 27'h0000018f, 32'h00000400,
  1'd1,  5'd22, 27'h000000ec, 5'd11, 27'h000000fa, 5'd9, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000013a, 5'd11, 27'h00000201, 5'd16, 27'h00000042, 32'h00000400,
  1'd1,  5'd25, 27'h0000007e, 5'd12, 27'h000002d3, 5'd26, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000309, 5'd22, 27'h0000038b, 5'd6, 27'h0000004f, 32'h00000400,
  1'd1,  5'd22, 27'h0000025e, 5'd22, 27'h0000013f, 5'd19, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000312, 5'd23, 27'h00000187, 5'd25, 27'h0000038a, 32'h00000400,
  1'd1,  5'd2, 27'h0000011b, 5'd7, 27'h000001c8, 5'd1, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000081, 5'd10, 27'h00000021, 5'd13, 27'h00000326, 32'h00000400,
  1'd1,  5'd3, 27'h00000108, 5'd5, 27'h00000261, 5'd21, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000002b, 5'd19, 27'h00000255, 5'd1, 27'h0000018d, 32'h00000400,
  1'd1,  5'd0, 27'h000000d6, 5'd17, 27'h0000003a, 5'd14, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000111, 5'd20, 27'h00000257, 5'd22, 27'h000003fe, 32'h00000400,
  1'd1,  5'd2, 27'h0000026f, 5'd30, 27'h000002cc, 5'd2, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000f3, 5'd28, 27'h00000110, 5'd11, 27'h00000259, 32'h00000400,
  1'd1,  5'd5, 27'h00000024, 5'd29, 27'h00000196, 5'd23, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000304, 5'd6, 27'h00000276, 5'd1, 27'h000001e9, 32'h00000400,
  1'd1,  5'd14, 27'h00000285, 5'd7, 27'h0000007c, 5'd12, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000013e, 5'd9, 27'h000001ad, 5'd23, 27'h000000cc, 32'h00000400,
  1'd1,  5'd14, 27'h00000274, 5'd17, 27'h000003c7, 5'd2, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000083, 5'd20, 27'h0000010d, 5'd11, 27'h00000274, 32'h00000400,
  1'd1,  5'd14, 27'h000003aa, 5'd15, 27'h000003e2, 5'd21, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000fe, 5'd30, 27'h000002c8, 5'd4, 27'h00000295, 32'h00000400,
  1'd1,  5'd14, 27'h00000009, 5'd30, 27'h000000ab, 5'd10, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000005d, 5'd29, 27'h000001eb, 5'd25, 27'h000000de, 32'h00000400,
  1'd1,  5'd24, 27'h0000009b, 5'd10, 27'h00000087, 5'd3, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000018c, 5'd7, 27'h000002d0, 5'd14, 27'h00000145, 32'h00000400,
  1'd1,  5'd22, 27'h00000272, 5'd9, 27'h00000309, 5'd23, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e6, 5'd18, 27'h000001e8, 5'd3, 27'h00000385, 32'h00000400,
  1'd1,  5'd25, 27'h00000332, 5'd20, 27'h0000017f, 5'd15, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ea, 5'd16, 27'h000002af, 5'd24, 27'h000000cb, 32'h00000400,
  1'd1,  5'd24, 27'h000001c7, 5'd28, 27'h000000fb, 5'd3, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001dd, 5'd30, 27'h00000249, 5'd11, 27'h00000018, 32'h00000400,
  1'd1,  5'd25, 27'h00000081, 5'd28, 27'h000002a4, 5'd25, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001fb, 5'd5, 27'h000000cc, 5'd6, 27'h000002c0, 32'h00000400,
  1'd1,  5'd4, 27'h000003e0, 5'd9, 27'h00000136, 5'd18, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000268, 5'd9, 27'h000000f2, 5'd29, 27'h00000378, 32'h00000400,
  1'd1,  5'd2, 27'h00000237, 5'd18, 27'h0000003f, 5'd10, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e7, 5'd17, 27'h000002f2, 5'd19, 27'h000000bb, 32'h00000400,
  1'd1,  5'd2, 27'h000001b0, 5'd16, 27'h00000295, 5'd25, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000fb, 5'd28, 27'h000003a5, 5'd7, 27'h000001d7, 32'h00000400,
  1'd1,  5'd3, 27'h00000118, 5'd30, 27'h0000030f, 5'd16, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ba, 5'd27, 27'h000001d2, 5'd27, 27'h0000039f, 32'h00000400,
  1'd1,  5'd11, 27'h00000108, 5'd5, 27'h000003d6, 5'd6, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d7, 5'd8, 27'h0000020c, 5'd15, 27'h00000354, 32'h00000400,
  1'd1,  5'd11, 27'h0000018a, 5'd5, 27'h0000011c, 5'd27, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000381, 5'd16, 27'h00000012, 5'd7, 27'h000003de, 32'h00000400,
  1'd1,  5'd10, 27'h000001e6, 5'd17, 27'h000000b1, 5'd16, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000038d, 5'd18, 27'h000000c9, 5'd27, 27'h00000154, 32'h00000400,
  1'd1,  5'd15, 27'h000001e8, 5'd27, 27'h0000033f, 5'd7, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e5, 5'd28, 27'h000002a6, 5'd18, 27'h00000065, 32'h00000400,
  1'd1,  5'd13, 27'h00000136, 5'd28, 27'h000002a8, 5'd28, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000138, 5'd8, 27'h0000007c, 5'd6, 27'h00000121, 32'h00000400,
  1'd1,  5'd20, 27'h0000035f, 5'd6, 27'h000002c7, 5'd18, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000023f, 5'd5, 27'h000001fd, 5'd30, 27'h00000270, 32'h00000400,
  1'd1,  5'd21, 27'h0000027f, 5'd18, 27'h00000239, 5'd8, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000225, 5'd18, 27'h0000006a, 5'd18, 27'h000003cd, 32'h00000400,
  1'd1,  5'd25, 27'h00000008, 5'd16, 27'h0000036b, 5'd25, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000002b, 5'd30, 27'h000002a8, 5'd7, 27'h000003d7, 32'h00000400,
  1'd1,  5'd20, 27'h000002be, 5'd26, 27'h0000034c, 5'd19, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003a0, 5'd30, 27'h0000029a, 5'd30, 27'h000001c4, 32'h00000400,
  1'd1,  5'd5, 27'h000002b1, 5'd0, 27'h000002a8, 5'd10, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e9, 5'd2, 27'h00000310, 5'd19, 27'h000000cf, 32'h00000400,
  1'd1,  5'd7, 27'h000001a9, 5'd3, 27'h00000220, 5'd29, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000175, 5'd13, 27'h00000230, 5'd2, 27'h00000063, 32'h00000400,
  1'd1,  5'd7, 27'h0000037c, 5'd14, 27'h000003d7, 5'd13, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000020e, 5'd11, 27'h0000007b, 5'd24, 27'h00000250, 32'h00000400,
  1'd1,  5'd9, 27'h00000089, 5'd24, 27'h0000025e, 5'd3, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002cb, 5'd20, 27'h00000394, 5'd14, 27'h00000274, 32'h00000400,
  1'd1,  5'd10, 27'h0000002d, 5'd24, 27'h000002a8, 5'd25, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000098, 5'd1, 27'h00000262, 5'd6, 27'h000002d2, 32'h00000400,
  1'd1,  5'd17, 27'h0000038d, 5'd3, 27'h0000003c, 5'd16, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000035b, 5'd3, 27'h000003cf, 5'd27, 27'h0000034f, 32'h00000400,
  1'd1,  5'd17, 27'h00000143, 5'd11, 27'h00000126, 5'd4, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000023d, 5'd12, 27'h00000007, 5'd11, 27'h000001e8, 32'h00000400,
  1'd1,  5'd16, 27'h000000ae, 5'd14, 27'h00000031, 5'd24, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000381, 5'd22, 27'h00000328, 5'd3, 27'h00000218, 32'h00000400,
  1'd1,  5'd18, 27'h000003e1, 5'd25, 27'h0000020b, 5'd12, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000092, 5'd21, 27'h00000221, 5'd21, 27'h00000319, 32'h00000400,
  1'd1,  5'd30, 27'h000001b0, 5'd3, 27'h00000133, 5'd4, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000061, 5'd3, 27'h00000069, 5'd11, 27'h00000071, 32'h00000400,
  1'd1,  5'd29, 27'h00000385, 5'd3, 27'h00000209, 5'd25, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000206, 5'd12, 27'h0000003c, 5'd1, 27'h0000029c, 32'h00000400,
  1'd1,  5'd26, 27'h0000005e, 5'd15, 27'h000001d0, 5'd12, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000339, 5'd15, 27'h00000061, 5'd22, 27'h0000004a, 32'h00000400,
  1'd1,  5'd26, 27'h00000235, 5'd22, 27'h000001f0, 5'd0, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f8, 5'd21, 27'h000001b0, 5'd13, 27'h00000238, 32'h00000400,
  1'd1,  5'd28, 27'h00000274, 5'd22, 27'h00000087, 5'd23, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000000b, 5'd2, 27'h000001ad, 5'd0, 27'h00000170, 32'h00000400,
  1'd1,  5'd7, 27'h000000b6, 5'd2, 27'h00000342, 5'd11, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d3, 5'd4, 27'h000003de, 5'd21, 27'h000003d5, 32'h00000400,
  1'd1,  5'd7, 27'h00000082, 5'd13, 27'h000003f0, 5'd6, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000095, 5'd15, 27'h000000d3, 5'd16, 27'h00000247, 32'h00000400,
  1'd1,  5'd8, 27'h00000385, 5'd12, 27'h00000380, 5'd27, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000142, 5'd22, 27'h00000280, 5'd6, 27'h000001fb, 32'h00000400,
  1'd1,  5'd6, 27'h00000066, 5'd23, 27'h00000156, 5'd17, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001b2, 5'd21, 27'h00000350, 5'd30, 27'h00000228, 32'h00000400,
  1'd1,  5'd16, 27'h000001f6, 5'd5, 27'h0000001a, 5'd1, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000037f, 5'd0, 27'h00000339, 5'd13, 27'h00000156, 32'h00000400,
  1'd1,  5'd18, 27'h00000234, 5'd2, 27'h000003b3, 5'd23, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000291, 5'd13, 27'h000001da, 5'd6, 27'h0000020c, 32'h00000400,
  1'd1,  5'd19, 27'h0000004d, 5'd14, 27'h0000018b, 5'd19, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c1, 5'd13, 27'h0000021a, 5'd30, 27'h00000208, 32'h00000400,
  1'd1,  5'd15, 27'h00000387, 5'd25, 27'h000002ad, 5'd7, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a5, 5'd25, 27'h000000e8, 5'd19, 27'h000003c8, 32'h00000400,
  1'd1,  5'd15, 27'h0000039b, 5'd23, 27'h000000bc, 5'd28, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000245, 5'd1, 27'h0000025b, 5'd8, 27'h000001a2, 32'h00000400,
  1'd1,  5'd26, 27'h000000cb, 5'd0, 27'h0000019f, 5'd16, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000364, 5'd4, 27'h000003fe, 5'd27, 27'h000003a5, 32'h00000400,
  1'd1,  5'd29, 27'h000003ae, 5'd14, 27'h000001c3, 5'd8, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000168, 5'd12, 27'h0000009d, 5'd16, 27'h00000345, 32'h00000400,
  1'd1,  5'd30, 27'h000000dd, 5'd13, 27'h00000160, 5'd30, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000023f, 5'd22, 27'h00000140, 5'd6, 27'h000000e2, 32'h00000400,
  1'd1,  5'd29, 27'h000002ac, 5'd25, 27'h00000111, 5'd19, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f6, 5'd22, 27'h000002af, 5'd27, 27'h00000273, 32'h00000400,
  1'd1,  5'd9, 27'h000000bd, 5'd8, 27'h0000015a, 5'd2, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000347, 5'd9, 27'h00000323, 5'd12, 27'h00000167, 32'h00000400,
  1'd1,  5'd9, 27'h000002df, 5'd7, 27'h000003a8, 5'd21, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000336, 5'd18, 27'h00000018, 5'd3, 27'h00000327, 32'h00000400,
  1'd1,  5'd8, 27'h00000270, 5'd18, 27'h0000025c, 5'd11, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000012f, 5'd17, 27'h00000213, 5'd20, 27'h000002e5, 32'h00000400,
  1'd1,  5'd6, 27'h000002fe, 5'd30, 27'h00000315, 5'd2, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000223, 5'd27, 27'h0000034e, 5'd13, 27'h00000381, 32'h00000400,
  1'd1,  5'd9, 27'h00000400, 5'd30, 27'h000000d2, 5'd21, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000e0, 5'd10, 27'h000000c8, 5'd3, 27'h0000024e, 32'h00000400,
  1'd1,  5'd16, 27'h00000369, 5'd6, 27'h00000294, 5'd12, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000125, 5'd9, 27'h0000000b, 5'd22, 27'h0000025f, 32'h00000400,
  1'd1,  5'd16, 27'h00000372, 5'd17, 27'h000001c2, 5'd2, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000215, 5'd15, 27'h000002a8, 5'd10, 27'h00000329, 32'h00000400,
  1'd1,  5'd19, 27'h000001db, 5'd20, 27'h0000003f, 5'd23, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000393, 5'd28, 27'h00000017, 5'd2, 27'h00000328, 32'h00000400,
  1'd1,  5'd18, 27'h000003d7, 5'd26, 27'h000003c9, 5'd10, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000025a, 5'd26, 27'h00000207, 5'd22, 27'h0000021d, 32'h00000400,
  1'd1,  5'd28, 27'h00000004, 5'd9, 27'h00000325, 5'd2, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001eb, 5'd8, 27'h0000034a, 5'd11, 27'h00000085, 32'h00000400,
  1'd1,  5'd26, 27'h000003c8, 5'd5, 27'h00000354, 5'd21, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000296, 5'd18, 27'h000002a3, 5'd4, 27'h00000234, 32'h00000400,
  1'd1,  5'd26, 27'h00000304, 5'd16, 27'h00000196, 5'd14, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003d3, 5'd20, 27'h0000000c, 5'd22, 27'h000003dc, 32'h00000400,
  1'd1,  5'd30, 27'h00000343, 5'd30, 27'h000001e6, 5'd4, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000361, 5'd30, 27'h0000037f, 5'd12, 27'h000002cc, 32'h00000400,
  1'd1,  5'd30, 27'h00000090, 5'd30, 27'h0000038d, 5'd25, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000306, 5'd9, 27'h0000020a, 5'd10, 27'h000000c8, 32'h00000400,
  1'd1,  5'd8, 27'h000003e8, 5'd8, 27'h0000035d, 5'd18, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e8, 5'd7, 27'h000000ec, 5'd26, 27'h0000019f, 32'h00000400,
  1'd1,  5'd8, 27'h0000001f, 5'd16, 27'h0000033d, 5'd8, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000e0, 5'd15, 27'h00000357, 5'd20, 27'h00000236, 32'h00000400,
  1'd1,  5'd8, 27'h000003bd, 5'd18, 27'h000001f4, 5'd28, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003e0, 5'd27, 27'h00000200, 5'd5, 27'h000002ad, 32'h00000400,
  1'd1,  5'd6, 27'h0000021f, 5'd26, 27'h00000001, 5'd16, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000091, 5'd28, 27'h00000021, 5'd28, 27'h00000166, 32'h00000400,
  1'd1,  5'd17, 27'h00000354, 5'd8, 27'h00000323, 5'd9, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000003c, 5'd8, 27'h000000e6, 5'd16, 27'h0000024d, 32'h00000400,
  1'd1,  5'd16, 27'h000003c1, 5'd7, 27'h0000016c, 5'd27, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000136, 5'd18, 27'h00000244, 5'd5, 27'h0000022b, 32'h00000400,
  1'd1,  5'd18, 27'h000000c2, 5'd16, 27'h00000209, 5'd17, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001c3, 5'd16, 27'h000001f2, 5'd26, 27'h00000104, 32'h00000400,
  1'd1,  5'd17, 27'h000000f7, 5'd30, 27'h0000002f, 5'd5, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000255, 5'd29, 27'h000001c8, 5'd20, 27'h00000291, 32'h00000400,
  1'd1,  5'd17, 27'h000003ef, 5'd29, 27'h00000306, 5'd27, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000034, 5'd9, 27'h00000296, 5'd6, 27'h000001a7, 32'h00000400,
  1'd1,  5'd30, 27'h0000018c, 5'd7, 27'h0000004c, 5'd16, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001c9, 5'd5, 27'h000000c2, 5'd30, 27'h00000361, 32'h00000400,
  1'd1,  5'd29, 27'h000001f2, 5'd17, 27'h0000000b, 5'd7, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003db, 5'd19, 27'h000000df, 5'd20, 27'h0000005b, 32'h00000400,
  1'd1,  5'd27, 27'h0000024f, 5'd20, 27'h000000ca, 5'd28, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000004, 5'd30, 27'h000000ce, 5'd7, 27'h000001c4, 32'h00000400,
  1'd1,  5'd28, 27'h0000005e, 5'd26, 27'h000000e6, 5'd19, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000046, 5'd30, 27'h000003ac, 5'd26, 27'h000003fc, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000058, 5'd4, 27'h0000003f, 5'd4, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000182, 5'd1, 27'h00000340, 5'd14, 27'h000001fc, 32'h00000400,
  1'd1,  5'd0, 27'h00000191, 5'd0, 27'h000000cb, 5'd21, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b1, 5'd14, 27'h000003cf, 5'd0, 27'h00000214, 32'h00000400,
  1'd1,  5'd1, 27'h0000030c, 5'd14, 27'h000002c1, 5'd12, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000339, 5'd10, 27'h00000300, 5'd23, 27'h0000002c, 32'h00000400,
  1'd1,  5'd2, 27'h000000ea, 5'd25, 27'h00000093, 5'd2, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003da, 5'd23, 27'h000000f5, 5'd13, 27'h0000038c, 32'h00000400,
  1'd1,  5'd3, 27'h00000150, 5'd22, 27'h00000344, 5'd22, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000297, 5'd1, 27'h00000351, 5'd4, 27'h000002c9, 32'h00000400,
  1'd1,  5'd15, 27'h00000155, 5'd2, 27'h0000010b, 5'd10, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000015b, 5'd5, 27'h00000063, 5'd21, 27'h00000010, 32'h00000400,
  1'd1,  5'd12, 27'h000002ce, 5'd10, 27'h000001ed, 5'd1, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000330, 5'd11, 27'h0000013c, 5'd13, 27'h00000130, 32'h00000400,
  1'd1,  5'd14, 27'h0000029c, 5'd12, 27'h00000231, 5'd25, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002fc, 5'd22, 27'h000002ac, 5'd4, 27'h000001dd, 32'h00000400,
  1'd1,  5'd10, 27'h000002ba, 5'd22, 27'h00000208, 5'd14, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ce, 5'd23, 27'h000000a8, 5'd25, 27'h00000111, 32'h00000400,
  1'd1,  5'd21, 27'h0000015a, 5'd0, 27'h00000335, 5'd2, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000014, 5'd3, 27'h0000002a, 5'd12, 27'h000001c6, 32'h00000400,
  1'd1,  5'd23, 27'h000001c8, 5'd4, 27'h000001d4, 5'd22, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000e5, 5'd10, 27'h0000038d, 5'd1, 27'h000000f5, 32'h00000400,
  1'd1,  5'd25, 27'h00000276, 5'd10, 27'h0000038a, 5'd13, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000149, 5'd13, 27'h00000085, 5'd22, 27'h000000f8, 32'h00000400,
  1'd1,  5'd23, 27'h000003d2, 5'd24, 27'h00000308, 5'd3, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b2, 5'd24, 27'h000003ae, 5'd13, 27'h00000332, 32'h00000400,
  1'd1,  5'd23, 27'h000001e9, 5'd22, 27'h00000037, 5'd21, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000386, 5'd2, 27'h00000275, 5'd7, 27'h00000352, 32'h00000400,
  1'd1,  5'd1, 27'h0000011f, 5'd1, 27'h000001af, 5'd16, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000d3, 5'd3, 27'h000003ac, 5'd27, 27'h00000043, 32'h00000400,
  1'd1,  5'd3, 27'h00000095, 5'd15, 27'h0000012d, 5'd8, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000126, 5'd12, 27'h000000b7, 5'd15, 27'h000002ca, 32'h00000400,
  1'd1,  5'd3, 27'h00000290, 5'd11, 27'h00000167, 5'd26, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000201, 5'd24, 27'h0000022c, 5'd6, 27'h000000e8, 32'h00000400,
  1'd1,  5'd3, 27'h00000332, 5'd21, 27'h000003a2, 5'd18, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000314, 5'd22, 27'h000001a9, 5'd26, 27'h000001cf, 32'h00000400,
  1'd1,  5'd14, 27'h000000d8, 5'd0, 27'h00000175, 5'd8, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003c7, 5'd0, 27'h000001c9, 5'd19, 27'h000003fd, 32'h00000400,
  1'd1,  5'd13, 27'h000000a8, 5'd3, 27'h0000027a, 5'd27, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000037b, 5'd13, 27'h00000221, 5'd9, 27'h00000172, 32'h00000400,
  1'd1,  5'd13, 27'h00000366, 5'd11, 27'h000003bc, 5'd15, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001fc, 5'd14, 27'h00000130, 5'd27, 27'h000000e6, 32'h00000400,
  1'd1,  5'd13, 27'h0000001e, 5'd25, 27'h000001bd, 5'd7, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000339, 5'd22, 27'h00000385, 5'd15, 27'h00000339, 32'h00000400,
  1'd1,  5'd12, 27'h0000022d, 5'd21, 27'h00000349, 5'd29, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000108, 5'd0, 27'h0000028f, 5'd9, 27'h0000012a, 32'h00000400,
  1'd1,  5'd22, 27'h00000101, 5'd0, 27'h0000014c, 5'd15, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000034d, 5'd1, 27'h00000379, 5'd27, 27'h000003de, 32'h00000400,
  1'd1,  5'd25, 27'h00000060, 5'd11, 27'h00000110, 5'd6, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000105, 5'd13, 27'h00000032, 5'd18, 27'h0000027c, 32'h00000400,
  1'd1,  5'd22, 27'h000000cb, 5'd11, 27'h000002a9, 5'd27, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000115, 5'd21, 27'h000000ae, 5'd9, 27'h000000a7, 32'h00000400,
  1'd1,  5'd21, 27'h0000034b, 5'd23, 27'h000000c5, 5'd20, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000bd, 5'd22, 27'h000001c5, 5'd29, 27'h00000290, 32'h00000400,
  1'd1,  5'd3, 27'h000002ad, 5'd10, 27'h00000024, 5'd4, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003ae, 5'd9, 27'h000001b1, 5'd14, 27'h00000060, 32'h00000400,
  1'd1,  5'd0, 27'h000003a3, 5'd7, 27'h00000244, 5'd24, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001cc, 5'd16, 27'h000002b6, 5'd4, 27'h0000034e, 32'h00000400,
  1'd1,  5'd0, 27'h00000192, 5'd17, 27'h00000001, 5'd14, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000004a, 5'd16, 27'h000002c1, 5'd21, 27'h0000036c, 32'h00000400,
  1'd1,  5'd4, 27'h000002b0, 5'd26, 27'h000000b0, 5'd3, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036d, 5'd27, 27'h000000d1, 5'd11, 27'h00000147, 32'h00000400,
  1'd1,  5'd0, 27'h00000020, 5'd27, 27'h000002be, 5'd24, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021c, 5'd7, 27'h000003f4, 5'd4, 27'h0000035f, 32'h00000400,
  1'd1,  5'd10, 27'h000001db, 5'd9, 27'h00000260, 5'd12, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003b6, 5'd10, 27'h0000010a, 5'd24, 27'h000000a9, 32'h00000400,
  1'd1,  5'd13, 27'h0000015d, 5'd16, 27'h000001f7, 5'd0, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000339, 5'd15, 27'h000002e8, 5'd11, 27'h00000320, 32'h00000400,
  1'd1,  5'd11, 27'h0000013b, 5'd16, 27'h0000037b, 5'd25, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003ba, 5'd26, 27'h000003fa, 5'd2, 27'h00000169, 32'h00000400,
  1'd1,  5'd12, 27'h000000b2, 5'd30, 27'h000001c9, 5'd15, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003dd, 5'd26, 27'h00000343, 5'd23, 27'h000003df, 32'h00000400,
  1'd1,  5'd25, 27'h00000034, 5'd6, 27'h00000118, 5'd3, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000358, 5'd7, 27'h0000037e, 5'd11, 27'h000003e5, 32'h00000400,
  1'd1,  5'd21, 27'h00000382, 5'd7, 27'h0000029f, 5'd20, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000034f, 5'd19, 27'h000002a1, 5'd2, 27'h000003bf, 32'h00000400,
  1'd1,  5'd22, 27'h000002a7, 5'd17, 27'h0000034b, 5'd10, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000055, 5'd19, 27'h000003e3, 5'd23, 27'h00000107, 32'h00000400,
  1'd1,  5'd20, 27'h000002ab, 5'd28, 27'h000001e1, 5'd2, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001ea, 5'd27, 27'h00000135, 5'd14, 27'h0000027f, 32'h00000400,
  1'd1,  5'd22, 27'h00000397, 5'd28, 27'h00000096, 5'd22, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000114, 5'd8, 27'h00000073, 5'd6, 27'h000000ed, 32'h00000400,
  1'd1,  5'd0, 27'h00000104, 5'd9, 27'h0000028c, 5'd18, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000006c, 5'd9, 27'h000002a9, 5'd26, 27'h00000396, 32'h00000400,
  1'd1,  5'd0, 27'h00000136, 5'd16, 27'h00000168, 5'd6, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000159, 5'd20, 27'h0000018b, 5'd19, 27'h00000044, 32'h00000400,
  1'd1,  5'd3, 27'h000001d8, 5'd17, 27'h0000030e, 5'd28, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f8, 5'd26, 27'h000000fe, 5'd9, 27'h00000033, 32'h00000400,
  1'd1,  5'd4, 27'h000002ac, 5'd27, 27'h000001ec, 5'd18, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000043, 5'd28, 27'h00000173, 5'd28, 27'h0000003d, 32'h00000400,
  1'd1,  5'd11, 27'h0000014d, 5'd10, 27'h00000112, 5'd7, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f7, 5'd7, 27'h000003e1, 5'd16, 27'h0000030c, 32'h00000400,
  1'd1,  5'd13, 27'h000000f5, 5'd5, 27'h0000028e, 5'd30, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000174, 5'd16, 27'h000002fa, 5'd6, 27'h000000cd, 32'h00000400,
  1'd1,  5'd15, 27'h0000017d, 5'd18, 27'h0000017d, 5'd16, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002b4, 5'd20, 27'h00000210, 5'd29, 27'h00000264, 32'h00000400,
  1'd1,  5'd11, 27'h0000022b, 5'd28, 27'h0000005c, 5'd7, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002e5, 5'd30, 27'h000003f9, 5'd16, 27'h000001ba, 32'h00000400,
  1'd1,  5'd15, 27'h000001f4, 5'd26, 27'h00000002, 5'd30, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000041, 5'd9, 27'h000001ac, 5'd7, 27'h000002b8, 32'h00000400,
  1'd1,  5'd24, 27'h000001a2, 5'd6, 27'h00000191, 5'd20, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000e8, 5'd9, 27'h0000015c, 5'd27, 27'h00000229, 32'h00000400,
  1'd1,  5'd23, 27'h00000121, 5'd19, 27'h0000026a, 5'd6, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000018a, 5'd17, 27'h00000067, 5'd18, 27'h000002f1, 32'h00000400,
  1'd1,  5'd23, 27'h00000090, 5'd17, 27'h000000ad, 5'd28, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035b, 5'd28, 27'h0000003e, 5'd8, 27'h000000e7, 32'h00000400,
  1'd1,  5'd24, 27'h000001b8, 5'd29, 27'h0000019f, 5'd19, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000bf, 5'd27, 27'h00000352, 5'd29, 27'h000002f9, 32'h00000400,
  1'd1,  5'd5, 27'h0000039d, 5'd4, 27'h0000031d, 5'd7, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003f9, 5'd3, 27'h000002ff, 5'd17, 27'h000001a5, 32'h00000400,
  1'd1,  5'd9, 27'h00000346, 5'd0, 27'h0000006b, 5'd30, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000265, 5'd12, 27'h000002b4, 5'd0, 27'h0000018b, 32'h00000400,
  1'd1,  5'd8, 27'h000003ec, 5'd10, 27'h000002f9, 5'd12, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000396, 5'd13, 27'h000003b1, 5'd23, 27'h00000143, 32'h00000400,
  1'd1,  5'd8, 27'h000001d5, 5'd20, 27'h000003fa, 5'd1, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000cf, 5'd25, 27'h000001ef, 5'd10, 27'h000002f2, 32'h00000400,
  1'd1,  5'd7, 27'h000001fc, 5'd21, 27'h00000022, 5'd25, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000028c, 5'd4, 27'h0000009d, 5'd6, 27'h000003f8, 32'h00000400,
  1'd1,  5'd16, 27'h00000381, 5'd0, 27'h00000115, 5'd20, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000075, 5'd5, 27'h00000038, 5'd29, 27'h00000337, 32'h00000400,
  1'd1,  5'd17, 27'h0000013e, 5'd13, 27'h00000027, 5'd0, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000028d, 5'd11, 27'h0000025e, 5'd15, 27'h00000152, 32'h00000400,
  1'd1,  5'd18, 27'h00000070, 5'd12, 27'h0000031e, 5'd21, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e0, 5'd24, 27'h000000cf, 5'd0, 27'h00000212, 32'h00000400,
  1'd1,  5'd18, 27'h000003a7, 5'd23, 27'h000000b2, 5'd10, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000eb, 5'd24, 27'h0000022d, 5'd22, 27'h000003e1, 32'h00000400,
  1'd1,  5'd28, 27'h00000369, 5'd4, 27'h0000031f, 5'd1, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003b1, 5'd3, 27'h000001e6, 5'd14, 27'h000001d2, 32'h00000400,
  1'd1,  5'd30, 27'h000001db, 5'd5, 27'h00000053, 5'd25, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000026a, 5'd10, 27'h000002ec, 5'd2, 27'h00000073, 32'h00000400,
  1'd1,  5'd30, 27'h0000003e, 5'd10, 27'h000003db, 5'd12, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a4, 5'd10, 27'h00000326, 5'd25, 27'h000001b4, 32'h00000400,
  1'd1,  5'd30, 27'h000003af, 5'd22, 27'h0000007c, 5'd1, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ad, 5'd22, 27'h00000214, 5'd11, 27'h00000006, 32'h00000400,
  1'd1,  5'd26, 27'h00000287, 5'd25, 27'h00000172, 5'd24, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000334, 5'd1, 27'h0000011c, 5'd4, 27'h000002dc, 32'h00000400,
  1'd1,  5'd9, 27'h000003e3, 5'd0, 27'h00000336, 5'd13, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018f, 5'd1, 27'h000003a6, 5'd25, 27'h00000114, 32'h00000400,
  1'd1,  5'd8, 27'h000003fb, 5'd14, 27'h000001b2, 5'd8, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000206, 5'd14, 27'h00000386, 5'd17, 27'h0000008b, 32'h00000400,
  1'd1,  5'd7, 27'h00000366, 5'd12, 27'h000000e3, 5'd26, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a1, 5'd21, 27'h0000022c, 5'd7, 27'h0000017a, 32'h00000400,
  1'd1,  5'd9, 27'h000001e5, 5'd21, 27'h0000000b, 5'd19, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000307, 5'd24, 27'h000002c2, 5'd26, 27'h00000226, 32'h00000400,
  1'd1,  5'd17, 27'h00000176, 5'd0, 27'h00000235, 5'd4, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000035e, 5'd3, 27'h0000024b, 5'd14, 27'h00000330, 32'h00000400,
  1'd1,  5'd17, 27'h00000358, 5'd1, 27'h000003b0, 5'd24, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d1, 5'd14, 27'h000003bf, 5'd7, 27'h000003ea, 32'h00000400,
  1'd1,  5'd15, 27'h00000207, 5'd14, 27'h000002bd, 5'd20, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000026c, 5'd11, 27'h00000376, 5'd29, 27'h00000260, 32'h00000400,
  1'd1,  5'd18, 27'h00000354, 5'd21, 27'h0000021f, 5'd7, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000104, 5'd22, 27'h000003f4, 5'd19, 27'h000003e6, 32'h00000400,
  1'd1,  5'd17, 27'h000003b2, 5'd23, 27'h0000019a, 5'd25, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c4, 5'd3, 27'h00000219, 5'd9, 27'h000001eb, 32'h00000400,
  1'd1,  5'd30, 27'h00000227, 5'd4, 27'h0000011f, 5'd19, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b9, 5'd2, 27'h0000032d, 5'd30, 27'h0000024c, 32'h00000400,
  1'd1,  5'd28, 27'h000000a6, 5'd14, 27'h000001e3, 5'd10, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000052, 5'd11, 27'h0000000a, 5'd18, 27'h0000035c, 32'h00000400,
  1'd1,  5'd26, 27'h0000006c, 5'd12, 27'h000000d0, 5'd30, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000158, 5'd22, 27'h000002ae, 5'd6, 27'h0000024b, 32'h00000400,
  1'd1,  5'd26, 27'h00000302, 5'd21, 27'h000002e5, 5'd18, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000003d, 5'd23, 27'h00000395, 5'd25, 27'h000003d2, 32'h00000400,
  1'd1,  5'd6, 27'h000001cb, 5'd5, 27'h00000267, 5'd2, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003b3, 5'd5, 27'h00000397, 5'd11, 27'h000002fa, 32'h00000400,
  1'd1,  5'd5, 27'h000001d5, 5'd8, 27'h00000049, 5'd25, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000015, 5'd19, 27'h000000ca, 5'd4, 27'h00000217, 32'h00000400,
  1'd1,  5'd7, 27'h00000357, 5'd17, 27'h000002dd, 5'd12, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c8, 5'd20, 27'h0000014b, 5'd21, 27'h0000007e, 32'h00000400,
  1'd1,  5'd9, 27'h00000083, 5'd29, 27'h000001a6, 5'd3, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b7, 5'd28, 27'h000002ac, 5'd15, 27'h0000017d, 32'h00000400,
  1'd1,  5'd7, 27'h000001fc, 5'd26, 27'h000003f5, 5'd22, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000366, 5'd5, 27'h00000282, 5'd2, 27'h000002d1, 32'h00000400,
  1'd1,  5'd17, 27'h000001a9, 5'd6, 27'h000002c2, 5'd10, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000fb, 5'd5, 27'h000003d9, 5'd22, 27'h00000300, 32'h00000400,
  1'd1,  5'd18, 27'h000003aa, 5'd16, 27'h000001c9, 5'd4, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000271, 5'd19, 27'h0000009f, 5'd12, 27'h00000260, 32'h00000400,
  1'd1,  5'd16, 27'h000002bc, 5'd19, 27'h00000287, 5'd21, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000038, 5'd28, 27'h000003f0, 5'd2, 27'h0000036e, 32'h00000400,
  1'd1,  5'd16, 27'h0000037c, 5'd26, 27'h000000a0, 5'd15, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f5, 5'd28, 27'h00000003, 5'd23, 27'h0000012b, 32'h00000400,
  1'd1,  5'd26, 27'h000003d9, 5'd9, 27'h00000069, 5'd4, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000036d, 5'd6, 27'h00000111, 5'd14, 27'h00000090, 32'h00000400,
  1'd1,  5'd27, 27'h00000108, 5'd6, 27'h0000009c, 5'd25, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b6, 5'd17, 27'h000001c9, 5'd2, 27'h00000188, 32'h00000400,
  1'd1,  5'd26, 27'h0000019c, 5'd15, 27'h00000230, 5'd14, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000301, 5'd20, 27'h00000152, 5'd24, 27'h000000dc, 32'h00000400,
  1'd1,  5'd28, 27'h0000007d, 5'd28, 27'h0000025d, 5'd0, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002b7, 5'd25, 27'h000003d0, 5'd11, 27'h0000018a, 32'h00000400,
  1'd1,  5'd29, 27'h000000bb, 5'd29, 27'h000003f5, 5'd23, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001af, 5'd8, 27'h00000217, 5'd6, 27'h0000009c, 32'h00000400,
  1'd1,  5'd9, 27'h000002c8, 5'd8, 27'h0000002d, 5'd19, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000031a, 5'd6, 27'h0000002b, 5'd30, 27'h00000305, 32'h00000400,
  1'd1,  5'd6, 27'h000001a6, 5'd16, 27'h00000220, 5'd6, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000234, 5'd18, 27'h0000005c, 5'd20, 27'h000000e5, 32'h00000400,
  1'd1,  5'd5, 27'h00000372, 5'd20, 27'h00000224, 5'd30, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000011b, 5'd29, 27'h00000077, 5'd7, 27'h000000a6, 32'h00000400,
  1'd1,  5'd8, 27'h000002b0, 5'd27, 27'h0000001c, 5'd19, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000400, 5'd30, 27'h0000011a, 5'd29, 27'h0000013e, 32'h00000400,
  1'd1,  5'd19, 27'h00000055, 5'd9, 27'h000000f8, 5'd5, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000298, 5'd8, 27'h00000223, 5'd18, 27'h00000032, 32'h00000400,
  1'd1,  5'd17, 27'h0000035c, 5'd7, 27'h000003a3, 5'd28, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e9, 5'd16, 27'h000001cb, 5'd6, 27'h0000011e, 32'h00000400,
  1'd1,  5'd16, 27'h0000018b, 5'd15, 27'h0000026e, 5'd15, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000011a, 5'd18, 27'h000000fa, 5'd29, 27'h00000114, 32'h00000400,
  1'd1,  5'd17, 27'h00000171, 5'd27, 27'h00000344, 5'd5, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ce, 5'd28, 27'h00000169, 5'd16, 27'h0000020e, 32'h00000400,
  1'd1,  5'd20, 27'h000000d3, 5'd28, 27'h000000c1, 5'd30, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000029a, 5'd8, 27'h000001e9, 5'd8, 27'h00000274, 32'h00000400,
  1'd1,  5'd30, 27'h00000379, 5'd7, 27'h00000081, 5'd16, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000397, 5'd6, 27'h000002fc, 5'd30, 27'h00000125, 32'h00000400,
  1'd1,  5'd26, 27'h00000382, 5'd15, 27'h00000236, 5'd9, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000023, 5'd19, 27'h0000034d, 5'd16, 27'h000002a4, 32'h00000400,
  1'd1,  5'd29, 27'h00000004, 5'd19, 27'h00000042, 5'd29, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000006a, 5'd27, 27'h00000173, 5'd10, 27'h00000107, 32'h00000400,
  1'd1,  5'd29, 27'h000001b2, 5'd30, 27'h0000010b, 5'd16, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a1, 5'd26, 27'h00000205, 5'd25, 27'h00000372, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000004f, 5'd2, 27'h000000aa, 5'd1, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ca, 5'd2, 27'h000001bb, 5'd11, 27'h00000382, 32'h00000400,
  1'd1,  5'd1, 27'h00000210, 5'd0, 27'h00000067, 5'd25, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c4, 5'd13, 27'h000002ce, 5'd0, 27'h0000009f, 32'h00000400,
  1'd1,  5'd4, 27'h000003c6, 5'd11, 27'h000000bd, 5'd15, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f7, 5'd13, 27'h0000022b, 5'd25, 27'h00000247, 32'h00000400,
  1'd1,  5'd1, 27'h000003cb, 5'd24, 27'h000001e4, 5'd2, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000019d, 5'd23, 27'h0000035f, 5'd10, 27'h0000034f, 32'h00000400,
  1'd1,  5'd2, 27'h00000225, 5'd21, 27'h00000224, 5'd25, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a9, 5'd2, 27'h00000077, 5'd4, 27'h0000002a, 32'h00000400,
  1'd1,  5'd13, 27'h0000031e, 5'd0, 27'h00000198, 5'd11, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000102, 5'd5, 27'h00000099, 5'd21, 27'h0000038a, 32'h00000400,
  1'd1,  5'd13, 27'h00000221, 5'd14, 27'h00000383, 5'd3, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000134, 5'd13, 27'h000001d8, 5'd10, 27'h000003fc, 32'h00000400,
  1'd1,  5'd13, 27'h0000007b, 5'd12, 27'h000001ea, 5'd23, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029d, 5'd25, 27'h000000c5, 5'd3, 27'h00000260, 32'h00000400,
  1'd1,  5'd13, 27'h00000155, 5'd20, 27'h00000303, 5'd15, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000022b, 5'd21, 27'h00000293, 5'd21, 27'h000002fc, 32'h00000400,
  1'd1,  5'd20, 27'h000002cb, 5'd0, 27'h00000336, 5'd3, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000214, 5'd5, 27'h00000046, 5'd11, 27'h00000031, 32'h00000400,
  1'd1,  5'd20, 27'h000002c0, 5'd0, 27'h00000318, 5'd25, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019e, 5'd13, 27'h0000031d, 5'd2, 27'h000003c1, 32'h00000400,
  1'd1,  5'd23, 27'h00000205, 5'd11, 27'h0000002c, 5'd10, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000199, 5'd10, 27'h00000368, 5'd21, 27'h00000095, 32'h00000400,
  1'd1,  5'd25, 27'h00000044, 5'd23, 27'h00000398, 5'd2, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001cc, 5'd21, 27'h000003db, 5'd14, 27'h0000005b, 32'h00000400,
  1'd1,  5'd24, 27'h00000053, 5'd24, 27'h000003be, 5'd22, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000272, 5'd3, 27'h000003e0, 5'd9, 27'h00000255, 32'h00000400,
  1'd1,  5'd1, 27'h000001c3, 5'd0, 27'h00000206, 5'd18, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000311, 5'd2, 27'h000000f9, 5'd27, 27'h00000395, 32'h00000400,
  1'd1,  5'd2, 27'h000003d0, 5'd12, 27'h00000180, 5'd5, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000b1, 5'd15, 27'h000001cf, 5'd18, 27'h000000be, 32'h00000400,
  1'd1,  5'd4, 27'h00000043, 5'd12, 27'h000000d2, 5'd30, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000b0, 5'd25, 27'h000000c6, 5'd7, 27'h00000311, 32'h00000400,
  1'd1,  5'd2, 27'h0000025b, 5'd21, 27'h00000041, 5'd16, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000060, 5'd22, 27'h000001b3, 5'd29, 27'h000001d8, 32'h00000400,
  1'd1,  5'd13, 27'h00000216, 5'd1, 27'h0000026e, 5'd5, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000015e, 5'd0, 27'h00000014, 5'd16, 27'h000002a6, 32'h00000400,
  1'd1,  5'd10, 27'h00000198, 5'd4, 27'h000002b1, 5'd26, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000df, 5'd12, 27'h000000ce, 5'd6, 27'h0000001e, 32'h00000400,
  1'd1,  5'd15, 27'h00000153, 5'd11, 27'h000003be, 5'd16, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000038c, 5'd14, 27'h00000338, 5'd26, 27'h00000148, 32'h00000400,
  1'd1,  5'd12, 27'h000003c2, 5'd20, 27'h000002bb, 5'd5, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000141, 5'd21, 27'h000000c9, 5'd20, 27'h00000080, 32'h00000400,
  1'd1,  5'd10, 27'h00000220, 5'd23, 27'h00000060, 5'd27, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ee, 5'd3, 27'h0000008c, 5'd10, 27'h000000a6, 32'h00000400,
  1'd1,  5'd25, 27'h00000057, 5'd3, 27'h0000011c, 5'd17, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000017c, 5'd0, 27'h00000078, 5'd28, 27'h00000268, 32'h00000400,
  1'd1,  5'd21, 27'h0000037c, 5'd15, 27'h000000f0, 5'd7, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b4, 5'd13, 27'h000001ca, 5'd18, 27'h000002af, 32'h00000400,
  1'd1,  5'd22, 27'h00000132, 5'd11, 27'h00000251, 5'd28, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a1, 5'd22, 27'h000000db, 5'd5, 27'h00000138, 32'h00000400,
  1'd1,  5'd22, 27'h000003ec, 5'd23, 27'h00000174, 5'd16, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002a2, 5'd24, 27'h00000355, 5'd29, 27'h0000036e, 32'h00000400,
  1'd1,  5'd2, 27'h000000ed, 5'd6, 27'h00000185, 5'd1, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001c1, 5'd8, 27'h0000002a, 5'd10, 27'h0000039f, 32'h00000400,
  1'd1,  5'd1, 27'h0000026e, 5'd6, 27'h00000021, 5'd23, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000331, 5'd19, 27'h000001e8, 5'd3, 27'h0000022e, 32'h00000400,
  1'd1,  5'd0, 27'h000003cb, 5'd17, 27'h0000007a, 5'd13, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000288, 5'd20, 27'h000001b7, 5'd25, 27'h000000c7, 32'h00000400,
  1'd1,  5'd1, 27'h000002e4, 5'd27, 27'h00000372, 5'd3, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000038d, 5'd30, 27'h000002be, 5'd14, 27'h00000318, 32'h00000400,
  1'd1,  5'd3, 27'h0000008b, 5'd30, 27'h000000f6, 5'd22, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029c, 5'd9, 27'h00000381, 5'd5, 27'h0000001e, 32'h00000400,
  1'd1,  5'd14, 27'h00000393, 5'd10, 27'h00000131, 5'd10, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000120, 5'd8, 27'h00000082, 5'd25, 27'h0000030c, 32'h00000400,
  1'd1,  5'd12, 27'h000003a5, 5'd16, 27'h0000006f, 5'd3, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003db, 5'd16, 27'h00000056, 5'd11, 27'h00000117, 32'h00000400,
  1'd1,  5'd11, 27'h000000a7, 5'd20, 27'h0000017b, 5'd25, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000146, 5'd30, 27'h0000027e, 5'd2, 27'h0000026e, 32'h00000400,
  1'd1,  5'd10, 27'h00000267, 5'd26, 27'h000003ac, 5'd10, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000333, 5'd26, 27'h0000008e, 5'd25, 27'h0000008e, 32'h00000400,
  1'd1,  5'd22, 27'h00000037, 5'd8, 27'h0000035f, 5'd2, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000176, 5'd6, 27'h00000198, 5'd12, 27'h00000124, 32'h00000400,
  1'd1,  5'd24, 27'h000002e9, 5'd7, 27'h000003f2, 5'd25, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000288, 5'd20, 27'h0000027c, 5'd3, 27'h00000160, 32'h00000400,
  1'd1,  5'd22, 27'h00000016, 5'd20, 27'h00000073, 5'd10, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001bb, 5'd19, 27'h00000228, 5'd25, 27'h00000039, 32'h00000400,
  1'd1,  5'd24, 27'h00000242, 5'd30, 27'h000002b8, 5'd3, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000039b, 5'd26, 27'h0000023e, 5'd15, 27'h0000008f, 32'h00000400,
  1'd1,  5'd21, 27'h00000073, 5'd27, 27'h0000021d, 5'd25, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000037f, 5'd5, 27'h00000200, 5'd7, 27'h00000111, 32'h00000400,
  1'd1,  5'd3, 27'h000003dc, 5'd9, 27'h00000072, 5'd18, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000398, 5'd9, 27'h000003fd, 5'd29, 27'h0000014c, 32'h00000400,
  1'd1,  5'd4, 27'h00000048, 5'd20, 27'h00000025, 5'd8, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014b, 5'd17, 27'h00000098, 5'd16, 27'h0000003c, 32'h00000400,
  1'd1,  5'd0, 27'h00000051, 5'd19, 27'h000003a7, 5'd30, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001e0, 5'd30, 27'h0000005c, 5'd6, 27'h00000316, 32'h00000400,
  1'd1,  5'd1, 27'h000002c6, 5'd27, 27'h00000269, 5'd16, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000120, 5'd29, 27'h0000011b, 5'd30, 27'h0000024d, 32'h00000400,
  1'd1,  5'd10, 27'h000003c7, 5'd8, 27'h00000003, 5'd6, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000033b, 5'd9, 27'h00000149, 5'd19, 27'h0000026c, 32'h00000400,
  1'd1,  5'd10, 27'h0000037a, 5'd6, 27'h00000106, 5'd30, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000028f, 5'd17, 27'h000002df, 5'd10, 27'h0000008c, 32'h00000400,
  1'd1,  5'd13, 27'h00000252, 5'd17, 27'h000002d5, 5'd17, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000244, 5'd20, 27'h000001cd, 5'd28, 27'h000000b4, 32'h00000400,
  1'd1,  5'd15, 27'h00000154, 5'd30, 27'h00000377, 5'd10, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000014c, 5'd25, 27'h000003f7, 5'd18, 27'h00000097, 32'h00000400,
  1'd1,  5'd10, 27'h000003be, 5'd26, 27'h00000127, 5'd27, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001fd, 5'd7, 27'h000002e3, 5'd9, 27'h000000a4, 32'h00000400,
  1'd1,  5'd25, 27'h00000216, 5'd6, 27'h00000049, 5'd19, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000020e, 5'd8, 27'h00000271, 5'd26, 27'h000002ae, 32'h00000400,
  1'd1,  5'd23, 27'h000000d9, 5'd19, 27'h0000025d, 5'd6, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000069, 5'd16, 27'h0000015c, 5'd18, 27'h0000008f, 32'h00000400,
  1'd1,  5'd24, 27'h000002b3, 5'd19, 27'h00000303, 5'd27, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000037b, 5'd28, 27'h00000134, 5'd5, 27'h000000c1, 32'h00000400,
  1'd1,  5'd22, 27'h00000302, 5'd28, 27'h000000c4, 5'd20, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003a8, 5'd30, 27'h000003ed, 5'd26, 27'h0000031f, 32'h00000400,
  1'd1,  5'd5, 27'h00000179, 5'd4, 27'h000001c8, 5'd7, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000105, 5'd2, 27'h00000037, 5'd17, 27'h00000297, 32'h00000400,
  1'd1,  5'd6, 27'h00000170, 5'd2, 27'h000002cf, 5'd29, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000231, 5'd10, 27'h000003e4, 5'd2, 27'h0000025e, 32'h00000400,
  1'd1,  5'd7, 27'h0000019b, 5'd12, 27'h00000093, 5'd13, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e7, 5'd15, 27'h0000017b, 5'd21, 27'h00000326, 32'h00000400,
  1'd1,  5'd6, 27'h00000276, 5'd22, 27'h000001a7, 5'd2, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000067, 5'd25, 27'h000001cd, 5'd11, 27'h00000387, 32'h00000400,
  1'd1,  5'd5, 27'h000002d0, 5'd22, 27'h000003cf, 5'd25, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000325, 5'd1, 27'h000000b8, 5'd9, 27'h000000e4, 32'h00000400,
  1'd1,  5'd16, 27'h00000015, 5'd3, 27'h0000022c, 5'd16, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d6, 5'd0, 27'h000000f8, 5'd26, 27'h000002f8, 32'h00000400,
  1'd1,  5'd16, 27'h00000304, 5'd13, 27'h0000023f, 5'd5, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000e5, 5'd15, 27'h000000f6, 5'd14, 27'h00000162, 32'h00000400,
  1'd1,  5'd19, 27'h0000006a, 5'd10, 27'h00000188, 5'd23, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000118, 5'd23, 27'h00000358, 5'd1, 27'h00000298, 32'h00000400,
  1'd1,  5'd18, 27'h0000038a, 5'd25, 27'h0000013c, 5'd10, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000003e, 5'd21, 27'h000000ab, 5'd22, 27'h0000013b, 32'h00000400,
  1'd1,  5'd29, 27'h00000227, 5'd4, 27'h000002ef, 5'd0, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000019d, 5'd3, 27'h00000226, 5'd11, 27'h00000194, 32'h00000400,
  1'd1,  5'd26, 27'h00000117, 5'd0, 27'h0000030e, 5'd24, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c1, 5'd13, 27'h000001fb, 5'd2, 27'h0000036a, 32'h00000400,
  1'd1,  5'd30, 27'h0000010d, 5'd13, 27'h00000108, 5'd14, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000014c, 5'd14, 27'h00000153, 5'd20, 27'h000002c0, 32'h00000400,
  1'd1,  5'd29, 27'h000000a3, 5'd25, 27'h000000ad, 5'd4, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000071, 5'd22, 27'h00000371, 5'd13, 27'h00000082, 32'h00000400,
  1'd1,  5'd28, 27'h000001cf, 5'd25, 27'h00000021, 5'd22, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000022f, 5'd2, 27'h000001e5, 5'd4, 27'h0000037d, 32'h00000400,
  1'd1,  5'd8, 27'h000001e5, 5'd3, 27'h000002eb, 5'd13, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000020d, 5'd4, 27'h00000090, 5'd24, 27'h0000032d, 32'h00000400,
  1'd1,  5'd6, 27'h000001f8, 5'd14, 27'h00000031, 5'd6, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003c4, 5'd15, 27'h00000073, 5'd18, 27'h0000008f, 32'h00000400,
  1'd1,  5'd5, 27'h000003d0, 5'd14, 27'h00000150, 5'd26, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001aa, 5'd22, 27'h000000c2, 5'd10, 27'h0000002c, 32'h00000400,
  1'd1,  5'd6, 27'h0000020e, 5'd22, 27'h00000284, 5'd19, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000325, 5'd24, 27'h00000099, 5'd28, 27'h00000355, 32'h00000400,
  1'd1,  5'd18, 27'h000002ad, 5'd4, 27'h00000077, 5'd4, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d0, 5'd4, 27'h000001c0, 5'd13, 27'h00000044, 32'h00000400,
  1'd1,  5'd17, 27'h000000bd, 5'd1, 27'h000001e4, 5'd22, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000139, 5'd14, 27'h000002f0, 5'd6, 27'h000001c9, 32'h00000400,
  1'd1,  5'd15, 27'h0000030e, 5'd11, 27'h00000107, 5'd16, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000028a, 5'd10, 27'h00000189, 5'd26, 27'h00000133, 32'h00000400,
  1'd1,  5'd19, 27'h0000030a, 5'd23, 27'h000001d1, 5'd9, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a8, 5'd21, 27'h00000189, 5'd16, 27'h000000c7, 32'h00000400,
  1'd1,  5'd19, 27'h0000022e, 5'd25, 27'h000000c4, 5'd30, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000229, 5'd2, 27'h00000373, 5'd7, 27'h0000025d, 32'h00000400,
  1'd1,  5'd29, 27'h00000268, 5'd3, 27'h00000034, 5'd16, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000bd, 5'd3, 27'h00000145, 5'd28, 27'h0000029b, 32'h00000400,
  1'd1,  5'd29, 27'h000001df, 5'd14, 27'h0000023f, 5'd8, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d8, 5'd13, 27'h000003c5, 5'd19, 27'h0000012c, 32'h00000400,
  1'd1,  5'd26, 27'h00000197, 5'd13, 27'h00000385, 5'd27, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ed, 5'd21, 27'h000001c6, 5'd8, 27'h0000011e, 32'h00000400,
  1'd1,  5'd30, 27'h00000227, 5'd24, 27'h0000036a, 5'd20, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000011e, 5'd23, 27'h000003f1, 5'd28, 27'h0000039a, 32'h00000400,
  1'd1,  5'd5, 27'h00000259, 5'd9, 27'h000002a1, 5'd2, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000267, 5'd9, 27'h000002b6, 5'd13, 27'h000000ef, 32'h00000400,
  1'd1,  5'd5, 27'h000000cc, 5'd8, 27'h000001ce, 5'd25, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000002e, 5'd19, 27'h0000036c, 5'd2, 27'h00000224, 32'h00000400,
  1'd1,  5'd5, 27'h00000292, 5'd17, 27'h000001a7, 5'd14, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000380, 5'd15, 27'h0000033c, 5'd25, 27'h0000026b, 32'h00000400,
  1'd1,  5'd5, 27'h0000036c, 5'd26, 27'h0000033b, 5'd4, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000332, 5'd29, 27'h000002c4, 5'd13, 27'h00000073, 32'h00000400,
  1'd1,  5'd6, 27'h0000034f, 5'd28, 27'h00000195, 5'd23, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000006a, 5'd9, 27'h00000289, 5'd3, 27'h0000036c, 32'h00000400,
  1'd1,  5'd20, 27'h00000137, 5'd6, 27'h000001a2, 5'd13, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003f8, 5'd8, 27'h000001c2, 5'd20, 27'h0000035d, 32'h00000400,
  1'd1,  5'd19, 27'h0000030e, 5'd17, 27'h00000049, 5'd3, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000b3, 5'd19, 27'h00000102, 5'd13, 27'h00000195, 32'h00000400,
  1'd1,  5'd16, 27'h00000334, 5'd18, 27'h00000307, 5'd24, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000084, 5'd26, 27'h000000a7, 5'd3, 27'h00000304, 32'h00000400,
  1'd1,  5'd15, 27'h000003e4, 5'd27, 27'h00000049, 5'd11, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000003, 5'd28, 27'h000001f2, 5'd20, 27'h0000036e, 32'h00000400,
  1'd1,  5'd30, 27'h000001e7, 5'd7, 27'h000000ef, 5'd1, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c8, 5'd8, 27'h0000034d, 5'd14, 27'h0000020c, 32'h00000400,
  1'd1,  5'd27, 27'h0000032a, 5'd9, 27'h000002ae, 5'd23, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000065, 5'd15, 27'h0000021d, 5'd0, 27'h00000042, 32'h00000400,
  1'd1,  5'd29, 27'h0000036e, 5'd19, 27'h0000020f, 5'd10, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000001c, 5'd17, 27'h000002ab, 5'd21, 27'h00000242, 32'h00000400,
  1'd1,  5'd27, 27'h000001e4, 5'd29, 27'h00000116, 5'd3, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001bb, 5'd30, 27'h000002f8, 5'd12, 27'h000002f7, 32'h00000400,
  1'd1,  5'd26, 27'h000000eb, 5'd27, 27'h000000dd, 5'd21, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c7, 5'd9, 27'h00000305, 5'd6, 27'h000001e9, 32'h00000400,
  1'd1,  5'd8, 27'h0000028f, 5'd9, 27'h000000d2, 5'd19, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000346, 5'd5, 27'h0000035c, 5'd26, 27'h0000017d, 32'h00000400,
  1'd1,  5'd5, 27'h00000186, 5'd16, 27'h000003fe, 5'd6, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005b, 5'd17, 27'h00000344, 5'd19, 27'h000000b0, 32'h00000400,
  1'd1,  5'd6, 27'h00000037, 5'd19, 27'h00000227, 5'd29, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000131, 5'd29, 27'h000000c5, 5'd5, 27'h000003dc, 32'h00000400,
  1'd1,  5'd7, 27'h00000222, 5'd28, 27'h00000319, 5'd16, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000031c, 5'd26, 27'h00000216, 5'd28, 27'h00000382, 32'h00000400,
  1'd1,  5'd19, 27'h000002ac, 5'd9, 27'h000002dc, 5'd9, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000f3, 5'd7, 27'h000003ce, 5'd17, 27'h00000130, 32'h00000400,
  1'd1,  5'd17, 27'h0000012a, 5'd9, 27'h00000229, 5'd28, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000047, 5'd15, 27'h0000034e, 5'd6, 27'h000003c1, 32'h00000400,
  1'd1,  5'd16, 27'h00000063, 5'd20, 27'h00000195, 5'd17, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000390, 5'd18, 27'h00000130, 5'd29, 27'h000001b6, 32'h00000400,
  1'd1,  5'd19, 27'h000002da, 5'd30, 27'h00000063, 5'd6, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000294, 5'd28, 27'h000001b6, 5'd16, 27'h0000007b, 32'h00000400,
  1'd1,  5'd17, 27'h00000244, 5'd28, 27'h000003fe, 5'd29, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000017e, 5'd6, 27'h0000027a, 5'd7, 27'h00000134, 32'h00000400,
  1'd1,  5'd29, 27'h000002e5, 5'd7, 27'h000002fa, 5'd18, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000169, 5'd9, 27'h000000be, 5'd28, 27'h00000222, 32'h00000400,
  1'd1,  5'd26, 27'h00000187, 5'd17, 27'h000003a5, 5'd7, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000382, 5'd16, 27'h000000c0, 5'd19, 27'h000001dd, 32'h00000400,
  1'd1,  5'd27, 27'h00000104, 5'd19, 27'h000002f7, 5'd29, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f2, 5'd29, 27'h000002c3, 5'd5, 27'h000002c3, 32'h00000400,
  1'd1,  5'd27, 27'h0000024c, 5'd27, 27'h000002f7, 5'd19, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000219, 5'd28, 27'h00000197, 5'd27, 27'h0000031a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000154, 5'd0, 27'h00000336, 5'd2, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000fc, 5'd2, 27'h0000004c, 5'd11, 27'h0000006d, 32'h00000400,
  1'd1,  5'd1, 27'h000002fd, 5'd2, 27'h00000330, 5'd24, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005c, 5'd12, 27'h000002bc, 5'd3, 27'h000000c7, 32'h00000400,
  1'd1,  5'd2, 27'h00000138, 5'd11, 27'h000003ed, 5'd15, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000001c, 5'd11, 27'h00000072, 5'd24, 27'h000001bd, 32'h00000400,
  1'd1,  5'd3, 27'h000003d6, 5'd25, 27'h00000297, 5'd4, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000257, 5'd20, 27'h0000031c, 5'd14, 27'h00000262, 32'h00000400,
  1'd1,  5'd2, 27'h000000ac, 5'd23, 27'h00000225, 5'd24, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000023b, 5'd3, 27'h000003e0, 5'd3, 27'h00000045, 32'h00000400,
  1'd1,  5'd13, 27'h00000258, 5'd4, 27'h000001b2, 5'd13, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f1, 5'd3, 27'h000000a2, 5'd21, 27'h00000255, 32'h00000400,
  1'd1,  5'd10, 27'h000002a6, 5'd15, 27'h00000009, 5'd0, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038e, 5'd10, 27'h00000165, 5'd12, 27'h0000023e, 32'h00000400,
  1'd1,  5'd11, 27'h00000003, 5'd15, 27'h0000005e, 5'd22, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000370, 5'd24, 27'h000002f5, 5'd3, 27'h00000025, 32'h00000400,
  1'd1,  5'd15, 27'h00000077, 5'd24, 27'h000000a6, 5'd13, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000000b, 5'd23, 27'h0000011c, 5'd22, 27'h00000218, 32'h00000400,
  1'd1,  5'd25, 27'h000000c1, 5'd4, 27'h0000023d, 5'd3, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003bd, 5'd0, 27'h0000004e, 5'd12, 27'h00000164, 32'h00000400,
  1'd1,  5'd23, 27'h0000010f, 5'd3, 27'h00000329, 5'd24, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000203, 5'd10, 27'h000002d0, 5'd2, 27'h000001b6, 32'h00000400,
  1'd1,  5'd21, 27'h00000062, 5'd13, 27'h000001b3, 5'd15, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000023, 5'd13, 27'h0000016c, 5'd22, 27'h00000283, 32'h00000400,
  1'd1,  5'd23, 27'h00000024, 5'd22, 27'h000001f4, 5'd2, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a1, 5'd21, 27'h000003dc, 5'd12, 27'h00000210, 32'h00000400,
  1'd1,  5'd23, 27'h000002e0, 5'd21, 27'h00000355, 5'd25, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000195, 5'd0, 27'h0000028d, 5'd10, 27'h00000035, 32'h00000400,
  1'd1,  5'd0, 27'h00000227, 5'd0, 27'h000002f6, 5'd19, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000196, 5'd3, 27'h00000178, 5'd26, 27'h000003a3, 32'h00000400,
  1'd1,  5'd4, 27'h00000173, 5'd12, 27'h00000161, 5'd7, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000282, 5'd10, 27'h000001da, 5'd16, 27'h00000317, 32'h00000400,
  1'd1,  5'd1, 27'h000000e9, 5'd12, 27'h00000119, 5'd26, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000e2, 5'd25, 27'h00000105, 5'd6, 27'h000003cd, 32'h00000400,
  1'd1,  5'd2, 27'h000002b8, 5'd25, 27'h000001ac, 5'd15, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000330, 5'd21, 27'h000002fa, 5'd27, 27'h0000005e, 32'h00000400,
  1'd1,  5'd13, 27'h00000159, 5'd2, 27'h000000ee, 5'd7, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000122, 5'd0, 27'h00000004, 5'd15, 27'h0000038b, 32'h00000400,
  1'd1,  5'd14, 27'h00000136, 5'd2, 27'h000003d4, 5'd29, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000017b, 5'd15, 27'h000000c1, 5'd7, 27'h000002ef, 32'h00000400,
  1'd1,  5'd14, 27'h00000361, 5'd12, 27'h0000014a, 5'd20, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001a2, 5'd14, 27'h0000017d, 5'd30, 27'h0000006e, 32'h00000400,
  1'd1,  5'd14, 27'h0000023e, 5'd23, 27'h0000004b, 5'd6, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000167, 5'd22, 27'h00000196, 5'd16, 27'h000003aa, 32'h00000400,
  1'd1,  5'd13, 27'h0000020f, 5'd20, 27'h000002dc, 5'd28, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000255, 5'd3, 27'h000000c7, 5'd9, 27'h000003aa, 32'h00000400,
  1'd1,  5'd21, 27'h00000179, 5'd3, 27'h00000033, 5'd16, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000a1, 5'd0, 27'h000000f9, 5'd30, 27'h000001f9, 32'h00000400,
  1'd1,  5'd23, 27'h0000039a, 5'd12, 27'h00000001, 5'd10, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001fa, 5'd15, 27'h00000131, 5'd16, 27'h00000207, 32'h00000400,
  1'd1,  5'd24, 27'h00000189, 5'd14, 27'h00000070, 5'd28, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001e7, 5'd20, 27'h00000332, 5'd6, 27'h0000025e, 32'h00000400,
  1'd1,  5'd23, 27'h00000247, 5'd21, 27'h000000c9, 5'd16, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ed, 5'd23, 27'h00000187, 5'd27, 27'h00000072, 32'h00000400,
  1'd1,  5'd0, 27'h00000103, 5'd9, 27'h0000018a, 5'd1, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001fe, 5'd7, 27'h000001c4, 5'd14, 27'h000002c3, 32'h00000400,
  1'd1,  5'd3, 27'h0000018c, 5'd9, 27'h00000326, 5'd24, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000031b, 5'd20, 27'h00000146, 5'd4, 27'h0000037c, 32'h00000400,
  1'd1,  5'd3, 27'h0000029f, 5'd16, 27'h0000009a, 5'd12, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000a2, 5'd20, 27'h000000b3, 5'd21, 27'h000002a9, 32'h00000400,
  1'd1,  5'd0, 27'h0000039f, 5'd28, 27'h00000213, 5'd3, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000050, 5'd28, 27'h0000017e, 5'd11, 27'h00000386, 32'h00000400,
  1'd1,  5'd4, 27'h000002e6, 5'd30, 27'h000000ec, 5'd22, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000018e, 5'd9, 27'h000002d3, 5'd3, 27'h00000257, 32'h00000400,
  1'd1,  5'd10, 27'h00000159, 5'd5, 27'h000002ea, 5'd11, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000028c, 5'd5, 27'h00000258, 5'd21, 27'h00000294, 32'h00000400,
  1'd1,  5'd13, 27'h000002bd, 5'd20, 27'h000000bc, 5'd0, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000032b, 5'd18, 27'h0000023f, 5'd11, 27'h0000001d, 32'h00000400,
  1'd1,  5'd13, 27'h0000005c, 5'd16, 27'h000001d4, 5'd25, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000175, 5'd27, 27'h0000013d, 5'd4, 27'h00000281, 32'h00000400,
  1'd1,  5'd14, 27'h0000002f, 5'd28, 27'h000000c4, 5'd13, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003ab, 5'd30, 27'h0000038f, 5'd25, 27'h00000068, 32'h00000400,
  1'd1,  5'd22, 27'h0000015e, 5'd7, 27'h0000008f, 5'd0, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ee, 5'd10, 27'h0000012b, 5'd11, 27'h000002bd, 32'h00000400,
  1'd1,  5'd20, 27'h000002d7, 5'd7, 27'h00000348, 5'd20, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002be, 5'd19, 27'h0000016e, 5'd1, 27'h00000314, 32'h00000400,
  1'd1,  5'd21, 27'h00000357, 5'd20, 27'h00000046, 5'd12, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ab, 5'd16, 27'h000000e8, 5'd22, 27'h00000071, 32'h00000400,
  1'd1,  5'd25, 27'h0000021c, 5'd30, 27'h000000df, 5'd1, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000007a, 5'd29, 27'h00000248, 5'd14, 27'h0000007c, 32'h00000400,
  1'd1,  5'd25, 27'h00000298, 5'd26, 27'h000001d4, 5'd24, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000038c, 5'd10, 27'h00000018, 5'd9, 27'h0000018f, 32'h00000400,
  1'd1,  5'd0, 27'h000001eb, 5'd10, 27'h000000d5, 5'd15, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f8, 5'd5, 27'h000001ae, 5'd27, 27'h0000035e, 32'h00000400,
  1'd1,  5'd1, 27'h00000336, 5'd15, 27'h00000344, 5'd9, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000150, 5'd18, 27'h00000087, 5'd19, 27'h00000288, 32'h00000400,
  1'd1,  5'd2, 27'h00000187, 5'd16, 27'h0000019b, 5'd26, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000020c, 5'd27, 27'h0000025c, 5'd9, 27'h000002e9, 32'h00000400,
  1'd1,  5'd4, 27'h00000065, 5'd30, 27'h0000004b, 5'd15, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000032e, 5'd30, 27'h0000014d, 5'd28, 27'h000002cc, 32'h00000400,
  1'd1,  5'd14, 27'h000001c2, 5'd5, 27'h000000e1, 5'd8, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000d0, 5'd7, 27'h0000033a, 5'd19, 27'h00000233, 32'h00000400,
  1'd1,  5'd12, 27'h00000302, 5'd6, 27'h00000092, 5'd26, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a5, 5'd20, 27'h000001ad, 5'd9, 27'h000001af, 32'h00000400,
  1'd1,  5'd10, 27'h00000228, 5'd18, 27'h000003be, 5'd19, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000256, 5'd15, 27'h00000256, 5'd30, 27'h00000056, 32'h00000400,
  1'd1,  5'd12, 27'h0000005c, 5'd26, 27'h0000011f, 5'd9, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031b, 5'd29, 27'h0000015f, 5'd19, 27'h00000129, 32'h00000400,
  1'd1,  5'd13, 27'h000001b4, 5'd29, 27'h000001c3, 5'd29, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000012e, 5'd7, 27'h000002fb, 5'd9, 27'h00000138, 32'h00000400,
  1'd1,  5'd22, 27'h000000da, 5'd9, 27'h0000019b, 5'd18, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000000a, 5'd8, 27'h00000398, 5'd30, 27'h000003df, 32'h00000400,
  1'd1,  5'd21, 27'h0000030b, 5'd19, 27'h000000ef, 5'd9, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000359, 5'd17, 27'h000002dc, 5'd17, 27'h0000020a, 32'h00000400,
  1'd1,  5'd23, 27'h000001cf, 5'd16, 27'h000002de, 5'd27, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000064, 5'd27, 27'h0000035a, 5'd9, 27'h000000a1, 32'h00000400,
  1'd1,  5'd23, 27'h0000039f, 5'd29, 27'h000000c7, 5'd16, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000259, 5'd30, 27'h0000001c, 5'd28, 27'h00000059, 32'h00000400,
  1'd1,  5'd7, 27'h0000035b, 5'd5, 27'h00000038, 5'd7, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000077, 5'd0, 27'h00000015, 5'd20, 27'h00000089, 32'h00000400,
  1'd1,  5'd9, 27'h00000259, 5'd1, 27'h000002c3, 5'd28, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000036a, 5'd12, 27'h0000009b, 5'd4, 27'h0000012e, 32'h00000400,
  1'd1,  5'd5, 27'h000001f0, 5'd14, 27'h00000368, 5'd13, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000002, 5'd14, 27'h000001d5, 5'd25, 27'h00000142, 32'h00000400,
  1'd1,  5'd5, 27'h0000032e, 5'd25, 27'h0000024e, 5'd0, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000132, 5'd24, 27'h00000104, 5'd15, 27'h00000195, 32'h00000400,
  1'd1,  5'd5, 27'h000001eb, 5'd25, 27'h0000019d, 5'd24, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000206, 5'd4, 27'h0000016b, 5'd5, 27'h000000de, 32'h00000400,
  1'd1,  5'd15, 27'h00000268, 5'd3, 27'h00000179, 5'd15, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a5, 5'd4, 27'h00000089, 5'd29, 27'h0000016f, 32'h00000400,
  1'd1,  5'd15, 27'h0000030b, 5'd12, 27'h000002ea, 5'd1, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000139, 5'd11, 27'h0000039d, 5'd13, 27'h0000035e, 32'h00000400,
  1'd1,  5'd18, 27'h000001a4, 5'd13, 27'h00000144, 5'd21, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000230, 5'd23, 27'h00000278, 5'd2, 27'h000002da, 32'h00000400,
  1'd1,  5'd15, 27'h00000399, 5'd25, 27'h000002f3, 5'd13, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000019c, 5'd21, 27'h000003ca, 5'd22, 27'h00000315, 32'h00000400,
  1'd1,  5'd26, 27'h000001a7, 5'd2, 27'h000000e6, 5'd0, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c1, 5'd4, 27'h000001e4, 5'd12, 27'h000001f5, 32'h00000400,
  1'd1,  5'd26, 27'h000000e4, 5'd0, 27'h00000104, 5'd24, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000071, 5'd14, 27'h00000075, 5'd4, 27'h0000003a, 32'h00000400,
  1'd1,  5'd27, 27'h000001b2, 5'd10, 27'h000002b3, 5'd10, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000003a, 5'd10, 27'h00000355, 5'd22, 27'h000002f9, 32'h00000400,
  1'd1,  5'd29, 27'h000002cb, 5'd24, 27'h00000370, 5'd0, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002af, 5'd23, 27'h000000d5, 5'd15, 27'h0000002d, 32'h00000400,
  1'd1,  5'd26, 27'h00000358, 5'd22, 27'h0000012c, 5'd21, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000069, 5'd4, 27'h0000032b, 5'd3, 27'h0000024a, 32'h00000400,
  1'd1,  5'd9, 27'h000000be, 5'd2, 27'h000001b8, 5'd11, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000207, 5'd5, 27'h0000000d, 5'd22, 27'h000000bf, 32'h00000400,
  1'd1,  5'd6, 27'h000001a0, 5'd12, 27'h0000031d, 5'd5, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000074, 5'd13, 27'h000003c2, 5'd20, 27'h000001bc, 32'h00000400,
  1'd1,  5'd10, 27'h000000cb, 5'd11, 27'h000000c9, 5'd30, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000288, 5'd21, 27'h0000030b, 5'd6, 27'h00000159, 32'h00000400,
  1'd1,  5'd7, 27'h000001dc, 5'd23, 27'h000003fb, 5'd18, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000127, 5'd25, 27'h000000c6, 5'd29, 27'h0000022d, 32'h00000400,
  1'd1,  5'd20, 27'h00000268, 5'd4, 27'h000002c2, 5'd3, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d3, 5'd1, 27'h000001bc, 5'd12, 27'h000003df, 32'h00000400,
  1'd1,  5'd19, 27'h00000322, 5'd3, 27'h000000d0, 5'd24, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000025a, 5'd12, 27'h000001ba, 5'd10, 27'h0000002e, 32'h00000400,
  1'd1,  5'd17, 27'h00000077, 5'd15, 27'h000001e4, 5'd16, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000264, 5'd14, 27'h000001eb, 5'd26, 27'h0000004c, 32'h00000400,
  1'd1,  5'd16, 27'h00000297, 5'd23, 27'h00000307, 5'd6, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f1, 5'd25, 27'h0000014b, 5'd16, 27'h0000008e, 32'h00000400,
  1'd1,  5'd20, 27'h00000119, 5'd24, 27'h0000021e, 5'd27, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000203, 5'd0, 27'h0000000b, 5'd10, 27'h00000123, 32'h00000400,
  1'd1,  5'd28, 27'h000003ed, 5'd3, 27'h000001d2, 5'd15, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000286, 5'd2, 27'h00000004, 5'd27, 27'h00000103, 32'h00000400,
  1'd1,  5'd29, 27'h000002e4, 5'd14, 27'h000001af, 5'd10, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036d, 5'd13, 27'h00000115, 5'd18, 27'h00000344, 32'h00000400,
  1'd1,  5'd29, 27'h00000217, 5'd12, 27'h0000004f, 5'd27, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000032f, 5'd20, 27'h00000397, 5'd6, 27'h000001f4, 32'h00000400,
  1'd1,  5'd29, 27'h00000010, 5'd24, 27'h000003dc, 5'd15, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000028f, 5'd22, 27'h000003e2, 5'd30, 27'h000003b6, 32'h00000400,
  1'd1,  5'd7, 27'h000000c7, 5'd8, 27'h0000037a, 5'd1, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000135, 5'd6, 27'h000003cc, 5'd10, 27'h0000038f, 32'h00000400,
  1'd1,  5'd7, 27'h000002b9, 5'd8, 27'h000002aa, 5'd24, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000020c, 5'd16, 27'h00000163, 5'd4, 27'h000001eb, 32'h00000400,
  1'd1,  5'd10, 27'h00000085, 5'd15, 27'h000003f4, 5'd14, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000a1, 5'd15, 27'h000002b8, 5'd21, 27'h0000005f, 32'h00000400,
  1'd1,  5'd9, 27'h000003f7, 5'd30, 27'h00000365, 5'd3, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000175, 5'd27, 27'h00000072, 5'd10, 27'h000002be, 32'h00000400,
  1'd1,  5'd8, 27'h000001ee, 5'd30, 27'h000000db, 5'd25, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002cc, 5'd7, 27'h000001f0, 5'd2, 27'h00000326, 32'h00000400,
  1'd1,  5'd16, 27'h00000150, 5'd6, 27'h000003e1, 5'd14, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000339, 5'd8, 27'h0000028d, 5'd24, 27'h00000221, 32'h00000400,
  1'd1,  5'd18, 27'h00000357, 5'd20, 27'h0000019e, 5'd4, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001e6, 5'd19, 27'h000002d0, 5'd14, 27'h000000e3, 32'h00000400,
  1'd1,  5'd16, 27'h00000104, 5'd18, 27'h00000339, 5'd21, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001f6, 5'd28, 27'h00000205, 5'd1, 27'h000003d8, 32'h00000400,
  1'd1,  5'd17, 27'h00000318, 5'd27, 27'h000003c6, 5'd10, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000022b, 5'd26, 27'h000003b3, 5'd25, 27'h0000023b, 32'h00000400,
  1'd1,  5'd28, 27'h000000fb, 5'd5, 27'h00000367, 5'd0, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000007a, 5'd8, 27'h00000346, 5'd14, 27'h00000221, 32'h00000400,
  1'd1,  5'd28, 27'h000003f9, 5'd8, 27'h00000303, 5'd24, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001d6, 5'd19, 27'h0000017c, 5'd3, 27'h00000006, 32'h00000400,
  1'd1,  5'd29, 27'h00000190, 5'd20, 27'h00000178, 5'd13, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000193, 5'd16, 27'h000001e3, 5'd22, 27'h0000032d, 32'h00000400,
  1'd1,  5'd26, 27'h0000035a, 5'd27, 27'h000002da, 5'd2, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000365, 5'd28, 27'h000003e7, 5'd12, 27'h000001bb, 32'h00000400,
  1'd1,  5'd28, 27'h00000061, 5'd28, 27'h00000118, 5'd24, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f7, 5'd7, 27'h000002ee, 5'd9, 27'h000002e7, 32'h00000400,
  1'd1,  5'd7, 27'h0000009a, 5'd7, 27'h000003ac, 5'd15, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000046, 5'd6, 27'h0000011f, 5'd29, 27'h00000289, 32'h00000400,
  1'd1,  5'd7, 27'h00000373, 5'd17, 27'h000002f0, 5'd9, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000103, 5'd16, 27'h00000334, 5'd16, 27'h000001dc, 32'h00000400,
  1'd1,  5'd7, 27'h00000046, 5'd18, 27'h00000308, 5'd26, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000218, 5'd27, 27'h0000011d, 5'd7, 27'h0000017c, 32'h00000400,
  1'd1,  5'd5, 27'h000000db, 5'd26, 27'h0000034a, 5'd16, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001c0, 5'd27, 27'h00000005, 5'd26, 27'h000002e8, 32'h00000400,
  1'd1,  5'd16, 27'h00000367, 5'd8, 27'h0000015f, 5'd5, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000300, 5'd10, 27'h00000112, 5'd19, 27'h000001fa, 32'h00000400,
  1'd1,  5'd18, 27'h000000d6, 5'd5, 27'h00000200, 5'd28, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000400, 5'd17, 27'h000000dc, 5'd6, 27'h00000106, 32'h00000400,
  1'd1,  5'd17, 27'h00000273, 5'd15, 27'h0000031e, 5'd19, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000f3, 5'd18, 27'h00000266, 5'd27, 27'h000000dc, 32'h00000400,
  1'd1,  5'd20, 27'h00000093, 5'd26, 27'h000002a9, 5'd9, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a7, 5'd29, 27'h000002d1, 5'd20, 27'h00000154, 32'h00000400,
  1'd1,  5'd20, 27'h000000b1, 5'd29, 27'h000000bf, 5'd27, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000115, 5'd5, 27'h000000bd, 5'd9, 27'h000003c9, 32'h00000400,
  1'd1,  5'd27, 27'h0000003e, 5'd7, 27'h0000030a, 5'd19, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000031c, 5'd6, 27'h00000249, 5'd30, 27'h00000131, 32'h00000400,
  1'd1,  5'd29, 27'h0000038b, 5'd17, 27'h0000019d, 5'd7, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034f, 5'd18, 27'h00000115, 5'd17, 27'h00000207, 32'h00000400,
  1'd1,  5'd26, 27'h00000002, 5'd17, 27'h0000025e, 5'd28, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000299, 5'd28, 27'h000000ca, 5'd5, 27'h00000108, 32'h00000400,
  1'd1,  5'd27, 27'h00000374, 5'd30, 27'h000000e2, 5'd18, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002b0, 5'd27, 27'h00000015, 5'd27, 27'h000002d3, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h0000034b, 5'd4, 27'h000003b7, 5'd1, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000000, 5'd3, 27'h0000028b, 5'd11, 27'h000003a2, 32'h00000400,
  1'd1,  5'd3, 27'h00000198, 5'd1, 27'h000003cf, 5'd25, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f9, 5'd10, 27'h00000308, 5'd2, 27'h0000026a, 32'h00000400,
  1'd1,  5'd4, 27'h0000016b, 5'd14, 27'h00000212, 5'd12, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000277, 5'd14, 27'h0000039d, 5'd23, 27'h000003c9, 32'h00000400,
  1'd1,  5'd4, 27'h00000234, 5'd23, 27'h00000250, 5'd4, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001cf, 5'd23, 27'h00000235, 5'd10, 27'h0000028c, 32'h00000400,
  1'd1,  5'd3, 27'h000003b7, 5'd22, 27'h00000050, 5'd24, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000004d, 5'd4, 27'h00000045, 5'd0, 27'h00000062, 32'h00000400,
  1'd1,  5'd12, 27'h000003e4, 5'd1, 27'h000000f2, 5'd12, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002e3, 5'd4, 27'h000003f0, 5'd23, 27'h00000206, 32'h00000400,
  1'd1,  5'd13, 27'h000002fc, 5'd11, 27'h000000ab, 5'd2, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000036, 5'd10, 27'h0000028e, 5'd14, 27'h000002e5, 32'h00000400,
  1'd1,  5'd11, 27'h000000b0, 5'd13, 27'h00000336, 5'd20, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025d, 5'd23, 27'h0000035c, 5'd3, 27'h00000204, 32'h00000400,
  1'd1,  5'd12, 27'h00000303, 5'd23, 27'h0000020b, 5'd14, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000084, 5'd22, 27'h0000016d, 5'd21, 27'h00000106, 32'h00000400,
  1'd1,  5'd21, 27'h00000092, 5'd3, 27'h000000e6, 5'd1, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000066, 5'd0, 27'h00000023, 5'd11, 27'h0000016b, 32'h00000400,
  1'd1,  5'd22, 27'h000001be, 5'd2, 27'h00000232, 5'd22, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000f7, 5'd14, 27'h0000013b, 5'd1, 27'h000000fb, 32'h00000400,
  1'd1,  5'd22, 27'h00000396, 5'd13, 27'h00000218, 5'd10, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000af, 5'd11, 27'h000001b0, 5'd24, 27'h000001d0, 32'h00000400,
  1'd1,  5'd24, 27'h00000141, 5'd23, 27'h00000039, 5'd3, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002e5, 5'd23, 27'h00000053, 5'd14, 27'h0000017a, 32'h00000400,
  1'd1,  5'd24, 27'h00000371, 5'd24, 27'h00000320, 5'd25, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b6, 5'd4, 27'h0000016e, 5'd7, 27'h00000392, 32'h00000400,
  1'd1,  5'd3, 27'h000000fd, 5'd1, 27'h00000213, 5'd19, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000124, 5'd1, 27'h0000025e, 5'd26, 27'h0000030b, 32'h00000400,
  1'd1,  5'd0, 27'h000003c1, 5'd10, 27'h000003ec, 5'd9, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000041, 5'd12, 27'h0000024c, 5'd17, 27'h00000386, 32'h00000400,
  1'd1,  5'd1, 27'h00000207, 5'd13, 27'h0000003a, 5'd26, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000263, 5'd23, 27'h000000de, 5'd7, 27'h00000360, 32'h00000400,
  1'd1,  5'd0, 27'h0000019b, 5'd24, 27'h00000061, 5'd19, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000020f, 5'd20, 27'h00000399, 5'd26, 27'h000001a9, 32'h00000400,
  1'd1,  5'd12, 27'h0000005a, 5'd3, 27'h000001bf, 5'd7, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001de, 5'd1, 27'h00000254, 5'd16, 27'h0000019f, 32'h00000400,
  1'd1,  5'd11, 27'h00000083, 5'd0, 27'h00000336, 5'd29, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003a5, 5'd11, 27'h00000238, 5'd6, 27'h000003c8, 32'h00000400,
  1'd1,  5'd14, 27'h000002b2, 5'd14, 27'h00000125, 5'd18, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000360, 5'd10, 27'h000003c2, 5'd30, 27'h000002bd, 32'h00000400,
  1'd1,  5'd12, 27'h00000200, 5'd23, 27'h00000179, 5'd7, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000109, 5'd25, 27'h000000e4, 5'd16, 27'h0000031d, 32'h00000400,
  1'd1,  5'd10, 27'h000003ae, 5'd24, 27'h0000022c, 5'd29, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000006f, 5'd4, 27'h000003bf, 5'd5, 27'h000002cd, 32'h00000400,
  1'd1,  5'd23, 27'h000000db, 5'd4, 27'h0000008c, 5'd17, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002af, 5'd4, 27'h000002e8, 5'd27, 27'h00000352, 32'h00000400,
  1'd1,  5'd23, 27'h00000063, 5'd13, 27'h00000288, 5'd7, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000282, 5'd12, 27'h0000025a, 5'd16, 27'h00000139, 32'h00000400,
  1'd1,  5'd24, 27'h000001c3, 5'd15, 27'h00000078, 5'd29, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001d1, 5'd23, 27'h000003c8, 5'd7, 27'h000000a6, 32'h00000400,
  1'd1,  5'd22, 27'h0000028c, 5'd24, 27'h000003d4, 5'd15, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f9, 5'd21, 27'h000001c8, 5'd28, 27'h000003fe, 32'h00000400,
  1'd1,  5'd4, 27'h000002f2, 5'd8, 27'h00000029, 5'd1, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003e2, 5'd9, 27'h00000126, 5'd12, 27'h0000009e, 32'h00000400,
  1'd1,  5'd2, 27'h0000013b, 5'd8, 27'h0000015a, 5'd24, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000217, 5'd18, 27'h00000397, 5'd4, 27'h000003ed, 32'h00000400,
  1'd1,  5'd1, 27'h000001b3, 5'd17, 27'h000003e5, 5'd12, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000032d, 5'd16, 27'h0000001e, 5'd22, 27'h000000ba, 32'h00000400,
  1'd1,  5'd1, 27'h0000024f, 5'd26, 27'h000001cc, 5'd3, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003cc, 5'd25, 27'h0000036d, 5'd11, 27'h000000a0, 32'h00000400,
  1'd1,  5'd4, 27'h00000077, 5'd26, 27'h0000033c, 5'd20, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000070, 5'd5, 27'h0000038c, 5'd1, 27'h00000305, 32'h00000400,
  1'd1,  5'd10, 27'h0000018b, 5'd7, 27'h00000112, 5'd12, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a8, 5'd6, 27'h000002db, 5'd24, 27'h000001e5, 32'h00000400,
  1'd1,  5'd13, 27'h0000003d, 5'd16, 27'h00000002, 5'd3, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003c7, 5'd19, 27'h000000f7, 5'd10, 27'h0000017e, 32'h00000400,
  1'd1,  5'd13, 27'h00000101, 5'd16, 27'h00000089, 5'd21, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002dd, 5'd28, 27'h0000034b, 5'd0, 27'h0000019b, 32'h00000400,
  1'd1,  5'd10, 27'h000001bb, 5'd29, 27'h0000012d, 5'd14, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000018, 5'd30, 27'h0000025f, 5'd22, 27'h0000005f, 32'h00000400,
  1'd1,  5'd24, 27'h000001cf, 5'd5, 27'h000003d7, 5'd2, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000015d, 5'd5, 27'h00000234, 5'd12, 27'h00000171, 32'h00000400,
  1'd1,  5'd22, 27'h00000360, 5'd6, 27'h00000082, 5'd22, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000144, 5'd17, 27'h00000360, 5'd3, 27'h0000036a, 32'h00000400,
  1'd1,  5'd24, 27'h000003e9, 5'd17, 27'h0000016b, 5'd13, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000035, 5'd17, 27'h0000037a, 5'd21, 27'h00000207, 32'h00000400,
  1'd1,  5'd22, 27'h000003d8, 5'd26, 27'h000000fb, 5'd4, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000d3, 5'd26, 27'h000003a2, 5'd15, 27'h000000cd, 32'h00000400,
  1'd1,  5'd25, 27'h000002d1, 5'd29, 27'h000003c0, 5'd25, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d5, 5'd7, 27'h000002ae, 5'd6, 27'h000002b9, 32'h00000400,
  1'd1,  5'd2, 27'h000001f4, 5'd5, 27'h0000012c, 5'd17, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000022, 5'd7, 27'h00000333, 5'd28, 27'h00000306, 32'h00000400,
  1'd1,  5'd1, 27'h000002c5, 5'd19, 27'h00000231, 5'd9, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000175, 5'd16, 27'h000003fa, 5'd20, 27'h00000131, 32'h00000400,
  1'd1,  5'd1, 27'h0000038d, 5'd20, 27'h000000db, 5'd28, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000017f, 5'd28, 27'h000000e9, 5'd8, 27'h00000064, 32'h00000400,
  1'd1,  5'd3, 27'h00000294, 5'd27, 27'h000000c3, 5'd20, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ad, 5'd30, 27'h0000037e, 5'd30, 27'h0000025e, 32'h00000400,
  1'd1,  5'd11, 27'h000002c3, 5'd7, 27'h0000005c, 5'd6, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000013, 5'd7, 27'h000002a0, 5'd18, 27'h00000400, 32'h00000400,
  1'd1,  5'd12, 27'h000000ee, 5'd8, 27'h00000269, 5'd29, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000018a, 5'd20, 27'h00000260, 5'd5, 27'h000000ae, 32'h00000400,
  1'd1,  5'd11, 27'h000002df, 5'd19, 27'h000003e9, 5'd18, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000014, 5'd18, 27'h00000275, 5'd30, 27'h0000029b, 32'h00000400,
  1'd1,  5'd10, 27'h0000017a, 5'd26, 27'h000003ec, 5'd9, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001b1, 5'd29, 27'h000000b2, 5'd18, 27'h00000026, 32'h00000400,
  1'd1,  5'd15, 27'h00000088, 5'd25, 27'h000003ed, 5'd30, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034d, 5'd10, 27'h00000031, 5'd8, 27'h00000031, 32'h00000400,
  1'd1,  5'd23, 27'h000002aa, 5'd7, 27'h000001fa, 5'd19, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000232, 5'd8, 27'h000003d4, 5'd25, 27'h000003a7, 32'h00000400,
  1'd1,  5'd23, 27'h0000006a, 5'd18, 27'h0000010d, 5'd5, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000188, 5'd15, 27'h00000204, 5'd18, 27'h0000033a, 32'h00000400,
  1'd1,  5'd22, 27'h0000021b, 5'd15, 27'h000002bd, 5'd26, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000293, 5'd26, 27'h000003e9, 5'd6, 27'h000000b2, 32'h00000400,
  1'd1,  5'd22, 27'h00000038, 5'd29, 27'h00000267, 5'd16, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000272, 5'd27, 27'h0000035a, 5'd30, 27'h0000018e, 32'h00000400,
  1'd1,  5'd6, 27'h00000279, 5'd2, 27'h000003f0, 5'd7, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000035c, 5'd1, 27'h000002e9, 5'd17, 27'h000003b4, 32'h00000400,
  1'd1,  5'd5, 27'h00000337, 5'd2, 27'h000002cf, 5'd27, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000102, 5'd13, 27'h000002fe, 5'd1, 27'h000002ad, 32'h00000400,
  1'd1,  5'd6, 27'h00000246, 5'd11, 27'h0000005b, 5'd13, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000255, 5'd15, 27'h000001d6, 5'd22, 27'h000000b2, 32'h00000400,
  1'd1,  5'd7, 27'h0000020e, 5'd22, 27'h0000018a, 5'd1, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000190, 5'd22, 27'h000002b8, 5'd14, 27'h00000169, 32'h00000400,
  1'd1,  5'd6, 27'h0000023f, 5'd20, 27'h0000037b, 5'd25, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d8, 5'd3, 27'h0000000a, 5'd7, 27'h0000026f, 32'h00000400,
  1'd1,  5'd16, 27'h00000039, 5'd1, 27'h0000005f, 5'd17, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000009c, 5'd4, 27'h000001f2, 5'd28, 27'h000002e1, 32'h00000400,
  1'd1,  5'd17, 27'h0000022e, 5'd14, 27'h0000016e, 5'd2, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000108, 5'd11, 27'h00000180, 5'd15, 27'h00000192, 32'h00000400,
  1'd1,  5'd15, 27'h00000225, 5'd13, 27'h000001b4, 5'd25, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000176, 5'd21, 27'h000000a7, 5'd4, 27'h00000029, 32'h00000400,
  1'd1,  5'd15, 27'h0000032e, 5'd25, 27'h0000003f, 5'd14, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e5, 5'd25, 27'h000001c2, 5'd23, 27'h00000318, 32'h00000400,
  1'd1,  5'd29, 27'h00000254, 5'd0, 27'h000001ed, 5'd2, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000336, 5'd3, 27'h000001f0, 5'd13, 27'h00000315, 32'h00000400,
  1'd1,  5'd28, 27'h000002e6, 5'd0, 27'h000002d0, 5'd23, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c0, 5'd15, 27'h00000041, 5'd1, 27'h00000304, 32'h00000400,
  1'd1,  5'd29, 27'h000002a5, 5'd14, 27'h000003fd, 5'd14, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a6, 5'd12, 27'h00000018, 5'd24, 27'h0000008d, 32'h00000400,
  1'd1,  5'd27, 27'h0000033f, 5'd24, 27'h00000050, 5'd3, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000277, 5'd22, 27'h000001d1, 5'd15, 27'h00000178, 32'h00000400,
  1'd1,  5'd29, 27'h000000c8, 5'd22, 27'h0000039e, 5'd20, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000006a, 5'd1, 27'h000001b0, 5'd5, 27'h00000084, 32'h00000400,
  1'd1,  5'd6, 27'h0000034c, 5'd4, 27'h000003dc, 5'd13, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ac, 5'd0, 27'h000002cb, 5'd23, 27'h000003af, 32'h00000400,
  1'd1,  5'd9, 27'h00000051, 5'd14, 27'h000001a3, 5'd5, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002ef, 5'd10, 27'h00000166, 5'd19, 27'h000002da, 32'h00000400,
  1'd1,  5'd7, 27'h000000a6, 5'd15, 27'h000000b3, 5'd27, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000002c, 5'd21, 27'h0000030d, 5'd7, 27'h0000035c, 32'h00000400,
  1'd1,  5'd8, 27'h0000028e, 5'd23, 27'h000001d4, 5'd16, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002a7, 5'd24, 27'h0000003e, 5'd30, 27'h00000336, 32'h00000400,
  1'd1,  5'd17, 27'h000000d0, 5'd4, 27'h00000092, 5'd2, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000000, 5'd3, 27'h00000133, 5'd13, 27'h000001d5, 32'h00000400,
  1'd1,  5'd16, 27'h00000020, 5'd4, 27'h00000329, 5'd22, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f2, 5'd13, 27'h00000069, 5'd6, 27'h000003d0, 32'h00000400,
  1'd1,  5'd18, 27'h00000049, 5'd10, 27'h00000290, 5'd16, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000004f, 5'd11, 27'h00000372, 5'd28, 27'h0000022f, 32'h00000400,
  1'd1,  5'd19, 27'h0000021a, 5'd23, 27'h0000010c, 5'd8, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001c2, 5'd22, 27'h00000026, 5'd17, 27'h000002d1, 32'h00000400,
  1'd1,  5'd17, 27'h00000290, 5'd21, 27'h000001b1, 5'd27, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a9, 5'd0, 27'h00000179, 5'd6, 27'h00000248, 32'h00000400,
  1'd1,  5'd28, 27'h00000220, 5'd0, 27'h000001a8, 5'd17, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000043, 5'd4, 27'h00000364, 5'd30, 27'h00000142, 32'h00000400,
  1'd1,  5'd29, 27'h000003c9, 5'd12, 27'h000000c0, 5'd6, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000030, 5'd15, 27'h00000092, 5'd20, 27'h000000a4, 32'h00000400,
  1'd1,  5'd29, 27'h000003cd, 5'd14, 27'h000000f6, 5'd26, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000355, 5'd23, 27'h0000012c, 5'd9, 27'h0000037c, 32'h00000400,
  1'd1,  5'd27, 27'h00000249, 5'd21, 27'h000003d9, 5'd19, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000000e, 5'd22, 27'h0000010d, 5'd27, 27'h0000031e, 32'h00000400,
  1'd1,  5'd7, 27'h0000012f, 5'd9, 27'h000001f3, 5'd0, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001c1, 5'd7, 27'h00000397, 5'd14, 27'h00000287, 32'h00000400,
  1'd1,  5'd6, 27'h00000039, 5'd8, 27'h0000005f, 5'd23, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023b, 5'd18, 27'h000003f8, 5'd0, 27'h000000e5, 32'h00000400,
  1'd1,  5'd6, 27'h000000a2, 5'd16, 27'h000000e4, 5'd12, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012d, 5'd19, 27'h0000010b, 5'd22, 27'h00000099, 32'h00000400,
  1'd1,  5'd9, 27'h0000023e, 5'd28, 27'h00000109, 5'd0, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000a7, 5'd27, 27'h000003f0, 5'd11, 27'h00000228, 32'h00000400,
  1'd1,  5'd9, 27'h0000035b, 5'd27, 27'h000000ba, 5'd24, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000210, 5'd10, 27'h000000af, 5'd3, 27'h000000e6, 32'h00000400,
  1'd1,  5'd19, 27'h0000013d, 5'd9, 27'h00000155, 5'd14, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e8, 5'd7, 27'h000001e6, 5'd24, 27'h00000152, 32'h00000400,
  1'd1,  5'd19, 27'h00000090, 5'd18, 27'h000003b2, 5'd3, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000219, 5'd15, 27'h000002ec, 5'd13, 27'h00000284, 32'h00000400,
  1'd1,  5'd20, 27'h00000127, 5'd18, 27'h00000224, 5'd24, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000035, 5'd30, 27'h00000399, 5'd4, 27'h000000a4, 32'h00000400,
  1'd1,  5'd16, 27'h0000010f, 5'd27, 27'h000000f0, 5'd11, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000326, 5'd29, 27'h000001f2, 5'd24, 27'h00000087, 32'h00000400,
  1'd1,  5'd26, 27'h0000028e, 5'd5, 27'h000000b8, 5'd2, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a2, 5'd9, 27'h0000004d, 5'd12, 27'h00000084, 32'h00000400,
  1'd1,  5'd26, 27'h0000015c, 5'd9, 27'h000002ee, 5'd21, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000160, 5'd18, 27'h00000125, 5'd3, 27'h00000034, 32'h00000400,
  1'd1,  5'd25, 27'h00000396, 5'd16, 27'h000001cf, 5'd15, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000d2, 5'd17, 27'h00000256, 5'd24, 27'h00000085, 32'h00000400,
  1'd1,  5'd27, 27'h00000031, 5'd30, 27'h00000330, 5'd1, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000324, 5'd27, 27'h00000127, 5'd12, 27'h00000116, 32'h00000400,
  1'd1,  5'd26, 27'h000003fd, 5'd28, 27'h000003e4, 5'd25, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d0, 5'd9, 27'h00000103, 5'd8, 27'h000000f3, 32'h00000400,
  1'd1,  5'd9, 27'h00000273, 5'd7, 27'h00000197, 5'd17, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001f3, 5'd10, 27'h0000012c, 5'd26, 27'h0000037e, 32'h00000400,
  1'd1,  5'd10, 27'h00000135, 5'd18, 27'h000003f2, 5'd6, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000001c, 5'd15, 27'h000002ee, 5'd15, 27'h000002b5, 32'h00000400,
  1'd1,  5'd7, 27'h00000293, 5'd17, 27'h00000101, 5'd26, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003bb, 5'd30, 27'h000003ce, 5'd8, 27'h00000055, 32'h00000400,
  1'd1,  5'd6, 27'h000002ac, 5'd27, 27'h0000019c, 5'd19, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000152, 5'd27, 27'h00000004, 5'd28, 27'h000003d3, 32'h00000400,
  1'd1,  5'd18, 27'h00000108, 5'd10, 27'h00000146, 5'd6, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000008b, 5'd6, 27'h0000001c, 5'd17, 27'h000001d9, 32'h00000400,
  1'd1,  5'd16, 27'h00000154, 5'd7, 27'h00000292, 5'd29, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000027, 5'd18, 27'h000001f6, 5'd9, 27'h0000014b, 32'h00000400,
  1'd1,  5'd19, 27'h000003bb, 5'd16, 27'h00000118, 5'd18, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000294, 5'd15, 27'h000003e9, 5'd28, 27'h000001e7, 32'h00000400,
  1'd1,  5'd15, 27'h00000396, 5'd29, 27'h000003b2, 5'd7, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000210, 5'd29, 27'h0000024e, 5'd19, 27'h000003cf, 32'h00000400,
  1'd1,  5'd18, 27'h000003df, 5'd27, 27'h00000236, 5'd29, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ed, 5'd10, 27'h0000014e, 5'd8, 27'h00000056, 32'h00000400,
  1'd1,  5'd28, 27'h00000330, 5'd7, 27'h00000362, 5'd20, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000037e, 5'd8, 27'h000002df, 5'd27, 27'h0000026e, 32'h00000400,
  1'd1,  5'd29, 27'h00000299, 5'd20, 27'h00000009, 5'd8, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000383, 5'd19, 27'h0000023b, 5'd18, 27'h00000232, 32'h00000400,
  1'd1,  5'd28, 27'h000000b5, 5'd19, 27'h000002fa, 5'd29, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ae, 5'd29, 27'h00000374, 5'd6, 27'h000001b3, 32'h00000400,
  1'd1,  5'd29, 27'h00000023, 5'd28, 27'h000001ff, 5'd18, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000368, 5'd30, 27'h00000090, 5'd28, 27'h0000007c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h0000024a, 5'd3, 27'h000001c9, 5'd4, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ba, 5'd4, 27'h000003db, 5'd13, 27'h00000092, 32'h00000400,
  1'd1,  5'd1, 27'h000002a2, 5'd3, 27'h000001ee, 5'd23, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000022d, 5'd13, 27'h000000c6, 5'd0, 27'h000000be, 32'h00000400,
  1'd1,  5'd3, 27'h0000003f, 5'd11, 27'h00000209, 5'd12, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a4, 5'd14, 27'h00000111, 5'd20, 27'h00000374, 32'h00000400,
  1'd1,  5'd0, 27'h00000096, 5'd23, 27'h0000025f, 5'd2, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032a, 5'd25, 27'h00000281, 5'd13, 27'h00000250, 32'h00000400,
  1'd1,  5'd4, 27'h00000185, 5'd25, 27'h000001d4, 5'd22, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000034, 5'd0, 27'h00000253, 5'd0, 27'h0000038d, 32'h00000400,
  1'd1,  5'd11, 27'h0000011e, 5'd4, 27'h000001f4, 5'd10, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002d5, 5'd3, 27'h0000011d, 5'd25, 27'h000002e9, 32'h00000400,
  1'd1,  5'd15, 27'h00000055, 5'd10, 27'h00000361, 5'd3, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000355, 5'd14, 27'h00000337, 5'd11, 27'h00000141, 32'h00000400,
  1'd1,  5'd12, 27'h00000336, 5'd10, 27'h00000311, 5'd22, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000097, 5'd24, 27'h00000262, 5'd2, 27'h00000111, 32'h00000400,
  1'd1,  5'd10, 27'h00000390, 5'd24, 27'h00000049, 5'd15, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000179, 5'd22, 27'h00000109, 5'd20, 27'h000002b2, 32'h00000400,
  1'd1,  5'd25, 27'h000000dd, 5'd4, 27'h000003fc, 5'd2, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000034c, 5'd2, 27'h0000006a, 5'd12, 27'h000000c4, 32'h00000400,
  1'd1,  5'd21, 27'h000000d5, 5'd1, 27'h000001e3, 5'd21, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e7, 5'd14, 27'h000003e6, 5'd4, 27'h0000022d, 32'h00000400,
  1'd1,  5'd23, 27'h0000039e, 5'd11, 27'h00000198, 5'd13, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000363, 5'd11, 27'h00000267, 5'd22, 27'h0000015d, 32'h00000400,
  1'd1,  5'd23, 27'h0000016b, 5'd22, 27'h00000182, 5'd4, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000129, 5'd23, 27'h000003b4, 5'd10, 27'h0000034d, 32'h00000400,
  1'd1,  5'd22, 27'h000003ac, 5'd22, 27'h000000d8, 5'd24, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000080, 5'd1, 27'h00000088, 5'd5, 27'h0000025b, 32'h00000400,
  1'd1,  5'd4, 27'h00000216, 5'd4, 27'h000002f8, 5'd18, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002aa, 5'd0, 27'h000002a9, 5'd29, 27'h00000297, 32'h00000400,
  1'd1,  5'd1, 27'h000001aa, 5'd14, 27'h00000320, 5'd10, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000003f, 5'd14, 27'h000000c7, 5'd19, 27'h00000267, 32'h00000400,
  1'd1,  5'd0, 27'h000001a0, 5'd11, 27'h000003f5, 5'd30, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000bb, 5'd25, 27'h0000034d, 5'd5, 27'h00000271, 32'h00000400,
  1'd1,  5'd3, 27'h00000210, 5'd25, 27'h0000015a, 5'd18, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000340, 5'd21, 27'h00000211, 5'd27, 27'h00000196, 32'h00000400,
  1'd1,  5'd13, 27'h00000028, 5'd1, 27'h000003b2, 5'd8, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fe, 5'd4, 27'h0000021e, 5'd16, 27'h000001c7, 32'h00000400,
  1'd1,  5'd10, 27'h000002e2, 5'd5, 27'h0000005e, 5'd28, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000252, 5'd14, 27'h00000008, 5'd7, 27'h00000399, 32'h00000400,
  1'd1,  5'd12, 27'h000003e5, 5'd15, 27'h000001ad, 5'd17, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000012e, 5'd13, 27'h0000011a, 5'd28, 27'h000002ef, 32'h00000400,
  1'd1,  5'd13, 27'h000002bc, 5'd25, 27'h000000e7, 5'd6, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001bb, 5'd24, 27'h000002ff, 5'd16, 27'h000003e7, 32'h00000400,
  1'd1,  5'd14, 27'h0000013f, 5'd24, 27'h0000005b, 5'd28, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000147, 5'd2, 27'h000003aa, 5'd8, 27'h00000242, 32'h00000400,
  1'd1,  5'd22, 27'h0000011b, 5'd2, 27'h00000082, 5'd20, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003ff, 5'd4, 27'h00000117, 5'd27, 27'h000002a0, 32'h00000400,
  1'd1,  5'd20, 27'h00000321, 5'd13, 27'h0000004b, 5'd7, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000219, 5'd15, 27'h00000096, 5'd18, 27'h00000279, 32'h00000400,
  1'd1,  5'd25, 27'h000002b5, 5'd14, 27'h00000109, 5'd27, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d8, 5'd21, 27'h00000006, 5'd10, 27'h00000150, 32'h00000400,
  1'd1,  5'd23, 27'h000003d2, 5'd23, 27'h0000001e, 5'd17, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000004f, 5'd25, 27'h00000116, 5'd28, 27'h000000f4, 32'h00000400,
  1'd1,  5'd3, 27'h000002ad, 5'd5, 27'h00000241, 5'd1, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000121, 5'd6, 27'h00000050, 5'd12, 27'h000003ed, 32'h00000400,
  1'd1,  5'd0, 27'h000000cd, 5'd8, 27'h00000392, 5'd21, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000031b, 5'd15, 27'h0000029c, 5'd4, 27'h000000e8, 32'h00000400,
  1'd1,  5'd0, 27'h00000108, 5'd20, 27'h000000aa, 5'd15, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f0, 5'd19, 27'h000002fe, 5'd23, 27'h000003fb, 32'h00000400,
  1'd1,  5'd0, 27'h00000346, 5'd26, 27'h00000271, 5'd3, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000013f, 5'd28, 27'h000002b9, 5'd13, 27'h00000085, 32'h00000400,
  1'd1,  5'd3, 27'h0000021b, 5'd28, 27'h000000ae, 5'd21, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000085, 5'd7, 27'h0000030b, 5'd0, 27'h00000036, 32'h00000400,
  1'd1,  5'd15, 27'h000001be, 5'd7, 27'h00000270, 5'd12, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000323, 5'd6, 27'h00000222, 5'd23, 27'h000000d4, 32'h00000400,
  1'd1,  5'd12, 27'h000003a6, 5'd18, 27'h000001be, 5'd3, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000399, 5'd20, 27'h00000050, 5'd14, 27'h000000b1, 32'h00000400,
  1'd1,  5'd14, 27'h0000029b, 5'd20, 27'h000000ec, 5'd24, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000a6, 5'd30, 27'h0000029c, 5'd2, 27'h00000358, 32'h00000400,
  1'd1,  5'd10, 27'h000002b5, 5'd30, 27'h000003ff, 5'd14, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a6, 5'd27, 27'h000003a7, 5'd23, 27'h000002a5, 32'h00000400,
  1'd1,  5'd21, 27'h000002bd, 5'd8, 27'h0000015f, 5'd0, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000340, 5'd8, 27'h00000022, 5'd14, 27'h000000f4, 32'h00000400,
  1'd1,  5'd20, 27'h000002d6, 5'd7, 27'h00000212, 5'd23, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000038f, 5'd20, 27'h00000048, 5'd0, 27'h00000178, 32'h00000400,
  1'd1,  5'd22, 27'h0000018e, 5'd16, 27'h00000387, 5'd14, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000307, 5'd16, 27'h000003cb, 5'd23, 27'h00000367, 32'h00000400,
  1'd1,  5'd22, 27'h0000030a, 5'd28, 27'h00000075, 5'd0, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002c8, 5'd27, 27'h000002c6, 5'd13, 27'h00000214, 32'h00000400,
  1'd1,  5'd21, 27'h00000099, 5'd28, 27'h00000276, 5'd25, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d5, 5'd9, 27'h00000004, 5'd6, 27'h0000036c, 32'h00000400,
  1'd1,  5'd4, 27'h000001f9, 5'd8, 27'h0000016d, 5'd15, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000014, 5'd6, 27'h00000394, 5'd26, 27'h000003c3, 32'h00000400,
  1'd1,  5'd4, 27'h0000011d, 5'd17, 27'h0000035d, 5'd6, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000030f, 5'd18, 27'h0000030f, 5'd17, 27'h00000345, 32'h00000400,
  1'd1,  5'd4, 27'h0000004f, 5'd18, 27'h00000296, 5'd28, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000008a, 5'd29, 27'h00000123, 5'd7, 27'h0000012a, 32'h00000400,
  1'd1,  5'd3, 27'h00000081, 5'd26, 27'h0000025a, 5'd17, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018f, 5'd30, 27'h000000ba, 5'd29, 27'h00000370, 32'h00000400,
  1'd1,  5'd12, 27'h000000fa, 5'd9, 27'h000000b3, 5'd8, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000360, 5'd9, 27'h0000007f, 5'd17, 27'h000002ad, 32'h00000400,
  1'd1,  5'd10, 27'h00000293, 5'd8, 27'h00000048, 5'd29, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000192, 5'd18, 27'h00000320, 5'd7, 27'h00000222, 32'h00000400,
  1'd1,  5'd15, 27'h00000061, 5'd18, 27'h00000319, 5'd16, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000002d, 5'd19, 27'h0000003b, 5'd30, 27'h000000bc, 32'h00000400,
  1'd1,  5'd12, 27'h00000350, 5'd27, 27'h000001a1, 5'd8, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000074, 5'd30, 27'h000002ec, 5'd17, 27'h000000e9, 32'h00000400,
  1'd1,  5'd13, 27'h00000383, 5'd30, 27'h000001de, 5'd30, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000007b, 5'd7, 27'h0000007e, 5'd6, 27'h000003c6, 32'h00000400,
  1'd1,  5'd20, 27'h00000369, 5'd7, 27'h00000131, 5'd19, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000135, 5'd10, 27'h000000f5, 5'd27, 27'h000000e6, 32'h00000400,
  1'd1,  5'd23, 27'h00000278, 5'd18, 27'h00000043, 5'd7, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000025d, 5'd16, 27'h0000034e, 5'd20, 27'h00000114, 32'h00000400,
  1'd1,  5'd21, 27'h000001bc, 5'd17, 27'h00000076, 5'd28, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000026d, 5'd28, 27'h000002a0, 5'd5, 27'h0000035d, 32'h00000400,
  1'd1,  5'd22, 27'h0000000a, 5'd30, 27'h0000037b, 5'd16, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000377, 5'd29, 27'h00000136, 5'd27, 27'h000001fd, 32'h00000400,
  1'd1,  5'd8, 27'h00000164, 5'd2, 27'h0000012b, 5'd5, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000227, 5'd4, 27'h0000019a, 5'd18, 27'h000000f3, 32'h00000400,
  1'd1,  5'd5, 27'h000001f6, 5'd1, 27'h000003ab, 5'd26, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b3, 5'd11, 27'h0000033a, 5'd3, 27'h0000038e, 32'h00000400,
  1'd1,  5'd10, 27'h0000011d, 5'd15, 27'h0000010b, 5'd11, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003b8, 5'd10, 27'h00000348, 5'd22, 27'h0000002b, 32'h00000400,
  1'd1,  5'd8, 27'h0000012d, 5'd24, 27'h00000215, 5'd3, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f8, 5'd24, 27'h000000e8, 5'd11, 27'h00000178, 32'h00000400,
  1'd1,  5'd9, 27'h00000140, 5'd21, 27'h000003ee, 5'd25, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000007c, 5'd3, 27'h000001bf, 5'd7, 27'h00000061, 32'h00000400,
  1'd1,  5'd19, 27'h0000013c, 5'd3, 27'h000000ad, 5'd17, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000308, 5'd4, 27'h00000390, 5'd27, 27'h00000267, 32'h00000400,
  1'd1,  5'd19, 27'h00000220, 5'd10, 27'h00000203, 5'd2, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000019f, 5'd13, 27'h00000291, 5'd12, 27'h00000077, 32'h00000400,
  1'd1,  5'd18, 27'h000002fd, 5'd13, 27'h00000013, 5'd21, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d6, 5'd22, 27'h00000238, 5'd0, 27'h00000207, 32'h00000400,
  1'd1,  5'd19, 27'h0000000b, 5'd23, 27'h000001f6, 5'd11, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002e7, 5'd24, 27'h00000308, 5'd23, 27'h000002eb, 32'h00000400,
  1'd1,  5'd27, 27'h000000e2, 5'd4, 27'h000001ea, 5'd2, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000280, 5'd5, 27'h00000030, 5'd11, 27'h000000c0, 32'h00000400,
  1'd1,  5'd27, 27'h00000093, 5'd3, 27'h000002fc, 5'd24, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ca, 5'd12, 27'h000001fd, 5'd3, 27'h0000016c, 32'h00000400,
  1'd1,  5'd26, 27'h0000025a, 5'd12, 27'h00000377, 5'd10, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000023d, 5'd12, 27'h000001a0, 5'd21, 27'h000002c0, 32'h00000400,
  1'd1,  5'd28, 27'h00000254, 5'd24, 27'h000002b9, 5'd3, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000de, 5'd23, 27'h00000192, 5'd13, 27'h0000029b, 32'h00000400,
  1'd1,  5'd29, 27'h00000175, 5'd25, 27'h00000069, 5'd24, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000267, 5'd1, 27'h00000152, 5'd1, 27'h000002b5, 32'h00000400,
  1'd1,  5'd10, 27'h00000048, 5'd0, 27'h00000306, 5'd14, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000029c, 5'd4, 27'h000000e6, 5'd24, 27'h00000052, 32'h00000400,
  1'd1,  5'd8, 27'h00000375, 5'd11, 27'h0000005d, 5'd6, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000132, 5'd13, 27'h0000007f, 5'd19, 27'h0000027d, 32'h00000400,
  1'd1,  5'd7, 27'h0000029b, 5'd10, 27'h00000236, 5'd29, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000005f, 5'd20, 27'h000003e2, 5'd6, 27'h00000037, 32'h00000400,
  1'd1,  5'd6, 27'h0000031c, 5'd21, 27'h00000363, 5'd20, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000390, 5'd25, 27'h000001c7, 5'd29, 27'h000002d2, 32'h00000400,
  1'd1,  5'd19, 27'h0000021b, 5'd1, 27'h000003a2, 5'd2, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000029, 5'd4, 27'h000000b5, 5'd12, 27'h00000277, 32'h00000400,
  1'd1,  5'd15, 27'h000003e2, 5'd1, 27'h00000240, 5'd23, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000371, 5'd12, 27'h0000008e, 5'd8, 27'h00000174, 32'h00000400,
  1'd1,  5'd16, 27'h00000248, 5'd15, 27'h000001c8, 5'd18, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003dc, 5'd12, 27'h00000056, 5'd29, 27'h0000030b, 32'h00000400,
  1'd1,  5'd20, 27'h00000028, 5'd21, 27'h000001b0, 5'd6, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000296, 5'd24, 27'h00000191, 5'd16, 27'h00000096, 32'h00000400,
  1'd1,  5'd18, 27'h0000037e, 5'd25, 27'h0000014b, 5'd30, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000c1, 5'd2, 27'h000002d6, 5'd8, 27'h000002d4, 32'h00000400,
  1'd1,  5'd30, 27'h0000011a, 5'd4, 27'h0000004d, 5'd18, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000384, 5'd2, 27'h0000016a, 5'd28, 27'h0000001e, 32'h00000400,
  1'd1,  5'd26, 27'h000000bb, 5'd13, 27'h000003c2, 5'd8, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000035, 5'd11, 27'h00000002, 5'd19, 27'h0000016c, 32'h00000400,
  1'd1,  5'd30, 27'h000000cc, 5'd13, 27'h000001fc, 5'd26, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000132, 5'd23, 27'h00000299, 5'd9, 27'h000003fb, 32'h00000400,
  1'd1,  5'd26, 27'h000000df, 5'd23, 27'h000003f0, 5'd17, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c1, 5'd23, 27'h0000015c, 5'd29, 27'h0000023e, 32'h00000400,
  1'd1,  5'd5, 27'h000001e3, 5'd6, 27'h000000a4, 5'd2, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000236, 5'd9, 27'h0000007d, 5'd10, 27'h0000031e, 32'h00000400,
  1'd1,  5'd5, 27'h000003ec, 5'd8, 27'h00000291, 5'd20, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c0, 5'd19, 27'h0000034e, 5'd1, 27'h0000038e, 32'h00000400,
  1'd1,  5'd8, 27'h00000192, 5'd17, 27'h000000a5, 5'd12, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002bf, 5'd19, 27'h00000208, 5'd23, 27'h0000034d, 32'h00000400,
  1'd1,  5'd10, 27'h000000ea, 5'd27, 27'h00000091, 5'd2, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c0, 5'd27, 27'h000000fb, 5'd14, 27'h0000006b, 32'h00000400,
  1'd1,  5'd7, 27'h0000013e, 5'd28, 27'h00000257, 5'd25, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000235, 5'd6, 27'h00000379, 5'd3, 27'h0000001b, 32'h00000400,
  1'd1,  5'd16, 27'h0000021a, 5'd8, 27'h000002d8, 5'd11, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029b, 5'd5, 27'h00000133, 5'd20, 27'h000003cf, 32'h00000400,
  1'd1,  5'd18, 27'h0000021c, 5'd16, 27'h00000091, 5'd4, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000277, 5'd16, 27'h00000011, 5'd12, 27'h00000144, 32'h00000400,
  1'd1,  5'd19, 27'h000001ec, 5'd18, 27'h00000351, 5'd20, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f9, 5'd25, 27'h000003da, 5'd2, 27'h000001d0, 32'h00000400,
  1'd1,  5'd16, 27'h000003c8, 5'd29, 27'h00000374, 5'd13, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000285, 5'd29, 27'h0000017b, 5'd23, 27'h000001d1, 32'h00000400,
  1'd1,  5'd27, 27'h00000045, 5'd9, 27'h000003da, 5'd4, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000033e, 5'd6, 27'h00000332, 5'd14, 27'h0000020a, 32'h00000400,
  1'd1,  5'd28, 27'h00000061, 5'd6, 27'h000003e9, 5'd22, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001a9, 5'd19, 27'h0000027d, 5'd2, 27'h000003c5, 32'h00000400,
  1'd1,  5'd29, 27'h00000181, 5'd16, 27'h00000160, 5'd14, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000001a, 5'd18, 27'h0000018b, 5'd21, 27'h0000034c, 32'h00000400,
  1'd1,  5'd27, 27'h0000037e, 5'd30, 27'h000001d0, 5'd0, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000322, 5'd30, 27'h00000203, 5'd12, 27'h0000029d, 32'h00000400,
  1'd1,  5'd28, 27'h00000196, 5'd30, 27'h00000060, 5'd22, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000097, 5'd6, 27'h0000020e, 5'd7, 27'h000000e8, 32'h00000400,
  1'd1,  5'd5, 27'h000000e0, 5'd10, 27'h000000eb, 5'd20, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000082, 5'd8, 27'h00000269, 5'd30, 27'h000003f2, 32'h00000400,
  1'd1,  5'd5, 27'h000001c1, 5'd19, 27'h0000038f, 5'd7, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000077, 5'd19, 27'h0000010a, 5'd18, 27'h000000ac, 32'h00000400,
  1'd1,  5'd7, 27'h0000028d, 5'd17, 27'h000000e2, 5'd26, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000260, 5'd25, 27'h000003b6, 5'd9, 27'h00000049, 32'h00000400,
  1'd1,  5'd8, 27'h00000114, 5'd30, 27'h0000035d, 5'd17, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000078, 5'd30, 27'h00000225, 5'd28, 27'h000002de, 32'h00000400,
  1'd1,  5'd15, 27'h000002d1, 5'd8, 27'h000000f1, 5'd8, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001fd, 5'd7, 27'h000000d1, 5'd18, 27'h00000056, 32'h00000400,
  1'd1,  5'd16, 27'h0000000e, 5'd8, 27'h0000009a, 5'd30, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002ec, 5'd20, 27'h00000279, 5'd5, 27'h00000241, 32'h00000400,
  1'd1,  5'd16, 27'h000003d4, 5'd18, 27'h000003a5, 5'd20, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d1, 5'd19, 27'h000001ef, 5'd29, 27'h000003c9, 32'h00000400,
  1'd1,  5'd19, 27'h000003b7, 5'd26, 27'h00000245, 5'd6, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b5, 5'd29, 27'h00000359, 5'd20, 27'h000001be, 32'h00000400,
  1'd1,  5'd20, 27'h00000081, 5'd26, 27'h00000317, 5'd27, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000019b, 5'd8, 27'h000001cd, 5'd6, 27'h00000217, 32'h00000400,
  1'd1,  5'd28, 27'h000002a5, 5'd7, 27'h00000253, 5'd17, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a1, 5'd8, 27'h00000152, 5'd27, 27'h00000176, 32'h00000400,
  1'd1,  5'd29, 27'h000002ef, 5'd20, 27'h00000202, 5'd9, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e7, 5'd16, 27'h000001eb, 5'd16, 27'h00000092, 32'h00000400,
  1'd1,  5'd26, 27'h00000037, 5'd20, 27'h0000024b, 5'd29, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000023f, 5'd30, 27'h0000015b, 5'd6, 27'h0000019f, 32'h00000400,
  1'd1,  5'd29, 27'h0000037b, 5'd28, 27'h000003f5, 5'd18, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000030d, 5'd27, 27'h00000041, 5'd27, 27'h000001e9, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h00000070, 5'd4, 27'h0000010f, 5'd0, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003e1, 5'd1, 27'h000002f1, 5'd11, 27'h000002a7, 32'h00000400,
  1'd1,  5'd2, 27'h0000034a, 5'd4, 27'h0000009a, 5'd23, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000022, 5'd12, 27'h00000041, 5'd0, 27'h00000378, 32'h00000400,
  1'd1,  5'd3, 27'h000003aa, 5'd13, 27'h00000349, 5'd10, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d7, 5'd10, 27'h00000279, 5'd23, 27'h000003f7, 32'h00000400,
  1'd1,  5'd0, 27'h000002bb, 5'd23, 27'h000001e7, 5'd3, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002b7, 5'd22, 27'h00000266, 5'd14, 27'h00000339, 32'h00000400,
  1'd1,  5'd0, 27'h0000006d, 5'd25, 27'h00000104, 5'd21, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f6, 5'd1, 27'h000001b9, 5'd4, 27'h00000152, 32'h00000400,
  1'd1,  5'd14, 27'h000003c7, 5'd3, 27'h00000109, 5'd14, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c9, 5'd0, 27'h00000068, 5'd22, 27'h0000002e, 32'h00000400,
  1'd1,  5'd14, 27'h00000132, 5'd11, 27'h0000002d, 5'd1, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029f, 5'd12, 27'h000003e9, 5'd15, 27'h00000098, 32'h00000400,
  1'd1,  5'd14, 27'h00000286, 5'd13, 27'h00000068, 5'd25, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001fb, 5'd23, 27'h00000367, 5'd2, 27'h0000006b, 32'h00000400,
  1'd1,  5'd12, 27'h00000151, 5'd20, 27'h000003ea, 5'd10, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000035, 5'd25, 27'h00000305, 5'd23, 27'h000001c4, 32'h00000400,
  1'd1,  5'd24, 27'h00000210, 5'd2, 27'h0000028d, 5'd2, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001c5, 5'd3, 27'h000002f9, 5'd13, 27'h000000eb, 32'h00000400,
  1'd1,  5'd23, 27'h00000301, 5'd2, 27'h0000027f, 5'd24, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b6, 5'd11, 27'h000003a8, 5'd1, 27'h00000282, 32'h00000400,
  1'd1,  5'd23, 27'h000002d3, 5'd12, 27'h000002fc, 5'd14, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000a9, 5'd10, 27'h000003c4, 5'd23, 27'h0000028b, 32'h00000400,
  1'd1,  5'd22, 27'h00000110, 5'd22, 27'h00000223, 5'd4, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000017e, 5'd24, 27'h0000021e, 5'd12, 27'h000000f5, 32'h00000400,
  1'd1,  5'd21, 27'h0000020e, 5'd22, 27'h0000010d, 5'd24, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000054, 5'd4, 27'h000002bb, 5'd6, 27'h0000022e, 32'h00000400,
  1'd1,  5'd5, 27'h0000006e, 5'd1, 27'h0000006f, 5'd17, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000114, 5'd2, 27'h000002c5, 5'd30, 27'h000000a5, 32'h00000400,
  1'd1,  5'd5, 27'h00000013, 5'd12, 27'h000003c5, 5'd10, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001cb, 5'd12, 27'h000001ad, 5'd17, 27'h0000022f, 32'h00000400,
  1'd1,  5'd0, 27'h000003be, 5'd11, 27'h000001a2, 5'd27, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000a0, 5'd20, 27'h000002fd, 5'd6, 27'h000002e9, 32'h00000400,
  1'd1,  5'd3, 27'h000003e1, 5'd21, 27'h0000028d, 5'd16, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000290, 5'd21, 27'h0000028b, 5'd28, 27'h00000083, 32'h00000400,
  1'd1,  5'd14, 27'h000000ce, 5'd2, 27'h000002e6, 5'd6, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a6, 5'd4, 27'h000001f2, 5'd16, 27'h00000066, 32'h00000400,
  1'd1,  5'd14, 27'h0000034a, 5'd2, 27'h0000026c, 5'd27, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000350, 5'd14, 27'h000002f0, 5'd8, 27'h00000040, 32'h00000400,
  1'd1,  5'd14, 27'h00000067, 5'd12, 27'h000000cf, 5'd17, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000088, 5'd12, 27'h0000020c, 5'd27, 27'h000003f0, 32'h00000400,
  1'd1,  5'd13, 27'h000002ad, 5'd25, 27'h00000324, 5'd7, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b2, 5'd24, 27'h000001bc, 5'd18, 27'h0000025f, 32'h00000400,
  1'd1,  5'd14, 27'h000003d6, 5'd24, 27'h00000377, 5'd30, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003c4, 5'd1, 27'h00000218, 5'd9, 27'h000000b2, 32'h00000400,
  1'd1,  5'd23, 27'h0000007c, 5'd5, 27'h0000004d, 5'd15, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e2, 5'd2, 27'h0000034c, 5'd30, 27'h00000120, 32'h00000400,
  1'd1,  5'd23, 27'h000000ab, 5'd11, 27'h000001cf, 5'd6, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000009c, 5'd10, 27'h00000374, 5'd17, 27'h0000024a, 32'h00000400,
  1'd1,  5'd25, 27'h000001be, 5'd13, 27'h0000037c, 5'd27, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000010a, 5'd21, 27'h0000013d, 5'd6, 27'h0000036e, 32'h00000400,
  1'd1,  5'd23, 27'h0000019f, 5'd23, 27'h00000139, 5'd18, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000019f, 5'd24, 27'h00000211, 5'd30, 27'h00000242, 32'h00000400,
  1'd1,  5'd2, 27'h0000031d, 5'd8, 27'h0000033d, 5'd1, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003ef, 5'd8, 27'h0000017d, 5'd14, 27'h00000193, 32'h00000400,
  1'd1,  5'd4, 27'h00000177, 5'd8, 27'h0000037b, 5'd24, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d2, 5'd17, 27'h00000341, 5'd4, 27'h00000216, 32'h00000400,
  1'd1,  5'd0, 27'h00000038, 5'd19, 27'h0000035b, 5'd13, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000269, 5'd15, 27'h000003fb, 5'd23, 27'h000002f9, 32'h00000400,
  1'd1,  5'd4, 27'h00000242, 5'd28, 27'h000001f3, 5'd4, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000030f, 5'd26, 27'h00000245, 5'd11, 27'h0000002c, 32'h00000400,
  1'd1,  5'd2, 27'h0000014b, 5'd29, 27'h00000083, 5'd25, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000346, 5'd7, 27'h000003b6, 5'd1, 27'h0000027d, 32'h00000400,
  1'd1,  5'd14, 27'h0000024f, 5'd8, 27'h000000d3, 5'd12, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000010a, 5'd7, 27'h000003a1, 5'd23, 27'h000002ab, 32'h00000400,
  1'd1,  5'd11, 27'h00000207, 5'd18, 27'h00000272, 5'd3, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000165, 5'd16, 27'h00000342, 5'd11, 27'h00000268, 32'h00000400,
  1'd1,  5'd14, 27'h00000261, 5'd17, 27'h00000062, 5'd24, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000246, 5'd26, 27'h000001bb, 5'd0, 27'h0000015a, 32'h00000400,
  1'd1,  5'd12, 27'h0000028a, 5'd30, 27'h000003e5, 5'd15, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e1, 5'd29, 27'h000001e2, 5'd21, 27'h00000037, 32'h00000400,
  1'd1,  5'd24, 27'h00000317, 5'd7, 27'h000001bd, 5'd4, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000cd, 5'd6, 27'h00000163, 5'd11, 27'h000000f0, 32'h00000400,
  1'd1,  5'd21, 27'h000001bf, 5'd5, 27'h000003e7, 5'd23, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001d9, 5'd19, 27'h00000149, 5'd2, 27'h00000279, 32'h00000400,
  1'd1,  5'd22, 27'h000002ce, 5'd20, 27'h000000bc, 5'd12, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000352, 5'd16, 27'h000000d9, 5'd24, 27'h0000013a, 32'h00000400,
  1'd1,  5'd23, 27'h000002da, 5'd27, 27'h00000007, 5'd4, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003ac, 5'd26, 27'h000000c5, 5'd11, 27'h000002c6, 32'h00000400,
  1'd1,  5'd22, 27'h0000009a, 5'd29, 27'h00000348, 5'd21, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000006f, 5'd9, 27'h00000333, 5'd9, 27'h0000019b, 32'h00000400,
  1'd1,  5'd3, 27'h000001d8, 5'd7, 27'h0000027b, 5'd20, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002fd, 5'd6, 27'h0000033e, 5'd30, 27'h000000f5, 32'h00000400,
  1'd1,  5'd2, 27'h000001bb, 5'd19, 27'h000001f9, 5'd7, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ac, 5'd15, 27'h00000248, 5'd19, 27'h0000023e, 32'h00000400,
  1'd1,  5'd1, 27'h00000293, 5'd15, 27'h000002be, 5'd29, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000008d, 5'd28, 27'h00000357, 5'd9, 27'h00000196, 32'h00000400,
  1'd1,  5'd4, 27'h000003fe, 5'd30, 27'h000003e0, 5'd16, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022a, 5'd26, 27'h0000018f, 5'd27, 27'h00000331, 32'h00000400,
  1'd1,  5'd13, 27'h00000170, 5'd7, 27'h000001be, 5'd9, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000091, 5'd10, 27'h000000d0, 5'd20, 27'h0000006f, 32'h00000400,
  1'd1,  5'd10, 27'h00000175, 5'd7, 27'h00000190, 5'd27, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000245, 5'd19, 27'h000003a6, 5'd5, 27'h000002c7, 32'h00000400,
  1'd1,  5'd11, 27'h00000091, 5'd19, 27'h00000119, 5'd18, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000fc, 5'd19, 27'h000003be, 5'd26, 27'h000002b0, 32'h00000400,
  1'd1,  5'd14, 27'h000002ef, 5'd29, 27'h0000017c, 5'd7, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000071, 5'd29, 27'h0000034a, 5'd20, 27'h000000f0, 32'h00000400,
  1'd1,  5'd13, 27'h0000019e, 5'd30, 27'h000000c0, 5'd26, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000038f, 5'd7, 27'h000001c0, 5'd5, 27'h000003d9, 32'h00000400,
  1'd1,  5'd24, 27'h0000008d, 5'd5, 27'h00000380, 5'd19, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000312, 5'd6, 27'h000001dd, 5'd26, 27'h00000186, 32'h00000400,
  1'd1,  5'd23, 27'h000003df, 5'd20, 27'h00000272, 5'd6, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000394, 5'd15, 27'h000002ba, 5'd17, 27'h00000018, 32'h00000400,
  1'd1,  5'd22, 27'h0000011b, 5'd17, 27'h000002e1, 5'd28, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000373, 5'd25, 27'h000003a9, 5'd6, 27'h000001a1, 32'h00000400,
  1'd1,  5'd25, 27'h00000155, 5'd27, 27'h00000069, 5'd17, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000314, 5'd27, 27'h0000006b, 5'd27, 27'h0000027c, 32'h00000400,
  1'd1,  5'd8, 27'h00000262, 5'd4, 27'h000003ae, 5'd5, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001f3, 5'd2, 27'h00000125, 5'd19, 27'h00000051, 32'h00000400,
  1'd1,  5'd6, 27'h000000ad, 5'd2, 27'h00000080, 5'd30, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000096, 5'd14, 27'h000001de, 5'd3, 27'h00000296, 32'h00000400,
  1'd1,  5'd7, 27'h00000212, 5'd15, 27'h00000165, 5'd10, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000030a, 5'd13, 27'h00000128, 5'd23, 27'h0000039b, 32'h00000400,
  1'd1,  5'd9, 27'h00000246, 5'd24, 27'h00000335, 5'd3, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000019c, 5'd25, 27'h0000031e, 5'd13, 27'h000001ae, 32'h00000400,
  1'd1,  5'd7, 27'h00000104, 5'd21, 27'h00000397, 5'd24, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000361, 5'd0, 27'h000000dc, 5'd7, 27'h000002e3, 32'h00000400,
  1'd1,  5'd20, 27'h000000c8, 5'd5, 27'h00000062, 5'd16, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b6, 5'd2, 27'h00000268, 5'd25, 27'h00000376, 32'h00000400,
  1'd1,  5'd19, 27'h00000044, 5'd12, 27'h00000194, 5'd1, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000257, 5'd15, 27'h00000053, 5'd14, 27'h0000012a, 32'h00000400,
  1'd1,  5'd19, 27'h00000298, 5'd10, 27'h00000355, 5'd23, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000010, 5'd25, 27'h00000206, 5'd0, 27'h0000004f, 32'h00000400,
  1'd1,  5'd15, 27'h000002d6, 5'd24, 27'h000002cd, 5'd11, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000027f, 5'd22, 27'h00000284, 5'd21, 27'h00000047, 32'h00000400,
  1'd1,  5'd28, 27'h000001b1, 5'd5, 27'h00000008, 5'd0, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b2, 5'd1, 27'h000001a2, 5'd12, 27'h00000379, 32'h00000400,
  1'd1,  5'd29, 27'h00000306, 5'd4, 27'h00000372, 5'd24, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000091, 5'd14, 27'h000002b1, 5'd1, 27'h00000224, 32'h00000400,
  1'd1,  5'd28, 27'h00000276, 5'd12, 27'h000002bf, 5'd11, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001fd, 5'd10, 27'h00000226, 5'd20, 27'h00000344, 32'h00000400,
  1'd1,  5'd27, 27'h00000204, 5'd22, 27'h00000137, 5'd2, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003c1, 5'd25, 27'h00000006, 5'd12, 27'h0000021d, 32'h00000400,
  1'd1,  5'd30, 27'h000003de, 5'd23, 27'h0000005e, 5'd22, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f6, 5'd4, 27'h0000003c, 5'd1, 27'h0000021a, 32'h00000400,
  1'd1,  5'd7, 27'h000002f3, 5'd0, 27'h000001b9, 5'd14, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000032, 5'd1, 27'h000003e8, 5'd24, 27'h000003e0, 32'h00000400,
  1'd1,  5'd8, 27'h00000254, 5'd11, 27'h00000392, 5'd7, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003fc, 5'd10, 27'h0000034a, 5'd18, 27'h0000002c, 32'h00000400,
  1'd1,  5'd5, 27'h000000d4, 5'd14, 27'h000003eb, 5'd30, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b6, 5'd23, 27'h00000140, 5'd6, 27'h000000d2, 32'h00000400,
  1'd1,  5'd9, 27'h0000030d, 5'd24, 27'h00000088, 5'd17, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000387, 5'd23, 27'h00000388, 5'd28, 27'h0000034b, 32'h00000400,
  1'd1,  5'd19, 27'h0000000e, 5'd1, 27'h00000335, 5'd4, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000217, 5'd1, 27'h00000209, 5'd12, 27'h0000015b, 32'h00000400,
  1'd1,  5'd19, 27'h0000034f, 5'd0, 27'h000000dc, 5'd22, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002da, 5'd15, 27'h000001e4, 5'd7, 27'h0000007e, 32'h00000400,
  1'd1,  5'd17, 27'h00000160, 5'd11, 27'h0000000a, 5'd19, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000373, 5'd11, 27'h000000c5, 5'd27, 27'h000002cc, 32'h00000400,
  1'd1,  5'd19, 27'h000003ac, 5'd24, 27'h00000168, 5'd9, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003fd, 5'd23, 27'h00000390, 5'd15, 27'h00000363, 32'h00000400,
  1'd1,  5'd17, 27'h00000035, 5'd21, 27'h000001c3, 5'd30, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ac, 5'd1, 27'h00000202, 5'd7, 27'h000002d0, 32'h00000400,
  1'd1,  5'd27, 27'h000003c8, 5'd0, 27'h0000014e, 5'd16, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000021e, 5'd4, 27'h000003a8, 5'd26, 27'h00000112, 32'h00000400,
  1'd1,  5'd27, 27'h000000a6, 5'd14, 27'h00000023, 5'd8, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000015e, 5'd15, 27'h00000082, 5'd15, 27'h00000306, 32'h00000400,
  1'd1,  5'd28, 27'h000002bf, 5'd10, 27'h0000038c, 5'd26, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000063, 5'd22, 27'h00000046, 5'd8, 27'h0000000d, 32'h00000400,
  1'd1,  5'd26, 27'h00000357, 5'd25, 27'h00000082, 5'd20, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000013f, 5'd20, 27'h00000355, 5'd29, 27'h0000030e, 32'h00000400,
  1'd1,  5'd5, 27'h00000120, 5'd5, 27'h0000012c, 5'd3, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000027, 5'd6, 27'h00000373, 5'd11, 27'h0000008b, 32'h00000400,
  1'd1,  5'd8, 27'h00000046, 5'd10, 27'h0000013b, 5'd24, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000095, 5'd17, 27'h000002b0, 5'd0, 27'h00000328, 32'h00000400,
  1'd1,  5'd8, 27'h000002ad, 5'd20, 27'h0000017a, 5'd11, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000153, 5'd17, 27'h00000189, 5'd22, 27'h00000269, 32'h00000400,
  1'd1,  5'd9, 27'h000000fd, 5'd28, 27'h00000221, 5'd1, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000016, 5'd30, 27'h0000000d, 5'd14, 27'h0000030d, 32'h00000400,
  1'd1,  5'd5, 27'h00000261, 5'd27, 27'h00000157, 5'd21, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000189, 5'd6, 27'h0000025f, 5'd5, 27'h00000001, 32'h00000400,
  1'd1,  5'd18, 27'h00000368, 5'd7, 27'h00000304, 5'd13, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001a0, 5'd9, 27'h000002d2, 5'd24, 27'h00000337, 32'h00000400,
  1'd1,  5'd17, 27'h000002ef, 5'd20, 27'h00000253, 5'd3, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003b8, 5'd20, 27'h00000278, 5'd13, 27'h00000169, 32'h00000400,
  1'd1,  5'd17, 27'h00000376, 5'd15, 27'h00000343, 5'd21, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000162, 5'd28, 27'h000001aa, 5'd4, 27'h000001f1, 32'h00000400,
  1'd1,  5'd20, 27'h00000017, 5'd26, 27'h000001d0, 5'd14, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000049, 5'd26, 27'h000002d5, 5'd21, 27'h0000023b, 32'h00000400,
  1'd1,  5'd27, 27'h0000024c, 5'd6, 27'h0000010a, 5'd2, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000034, 5'd5, 27'h00000365, 5'd13, 27'h0000027d, 32'h00000400,
  1'd1,  5'd29, 27'h00000020, 5'd9, 27'h000002d7, 5'd25, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000028, 5'd20, 27'h000000b5, 5'd5, 27'h00000092, 32'h00000400,
  1'd1,  5'd29, 27'h00000366, 5'd18, 27'h000002ad, 5'd11, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000312, 5'd18, 27'h000002a9, 5'd24, 27'h00000239, 32'h00000400,
  1'd1,  5'd27, 27'h00000108, 5'd28, 27'h00000325, 5'd2, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000015c, 5'd29, 27'h000002d4, 5'd11, 27'h00000338, 32'h00000400,
  1'd1,  5'd28, 27'h0000021a, 5'd28, 27'h00000024, 5'd21, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005c, 5'd5, 27'h0000027c, 5'd9, 27'h0000037c, 32'h00000400,
  1'd1,  5'd9, 27'h000000f2, 5'd5, 27'h00000349, 5'd17, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000014a, 5'd9, 27'h0000006d, 5'd29, 27'h00000360, 32'h00000400,
  1'd1,  5'd9, 27'h0000003a, 5'd17, 27'h00000147, 5'd5, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a3, 5'd16, 27'h0000025a, 5'd20, 27'h000000af, 32'h00000400,
  1'd1,  5'd5, 27'h000000be, 5'd15, 27'h000002f7, 5'd30, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000033, 5'd27, 27'h0000001c, 5'd7, 27'h00000182, 32'h00000400,
  1'd1,  5'd9, 27'h00000022, 5'd29, 27'h000001b1, 5'd16, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000015d, 5'd26, 27'h000003e1, 5'd29, 27'h00000267, 32'h00000400,
  1'd1,  5'd17, 27'h00000272, 5'd7, 27'h00000293, 5'd6, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009a, 5'd7, 27'h0000001e, 5'd18, 27'h0000026e, 32'h00000400,
  1'd1,  5'd19, 27'h0000018c, 5'd9, 27'h00000221, 5'd27, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029b, 5'd19, 27'h00000390, 5'd6, 27'h0000035f, 32'h00000400,
  1'd1,  5'd16, 27'h000002d8, 5'd18, 27'h000001cf, 5'd20, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000102, 5'd19, 27'h00000282, 5'd26, 27'h0000039e, 32'h00000400,
  1'd1,  5'd19, 27'h00000364, 5'd29, 27'h000002a8, 5'd6, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f9, 5'd25, 27'h0000038c, 5'd15, 27'h0000028e, 32'h00000400,
  1'd1,  5'd18, 27'h0000029e, 5'd27, 27'h0000035c, 5'd26, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003ec, 5'd6, 27'h00000033, 5'd9, 27'h000003a0, 32'h00000400,
  1'd1,  5'd29, 27'h00000137, 5'd6, 27'h00000369, 5'd16, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000212, 5'd5, 27'h00000181, 5'd30, 27'h000000ab, 32'h00000400,
  1'd1,  5'd30, 27'h00000172, 5'd16, 27'h000003aa, 5'd8, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a6, 5'd18, 27'h0000033e, 5'd18, 27'h000003d4, 32'h00000400,
  1'd1,  5'd30, 27'h0000019b, 5'd17, 27'h00000359, 5'd28, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c2, 5'd27, 27'h00000173, 5'd9, 27'h00000077, 32'h00000400,
  1'd1,  5'd30, 27'h00000363, 5'd29, 27'h0000022c, 5'd20, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000003d, 5'd27, 27'h0000015b, 5'd30, 27'h00000102, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000100, 5'd1, 27'h0000034f, 5'd4, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000f2, 5'd0, 27'h0000015d, 5'd11, 27'h0000014b, 32'h00000400,
  1'd1,  5'd1, 27'h000003e7, 5'd4, 27'h0000027d, 5'd25, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ce, 5'd11, 27'h000003ff, 5'd4, 27'h00000070, 32'h00000400,
  1'd1,  5'd2, 27'h00000034, 5'd14, 27'h000000ed, 5'd10, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002e3, 5'd12, 27'h000003e0, 5'd21, 27'h000002a9, 32'h00000400,
  1'd1,  5'd1, 27'h00000240, 5'd22, 27'h0000018a, 5'd3, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a0, 5'd25, 27'h00000338, 5'd10, 27'h000003b6, 32'h00000400,
  1'd1,  5'd0, 27'h00000299, 5'd21, 27'h000000a1, 5'd24, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000020, 5'd3, 27'h00000231, 5'd5, 27'h00000038, 32'h00000400,
  1'd1,  5'd11, 27'h0000013e, 5'd0, 27'h000002d2, 5'd14, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000006d, 5'd2, 27'h00000249, 5'd25, 27'h000001e7, 32'h00000400,
  1'd1,  5'd12, 27'h00000199, 5'd15, 27'h00000154, 5'd2, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002fa, 5'd15, 27'h000001d3, 5'd12, 27'h000001ff, 32'h00000400,
  1'd1,  5'd14, 27'h0000015b, 5'd11, 27'h00000329, 5'd22, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000166, 5'd22, 27'h000002a2, 5'd0, 27'h00000335, 32'h00000400,
  1'd1,  5'd11, 27'h00000014, 5'd23, 27'h00000139, 5'd15, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000306, 5'd23, 27'h0000020e, 5'd21, 27'h00000071, 32'h00000400,
  1'd1,  5'd23, 27'h000001d9, 5'd3, 27'h0000032b, 5'd0, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000103, 5'd1, 27'h000003bd, 5'd13, 27'h0000020a, 32'h00000400,
  1'd1,  5'd24, 27'h000000c8, 5'd4, 27'h000003f2, 5'd25, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000309, 5'd10, 27'h000002b2, 5'd2, 27'h00000363, 32'h00000400,
  1'd1,  5'd23, 27'h0000012e, 5'd10, 27'h000003d3, 5'd13, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002df, 5'd13, 27'h00000186, 5'd23, 27'h0000011b, 32'h00000400,
  1'd1,  5'd23, 27'h000002d5, 5'd21, 27'h000002a7, 5'd2, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000365, 5'd24, 27'h0000009a, 5'd13, 27'h00000063, 32'h00000400,
  1'd1,  5'd22, 27'h0000019b, 5'd24, 27'h0000035d, 5'd25, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000035c, 5'd4, 27'h00000315, 5'd7, 27'h000003f9, 32'h00000400,
  1'd1,  5'd2, 27'h0000026d, 5'd4, 27'h00000205, 5'd15, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000eb, 5'd0, 27'h0000028a, 5'd26, 27'h000002af, 32'h00000400,
  1'd1,  5'd4, 27'h00000196, 5'd15, 27'h000001e8, 5'd8, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000235, 5'd13, 27'h000003d1, 5'd17, 27'h0000029c, 32'h00000400,
  1'd1,  5'd3, 27'h00000110, 5'd15, 27'h0000006b, 5'd29, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000148, 5'd21, 27'h0000027f, 5'd8, 27'h000002aa, 32'h00000400,
  1'd1,  5'd3, 27'h00000265, 5'd21, 27'h0000031f, 5'd18, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e9, 5'd25, 27'h00000204, 5'd28, 27'h000000d4, 32'h00000400,
  1'd1,  5'd11, 27'h0000021c, 5'd4, 27'h00000143, 5'd9, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001cd, 5'd4, 27'h0000002f, 5'd17, 27'h00000263, 32'h00000400,
  1'd1,  5'd15, 27'h0000013d, 5'd0, 27'h0000015f, 5'd27, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001ce, 5'd11, 27'h00000192, 5'd7, 27'h00000110, 32'h00000400,
  1'd1,  5'd14, 27'h000002a9, 5'd14, 27'h000000d2, 5'd18, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000143, 5'd11, 27'h00000245, 5'd27, 27'h00000160, 32'h00000400,
  1'd1,  5'd10, 27'h000003c1, 5'd25, 27'h0000033b, 5'd6, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b8, 5'd25, 27'h00000068, 5'd18, 27'h000000bd, 32'h00000400,
  1'd1,  5'd13, 27'h0000007e, 5'd21, 27'h000002fc, 5'd27, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021f, 5'd1, 27'h0000029d, 5'd7, 27'h00000320, 32'h00000400,
  1'd1,  5'd22, 27'h0000013c, 5'd2, 27'h00000331, 5'd19, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000fd, 5'd2, 27'h0000000e, 5'd30, 27'h00000095, 32'h00000400,
  1'd1,  5'd24, 27'h00000102, 5'd11, 27'h000002c7, 5'd8, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000007e, 5'd15, 27'h00000095, 5'd15, 27'h0000021f, 32'h00000400,
  1'd1,  5'd25, 27'h000001f9, 5'd10, 27'h00000237, 5'd29, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000159, 5'd21, 27'h0000009e, 5'd9, 27'h00000126, 32'h00000400,
  1'd1,  5'd24, 27'h00000232, 5'd23, 27'h00000209, 5'd20, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001e8, 5'd20, 27'h000003c3, 5'd29, 27'h0000030d, 32'h00000400,
  1'd1,  5'd2, 27'h0000005b, 5'd5, 27'h0000018d, 5'd2, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000142, 5'd9, 27'h000000be, 5'd13, 27'h0000037b, 32'h00000400,
  1'd1,  5'd1, 27'h00000166, 5'd10, 27'h00000051, 5'd23, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d4, 5'd15, 27'h0000025d, 5'd2, 27'h000000a6, 32'h00000400,
  1'd1,  5'd2, 27'h00000012, 5'd19, 27'h000003e0, 5'd13, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000025a, 5'd17, 27'h000000c7, 5'd23, 27'h0000031d, 32'h00000400,
  1'd1,  5'd4, 27'h0000006a, 5'd29, 27'h00000200, 5'd3, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000028b, 5'd28, 27'h000002e0, 5'd14, 27'h00000087, 32'h00000400,
  1'd1,  5'd1, 27'h0000007b, 5'd30, 27'h000002e4, 5'd21, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003eb, 5'd9, 27'h000003c2, 5'd4, 27'h00000244, 32'h00000400,
  1'd1,  5'd15, 27'h00000042, 5'd10, 27'h00000142, 5'd13, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000287, 5'd10, 27'h00000006, 5'd24, 27'h000001ca, 32'h00000400,
  1'd1,  5'd12, 27'h000003ca, 5'd18, 27'h00000065, 5'd3, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000170, 5'd19, 27'h000002ba, 5'd14, 27'h00000155, 32'h00000400,
  1'd1,  5'd15, 27'h00000129, 5'd17, 27'h000003ae, 5'd20, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000233, 5'd30, 27'h0000007e, 5'd2, 27'h00000157, 32'h00000400,
  1'd1,  5'd12, 27'h00000111, 5'd28, 27'h0000022a, 5'd10, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ec, 5'd26, 27'h0000026b, 5'd23, 27'h00000343, 32'h00000400,
  1'd1,  5'd24, 27'h000002f4, 5'd5, 27'h000002d6, 5'd0, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000014f, 5'd6, 27'h00000383, 5'd13, 27'h00000108, 32'h00000400,
  1'd1,  5'd25, 27'h00000072, 5'd10, 27'h0000002e, 5'd24, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000073, 5'd20, 27'h000001f1, 5'd3, 27'h0000004a, 32'h00000400,
  1'd1,  5'd24, 27'h000003a2, 5'd15, 27'h00000301, 5'd14, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000236, 5'd19, 27'h00000353, 5'd23, 27'h0000034a, 32'h00000400,
  1'd1,  5'd24, 27'h00000126, 5'd29, 27'h000000d6, 5'd2, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000054, 5'd28, 27'h00000050, 5'd15, 27'h000001b8, 32'h00000400,
  1'd1,  5'd23, 27'h00000138, 5'd30, 27'h000003bd, 5'd25, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000012c, 5'd7, 27'h000003dc, 5'd10, 27'h000000e7, 32'h00000400,
  1'd1,  5'd1, 27'h00000058, 5'd6, 27'h000003b6, 5'd20, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000281, 5'd9, 27'h000000b1, 5'd28, 27'h00000353, 32'h00000400,
  1'd1,  5'd1, 27'h00000030, 5'd19, 27'h00000371, 5'd10, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d9, 5'd16, 27'h000002ce, 5'd20, 27'h000001b1, 32'h00000400,
  1'd1,  5'd3, 27'h000000bf, 5'd17, 27'h000002b6, 5'd29, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000026, 5'd27, 27'h000003a1, 5'd6, 27'h000000be, 32'h00000400,
  1'd1,  5'd3, 27'h00000358, 5'd29, 27'h0000030e, 5'd17, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000246, 5'd30, 27'h0000005e, 5'd30, 27'h000000a8, 32'h00000400,
  1'd1,  5'd13, 27'h00000208, 5'd8, 27'h000002a3, 5'd8, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003e6, 5'd6, 27'h00000267, 5'd15, 27'h0000027b, 32'h00000400,
  1'd1,  5'd14, 27'h000002c5, 5'd9, 27'h00000378, 5'd30, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000024b, 5'd16, 27'h00000381, 5'd6, 27'h00000086, 32'h00000400,
  1'd1,  5'd12, 27'h00000123, 5'd18, 27'h00000276, 5'd18, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003ca, 5'd19, 27'h00000153, 5'd26, 27'h0000003d, 32'h00000400,
  1'd1,  5'd13, 27'h000001ac, 5'd28, 27'h0000005b, 5'd7, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000019b, 5'd29, 27'h0000018a, 5'd19, 27'h0000029e, 32'h00000400,
  1'd1,  5'd14, 27'h000000ef, 5'd29, 27'h000000b4, 5'd29, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000da, 5'd6, 27'h000002d3, 5'd7, 27'h000000c9, 32'h00000400,
  1'd1,  5'd24, 27'h0000009f, 5'd5, 27'h000003b0, 5'd20, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000396, 5'd5, 27'h0000017b, 5'd27, 27'h000002c3, 32'h00000400,
  1'd1,  5'd25, 27'h00000351, 5'd20, 27'h000001ac, 5'd8, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000018, 5'd16, 27'h00000266, 5'd20, 27'h00000106, 32'h00000400,
  1'd1,  5'd25, 27'h0000000e, 5'd16, 27'h000003c5, 5'd27, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000102, 5'd29, 27'h000001c2, 5'd7, 27'h00000350, 32'h00000400,
  1'd1,  5'd23, 27'h0000039a, 5'd28, 27'h00000105, 5'd19, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b6, 5'd30, 27'h00000098, 5'd27, 27'h000001ce, 32'h00000400,
  1'd1,  5'd8, 27'h00000100, 5'd0, 27'h000002a8, 5'd5, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002eb, 5'd4, 27'h00000006, 5'd19, 27'h00000371, 32'h00000400,
  1'd1,  5'd7, 27'h0000024b, 5'd2, 27'h00000059, 5'd26, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000d6, 5'd14, 27'h0000024b, 5'd2, 27'h000003af, 32'h00000400,
  1'd1,  5'd10, 27'h00000012, 5'd10, 27'h00000242, 5'd14, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000156, 5'd14, 27'h0000010e, 5'd22, 27'h00000226, 32'h00000400,
  1'd1,  5'd5, 27'h000002be, 5'd20, 27'h0000034c, 5'd0, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034b, 5'd25, 27'h000002dd, 5'd14, 27'h00000202, 32'h00000400,
  1'd1,  5'd9, 27'h0000029f, 5'd24, 27'h0000028d, 5'd23, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000009e, 5'd4, 27'h000001b5, 5'd8, 27'h00000194, 32'h00000400,
  1'd1,  5'd20, 27'h000000e6, 5'd1, 27'h00000236, 5'd20, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000300, 5'd3, 27'h000001d3, 5'd30, 27'h0000024c, 32'h00000400,
  1'd1,  5'd19, 27'h00000101, 5'd13, 27'h000003c8, 5'd2, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ef, 5'd12, 27'h00000159, 5'd14, 27'h0000022d, 32'h00000400,
  1'd1,  5'd17, 27'h000002e2, 5'd12, 27'h00000058, 5'd24, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000019e, 5'd23, 27'h00000289, 5'd1, 27'h00000018, 32'h00000400,
  1'd1,  5'd16, 27'h000002cb, 5'd20, 27'h000002e0, 5'd11, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003cf, 5'd22, 27'h00000053, 5'd23, 27'h00000133, 32'h00000400,
  1'd1,  5'd30, 27'h00000264, 5'd3, 27'h000003ad, 5'd2, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000165, 5'd2, 27'h00000176, 5'd14, 27'h000000b5, 32'h00000400,
  1'd1,  5'd26, 27'h000000eb, 5'd0, 27'h00000212, 5'd25, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000272, 5'd14, 27'h000000b4, 5'd4, 27'h00000087, 32'h00000400,
  1'd1,  5'd27, 27'h000002fc, 5'd12, 27'h00000260, 5'd13, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000011c, 5'd13, 27'h0000012d, 5'd20, 27'h000002b4, 32'h00000400,
  1'd1,  5'd29, 27'h00000352, 5'd24, 27'h0000005e, 5'd3, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d2, 5'd22, 27'h00000038, 5'd13, 27'h000002bf, 32'h00000400,
  1'd1,  5'd29, 27'h00000140, 5'd24, 27'h000003bd, 5'd24, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ab, 5'd4, 27'h000000a4, 5'd4, 27'h0000012c, 32'h00000400,
  1'd1,  5'd8, 27'h000001d5, 5'd4, 27'h00000096, 5'd13, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ef, 5'd4, 27'h000001eb, 5'd24, 27'h00000055, 32'h00000400,
  1'd1,  5'd6, 27'h000003ab, 5'd13, 27'h0000010d, 5'd5, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000033c, 5'd11, 27'h00000328, 5'd18, 27'h0000031a, 32'h00000400,
  1'd1,  5'd6, 27'h000000c1, 5'd11, 27'h00000250, 5'd27, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003fd, 5'd25, 27'h00000050, 5'd6, 27'h00000329, 32'h00000400,
  1'd1,  5'd7, 27'h000000e7, 5'd22, 27'h0000002b, 5'd18, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000216, 5'd22, 27'h0000018c, 5'd30, 27'h00000246, 32'h00000400,
  1'd1,  5'd18, 27'h0000031b, 5'd4, 27'h00000280, 5'd5, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000024, 5'd2, 27'h0000024c, 5'd13, 27'h000001fe, 32'h00000400,
  1'd1,  5'd20, 27'h000000e3, 5'd3, 27'h0000038a, 5'd21, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000362, 5'd15, 27'h0000019b, 5'd10, 27'h0000013f, 32'h00000400,
  1'd1,  5'd16, 27'h000002b8, 5'd14, 27'h000002fd, 5'd17, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001dc, 5'd13, 27'h0000038f, 5'd29, 27'h0000031a, 32'h00000400,
  1'd1,  5'd16, 27'h00000258, 5'd22, 27'h00000002, 5'd6, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000066, 5'd22, 27'h000002c7, 5'd19, 27'h0000013e, 32'h00000400,
  1'd1,  5'd17, 27'h00000354, 5'd25, 27'h00000033, 5'd28, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003cf, 5'd2, 27'h00000210, 5'd9, 27'h000001cf, 32'h00000400,
  1'd1,  5'd29, 27'h0000015d, 5'd2, 27'h0000017e, 5'd16, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000140, 5'd5, 27'h00000033, 5'd30, 27'h00000371, 32'h00000400,
  1'd1,  5'd30, 27'h00000276, 5'd13, 27'h00000174, 5'd7, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000215, 5'd13, 27'h000000e1, 5'd18, 27'h000003d7, 32'h00000400,
  1'd1,  5'd29, 27'h000001f4, 5'd13, 27'h00000194, 5'd26, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002ee, 5'd21, 27'h000000c4, 5'd7, 27'h00000033, 32'h00000400,
  1'd1,  5'd27, 27'h00000123, 5'd23, 27'h000000d4, 5'd19, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000306, 5'd21, 27'h000001fb, 5'd26, 27'h00000218, 32'h00000400,
  1'd1,  5'd9, 27'h00000314, 5'd6, 27'h00000131, 5'd2, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000283, 5'd7, 27'h00000080, 5'd12, 27'h00000368, 32'h00000400,
  1'd1,  5'd9, 27'h0000010f, 5'd6, 27'h00000373, 5'd25, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000007, 5'd20, 27'h0000008f, 5'd4, 27'h00000209, 32'h00000400,
  1'd1,  5'd9, 27'h00000167, 5'd18, 27'h00000395, 5'd14, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000027f, 5'd16, 27'h000003ea, 5'd24, 27'h00000223, 32'h00000400,
  1'd1,  5'd9, 27'h0000021f, 5'd26, 27'h000002d9, 5'd4, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000165, 5'd29, 27'h00000346, 5'd10, 27'h000003b0, 32'h00000400,
  1'd1,  5'd7, 27'h0000012e, 5'd30, 27'h00000099, 5'd25, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000384, 5'd5, 27'h000003b8, 5'd3, 27'h000001e5, 32'h00000400,
  1'd1,  5'd16, 27'h0000010e, 5'd8, 27'h000000cf, 5'd12, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a7, 5'd7, 27'h00000251, 5'd21, 27'h00000075, 32'h00000400,
  1'd1,  5'd19, 27'h00000014, 5'd18, 27'h000000ea, 5'd3, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ba, 5'd17, 27'h00000065, 5'd12, 27'h00000083, 32'h00000400,
  1'd1,  5'd18, 27'h00000068, 5'd19, 27'h0000002e, 5'd23, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003bf, 5'd29, 27'h000002f4, 5'd4, 27'h0000005f, 32'h00000400,
  1'd1,  5'd18, 27'h00000330, 5'd30, 27'h0000033f, 5'd12, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000249, 5'd27, 27'h00000228, 5'd22, 27'h00000073, 32'h00000400,
  1'd1,  5'd29, 27'h0000017b, 5'd8, 27'h0000019c, 5'd3, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000025f, 5'd7, 27'h00000014, 5'd14, 27'h0000016d, 32'h00000400,
  1'd1,  5'd28, 27'h00000267, 5'd7, 27'h00000073, 5'd25, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c2, 5'd16, 27'h000002d3, 5'd0, 27'h00000245, 32'h00000400,
  1'd1,  5'd28, 27'h0000006e, 5'd17, 27'h00000063, 5'd11, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001fb, 5'd20, 27'h000001e7, 5'd21, 27'h000003c8, 32'h00000400,
  1'd1,  5'd28, 27'h0000029e, 5'd28, 27'h00000057, 5'd0, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003e4, 5'd26, 27'h00000040, 5'd14, 27'h000000c4, 32'h00000400,
  1'd1,  5'd29, 27'h0000016d, 5'd28, 27'h0000020f, 5'd25, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fa, 5'd8, 27'h000002ae, 5'd6, 27'h00000053, 32'h00000400,
  1'd1,  5'd10, 27'h000000cf, 5'd8, 27'h0000028b, 5'd19, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020c, 5'd7, 27'h00000122, 5'd29, 27'h0000024f, 32'h00000400,
  1'd1,  5'd6, 27'h0000030b, 5'd20, 27'h000001e3, 5'd6, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000026e, 5'd17, 27'h00000208, 5'd18, 27'h000000fd, 32'h00000400,
  1'd1,  5'd8, 27'h00000086, 5'd20, 27'h0000002b, 5'd27, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021d, 5'd26, 27'h00000298, 5'd7, 27'h00000311, 32'h00000400,
  1'd1,  5'd8, 27'h00000154, 5'd30, 27'h000001d3, 5'd20, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003b4, 5'd27, 27'h0000007a, 5'd29, 27'h0000032d, 32'h00000400,
  1'd1,  5'd17, 27'h0000015f, 5'd5, 27'h000003a6, 5'd6, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002bf, 5'd8, 27'h00000288, 5'd15, 27'h00000322, 32'h00000400,
  1'd1,  5'd17, 27'h0000021e, 5'd8, 27'h0000033f, 5'd30, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000393, 5'd19, 27'h00000350, 5'd10, 27'h00000113, 32'h00000400,
  1'd1,  5'd19, 27'h000001fa, 5'd20, 27'h00000259, 5'd20, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000031e, 5'd16, 27'h000001f2, 5'd30, 27'h000001f5, 32'h00000400,
  1'd1,  5'd15, 27'h000003d1, 5'd30, 27'h0000011d, 5'd9, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b7, 5'd30, 27'h00000140, 5'd20, 27'h0000008a, 32'h00000400,
  1'd1,  5'd17, 27'h000003de, 5'd26, 27'h00000055, 5'd28, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000023f, 5'd9, 27'h000000b5, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd28, 27'h000000c8, 5'd8, 27'h00000053, 5'd17, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000343, 5'd6, 27'h00000100, 5'd28, 27'h0000034c, 32'h00000400,
  1'd1,  5'd29, 27'h00000339, 5'd17, 27'h000000cf, 5'd7, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000002e, 5'd17, 27'h00000218, 5'd17, 27'h00000145, 32'h00000400,
  1'd1,  5'd28, 27'h000000fb, 5'd19, 27'h0000034e, 5'd27, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000124, 5'd30, 27'h00000208, 5'd10, 27'h0000014f, 32'h00000400,
  1'd1,  5'd30, 27'h0000022c, 5'd29, 27'h0000013e, 5'd17, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b8, 5'd27, 27'h0000006d, 5'd27, 27'h00000129, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003b6, 5'd1, 27'h000002d2, 5'd4, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000011e, 5'd0, 27'h0000001f, 5'd14, 27'h00000307, 32'h00000400,
  1'd1,  5'd1, 27'h000001c1, 5'd0, 27'h0000029b, 5'd25, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000279, 5'd13, 27'h0000010b, 5'd1, 27'h000003f8, 32'h00000400,
  1'd1,  5'd4, 27'h00000283, 5'd10, 27'h000001e3, 5'd13, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000294, 5'd13, 27'h000003ef, 5'd23, 27'h00000177, 32'h00000400,
  1'd1,  5'd4, 27'h00000219, 5'd23, 27'h0000011a, 5'd2, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001aa, 5'd20, 27'h00000373, 5'd14, 27'h000002a1, 32'h00000400,
  1'd1,  5'd4, 27'h000002bd, 5'd23, 27'h00000091, 5'd21, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013e, 5'd3, 27'h0000017b, 5'd3, 27'h000003a4, 32'h00000400,
  1'd1,  5'd11, 27'h00000311, 5'd2, 27'h00000040, 5'd12, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000287, 5'd2, 27'h00000091, 5'd20, 27'h000002b9, 32'h00000400,
  1'd1,  5'd10, 27'h000002e7, 5'd14, 27'h00000161, 5'd5, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000d2, 5'd11, 27'h00000204, 5'd14, 27'h0000003f, 32'h00000400,
  1'd1,  5'd14, 27'h00000302, 5'd12, 27'h00000071, 5'd24, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000021d, 5'd22, 27'h0000005c, 5'd4, 27'h000003de, 32'h00000400,
  1'd1,  5'd11, 27'h000003b6, 5'd20, 27'h000002ae, 5'd15, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000368, 5'd23, 27'h00000280, 5'd21, 27'h0000015c, 32'h00000400,
  1'd1,  5'd25, 27'h00000004, 5'd1, 27'h00000282, 5'd4, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001c9, 5'd3, 27'h00000156, 5'd14, 27'h000002e8, 32'h00000400,
  1'd1,  5'd22, 27'h000001f2, 5'd4, 27'h000001b0, 5'd22, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000023c, 5'd14, 27'h00000020, 5'd1, 27'h000001e1, 32'h00000400,
  1'd1,  5'd24, 27'h00000269, 5'd15, 27'h00000092, 5'd12, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001cc, 5'd11, 27'h00000202, 5'd23, 27'h00000032, 32'h00000400,
  1'd1,  5'd22, 27'h00000261, 5'd25, 27'h00000041, 5'd3, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ab, 5'd25, 27'h00000157, 5'd12, 27'h00000388, 32'h00000400,
  1'd1,  5'd25, 27'h00000229, 5'd21, 27'h00000072, 5'd24, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b8, 5'd2, 27'h000000d2, 5'd7, 27'h00000085, 32'h00000400,
  1'd1,  5'd0, 27'h00000033, 5'd3, 27'h000003aa, 5'd20, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000338, 5'd2, 27'h000003a3, 5'd29, 27'h000003ed, 32'h00000400,
  1'd1,  5'd1, 27'h000000e1, 5'd13, 27'h00000335, 5'd5, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d6, 5'd12, 27'h00000189, 5'd19, 27'h0000005d, 32'h00000400,
  1'd1,  5'd2, 27'h00000400, 5'd14, 27'h00000151, 5'd28, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003c0, 5'd22, 27'h000000c6, 5'd5, 27'h000001f0, 32'h00000400,
  1'd1,  5'd5, 27'h0000007f, 5'd23, 27'h0000001e, 5'd19, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000343, 5'd22, 27'h00000062, 5'd30, 27'h000002ee, 32'h00000400,
  1'd1,  5'd10, 27'h0000032f, 5'd3, 27'h00000244, 5'd6, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b0, 5'd1, 27'h000002ad, 5'd17, 27'h000001c4, 32'h00000400,
  1'd1,  5'd10, 27'h000001ee, 5'd2, 27'h00000158, 5'd29, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000bd, 5'd12, 27'h000003be, 5'd8, 27'h000001fb, 32'h00000400,
  1'd1,  5'd15, 27'h000001b4, 5'd10, 27'h0000029a, 5'd16, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000083, 5'd14, 27'h0000035b, 5'd26, 27'h000002e3, 32'h00000400,
  1'd1,  5'd15, 27'h000001c2, 5'd21, 27'h00000064, 5'd5, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002dd, 5'd22, 27'h0000032d, 5'd19, 27'h0000008f, 32'h00000400,
  1'd1,  5'd13, 27'h0000031e, 5'd21, 27'h000000e2, 5'd30, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000289, 5'd0, 27'h00000316, 5'd5, 27'h000002e4, 32'h00000400,
  1'd1,  5'd24, 27'h00000017, 5'd2, 27'h000002a2, 5'd20, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000159, 5'd1, 27'h00000388, 5'd28, 27'h00000049, 32'h00000400,
  1'd1,  5'd24, 27'h0000011f, 5'd15, 27'h0000000b, 5'd8, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000234, 5'd14, 27'h000000c4, 5'd16, 27'h000000d2, 32'h00000400,
  1'd1,  5'd24, 27'h0000025e, 5'd10, 27'h000003a5, 5'd29, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fa, 5'd23, 27'h0000015b, 5'd7, 27'h00000292, 32'h00000400,
  1'd1,  5'd20, 27'h000003f0, 5'd21, 27'h0000028f, 5'd16, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e1, 5'd24, 27'h0000039d, 5'd30, 27'h000003eb, 32'h00000400,
  1'd1,  5'd4, 27'h000000e1, 5'd9, 27'h00000130, 5'd3, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000347, 5'd5, 27'h000002f3, 5'd10, 27'h0000037a, 32'h00000400,
  1'd1,  5'd1, 27'h000001d0, 5'd6, 27'h000002a4, 5'd23, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000066, 5'd19, 27'h0000000b, 5'd1, 27'h0000012d, 32'h00000400,
  1'd1,  5'd0, 27'h00000152, 5'd15, 27'h00000270, 5'd11, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001c7, 5'd20, 27'h00000048, 5'd21, 27'h00000366, 32'h00000400,
  1'd1,  5'd3, 27'h0000022c, 5'd30, 27'h000000a8, 5'd0, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003af, 5'd29, 27'h00000114, 5'd14, 27'h0000019f, 32'h00000400,
  1'd1,  5'd4, 27'h00000254, 5'd28, 27'h0000029e, 5'd21, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000011e, 5'd5, 27'h0000031d, 5'd1, 27'h00000188, 32'h00000400,
  1'd1,  5'd10, 27'h000003dd, 5'd8, 27'h000001a7, 5'd14, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000019d, 5'd9, 27'h0000004e, 5'd24, 27'h000003e9, 32'h00000400,
  1'd1,  5'd14, 27'h000003fd, 5'd15, 27'h000002bc, 5'd4, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ef, 5'd20, 27'h0000011b, 5'd10, 27'h000001d4, 32'h00000400,
  1'd1,  5'd11, 27'h00000078, 5'd18, 27'h000003d7, 5'd21, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f6, 5'd30, 27'h000002ec, 5'd1, 27'h00000183, 32'h00000400,
  1'd1,  5'd14, 27'h000001e9, 5'd30, 27'h000003dc, 5'd14, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000217, 5'd29, 27'h000003e3, 5'd25, 27'h0000012f, 32'h00000400,
  1'd1,  5'd23, 27'h0000019f, 5'd6, 27'h000002e3, 5'd1, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000223, 5'd9, 27'h000003fb, 5'd15, 27'h00000198, 32'h00000400,
  1'd1,  5'd25, 27'h000002b8, 5'd9, 27'h00000331, 5'd24, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000bb, 5'd20, 27'h00000132, 5'd4, 27'h000000fe, 32'h00000400,
  1'd1,  5'd21, 27'h000002ef, 5'd19, 27'h0000018e, 5'd11, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002c2, 5'd16, 27'h00000338, 5'd25, 27'h00000091, 32'h00000400,
  1'd1,  5'd23, 27'h000001d9, 5'd30, 27'h00000041, 5'd3, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f8, 5'd27, 27'h0000035b, 5'd12, 27'h00000085, 32'h00000400,
  1'd1,  5'd23, 27'h0000005f, 5'd29, 27'h00000141, 5'd22, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000002, 5'd10, 27'h000000ee, 5'd9, 27'h0000007d, 32'h00000400,
  1'd1,  5'd0, 27'h00000073, 5'd8, 27'h000001f3, 5'd15, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002fa, 5'd6, 27'h00000364, 5'd27, 27'h0000035a, 32'h00000400,
  1'd1,  5'd4, 27'h0000029a, 5'd17, 27'h000003ab, 5'd10, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000195, 5'd18, 27'h00000323, 5'd16, 27'h000003f7, 32'h00000400,
  1'd1,  5'd4, 27'h000002f7, 5'd19, 27'h000003bc, 5'd26, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000216, 5'd27, 27'h00000009, 5'd9, 27'h000003f6, 32'h00000400,
  1'd1,  5'd1, 27'h000002ef, 5'd30, 27'h00000027, 5'd15, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039b, 5'd26, 27'h00000395, 5'd27, 27'h0000008b, 32'h00000400,
  1'd1,  5'd10, 27'h000002f6, 5'd8, 27'h00000358, 5'd9, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ca, 5'd7, 27'h0000025f, 5'd20, 27'h0000019e, 32'h00000400,
  1'd1,  5'd12, 27'h000003d0, 5'd10, 27'h000000da, 5'd30, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000333, 5'd16, 27'h0000008f, 5'd5, 27'h0000036e, 32'h00000400,
  1'd1,  5'd12, 27'h0000035e, 5'd18, 27'h000000f8, 5'd18, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c4, 5'd18, 27'h0000039f, 5'd26, 27'h00000172, 32'h00000400,
  1'd1,  5'd12, 27'h0000037f, 5'd29, 27'h000002a2, 5'd8, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000319, 5'd26, 27'h000002c7, 5'd20, 27'h00000121, 32'h00000400,
  1'd1,  5'd15, 27'h0000004a, 5'd27, 27'h000001ff, 5'd26, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000039e, 5'd6, 27'h0000019f, 5'd8, 27'h000002cc, 32'h00000400,
  1'd1,  5'd23, 27'h0000013e, 5'd6, 27'h000002d9, 5'd17, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000037a, 5'd6, 27'h00000155, 5'd30, 27'h00000147, 32'h00000400,
  1'd1,  5'd24, 27'h0000029b, 5'd20, 27'h0000023b, 5'd9, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001e0, 5'd18, 27'h00000012, 5'd15, 27'h000002cd, 32'h00000400,
  1'd1,  5'd21, 27'h0000014f, 5'd16, 27'h000002ca, 5'd25, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003fc, 5'd28, 27'h00000315, 5'd8, 27'h00000262, 32'h00000400,
  1'd1,  5'd24, 27'h000000ea, 5'd30, 27'h000001c1, 5'd20, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000017a, 5'd26, 27'h0000039d, 5'd28, 27'h0000034c, 32'h00000400,
  1'd1,  5'd10, 27'h00000081, 5'd1, 27'h000003d5, 5'd5, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b0, 5'd4, 27'h000000fa, 5'd19, 27'h00000343, 32'h00000400,
  1'd1,  5'd7, 27'h000003e2, 5'd3, 27'h000003af, 5'd28, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003c0, 5'd11, 27'h000002aa, 5'd0, 27'h00000064, 32'h00000400,
  1'd1,  5'd6, 27'h000003f5, 5'd15, 27'h000000e4, 5'd11, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000014, 5'd14, 27'h000000fc, 5'd23, 27'h000003d9, 32'h00000400,
  1'd1,  5'd9, 27'h000003da, 5'd24, 27'h0000007c, 5'd1, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000382, 5'd22, 27'h00000315, 5'd12, 27'h0000035b, 32'h00000400,
  1'd1,  5'd6, 27'h000002af, 5'd20, 27'h0000035a, 5'd24, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003c1, 5'd2, 27'h00000304, 5'd10, 27'h000000bd, 32'h00000400,
  1'd1,  5'd16, 27'h0000032c, 5'd3, 27'h00000340, 5'd16, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f7, 5'd3, 27'h00000176, 5'd28, 27'h000002ac, 32'h00000400,
  1'd1,  5'd19, 27'h00000017, 5'd12, 27'h00000281, 5'd1, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000022, 5'd11, 27'h000003c4, 5'd12, 27'h000002c1, 32'h00000400,
  1'd1,  5'd18, 27'h00000114, 5'd14, 27'h00000313, 5'd22, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000286, 5'd20, 27'h00000335, 5'd0, 27'h00000248, 32'h00000400,
  1'd1,  5'd17, 27'h0000033e, 5'd22, 27'h00000167, 5'd11, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000087, 5'd20, 27'h000002ce, 5'd24, 27'h000001d3, 32'h00000400,
  1'd1,  5'd28, 27'h0000002c, 5'd3, 27'h0000015a, 5'd3, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000256, 5'd0, 27'h00000093, 5'd13, 27'h00000271, 32'h00000400,
  1'd1,  5'd28, 27'h000002e3, 5'd0, 27'h00000144, 5'd23, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000262, 5'd12, 27'h0000033e, 5'd0, 27'h000001e1, 32'h00000400,
  1'd1,  5'd30, 27'h0000020f, 5'd14, 27'h000000b3, 5'd14, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a2, 5'd14, 27'h0000003b, 5'd21, 27'h000001a5, 32'h00000400,
  1'd1,  5'd26, 27'h000001f4, 5'd22, 27'h000003e5, 5'd2, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000274, 5'd25, 27'h00000347, 5'd12, 27'h0000007d, 32'h00000400,
  1'd1,  5'd28, 27'h00000044, 5'd25, 27'h000000f7, 5'd23, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b7, 5'd1, 27'h000003f2, 5'd3, 27'h000000fc, 32'h00000400,
  1'd1,  5'd5, 27'h000001a1, 5'd1, 27'h000000a1, 5'd11, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000f5, 5'd4, 27'h000002d0, 5'd21, 27'h000000c7, 32'h00000400,
  1'd1,  5'd7, 27'h000002c6, 5'd12, 27'h000000a1, 5'd5, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000027b, 5'd12, 27'h0000034c, 5'd17, 27'h00000033, 32'h00000400,
  1'd1,  5'd6, 27'h0000030f, 5'd13, 27'h00000123, 5'd26, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000395, 5'd23, 27'h00000215, 5'd6, 27'h0000004c, 32'h00000400,
  1'd1,  5'd6, 27'h00000032, 5'd24, 27'h00000083, 5'd19, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000117, 5'd24, 27'h000003d5, 5'd28, 27'h00000139, 32'h00000400,
  1'd1,  5'd19, 27'h000003e8, 5'd3, 27'h0000011b, 5'd0, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000023d, 5'd3, 27'h0000018c, 5'd14, 27'h000003dd, 32'h00000400,
  1'd1,  5'd16, 27'h000003ce, 5'd0, 27'h00000196, 5'd24, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000373, 5'd13, 27'h000001a4, 5'd7, 27'h0000029a, 32'h00000400,
  1'd1,  5'd17, 27'h000003f5, 5'd15, 27'h000001f1, 5'd18, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000002d, 5'd12, 27'h00000011, 5'd26, 27'h000000c2, 32'h00000400,
  1'd1,  5'd20, 27'h000000e6, 5'd25, 27'h00000063, 5'd5, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001cc, 5'd21, 27'h000003b6, 5'd18, 27'h000002a6, 32'h00000400,
  1'd1,  5'd16, 27'h00000122, 5'd22, 27'h000003ff, 5'd26, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d1, 5'd5, 27'h0000009a, 5'd5, 27'h0000010e, 32'h00000400,
  1'd1,  5'd30, 27'h0000000d, 5'd5, 27'h0000002e, 5'd15, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000026a, 5'd5, 27'h00000057, 5'd27, 27'h00000017, 32'h00000400,
  1'd1,  5'd26, 27'h000000c4, 5'd13, 27'h0000025e, 5'd6, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000353, 5'd11, 27'h000001b0, 5'd20, 27'h000000a5, 32'h00000400,
  1'd1,  5'd28, 27'h0000012d, 5'd14, 27'h0000008a, 5'd25, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025d, 5'd21, 27'h0000010f, 5'd6, 27'h00000249, 32'h00000400,
  1'd1,  5'd27, 27'h00000109, 5'd25, 27'h0000013d, 5'd17, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038c, 5'd22, 27'h00000187, 5'd27, 27'h00000245, 32'h00000400,
  1'd1,  5'd6, 27'h00000165, 5'd9, 27'h000001df, 5'd2, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e5, 5'd9, 27'h00000259, 5'd10, 27'h000002df, 32'h00000400,
  1'd1,  5'd5, 27'h000002d7, 5'd6, 27'h00000137, 5'd23, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e7, 5'd20, 27'h00000038, 5'd2, 27'h000000a2, 32'h00000400,
  1'd1,  5'd9, 27'h00000222, 5'd16, 27'h00000017, 5'd10, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000003e, 5'd18, 27'h000002f3, 5'd21, 27'h000000e5, 32'h00000400,
  1'd1,  5'd6, 27'h000000ba, 5'd27, 27'h00000362, 5'd1, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003fb, 5'd29, 27'h00000130, 5'd12, 27'h0000009f, 32'h00000400,
  1'd1,  5'd8, 27'h000002ee, 5'd28, 27'h000002c4, 5'd21, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000337, 5'd9, 27'h0000036b, 5'd2, 27'h00000396, 32'h00000400,
  1'd1,  5'd17, 27'h0000038e, 5'd8, 27'h00000373, 5'd13, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003cd, 5'd6, 27'h0000012c, 5'd24, 27'h000002c9, 32'h00000400,
  1'd1,  5'd16, 27'h0000020e, 5'd16, 27'h000002c3, 5'd0, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a3, 5'd18, 27'h000002cd, 5'd15, 27'h00000159, 32'h00000400,
  1'd1,  5'd16, 27'h000001ab, 5'd17, 27'h000002ff, 5'd21, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000305, 5'd26, 27'h000003c6, 5'd1, 27'h0000005b, 32'h00000400,
  1'd1,  5'd16, 27'h000000d4, 5'd28, 27'h00000394, 5'd14, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000094, 5'd26, 27'h0000011d, 5'd21, 27'h00000150, 32'h00000400,
  1'd1,  5'd27, 27'h000001f8, 5'd7, 27'h0000028d, 5'd3, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b1, 5'd8, 27'h000003dc, 5'd14, 27'h000000cf, 32'h00000400,
  1'd1,  5'd30, 27'h00000257, 5'd7, 27'h0000027c, 5'd23, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000009, 5'd19, 27'h000001af, 5'd1, 27'h000001f8, 32'h00000400,
  1'd1,  5'd28, 27'h00000354, 5'd19, 27'h000003fd, 5'd14, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000295, 5'd19, 27'h00000380, 5'd25, 27'h000001be, 32'h00000400,
  1'd1,  5'd28, 27'h0000013f, 5'd30, 27'h00000117, 5'd0, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000305, 5'd28, 27'h000001ed, 5'd10, 27'h000003fd, 32'h00000400,
  1'd1,  5'd27, 27'h00000294, 5'd29, 27'h00000021, 5'd24, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000096, 5'd8, 27'h000000f3, 5'd5, 27'h000001c5, 32'h00000400,
  1'd1,  5'd8, 27'h000002da, 5'd7, 27'h0000011d, 5'd18, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000000e, 5'd7, 27'h0000018f, 5'd28, 27'h0000011a, 32'h00000400,
  1'd1,  5'd8, 27'h00000015, 5'd19, 27'h00000018, 5'd6, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000ef, 5'd16, 27'h00000140, 5'd16, 27'h0000038a, 32'h00000400,
  1'd1,  5'd9, 27'h0000024d, 5'd17, 27'h0000035c, 5'd28, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001cf, 5'd29, 27'h000000f5, 5'd9, 27'h00000330, 32'h00000400,
  1'd1,  5'd10, 27'h00000123, 5'd30, 27'h000001d0, 5'd15, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f4, 5'd30, 27'h00000228, 5'd28, 27'h00000083, 32'h00000400,
  1'd1,  5'd16, 27'h00000296, 5'd9, 27'h00000127, 5'd6, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000012f, 5'd9, 27'h00000083, 5'd19, 27'h00000117, 32'h00000400,
  1'd1,  5'd15, 27'h000002da, 5'd8, 27'h0000036f, 5'd25, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000398, 5'd16, 27'h00000019, 5'd8, 27'h0000004e, 32'h00000400,
  1'd1,  5'd15, 27'h000002d5, 5'd18, 27'h000001f1, 5'd20, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000015f, 5'd16, 27'h0000005c, 5'd29, 27'h000003b6, 32'h00000400,
  1'd1,  5'd17, 27'h00000308, 5'd27, 27'h000001f2, 5'd6, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000008c, 5'd26, 27'h00000210, 5'd16, 27'h000001bc, 32'h00000400,
  1'd1,  5'd18, 27'h00000103, 5'd26, 27'h00000208, 5'd27, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000011b, 5'd10, 27'h00000055, 5'd9, 27'h00000220, 32'h00000400,
  1'd1,  5'd30, 27'h0000025f, 5'd6, 27'h00000315, 5'd19, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a8, 5'd10, 27'h00000093, 5'd29, 27'h000000ef, 32'h00000400,
  1'd1,  5'd28, 27'h0000031b, 5'd18, 27'h00000341, 5'd5, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003ce, 5'd17, 27'h00000293, 5'd20, 27'h0000026c, 32'h00000400,
  1'd1,  5'd27, 27'h000002b4, 5'd20, 27'h00000078, 5'd26, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000302, 5'd30, 27'h0000014e, 5'd9, 27'h0000038f, 32'h00000400,
  1'd1,  5'd27, 27'h000000bc, 5'd27, 27'h0000026d, 5'd17, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ef, 5'd29, 27'h000003f6, 5'd29, 27'h00000379, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000293, 5'd4, 27'h000000b3, 5'd3, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000055, 5'd2, 27'h000001d5, 5'd12, 27'h00000344, 32'h00000400,
  1'd1,  5'd2, 27'h00000389, 5'd4, 27'h000002d5, 5'd21, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000083, 5'd10, 27'h000003c1, 5'd2, 27'h00000279, 32'h00000400,
  1'd1,  5'd0, 27'h000000bf, 5'd13, 27'h00000138, 5'd15, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002b4, 5'd14, 27'h000001f1, 5'd21, 27'h00000061, 32'h00000400,
  1'd1,  5'd0, 27'h000001fd, 5'd24, 27'h0000014b, 5'd2, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000231, 5'd25, 27'h000000e5, 5'd12, 27'h000001e6, 32'h00000400,
  1'd1,  5'd3, 27'h000003f5, 5'd25, 27'h000000c8, 5'd23, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000013b, 5'd4, 27'h000001c5, 5'd2, 27'h00000068, 32'h00000400,
  1'd1,  5'd12, 27'h000001b2, 5'd1, 27'h000000e8, 5'd10, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000330, 5'd1, 27'h000002f9, 5'd21, 27'h000001bd, 32'h00000400,
  1'd1,  5'd11, 27'h00000028, 5'd11, 27'h00000224, 5'd2, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000055, 5'd13, 27'h00000217, 5'd11, 27'h00000184, 32'h00000400,
  1'd1,  5'd12, 27'h00000195, 5'd10, 27'h00000254, 5'd23, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000304, 5'd23, 27'h000001da, 5'd3, 27'h00000357, 32'h00000400,
  1'd1,  5'd14, 27'h000001ad, 5'd22, 27'h000002f2, 5'd13, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008d, 5'd22, 27'h00000220, 5'd23, 27'h00000400, 32'h00000400,
  1'd1,  5'd24, 27'h000001e6, 5'd3, 27'h0000028b, 5'd1, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a1, 5'd4, 27'h0000006a, 5'd13, 27'h0000023d, 32'h00000400,
  1'd1,  5'd22, 27'h000000a8, 5'd3, 27'h00000128, 5'd24, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001a2, 5'd15, 27'h0000018c, 5'd1, 27'h00000286, 32'h00000400,
  1'd1,  5'd21, 27'h00000077, 5'd13, 27'h000000ac, 5'd11, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e4, 5'd13, 27'h000000fe, 5'd23, 27'h00000032, 32'h00000400,
  1'd1,  5'd25, 27'h000001d8, 5'd22, 27'h000003bb, 5'd2, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000038e, 5'd25, 27'h00000279, 5'd10, 27'h0000039a, 32'h00000400,
  1'd1,  5'd25, 27'h000000ff, 5'd24, 27'h0000022c, 5'd24, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f6, 5'd2, 27'h00000284, 5'd8, 27'h000001e2, 32'h00000400,
  1'd1,  5'd2, 27'h00000201, 5'd3, 27'h000000a5, 5'd19, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000020e, 5'd4, 27'h00000090, 5'd30, 27'h00000360, 32'h00000400,
  1'd1,  5'd4, 27'h00000223, 5'd13, 27'h0000025e, 5'd7, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000113, 5'd14, 27'h00000380, 5'd15, 27'h0000027d, 32'h00000400,
  1'd1,  5'd0, 27'h000003db, 5'd11, 27'h00000205, 5'd28, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f4, 5'd22, 27'h000002b0, 5'd8, 27'h000002fe, 32'h00000400,
  1'd1,  5'd2, 27'h000001a2, 5'd24, 27'h000003f5, 5'd20, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000035e, 5'd23, 27'h000001e2, 5'd30, 27'h00000092, 32'h00000400,
  1'd1,  5'd11, 27'h000001a6, 5'd1, 27'h00000079, 5'd8, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d4, 5'd0, 27'h00000250, 5'd16, 27'h0000011e, 32'h00000400,
  1'd1,  5'd11, 27'h00000084, 5'd4, 27'h000003c6, 5'd29, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000b5, 5'd11, 27'h00000258, 5'd6, 27'h0000001f, 32'h00000400,
  1'd1,  5'd10, 27'h00000224, 5'd11, 27'h00000067, 5'd16, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003f9, 5'd14, 27'h00000044, 5'd26, 27'h00000222, 32'h00000400,
  1'd1,  5'd14, 27'h000000db, 5'd22, 27'h0000027e, 5'd8, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000039b, 5'd21, 27'h000002e9, 5'd19, 27'h000003c5, 32'h00000400,
  1'd1,  5'd14, 27'h00000310, 5'd20, 27'h00000375, 5'd29, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000026c, 5'd4, 27'h00000344, 5'd6, 27'h000001ac, 32'h00000400,
  1'd1,  5'd22, 27'h0000012d, 5'd5, 27'h00000017, 5'd17, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000134, 5'd4, 27'h00000367, 5'd29, 27'h000000d3, 32'h00000400,
  1'd1,  5'd23, 27'h00000330, 5'd15, 27'h0000008e, 5'd8, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000006c, 5'd11, 27'h000002ed, 5'd20, 27'h0000002e, 32'h00000400,
  1'd1,  5'd22, 27'h000000b0, 5'd13, 27'h0000025d, 5'd27, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000033a, 5'd23, 27'h000001db, 5'd9, 27'h00000078, 32'h00000400,
  1'd1,  5'd23, 27'h000000ca, 5'd24, 27'h00000215, 5'd18, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000094, 5'd21, 27'h0000035a, 5'd25, 27'h000003a6, 32'h00000400,
  1'd1,  5'd2, 27'h000001d2, 5'd9, 27'h00000128, 5'd2, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000af, 5'd6, 27'h00000269, 5'd11, 27'h000000f8, 32'h00000400,
  1'd1,  5'd4, 27'h00000388, 5'd6, 27'h000003c0, 5'd24, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000249, 5'd17, 27'h0000010b, 5'd5, 27'h000000a1, 32'h00000400,
  1'd1,  5'd3, 27'h00000189, 5'd16, 27'h00000081, 5'd11, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000336, 5'd15, 27'h00000203, 5'd24, 27'h0000017a, 32'h00000400,
  1'd1,  5'd3, 27'h0000000a, 5'd26, 27'h00000027, 5'd0, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ed, 5'd28, 27'h0000012b, 5'd12, 27'h000001cc, 32'h00000400,
  1'd1,  5'd2, 27'h0000033f, 5'd27, 27'h00000026, 5'd22, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000036f, 5'd9, 27'h000003bc, 5'd1, 27'h000000b1, 32'h00000400,
  1'd1,  5'd11, 27'h00000323, 5'd7, 27'h000001b1, 5'd15, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003d8, 5'd9, 27'h000000f7, 5'd22, 27'h0000005c, 32'h00000400,
  1'd1,  5'd15, 27'h000000ae, 5'd19, 27'h000001d4, 5'd1, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000060, 5'd20, 27'h0000021a, 5'd11, 27'h0000025f, 32'h00000400,
  1'd1,  5'd13, 27'h000003ae, 5'd19, 27'h0000021e, 5'd24, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000034b, 5'd29, 27'h000001b4, 5'd3, 27'h00000225, 32'h00000400,
  1'd1,  5'd13, 27'h000003c3, 5'd26, 27'h00000277, 5'd11, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000339, 5'd26, 27'h00000181, 5'd22, 27'h000000e4, 32'h00000400,
  1'd1,  5'd23, 27'h00000354, 5'd6, 27'h000002bd, 5'd4, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000030f, 5'd6, 27'h0000023e, 5'd14, 27'h0000038a, 32'h00000400,
  1'd1,  5'd24, 27'h000000dd, 5'd9, 27'h0000014f, 5'd24, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000294, 5'd17, 27'h00000384, 5'd0, 27'h000000eb, 32'h00000400,
  1'd1,  5'd25, 27'h0000009d, 5'd20, 27'h00000253, 5'd13, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000363, 5'd16, 27'h000003d3, 5'd21, 27'h0000030a, 32'h00000400,
  1'd1,  5'd25, 27'h00000316, 5'd30, 27'h000001d9, 5'd4, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000009a, 5'd28, 27'h000003b5, 5'd11, 27'h00000177, 32'h00000400,
  1'd1,  5'd20, 27'h000002ea, 5'd27, 27'h000000f5, 5'd24, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003ad, 5'd9, 27'h0000014c, 5'd9, 27'h000003b9, 32'h00000400,
  1'd1,  5'd3, 27'h00000108, 5'd5, 27'h0000013e, 5'd19, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000aa, 5'd9, 27'h00000055, 5'd29, 27'h00000034, 32'h00000400,
  1'd1,  5'd0, 27'h00000262, 5'd18, 27'h00000269, 5'd6, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000aa, 5'd18, 27'h00000276, 5'd16, 27'h000002a3, 32'h00000400,
  1'd1,  5'd2, 27'h00000317, 5'd20, 27'h0000012f, 5'd28, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000011b, 5'd30, 27'h00000133, 5'd7, 27'h000003ca, 32'h00000400,
  1'd1,  5'd0, 27'h0000021a, 5'd29, 27'h00000009, 5'd18, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000345, 5'd29, 27'h0000006b, 5'd29, 27'h00000037, 32'h00000400,
  1'd1,  5'd14, 27'h00000118, 5'd6, 27'h00000061, 5'd10, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f7, 5'd9, 27'h0000032d, 5'd16, 27'h0000008d, 32'h00000400,
  1'd1,  5'd11, 27'h000001ca, 5'd9, 27'h00000337, 5'd26, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b4, 5'd16, 27'h000002ca, 5'd6, 27'h000000f2, 32'h00000400,
  1'd1,  5'd14, 27'h0000007a, 5'd20, 27'h000002a7, 5'd17, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001c7, 5'd15, 27'h000003f2, 5'd28, 27'h00000037, 32'h00000400,
  1'd1,  5'd13, 27'h0000003f, 5'd30, 27'h00000341, 5'd10, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000000c, 5'd29, 27'h00000337, 5'd17, 27'h0000018c, 32'h00000400,
  1'd1,  5'd13, 27'h000000ed, 5'd30, 27'h000003be, 5'd27, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000014, 5'd8, 27'h00000007, 5'd8, 27'h00000146, 32'h00000400,
  1'd1,  5'd24, 27'h00000039, 5'd9, 27'h000001cc, 5'd15, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003f7, 5'd8, 27'h000000d7, 5'd26, 27'h0000027f, 32'h00000400,
  1'd1,  5'd25, 27'h00000030, 5'd15, 27'h000002ca, 5'd6, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000003a, 5'd15, 27'h00000225, 5'd17, 27'h00000251, 32'h00000400,
  1'd1,  5'd21, 27'h000002a6, 5'd17, 27'h00000085, 5'd27, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a9, 5'd28, 27'h00000171, 5'd9, 27'h00000295, 32'h00000400,
  1'd1,  5'd23, 27'h00000120, 5'd27, 27'h00000374, 5'd18, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000018c, 5'd27, 27'h00000285, 5'd26, 27'h0000029a, 32'h00000400,
  1'd1,  5'd5, 27'h0000035c, 5'd1, 27'h0000026c, 5'd8, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001fb, 5'd3, 27'h000001f0, 5'd19, 27'h000003a7, 32'h00000400,
  1'd1,  5'd9, 27'h000000d3, 5'd2, 27'h0000039f, 5'd28, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000209, 5'd11, 27'h0000038e, 5'd1, 27'h00000058, 32'h00000400,
  1'd1,  5'd5, 27'h0000024d, 5'd14, 27'h000001dc, 5'd13, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003bf, 5'd13, 27'h00000156, 5'd20, 27'h00000354, 32'h00000400,
  1'd1,  5'd9, 27'h00000104, 5'd22, 27'h000000e6, 5'd1, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000396, 5'd21, 27'h000001e9, 5'd14, 27'h000001e2, 32'h00000400,
  1'd1,  5'd8, 27'h000000cf, 5'd20, 27'h0000036c, 5'd24, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c0, 5'd2, 27'h0000019c, 5'd9, 27'h00000325, 32'h00000400,
  1'd1,  5'd18, 27'h00000128, 5'd1, 27'h000000b6, 5'd18, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000189, 5'd1, 27'h0000035f, 5'd28, 27'h00000053, 32'h00000400,
  1'd1,  5'd19, 27'h00000395, 5'd11, 27'h0000020e, 5'd2, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b4, 5'd14, 27'h00000234, 5'd13, 27'h00000271, 32'h00000400,
  1'd1,  5'd16, 27'h0000007f, 5'd12, 27'h000002ed, 5'd22, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000112, 5'd24, 27'h000002f7, 5'd1, 27'h000002ae, 32'h00000400,
  1'd1,  5'd16, 27'h000000a0, 5'd21, 27'h00000251, 5'd10, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000020, 5'd21, 27'h0000009b, 5'd25, 27'h00000319, 32'h00000400,
  1'd1,  5'd26, 27'h00000371, 5'd4, 27'h000001d2, 5'd2, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000ce, 5'd0, 27'h00000164, 5'd14, 27'h00000015, 32'h00000400,
  1'd1,  5'd26, 27'h00000392, 5'd3, 27'h00000258, 5'd23, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002a0, 5'd10, 27'h000002f0, 5'd0, 27'h000002b6, 32'h00000400,
  1'd1,  5'd27, 27'h00000388, 5'd10, 27'h000002af, 5'd12, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002d4, 5'd14, 27'h0000031a, 5'd24, 27'h00000369, 32'h00000400,
  1'd1,  5'd26, 27'h00000054, 5'd20, 27'h000003f0, 5'd4, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e1, 5'd23, 27'h00000238, 5'd10, 27'h000003f2, 32'h00000400,
  1'd1,  5'd29, 27'h00000325, 5'd25, 27'h00000185, 5'd22, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000205, 5'd2, 27'h00000238, 5'd3, 27'h0000026b, 32'h00000400,
  1'd1,  5'd7, 27'h000003dd, 5'd3, 27'h00000309, 5'd11, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003df, 5'd3, 27'h00000079, 5'd21, 27'h000002f5, 32'h00000400,
  1'd1,  5'd6, 27'h000001a0, 5'd13, 27'h000002ab, 5'd5, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000209, 5'd15, 27'h00000140, 5'd15, 27'h00000362, 32'h00000400,
  1'd1,  5'd5, 27'h0000035d, 5'd13, 27'h00000362, 5'd28, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ac, 5'd20, 27'h000002e7, 5'd6, 27'h00000364, 32'h00000400,
  1'd1,  5'd5, 27'h000001c6, 5'd22, 27'h00000018, 5'd17, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000128, 5'd25, 27'h000002f1, 5'd29, 27'h000003d5, 32'h00000400,
  1'd1,  5'd16, 27'h000000fd, 5'd4, 27'h0000020f, 5'd2, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ca, 5'd3, 27'h000001bf, 5'd13, 27'h000002a6, 32'h00000400,
  1'd1,  5'd17, 27'h00000341, 5'd2, 27'h0000035e, 5'd22, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000061, 5'd14, 27'h000003cc, 5'd9, 27'h0000027b, 32'h00000400,
  1'd1,  5'd15, 27'h0000026b, 5'd11, 27'h000003f0, 5'd16, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b2, 5'd11, 27'h00000062, 5'd30, 27'h00000090, 32'h00000400,
  1'd1,  5'd20, 27'h00000207, 5'd22, 27'h000001b0, 5'd6, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000390, 5'd25, 27'h000001c4, 5'd16, 27'h0000026d, 32'h00000400,
  1'd1,  5'd16, 27'h000003cd, 5'd20, 27'h000003b3, 5'd30, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000195, 5'd4, 27'h0000009a, 5'd7, 27'h000002ac, 32'h00000400,
  1'd1,  5'd26, 27'h000003e6, 5'd1, 27'h0000031a, 5'd15, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000373, 5'd2, 27'h00000044, 5'd28, 27'h00000238, 32'h00000400,
  1'd1,  5'd29, 27'h00000204, 5'd11, 27'h000002fa, 5'd10, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000240, 5'd12, 27'h0000018b, 5'd17, 27'h00000054, 32'h00000400,
  1'd1,  5'd30, 27'h00000221, 5'd11, 27'h000003a6, 5'd30, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000da, 5'd21, 27'h0000015e, 5'd5, 27'h000002df, 32'h00000400,
  1'd1,  5'd27, 27'h000003e2, 5'd21, 27'h000002b0, 5'd17, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000012e, 5'd20, 27'h00000388, 5'd27, 27'h00000296, 32'h00000400,
  1'd1,  5'd7, 27'h000000db, 5'd9, 27'h0000013a, 5'd4, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000187, 5'd6, 27'h00000313, 5'd14, 27'h0000010a, 32'h00000400,
  1'd1,  5'd5, 27'h000002f5, 5'd7, 27'h0000026f, 5'd22, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e9, 5'd16, 27'h00000038, 5'd0, 27'h00000110, 32'h00000400,
  1'd1,  5'd9, 27'h000002a2, 5'd20, 27'h000002a6, 5'd14, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000200, 5'd16, 27'h00000313, 5'd24, 27'h00000291, 32'h00000400,
  1'd1,  5'd7, 27'h00000218, 5'd30, 27'h000001fb, 5'd1, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000032b, 5'd27, 27'h0000037f, 5'd15, 27'h000000c5, 32'h00000400,
  1'd1,  5'd9, 27'h0000028c, 5'd30, 27'h000001cf, 5'd25, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000b7, 5'd6, 27'h00000169, 5'd1, 27'h000003b9, 32'h00000400,
  1'd1,  5'd16, 27'h0000007a, 5'd8, 27'h000003c7, 5'd12, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000022b, 5'd8, 27'h00000131, 5'd20, 27'h00000316, 32'h00000400,
  1'd1,  5'd16, 27'h00000100, 5'd18, 27'h0000010c, 5'd5, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ec, 5'd17, 27'h000001d1, 5'd12, 27'h00000102, 32'h00000400,
  1'd1,  5'd19, 27'h000000fd, 5'd17, 27'h00000334, 5'd23, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000f5, 5'd28, 27'h000001fd, 5'd3, 27'h00000012, 32'h00000400,
  1'd1,  5'd19, 27'h000003eb, 5'd26, 27'h000003e6, 5'd11, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000330, 5'd30, 27'h000003e3, 5'd25, 27'h000000ef, 32'h00000400,
  1'd1,  5'd29, 27'h000003b4, 5'd5, 27'h0000038a, 5'd2, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000330, 5'd7, 27'h000003c4, 5'd12, 27'h00000015, 32'h00000400,
  1'd1,  5'd28, 27'h00000108, 5'd5, 27'h0000030b, 5'd23, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003b2, 5'd18, 27'h00000290, 5'd4, 27'h000001de, 32'h00000400,
  1'd1,  5'd26, 27'h00000075, 5'd18, 27'h0000012f, 5'd14, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000213, 5'd20, 27'h00000167, 5'd24, 27'h00000303, 32'h00000400,
  1'd1,  5'd28, 27'h000003c6, 5'd30, 27'h000002fe, 5'd0, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001dd, 5'd28, 27'h000002ae, 5'd12, 27'h0000015d, 32'h00000400,
  1'd1,  5'd27, 27'h000002af, 5'd25, 27'h0000039d, 5'd25, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e4, 5'd9, 27'h00000143, 5'd5, 27'h000001fb, 32'h00000400,
  1'd1,  5'd6, 27'h0000015e, 5'd9, 27'h000002b5, 5'd17, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ab, 5'd9, 27'h00000273, 5'd30, 27'h0000039a, 32'h00000400,
  1'd1,  5'd10, 27'h0000008d, 5'd17, 27'h00000029, 5'd7, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000008f, 5'd18, 27'h000000a2, 5'd19, 27'h00000400, 32'h00000400,
  1'd1,  5'd9, 27'h00000262, 5'd18, 27'h000003cd, 5'd30, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034c, 5'd28, 27'h000000dd, 5'd6, 27'h000003cd, 32'h00000400,
  1'd1,  5'd8, 27'h00000210, 5'd29, 27'h000002b8, 5'd18, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000004f, 5'd26, 27'h00000088, 5'd28, 27'h000000b6, 32'h00000400,
  1'd1,  5'd17, 27'h00000316, 5'd8, 27'h00000060, 5'd7, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000281, 5'd6, 27'h000001b7, 5'd16, 27'h000000d4, 32'h00000400,
  1'd1,  5'd19, 27'h0000010b, 5'd6, 27'h00000294, 5'd27, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002a4, 5'd19, 27'h00000056, 5'd8, 27'h000000af, 32'h00000400,
  1'd1,  5'd20, 27'h0000011b, 5'd19, 27'h00000360, 5'd17, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000130, 5'd15, 27'h00000319, 5'd26, 27'h000002a8, 32'h00000400,
  1'd1,  5'd15, 27'h000002c6, 5'd26, 27'h00000396, 5'd9, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000008d, 5'd28, 27'h0000033b, 5'd15, 27'h000002cb, 32'h00000400,
  1'd1,  5'd18, 27'h00000111, 5'd26, 27'h00000310, 5'd29, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d6, 5'd9, 27'h00000072, 5'd6, 27'h000002b2, 32'h00000400,
  1'd1,  5'd26, 27'h0000009d, 5'd6, 27'h0000005d, 5'd16, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000175, 5'd8, 27'h000003f1, 5'd29, 27'h00000360, 32'h00000400,
  1'd1,  5'd26, 27'h00000327, 5'd18, 27'h00000071, 5'd5, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d1, 5'd15, 27'h000002b7, 5'd15, 27'h000003cc, 32'h00000400,
  1'd1,  5'd29, 27'h000003e9, 5'd16, 27'h00000340, 5'd29, 27'h000001e2, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000259, 5'd26, 27'h0000025c, 5'd9, 27'h00000110, 32'h00000400,
  1'd1,  5'd27, 27'h000001b2, 5'd27, 27'h00000312, 5'd17, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002fa, 5'd28, 27'h00000297, 5'd29, 27'h000001da, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000004d, 5'd0, 27'h000000b1, 5'd0, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000197, 5'd2, 27'h000000ed, 5'd12, 27'h00000117, 32'h00000400,
  1'd1,  5'd3, 27'h00000082, 5'd0, 27'h0000018c, 5'd25, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000344, 5'd10, 27'h000001f1, 5'd4, 27'h0000008e, 32'h00000400,
  1'd1,  5'd5, 27'h0000002c, 5'd12, 27'h000000f3, 5'd12, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000021c, 5'd12, 27'h00000334, 5'd22, 27'h00000236, 32'h00000400,
  1'd1,  5'd0, 27'h0000000e, 5'd22, 27'h0000008b, 5'd1, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d2, 5'd22, 27'h000001d8, 5'd14, 27'h00000330, 32'h00000400,
  1'd1,  5'd3, 27'h000002d7, 5'd20, 27'h00000364, 5'd24, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000108, 5'd1, 27'h0000034c, 5'd5, 27'h00000043, 32'h00000400,
  1'd1,  5'd13, 27'h00000369, 5'd1, 27'h000003a4, 5'd12, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ab, 5'd1, 27'h0000033e, 5'd24, 27'h00000217, 32'h00000400,
  1'd1,  5'd14, 27'h00000399, 5'd15, 27'h00000099, 5'd0, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000014d, 5'd12, 27'h000003d6, 5'd11, 27'h000003c1, 32'h00000400,
  1'd1,  5'd11, 27'h000000be, 5'd11, 27'h000003d9, 5'd23, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003aa, 5'd24, 27'h00000349, 5'd4, 27'h00000038, 32'h00000400,
  1'd1,  5'd13, 27'h0000001d, 5'd25, 27'h0000010a, 5'd14, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000142, 5'd24, 27'h0000001a, 5'd25, 27'h000001ab, 32'h00000400,
  1'd1,  5'd24, 27'h00000357, 5'd4, 27'h00000003, 5'd2, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ae, 5'd1, 27'h000002d3, 5'd15, 27'h00000001, 32'h00000400,
  1'd1,  5'd24, 27'h00000105, 5'd0, 27'h000000cf, 5'd22, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e8, 5'd14, 27'h000002b3, 5'd3, 27'h00000385, 32'h00000400,
  1'd1,  5'd22, 27'h00000053, 5'd13, 27'h000003a5, 5'd14, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000004f, 5'd14, 27'h0000020e, 5'd23, 27'h000002a7, 32'h00000400,
  1'd1,  5'd23, 27'h00000395, 5'd24, 27'h000002b7, 5'd2, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000328, 5'd24, 27'h00000234, 5'd12, 27'h0000013d, 32'h00000400,
  1'd1,  5'd23, 27'h00000014, 5'd23, 27'h0000001d, 5'd24, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000346, 5'd4, 27'h000002b0, 5'd6, 27'h000002ac, 32'h00000400,
  1'd1,  5'd2, 27'h000002b5, 5'd1, 27'h00000314, 5'd19, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fc, 5'd4, 27'h00000011, 5'd30, 27'h00000051, 32'h00000400,
  1'd1,  5'd0, 27'h0000010e, 5'd13, 27'h000003c2, 5'd9, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000003b, 5'd12, 27'h000000a5, 5'd16, 27'h00000023, 32'h00000400,
  1'd1,  5'd5, 27'h0000004e, 5'd10, 27'h000003a6, 5'd25, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000001, 5'd21, 27'h000001c4, 5'd8, 27'h0000032a, 32'h00000400,
  1'd1,  5'd3, 27'h00000348, 5'd23, 27'h000001c1, 5'd18, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000007f, 5'd20, 27'h000002b2, 5'd28, 27'h0000010d, 32'h00000400,
  1'd1,  5'd10, 27'h00000314, 5'd3, 27'h00000075, 5'd9, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003f, 5'd4, 27'h00000214, 5'd20, 27'h0000007f, 32'h00000400,
  1'd1,  5'd13, 27'h00000323, 5'd1, 27'h000000b2, 5'd28, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000016f, 5'd12, 27'h0000016c, 5'd9, 27'h0000038b, 32'h00000400,
  1'd1,  5'd12, 27'h0000004c, 5'd12, 27'h00000007, 5'd16, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000148, 5'd14, 27'h00000038, 5'd30, 27'h000000eb, 32'h00000400,
  1'd1,  5'd14, 27'h00000016, 5'd21, 27'h0000033b, 5'd9, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000352, 5'd25, 27'h00000119, 5'd16, 27'h0000005c, 32'h00000400,
  1'd1,  5'd12, 27'h0000021b, 5'd21, 27'h000000de, 5'd27, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000023c, 5'd2, 27'h0000023b, 5'd6, 27'h0000003a, 32'h00000400,
  1'd1,  5'd24, 27'h000001d4, 5'd5, 27'h000000a3, 5'd17, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003d0, 5'd2, 27'h00000189, 5'd30, 27'h00000078, 32'h00000400,
  1'd1,  5'd21, 27'h000002ff, 5'd13, 27'h00000235, 5'd5, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000228, 5'd12, 27'h00000114, 5'd18, 27'h000002c7, 32'h00000400,
  1'd1,  5'd24, 27'h0000035a, 5'd14, 27'h0000009a, 5'd26, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000024a, 5'd23, 27'h00000278, 5'd6, 27'h000001d7, 32'h00000400,
  1'd1,  5'd22, 27'h000001a9, 5'd21, 27'h000000ee, 5'd16, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000240, 5'd23, 27'h000001a1, 5'd30, 27'h0000001e, 32'h00000400,
  1'd1,  5'd2, 27'h000002db, 5'd6, 27'h000002bd, 5'd2, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000146, 5'd5, 27'h00000246, 5'd14, 27'h00000076, 32'h00000400,
  1'd1,  5'd4, 27'h00000227, 5'd7, 27'h00000186, 5'd25, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000087, 5'd17, 27'h000003ac, 5'd4, 27'h0000002f, 32'h00000400,
  1'd1,  5'd3, 27'h00000196, 5'd17, 27'h00000150, 5'd10, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f0, 5'd19, 27'h0000023a, 5'd20, 27'h000002b7, 32'h00000400,
  1'd1,  5'd1, 27'h00000345, 5'd29, 27'h00000024, 5'd1, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000036a, 5'd30, 27'h00000212, 5'd12, 27'h00000054, 32'h00000400,
  1'd1,  5'd2, 27'h00000219, 5'd29, 27'h0000015c, 5'd24, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000264, 5'd6, 27'h0000038c, 5'd5, 27'h00000042, 32'h00000400,
  1'd1,  5'd13, 27'h00000144, 5'd5, 27'h00000281, 5'd10, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000013, 5'd7, 27'h0000032f, 5'd24, 27'h00000267, 32'h00000400,
  1'd1,  5'd12, 27'h0000001e, 5'd20, 27'h00000239, 5'd2, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023b, 5'd15, 27'h0000039b, 5'd14, 27'h0000013c, 32'h00000400,
  1'd1,  5'd13, 27'h00000122, 5'd15, 27'h000003ba, 5'd21, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000047, 5'd27, 27'h00000276, 5'd3, 27'h00000173, 32'h00000400,
  1'd1,  5'd11, 27'h00000348, 5'd27, 27'h0000023c, 5'd13, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a7, 5'd28, 27'h00000377, 5'd21, 27'h000001d6, 32'h00000400,
  1'd1,  5'd23, 27'h0000017e, 5'd8, 27'h000001d0, 5'd1, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002f1, 5'd5, 27'h00000389, 5'd12, 27'h0000035c, 32'h00000400,
  1'd1,  5'd21, 27'h000000a2, 5'd7, 27'h000000dd, 5'd21, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000025, 5'd18, 27'h0000021a, 5'd2, 27'h0000038c, 32'h00000400,
  1'd1,  5'd25, 27'h00000267, 5'd15, 27'h000003c3, 5'd12, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000128, 5'd18, 27'h00000344, 5'd22, 27'h0000028b, 32'h00000400,
  1'd1,  5'd21, 27'h00000270, 5'd27, 27'h00000318, 5'd2, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000051, 5'd30, 27'h00000035, 5'd15, 27'h000000d7, 32'h00000400,
  1'd1,  5'd21, 27'h0000032f, 5'd28, 27'h00000150, 5'd23, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000157, 5'd5, 27'h0000036f, 5'd6, 27'h00000168, 32'h00000400,
  1'd1,  5'd0, 27'h00000338, 5'd6, 27'h00000056, 5'd19, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000020c, 5'd5, 27'h000000ad, 5'd27, 27'h000001fa, 32'h00000400,
  1'd1,  5'd3, 27'h0000028d, 5'd17, 27'h0000011e, 5'd6, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000387, 5'd15, 27'h00000345, 5'd15, 27'h000003c9, 32'h00000400,
  1'd1,  5'd3, 27'h0000018f, 5'd18, 27'h00000104, 5'd26, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002a5, 5'd27, 27'h000001eb, 5'd9, 27'h000000ca, 32'h00000400,
  1'd1,  5'd4, 27'h000003e4, 5'd28, 27'h0000013d, 5'd15, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001d2, 5'd26, 27'h00000165, 5'd28, 27'h000002ef, 32'h00000400,
  1'd1,  5'd13, 27'h0000029c, 5'd7, 27'h00000096, 5'd10, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000037f, 5'd10, 27'h0000000f, 5'd16, 27'h00000164, 32'h00000400,
  1'd1,  5'd13, 27'h00000242, 5'd6, 27'h00000118, 5'd26, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000051, 5'd15, 27'h00000308, 5'd8, 27'h000000c6, 32'h00000400,
  1'd1,  5'd12, 27'h0000034b, 5'd15, 27'h00000251, 5'd20, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000031d, 5'd16, 27'h000000b7, 5'd26, 27'h0000037d, 32'h00000400,
  1'd1,  5'd12, 27'h0000019b, 5'd30, 27'h0000030a, 5'd9, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f3, 5'd27, 27'h000003ca, 5'd15, 27'h00000249, 32'h00000400,
  1'd1,  5'd13, 27'h00000199, 5'd26, 27'h000002b2, 5'd29, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000002b, 5'd8, 27'h000002fc, 5'd10, 27'h000000e5, 32'h00000400,
  1'd1,  5'd21, 27'h00000058, 5'd8, 27'h00000391, 5'd16, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003af, 5'd5, 27'h000002c6, 5'd29, 27'h00000267, 32'h00000400,
  1'd1,  5'd22, 27'h000002cd, 5'd16, 27'h000001cf, 5'd8, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000145, 5'd17, 27'h00000399, 5'd18, 27'h0000020a, 32'h00000400,
  1'd1,  5'd22, 27'h000000e4, 5'd18, 27'h0000014c, 5'd28, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001e0, 5'd27, 27'h0000004a, 5'd10, 27'h00000010, 32'h00000400,
  1'd1,  5'd25, 27'h0000033f, 5'd29, 27'h00000124, 5'd17, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000129, 5'd29, 27'h0000029b, 5'd28, 27'h000003d7, 32'h00000400,
  1'd1,  5'd8, 27'h00000276, 5'd4, 27'h000002f5, 5'd5, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c2, 5'd3, 27'h00000012, 5'd16, 27'h000003ed, 32'h00000400,
  1'd1,  5'd5, 27'h00000392, 5'd2, 27'h00000094, 5'd25, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002b4, 5'd14, 27'h00000048, 5'd1, 27'h0000030c, 32'h00000400,
  1'd1,  5'd8, 27'h000001b7, 5'd14, 27'h00000372, 5'd10, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000010f, 5'd12, 27'h00000060, 5'd22, 27'h00000072, 32'h00000400,
  1'd1,  5'd5, 27'h00000382, 5'd20, 27'h00000344, 5'd3, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000160, 5'd22, 27'h00000375, 5'd15, 27'h000001eb, 32'h00000400,
  1'd1,  5'd10, 27'h0000013b, 5'd22, 27'h00000394, 5'd23, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000219, 5'd0, 27'h00000198, 5'd8, 27'h00000173, 32'h00000400,
  1'd1,  5'd15, 27'h0000038b, 5'd2, 27'h00000154, 5'd17, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000169, 5'd5, 27'h00000082, 5'd29, 27'h000001f3, 32'h00000400,
  1'd1,  5'd19, 27'h00000225, 5'd11, 27'h00000051, 5'd1, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000232, 5'd14, 27'h0000021b, 5'd14, 27'h000003e3, 32'h00000400,
  1'd1,  5'd19, 27'h00000106, 5'd14, 27'h0000021b, 5'd24, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000017c, 5'd23, 27'h00000073, 5'd3, 27'h000000da, 32'h00000400,
  1'd1,  5'd16, 27'h00000043, 5'd21, 27'h0000001e, 5'd11, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009c, 5'd21, 27'h00000138, 5'd22, 27'h00000127, 32'h00000400,
  1'd1,  5'd29, 27'h00000051, 5'd3, 27'h000003f8, 5'd2, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000028a, 5'd0, 27'h00000378, 5'd12, 27'h00000206, 32'h00000400,
  1'd1,  5'd27, 27'h00000049, 5'd2, 27'h000003ea, 5'd25, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000211, 5'd11, 27'h0000036c, 5'd2, 27'h0000039d, 32'h00000400,
  1'd1,  5'd29, 27'h00000313, 5'd12, 27'h000000d0, 5'd14, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003f0, 5'd15, 27'h00000145, 5'd21, 27'h00000332, 32'h00000400,
  1'd1,  5'd26, 27'h000001ea, 5'd22, 27'h00000233, 5'd2, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a8, 5'd24, 27'h0000028c, 5'd12, 27'h000000ba, 32'h00000400,
  1'd1,  5'd29, 27'h000000c0, 5'd22, 27'h0000003f, 5'd24, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000001b, 5'd2, 27'h0000030d, 5'd1, 27'h000000f1, 32'h00000400,
  1'd1,  5'd6, 27'h00000363, 5'd1, 27'h000002b9, 5'd13, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000211, 5'd5, 27'h00000076, 5'd23, 27'h000001be, 32'h00000400,
  1'd1,  5'd8, 27'h0000004b, 5'd14, 27'h000000dd, 5'd6, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000040, 5'd14, 27'h000000bc, 5'd18, 27'h00000336, 32'h00000400,
  1'd1,  5'd10, 27'h000000cc, 5'd11, 27'h0000016a, 5'd27, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e2, 5'd23, 27'h000002a5, 5'd9, 27'h0000021e, 32'h00000400,
  1'd1,  5'd8, 27'h000003ad, 5'd21, 27'h000002ff, 5'd18, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000037c, 5'd21, 27'h0000000e, 5'd30, 27'h000001e2, 32'h00000400,
  1'd1,  5'd16, 27'h0000007a, 5'd1, 27'h0000021b, 5'd0, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000fa, 5'd4, 27'h00000008, 5'd13, 27'h00000105, 32'h00000400,
  1'd1,  5'd15, 27'h00000374, 5'd4, 27'h000001f8, 5'd22, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000114, 5'd10, 27'h0000025d, 5'd6, 27'h0000032d, 32'h00000400,
  1'd1,  5'd20, 27'h000001f7, 5'd14, 27'h00000128, 5'd15, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000172, 5'd14, 27'h00000217, 5'd29, 27'h000003a6, 32'h00000400,
  1'd1,  5'd17, 27'h0000004a, 5'd21, 27'h000002ef, 5'd5, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002cb, 5'd24, 27'h000001d6, 5'd16, 27'h000000cd, 32'h00000400,
  1'd1,  5'd18, 27'h000000c0, 5'd20, 27'h0000037b, 5'd28, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000064, 5'd0, 27'h00000034, 5'd6, 27'h00000014, 32'h00000400,
  1'd1,  5'd28, 27'h00000131, 5'd1, 27'h00000259, 5'd15, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000036b, 5'd0, 27'h000000a9, 5'd29, 27'h0000005a, 32'h00000400,
  1'd1,  5'd28, 27'h000001d5, 5'd14, 27'h000002ed, 5'd7, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002c3, 5'd11, 27'h0000029c, 5'd15, 27'h00000259, 32'h00000400,
  1'd1,  5'd26, 27'h000001c0, 5'd10, 27'h00000388, 5'd27, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000128, 5'd20, 27'h00000309, 5'd9, 27'h0000008e, 32'h00000400,
  1'd1,  5'd28, 27'h00000215, 5'd20, 27'h00000322, 5'd15, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000053, 5'd22, 27'h0000037a, 5'd27, 27'h00000159, 32'h00000400,
  1'd1,  5'd5, 27'h0000018e, 5'd6, 27'h000000d3, 5'd0, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000186, 5'd8, 27'h000002d1, 5'd12, 27'h000002f5, 32'h00000400,
  1'd1,  5'd8, 27'h00000262, 5'd6, 27'h00000061, 5'd21, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000033f, 5'd17, 27'h00000053, 5'd4, 27'h0000004e, 32'h00000400,
  1'd1,  5'd7, 27'h000000e6, 5'd17, 27'h00000353, 5'd10, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000057, 5'd20, 27'h0000025b, 5'd23, 27'h000003c6, 32'h00000400,
  1'd1,  5'd8, 27'h00000367, 5'd30, 27'h00000020, 5'd2, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002fb, 5'd30, 27'h000000ea, 5'd14, 27'h00000347, 32'h00000400,
  1'd1,  5'd8, 27'h0000022f, 5'd26, 27'h00000042, 5'd25, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000016c, 5'd9, 27'h000003a9, 5'd5, 27'h00000037, 32'h00000400,
  1'd1,  5'd18, 27'h000002a1, 5'd6, 27'h000001fe, 5'd11, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000187, 5'd8, 27'h000002dd, 5'd25, 27'h000001d2, 32'h00000400,
  1'd1,  5'd20, 27'h00000036, 5'd19, 27'h00000088, 5'd4, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000349, 5'd17, 27'h000000c1, 5'd11, 27'h0000014c, 32'h00000400,
  1'd1,  5'd16, 27'h000002d6, 5'd19, 27'h000002b3, 5'd23, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e7, 5'd30, 27'h000001c0, 5'd3, 27'h0000011b, 32'h00000400,
  1'd1,  5'd19, 27'h000001cf, 5'd29, 27'h000002c6, 5'd13, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000257, 5'd29, 27'h000000b8, 5'd23, 27'h00000320, 32'h00000400,
  1'd1,  5'd25, 27'h000003c7, 5'd7, 27'h0000018a, 5'd3, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000099, 5'd9, 27'h000003e4, 5'd12, 27'h00000364, 32'h00000400,
  1'd1,  5'd26, 27'h000000ad, 5'd7, 27'h0000001c, 5'd23, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000029a, 5'd17, 27'h00000182, 5'd3, 27'h000002c7, 32'h00000400,
  1'd1,  5'd26, 27'h00000319, 5'd19, 27'h000000cf, 5'd13, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000251, 5'd17, 27'h000001ca, 5'd24, 27'h00000150, 32'h00000400,
  1'd1,  5'd25, 27'h000003ba, 5'd28, 27'h00000110, 5'd5, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000006d, 5'd27, 27'h00000280, 5'd10, 27'h0000018a, 32'h00000400,
  1'd1,  5'd28, 27'h000001f2, 5'd30, 27'h000001c9, 5'd22, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000322, 5'd7, 27'h0000017a, 5'd5, 27'h000001cc, 32'h00000400,
  1'd1,  5'd8, 27'h0000016c, 5'd6, 27'h00000008, 5'd17, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000137, 5'd9, 27'h00000267, 5'd27, 27'h00000057, 32'h00000400,
  1'd1,  5'd6, 27'h00000130, 5'd18, 27'h00000277, 5'd7, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000004d, 5'd19, 27'h00000245, 5'd18, 27'h000001db, 32'h00000400,
  1'd1,  5'd8, 27'h00000045, 5'd17, 27'h00000039, 5'd29, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000124, 5'd30, 27'h000000de, 5'd6, 27'h0000037e, 32'h00000400,
  1'd1,  5'd9, 27'h00000206, 5'd26, 27'h00000369, 5'd16, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000104, 5'd30, 27'h0000031a, 5'd28, 27'h000002a9, 32'h00000400,
  1'd1,  5'd20, 27'h00000007, 5'd8, 27'h0000034b, 5'd5, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000026a, 5'd5, 27'h0000011d, 5'd18, 27'h000002f0, 32'h00000400,
  1'd1,  5'd18, 27'h000001e8, 5'd6, 27'h000002e8, 5'd29, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002cc, 5'd19, 27'h000001ea, 5'd9, 27'h0000006e, 32'h00000400,
  1'd1,  5'd18, 27'h000001af, 5'd18, 27'h0000003c, 5'd16, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000003d, 5'd20, 27'h000000b6, 5'd26, 27'h000003ba, 32'h00000400,
  1'd1,  5'd19, 27'h000000d9, 5'd29, 27'h0000029d, 5'd7, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000038d, 5'd26, 27'h000000c4, 5'd15, 27'h00000314, 32'h00000400,
  1'd1,  5'd15, 27'h000003dc, 5'd29, 27'h00000378, 5'd27, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000018d, 5'd8, 27'h00000372, 5'd9, 27'h000002c0, 32'h00000400,
  1'd1,  5'd27, 27'h00000399, 5'd10, 27'h0000012a, 5'd19, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000241, 5'd9, 27'h000003d0, 5'd30, 27'h0000021e, 32'h00000400,
  1'd1,  5'd30, 27'h000003bb, 5'd16, 27'h00000367, 5'd6, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000008a, 5'd17, 27'h00000090, 5'd17, 27'h000001e3, 32'h00000400,
  1'd1,  5'd30, 27'h00000122, 5'd18, 27'h000002b0, 5'd27, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000036d, 5'd27, 27'h00000370, 5'd9, 27'h00000293, 32'h00000400,
  1'd1,  5'd26, 27'h0000009a, 5'd27, 27'h000003dc, 5'd17, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000dd, 5'd27, 27'h0000038c, 5'd30, 27'h000001b1, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000058, 5'd0, 27'h000000d5, 5'd1, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000038a, 5'd1, 27'h0000031a, 5'd15, 27'h0000000b, 32'h00000400,
  1'd1,  5'd1, 27'h0000003f, 5'd5, 27'h00000002, 5'd24, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000186, 5'd14, 27'h000002a4, 5'd3, 27'h0000011d, 32'h00000400,
  1'd1,  5'd0, 27'h0000005c, 5'd13, 27'h00000080, 5'd10, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000dc, 5'd13, 27'h00000209, 5'd24, 27'h00000017, 32'h00000400,
  1'd1,  5'd0, 27'h0000033b, 5'd22, 27'h0000035b, 5'd1, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000002a, 5'd21, 27'h000001af, 5'd13, 27'h00000305, 32'h00000400,
  1'd1,  5'd1, 27'h00000157, 5'd22, 27'h0000031d, 5'd24, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000004e, 5'd1, 27'h000002ae, 5'd0, 27'h0000015d, 32'h00000400,
  1'd1,  5'd11, 27'h000003f2, 5'd2, 27'h000000ad, 5'd14, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000206, 5'd1, 27'h0000001f, 5'd24, 27'h000000d6, 32'h00000400,
  1'd1,  5'd13, 27'h000000b2, 5'd14, 27'h000000b4, 5'd0, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000db, 5'd11, 27'h00000187, 5'd11, 27'h00000329, 32'h00000400,
  1'd1,  5'd15, 27'h000000e7, 5'd13, 27'h00000212, 5'd22, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000029, 5'd21, 27'h0000013c, 5'd3, 27'h00000230, 32'h00000400,
  1'd1,  5'd13, 27'h000001dd, 5'd24, 27'h00000088, 5'd12, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c7, 5'd24, 27'h0000022c, 5'd25, 27'h00000123, 32'h00000400,
  1'd1,  5'd22, 27'h00000075, 5'd4, 27'h00000248, 5'd5, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000132, 5'd3, 27'h000002f8, 5'd11, 27'h000000fc, 32'h00000400,
  1'd1,  5'd24, 27'h000002d2, 5'd1, 27'h000003cb, 5'd23, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000006, 5'd12, 27'h000000c0, 5'd1, 27'h000000e9, 32'h00000400,
  1'd1,  5'd22, 27'h00000359, 5'd14, 27'h0000035d, 5'd13, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000231, 5'd12, 27'h00000309, 5'd23, 27'h00000263, 32'h00000400,
  1'd1,  5'd22, 27'h0000038c, 5'd25, 27'h00000315, 5'd2, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000122, 5'd23, 27'h00000096, 5'd11, 27'h00000382, 32'h00000400,
  1'd1,  5'd22, 27'h0000014c, 5'd21, 27'h000003b9, 5'd23, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d9, 5'd2, 27'h000001bd, 5'd8, 27'h00000059, 32'h00000400,
  1'd1,  5'd1, 27'h0000009c, 5'd3, 27'h0000014a, 5'd19, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000009d, 5'd3, 27'h0000039a, 5'd27, 27'h000000eb, 32'h00000400,
  1'd1,  5'd2, 27'h000001d3, 5'd13, 27'h00000193, 5'd7, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000014c, 5'd15, 27'h00000013, 5'd20, 27'h000001f9, 32'h00000400,
  1'd1,  5'd2, 27'h000001c7, 5'd14, 27'h00000049, 5'd29, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000035d, 5'd23, 27'h00000348, 5'd8, 27'h000001e7, 32'h00000400,
  1'd1,  5'd4, 27'h000002a5, 5'd25, 27'h0000025a, 5'd18, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000037, 5'd21, 27'h000003f0, 5'd28, 27'h0000010f, 32'h00000400,
  1'd1,  5'd10, 27'h000003c7, 5'd5, 27'h00000008, 5'd5, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000006e, 5'd4, 27'h00000016, 5'd19, 27'h000002e4, 32'h00000400,
  1'd1,  5'd12, 27'h0000001a, 5'd2, 27'h000003db, 5'd30, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000030c, 5'd10, 27'h0000022b, 5'd9, 27'h00000223, 32'h00000400,
  1'd1,  5'd11, 27'h000001b0, 5'd11, 27'h00000315, 5'd17, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000025d, 5'd15, 27'h000001ca, 5'd28, 27'h000000ef, 32'h00000400,
  1'd1,  5'd14, 27'h0000024e, 5'd25, 27'h00000017, 5'd6, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011f, 5'd21, 27'h00000165, 5'd19, 27'h000002f8, 32'h00000400,
  1'd1,  5'd15, 27'h0000008f, 5'd20, 27'h0000037b, 5'd29, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d6, 5'd2, 27'h00000130, 5'd9, 27'h0000034e, 32'h00000400,
  1'd1,  5'd25, 27'h000001a2, 5'd2, 27'h000002c6, 5'd20, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000344, 5'd2, 27'h0000023c, 5'd29, 27'h00000398, 32'h00000400,
  1'd1,  5'd22, 27'h000000d6, 5'd15, 27'h0000013e, 5'd6, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000026a, 5'd11, 27'h00000290, 5'd16, 27'h0000030c, 32'h00000400,
  1'd1,  5'd24, 27'h000000ec, 5'd12, 27'h0000015b, 5'd25, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000090, 5'd21, 27'h000003a9, 5'd7, 27'h000000ab, 32'h00000400,
  1'd1,  5'd23, 27'h0000011e, 5'd25, 27'h0000012a, 5'd19, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e4, 5'd24, 27'h000000e5, 5'd30, 27'h0000039f, 32'h00000400,
  1'd1,  5'd0, 27'h0000034d, 5'd10, 27'h00000116, 5'd2, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f4, 5'd6, 27'h00000362, 5'd12, 27'h000001f9, 32'h00000400,
  1'd1,  5'd2, 27'h0000012c, 5'd7, 27'h00000051, 5'd21, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000367, 5'd19, 27'h000001b0, 5'd1, 27'h000001ba, 32'h00000400,
  1'd1,  5'd0, 27'h0000003a, 5'd17, 27'h000001ce, 5'd12, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000014f, 5'd18, 27'h00000223, 5'd22, 27'h0000026f, 32'h00000400,
  1'd1,  5'd4, 27'h000002f6, 5'd29, 27'h000001f9, 5'd4, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000023a, 5'd27, 27'h00000112, 5'd12, 27'h000000f1, 32'h00000400,
  1'd1,  5'd0, 27'h0000012c, 5'd26, 27'h0000007e, 5'd22, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000026a, 5'd6, 27'h0000035b, 5'd3, 27'h0000027e, 32'h00000400,
  1'd1,  5'd11, 27'h000002c4, 5'd7, 27'h00000060, 5'd13, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d3, 5'd6, 27'h0000019e, 5'd25, 27'h0000034a, 32'h00000400,
  1'd1,  5'd12, 27'h0000019f, 5'd19, 27'h000001c3, 5'd1, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d1, 5'd17, 27'h00000151, 5'd15, 27'h00000149, 32'h00000400,
  1'd1,  5'd13, 27'h000000df, 5'd19, 27'h0000029a, 5'd21, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000f2, 5'd27, 27'h0000010f, 5'd1, 27'h00000396, 32'h00000400,
  1'd1,  5'd13, 27'h000002c1, 5'd30, 27'h00000267, 5'd13, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000018c, 5'd28, 27'h00000323, 5'd22, 27'h000003ca, 32'h00000400,
  1'd1,  5'd25, 27'h000002fa, 5'd9, 27'h00000215, 5'd1, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001a1, 5'd6, 27'h00000064, 5'd12, 27'h000000a4, 32'h00000400,
  1'd1,  5'd22, 27'h0000023f, 5'd8, 27'h00000378, 5'd20, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002c5, 5'd19, 27'h00000077, 5'd4, 27'h0000008e, 32'h00000400,
  1'd1,  5'd22, 27'h00000032, 5'd17, 27'h000001d9, 5'd15, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000070, 5'd17, 27'h00000264, 5'd25, 27'h0000024a, 32'h00000400,
  1'd1,  5'd21, 27'h000001a1, 5'd29, 27'h000002e8, 5'd1, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000182, 5'd27, 27'h00000086, 5'd14, 27'h000000da, 32'h00000400,
  1'd1,  5'd25, 27'h00000082, 5'd28, 27'h000000f4, 5'd25, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f8, 5'd8, 27'h00000000, 5'd9, 27'h0000031a, 32'h00000400,
  1'd1,  5'd0, 27'h00000185, 5'd8, 27'h00000226, 5'd19, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000284, 5'd5, 27'h000000fa, 5'd26, 27'h00000165, 32'h00000400,
  1'd1,  5'd1, 27'h000001f1, 5'd15, 27'h0000031f, 5'd6, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000b0, 5'd16, 27'h00000363, 5'd18, 27'h000003aa, 32'h00000400,
  1'd1,  5'd3, 27'h000000b0, 5'd17, 27'h00000149, 5'd29, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000005c, 5'd29, 27'h00000284, 5'd6, 27'h000003ce, 32'h00000400,
  1'd1,  5'd0, 27'h000001f0, 5'd30, 27'h000002ca, 5'd18, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000220, 5'd29, 27'h00000072, 5'd30, 27'h000002ef, 32'h00000400,
  1'd1,  5'd12, 27'h00000118, 5'd6, 27'h000001c0, 5'd6, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000177, 5'd5, 27'h000001d2, 5'd19, 27'h00000066, 32'h00000400,
  1'd1,  5'd13, 27'h00000321, 5'd6, 27'h00000389, 5'd27, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000162, 5'd15, 27'h0000033c, 5'd8, 27'h000001c6, 32'h00000400,
  1'd1,  5'd12, 27'h0000000f, 5'd15, 27'h0000024b, 5'd20, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b9, 5'd19, 27'h000003d9, 5'd29, 27'h00000114, 32'h00000400,
  1'd1,  5'd10, 27'h000001ed, 5'd26, 27'h00000001, 5'd5, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000039d, 5'd26, 27'h00000093, 5'd17, 27'h000001f9, 32'h00000400,
  1'd1,  5'd12, 27'h0000003d, 5'd26, 27'h000001b3, 5'd29, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000234, 5'd5, 27'h00000144, 5'd9, 27'h00000380, 32'h00000400,
  1'd1,  5'd20, 27'h000003a5, 5'd6, 27'h000000eb, 5'd17, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000074, 5'd8, 27'h00000092, 5'd30, 27'h00000365, 32'h00000400,
  1'd1,  5'd23, 27'h0000037a, 5'd17, 27'h000003fa, 5'd7, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000007e, 5'd18, 27'h000002a6, 5'd19, 27'h000000ec, 32'h00000400,
  1'd1,  5'd25, 27'h0000002b, 5'd16, 27'h00000159, 5'd28, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000168, 5'd27, 27'h000000fe, 5'd9, 27'h0000012d, 32'h00000400,
  1'd1,  5'd21, 27'h0000003a, 5'd29, 27'h000001b9, 5'd17, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003b4, 5'd30, 27'h000002f2, 5'd30, 27'h000000a8, 32'h00000400,
  1'd1,  5'd7, 27'h00000264, 5'd1, 27'h0000003e, 5'd8, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000055, 5'd1, 27'h000003bb, 5'd18, 27'h000002d8, 32'h00000400,
  1'd1,  5'd9, 27'h00000210, 5'd4, 27'h000000b4, 5'd29, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033a, 5'd13, 27'h00000317, 5'd3, 27'h000002dc, 32'h00000400,
  1'd1,  5'd7, 27'h0000037f, 5'd11, 27'h000001de, 5'd15, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002b8, 5'd10, 27'h00000356, 5'd21, 27'h00000278, 32'h00000400,
  1'd1,  5'd7, 27'h00000323, 5'd25, 27'h0000011e, 5'd2, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ec, 5'd23, 27'h00000199, 5'd13, 27'h0000021c, 32'h00000400,
  1'd1,  5'd7, 27'h00000359, 5'd23, 27'h0000018d, 5'd23, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000065, 5'd4, 27'h000001c8, 5'd8, 27'h00000210, 32'h00000400,
  1'd1,  5'd19, 27'h0000017c, 5'd4, 27'h00000139, 5'd15, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000156, 5'd1, 27'h000003e1, 5'd27, 27'h0000015e, 32'h00000400,
  1'd1,  5'd19, 27'h00000020, 5'd12, 27'h00000038, 5'd1, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002a4, 5'd11, 27'h00000129, 5'd11, 27'h00000134, 32'h00000400,
  1'd1,  5'd19, 27'h0000010d, 5'd10, 27'h0000029e, 5'd23, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ec, 5'd25, 27'h0000015b, 5'd3, 27'h0000003a, 32'h00000400,
  1'd1,  5'd17, 27'h000001e2, 5'd24, 27'h00000290, 5'd12, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000017d, 5'd22, 27'h000001f5, 5'd22, 27'h00000233, 32'h00000400,
  1'd1,  5'd29, 27'h0000016a, 5'd3, 27'h000002a3, 5'd3, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000004f, 5'd2, 27'h00000085, 5'd11, 27'h00000307, 32'h00000400,
  1'd1,  5'd29, 27'h00000065, 5'd3, 27'h0000015c, 5'd25, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000dc, 5'd10, 27'h000003f8, 5'd3, 27'h0000004a, 32'h00000400,
  1'd1,  5'd29, 27'h00000065, 5'd11, 27'h00000200, 5'd14, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000036c, 5'd11, 27'h000002bc, 5'd25, 27'h000002fa, 32'h00000400,
  1'd1,  5'd28, 27'h00000041, 5'd25, 27'h0000013c, 5'd3, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d2, 5'd25, 27'h00000323, 5'd10, 27'h00000257, 32'h00000400,
  1'd1,  5'd26, 27'h0000008a, 5'd25, 27'h00000129, 5'd23, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c1, 5'd3, 27'h000002dd, 5'd0, 27'h000002a5, 32'h00000400,
  1'd1,  5'd6, 27'h000003f8, 5'd4, 27'h00000242, 5'd13, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a2, 5'd5, 27'h0000001a, 5'd21, 27'h00000347, 32'h00000400,
  1'd1,  5'd9, 27'h00000265, 5'd13, 27'h00000063, 5'd5, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000fc, 5'd11, 27'h000002ec, 5'd19, 27'h000001df, 32'h00000400,
  1'd1,  5'd8, 27'h0000004c, 5'd13, 27'h000001b6, 5'd26, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021c, 5'd24, 27'h000001bd, 5'd5, 27'h000001a3, 32'h00000400,
  1'd1,  5'd7, 27'h00000331, 5'd22, 27'h0000037a, 5'd19, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000008a, 5'd25, 27'h0000020a, 5'd26, 27'h00000217, 32'h00000400,
  1'd1,  5'd18, 27'h000003a4, 5'd0, 27'h000002cc, 5'd1, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000311, 5'd3, 27'h000003ab, 5'd12, 27'h000003aa, 32'h00000400,
  1'd1,  5'd17, 27'h000001f3, 5'd0, 27'h000000b8, 5'd23, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000225, 5'd13, 27'h0000037a, 5'd7, 27'h00000102, 32'h00000400,
  1'd1,  5'd20, 27'h00000057, 5'd10, 27'h000002fb, 5'd17, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003b3, 5'd10, 27'h00000176, 5'd26, 27'h000001ff, 32'h00000400,
  1'd1,  5'd19, 27'h00000150, 5'd22, 27'h0000016f, 5'd7, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001be, 5'd21, 27'h000002e7, 5'd17, 27'h00000388, 32'h00000400,
  1'd1,  5'd20, 27'h000000c0, 5'd21, 27'h00000387, 5'd26, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000006a, 5'd4, 27'h00000286, 5'd10, 27'h00000105, 32'h00000400,
  1'd1,  5'd28, 27'h00000302, 5'd4, 27'h00000099, 5'd17, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000039c, 5'd3, 27'h000001e6, 5'd29, 27'h00000107, 32'h00000400,
  1'd1,  5'd30, 27'h000001f8, 5'd12, 27'h000000c8, 5'd8, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000031c, 5'd13, 27'h0000017a, 5'd20, 27'h00000265, 32'h00000400,
  1'd1,  5'd29, 27'h0000029b, 5'd10, 27'h0000037d, 5'd28, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000042, 5'd25, 27'h00000048, 5'd6, 27'h00000090, 32'h00000400,
  1'd1,  5'd28, 27'h0000008b, 5'd22, 27'h000002f2, 5'd16, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000039d, 5'd24, 27'h00000275, 5'd27, 27'h0000019a, 32'h00000400,
  1'd1,  5'd8, 27'h00000197, 5'd5, 27'h00000287, 5'd0, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000005c, 5'd8, 27'h000001d3, 5'd14, 27'h0000007b, 32'h00000400,
  1'd1,  5'd7, 27'h000002bc, 5'd8, 27'h000000de, 5'd23, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000243, 5'd15, 27'h00000227, 5'd1, 27'h000001ae, 32'h00000400,
  1'd1,  5'd7, 27'h00000107, 5'd15, 27'h00000297, 5'd11, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000c, 5'd20, 27'h00000237, 5'd21, 27'h0000016b, 32'h00000400,
  1'd1,  5'd9, 27'h000003de, 5'd28, 27'h0000029d, 5'd1, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000299, 5'd26, 27'h000000a6, 5'd14, 27'h00000243, 32'h00000400,
  1'd1,  5'd8, 27'h0000021c, 5'd27, 27'h00000023, 5'd25, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e7, 5'd5, 27'h00000123, 5'd1, 27'h00000201, 32'h00000400,
  1'd1,  5'd18, 27'h00000272, 5'd7, 27'h0000026a, 5'd15, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002b4, 5'd9, 27'h000001c7, 5'd22, 27'h00000284, 32'h00000400,
  1'd1,  5'd16, 27'h000000ba, 5'd16, 27'h0000009c, 5'd2, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000112, 5'd20, 27'h0000022d, 5'd14, 27'h000001c3, 32'h00000400,
  1'd1,  5'd16, 27'h000002da, 5'd16, 27'h00000309, 5'd23, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b2, 5'd26, 27'h00000381, 5'd1, 27'h000003db, 32'h00000400,
  1'd1,  5'd18, 27'h00000115, 5'd29, 27'h0000029d, 5'd13, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000155, 5'd28, 27'h00000142, 5'd25, 27'h000000d3, 32'h00000400,
  1'd1,  5'd26, 27'h000000a3, 5'd6, 27'h00000188, 5'd1, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000299, 5'd9, 27'h00000231, 5'd13, 27'h00000320, 32'h00000400,
  1'd1,  5'd29, 27'h0000016a, 5'd7, 27'h000002a3, 5'd22, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000269, 5'd20, 27'h000001b8, 5'd4, 27'h0000038e, 32'h00000400,
  1'd1,  5'd27, 27'h00000291, 5'd17, 27'h00000082, 5'd11, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000081, 5'd19, 27'h0000024f, 5'd22, 27'h000000ef, 32'h00000400,
  1'd1,  5'd28, 27'h00000200, 5'd26, 27'h0000001e, 5'd1, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000317, 5'd29, 27'h000001ec, 5'd12, 27'h000003fc, 32'h00000400,
  1'd1,  5'd26, 27'h00000358, 5'd30, 27'h000002f9, 5'd21, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ed, 5'd9, 27'h0000022e, 5'd8, 27'h0000009b, 32'h00000400,
  1'd1,  5'd7, 27'h000001c0, 5'd8, 27'h000003ed, 5'd17, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003c1, 5'd10, 27'h00000007, 5'd27, 27'h0000018a, 32'h00000400,
  1'd1,  5'd9, 27'h00000272, 5'd16, 27'h00000152, 5'd9, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000094, 5'd15, 27'h00000374, 5'd17, 27'h000001d9, 32'h00000400,
  1'd1,  5'd8, 27'h000002c0, 5'd16, 27'h000000bd, 5'd29, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000375, 5'd28, 27'h000002f7, 5'd10, 27'h0000014d, 32'h00000400,
  1'd1,  5'd9, 27'h000001d8, 5'd27, 27'h000000c8, 5'd17, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000263, 5'd26, 27'h00000273, 5'd27, 27'h00000278, 32'h00000400,
  1'd1,  5'd17, 27'h000000d2, 5'd8, 27'h000002d7, 5'd9, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000025, 5'd7, 27'h00000249, 5'd17, 27'h0000010e, 32'h00000400,
  1'd1,  5'd15, 27'h00000252, 5'd5, 27'h0000030c, 5'd28, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000033d, 5'd18, 27'h000000ba, 5'd7, 27'h00000144, 32'h00000400,
  1'd1,  5'd19, 27'h000002ea, 5'd15, 27'h0000033b, 5'd17, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000006b, 5'd20, 27'h000001ea, 5'd28, 27'h00000123, 32'h00000400,
  1'd1,  5'd16, 27'h0000034d, 5'd27, 27'h000001c0, 5'd9, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000028d, 5'd28, 27'h00000110, 5'd18, 27'h00000154, 32'h00000400,
  1'd1,  5'd17, 27'h000002de, 5'd29, 27'h00000102, 5'd29, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023b, 5'd7, 27'h00000316, 5'd8, 27'h000001cc, 32'h00000400,
  1'd1,  5'd28, 27'h000000ad, 5'd8, 27'h000001f3, 5'd18, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000030a, 5'd8, 27'h000002cb, 5'd28, 27'h00000221, 32'h00000400,
  1'd1,  5'd27, 27'h000002e5, 5'd16, 27'h000003a6, 5'd5, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f1, 5'd17, 27'h000001ac, 5'd20, 27'h00000004, 32'h00000400,
  1'd1,  5'd30, 27'h0000036b, 5'd18, 27'h000003f3, 5'd28, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000018b, 5'd30, 27'h000001cb, 5'd6, 27'h00000331, 32'h00000400,
  1'd1,  5'd28, 27'h000002f6, 5'd30, 27'h000000aa, 5'd17, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000094, 5'd29, 27'h0000027d, 5'd26, 27'h000002fb, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000360, 5'd0, 27'h000002e9, 5'd3, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000fd, 5'd2, 27'h0000026f, 5'd14, 27'h0000029f, 32'h00000400,
  1'd1,  5'd3, 27'h000001c0, 5'd1, 27'h0000027e, 5'd24, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000286, 5'd13, 27'h00000233, 5'd0, 27'h00000277, 32'h00000400,
  1'd1,  5'd4, 27'h000001c6, 5'd10, 27'h00000168, 5'd14, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000162, 5'd12, 27'h000000e6, 5'd23, 27'h000000c6, 32'h00000400,
  1'd1,  5'd2, 27'h00000002, 5'd25, 27'h0000030e, 5'd2, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000150, 5'd20, 27'h0000036a, 5'd11, 27'h00000319, 32'h00000400,
  1'd1,  5'd1, 27'h000001f6, 5'd20, 27'h000003d3, 5'd22, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000390, 5'd4, 27'h000002fb, 5'd2, 27'h00000002, 32'h00000400,
  1'd1,  5'd10, 27'h00000363, 5'd1, 27'h000003ce, 5'd10, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001e8, 5'd4, 27'h000003c8, 5'd23, 27'h000001ef, 32'h00000400,
  1'd1,  5'd15, 27'h00000017, 5'd10, 27'h0000027d, 5'd0, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000146, 5'd13, 27'h00000107, 5'd15, 27'h0000003a, 32'h00000400,
  1'd1,  5'd11, 27'h00000306, 5'd11, 27'h000001e7, 5'd21, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f5, 5'd24, 27'h00000102, 5'd4, 27'h000000d9, 32'h00000400,
  1'd1,  5'd14, 27'h00000301, 5'd25, 27'h00000210, 5'd10, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000249, 5'd23, 27'h000000aa, 5'd23, 27'h000002f9, 32'h00000400,
  1'd1,  5'd23, 27'h00000234, 5'd4, 27'h00000280, 5'd3, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001e8, 5'd1, 27'h000002b9, 5'd11, 27'h000003d9, 32'h00000400,
  1'd1,  5'd22, 27'h0000032b, 5'd2, 27'h00000081, 5'd25, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003cb, 5'd12, 27'h00000088, 5'd3, 27'h00000337, 32'h00000400,
  1'd1,  5'd20, 27'h00000324, 5'd12, 27'h000000f5, 5'd11, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000120, 5'd13, 27'h000002e7, 5'd24, 27'h00000025, 32'h00000400,
  1'd1,  5'd21, 27'h000002d1, 5'd23, 27'h00000241, 5'd4, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f9, 5'd24, 27'h00000333, 5'd15, 27'h00000068, 32'h00000400,
  1'd1,  5'd22, 27'h000001f6, 5'd21, 27'h000003e2, 5'd21, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000be, 5'd4, 27'h000003aa, 5'd7, 27'h00000192, 32'h00000400,
  1'd1,  5'd4, 27'h000000c2, 5'd3, 27'h00000291, 5'd19, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b2, 5'd2, 27'h000002c2, 5'd27, 27'h000003a2, 32'h00000400,
  1'd1,  5'd2, 27'h0000030b, 5'd15, 27'h00000149, 5'd5, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000028b, 5'd12, 27'h0000005d, 5'd19, 27'h0000039f, 32'h00000400,
  1'd1,  5'd1, 27'h0000020a, 5'd14, 27'h0000001d, 5'd28, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000f5, 5'd25, 27'h000002fa, 5'd8, 27'h00000396, 32'h00000400,
  1'd1,  5'd1, 27'h00000067, 5'd22, 27'h00000083, 5'd19, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000009a, 5'd22, 27'h000003ea, 5'd29, 27'h000003bc, 32'h00000400,
  1'd1,  5'd12, 27'h00000160, 5'd1, 27'h000000aa, 5'd10, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000131, 5'd4, 27'h00000339, 5'd20, 27'h000002a1, 32'h00000400,
  1'd1,  5'd12, 27'h000000e7, 5'd2, 27'h00000100, 5'd30, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000012f, 5'd11, 27'h000000d4, 5'd7, 27'h0000017f, 32'h00000400,
  1'd1,  5'd15, 27'h0000012b, 5'd14, 27'h00000262, 5'd19, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000113, 5'd10, 27'h000003da, 5'd26, 27'h000002fc, 32'h00000400,
  1'd1,  5'd10, 27'h000002b2, 5'd22, 27'h0000023c, 5'd9, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000390, 5'd25, 27'h00000352, 5'd19, 27'h000001de, 32'h00000400,
  1'd1,  5'd12, 27'h00000385, 5'd22, 27'h00000306, 5'd26, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002cb, 5'd3, 27'h0000011c, 5'd8, 27'h00000360, 32'h00000400,
  1'd1,  5'd24, 27'h00000107, 5'd4, 27'h0000008e, 5'd19, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000140, 5'd1, 27'h000003d2, 5'd26, 27'h000003d5, 32'h00000400,
  1'd1,  5'd25, 27'h0000014b, 5'd12, 27'h000002dc, 5'd8, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a2, 5'd13, 27'h000001c0, 5'd20, 27'h000000ab, 32'h00000400,
  1'd1,  5'd23, 27'h0000011b, 5'd13, 27'h00000129, 5'd27, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003f8, 5'd24, 27'h00000266, 5'd6, 27'h0000015d, 32'h00000400,
  1'd1,  5'd23, 27'h00000389, 5'd23, 27'h0000019d, 5'd18, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000024, 5'd25, 27'h00000063, 5'd26, 27'h000001dd, 32'h00000400,
  1'd1,  5'd3, 27'h00000358, 5'd7, 27'h00000062, 5'd5, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003ad, 5'd5, 27'h00000339, 5'd14, 27'h00000251, 32'h00000400,
  1'd1,  5'd1, 27'h0000016d, 5'd8, 27'h00000035, 5'd21, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000031b, 5'd17, 27'h000001f4, 5'd3, 27'h00000027, 32'h00000400,
  1'd1,  5'd0, 27'h0000038c, 5'd15, 27'h0000032a, 5'd10, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e5, 5'd18, 27'h0000014c, 5'd21, 27'h0000004d, 32'h00000400,
  1'd1,  5'd3, 27'h00000146, 5'd26, 27'h000003d8, 5'd2, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000341, 5'd27, 27'h0000028a, 5'd15, 27'h000000ab, 32'h00000400,
  1'd1,  5'd2, 27'h000002ce, 5'd27, 27'h000002cd, 5'd25, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000c7, 5'd9, 27'h000001bc, 5'd2, 27'h000002b5, 32'h00000400,
  1'd1,  5'd10, 27'h0000022a, 5'd9, 27'h000002fb, 5'd15, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000247, 5'd9, 27'h000002f3, 5'd21, 27'h000002c4, 32'h00000400,
  1'd1,  5'd14, 27'h0000019c, 5'd16, 27'h000001f3, 5'd4, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001af, 5'd17, 27'h000002b5, 5'd15, 27'h000000cd, 32'h00000400,
  1'd1,  5'd12, 27'h00000140, 5'd20, 27'h000000d7, 5'd25, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000192, 5'd29, 27'h000001ef, 5'd3, 27'h0000004b, 32'h00000400,
  1'd1,  5'd13, 27'h000003af, 5'd26, 27'h0000019b, 5'd11, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c0, 5'd27, 27'h00000178, 5'd21, 27'h0000015b, 32'h00000400,
  1'd1,  5'd20, 27'h000003ad, 5'd9, 27'h000001a9, 5'd4, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001d6, 5'd8, 27'h000001be, 5'd13, 27'h000003ee, 32'h00000400,
  1'd1,  5'd23, 27'h0000034b, 5'd8, 27'h0000013d, 5'd22, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001eb, 5'd19, 27'h000003a3, 5'd0, 27'h0000037a, 32'h00000400,
  1'd1,  5'd25, 27'h0000005f, 5'd20, 27'h00000218, 5'd15, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000392, 5'd19, 27'h000003b2, 5'd22, 27'h00000332, 32'h00000400,
  1'd1,  5'd25, 27'h000001d7, 5'd29, 27'h00000287, 5'd2, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b2, 5'd27, 27'h00000255, 5'd14, 27'h0000036e, 32'h00000400,
  1'd1,  5'd21, 27'h0000039d, 5'd25, 27'h0000036b, 5'd22, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000067, 5'd9, 27'h0000036f, 5'd6, 27'h000002d8, 32'h00000400,
  1'd1,  5'd3, 27'h000003e8, 5'd7, 27'h00000209, 5'd16, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000003a, 5'd9, 27'h00000118, 5'd29, 27'h00000130, 32'h00000400,
  1'd1,  5'd0, 27'h00000259, 5'd19, 27'h00000226, 5'd6, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000114, 5'd20, 27'h00000144, 5'd17, 27'h00000224, 32'h00000400,
  1'd1,  5'd2, 27'h00000362, 5'd20, 27'h000001eb, 5'd30, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002cb, 5'd30, 27'h000002da, 5'd6, 27'h000002a2, 32'h00000400,
  1'd1,  5'd2, 27'h000001c6, 5'd30, 27'h0000000c, 5'd19, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000006b, 5'd26, 27'h000000e4, 5'd30, 27'h00000190, 32'h00000400,
  1'd1,  5'd15, 27'h0000002a, 5'd5, 27'h00000193, 5'd7, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003f9, 5'd7, 27'h00000133, 5'd16, 27'h0000022c, 32'h00000400,
  1'd1,  5'd12, 27'h00000145, 5'd6, 27'h00000387, 5'd28, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000b0, 5'd19, 27'h0000006b, 5'd7, 27'h00000251, 32'h00000400,
  1'd1,  5'd11, 27'h00000232, 5'd19, 27'h000000b8, 5'd16, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000123, 5'd19, 27'h000003d7, 5'd29, 27'h000000f9, 32'h00000400,
  1'd1,  5'd15, 27'h000000ec, 5'd29, 27'h00000129, 5'd9, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000017e, 5'd25, 27'h00000389, 5'd20, 27'h0000025d, 32'h00000400,
  1'd1,  5'd14, 27'h000002b1, 5'd26, 27'h00000322, 5'd30, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003b5, 5'd9, 27'h0000019d, 5'd9, 27'h00000382, 32'h00000400,
  1'd1,  5'd21, 27'h000001c2, 5'd6, 27'h0000039f, 5'd18, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000311, 5'd9, 27'h0000039b, 5'd30, 27'h000000e3, 32'h00000400,
  1'd1,  5'd22, 27'h000003f8, 5'd15, 27'h00000244, 5'd9, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000029c, 5'd17, 27'h00000398, 5'd20, 27'h0000018c, 32'h00000400,
  1'd1,  5'd21, 27'h0000006f, 5'd18, 27'h00000060, 5'd27, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001b4, 5'd26, 27'h000001ad, 5'd6, 27'h00000053, 32'h00000400,
  1'd1,  5'd23, 27'h00000140, 5'd28, 27'h00000148, 5'd18, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002cc, 5'd30, 27'h000002fb, 5'd27, 27'h00000033, 32'h00000400,
  1'd1,  5'd6, 27'h000003c2, 5'd2, 27'h000002d7, 5'd9, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000028b, 5'd0, 27'h000002af, 5'd18, 27'h00000293, 32'h00000400,
  1'd1,  5'd6, 27'h00000349, 5'd1, 27'h000003c5, 5'd30, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000291, 5'd10, 27'h00000335, 5'd0, 27'h000001a6, 32'h00000400,
  1'd1,  5'd9, 27'h000001c5, 5'd11, 27'h00000376, 5'd12, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000320, 5'd13, 27'h000001f9, 5'd25, 27'h000002a3, 32'h00000400,
  1'd1,  5'd8, 27'h000002fd, 5'd22, 27'h0000038d, 5'd3, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000276, 5'd23, 27'h000003be, 5'd11, 27'h000001c8, 32'h00000400,
  1'd1,  5'd7, 27'h000001cd, 5'd23, 27'h00000381, 5'd23, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003c4, 5'd2, 27'h0000016b, 5'd9, 27'h000002c8, 32'h00000400,
  1'd1,  5'd20, 27'h0000010f, 5'd0, 27'h000001fe, 5'd15, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000011b, 5'd0, 27'h0000022e, 5'd30, 27'h00000294, 32'h00000400,
  1'd1,  5'd18, 27'h00000053, 5'd10, 27'h00000215, 5'd4, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000198, 5'd12, 27'h000000f2, 5'd13, 27'h000000a4, 32'h00000400,
  1'd1,  5'd19, 27'h000001ac, 5'd14, 27'h0000033b, 5'd25, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000059, 5'd21, 27'h00000060, 5'd4, 27'h00000351, 32'h00000400,
  1'd1,  5'd20, 27'h000000bb, 5'd21, 27'h0000035d, 5'd13, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ba, 5'd25, 27'h000000f7, 5'd25, 27'h0000005b, 32'h00000400,
  1'd1,  5'd26, 27'h000002e9, 5'd0, 27'h0000000d, 5'd5, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000017f, 5'd3, 27'h00000353, 5'd13, 27'h000001b0, 32'h00000400,
  1'd1,  5'd25, 27'h0000038f, 5'd0, 27'h0000008e, 5'd21, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001fb, 5'd14, 27'h000001f1, 5'd3, 27'h0000038d, 32'h00000400,
  1'd1,  5'd28, 27'h0000028d, 5'd13, 27'h000002aa, 5'd14, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000137, 5'd12, 27'h00000315, 5'd22, 27'h0000008c, 32'h00000400,
  1'd1,  5'd29, 27'h0000008d, 5'd25, 27'h000002c5, 5'd3, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002d1, 5'd23, 27'h00000162, 5'd14, 27'h00000237, 32'h00000400,
  1'd1,  5'd29, 27'h00000375, 5'd22, 27'h0000003f, 5'd21, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000120, 5'd3, 27'h000000fc, 5'd3, 27'h000003dc, 32'h00000400,
  1'd1,  5'd8, 27'h000000f0, 5'd3, 27'h00000292, 5'd11, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000311, 5'd0, 27'h00000113, 5'd24, 27'h000001d0, 32'h00000400,
  1'd1,  5'd6, 27'h0000012d, 5'd11, 27'h000001dc, 5'd9, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000188, 5'd12, 27'h000002ff, 5'd18, 27'h00000264, 32'h00000400,
  1'd1,  5'd5, 27'h00000277, 5'd11, 27'h00000101, 5'd29, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002ed, 5'd21, 27'h00000135, 5'd6, 27'h000003cb, 32'h00000400,
  1'd1,  5'd8, 27'h00000016, 5'd22, 27'h00000165, 5'd16, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000065, 5'd20, 27'h00000396, 5'd27, 27'h000003d4, 32'h00000400,
  1'd1,  5'd16, 27'h00000327, 5'd2, 27'h000001e0, 5'd3, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000107, 5'd4, 27'h0000039a, 5'd11, 27'h00000213, 32'h00000400,
  1'd1,  5'd18, 27'h00000349, 5'd1, 27'h00000322, 5'd22, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000026d, 5'd10, 27'h0000021a, 5'd6, 27'h0000016b, 32'h00000400,
  1'd1,  5'd19, 27'h00000270, 5'd12, 27'h000002a2, 5'd15, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000071, 5'd14, 27'h000000ab, 5'd28, 27'h00000379, 32'h00000400,
  1'd1,  5'd15, 27'h0000028b, 5'd24, 27'h00000246, 5'd6, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a4, 5'd20, 27'h000002bd, 5'd15, 27'h000002ff, 32'h00000400,
  1'd1,  5'd20, 27'h0000028c, 5'd25, 27'h00000350, 5'd27, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000314, 5'd4, 27'h000000ac, 5'd7, 27'h000003e3, 32'h00000400,
  1'd1,  5'd28, 27'h00000390, 5'd1, 27'h0000002a, 5'd18, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c9, 5'd0, 27'h000003ea, 5'd27, 27'h00000185, 32'h00000400,
  1'd1,  5'd27, 27'h0000025d, 5'd13, 27'h00000328, 5'd7, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000368, 5'd13, 27'h00000339, 5'd17, 27'h00000047, 32'h00000400,
  1'd1,  5'd28, 27'h00000221, 5'd11, 27'h000001f3, 5'd28, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a3, 5'd22, 27'h000003fd, 5'd7, 27'h00000006, 32'h00000400,
  1'd1,  5'd30, 27'h000001df, 5'd24, 27'h000001b0, 5'd19, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001e6, 5'd23, 27'h000000da, 5'd29, 27'h00000348, 32'h00000400,
  1'd1,  5'd7, 27'h0000012e, 5'd5, 27'h00000350, 5'd1, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000006d, 5'd5, 27'h000000ec, 5'd14, 27'h000003e5, 32'h00000400,
  1'd1,  5'd6, 27'h00000220, 5'd8, 27'h00000004, 5'd23, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000159, 5'd18, 27'h00000099, 5'd1, 27'h000001b5, 32'h00000400,
  1'd1,  5'd9, 27'h00000071, 5'd17, 27'h000003b3, 5'd15, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c5, 5'd18, 27'h0000014a, 5'd24, 27'h0000014e, 32'h00000400,
  1'd1,  5'd7, 27'h0000016f, 5'd27, 27'h00000122, 5'd4, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001af, 5'd28, 27'h0000013a, 5'd13, 27'h00000022, 32'h00000400,
  1'd1,  5'd9, 27'h00000249, 5'd30, 27'h00000123, 5'd23, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000357, 5'd6, 27'h0000014e, 5'd2, 27'h0000012c, 32'h00000400,
  1'd1,  5'd15, 27'h00000200, 5'd8, 27'h00000246, 5'd11, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003fb, 5'd9, 27'h000002f5, 5'd21, 27'h000001e6, 32'h00000400,
  1'd1,  5'd16, 27'h000001c9, 5'd15, 27'h000003ac, 5'd2, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000357, 5'd19, 27'h00000207, 5'd12, 27'h000003e4, 32'h00000400,
  1'd1,  5'd19, 27'h00000337, 5'd16, 27'h0000009e, 5'd21, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000210, 5'd29, 27'h00000382, 5'd5, 27'h0000003a, 32'h00000400,
  1'd1,  5'd16, 27'h000003e6, 5'd30, 27'h00000292, 5'd13, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000245, 5'd29, 27'h0000035e, 5'd25, 27'h000002c7, 32'h00000400,
  1'd1,  5'd30, 27'h000002f0, 5'd8, 27'h00000204, 5'd0, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e3, 5'd6, 27'h0000031a, 5'd11, 27'h0000016c, 32'h00000400,
  1'd1,  5'd26, 27'h0000029b, 5'd9, 27'h0000027c, 5'd20, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002be, 5'd20, 27'h00000066, 5'd4, 27'h00000143, 32'h00000400,
  1'd1,  5'd30, 27'h0000000d, 5'd20, 27'h00000238, 5'd12, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000023c, 5'd18, 27'h000002a2, 5'd25, 27'h00000028, 32'h00000400,
  1'd1,  5'd28, 27'h000001fe, 5'd27, 27'h000003ea, 5'd4, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012a, 5'd26, 27'h00000072, 5'd13, 27'h000003c9, 32'h00000400,
  1'd1,  5'd25, 27'h000003d3, 5'd28, 27'h00000333, 5'd23, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000007b, 5'd7, 27'h00000082, 5'd8, 27'h0000000b, 32'h00000400,
  1'd1,  5'd7, 27'h00000246, 5'd8, 27'h00000031, 5'd17, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000211, 5'd9, 27'h0000036e, 5'd26, 27'h00000358, 32'h00000400,
  1'd1,  5'd5, 27'h000002a7, 5'd16, 27'h00000212, 5'd7, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000354, 5'd16, 27'h00000128, 5'd19, 27'h0000039b, 32'h00000400,
  1'd1,  5'd7, 27'h0000021b, 5'd18, 27'h000002dd, 5'd29, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012d, 5'd28, 27'h000000d7, 5'd7, 27'h000002d0, 32'h00000400,
  1'd1,  5'd6, 27'h00000191, 5'd27, 27'h0000010b, 5'd18, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b8, 5'd30, 27'h00000372, 5'd30, 27'h000002d8, 32'h00000400,
  1'd1,  5'd15, 27'h0000025b, 5'd6, 27'h00000201, 5'd7, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000280, 5'd10, 27'h0000000d, 5'd19, 27'h00000290, 32'h00000400,
  1'd1,  5'd18, 27'h00000132, 5'd5, 27'h00000352, 5'd27, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000be, 5'd20, 27'h0000018d, 5'd8, 27'h0000029d, 32'h00000400,
  1'd1,  5'd18, 27'h000000ee, 5'd19, 27'h00000159, 5'd19, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003cd, 5'd18, 27'h00000311, 5'd30, 27'h0000016e, 32'h00000400,
  1'd1,  5'd18, 27'h00000225, 5'd26, 27'h00000259, 5'd8, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000239, 5'd28, 27'h000001ff, 5'd17, 27'h000000ce, 32'h00000400,
  1'd1,  5'd16, 27'h000003ba, 5'd29, 27'h0000018e, 5'd25, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e0, 5'd7, 27'h00000096, 5'd9, 27'h000003a6, 32'h00000400,
  1'd1,  5'd29, 27'h00000012, 5'd6, 27'h00000157, 5'd19, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000307, 5'd8, 27'h00000171, 5'd28, 27'h00000105, 32'h00000400,
  1'd1,  5'd29, 27'h000000f8, 5'd19, 27'h000000a3, 5'd5, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000394, 5'd17, 27'h000001bc, 5'd19, 27'h0000008a, 32'h00000400,
  1'd1,  5'd28, 27'h000000f0, 5'd15, 27'h000002de, 5'd27, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000056, 5'd28, 27'h000002a0, 5'd5, 27'h000001cc, 32'h00000400,
  1'd1,  5'd30, 27'h000000ea, 5'd27, 27'h00000011, 5'd17, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019d, 5'd30, 27'h000001d6, 5'd30, 27'h0000027c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000231, 5'd0, 27'h00000319, 5'd4, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000322, 5'd0, 27'h000000af, 5'd13, 27'h00000125, 32'h00000400,
  1'd1,  5'd1, 27'h0000019d, 5'd1, 27'h000003a3, 5'd22, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000128, 5'd10, 27'h00000165, 5'd2, 27'h00000318, 32'h00000400,
  1'd1,  5'd3, 27'h000002ab, 5'd11, 27'h0000020d, 5'd10, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e1, 5'd13, 27'h00000204, 5'd24, 27'h000003a7, 32'h00000400,
  1'd1,  5'd2, 27'h0000021b, 5'd24, 27'h000003a7, 5'd4, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000094, 5'd24, 27'h0000021e, 5'd10, 27'h000003c2, 32'h00000400,
  1'd1,  5'd2, 27'h000001a6, 5'd24, 27'h00000253, 5'd23, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000255, 5'd3, 27'h0000036d, 5'd2, 27'h0000031e, 32'h00000400,
  1'd1,  5'd12, 27'h000001b5, 5'd1, 27'h00000303, 5'd11, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000187, 5'd3, 27'h00000008, 5'd24, 27'h000003f1, 32'h00000400,
  1'd1,  5'd13, 27'h00000374, 5'd12, 27'h0000007f, 5'd2, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000008a, 5'd15, 27'h000001a6, 5'd15, 27'h00000024, 32'h00000400,
  1'd1,  5'd11, 27'h0000018d, 5'd15, 27'h000000eb, 5'd24, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000366, 5'd23, 27'h000002ab, 5'd3, 27'h00000019, 32'h00000400,
  1'd1,  5'd12, 27'h00000051, 5'd21, 27'h00000216, 5'd11, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a0, 5'd20, 27'h00000381, 5'd24, 27'h000001f1, 32'h00000400,
  1'd1,  5'd25, 27'h00000018, 5'd0, 27'h0000039e, 5'd2, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000108, 5'd3, 27'h00000308, 5'd12, 27'h00000328, 32'h00000400,
  1'd1,  5'd22, 27'h00000022, 5'd2, 27'h000003c1, 5'd23, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000147, 5'd14, 27'h0000020a, 5'd2, 27'h000001c3, 32'h00000400,
  1'd1,  5'd23, 27'h00000055, 5'd10, 27'h00000180, 5'd14, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000329, 5'd10, 27'h000002b0, 5'd24, 27'h00000378, 32'h00000400,
  1'd1,  5'd24, 27'h0000039d, 5'd21, 27'h00000265, 5'd1, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003c4, 5'd23, 27'h000002da, 5'd11, 27'h000001f0, 32'h00000400,
  1'd1,  5'd22, 27'h000000ff, 5'd23, 27'h0000010c, 5'd21, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000360, 5'd1, 27'h00000328, 5'd9, 27'h00000223, 32'h00000400,
  1'd1,  5'd2, 27'h000002e3, 5'd4, 27'h00000300, 5'd20, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000195, 5'd4, 27'h0000035d, 5'd27, 27'h000002d6, 32'h00000400,
  1'd1,  5'd2, 27'h00000023, 5'd14, 27'h000002b1, 5'd8, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a3, 5'd10, 27'h000003f0, 5'd16, 27'h000002ec, 32'h00000400,
  1'd1,  5'd2, 27'h00000379, 5'd15, 27'h000000b4, 5'd26, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000218, 5'd25, 27'h00000042, 5'd5, 27'h00000199, 32'h00000400,
  1'd1,  5'd2, 27'h000001ae, 5'd22, 27'h0000017a, 5'd18, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000031e, 5'd24, 27'h00000271, 5'd25, 27'h00000379, 32'h00000400,
  1'd1,  5'd10, 27'h000001c7, 5'd0, 27'h0000034f, 5'd6, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000350, 5'd1, 27'h0000027b, 5'd15, 27'h00000213, 32'h00000400,
  1'd1,  5'd14, 27'h00000346, 5'd5, 27'h00000026, 5'd29, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ac, 5'd14, 27'h000000ab, 5'd6, 27'h0000004b, 32'h00000400,
  1'd1,  5'd13, 27'h0000004a, 5'd12, 27'h00000151, 5'd20, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017f, 5'd14, 27'h000003b2, 5'd28, 27'h00000165, 32'h00000400,
  1'd1,  5'd13, 27'h00000094, 5'd24, 27'h000003c1, 5'd8, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000010d, 5'd25, 27'h0000001f, 5'd16, 27'h000003ea, 32'h00000400,
  1'd1,  5'd14, 27'h000001fc, 5'd23, 27'h00000338, 5'd27, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000fc, 5'd4, 27'h0000011b, 5'd7, 27'h000002a4, 32'h00000400,
  1'd1,  5'd24, 27'h00000217, 5'd2, 27'h000003ff, 5'd17, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000271, 5'd0, 27'h000003f6, 5'd27, 27'h0000018b, 32'h00000400,
  1'd1,  5'd25, 27'h000002c7, 5'd11, 27'h00000086, 5'd9, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000121, 5'd10, 27'h00000199, 5'd18, 27'h0000025c, 32'h00000400,
  1'd1,  5'd20, 27'h000002c6, 5'd14, 27'h000001a1, 5'd30, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000c5, 5'd22, 27'h0000028c, 5'd9, 27'h0000012c, 32'h00000400,
  1'd1,  5'd21, 27'h00000117, 5'd23, 27'h00000137, 5'd20, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000ba, 5'd22, 27'h000001e1, 5'd28, 27'h000003fd, 32'h00000400,
  1'd1,  5'd4, 27'h000000ed, 5'd6, 27'h000003e0, 5'd0, 27'h000003ee, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000199, 5'd6, 27'h000001e4, 5'd11, 27'h000003a6, 32'h00000400,
  1'd1,  5'd4, 27'h000003d7, 5'd7, 27'h000000b9, 5'd22, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000003a, 5'd20, 27'h00000250, 5'd4, 27'h000003f1, 32'h00000400,
  1'd1,  5'd3, 27'h000000f8, 5'd16, 27'h0000000b, 5'd13, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000004, 5'd15, 27'h0000021b, 5'd22, 27'h00000114, 32'h00000400,
  1'd1,  5'd0, 27'h00000344, 5'd26, 27'h000002eb, 5'd2, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003fa, 5'd30, 27'h0000032b, 5'd11, 27'h00000161, 32'h00000400,
  1'd1,  5'd3, 27'h00000175, 5'd27, 27'h000001e3, 5'd24, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002be, 5'd5, 27'h000001e5, 5'd1, 27'h000002ce, 32'h00000400,
  1'd1,  5'd11, 27'h0000000b, 5'd6, 27'h0000031a, 5'd13, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000108, 5'd5, 27'h000001dc, 5'd24, 27'h0000014a, 32'h00000400,
  1'd1,  5'd15, 27'h000001c3, 5'd18, 27'h0000012f, 5'd1, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000208, 5'd18, 27'h0000024d, 5'd14, 27'h000002ab, 32'h00000400,
  1'd1,  5'd11, 27'h0000007b, 5'd16, 27'h000001d2, 5'd24, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002a9, 5'd30, 27'h0000031f, 5'd2, 27'h000002a8, 32'h00000400,
  1'd1,  5'd14, 27'h000001e2, 5'd28, 27'h00000228, 5'd11, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000078, 5'd30, 27'h00000050, 5'd24, 27'h00000098, 32'h00000400,
  1'd1,  5'd24, 27'h00000272, 5'd8, 27'h000001b8, 5'd4, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006c, 5'd9, 27'h00000178, 5'd11, 27'h000003d3, 32'h00000400,
  1'd1,  5'd21, 27'h0000012a, 5'd8, 27'h00000198, 5'd25, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000017, 5'd19, 27'h000002a1, 5'd1, 27'h00000105, 32'h00000400,
  1'd1,  5'd25, 27'h00000335, 5'd15, 27'h00000295, 5'd11, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000008, 5'd19, 27'h000003c7, 5'd23, 27'h0000020e, 32'h00000400,
  1'd1,  5'd23, 27'h00000373, 5'd26, 27'h000001c4, 5'd5, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000052, 5'd29, 27'h000002cc, 5'd13, 27'h0000008c, 32'h00000400,
  1'd1,  5'd23, 27'h00000368, 5'd26, 27'h0000019a, 5'd20, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002ba, 5'd6, 27'h000001c8, 5'd6, 27'h00000039, 32'h00000400,
  1'd1,  5'd4, 27'h00000347, 5'd7, 27'h00000200, 5'd17, 27'h000002a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000216, 5'd5, 27'h000002a0, 5'd28, 27'h00000167, 32'h00000400,
  1'd1,  5'd3, 27'h0000003d, 5'd17, 27'h00000164, 5'd7, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000019, 5'd17, 27'h000002d6, 5'd19, 27'h00000309, 32'h00000400,
  1'd1,  5'd4, 27'h000001cb, 5'd15, 27'h00000353, 5'd30, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003eb, 5'd26, 27'h000002b6, 5'd6, 27'h00000170, 32'h00000400,
  1'd1,  5'd1, 27'h00000078, 5'd26, 27'h000000e7, 5'd18, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f1, 5'd28, 27'h00000300, 5'd29, 27'h00000395, 32'h00000400,
  1'd1,  5'd12, 27'h00000317, 5'd8, 27'h0000038f, 5'd7, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000112, 5'd7, 27'h00000174, 5'd17, 27'h000000f8, 32'h00000400,
  1'd1,  5'd15, 27'h000000a7, 5'd9, 27'h000001de, 5'd29, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000a9, 5'd20, 27'h000000c6, 5'd9, 27'h000001ea, 32'h00000400,
  1'd1,  5'd12, 27'h00000225, 5'd15, 27'h00000264, 5'd19, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000223, 5'd19, 27'h000001ac, 5'd29, 27'h0000021c, 32'h00000400,
  1'd1,  5'd11, 27'h000003dd, 5'd30, 27'h0000031d, 5'd7, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000255, 5'd26, 27'h000003d1, 5'd18, 27'h0000011b, 32'h00000400,
  1'd1,  5'd12, 27'h0000030a, 5'd28, 27'h00000322, 5'd29, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000219, 5'd7, 27'h000001b3, 5'd8, 27'h000000d2, 32'h00000400,
  1'd1,  5'd25, 27'h0000021b, 5'd9, 27'h000002b1, 5'd18, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000319, 5'd9, 27'h000001f7, 5'd29, 27'h0000007e, 32'h00000400,
  1'd1,  5'd21, 27'h000001a5, 5'd18, 27'h0000027e, 5'd7, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000008, 5'd18, 27'h00000353, 5'd16, 27'h0000006c, 32'h00000400,
  1'd1,  5'd25, 27'h000002fd, 5'd18, 27'h000002ef, 5'd30, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000326, 5'd30, 27'h00000147, 5'd5, 27'h0000029d, 32'h00000400,
  1'd1,  5'd21, 27'h000002ca, 5'd28, 27'h000000ac, 5'd17, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000333, 5'd27, 27'h00000049, 5'd29, 27'h0000035d, 32'h00000400,
  1'd1,  5'd8, 27'h00000326, 5'd2, 27'h000001a1, 5'd7, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000184, 5'd2, 27'h00000020, 5'd18, 27'h0000013a, 32'h00000400,
  1'd1,  5'd5, 27'h000003bf, 5'd2, 27'h00000102, 5'd29, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003d5, 5'd12, 27'h00000002, 5'd1, 27'h000000f3, 32'h00000400,
  1'd1,  5'd6, 27'h000002c9, 5'd14, 27'h00000343, 5'd12, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009a, 5'd11, 27'h00000271, 5'd22, 27'h0000005e, 32'h00000400,
  1'd1,  5'd9, 27'h000002dd, 5'd24, 27'h0000003b, 5'd2, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001e4, 5'd25, 27'h0000006f, 5'd10, 27'h000002a6, 32'h00000400,
  1'd1,  5'd6, 27'h0000001f, 5'd22, 27'h000001cc, 5'd21, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000009b, 5'd2, 27'h000000d9, 5'd7, 27'h000003c2, 32'h00000400,
  1'd1,  5'd17, 27'h000000de, 5'd0, 27'h000003bc, 5'd18, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000215, 5'd1, 27'h000000b4, 5'd26, 27'h000001a3, 32'h00000400,
  1'd1,  5'd17, 27'h0000032b, 5'd10, 27'h0000030f, 5'd0, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000241, 5'd10, 27'h00000399, 5'd10, 27'h000001e2, 32'h00000400,
  1'd1,  5'd16, 27'h00000376, 5'd13, 27'h00000324, 5'd25, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d3, 5'd22, 27'h0000002b, 5'd3, 27'h0000028d, 32'h00000400,
  1'd1,  5'd17, 27'h0000027d, 5'd25, 27'h00000149, 5'd11, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e8, 5'd22, 27'h0000020c, 5'd24, 27'h00000337, 32'h00000400,
  1'd1,  5'd26, 27'h0000001a, 5'd1, 27'h000002dd, 5'd4, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000112, 5'd2, 27'h00000022, 5'd12, 27'h000002f7, 32'h00000400,
  1'd1,  5'd27, 27'h000002a9, 5'd1, 27'h00000287, 5'd24, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001bc, 5'd11, 27'h000003a4, 5'd2, 27'h0000026f, 32'h00000400,
  1'd1,  5'd29, 27'h00000357, 5'd12, 27'h00000379, 5'd11, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000248, 5'd12, 27'h0000031e, 5'd23, 27'h00000068, 32'h00000400,
  1'd1,  5'd28, 27'h00000350, 5'd25, 27'h000001da, 5'd0, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000271, 5'd25, 27'h00000327, 5'd11, 27'h00000150, 32'h00000400,
  1'd1,  5'd26, 27'h000000f8, 5'd21, 27'h000000d2, 5'd24, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000035f, 5'd1, 27'h00000378, 5'd1, 27'h00000062, 32'h00000400,
  1'd1,  5'd5, 27'h0000023f, 5'd5, 27'h0000006b, 5'd11, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b9, 5'd2, 27'h00000105, 5'd20, 27'h0000030a, 32'h00000400,
  1'd1,  5'd10, 27'h0000013e, 5'd11, 27'h000002ba, 5'd6, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000068, 5'd11, 27'h00000006, 5'd16, 27'h00000015, 32'h00000400,
  1'd1,  5'd7, 27'h000002f8, 5'd13, 27'h000002ae, 5'd30, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000000c, 5'd24, 27'h000001c5, 5'd8, 27'h000003ee, 32'h00000400,
  1'd1,  5'd9, 27'h0000033a, 5'd22, 27'h000002f9, 5'd15, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003fb, 5'd21, 27'h00000178, 5'd30, 27'h000001eb, 32'h00000400,
  1'd1,  5'd17, 27'h00000221, 5'd0, 27'h000003f4, 5'd4, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000011, 5'd1, 27'h000001b2, 5'd11, 27'h000003ea, 32'h00000400,
  1'd1,  5'd19, 27'h000001c6, 5'd4, 27'h0000002d, 5'd23, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000029, 5'd14, 27'h000003a9, 5'd9, 27'h000000b3, 32'h00000400,
  1'd1,  5'd17, 27'h000000f0, 5'd12, 27'h0000038e, 5'd16, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000117, 5'd11, 27'h000001b0, 5'd30, 27'h00000293, 32'h00000400,
  1'd1,  5'd19, 27'h00000068, 5'd23, 27'h000000ac, 5'd8, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000296, 5'd21, 27'h00000092, 5'd18, 27'h0000022c, 32'h00000400,
  1'd1,  5'd16, 27'h0000012c, 5'd23, 27'h0000000a, 5'd27, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000211, 5'd1, 27'h000002ba, 5'd6, 27'h00000129, 32'h00000400,
  1'd1,  5'd28, 27'h000000b5, 5'd1, 27'h00000235, 5'd16, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b1, 5'd1, 27'h000001b9, 5'd25, 27'h000003e2, 32'h00000400,
  1'd1,  5'd28, 27'h000003c8, 5'd11, 27'h0000002a, 5'd5, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000129, 5'd12, 27'h000002d1, 5'd18, 27'h000001f4, 32'h00000400,
  1'd1,  5'd30, 27'h0000012e, 5'd11, 27'h000000bb, 5'd30, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000156, 5'd23, 27'h0000013e, 5'd8, 27'h00000213, 32'h00000400,
  1'd1,  5'd29, 27'h000000a4, 5'd21, 27'h000000fc, 5'd18, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003d6, 5'd25, 27'h00000301, 5'd29, 27'h0000014b, 32'h00000400,
  1'd1,  5'd10, 27'h000000be, 5'd7, 27'h00000164, 5'd0, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000361, 5'd6, 27'h000000db, 5'd15, 27'h00000059, 32'h00000400,
  1'd1,  5'd7, 27'h000003c8, 5'd6, 27'h0000035b, 5'd22, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000022e, 5'd20, 27'h0000025b, 5'd4, 27'h00000305, 32'h00000400,
  1'd1,  5'd5, 27'h00000328, 5'd17, 27'h0000024a, 5'd14, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000339, 5'd18, 27'h000001c0, 5'd23, 27'h000002a7, 32'h00000400,
  1'd1,  5'd6, 27'h000002ab, 5'd30, 27'h000001e0, 5'd1, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000012f, 5'd29, 27'h00000224, 5'd11, 27'h000003d8, 32'h00000400,
  1'd1,  5'd6, 27'h0000013e, 5'd28, 27'h000000e7, 5'd25, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000241, 5'd5, 27'h00000365, 5'd0, 27'h000002d1, 32'h00000400,
  1'd1,  5'd18, 27'h00000108, 5'd9, 27'h00000256, 5'd12, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000f1, 5'd7, 27'h000000ae, 5'd23, 27'h000001dc, 32'h00000400,
  1'd1,  5'd19, 27'h000000f8, 5'd18, 27'h00000003, 5'd0, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c2, 5'd18, 27'h000003ec, 5'd10, 27'h00000319, 32'h00000400,
  1'd1,  5'd19, 27'h00000085, 5'd16, 27'h0000005a, 5'd23, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000011b, 5'd27, 27'h00000202, 5'd0, 27'h000001ec, 32'h00000400,
  1'd1,  5'd17, 27'h000003cf, 5'd27, 27'h0000023d, 5'd13, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000141, 5'd28, 27'h000003ce, 5'd21, 27'h000002dd, 32'h00000400,
  1'd1,  5'd28, 27'h00000097, 5'd7, 27'h000000e8, 5'd0, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000209, 5'd6, 27'h0000028e, 5'd10, 27'h00000283, 32'h00000400,
  1'd1,  5'd30, 27'h00000094, 5'd9, 27'h0000027f, 5'd21, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000026a, 5'd16, 27'h000003cc, 5'd2, 27'h00000092, 32'h00000400,
  1'd1,  5'd27, 27'h00000238, 5'd19, 27'h0000038b, 5'd13, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000394, 5'd16, 27'h0000025a, 5'd21, 27'h000003d5, 32'h00000400,
  1'd1,  5'd26, 27'h0000020e, 5'd28, 27'h00000183, 5'd3, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001af, 5'd27, 27'h0000023e, 5'd13, 27'h0000019a, 32'h00000400,
  1'd1,  5'd25, 27'h00000386, 5'd28, 27'h00000371, 5'd24, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000061, 5'd5, 27'h000000d3, 5'd7, 27'h0000014e, 32'h00000400,
  1'd1,  5'd10, 27'h00000002, 5'd6, 27'h000003ff, 5'd16, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000d0, 5'd10, 27'h00000040, 5'd29, 27'h0000015c, 32'h00000400,
  1'd1,  5'd6, 27'h00000214, 5'd16, 27'h00000400, 5'd10, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002e2, 5'd18, 27'h0000020c, 5'd16, 27'h000001b3, 32'h00000400,
  1'd1,  5'd8, 27'h000000e5, 5'd19, 27'h00000112, 5'd30, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000322, 5'd30, 27'h0000024f, 5'd10, 27'h0000012b, 32'h00000400,
  1'd1,  5'd8, 27'h0000001a, 5'd28, 27'h00000004, 5'd19, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000cd, 5'd27, 27'h00000148, 5'd28, 27'h000000eb, 32'h00000400,
  1'd1,  5'd18, 27'h00000285, 5'd9, 27'h00000077, 5'd9, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000287, 5'd9, 27'h00000142, 5'd15, 27'h000002e6, 32'h00000400,
  1'd1,  5'd17, 27'h000001ca, 5'd5, 27'h00000284, 5'd30, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b2, 5'd15, 27'h0000030e, 5'd5, 27'h0000018e, 32'h00000400,
  1'd1,  5'd15, 27'h000002dd, 5'd17, 27'h00000275, 5'd18, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000362, 5'd18, 27'h00000341, 5'd29, 27'h000000f6, 32'h00000400,
  1'd1,  5'd16, 27'h00000053, 5'd29, 27'h000003d5, 5'd7, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000009e, 5'd30, 27'h000001d9, 5'd16, 27'h0000006d, 32'h00000400,
  1'd1,  5'd17, 27'h000000f1, 5'd29, 27'h00000137, 5'd28, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c1, 5'd5, 27'h000002b7, 5'd5, 27'h00000207, 32'h00000400,
  1'd1,  5'd26, 27'h00000155, 5'd9, 27'h000002f3, 5'd19, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000035f, 5'd5, 27'h0000022d, 5'd28, 27'h00000276, 32'h00000400,
  1'd1,  5'd30, 27'h00000124, 5'd17, 27'h00000319, 5'd6, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000299, 5'd16, 27'h00000193, 5'd18, 27'h000001fa, 32'h00000400,
  1'd1,  5'd26, 27'h000001f7, 5'd16, 27'h0000009b, 5'd28, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000014, 5'd26, 27'h0000010b, 5'd7, 27'h0000023c, 32'h00000400,
  1'd1,  5'd30, 27'h000001f3, 5'd28, 27'h00000249, 5'd19, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a4, 5'd28, 27'h000000cf, 5'd29, 27'h0000020c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h0000021a, 5'd0, 27'h000000a2, 5'd3, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000007c, 5'd2, 27'h000002fa, 5'd15, 27'h000000d8, 32'h00000400,
  1'd1,  5'd2, 27'h00000100, 5'd2, 27'h00000301, 5'd22, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000191, 5'd11, 27'h0000035c, 5'd0, 27'h0000015c, 32'h00000400,
  1'd1,  5'd2, 27'h00000114, 5'd13, 27'h0000016e, 5'd12, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002b4, 5'd10, 27'h00000365, 5'd24, 27'h000003c3, 32'h00000400,
  1'd1,  5'd3, 27'h0000033c, 5'd21, 27'h0000022b, 5'd4, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f6, 5'd23, 27'h00000037, 5'd15, 27'h0000005d, 32'h00000400,
  1'd1,  5'd0, 27'h00000007, 5'd21, 27'h00000244, 5'd24, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000201, 5'd1, 27'h0000032a, 5'd2, 27'h000001ca, 32'h00000400,
  1'd1,  5'd13, 27'h000000e3, 5'd3, 27'h00000304, 5'd11, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000000, 5'd2, 27'h000002df, 5'd24, 27'h0000016e, 32'h00000400,
  1'd1,  5'd10, 27'h00000287, 5'd12, 27'h000001bf, 5'd0, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000241, 5'd10, 27'h0000035d, 5'd15, 27'h000000f5, 32'h00000400,
  1'd1,  5'd11, 27'h00000015, 5'd12, 27'h000002ab, 5'd20, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000b9, 5'd21, 27'h000000d4, 5'd1, 27'h000001f6, 32'h00000400,
  1'd1,  5'd13, 27'h0000026e, 5'd23, 27'h00000090, 5'd12, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001dd, 5'd23, 27'h000003a8, 5'd24, 27'h000000d4, 32'h00000400,
  1'd1,  5'd23, 27'h0000018f, 5'd2, 27'h00000348, 5'd2, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000012d, 5'd4, 27'h000001a1, 5'd12, 27'h00000154, 32'h00000400,
  1'd1,  5'd25, 27'h0000010a, 5'd3, 27'h000001cf, 5'd22, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c8, 5'd10, 27'h000002da, 5'd4, 27'h00000169, 32'h00000400,
  1'd1,  5'd23, 27'h000003b2, 5'd12, 27'h00000113, 5'd10, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d2, 5'd13, 27'h00000036, 5'd25, 27'h00000168, 32'h00000400,
  1'd1,  5'd24, 27'h00000123, 5'd22, 27'h0000002f, 5'd3, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002f2, 5'd21, 27'h00000103, 5'd12, 27'h000001ea, 32'h00000400,
  1'd1,  5'd22, 27'h00000071, 5'd24, 27'h00000151, 5'd23, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002a1, 5'd1, 27'h000002b9, 5'd8, 27'h00000312, 32'h00000400,
  1'd1,  5'd0, 27'h0000019e, 5'd0, 27'h00000344, 5'd15, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a0, 5'd4, 27'h000003a2, 5'd28, 27'h000003b7, 32'h00000400,
  1'd1,  5'd3, 27'h000003cf, 5'd14, 27'h000002cf, 5'd7, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000bb, 5'd15, 27'h00000033, 5'd19, 27'h00000315, 32'h00000400,
  1'd1,  5'd3, 27'h000001ac, 5'd12, 27'h00000091, 5'd27, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000221, 5'd21, 27'h000001bb, 5'd8, 27'h00000279, 32'h00000400,
  1'd1,  5'd0, 27'h00000106, 5'd24, 27'h000001be, 5'd20, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000165, 5'd20, 27'h0000030c, 5'd30, 27'h000001d1, 32'h00000400,
  1'd1,  5'd12, 27'h0000012c, 5'd1, 27'h0000013d, 5'd10, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000019c, 5'd0, 27'h000000e3, 5'd19, 27'h0000034f, 32'h00000400,
  1'd1,  5'd13, 27'h00000041, 5'd0, 27'h0000006b, 5'd29, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000017e, 5'd10, 27'h0000032d, 5'd6, 27'h000001e1, 32'h00000400,
  1'd1,  5'd13, 27'h000002dc, 5'd14, 27'h000000cb, 5'd17, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000378, 5'd12, 27'h00000334, 5'd30, 27'h000000bb, 32'h00000400,
  1'd1,  5'd13, 27'h0000002b, 5'd23, 27'h000003c5, 5'd7, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000a6, 5'd22, 27'h0000021c, 5'd18, 27'h000000ae, 32'h00000400,
  1'd1,  5'd13, 27'h00000114, 5'd23, 27'h0000027d, 5'd29, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000062, 5'd3, 27'h0000021e, 5'd9, 27'h00000097, 32'h00000400,
  1'd1,  5'd23, 27'h000000eb, 5'd0, 27'h000002de, 5'd18, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000136, 5'd4, 27'h000002e2, 5'd26, 27'h00000060, 32'h00000400,
  1'd1,  5'd25, 27'h00000099, 5'd14, 27'h0000016a, 5'd6, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ed, 5'd14, 27'h00000260, 5'd15, 27'h000002a6, 32'h00000400,
  1'd1,  5'd21, 27'h000002da, 5'd12, 27'h000001d3, 5'd29, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000003b, 5'd21, 27'h000003ab, 5'd7, 27'h0000020f, 32'h00000400,
  1'd1,  5'd21, 27'h000003ea, 5'd23, 27'h000002e5, 5'd17, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000016c, 5'd23, 27'h00000294, 5'd27, 27'h000000d7, 32'h00000400,
  1'd1,  5'd4, 27'h000003d0, 5'd8, 27'h0000039b, 5'd1, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000006b, 5'd6, 27'h000003c3, 5'd10, 27'h00000377, 32'h00000400,
  1'd1,  5'd1, 27'h000002ec, 5'd8, 27'h00000061, 5'd24, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c6, 5'd19, 27'h000002f3, 5'd2, 27'h00000385, 32'h00000400,
  1'd1,  5'd0, 27'h0000023d, 5'd19, 27'h00000224, 5'd15, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027c, 5'd18, 27'h00000218, 5'd23, 27'h0000003a, 32'h00000400,
  1'd1,  5'd5, 27'h00000037, 5'd26, 27'h00000373, 5'd2, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000100, 5'd29, 27'h00000354, 5'd15, 27'h00000028, 32'h00000400,
  1'd1,  5'd0, 27'h0000014a, 5'd26, 27'h00000348, 5'd21, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000362, 5'd8, 27'h00000126, 5'd0, 27'h000003a8, 32'h00000400,
  1'd1,  5'd11, 27'h000002d9, 5'd5, 27'h00000235, 5'd10, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000009a, 5'd10, 27'h0000000c, 5'd23, 27'h000000a0, 32'h00000400,
  1'd1,  5'd14, 27'h000003e6, 5'd16, 27'h00000047, 5'd4, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d8, 5'd18, 27'h0000008a, 5'd12, 27'h000002fc, 32'h00000400,
  1'd1,  5'd14, 27'h00000223, 5'd18, 27'h00000213, 5'd24, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000187, 5'd28, 27'h00000184, 5'd0, 27'h00000092, 32'h00000400,
  1'd1,  5'd12, 27'h0000031f, 5'd28, 27'h00000140, 5'd12, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000e4, 5'd27, 27'h0000007d, 5'd22, 27'h0000011b, 32'h00000400,
  1'd1,  5'd25, 27'h0000008e, 5'd7, 27'h000001d2, 5'd2, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000168, 5'd8, 27'h000000cc, 5'd15, 27'h000000bd, 32'h00000400,
  1'd1,  5'd25, 27'h00000096, 5'd7, 27'h00000122, 5'd22, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000081, 5'd19, 27'h0000021e, 5'd0, 27'h000003df, 32'h00000400,
  1'd1,  5'd22, 27'h00000275, 5'd17, 27'h000002bc, 5'd14, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000162, 5'd17, 27'h0000032f, 5'd20, 27'h00000324, 32'h00000400,
  1'd1,  5'd23, 27'h0000016c, 5'd26, 27'h00000148, 5'd0, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000065, 5'd29, 27'h00000137, 5'd15, 27'h000000c1, 32'h00000400,
  1'd1,  5'd24, 27'h0000010d, 5'd27, 27'h000001a5, 5'd25, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000027b, 5'd6, 27'h00000021, 5'd9, 27'h000002ca, 32'h00000400,
  1'd1,  5'd3, 27'h00000114, 5'd9, 27'h0000004c, 5'd19, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d9, 5'd9, 27'h00000021, 5'd29, 27'h00000017, 32'h00000400,
  1'd1,  5'd1, 27'h000001de, 5'd18, 27'h00000344, 5'd8, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000010a, 5'd15, 27'h00000292, 5'd17, 27'h0000031f, 32'h00000400,
  1'd1,  5'd4, 27'h000003c5, 5'd19, 27'h000003c5, 5'd26, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000397, 5'd29, 27'h000002d4, 5'd10, 27'h00000023, 32'h00000400,
  1'd1,  5'd2, 27'h00000064, 5'd29, 27'h000000c3, 5'd15, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000227, 5'd30, 27'h000002c9, 5'd30, 27'h00000159, 32'h00000400,
  1'd1,  5'd12, 27'h00000157, 5'd10, 27'h00000110, 5'd5, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f1, 5'd6, 27'h0000001a, 5'd20, 27'h0000004f, 32'h00000400,
  1'd1,  5'd11, 27'h00000283, 5'd7, 27'h00000361, 5'd30, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000229, 5'd18, 27'h00000002, 5'd7, 27'h0000036e, 32'h00000400,
  1'd1,  5'd13, 27'h00000274, 5'd16, 27'h00000304, 5'd20, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000378, 5'd17, 27'h000002c9, 5'd26, 27'h000001cd, 32'h00000400,
  1'd1,  5'd10, 27'h000001b7, 5'd26, 27'h000002af, 5'd7, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fe, 5'd30, 27'h000002f0, 5'd17, 27'h000003d8, 32'h00000400,
  1'd1,  5'd13, 27'h000001db, 5'd30, 27'h00000194, 5'd27, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000299, 5'd10, 27'h00000093, 5'd8, 27'h000002c3, 32'h00000400,
  1'd1,  5'd24, 27'h000000d1, 5'd7, 27'h00000168, 5'd18, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000023c, 5'd10, 27'h00000122, 5'd26, 27'h00000354, 32'h00000400,
  1'd1,  5'd22, 27'h00000320, 5'd16, 27'h00000129, 5'd8, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000388, 5'd17, 27'h00000385, 5'd16, 27'h00000099, 32'h00000400,
  1'd1,  5'd23, 27'h000000b8, 5'd15, 27'h000002ed, 5'd28, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fe, 5'd27, 27'h00000170, 5'd6, 27'h000001c1, 32'h00000400,
  1'd1,  5'd23, 27'h00000090, 5'd29, 27'h00000164, 5'd19, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000005, 5'd27, 27'h0000001e, 5'd30, 27'h0000039e, 32'h00000400,
  1'd1,  5'd8, 27'h00000056, 5'd4, 27'h000003c3, 5'd8, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ee, 5'd4, 27'h00000080, 5'd16, 27'h000001d2, 32'h00000400,
  1'd1,  5'd9, 27'h00000136, 5'd1, 27'h00000034, 5'd27, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000025d, 5'd11, 27'h000003c0, 5'd5, 27'h000000aa, 32'h00000400,
  1'd1,  5'd9, 27'h00000302, 5'd11, 27'h00000071, 5'd13, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003fb, 5'd13, 27'h000000ee, 5'd23, 27'h0000002e, 32'h00000400,
  1'd1,  5'd10, 27'h00000135, 5'd22, 27'h0000026d, 5'd2, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007c, 5'd24, 27'h0000015e, 5'd13, 27'h00000118, 32'h00000400,
  1'd1,  5'd7, 27'h000002b1, 5'd21, 27'h0000027b, 5'd20, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000dc, 5'd2, 27'h00000381, 5'd8, 27'h00000331, 32'h00000400,
  1'd1,  5'd18, 27'h000000dc, 5'd0, 27'h0000037d, 5'd17, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000338, 5'd3, 27'h0000011f, 5'd28, 27'h0000001f, 32'h00000400,
  1'd1,  5'd20, 27'h00000090, 5'd13, 27'h00000189, 5'd0, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d9, 5'd11, 27'h000003a4, 5'd12, 27'h00000272, 32'h00000400,
  1'd1,  5'd15, 27'h00000280, 5'd11, 27'h000002aa, 5'd24, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000288, 5'd22, 27'h000001d3, 5'd4, 27'h0000004d, 32'h00000400,
  1'd1,  5'd19, 27'h00000385, 5'd24, 27'h00000218, 5'd12, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000027, 5'd23, 27'h00000242, 5'd20, 27'h000003bb, 32'h00000400,
  1'd1,  5'd28, 27'h000000de, 5'd4, 27'h00000015, 5'd4, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003df, 5'd1, 27'h00000162, 5'd14, 27'h000001e7, 32'h00000400,
  1'd1,  5'd27, 27'h000000aa, 5'd1, 27'h000001bd, 5'd23, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000065, 5'd15, 27'h00000066, 5'd4, 27'h000003c5, 32'h00000400,
  1'd1,  5'd27, 27'h000002e1, 5'd12, 27'h00000196, 5'd14, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000031d, 5'd14, 27'h00000288, 5'd22, 27'h00000263, 32'h00000400,
  1'd1,  5'd26, 27'h0000011f, 5'd20, 27'h00000375, 5'd3, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000306, 5'd23, 27'h00000098, 5'd13, 27'h0000024f, 32'h00000400,
  1'd1,  5'd28, 27'h00000220, 5'd24, 27'h000002e4, 5'd24, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000036c, 5'd2, 27'h0000030b, 5'd3, 27'h00000217, 32'h00000400,
  1'd1,  5'd8, 27'h000001da, 5'd3, 27'h00000297, 5'd12, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003db, 5'd2, 27'h00000243, 5'd24, 27'h00000374, 32'h00000400,
  1'd1,  5'd6, 27'h000000bf, 5'd11, 27'h00000302, 5'd6, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e8, 5'd13, 27'h00000395, 5'd18, 27'h0000019c, 32'h00000400,
  1'd1,  5'd5, 27'h000002e8, 5'd11, 27'h00000247, 5'd27, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000023f, 5'd23, 27'h000000f4, 5'd7, 27'h00000313, 32'h00000400,
  1'd1,  5'd8, 27'h0000016c, 5'd23, 27'h000001b0, 5'd17, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000022, 5'd24, 27'h00000312, 5'd29, 27'h00000233, 32'h00000400,
  1'd1,  5'd15, 27'h0000027d, 5'd3, 27'h00000179, 5'd2, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000007e, 5'd2, 27'h000003ae, 5'd14, 27'h0000016e, 32'h00000400,
  1'd1,  5'd15, 27'h00000310, 5'd2, 27'h000001f5, 5'd22, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000291, 5'd14, 27'h000001da, 5'd7, 27'h000001be, 32'h00000400,
  1'd1,  5'd16, 27'h000003f1, 5'd10, 27'h0000022c, 5'd19, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000106, 5'd12, 27'h000002e0, 5'd30, 27'h000001dc, 32'h00000400,
  1'd1,  5'd18, 27'h0000028d, 5'd22, 27'h0000036a, 5'd9, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000038, 5'd24, 27'h0000033d, 5'd18, 27'h000003e3, 32'h00000400,
  1'd1,  5'd16, 27'h000003d1, 5'd23, 27'h00000273, 5'd28, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003d0, 5'd4, 27'h00000077, 5'd6, 27'h000001d3, 32'h00000400,
  1'd1,  5'd29, 27'h00000036, 5'd4, 27'h0000005a, 5'd18, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000034b, 5'd1, 27'h00000189, 5'd26, 27'h000002ce, 32'h00000400,
  1'd1,  5'd27, 27'h0000012f, 5'd13, 27'h00000386, 5'd8, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000b0, 5'd11, 27'h00000384, 5'd16, 27'h000001bd, 32'h00000400,
  1'd1,  5'd29, 27'h0000009b, 5'd12, 27'h000001f0, 5'd26, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001f, 5'd23, 27'h000001a4, 5'd10, 27'h0000000c, 32'h00000400,
  1'd1,  5'd28, 27'h00000244, 5'd25, 27'h0000006e, 5'd20, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ef, 5'd21, 27'h00000244, 5'd26, 27'h00000392, 32'h00000400,
  1'd1,  5'd5, 27'h000002c0, 5'd7, 27'h0000035b, 5'd4, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000042, 5'd7, 27'h00000036, 5'd12, 27'h0000016d, 32'h00000400,
  1'd1,  5'd7, 27'h00000323, 5'd7, 27'h00000322, 5'd23, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000024c, 5'd19, 27'h0000015e, 5'd4, 27'h000002df, 32'h00000400,
  1'd1,  5'd7, 27'h00000003, 5'd16, 27'h0000018e, 5'd15, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000031b, 5'd18, 27'h000000ac, 5'd25, 27'h00000050, 32'h00000400,
  1'd1,  5'd9, 27'h00000245, 5'd28, 27'h0000010a, 5'd0, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000f8, 5'd28, 27'h00000397, 5'd12, 27'h0000024c, 32'h00000400,
  1'd1,  5'd8, 27'h000003d8, 5'd27, 27'h0000005f, 5'd25, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e2, 5'd6, 27'h000003f4, 5'd3, 27'h000000db, 32'h00000400,
  1'd1,  5'd17, 27'h000003a4, 5'd9, 27'h000003c3, 5'd11, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c9, 5'd7, 27'h00000041, 5'd24, 27'h0000025e, 32'h00000400,
  1'd1,  5'd17, 27'h00000209, 5'd19, 27'h000003fe, 5'd1, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001f9, 5'd17, 27'h0000016c, 5'd15, 27'h000000b5, 32'h00000400,
  1'd1,  5'd15, 27'h00000225, 5'd18, 27'h00000230, 5'd25, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002b1, 5'd28, 27'h00000351, 5'd1, 27'h000002a6, 32'h00000400,
  1'd1,  5'd20, 27'h00000025, 5'd30, 27'h000000a1, 5'd15, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000012, 5'd30, 27'h000003f7, 5'd22, 27'h000003ea, 32'h00000400,
  1'd1,  5'd30, 27'h00000360, 5'd5, 27'h000002cf, 5'd4, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000031c, 5'd10, 27'h0000012c, 5'd15, 27'h000000b5, 32'h00000400,
  1'd1,  5'd29, 27'h00000116, 5'd5, 27'h000000ea, 5'd23, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000282, 5'd20, 27'h000000fb, 5'd3, 27'h000003d1, 32'h00000400,
  1'd1,  5'd27, 27'h00000154, 5'd20, 27'h00000108, 5'd11, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000362, 5'd17, 27'h000002c3, 5'd21, 27'h000001c1, 32'h00000400,
  1'd1,  5'd28, 27'h00000050, 5'd27, 27'h000002b8, 5'd1, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002a3, 5'd26, 27'h000002b0, 5'd11, 27'h000000f2, 32'h00000400,
  1'd1,  5'd26, 27'h00000249, 5'd26, 27'h000001e8, 5'd20, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000225, 5'd7, 27'h00000006, 5'd9, 27'h00000124, 32'h00000400,
  1'd1,  5'd8, 27'h000000f3, 5'd5, 27'h00000354, 5'd18, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000008e, 5'd5, 27'h000000c7, 5'd26, 27'h0000031f, 32'h00000400,
  1'd1,  5'd5, 27'h00000224, 5'd16, 27'h00000022, 5'd7, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000019e, 5'd18, 27'h00000341, 5'd18, 27'h00000000, 32'h00000400,
  1'd1,  5'd6, 27'h000000b4, 5'd20, 27'h000000fc, 5'd30, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000030c, 5'd30, 27'h000003d5, 5'd7, 27'h000000ec, 32'h00000400,
  1'd1,  5'd8, 27'h000001aa, 5'd26, 27'h00000101, 5'd18, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c0, 5'd27, 27'h00000323, 5'd26, 27'h000000c6, 32'h00000400,
  1'd1,  5'd16, 27'h000000a4, 5'd7, 27'h000000f2, 5'd7, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000359, 5'd6, 27'h000001bb, 5'd18, 27'h0000012d, 32'h00000400,
  1'd1,  5'd17, 27'h000000a0, 5'd6, 27'h00000038, 5'd28, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000383, 5'd20, 27'h0000028b, 5'd8, 27'h0000039e, 32'h00000400,
  1'd1,  5'd18, 27'h000003c0, 5'd19, 27'h000000e4, 5'd19, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002e3, 5'd20, 27'h00000115, 5'd30, 27'h000002f1, 32'h00000400,
  1'd1,  5'd17, 27'h00000210, 5'd29, 27'h0000033c, 5'd6, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000207, 5'd30, 27'h00000254, 5'd19, 27'h000002fe, 32'h00000400,
  1'd1,  5'd18, 27'h0000008b, 5'd28, 27'h00000211, 5'd26, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001a1, 5'd9, 27'h000000c8, 5'd10, 27'h0000008c, 32'h00000400,
  1'd1,  5'd28, 27'h000000a9, 5'd8, 27'h0000038e, 5'd19, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000154, 5'd8, 27'h0000000c, 5'd27, 27'h0000025e, 32'h00000400,
  1'd1,  5'd28, 27'h00000011, 5'd17, 27'h00000015, 5'd9, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000003f, 5'd17, 27'h00000120, 5'd18, 27'h0000028d, 32'h00000400,
  1'd1,  5'd30, 27'h000002ab, 5'd16, 27'h00000171, 5'd29, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ad, 5'd28, 27'h00000301, 5'd9, 27'h0000010f, 32'h00000400,
  1'd1,  5'd28, 27'h0000011e, 5'd27, 27'h000000bc, 5'd20, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b7, 5'd27, 27'h00000165, 5'd26, 27'h000001eb, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000025, 5'd3, 27'h0000026b, 5'd3, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000a1, 5'd4, 27'h0000026f, 5'd15, 27'h0000014e, 32'h00000400,
  1'd1,  5'd1, 27'h0000009f, 5'd0, 27'h00000102, 5'd24, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002a1, 5'd13, 27'h000000ef, 5'd0, 27'h000003ef, 32'h00000400,
  1'd1,  5'd1, 27'h000002a0, 5'd10, 27'h000002b9, 5'd13, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000334, 5'd15, 27'h000000e8, 5'd22, 27'h0000026c, 32'h00000400,
  1'd1,  5'd3, 27'h00000063, 5'd21, 27'h000002df, 5'd1, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023a, 5'd21, 27'h00000132, 5'd13, 27'h00000016, 32'h00000400,
  1'd1,  5'd1, 27'h000003c3, 5'd25, 27'h000002f7, 5'd22, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003dd, 5'd2, 27'h000000e2, 5'd0, 27'h00000136, 32'h00000400,
  1'd1,  5'd14, 27'h000002d8, 5'd2, 27'h000000fa, 5'd15, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000301, 5'd3, 27'h000002fd, 5'd21, 27'h000003cf, 32'h00000400,
  1'd1,  5'd12, 27'h000002fa, 5'd12, 27'h00000380, 5'd4, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000355, 5'd14, 27'h000000b9, 5'd12, 27'h0000016f, 32'h00000400,
  1'd1,  5'd12, 27'h000001c5, 5'd12, 27'h0000036c, 5'd23, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d1, 5'd21, 27'h00000369, 5'd0, 27'h000002e8, 32'h00000400,
  1'd1,  5'd10, 27'h000001df, 5'd24, 27'h00000121, 5'd14, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d8, 5'd24, 27'h0000012d, 5'd20, 27'h000002fa, 32'h00000400,
  1'd1,  5'd24, 27'h00000200, 5'd1, 27'h000001a4, 5'd3, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000047, 5'd1, 27'h00000118, 5'd15, 27'h0000006c, 32'h00000400,
  1'd1,  5'd21, 27'h00000216, 5'd3, 27'h000000eb, 5'd21, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d2, 5'd13, 27'h000003f9, 5'd3, 27'h00000075, 32'h00000400,
  1'd1,  5'd23, 27'h000002b1, 5'd15, 27'h00000145, 5'd13, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000039c, 5'd10, 27'h0000018f, 5'd24, 27'h00000053, 32'h00000400,
  1'd1,  5'd22, 27'h00000106, 5'd25, 27'h00000238, 5'd0, 27'h00000242, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003b1, 5'd20, 27'h000003dc, 5'd14, 27'h000000b9, 32'h00000400,
  1'd1,  5'd23, 27'h00000138, 5'd23, 27'h0000019d, 5'd25, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ea, 5'd1, 27'h00000009, 5'd5, 27'h000001c8, 32'h00000400,
  1'd1,  5'd3, 27'h00000136, 5'd1, 27'h000003b3, 5'd17, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d4, 5'd1, 27'h0000018b, 5'd27, 27'h00000334, 32'h00000400,
  1'd1,  5'd0, 27'h0000009c, 5'd13, 27'h000003cc, 5'd8, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000297, 5'd10, 27'h000003ab, 5'd17, 27'h000001b4, 32'h00000400,
  1'd1,  5'd1, 27'h000003e7, 5'd11, 27'h00000062, 5'd29, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000102, 5'd25, 27'h0000016f, 5'd9, 27'h0000020b, 32'h00000400,
  1'd1,  5'd3, 27'h000003b5, 5'd21, 27'h00000084, 5'd20, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000009e, 5'd21, 27'h000001fd, 5'd26, 27'h0000018d, 32'h00000400,
  1'd1,  5'd12, 27'h000001e4, 5'd3, 27'h0000025d, 5'd5, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b0, 5'd4, 27'h000000ef, 5'd17, 27'h000001b8, 32'h00000400,
  1'd1,  5'd14, 27'h000002cf, 5'd5, 27'h0000009e, 5'd26, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e7, 5'd13, 27'h000002cf, 5'd9, 27'h00000243, 32'h00000400,
  1'd1,  5'd10, 27'h00000158, 5'd14, 27'h00000337, 5'd19, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000032b, 5'd11, 27'h0000020f, 5'd27, 27'h000000d4, 32'h00000400,
  1'd1,  5'd14, 27'h0000032c, 5'd23, 27'h000002db, 5'd8, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000008e, 5'd24, 27'h000002ae, 5'd20, 27'h0000025e, 32'h00000400,
  1'd1,  5'd12, 27'h000001ae, 5'd21, 27'h00000351, 5'd30, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000321, 5'd1, 27'h0000032a, 5'd7, 27'h000000cb, 32'h00000400,
  1'd1,  5'd24, 27'h00000113, 5'd0, 27'h00000098, 5'd15, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000d0, 5'd1, 27'h0000023d, 5'd26, 27'h000002db, 32'h00000400,
  1'd1,  5'd21, 27'h00000024, 5'd12, 27'h000000ed, 5'd8, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003df, 5'd12, 27'h000001e1, 5'd16, 27'h000002b0, 32'h00000400,
  1'd1,  5'd25, 27'h000000f9, 5'd14, 27'h000003e1, 5'd27, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ed, 5'd21, 27'h00000035, 5'd8, 27'h000001cc, 32'h00000400,
  1'd1,  5'd22, 27'h00000123, 5'd22, 27'h0000015b, 5'd15, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d9, 5'd24, 27'h00000376, 5'd27, 27'h00000392, 32'h00000400,
  1'd1,  5'd0, 27'h000001d7, 5'd5, 27'h0000018f, 5'd3, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012e, 5'd9, 27'h00000075, 5'd14, 27'h00000024, 32'h00000400,
  1'd1,  5'd0, 27'h00000209, 5'd9, 27'h00000263, 5'd24, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000231, 5'd20, 27'h00000238, 5'd0, 27'h00000114, 32'h00000400,
  1'd1,  5'd1, 27'h000003d9, 5'd18, 27'h00000272, 5'd15, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000015d, 5'd17, 27'h00000003, 5'd23, 27'h000002fa, 32'h00000400,
  1'd1,  5'd3, 27'h00000315, 5'd29, 27'h00000115, 5'd2, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ba, 5'd30, 27'h00000047, 5'd14, 27'h000000ab, 32'h00000400,
  1'd1,  5'd0, 27'h000002d3, 5'd27, 27'h000001d5, 5'd24, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003d0, 5'd7, 27'h000001e5, 5'd3, 27'h0000038c, 32'h00000400,
  1'd1,  5'd14, 27'h0000037c, 5'd8, 27'h000000c5, 5'd10, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000235, 5'd5, 27'h000003bb, 5'd24, 27'h00000245, 32'h00000400,
  1'd1,  5'd13, 27'h00000047, 5'd17, 27'h00000197, 5'd4, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002aa, 5'd19, 27'h0000021d, 5'd11, 27'h0000007b, 32'h00000400,
  1'd1,  5'd12, 27'h000000c3, 5'd18, 27'h0000038a, 5'd21, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000182, 5'd29, 27'h00000334, 5'd4, 27'h000003ff, 32'h00000400,
  1'd1,  5'd14, 27'h000003c1, 5'd26, 27'h00000306, 5'd15, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000191, 5'd26, 27'h000000d5, 5'd23, 27'h000003f8, 32'h00000400,
  1'd1,  5'd23, 27'h000000e3, 5'd7, 27'h0000013a, 5'd0, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000367, 5'd8, 27'h000000a2, 5'd13, 27'h0000034c, 32'h00000400,
  1'd1,  5'd24, 27'h00000392, 5'd8, 27'h000002ec, 5'd25, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000311, 5'd17, 27'h0000037f, 5'd1, 27'h000003a1, 32'h00000400,
  1'd1,  5'd25, 27'h0000015c, 5'd19, 27'h000003e1, 5'd13, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000025, 5'd19, 27'h00000025, 5'd21, 27'h000002bd, 32'h00000400,
  1'd1,  5'd23, 27'h00000051, 5'd28, 27'h00000301, 5'd0, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e4, 5'd30, 27'h000001fc, 5'd13, 27'h00000380, 32'h00000400,
  1'd1,  5'd23, 27'h00000214, 5'd29, 27'h000002de, 5'd25, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000034a, 5'd7, 27'h000001ae, 5'd5, 27'h00000107, 32'h00000400,
  1'd1,  5'd0, 27'h0000029f, 5'd5, 27'h00000267, 5'd15, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000012, 5'd7, 27'h000000bf, 5'd26, 27'h00000064, 32'h00000400,
  1'd1,  5'd1, 27'h00000257, 5'd16, 27'h0000001a, 5'd6, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ea, 5'd18, 27'h0000007a, 5'd20, 27'h00000022, 32'h00000400,
  1'd1,  5'd4, 27'h000003c4, 5'd16, 27'h0000034c, 5'd26, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000039e, 5'd26, 27'h000000e3, 5'd7, 27'h00000363, 32'h00000400,
  1'd1,  5'd1, 27'h00000325, 5'd25, 27'h000003d4, 5'd16, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000149, 5'd29, 27'h000000d9, 5'd27, 27'h0000000f, 32'h00000400,
  1'd1,  5'd13, 27'h0000022e, 5'd6, 27'h00000382, 5'd5, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000096, 5'd5, 27'h000000c7, 5'd20, 27'h00000280, 32'h00000400,
  1'd1,  5'd15, 27'h000001ad, 5'd8, 27'h000002ce, 5'd27, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000093, 5'd15, 27'h00000311, 5'd6, 27'h0000003f, 32'h00000400,
  1'd1,  5'd10, 27'h00000357, 5'd18, 27'h0000013e, 5'd17, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000001d, 5'd18, 27'h000002f9, 5'd29, 27'h000002d2, 32'h00000400,
  1'd1,  5'd13, 27'h0000027d, 5'd27, 27'h00000111, 5'd9, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000102, 5'd28, 27'h0000031b, 5'd15, 27'h0000027c, 32'h00000400,
  1'd1,  5'd13, 27'h0000003c, 5'd26, 27'h000003f6, 5'd29, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000033f, 5'd8, 27'h000001eb, 5'd6, 27'h000002a9, 32'h00000400,
  1'd1,  5'd20, 27'h000003d3, 5'd7, 27'h000003b5, 5'd20, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000295, 5'd6, 27'h000002cf, 5'd26, 27'h000000ed, 32'h00000400,
  1'd1,  5'd21, 27'h000001e2, 5'd18, 27'h000002c4, 5'd7, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000000d, 5'd18, 27'h000002e6, 5'd19, 27'h00000230, 32'h00000400,
  1'd1,  5'd24, 27'h000000d1, 5'd17, 27'h0000036b, 5'd26, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000044, 5'd27, 27'h000002df, 5'd5, 27'h000003e3, 32'h00000400,
  1'd1,  5'd25, 27'h000002c6, 5'd28, 27'h0000004d, 5'd18, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000103, 5'd30, 27'h00000022, 5'd25, 27'h0000039c, 32'h00000400,
  1'd1,  5'd6, 27'h00000086, 5'd0, 27'h0000026b, 5'd5, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000171, 5'd0, 27'h000000ae, 5'd18, 27'h000000a8, 32'h00000400,
  1'd1,  5'd5, 27'h00000355, 5'd5, 27'h00000050, 5'd25, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000190, 5'd10, 27'h00000278, 5'd1, 27'h00000177, 32'h00000400,
  1'd1,  5'd5, 27'h00000229, 5'd15, 27'h00000168, 5'd14, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021c, 5'd10, 27'h000002da, 5'd25, 27'h00000162, 32'h00000400,
  1'd1,  5'd7, 27'h000002cd, 5'd24, 27'h0000022f, 5'd3, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000008e, 5'd25, 27'h0000032d, 5'd14, 27'h0000016b, 32'h00000400,
  1'd1,  5'd9, 27'h00000153, 5'd20, 27'h000002c3, 5'd25, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000312, 5'd1, 27'h000001b4, 5'd6, 27'h00000189, 32'h00000400,
  1'd1,  5'd17, 27'h0000025f, 5'd2, 27'h0000001c, 5'd18, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000228, 5'd0, 27'h00000372, 5'd26, 27'h000002f0, 32'h00000400,
  1'd1,  5'd17, 27'h000000cb, 5'd13, 27'h000002fa, 5'd0, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002cb, 5'd14, 27'h00000167, 5'd15, 27'h000000c0, 32'h00000400,
  1'd1,  5'd17, 27'h000003a7, 5'd12, 27'h00000012, 5'd24, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000022b, 5'd24, 27'h00000202, 5'd4, 27'h000002ac, 32'h00000400,
  1'd1,  5'd15, 27'h000002bd, 5'd21, 27'h000002cf, 5'd15, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000245, 5'd22, 27'h00000023, 5'd23, 27'h0000029c, 32'h00000400,
  1'd1,  5'd30, 27'h000003e5, 5'd3, 27'h000003c4, 5'd0, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b6, 5'd4, 27'h000002b6, 5'd15, 27'h000000f7, 32'h00000400,
  1'd1,  5'd29, 27'h00000315, 5'd3, 27'h000003de, 5'd23, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000098, 5'd13, 27'h0000039c, 5'd1, 27'h00000115, 32'h00000400,
  1'd1,  5'd28, 27'h00000114, 5'd13, 27'h000000db, 5'd11, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c9, 5'd13, 27'h000000dd, 5'd25, 27'h000000ad, 32'h00000400,
  1'd1,  5'd27, 27'h00000366, 5'd21, 27'h00000078, 5'd0, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000026, 5'd24, 27'h000003af, 5'd13, 27'h00000087, 32'h00000400,
  1'd1,  5'd27, 27'h000001a7, 5'd22, 27'h00000319, 5'd22, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b5, 5'd4, 27'h00000207, 5'd3, 27'h00000115, 32'h00000400,
  1'd1,  5'd10, 27'h00000017, 5'd4, 27'h00000365, 5'd14, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000313, 5'd0, 27'h0000024f, 5'd24, 27'h000003ba, 32'h00000400,
  1'd1,  5'd8, 27'h000002ca, 5'd13, 27'h0000018c, 5'd6, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000051, 5'd13, 27'h000003a0, 5'd20, 27'h00000036, 32'h00000400,
  1'd1,  5'd9, 27'h00000183, 5'd10, 27'h00000166, 5'd28, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ad, 5'd20, 27'h000003fc, 5'd8, 27'h0000025f, 32'h00000400,
  1'd1,  5'd9, 27'h00000061, 5'd23, 27'h000001fc, 5'd15, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000136, 5'd25, 27'h0000030a, 5'd29, 27'h00000064, 32'h00000400,
  1'd1,  5'd19, 27'h000000a0, 5'd4, 27'h0000025b, 5'd0, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ff, 5'd2, 27'h00000082, 5'd12, 27'h0000002f, 32'h00000400,
  1'd1,  5'd20, 27'h00000294, 5'd5, 27'h00000012, 5'd24, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002a8, 5'd15, 27'h00000145, 5'd9, 27'h000003e9, 32'h00000400,
  1'd1,  5'd19, 27'h00000148, 5'd11, 27'h00000098, 5'd18, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e4, 5'd12, 27'h000000d8, 5'd27, 27'h000003ac, 32'h00000400,
  1'd1,  5'd18, 27'h00000029, 5'd22, 27'h0000013c, 5'd8, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016b, 5'd24, 27'h000002bf, 5'd19, 27'h000001ee, 32'h00000400,
  1'd1,  5'd18, 27'h00000020, 5'd24, 27'h000002ad, 5'd28, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038e, 5'd0, 27'h000000b9, 5'd9, 27'h0000012e, 32'h00000400,
  1'd1,  5'd27, 27'h000002e7, 5'd0, 27'h00000152, 5'd18, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000233, 5'd0, 27'h0000036e, 5'd30, 27'h000003d3, 32'h00000400,
  1'd1,  5'd28, 27'h000003bd, 5'd14, 27'h000003ac, 5'd6, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002c6, 5'd10, 27'h00000234, 5'd16, 27'h000001cd, 32'h00000400,
  1'd1,  5'd27, 27'h000001d5, 5'd12, 27'h0000021b, 5'd29, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000013e, 5'd21, 27'h00000220, 5'd8, 27'h00000177, 32'h00000400,
  1'd1,  5'd30, 27'h0000025f, 5'd21, 27'h0000001d, 5'd19, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000106, 5'd22, 27'h000000ec, 5'd26, 27'h00000370, 32'h00000400,
  1'd1,  5'd9, 27'h00000262, 5'd7, 27'h00000015, 5'd1, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000225, 5'd5, 27'h0000025a, 5'd15, 27'h00000055, 32'h00000400,
  1'd1,  5'd6, 27'h000002f3, 5'd5, 27'h0000012b, 5'd22, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000025a, 5'd16, 27'h0000016a, 5'd4, 27'h00000389, 32'h00000400,
  1'd1,  5'd7, 27'h0000000b, 5'd19, 27'h0000026b, 5'd12, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000039b, 5'd17, 27'h000003cf, 5'd23, 27'h00000384, 32'h00000400,
  1'd1,  5'd8, 27'h0000020f, 5'd27, 27'h00000273, 5'd1, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000009c, 5'd29, 27'h000002de, 5'd12, 27'h0000036a, 32'h00000400,
  1'd1,  5'd7, 27'h000001e8, 5'd27, 27'h00000088, 5'd21, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001e4, 5'd10, 27'h00000012, 5'd1, 27'h00000001, 32'h00000400,
  1'd1,  5'd20, 27'h000001e9, 5'd7, 27'h000002bb, 5'd13, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000205, 5'd9, 27'h000000c8, 5'd24, 27'h000002c4, 32'h00000400,
  1'd1,  5'd17, 27'h00000192, 5'd18, 27'h00000218, 5'd3, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ee, 5'd19, 27'h000001ac, 5'd12, 27'h00000203, 32'h00000400,
  1'd1,  5'd16, 27'h000003ab, 5'd16, 27'h000002f9, 5'd21, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000018e, 5'd29, 27'h00000016, 5'd3, 27'h0000030c, 32'h00000400,
  1'd1,  5'd17, 27'h000002da, 5'd29, 27'h00000287, 5'd14, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a8, 5'd28, 27'h000001f5, 5'd20, 27'h0000036b, 32'h00000400,
  1'd1,  5'd26, 27'h000000d0, 5'd8, 27'h0000030e, 5'd0, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003c4, 5'd8, 27'h000003fc, 5'd15, 27'h000001b5, 32'h00000400,
  1'd1,  5'd28, 27'h00000216, 5'd8, 27'h000003b2, 5'd21, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002bd, 5'd17, 27'h00000254, 5'd3, 27'h00000316, 32'h00000400,
  1'd1,  5'd26, 27'h0000039d, 5'd19, 27'h000001f2, 5'd15, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000016f, 5'd19, 27'h000000e4, 5'd25, 27'h00000311, 32'h00000400,
  1'd1,  5'd29, 27'h0000019a, 5'd28, 27'h0000014c, 5'd3, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007b, 5'd26, 27'h000003c5, 5'd12, 27'h0000026b, 32'h00000400,
  1'd1,  5'd29, 27'h00000169, 5'd25, 27'h0000037e, 5'd25, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000000b, 5'd9, 27'h00000333, 5'd9, 27'h00000098, 32'h00000400,
  1'd1,  5'd6, 27'h0000014f, 5'd9, 27'h000002c0, 5'd18, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000290, 5'd10, 27'h00000038, 5'd30, 27'h000001fe, 32'h00000400,
  1'd1,  5'd6, 27'h000002c5, 5'd17, 27'h000001a3, 5'd9, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b8, 5'd20, 27'h00000126, 5'd16, 27'h0000020f, 32'h00000400,
  1'd1,  5'd10, 27'h00000079, 5'd16, 27'h00000387, 5'd30, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000188, 5'd29, 27'h000000de, 5'd5, 27'h000000f0, 32'h00000400,
  1'd1,  5'd5, 27'h00000129, 5'd30, 27'h0000001a, 5'd20, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e9, 5'd28, 27'h000002a3, 5'd28, 27'h00000140, 32'h00000400,
  1'd1,  5'd16, 27'h0000038b, 5'd9, 27'h000002e8, 5'd5, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000286, 5'd8, 27'h00000155, 5'd20, 27'h00000295, 32'h00000400,
  1'd1,  5'd20, 27'h00000053, 5'd7, 27'h00000171, 5'd30, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001f4, 5'd15, 27'h00000293, 5'd5, 27'h00000187, 32'h00000400,
  1'd1,  5'd19, 27'h0000004c, 5'd15, 27'h000003d7, 5'd16, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000006f, 5'd15, 27'h0000022d, 5'd26, 27'h000000e0, 32'h00000400,
  1'd1,  5'd17, 27'h00000117, 5'd26, 27'h00000296, 5'd7, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000057, 5'd28, 27'h000000fa, 5'd19, 27'h000002de, 32'h00000400,
  1'd1,  5'd18, 27'h0000023c, 5'd29, 27'h000001af, 5'd28, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003be, 5'd5, 27'h00000274, 5'd7, 27'h00000263, 32'h00000400,
  1'd1,  5'd28, 27'h00000138, 5'd10, 27'h00000086, 5'd17, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000008a, 5'd7, 27'h000002fd, 5'd27, 27'h0000001f, 32'h00000400,
  1'd1,  5'd29, 27'h000000e5, 5'd20, 27'h000000d4, 5'd6, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e5, 5'd18, 27'h000003d3, 5'd16, 27'h00000337, 32'h00000400,
  1'd1,  5'd30, 27'h0000007d, 5'd16, 27'h0000019c, 5'd28, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e1, 5'd27, 27'h00000314, 5'd9, 27'h000000d2, 32'h00000400,
  1'd1,  5'd30, 27'h00000090, 5'd26, 27'h00000383, 5'd19, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000202, 5'd30, 27'h00000374, 5'd29, 27'h00000030, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000022f, 5'd0, 27'h000000ac, 5'd0, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c6, 5'd3, 27'h000000a9, 5'd15, 27'h000000c8, 32'h00000400,
  1'd1,  5'd2, 27'h0000034f, 5'd1, 27'h0000003c, 5'd21, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000195, 5'd11, 27'h000000bc, 5'd4, 27'h00000278, 32'h00000400,
  1'd1,  5'd0, 27'h00000121, 5'd13, 27'h0000025c, 5'd11, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000039, 5'd15, 27'h00000036, 5'd22, 27'h00000267, 32'h00000400,
  1'd1,  5'd2, 27'h00000376, 5'd23, 27'h0000001e, 5'd3, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c1, 5'd23, 27'h000002a0, 5'd11, 27'h0000039c, 32'h00000400,
  1'd1,  5'd0, 27'h000000a5, 5'd21, 27'h00000329, 5'd25, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000033, 5'd2, 27'h0000027f, 5'd0, 27'h000000c5, 32'h00000400,
  1'd1,  5'd12, 27'h000001ee, 5'd1, 27'h0000027c, 5'd13, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035d, 5'd2, 27'h0000009f, 5'd25, 27'h000002ce, 32'h00000400,
  1'd1,  5'd12, 27'h0000027b, 5'd14, 27'h00000238, 5'd4, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002a6, 5'd15, 27'h000001ab, 5'd13, 27'h00000129, 32'h00000400,
  1'd1,  5'd12, 27'h00000323, 5'd13, 27'h00000185, 5'd25, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000037a, 5'd20, 27'h0000037c, 5'd4, 27'h00000098, 32'h00000400,
  1'd1,  5'd12, 27'h0000024b, 5'd20, 27'h00000358, 5'd14, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b1, 5'd20, 27'h00000360, 5'd21, 27'h00000268, 32'h00000400,
  1'd1,  5'd21, 27'h00000085, 5'd0, 27'h000002ac, 5'd3, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000002f, 5'd3, 27'h00000062, 5'd11, 27'h0000038c, 32'h00000400,
  1'd1,  5'd24, 27'h00000033, 5'd4, 27'h00000094, 5'd22, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000181, 5'd10, 27'h00000347, 5'd4, 27'h00000056, 32'h00000400,
  1'd1,  5'd23, 27'h00000393, 5'd11, 27'h00000039, 5'd10, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000333, 5'd14, 27'h00000122, 5'd22, 27'h00000105, 32'h00000400,
  1'd1,  5'd25, 27'h00000055, 5'd22, 27'h00000389, 5'd3, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002d4, 5'd25, 27'h00000058, 5'd10, 27'h0000034c, 32'h00000400,
  1'd1,  5'd23, 27'h00000087, 5'd22, 27'h00000255, 5'd21, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001a7, 5'd2, 27'h000001df, 5'd8, 27'h00000028, 32'h00000400,
  1'd1,  5'd2, 27'h00000001, 5'd1, 27'h00000312, 5'd20, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000214, 5'd1, 27'h00000239, 5'd26, 27'h00000305, 32'h00000400,
  1'd1,  5'd3, 27'h00000070, 5'd12, 27'h00000389, 5'd6, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000070, 5'd13, 27'h00000056, 5'd15, 27'h0000036b, 32'h00000400,
  1'd1,  5'd1, 27'h0000015c, 5'd14, 27'h0000008d, 5'd26, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000025b, 5'd20, 27'h000003b6, 5'd6, 27'h000003aa, 32'h00000400,
  1'd1,  5'd2, 27'h0000039b, 5'd24, 27'h00000195, 5'd16, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039c, 5'd21, 27'h0000003a, 5'd30, 27'h0000019b, 32'h00000400,
  1'd1,  5'd13, 27'h000003d7, 5'd2, 27'h00000366, 5'd6, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e0, 5'd4, 27'h000002de, 5'd20, 27'h000000d3, 32'h00000400,
  1'd1,  5'd15, 27'h00000015, 5'd1, 27'h0000023f, 5'd27, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001cd, 5'd14, 27'h0000034a, 5'd6, 27'h000002c6, 32'h00000400,
  1'd1,  5'd15, 27'h00000074, 5'd14, 27'h00000343, 5'd20, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000217, 5'd14, 27'h000001b5, 5'd26, 27'h000001c9, 32'h00000400,
  1'd1,  5'd11, 27'h000001fe, 5'd21, 27'h0000010e, 5'd9, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000342, 5'd22, 27'h000000fb, 5'd16, 27'h00000249, 32'h00000400,
  1'd1,  5'd14, 27'h0000006e, 5'd21, 27'h00000081, 5'd28, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ec, 5'd4, 27'h000003bc, 5'd7, 27'h00000138, 32'h00000400,
  1'd1,  5'd22, 27'h0000028b, 5'd4, 27'h00000272, 5'd20, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003a1, 5'd2, 27'h000003cb, 5'd29, 27'h000001f8, 32'h00000400,
  1'd1,  5'd25, 27'h000000ca, 5'd13, 27'h0000028d, 5'd7, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ed, 5'd13, 27'h000003a1, 5'd18, 27'h000001fa, 32'h00000400,
  1'd1,  5'd24, 27'h000003a9, 5'd11, 27'h000002a5, 5'd30, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000016, 5'd24, 27'h000000c4, 5'd8, 27'h00000143, 32'h00000400,
  1'd1,  5'd21, 27'h000003b8, 5'd21, 27'h000002c8, 5'd17, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000032b, 5'd20, 27'h000002b8, 5'd28, 27'h00000100, 32'h00000400,
  1'd1,  5'd4, 27'h0000011a, 5'd6, 27'h000003e6, 5'd2, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a3, 5'd8, 27'h00000010, 5'd14, 27'h000003f5, 32'h00000400,
  1'd1,  5'd2, 27'h00000030, 5'd7, 27'h00000046, 5'd23, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000fe, 5'd16, 27'h000002db, 5'd2, 27'h000003ab, 32'h00000400,
  1'd1,  5'd5, 27'h0000006c, 5'd20, 27'h00000002, 5'd11, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000385, 5'd15, 27'h00000348, 5'd21, 27'h00000113, 32'h00000400,
  1'd1,  5'd0, 27'h00000024, 5'd27, 27'h0000035d, 5'd1, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000f2, 5'd29, 27'h000003d0, 5'd15, 27'h000000f7, 32'h00000400,
  1'd1,  5'd0, 27'h000002dd, 5'd27, 27'h00000249, 5'd23, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000397, 5'd9, 27'h0000024d, 5'd4, 27'h00000064, 32'h00000400,
  1'd1,  5'd10, 27'h000002a2, 5'd8, 27'h0000000f, 5'd14, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f6, 5'd8, 27'h0000036e, 5'd23, 27'h000003a0, 32'h00000400,
  1'd1,  5'd10, 27'h0000023e, 5'd18, 27'h000001bb, 5'd2, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000037d, 5'd19, 27'h00000336, 5'd15, 27'h0000014a, 32'h00000400,
  1'd1,  5'd13, 27'h00000379, 5'd15, 27'h00000384, 5'd24, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003fb, 5'd29, 27'h0000030e, 5'd3, 27'h000001dc, 32'h00000400,
  1'd1,  5'd12, 27'h000000d8, 5'd26, 27'h0000000e, 5'd13, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003f9, 5'd28, 27'h000001af, 5'd23, 27'h00000155, 32'h00000400,
  1'd1,  5'd21, 27'h00000369, 5'd6, 27'h00000125, 5'd3, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000008, 5'd7, 27'h00000199, 5'd13, 27'h000000bb, 32'h00000400,
  1'd1,  5'd20, 27'h00000325, 5'd9, 27'h0000031f, 5'd22, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c4, 5'd19, 27'h00000015, 5'd0, 27'h000003a9, 32'h00000400,
  1'd1,  5'd23, 27'h000001b4, 5'd19, 27'h0000037c, 5'd14, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000f9, 5'd17, 27'h00000396, 5'd25, 27'h0000025f, 32'h00000400,
  1'd1,  5'd25, 27'h000000e8, 5'd28, 27'h000003cf, 5'd4, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000160, 5'd28, 27'h00000081, 5'd14, 27'h000001d4, 32'h00000400,
  1'd1,  5'd25, 27'h00000244, 5'd30, 27'h000003e6, 5'd22, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ce, 5'd10, 27'h000000c6, 5'd7, 27'h000002d4, 32'h00000400,
  1'd1,  5'd1, 27'h000001da, 5'd9, 27'h000000a1, 5'd19, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000347, 5'd6, 27'h00000181, 5'd28, 27'h0000025b, 32'h00000400,
  1'd1,  5'd2, 27'h0000028a, 5'd20, 27'h000001fa, 5'd5, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000116, 5'd17, 27'h0000008d, 5'd16, 27'h00000344, 32'h00000400,
  1'd1,  5'd1, 27'h00000307, 5'd17, 27'h00000001, 5'd27, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000024e, 5'd26, 27'h00000099, 5'd8, 27'h0000027c, 32'h00000400,
  1'd1,  5'd0, 27'h00000369, 5'd27, 27'h000003a4, 5'd18, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002a9, 5'd28, 27'h00000381, 5'd27, 27'h00000197, 32'h00000400,
  1'd1,  5'd11, 27'h00000189, 5'd9, 27'h00000140, 5'd6, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000038d, 5'd5, 27'h000001ae, 5'd16, 27'h000000cd, 32'h00000400,
  1'd1,  5'd12, 27'h0000010d, 5'd7, 27'h000003a5, 5'd27, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000384, 5'd20, 27'h0000010c, 5'd6, 27'h00000267, 32'h00000400,
  1'd1,  5'd13, 27'h000003e8, 5'd15, 27'h000003e1, 5'd15, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000013e, 5'd19, 27'h00000180, 5'd27, 27'h00000105, 32'h00000400,
  1'd1,  5'd14, 27'h00000123, 5'd27, 27'h0000018d, 5'd10, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a2, 5'd27, 27'h0000025a, 5'd18, 27'h000001d4, 32'h00000400,
  1'd1,  5'd10, 27'h000003ad, 5'd28, 27'h00000224, 5'd30, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e4, 5'd8, 27'h0000033d, 5'd6, 27'h00000174, 32'h00000400,
  1'd1,  5'd22, 27'h00000131, 5'd10, 27'h000000f4, 5'd19, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d4, 5'd6, 27'h00000315, 5'd30, 27'h00000220, 32'h00000400,
  1'd1,  5'd21, 27'h000001f9, 5'd19, 27'h00000302, 5'd7, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b2, 5'd18, 27'h000001ff, 5'd15, 27'h00000372, 32'h00000400,
  1'd1,  5'd24, 27'h0000024b, 5'd19, 27'h000003b1, 5'd28, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000237, 5'd26, 27'h00000052, 5'd8, 27'h000000b2, 32'h00000400,
  1'd1,  5'd23, 27'h00000264, 5'd28, 27'h000001cf, 5'd16, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000033b, 5'd27, 27'h0000033e, 5'd28, 27'h0000025d, 32'h00000400,
  1'd1,  5'd8, 27'h00000010, 5'd4, 27'h0000027b, 5'd5, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000092, 5'd2, 27'h000002b6, 5'd19, 27'h00000336, 32'h00000400,
  1'd1,  5'd6, 27'h0000011a, 5'd0, 27'h0000038f, 5'd29, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000f3, 5'd11, 27'h000001ab, 5'd4, 27'h000001e7, 32'h00000400,
  1'd1,  5'd9, 27'h000003a9, 5'd14, 27'h0000014e, 5'd10, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002cb, 5'd14, 27'h00000025, 5'd22, 27'h00000060, 32'h00000400,
  1'd1,  5'd8, 27'h00000203, 5'd25, 27'h00000076, 5'd1, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000022c, 5'd25, 27'h0000002b, 5'd12, 27'h00000044, 32'h00000400,
  1'd1,  5'd9, 27'h000001e5, 5'd22, 27'h000000ee, 5'd24, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c8, 5'd0, 27'h00000349, 5'd10, 27'h00000014, 32'h00000400,
  1'd1,  5'd19, 27'h0000010f, 5'd4, 27'h000001ce, 5'd20, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000082, 5'd2, 27'h000002cf, 5'd28, 27'h00000138, 32'h00000400,
  1'd1,  5'd16, 27'h0000018d, 5'd10, 27'h0000027a, 5'd1, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000294, 5'd13, 27'h000000c0, 5'd12, 27'h00000172, 32'h00000400,
  1'd1,  5'd20, 27'h000000cd, 5'd11, 27'h000001bf, 5'd24, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000211, 5'd22, 27'h0000037d, 5'd3, 27'h00000241, 32'h00000400,
  1'd1,  5'd17, 27'h00000020, 5'd22, 27'h000000d2, 5'd14, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000080, 5'd21, 27'h000003bc, 5'd21, 27'h0000032c, 32'h00000400,
  1'd1,  5'd28, 27'h000001e3, 5'd3, 27'h000003fa, 5'd0, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000043, 5'd2, 27'h00000317, 5'd15, 27'h00000141, 32'h00000400,
  1'd1,  5'd30, 27'h00000174, 5'd4, 27'h00000033, 5'd23, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003df, 5'd15, 27'h0000002f, 5'd3, 27'h00000100, 32'h00000400,
  1'd1,  5'd28, 27'h00000247, 5'd15, 27'h000000bd, 5'd12, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000245, 5'd11, 27'h000003e0, 5'd22, 27'h000003ce, 32'h00000400,
  1'd1,  5'd30, 27'h000002fb, 5'd25, 27'h000002ed, 5'd0, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003dc, 5'd21, 27'h000000b2, 5'd11, 27'h0000012a, 32'h00000400,
  1'd1,  5'd29, 27'h00000163, 5'd21, 27'h00000109, 5'd23, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000389, 5'd1, 27'h000001f5, 5'd3, 27'h000003df, 32'h00000400,
  1'd1,  5'd5, 27'h000003e5, 5'd2, 27'h0000016e, 5'd11, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000008, 5'd3, 27'h00000320, 5'd22, 27'h00000298, 32'h00000400,
  1'd1,  5'd5, 27'h000002db, 5'd11, 27'h0000001a, 5'd7, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001b3, 5'd11, 27'h0000032c, 5'd20, 27'h00000136, 32'h00000400,
  1'd1,  5'd7, 27'h00000015, 5'd10, 27'h000002ac, 5'd28, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000076, 5'd22, 27'h0000027b, 5'd9, 27'h00000271, 32'h00000400,
  1'd1,  5'd8, 27'h000001e7, 5'd23, 27'h0000039d, 5'd18, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000011c, 5'd24, 27'h0000005d, 5'd26, 27'h00000321, 32'h00000400,
  1'd1,  5'd17, 27'h00000141, 5'd1, 27'h000003a6, 5'd5, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000b3, 5'd4, 27'h00000343, 5'd14, 27'h00000264, 32'h00000400,
  1'd1,  5'd18, 27'h000000b3, 5'd2, 27'h000003ee, 5'd22, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000079, 5'd11, 27'h000002bb, 5'd5, 27'h00000114, 32'h00000400,
  1'd1,  5'd17, 27'h0000022a, 5'd14, 27'h000003ad, 5'd18, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000234, 5'd10, 27'h00000269, 5'd30, 27'h0000029c, 32'h00000400,
  1'd1,  5'd19, 27'h0000000f, 5'd22, 27'h000000c0, 5'd7, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000002c, 5'd25, 27'h000002fb, 5'd16, 27'h00000111, 32'h00000400,
  1'd1,  5'd17, 27'h00000362, 5'd22, 27'h000002b0, 5'd26, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000157, 5'd0, 27'h00000031, 5'd7, 27'h000003b0, 32'h00000400,
  1'd1,  5'd27, 27'h000003da, 5'd4, 27'h000000d0, 5'd20, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000316, 5'd1, 27'h000002f9, 5'd30, 27'h000003c5, 32'h00000400,
  1'd1,  5'd25, 27'h00000382, 5'd10, 27'h000001b4, 5'd9, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000026e, 5'd11, 27'h000000a7, 5'd20, 27'h00000046, 32'h00000400,
  1'd1,  5'd27, 27'h0000025c, 5'd11, 27'h00000303, 5'd29, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000323, 5'd23, 27'h0000031f, 5'd5, 27'h000000c2, 32'h00000400,
  1'd1,  5'd29, 27'h0000017d, 5'd21, 27'h00000036, 5'd20, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000203, 5'd21, 27'h0000033c, 5'd26, 27'h00000291, 32'h00000400,
  1'd1,  5'd8, 27'h00000275, 5'd10, 27'h0000013b, 5'd4, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000211, 5'd7, 27'h00000332, 5'd14, 27'h0000011e, 32'h00000400,
  1'd1,  5'd6, 27'h00000005, 5'd8, 27'h00000151, 5'd23, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e7, 5'd20, 27'h0000011e, 5'd2, 27'h000003af, 32'h00000400,
  1'd1,  5'd9, 27'h0000020a, 5'd19, 27'h000003ae, 5'd11, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000165, 5'd15, 27'h000003a6, 5'd25, 27'h0000021b, 32'h00000400,
  1'd1,  5'd9, 27'h00000120, 5'd27, 27'h000002b5, 5'd2, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000307, 5'd29, 27'h000003c7, 5'd12, 27'h00000244, 32'h00000400,
  1'd1,  5'd8, 27'h00000371, 5'd26, 27'h000003c5, 5'd25, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000296, 5'd8, 27'h00000117, 5'd2, 27'h00000219, 32'h00000400,
  1'd1,  5'd19, 27'h000000d2, 5'd7, 27'h00000013, 5'd12, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000002d, 5'd6, 27'h000002c8, 5'd22, 27'h00000057, 32'h00000400,
  1'd1,  5'd20, 27'h0000014b, 5'd19, 27'h00000266, 5'd2, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000190, 5'd20, 27'h0000006c, 5'd12, 27'h00000214, 32'h00000400,
  1'd1,  5'd17, 27'h0000020d, 5'd15, 27'h0000036e, 5'd20, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ac, 5'd29, 27'h00000295, 5'd2, 27'h00000376, 32'h00000400,
  1'd1,  5'd18, 27'h00000184, 5'd29, 27'h000001ea, 5'd14, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000192, 5'd30, 27'h000000b5, 5'd25, 27'h000002ef, 32'h00000400,
  1'd1,  5'd29, 27'h0000013d, 5'd6, 27'h00000020, 5'd4, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000009b, 5'd6, 27'h00000273, 5'd15, 27'h00000194, 32'h00000400,
  1'd1,  5'd27, 27'h00000256, 5'd5, 27'h00000215, 5'd22, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000019f, 5'd16, 27'h000002cb, 5'd3, 27'h00000375, 32'h00000400,
  1'd1,  5'd27, 27'h0000023e, 5'd18, 27'h0000032c, 5'd13, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000356, 5'd17, 27'h000002a2, 5'd24, 27'h00000003, 32'h00000400,
  1'd1,  5'd27, 27'h000000ff, 5'd28, 27'h0000009d, 5'd3, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003ef, 5'd28, 27'h0000009b, 5'd15, 27'h00000074, 32'h00000400,
  1'd1,  5'd28, 27'h00000241, 5'd29, 27'h000003b5, 5'd24, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000218, 5'd9, 27'h0000006a, 5'd7, 27'h000003df, 32'h00000400,
  1'd1,  5'd10, 27'h00000093, 5'd6, 27'h0000004f, 5'd19, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000014, 5'd8, 27'h0000010e, 5'd26, 27'h00000044, 32'h00000400,
  1'd1,  5'd6, 27'h00000376, 5'd15, 27'h000002c8, 5'd5, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000147, 5'd17, 27'h0000008f, 5'd16, 27'h00000074, 32'h00000400,
  1'd1,  5'd7, 27'h0000027d, 5'd15, 27'h000002e9, 5'd28, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000030d, 5'd30, 27'h000002f9, 5'd8, 27'h00000153, 32'h00000400,
  1'd1,  5'd8, 27'h00000051, 5'd28, 27'h00000263, 5'd19, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c7, 5'd29, 27'h0000017b, 5'd26, 27'h000003eb, 32'h00000400,
  1'd1,  5'd18, 27'h0000030c, 5'd9, 27'h0000036a, 5'd9, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000010, 5'd6, 27'h00000397, 5'd20, 27'h0000015c, 32'h00000400,
  1'd1,  5'd18, 27'h0000001f, 5'd8, 27'h000000a4, 5'd27, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000022b, 5'd17, 27'h000002fc, 5'd9, 27'h00000015, 32'h00000400,
  1'd1,  5'd16, 27'h00000289, 5'd17, 27'h0000006f, 5'd16, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000051, 5'd18, 27'h00000262, 5'd30, 27'h00000350, 32'h00000400,
  1'd1,  5'd19, 27'h0000010d, 5'd25, 27'h0000036c, 5'd8, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000fe, 5'd30, 27'h0000014d, 5'd20, 27'h000000f0, 32'h00000400,
  1'd1,  5'd19, 27'h000003f1, 5'd28, 27'h000001bd, 5'd27, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000006f, 5'd6, 27'h000003c6, 5'd9, 27'h00000283, 32'h00000400,
  1'd1,  5'd28, 27'h000003fc, 5'd7, 27'h0000025c, 5'd18, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000151, 5'd5, 27'h0000021e, 5'd26, 27'h000001fd, 32'h00000400,
  1'd1,  5'd28, 27'h00000065, 5'd20, 27'h00000136, 5'd9, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002af, 5'd19, 27'h000001e4, 5'd19, 27'h0000000a, 32'h00000400,
  1'd1,  5'd29, 27'h00000090, 5'd18, 27'h0000012a, 5'd28, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000025f, 5'd29, 27'h0000039e, 5'd5, 27'h000002e2, 32'h00000400,
  1'd1,  5'd29, 27'h00000355, 5'd29, 27'h000001ec, 5'd17, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000031f, 5'd29, 27'h00000376, 5'd28, 27'h0000022e, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h0000038f, 5'd4, 27'h00000116, 5'd1, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000101, 5'd3, 27'h0000019b, 5'd12, 27'h000002b5, 32'h00000400,
  1'd1,  5'd2, 27'h00000365, 5'd4, 27'h000002a2, 5'd23, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001cc, 5'd10, 27'h0000024e, 5'd4, 27'h00000186, 32'h00000400,
  1'd1,  5'd2, 27'h0000027f, 5'd14, 27'h000002e0, 5'd11, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001de, 5'd11, 27'h0000031c, 5'd22, 27'h000001c9, 32'h00000400,
  1'd1,  5'd1, 27'h000001c0, 5'd23, 27'h00000325, 5'd4, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000100, 5'd21, 27'h000001ba, 5'd10, 27'h000003f9, 32'h00000400,
  1'd1,  5'd2, 27'h000003fe, 5'd21, 27'h000003db, 5'd20, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000067, 5'd1, 27'h0000023a, 5'd0, 27'h00000309, 32'h00000400,
  1'd1,  5'd12, 27'h0000002b, 5'd0, 27'h00000328, 5'd10, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000017f, 5'd0, 27'h0000028c, 5'd20, 27'h000003ac, 32'h00000400,
  1'd1,  5'd13, 27'h000001b2, 5'd11, 27'h00000131, 5'd0, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000083, 5'd13, 27'h0000010d, 5'd13, 27'h00000327, 32'h00000400,
  1'd1,  5'd11, 27'h000003a8, 5'd12, 27'h00000206, 5'd24, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ec, 5'd23, 27'h0000006f, 5'd3, 27'h00000035, 32'h00000400,
  1'd1,  5'd12, 27'h0000033f, 5'd24, 27'h0000037b, 5'd11, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c0, 5'd21, 27'h00000303, 5'd23, 27'h0000000a, 32'h00000400,
  1'd1,  5'd25, 27'h0000012f, 5'd1, 27'h0000022c, 5'd0, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000092, 5'd2, 27'h000003c8, 5'd14, 27'h00000183, 32'h00000400,
  1'd1,  5'd24, 27'h000001b8, 5'd4, 27'h00000192, 5'd25, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000136, 5'd12, 27'h000003c7, 5'd0, 27'h00000217, 32'h00000400,
  1'd1,  5'd25, 27'h00000006, 5'd13, 27'h00000034, 5'd10, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000354, 5'd11, 27'h00000230, 5'd21, 27'h000003c3, 32'h00000400,
  1'd1,  5'd25, 27'h00000061, 5'd24, 27'h00000263, 5'd4, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000267, 5'd24, 27'h00000318, 5'd14, 27'h000002d2, 32'h00000400,
  1'd1,  5'd24, 27'h00000313, 5'd20, 27'h00000351, 5'd22, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a4, 5'd1, 27'h0000025e, 5'd7, 27'h00000181, 32'h00000400,
  1'd1,  5'd2, 27'h0000004c, 5'd4, 27'h0000018e, 5'd16, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000018f, 5'd3, 27'h00000270, 5'd27, 27'h000003e4, 32'h00000400,
  1'd1,  5'd4, 27'h0000010f, 5'd14, 27'h000001d9, 5'd9, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000016c, 5'd14, 27'h000002a9, 5'd17, 27'h0000001d, 32'h00000400,
  1'd1,  5'd3, 27'h000001bf, 5'd15, 27'h000001fd, 5'd29, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003ce, 5'd23, 27'h000002cc, 5'd5, 27'h000002b0, 32'h00000400,
  1'd1,  5'd0, 27'h0000030e, 5'd22, 27'h0000014c, 5'd19, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000022e, 5'd23, 27'h000003bc, 5'd30, 27'h0000005a, 32'h00000400,
  1'd1,  5'd12, 27'h0000001a, 5'd4, 27'h0000024e, 5'd7, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000019f, 5'd0, 27'h000002fc, 5'd19, 27'h0000015f, 32'h00000400,
  1'd1,  5'd13, 27'h00000153, 5'd0, 27'h00000138, 5'd30, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003d4, 5'd14, 27'h000003e1, 5'd8, 27'h00000062, 32'h00000400,
  1'd1,  5'd11, 27'h00000248, 5'd11, 27'h00000112, 5'd17, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d9, 5'd12, 27'h0000030c, 5'd26, 27'h00000283, 32'h00000400,
  1'd1,  5'd11, 27'h000003e2, 5'd22, 27'h00000273, 5'd7, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002bc, 5'd21, 27'h00000331, 5'd20, 27'h000000bc, 32'h00000400,
  1'd1,  5'd12, 27'h000003f4, 5'd24, 27'h00000036, 5'd28, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000027d, 5'd0, 27'h000000ea, 5'd8, 27'h0000036b, 32'h00000400,
  1'd1,  5'd23, 27'h000002a7, 5'd1, 27'h0000029b, 5'd20, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003aa, 5'd4, 27'h000001e8, 5'd28, 27'h000000d9, 32'h00000400,
  1'd1,  5'd23, 27'h00000156, 5'd14, 27'h00000342, 5'd7, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000274, 5'd15, 27'h00000128, 5'd18, 27'h000003e0, 32'h00000400,
  1'd1,  5'd25, 27'h00000328, 5'd14, 27'h0000019b, 5'd26, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001ac, 5'd23, 27'h0000031b, 5'd8, 27'h00000265, 32'h00000400,
  1'd1,  5'd25, 27'h000002d3, 5'd20, 27'h000003cc, 5'd19, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000027c, 5'd24, 27'h0000002f, 5'd27, 27'h00000338, 32'h00000400,
  1'd1,  5'd0, 27'h000003f4, 5'd7, 27'h0000017b, 5'd0, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000270, 5'd8, 27'h000000bb, 5'd11, 27'h0000034a, 32'h00000400,
  1'd1,  5'd4, 27'h000000fa, 5'd8, 27'h000002d4, 5'd21, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039d, 5'd19, 27'h000002bd, 5'd0, 27'h00000169, 32'h00000400,
  1'd1,  5'd3, 27'h0000036f, 5'd20, 27'h000001f2, 5'd11, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000270, 5'd19, 27'h000001c4, 5'd21, 27'h000001f6, 32'h00000400,
  1'd1,  5'd1, 27'h000003a7, 5'd30, 27'h00000184, 5'd2, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001d6, 5'd28, 27'h000000a3, 5'd13, 27'h000003f5, 32'h00000400,
  1'd1,  5'd3, 27'h000001b8, 5'd26, 27'h000002e4, 5'd21, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000002f, 5'd8, 27'h000001c8, 5'd3, 27'h000000d2, 32'h00000400,
  1'd1,  5'd11, 27'h0000015d, 5'd7, 27'h0000004a, 5'd10, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000033c, 5'd8, 27'h0000003e, 5'd24, 27'h00000293, 32'h00000400,
  1'd1,  5'd13, 27'h0000012d, 5'd17, 27'h0000017f, 5'd3, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002aa, 5'd16, 27'h0000035f, 5'd10, 27'h000001fd, 32'h00000400,
  1'd1,  5'd11, 27'h00000097, 5'd18, 27'h000001b4, 5'd25, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000027f, 5'd27, 27'h000003ca, 5'd0, 27'h00000258, 32'h00000400,
  1'd1,  5'd14, 27'h000003d0, 5'd27, 27'h000001dc, 5'd12, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000028c, 5'd30, 27'h000002cc, 5'd20, 27'h000003a3, 32'h00000400,
  1'd1,  5'd24, 27'h00000043, 5'd10, 27'h00000117, 5'd2, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f2, 5'd6, 27'h00000363, 5'd13, 27'h00000236, 32'h00000400,
  1'd1,  5'd25, 27'h0000023e, 5'd6, 27'h00000181, 5'd22, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000186, 5'd19, 27'h000003d4, 5'd4, 27'h000003d9, 32'h00000400,
  1'd1,  5'd22, 27'h000002dd, 5'd20, 27'h00000194, 5'd11, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000233, 5'd15, 27'h00000237, 5'd22, 27'h0000002f, 32'h00000400,
  1'd1,  5'd24, 27'h000001bb, 5'd28, 27'h00000291, 5'd3, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000012d, 5'd28, 27'h00000239, 5'd11, 27'h0000018e, 32'h00000400,
  1'd1,  5'd21, 27'h00000383, 5'd30, 27'h000000ea, 5'd21, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000fa, 5'd5, 27'h00000267, 5'd9, 27'h00000323, 32'h00000400,
  1'd1,  5'd4, 27'h000002c2, 5'd10, 27'h0000003d, 5'd20, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ce, 5'd8, 27'h00000079, 5'd25, 27'h00000389, 32'h00000400,
  1'd1,  5'd2, 27'h00000067, 5'd17, 27'h0000035f, 5'd5, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f3, 5'd19, 27'h000002b6, 5'd20, 27'h00000196, 32'h00000400,
  1'd1,  5'd4, 27'h00000326, 5'd20, 27'h00000090, 5'd30, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000022f, 5'd28, 27'h000001e0, 5'd9, 27'h00000039, 32'h00000400,
  1'd1,  5'd0, 27'h0000038e, 5'd26, 27'h000001f1, 5'd17, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000007a, 5'd26, 27'h00000221, 5'd27, 27'h000000c9, 32'h00000400,
  1'd1,  5'd14, 27'h00000317, 5'd8, 27'h000001d8, 5'd8, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000016d, 5'd8, 27'h0000010c, 5'd19, 27'h00000386, 32'h00000400,
  1'd1,  5'd15, 27'h00000061, 5'd6, 27'h000000bb, 5'd28, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000018f, 5'd17, 27'h000002dc, 5'd6, 27'h000002a2, 32'h00000400,
  1'd1,  5'd12, 27'h000002dc, 5'd19, 27'h000002ca, 5'd18, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000226, 5'd17, 27'h0000033f, 5'd30, 27'h00000047, 32'h00000400,
  1'd1,  5'd12, 27'h00000153, 5'd29, 27'h000000b5, 5'd7, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000174, 5'd28, 27'h00000095, 5'd19, 27'h000003d9, 32'h00000400,
  1'd1,  5'd13, 27'h00000240, 5'd29, 27'h000003f4, 5'd27, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000350, 5'd7, 27'h0000013f, 5'd5, 27'h0000022e, 32'h00000400,
  1'd1,  5'd25, 27'h000001a3, 5'd6, 27'h000003d6, 5'd20, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000069, 5'd8, 27'h00000046, 5'd26, 27'h00000273, 32'h00000400,
  1'd1,  5'd25, 27'h000002d9, 5'd18, 27'h0000033d, 5'd7, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003df, 5'd19, 27'h00000118, 5'd20, 27'h000000db, 32'h00000400,
  1'd1,  5'd25, 27'h00000092, 5'd18, 27'h00000294, 5'd30, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000184, 5'd25, 27'h000003b9, 5'd9, 27'h0000005d, 32'h00000400,
  1'd1,  5'd22, 27'h0000010e, 5'd28, 27'h000001ab, 5'd20, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000129, 5'd29, 27'h000002b3, 5'd29, 27'h000001ab, 32'h00000400,
  1'd1,  5'd9, 27'h0000013c, 5'd3, 27'h00000036, 5'd6, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000153, 5'd3, 27'h000001c3, 5'd18, 27'h000003ce, 32'h00000400,
  1'd1,  5'd8, 27'h000001f8, 5'd1, 27'h000003a8, 5'd29, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000034, 5'd13, 27'h00000068, 5'd4, 27'h000002ce, 32'h00000400,
  1'd1,  5'd5, 27'h0000033a, 5'd13, 27'h00000236, 5'd12, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e1, 5'd12, 27'h00000107, 5'd22, 27'h00000380, 32'h00000400,
  1'd1,  5'd7, 27'h000001f2, 5'd22, 27'h000002d0, 5'd3, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ad, 5'd24, 27'h0000017c, 5'd11, 27'h000002d1, 32'h00000400,
  1'd1,  5'd8, 27'h000000bc, 5'd24, 27'h000003cc, 5'd23, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000024b, 5'd1, 27'h00000396, 5'd7, 27'h000002ab, 32'h00000400,
  1'd1,  5'd16, 27'h000003c7, 5'd3, 27'h000001f7, 5'd18, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c2, 5'd1, 27'h000001ff, 5'd26, 27'h0000033e, 32'h00000400,
  1'd1,  5'd19, 27'h000001d4, 5'd11, 27'h00000294, 5'd4, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000038e, 5'd10, 27'h0000033e, 5'd14, 27'h000002e4, 32'h00000400,
  1'd1,  5'd17, 27'h000000f2, 5'd11, 27'h000000af, 5'd24, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000099, 5'd25, 27'h00000091, 5'd2, 27'h000001c6, 32'h00000400,
  1'd1,  5'd18, 27'h000002af, 5'd21, 27'h000001ba, 5'd13, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ba, 5'd24, 27'h000003c8, 5'd24, 27'h00000242, 32'h00000400,
  1'd1,  5'd27, 27'h000003cd, 5'd0, 27'h000003b8, 5'd2, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000035f, 5'd1, 27'h00000055, 5'd11, 27'h00000363, 32'h00000400,
  1'd1,  5'd25, 27'h00000365, 5'd0, 27'h000003ee, 5'd22, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000009a, 5'd12, 27'h00000323, 5'd2, 27'h00000169, 32'h00000400,
  1'd1,  5'd28, 27'h0000008d, 5'd12, 27'h000003dd, 5'd13, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000032b, 5'd10, 27'h000002b6, 5'd24, 27'h000003ea, 32'h00000400,
  1'd1,  5'd27, 27'h0000030c, 5'd24, 27'h0000039e, 5'd3, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001d8, 5'd25, 27'h0000001c, 5'd11, 27'h00000143, 32'h00000400,
  1'd1,  5'd27, 27'h00000031, 5'd25, 27'h000000da, 5'd25, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000206, 5'd3, 27'h00000381, 5'd2, 27'h000000ff, 32'h00000400,
  1'd1,  5'd8, 27'h00000071, 5'd5, 27'h0000006e, 5'd13, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000007e, 5'd0, 27'h0000016e, 5'd25, 27'h00000013, 32'h00000400,
  1'd1,  5'd5, 27'h00000343, 5'd14, 27'h000002dc, 5'd8, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003de, 5'd13, 27'h000000b2, 5'd16, 27'h0000037e, 32'h00000400,
  1'd1,  5'd7, 27'h000003a4, 5'd12, 27'h000001e8, 5'd28, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002e2, 5'd24, 27'h000003f3, 5'd9, 27'h0000004d, 32'h00000400,
  1'd1,  5'd6, 27'h000003dd, 5'd21, 27'h0000004e, 5'd18, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000257, 5'd20, 27'h000003cd, 5'd29, 27'h000001aa, 32'h00000400,
  1'd1,  5'd19, 27'h000001e8, 5'd2, 27'h00000215, 5'd4, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000156, 5'd3, 27'h0000039c, 5'd10, 27'h00000297, 32'h00000400,
  1'd1,  5'd20, 27'h00000029, 5'd2, 27'h000000bc, 5'd25, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000174, 5'd15, 27'h00000099, 5'd7, 27'h000000bd, 32'h00000400,
  1'd1,  5'd18, 27'h00000270, 5'd11, 27'h00000342, 5'd17, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d9, 5'd13, 27'h000001ca, 5'd29, 27'h00000357, 32'h00000400,
  1'd1,  5'd16, 27'h000001ca, 5'd23, 27'h00000152, 5'd6, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000029, 5'd22, 27'h000002e3, 5'd16, 27'h0000007b, 32'h00000400,
  1'd1,  5'd16, 27'h000002c0, 5'd23, 27'h00000312, 5'd26, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c3, 5'd0, 27'h00000241, 5'd9, 27'h000003f0, 32'h00000400,
  1'd1,  5'd30, 27'h00000044, 5'd2, 27'h000002f2, 5'd16, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003f0, 5'd2, 27'h000002ae, 5'd26, 27'h00000136, 32'h00000400,
  1'd1,  5'd28, 27'h000001c1, 5'd10, 27'h00000205, 5'd10, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002fe, 5'd15, 27'h00000199, 5'd19, 27'h000003db, 32'h00000400,
  1'd1,  5'd28, 27'h00000131, 5'd15, 27'h0000003e, 5'd29, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000231, 5'd21, 27'h000003a9, 5'd6, 27'h00000097, 32'h00000400,
  1'd1,  5'd30, 27'h000002f3, 5'd24, 27'h000000b5, 5'd16, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000265, 5'd25, 27'h00000320, 5'd30, 27'h000003f8, 32'h00000400,
  1'd1,  5'd8, 27'h00000153, 5'd8, 27'h000001e0, 5'd4, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000187, 5'd9, 27'h000001c1, 5'd14, 27'h00000355, 32'h00000400,
  1'd1,  5'd5, 27'h000002d6, 5'd9, 27'h000002a1, 5'd25, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000126, 5'd20, 27'h000000df, 5'd4, 27'h000001d5, 32'h00000400,
  1'd1,  5'd5, 27'h0000030b, 5'd17, 27'h000002fc, 5'd14, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e7, 5'd16, 27'h000003a5, 5'd24, 27'h000003bc, 32'h00000400,
  1'd1,  5'd5, 27'h00000342, 5'd29, 27'h00000217, 5'd2, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000037d, 5'd29, 27'h0000005a, 5'd11, 27'h0000038f, 32'h00000400,
  1'd1,  5'd9, 27'h00000252, 5'd28, 27'h000000b6, 5'd24, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000269, 5'd6, 27'h00000392, 5'd3, 27'h000001cd, 32'h00000400,
  1'd1,  5'd20, 27'h00000042, 5'd6, 27'h00000395, 5'd15, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019b, 5'd9, 27'h00000355, 5'd25, 27'h00000083, 32'h00000400,
  1'd1,  5'd17, 27'h0000012d, 5'd20, 27'h00000082, 5'd4, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000043, 5'd16, 27'h0000020c, 5'd11, 27'h000001d8, 32'h00000400,
  1'd1,  5'd17, 27'h000002cc, 5'd19, 27'h000003da, 5'd21, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003bb, 5'd27, 27'h000003cf, 5'd0, 27'h000001a8, 32'h00000400,
  1'd1,  5'd20, 27'h00000087, 5'd30, 27'h000003e9, 5'd11, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000323, 5'd27, 27'h000003c0, 5'd24, 27'h000000ed, 32'h00000400,
  1'd1,  5'd30, 27'h00000212, 5'd9, 27'h00000072, 5'd1, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000306, 5'd9, 27'h0000015c, 5'd10, 27'h0000019e, 32'h00000400,
  1'd1,  5'd30, 27'h00000084, 5'd9, 27'h00000270, 5'd24, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000140, 5'd15, 27'h000002b7, 5'd4, 27'h0000022b, 32'h00000400,
  1'd1,  5'd27, 27'h0000003d, 5'd15, 27'h0000021e, 5'd12, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000309, 5'd16, 27'h000000bb, 5'd24, 27'h00000218, 32'h00000400,
  1'd1,  5'd29, 27'h000002b8, 5'd29, 27'h00000087, 5'd2, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b9, 5'd30, 27'h00000372, 5'd13, 27'h000001a0, 32'h00000400,
  1'd1,  5'd25, 27'h000003fb, 5'd26, 27'h00000282, 5'd23, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000029b, 5'd6, 27'h000003ad, 5'd7, 27'h00000274, 32'h00000400,
  1'd1,  5'd9, 27'h0000023a, 5'd7, 27'h000002c7, 5'd18, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000026e, 5'd5, 27'h000003f6, 5'd27, 27'h0000036c, 32'h00000400,
  1'd1,  5'd5, 27'h0000023c, 5'd17, 27'h00000074, 5'd10, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ab, 5'd15, 27'h00000235, 5'd18, 27'h00000225, 32'h00000400,
  1'd1,  5'd7, 27'h0000025f, 5'd19, 27'h000001ec, 5'd29, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000234, 5'd26, 27'h00000142, 5'd7, 27'h00000031, 32'h00000400,
  1'd1,  5'd8, 27'h0000034b, 5'd27, 27'h0000031a, 5'd15, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b7, 5'd27, 27'h0000001a, 5'd30, 27'h000003d0, 32'h00000400,
  1'd1,  5'd17, 27'h00000149, 5'd8, 27'h00000015, 5'd9, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000104, 5'd5, 27'h000001f5, 5'd19, 27'h0000020d, 32'h00000400,
  1'd1,  5'd17, 27'h00000024, 5'd10, 27'h0000004b, 5'd28, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ae, 5'd18, 27'h0000021d, 5'd9, 27'h000001cc, 32'h00000400,
  1'd1,  5'd16, 27'h00000258, 5'd19, 27'h000000aa, 5'd16, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000115, 5'd18, 27'h00000244, 5'd28, 27'h000003c1, 32'h00000400,
  1'd1,  5'd16, 27'h0000022e, 5'd30, 27'h00000321, 5'd7, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000223, 5'd30, 27'h00000079, 5'd19, 27'h000000a7, 32'h00000400,
  1'd1,  5'd19, 27'h000002fd, 5'd27, 27'h00000282, 5'd27, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000025, 5'd9, 27'h00000235, 5'd5, 27'h00000251, 32'h00000400,
  1'd1,  5'd27, 27'h00000126, 5'd9, 27'h00000312, 5'd18, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000e1, 5'd9, 27'h000001b4, 5'd29, 27'h00000061, 32'h00000400,
  1'd1,  5'd28, 27'h000002b3, 5'd18, 27'h000000f8, 5'd6, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000011d, 5'd16, 27'h0000005d, 5'd18, 27'h000000b2, 32'h00000400,
  1'd1,  5'd29, 27'h00000167, 5'd17, 27'h0000034b, 5'd28, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e6, 5'd30, 27'h00000189, 5'd8, 27'h000003f0, 32'h00000400,
  1'd1,  5'd28, 27'h000003a8, 5'd28, 27'h000001f2, 5'd15, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000299, 5'd29, 27'h000002ac, 5'd26, 27'h00000036, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000034, 5'd3, 27'h0000032b, 5'd0, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000019d, 5'd4, 27'h0000032c, 5'd14, 27'h00000165, 32'h00000400,
  1'd1,  5'd0, 27'h000003e4, 5'd2, 27'h00000325, 5'd21, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ee, 5'd11, 27'h00000340, 5'd0, 27'h00000299, 32'h00000400,
  1'd1,  5'd4, 27'h000003b0, 5'd12, 27'h00000027, 5'd10, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000028f, 5'd13, 27'h000001b4, 5'd23, 27'h00000360, 32'h00000400,
  1'd1,  5'd3, 27'h00000171, 5'd20, 27'h000002f2, 5'd2, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000025b, 5'd21, 27'h00000301, 5'd14, 27'h0000027e, 32'h00000400,
  1'd1,  5'd0, 27'h0000000a, 5'd22, 27'h000001cb, 5'd21, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000033e, 5'd2, 27'h000000fa, 5'd4, 27'h000003fc, 32'h00000400,
  1'd1,  5'd10, 27'h00000361, 5'd2, 27'h000003a4, 5'd12, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000097, 5'd1, 27'h0000009a, 5'd20, 27'h000003da, 32'h00000400,
  1'd1,  5'd11, 27'h0000035d, 5'd15, 27'h0000007f, 5'd0, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000204, 5'd11, 27'h0000038c, 5'd12, 27'h0000021c, 32'h00000400,
  1'd1,  5'd12, 27'h00000029, 5'd13, 27'h000003b9, 5'd25, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000190, 5'd23, 27'h00000359, 5'd0, 27'h00000340, 32'h00000400,
  1'd1,  5'd14, 27'h000002f7, 5'd23, 27'h0000029e, 5'd11, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000132, 5'd24, 27'h000002fa, 5'd21, 27'h000001d1, 32'h00000400,
  1'd1,  5'd24, 27'h000002b4, 5'd2, 27'h0000034c, 5'd2, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002dd, 5'd2, 27'h0000010e, 5'd14, 27'h000003e7, 32'h00000400,
  1'd1,  5'd23, 27'h00000218, 5'd4, 27'h00000222, 5'd24, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000184, 5'd11, 27'h00000101, 5'd0, 27'h0000010d, 32'h00000400,
  1'd1,  5'd24, 27'h0000035a, 5'd15, 27'h0000019b, 5'd15, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c8, 5'd11, 27'h0000022d, 5'd21, 27'h0000031f, 32'h00000400,
  1'd1,  5'd21, 27'h00000201, 5'd23, 27'h00000231, 5'd2, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001c, 5'd22, 27'h0000002b, 5'd12, 27'h00000396, 32'h00000400,
  1'd1,  5'd24, 27'h00000242, 5'd25, 27'h00000227, 5'd22, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002eb, 5'd2, 27'h0000005e, 5'd10, 27'h00000132, 32'h00000400,
  1'd1,  5'd1, 27'h000000d9, 5'd3, 27'h0000010f, 5'd16, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000142, 5'd3, 27'h00000177, 5'd26, 27'h000000c5, 32'h00000400,
  1'd1,  5'd0, 27'h0000017e, 5'd13, 27'h000001f0, 5'd7, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000029f, 5'd13, 27'h000001f0, 5'd17, 27'h00000085, 32'h00000400,
  1'd1,  5'd1, 27'h0000016b, 5'd10, 27'h000002e8, 5'd25, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d5, 5'd23, 27'h0000027f, 5'd6, 27'h000003b1, 32'h00000400,
  1'd1,  5'd2, 27'h000003e3, 5'd24, 27'h00000315, 5'd16, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000158, 5'd20, 27'h000003f0, 5'd25, 27'h00000378, 32'h00000400,
  1'd1,  5'd14, 27'h000002f4, 5'd1, 27'h00000167, 5'd9, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000190, 5'd1, 27'h00000118, 5'd16, 27'h000001f3, 32'h00000400,
  1'd1,  5'd10, 27'h0000039a, 5'd4, 27'h000001aa, 5'd29, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000181, 5'd14, 27'h000003f8, 5'd9, 27'h0000012c, 32'h00000400,
  1'd1,  5'd14, 27'h0000005f, 5'd13, 27'h000002df, 5'd19, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000da, 5'd10, 27'h000002e4, 5'd28, 27'h0000037c, 32'h00000400,
  1'd1,  5'd14, 27'h000002a8, 5'd25, 27'h000002e3, 5'd7, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000314, 5'd23, 27'h0000011c, 5'd18, 27'h00000105, 32'h00000400,
  1'd1,  5'd13, 27'h000002ed, 5'd22, 27'h00000275, 5'd27, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f1, 5'd2, 27'h00000118, 5'd8, 27'h000000c7, 32'h00000400,
  1'd1,  5'd21, 27'h0000013f, 5'd1, 27'h00000372, 5'd20, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002bb, 5'd1, 27'h00000339, 5'd28, 27'h00000226, 32'h00000400,
  1'd1,  5'd24, 27'h00000349, 5'd11, 27'h000003c6, 5'd6, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002ae, 5'd11, 27'h00000273, 5'd18, 27'h00000391, 32'h00000400,
  1'd1,  5'd21, 27'h000003a6, 5'd11, 27'h000002f6, 5'd27, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021d, 5'd22, 27'h00000316, 5'd5, 27'h000002cf, 32'h00000400,
  1'd1,  5'd24, 27'h00000346, 5'd22, 27'h0000028b, 5'd16, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000167, 5'd22, 27'h0000039b, 5'd28, 27'h0000008e, 32'h00000400,
  1'd1,  5'd3, 27'h0000007b, 5'd8, 27'h0000024e, 5'd2, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000011d, 5'd5, 27'h000003b2, 5'd14, 27'h0000006b, 32'h00000400,
  1'd1,  5'd4, 27'h0000027c, 5'd5, 27'h000000c6, 5'd21, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003b0, 5'd19, 27'h00000025, 5'd0, 27'h000001ee, 32'h00000400,
  1'd1,  5'd4, 27'h000001db, 5'd19, 27'h00000093, 5'd10, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003df, 5'd20, 27'h00000272, 5'd22, 27'h0000029c, 32'h00000400,
  1'd1,  5'd5, 27'h0000004e, 5'd26, 27'h000000f7, 5'd4, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000085, 5'd27, 27'h00000149, 5'd12, 27'h0000007c, 32'h00000400,
  1'd1,  5'd2, 27'h00000321, 5'd26, 27'h000000e6, 5'd23, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002d4, 5'd7, 27'h000003c6, 5'd5, 27'h0000007d, 32'h00000400,
  1'd1,  5'd14, 27'h00000021, 5'd5, 27'h00000153, 5'd12, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000000a, 5'd5, 27'h00000388, 5'd22, 27'h000003e5, 32'h00000400,
  1'd1,  5'd11, 27'h00000123, 5'd16, 27'h00000132, 5'd1, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000014, 5'd20, 27'h000001c0, 5'd14, 27'h0000011d, 32'h00000400,
  1'd1,  5'd10, 27'h00000178, 5'd15, 27'h0000021c, 5'd25, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001fa, 5'd26, 27'h00000234, 5'd1, 27'h000001d6, 32'h00000400,
  1'd1,  5'd10, 27'h00000178, 5'd26, 27'h00000198, 5'd14, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001da, 5'd30, 27'h0000027e, 5'd22, 27'h000002c4, 32'h00000400,
  1'd1,  5'd24, 27'h0000035f, 5'd9, 27'h000003f8, 5'd4, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000130, 5'd8, 27'h000003c1, 5'd12, 27'h00000302, 32'h00000400,
  1'd1,  5'd23, 27'h0000033d, 5'd8, 27'h000003f2, 5'd23, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000d6, 5'd16, 27'h00000207, 5'd0, 27'h0000035e, 32'h00000400,
  1'd1,  5'd22, 27'h00000310, 5'd16, 27'h00000334, 5'd12, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000023f, 5'd15, 27'h00000212, 5'd23, 27'h00000062, 32'h00000400,
  1'd1,  5'd23, 27'h00000331, 5'd30, 27'h0000010a, 5'd3, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000027d, 5'd29, 27'h0000029e, 5'd12, 27'h0000026a, 32'h00000400,
  1'd1,  5'd25, 27'h0000030a, 5'd27, 27'h0000004e, 5'd23, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000130, 5'd7, 27'h000003e1, 5'd6, 27'h000000ed, 32'h00000400,
  1'd1,  5'd3, 27'h000002e7, 5'd5, 27'h00000365, 5'd16, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000158, 5'd5, 27'h00000253, 5'd30, 27'h0000026d, 32'h00000400,
  1'd1,  5'd2, 27'h000002ad, 5'd17, 27'h00000197, 5'd9, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b4, 5'd17, 27'h000002c9, 5'd18, 27'h000003a7, 32'h00000400,
  1'd1,  5'd2, 27'h000000cb, 5'd19, 27'h000000ef, 5'd26, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d2, 5'd27, 27'h00000206, 5'd7, 27'h0000029c, 32'h00000400,
  1'd1,  5'd0, 27'h00000010, 5'd28, 27'h000003fe, 5'd17, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a6, 5'd28, 27'h000002c8, 5'd30, 27'h000000f6, 32'h00000400,
  1'd1,  5'd15, 27'h00000003, 5'd9, 27'h00000273, 5'd7, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000001b, 5'd6, 27'h0000018b, 5'd15, 27'h00000285, 32'h00000400,
  1'd1,  5'd12, 27'h00000178, 5'd9, 27'h00000184, 5'd28, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000258, 5'd20, 27'h000000f2, 5'd9, 27'h0000029e, 32'h00000400,
  1'd1,  5'd10, 27'h000002fd, 5'd15, 27'h000002f5, 5'd17, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000096, 5'd18, 27'h00000279, 5'd27, 27'h000003e8, 32'h00000400,
  1'd1,  5'd12, 27'h00000057, 5'd26, 27'h0000003e, 5'd7, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000a9, 5'd26, 27'h000002f3, 5'd19, 27'h000000f1, 32'h00000400,
  1'd1,  5'd11, 27'h000002c4, 5'd30, 27'h0000034c, 5'd29, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f6, 5'd9, 27'h0000001e, 5'd6, 27'h00000111, 32'h00000400,
  1'd1,  5'd21, 27'h0000002a, 5'd8, 27'h000002e6, 5'd17, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000393, 5'd7, 27'h00000105, 5'd27, 27'h0000024f, 32'h00000400,
  1'd1,  5'd23, 27'h0000026c, 5'd17, 27'h0000036d, 5'd9, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000190, 5'd17, 27'h00000379, 5'd17, 27'h00000234, 32'h00000400,
  1'd1,  5'd24, 27'h0000017e, 5'd20, 27'h000001f4, 5'd28, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b1, 5'd28, 27'h0000028d, 5'd8, 27'h0000001e, 32'h00000400,
  1'd1,  5'd24, 27'h00000353, 5'd26, 27'h000000b7, 5'd15, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000032, 5'd29, 27'h000002a4, 5'd27, 27'h00000116, 32'h00000400,
  1'd1,  5'd8, 27'h000000a6, 5'd1, 27'h000000b9, 5'd7, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000306, 5'd3, 27'h000003da, 5'd17, 27'h000002b6, 32'h00000400,
  1'd1,  5'd5, 27'h000001c1, 5'd3, 27'h00000236, 5'd28, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002c8, 5'd15, 27'h00000179, 5'd0, 27'h00000388, 32'h00000400,
  1'd1,  5'd5, 27'h000001e5, 5'd15, 27'h00000092, 5'd11, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002bd, 5'd11, 27'h000000ca, 5'd23, 27'h0000018b, 32'h00000400,
  1'd1,  5'd5, 27'h0000019a, 5'd24, 27'h00000121, 5'd1, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002c7, 5'd22, 27'h000001de, 5'd14, 27'h0000032d, 32'h00000400,
  1'd1,  5'd8, 27'h00000142, 5'd25, 27'h000001bb, 5'd25, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000111, 5'd0, 27'h000002ec, 5'd7, 27'h000000dd, 32'h00000400,
  1'd1,  5'd16, 27'h00000297, 5'd1, 27'h00000034, 5'd18, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001d4, 5'd3, 27'h00000398, 5'd29, 27'h00000128, 32'h00000400,
  1'd1,  5'd18, 27'h000003d3, 5'd12, 27'h00000295, 5'd3, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000001f, 5'd10, 27'h00000217, 5'd12, 27'h000001cf, 32'h00000400,
  1'd1,  5'd16, 27'h000002dd, 5'd12, 27'h0000024c, 5'd22, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000338, 5'd22, 27'h00000233, 5'd4, 27'h0000031f, 32'h00000400,
  1'd1,  5'd18, 27'h00000257, 5'd24, 27'h000003ab, 5'd13, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c4, 5'd22, 27'h00000369, 5'd23, 27'h00000136, 32'h00000400,
  1'd1,  5'd27, 27'h000000d0, 5'd1, 27'h00000294, 5'd4, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000023c, 5'd1, 27'h0000000f, 5'd11, 27'h00000018, 32'h00000400,
  1'd1,  5'd30, 27'h000000d1, 5'd4, 27'h0000023a, 5'd24, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f7, 5'd14, 27'h0000008f, 5'd1, 27'h000001ce, 32'h00000400,
  1'd1,  5'd26, 27'h00000066, 5'd14, 27'h00000126, 5'd12, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ef, 5'd10, 27'h00000270, 5'd25, 27'h00000317, 32'h00000400,
  1'd1,  5'd25, 27'h00000380, 5'd25, 27'h00000247, 5'd0, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a7, 5'd21, 27'h000001cf, 5'd12, 27'h000000cb, 32'h00000400,
  1'd1,  5'd28, 27'h0000037a, 5'd24, 27'h00000207, 5'd23, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000aa, 5'd0, 27'h00000223, 5'd2, 27'h00000332, 32'h00000400,
  1'd1,  5'd7, 27'h00000303, 5'd3, 27'h0000036d, 5'd14, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000185, 5'd0, 27'h00000132, 5'd21, 27'h000001c7, 32'h00000400,
  1'd1,  5'd8, 27'h00000197, 5'd11, 27'h00000136, 5'd8, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000285, 5'd10, 27'h000002e8, 5'd19, 27'h000002da, 32'h00000400,
  1'd1,  5'd9, 27'h000000a7, 5'd10, 27'h00000174, 5'd27, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d3, 5'd22, 27'h0000012d, 5'd7, 27'h00000324, 32'h00000400,
  1'd1,  5'd10, 27'h0000007d, 5'd21, 27'h00000049, 5'd17, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c9, 5'd20, 27'h00000359, 5'd26, 27'h00000342, 32'h00000400,
  1'd1,  5'd20, 27'h00000068, 5'd1, 27'h00000300, 5'd2, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003df, 5'd0, 27'h00000069, 5'd12, 27'h00000141, 32'h00000400,
  1'd1,  5'd20, 27'h0000007d, 5'd0, 27'h00000112, 5'd20, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c3, 5'd14, 27'h000000e0, 5'd9, 27'h000003ad, 32'h00000400,
  1'd1,  5'd19, 27'h00000382, 5'd14, 27'h00000217, 5'd17, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000219, 5'd10, 27'h00000360, 5'd27, 27'h0000000f, 32'h00000400,
  1'd1,  5'd16, 27'h000001a2, 5'd21, 27'h000003b4, 5'd9, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025a, 5'd21, 27'h00000018, 5'd18, 27'h00000145, 32'h00000400,
  1'd1,  5'd19, 27'h00000214, 5'd22, 27'h0000001d, 5'd27, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000048, 5'd1, 27'h00000304, 5'd7, 27'h00000146, 32'h00000400,
  1'd1,  5'd29, 27'h000002ce, 5'd0, 27'h000000f1, 5'd19, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024d, 5'd3, 27'h00000079, 5'd30, 27'h00000024, 32'h00000400,
  1'd1,  5'd27, 27'h000003a3, 5'd12, 27'h0000009a, 5'd9, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ae, 5'd14, 27'h00000388, 5'd16, 27'h000003ed, 32'h00000400,
  1'd1,  5'd27, 27'h00000170, 5'd11, 27'h00000135, 5'd28, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000138, 5'd25, 27'h000002fd, 5'd5, 27'h000003cc, 32'h00000400,
  1'd1,  5'd28, 27'h000001f4, 5'd22, 27'h0000036e, 5'd17, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000120, 5'd22, 27'h000003d6, 5'd30, 27'h00000168, 32'h00000400,
  1'd1,  5'd6, 27'h00000239, 5'd7, 27'h000000a9, 5'd1, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000350, 5'd6, 27'h00000004, 5'd10, 27'h000003f4, 32'h00000400,
  1'd1,  5'd6, 27'h0000014b, 5'd6, 27'h00000256, 5'd24, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000130, 5'd16, 27'h0000016e, 5'd2, 27'h0000039c, 32'h00000400,
  1'd1,  5'd10, 27'h0000002b, 5'd20, 27'h00000283, 5'd14, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000167, 5'd20, 27'h000001e6, 5'd25, 27'h00000134, 32'h00000400,
  1'd1,  5'd5, 27'h000003f2, 5'd29, 27'h000001c2, 5'd1, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001b5, 5'd26, 27'h00000260, 5'd11, 27'h00000372, 32'h00000400,
  1'd1,  5'd9, 27'h00000175, 5'd25, 27'h00000387, 5'd23, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000094, 5'd6, 27'h000003fe, 5'd3, 27'h0000002f, 32'h00000400,
  1'd1,  5'd20, 27'h000000a1, 5'd5, 27'h000000fc, 5'd11, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003b6, 5'd6, 27'h00000177, 5'd24, 27'h00000309, 32'h00000400,
  1'd1,  5'd19, 27'h000002d1, 5'd18, 27'h000001e8, 5'd2, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000013b, 5'd16, 27'h000000d7, 5'd10, 27'h000001e2, 32'h00000400,
  1'd1,  5'd19, 27'h0000009f, 5'd16, 27'h00000100, 5'd23, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001cc, 5'd25, 27'h0000036a, 5'd3, 27'h000003e4, 32'h00000400,
  1'd1,  5'd15, 27'h00000373, 5'd29, 27'h00000055, 5'd11, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000308, 5'd28, 27'h00000373, 5'd21, 27'h0000005d, 32'h00000400,
  1'd1,  5'd28, 27'h0000004c, 5'd9, 27'h000000eb, 5'd0, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000021c, 5'd8, 27'h00000242, 5'd11, 27'h0000000e, 32'h00000400,
  1'd1,  5'd27, 27'h0000007e, 5'd7, 27'h000001c1, 5'd21, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c5, 5'd19, 27'h000000ad, 5'd0, 27'h000001b2, 32'h00000400,
  1'd1,  5'd26, 27'h000001f1, 5'd17, 27'h00000359, 5'd11, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000014b, 5'd18, 27'h0000018e, 5'd23, 27'h00000119, 32'h00000400,
  1'd1,  5'd26, 27'h000001ef, 5'd28, 27'h00000108, 5'd5, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000001e, 5'd27, 27'h000000fd, 5'd11, 27'h000003c4, 32'h00000400,
  1'd1,  5'd25, 27'h0000037d, 5'd29, 27'h0000032d, 5'd22, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000017f, 5'd9, 27'h00000005, 5'd7, 27'h000000ca, 32'h00000400,
  1'd1,  5'd10, 27'h0000008d, 5'd8, 27'h0000009b, 5'd16, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000025a, 5'd5, 27'h000002d6, 5'd29, 27'h00000296, 32'h00000400,
  1'd1,  5'd10, 27'h00000111, 5'd20, 27'h000001b6, 5'd9, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003f, 5'd19, 27'h00000196, 5'd19, 27'h00000172, 32'h00000400,
  1'd1,  5'd10, 27'h00000011, 5'd17, 27'h00000342, 5'd29, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000277, 5'd26, 27'h00000210, 5'd5, 27'h000000b3, 32'h00000400,
  1'd1,  5'd7, 27'h00000076, 5'd30, 27'h000003fe, 5'd15, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c2, 5'd30, 27'h0000011c, 5'd29, 27'h000002de, 32'h00000400,
  1'd1,  5'd20, 27'h0000024a, 5'd5, 27'h00000163, 5'd6, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003d3, 5'd5, 27'h000001e1, 5'd20, 27'h000002aa, 32'h00000400,
  1'd1,  5'd17, 27'h0000020f, 5'd7, 27'h000002b9, 5'd29, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000df, 5'd17, 27'h0000020e, 5'd9, 27'h00000101, 32'h00000400,
  1'd1,  5'd15, 27'h00000297, 5'd19, 27'h00000170, 5'd16, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a6, 5'd18, 27'h00000087, 5'd30, 27'h000001d0, 32'h00000400,
  1'd1,  5'd16, 27'h00000281, 5'd27, 27'h000003a1, 5'd9, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000023d, 5'd28, 27'h000002d0, 5'd16, 27'h00000000, 32'h00000400,
  1'd1,  5'd17, 27'h0000024f, 5'd29, 27'h00000175, 5'd29, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000039c, 5'd5, 27'h0000029d, 5'd8, 27'h0000007a, 32'h00000400,
  1'd1,  5'd29, 27'h000000ac, 5'd8, 27'h0000004f, 5'd16, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000250, 5'd9, 27'h00000137, 5'd29, 27'h00000040, 32'h00000400,
  1'd1,  5'd29, 27'h000001e9, 5'd15, 27'h0000037f, 5'd7, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000ea, 5'd16, 27'h000003a5, 5'd19, 27'h000003e2, 32'h00000400,
  1'd1,  5'd27, 27'h00000045, 5'd17, 27'h00000252, 5'd29, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000010e, 5'd30, 27'h0000007d, 5'd6, 27'h00000293, 32'h00000400,
  1'd1,  5'd29, 27'h000003f7, 5'd26, 27'h00000012, 5'd16, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003af, 5'd30, 27'h00000076, 5'd26, 27'h00000364, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000292, 5'd4, 27'h000003be, 5'd4, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000259, 5'd3, 27'h00000179, 5'd13, 27'h00000293, 32'h00000400,
  1'd1,  5'd3, 27'h00000139, 5'd1, 27'h0000013c, 5'd22, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000038, 5'd11, 27'h0000016f, 5'd3, 27'h0000016d, 32'h00000400,
  1'd1,  5'd0, 27'h0000038d, 5'd11, 27'h00000083, 5'd11, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d5, 5'd11, 27'h00000325, 5'd24, 27'h0000024b, 32'h00000400,
  1'd1,  5'd2, 27'h0000034c, 5'd21, 27'h00000067, 5'd2, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000038f, 5'd25, 27'h0000004f, 5'd13, 27'h000003b0, 32'h00000400,
  1'd1,  5'd3, 27'h000002ea, 5'd20, 27'h000003a7, 5'd23, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e4, 5'd1, 27'h00000268, 5'd0, 27'h0000036e, 32'h00000400,
  1'd1,  5'd12, 27'h00000109, 5'd3, 27'h0000004d, 5'd15, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000340, 5'd3, 27'h0000001c, 5'd23, 27'h00000355, 32'h00000400,
  1'd1,  5'd12, 27'h0000023d, 5'd15, 27'h0000012e, 5'd0, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000011, 5'd11, 27'h00000132, 5'd15, 27'h00000082, 32'h00000400,
  1'd1,  5'd11, 27'h000000fe, 5'd12, 27'h000001a3, 5'd23, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000337, 5'd22, 27'h00000357, 5'd0, 27'h00000146, 32'h00000400,
  1'd1,  5'd14, 27'h0000039b, 5'd25, 27'h000002c9, 5'd12, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a2, 5'd24, 27'h00000179, 5'd20, 27'h00000311, 32'h00000400,
  1'd1,  5'd21, 27'h000001d9, 5'd1, 27'h0000028a, 5'd4, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000037a, 5'd5, 27'h0000008b, 5'd11, 27'h00000313, 32'h00000400,
  1'd1,  5'd23, 27'h00000154, 5'd3, 27'h000002d2, 5'd25, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000037d, 5'd14, 27'h000000cf, 5'd3, 27'h0000039f, 32'h00000400,
  1'd1,  5'd23, 27'h0000005d, 5'd10, 27'h00000244, 5'd14, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003eb, 5'd11, 27'h000001fb, 5'd21, 27'h0000010e, 32'h00000400,
  1'd1,  5'd25, 27'h000000ca, 5'd24, 27'h0000028e, 5'd3, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d7, 5'd24, 27'h00000021, 5'd11, 27'h00000284, 32'h00000400,
  1'd1,  5'd24, 27'h00000050, 5'd25, 27'h00000181, 5'd25, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001bc, 5'd0, 27'h000003d5, 5'd9, 27'h000002fe, 32'h00000400,
  1'd1,  5'd3, 27'h0000028c, 5'd2, 27'h000002c0, 5'd18, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000021e, 5'd4, 27'h00000133, 5'd28, 27'h0000020f, 32'h00000400,
  1'd1,  5'd4, 27'h0000031f, 5'd12, 27'h00000113, 5'd9, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002bc, 5'd14, 27'h00000373, 5'd17, 27'h00000318, 32'h00000400,
  1'd1,  5'd1, 27'h000001ca, 5'd12, 27'h00000342, 5'd29, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000030b, 5'd22, 27'h00000172, 5'd7, 27'h000000c2, 32'h00000400,
  1'd1,  5'd4, 27'h0000016d, 5'd22, 27'h000002ed, 5'd19, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000032f, 5'd23, 27'h0000015a, 5'd28, 27'h00000335, 32'h00000400,
  1'd1,  5'd13, 27'h00000172, 5'd3, 27'h00000057, 5'd9, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000036, 5'd5, 27'h0000004e, 5'd20, 27'h0000026f, 32'h00000400,
  1'd1,  5'd11, 27'h000002e4, 5'd1, 27'h0000004e, 5'd29, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000126, 5'd15, 27'h00000053, 5'd9, 27'h0000015f, 32'h00000400,
  1'd1,  5'd12, 27'h00000381, 5'd12, 27'h00000194, 5'd20, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000061, 5'd12, 27'h000003bb, 5'd27, 27'h000003be, 32'h00000400,
  1'd1,  5'd14, 27'h000002b4, 5'd24, 27'h0000029a, 5'd9, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f0, 5'd25, 27'h0000012c, 5'd19, 27'h0000015d, 32'h00000400,
  1'd1,  5'd12, 27'h000002ae, 5'd25, 27'h0000017d, 5'd29, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000190, 5'd2, 27'h00000054, 5'd6, 27'h0000010f, 32'h00000400,
  1'd1,  5'd25, 27'h000002f6, 5'd4, 27'h00000372, 5'd16, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000017c, 5'd2, 27'h0000037d, 5'd30, 27'h00000188, 32'h00000400,
  1'd1,  5'd24, 27'h00000352, 5'd14, 27'h000000d5, 5'd5, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000029c, 5'd13, 27'h00000302, 5'd16, 27'h000000a4, 32'h00000400,
  1'd1,  5'd22, 27'h000000cf, 5'd13, 27'h0000033b, 5'd26, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000057, 5'd23, 27'h00000307, 5'd5, 27'h0000012e, 32'h00000400,
  1'd1,  5'd22, 27'h00000035, 5'd24, 27'h0000006b, 5'd18, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e6, 5'd25, 27'h000001d7, 5'd27, 27'h00000314, 32'h00000400,
  1'd1,  5'd1, 27'h0000028a, 5'd8, 27'h000002b2, 5'd1, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000012f, 5'd6, 27'h000002df, 5'd10, 27'h00000252, 32'h00000400,
  1'd1,  5'd2, 27'h0000036a, 5'd10, 27'h00000096, 5'd22, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000111, 5'd18, 27'h000001ed, 5'd5, 27'h00000029, 32'h00000400,
  1'd1,  5'd2, 27'h0000013a, 5'd16, 27'h00000306, 5'd10, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000259, 5'd19, 27'h000001ca, 5'd24, 27'h000001c0, 32'h00000400,
  1'd1,  5'd2, 27'h0000017e, 5'd27, 27'h000000fb, 5'd1, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000033f, 5'd29, 27'h0000003c, 5'd13, 27'h0000016b, 32'h00000400,
  1'd1,  5'd0, 27'h00000385, 5'd30, 27'h000002a7, 5'd24, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c4, 5'd5, 27'h00000135, 5'd5, 27'h00000035, 32'h00000400,
  1'd1,  5'd11, 27'h0000026f, 5'd6, 27'h0000031d, 5'd11, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003cf, 5'd9, 27'h00000234, 5'd21, 27'h00000176, 32'h00000400,
  1'd1,  5'd15, 27'h000000fa, 5'd18, 27'h0000020d, 5'd1, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000088, 5'd19, 27'h00000058, 5'd15, 27'h00000135, 32'h00000400,
  1'd1,  5'd14, 27'h000003f1, 5'd19, 27'h00000253, 5'd24, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003fd, 5'd29, 27'h0000017a, 5'd0, 27'h0000007e, 32'h00000400,
  1'd1,  5'd14, 27'h0000031c, 5'd26, 27'h0000023d, 5'd12, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000343, 5'd27, 27'h00000303, 5'd21, 27'h00000061, 32'h00000400,
  1'd1,  5'd24, 27'h0000013e, 5'd7, 27'h000000e3, 5'd5, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003e1, 5'd8, 27'h00000330, 5'd13, 27'h000002e4, 32'h00000400,
  1'd1,  5'd24, 27'h000000d5, 5'd7, 27'h000000b3, 5'd22, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006a, 5'd19, 27'h0000037d, 5'd3, 27'h00000248, 32'h00000400,
  1'd1,  5'd21, 27'h000003c1, 5'd16, 27'h000001b3, 5'd12, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002f7, 5'd17, 27'h00000313, 5'd23, 27'h000001e4, 32'h00000400,
  1'd1,  5'd24, 27'h00000018, 5'd26, 27'h00000376, 5'd4, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003bd, 5'd29, 27'h00000052, 5'd12, 27'h0000020c, 32'h00000400,
  1'd1,  5'd21, 27'h0000033e, 5'd28, 27'h0000013e, 5'd22, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039d, 5'd7, 27'h000000a5, 5'd6, 27'h00000051, 32'h00000400,
  1'd1,  5'd4, 27'h000002ac, 5'd8, 27'h000002d0, 5'd17, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000004f, 5'd8, 27'h000003ab, 5'd30, 27'h00000370, 32'h00000400,
  1'd1,  5'd0, 27'h00000275, 5'd17, 27'h00000221, 5'd8, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000007e, 5'd18, 27'h000001d8, 5'd15, 27'h0000037c, 32'h00000400,
  1'd1,  5'd1, 27'h0000010d, 5'd19, 27'h000000bf, 5'd29, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000024a, 5'd26, 27'h00000215, 5'd7, 27'h00000232, 32'h00000400,
  1'd1,  5'd2, 27'h00000148, 5'd30, 27'h00000037, 5'd16, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f1, 5'd27, 27'h000000ab, 5'd28, 27'h000002f3, 32'h00000400,
  1'd1,  5'd14, 27'h000003e2, 5'd7, 27'h00000065, 5'd10, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001bc, 5'd5, 27'h000002eb, 5'd17, 27'h00000233, 32'h00000400,
  1'd1,  5'd11, 27'h00000013, 5'd6, 27'h00000088, 5'd30, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000242, 5'd17, 27'h000000e3, 5'd7, 27'h0000005b, 32'h00000400,
  1'd1,  5'd12, 27'h000000d4, 5'd18, 27'h000000c2, 5'd18, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000019d, 5'd18, 27'h0000012a, 5'd29, 27'h0000014e, 32'h00000400,
  1'd1,  5'd13, 27'h000001ae, 5'd27, 27'h00000044, 5'd7, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000009, 5'd26, 27'h000001e8, 5'd17, 27'h000001d4, 32'h00000400,
  1'd1,  5'd15, 27'h00000183, 5'd26, 27'h000001a6, 5'd30, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e6, 5'd5, 27'h0000024f, 5'd5, 27'h000001f3, 32'h00000400,
  1'd1,  5'd25, 27'h000002ac, 5'd7, 27'h00000013, 5'd20, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000030c, 5'd8, 27'h00000369, 5'd27, 27'h00000276, 32'h00000400,
  1'd1,  5'd21, 27'h0000008f, 5'd16, 27'h00000218, 5'd9, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000005f, 5'd18, 27'h000003bb, 5'd20, 27'h0000000d, 32'h00000400,
  1'd1,  5'd23, 27'h0000027d, 5'd17, 27'h000003ff, 5'd30, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002dd, 5'd29, 27'h000000b9, 5'd9, 27'h00000309, 32'h00000400,
  1'd1,  5'd23, 27'h000002d8, 5'd27, 27'h000001ff, 5'd19, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d7, 5'd28, 27'h000000b1, 5'd26, 27'h000002cd, 32'h00000400,
  1'd1,  5'd8, 27'h000003eb, 5'd3, 27'h00000115, 5'd8, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000185, 5'd2, 27'h0000005e, 5'd16, 27'h00000166, 32'h00000400,
  1'd1,  5'd9, 27'h00000036, 5'd1, 27'h0000024f, 5'd27, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000075, 5'd13, 27'h000000b2, 5'd0, 27'h00000395, 32'h00000400,
  1'd1,  5'd6, 27'h000000ff, 5'd13, 27'h00000300, 5'd14, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000063, 5'd15, 27'h00000132, 5'd23, 27'h000001ef, 32'h00000400,
  1'd1,  5'd7, 27'h0000017e, 5'd21, 27'h000000f1, 5'd3, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000089, 5'd24, 27'h0000010b, 5'd14, 27'h00000004, 32'h00000400,
  1'd1,  5'd7, 27'h0000002a, 5'd23, 27'h00000246, 5'd21, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000037c, 5'd1, 27'h00000217, 5'd8, 27'h000002b2, 32'h00000400,
  1'd1,  5'd19, 27'h000003a6, 5'd3, 27'h000002a0, 5'd15, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d3, 5'd5, 27'h00000080, 5'd29, 27'h00000005, 32'h00000400,
  1'd1,  5'd20, 27'h00000115, 5'd15, 27'h00000191, 5'd3, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003a0, 5'd11, 27'h00000148, 5'd10, 27'h0000032b, 32'h00000400,
  1'd1,  5'd20, 27'h0000027b, 5'd15, 27'h00000131, 5'd23, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002b5, 5'd22, 27'h00000188, 5'd1, 27'h0000011b, 32'h00000400,
  1'd1,  5'd17, 27'h0000017d, 5'd23, 27'h000002be, 5'd10, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000103, 5'd24, 27'h00000271, 5'd24, 27'h00000132, 32'h00000400,
  1'd1,  5'd29, 27'h000002d4, 5'd2, 27'h000003bb, 5'd1, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000d9, 5'd3, 27'h0000003c, 5'd13, 27'h00000354, 32'h00000400,
  1'd1,  5'd28, 27'h000002c7, 5'd3, 27'h000001f6, 5'd22, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000072, 5'd12, 27'h00000032, 5'd1, 27'h00000023, 32'h00000400,
  1'd1,  5'd26, 27'h000000b2, 5'd14, 27'h00000243, 5'd15, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000cb, 5'd13, 27'h00000107, 5'd20, 27'h000002ab, 32'h00000400,
  1'd1,  5'd27, 27'h0000039b, 5'd22, 27'h000000b3, 5'd0, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000398, 5'd25, 27'h00000047, 5'd14, 27'h00000169, 32'h00000400,
  1'd1,  5'd30, 27'h0000030e, 5'd25, 27'h00000047, 5'd20, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000021, 5'd1, 27'h00000025, 5'd3, 27'h00000006, 32'h00000400,
  1'd1,  5'd5, 27'h000000d3, 5'd0, 27'h000002e1, 5'd14, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000212, 5'd1, 27'h000001d8, 5'd23, 27'h00000257, 32'h00000400,
  1'd1,  5'd9, 27'h000003e8, 5'd15, 27'h000000cd, 5'd7, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000288, 5'd15, 27'h00000089, 5'd18, 27'h0000017c, 32'h00000400,
  1'd1,  5'd5, 27'h00000280, 5'd10, 27'h0000017d, 5'd28, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000182, 5'd25, 27'h000002de, 5'd6, 27'h00000067, 32'h00000400,
  1'd1,  5'd8, 27'h00000032, 5'd23, 27'h000003af, 5'd19, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000004, 5'd21, 27'h000001d3, 5'd30, 27'h00000205, 32'h00000400,
  1'd1,  5'd19, 27'h00000237, 5'd0, 27'h00000089, 5'd3, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ff, 5'd5, 27'h00000076, 5'd11, 27'h0000008c, 32'h00000400,
  1'd1,  5'd20, 27'h000001fd, 5'd4, 27'h0000007d, 5'd23, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ff, 5'd12, 27'h0000022e, 5'd7, 27'h0000032e, 32'h00000400,
  1'd1,  5'd18, 27'h0000018d, 5'd14, 27'h00000315, 5'd17, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000132, 5'd14, 27'h000000ab, 5'd25, 27'h000003a1, 32'h00000400,
  1'd1,  5'd20, 27'h0000010e, 5'd20, 27'h000002c0, 5'd6, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000257, 5'd24, 27'h00000204, 5'd18, 27'h000001fc, 32'h00000400,
  1'd1,  5'd15, 27'h00000397, 5'd20, 27'h00000324, 5'd29, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001cd, 5'd2, 27'h00000081, 5'd5, 27'h00000202, 32'h00000400,
  1'd1,  5'd30, 27'h000001bb, 5'd1, 27'h0000037e, 5'd19, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003c2, 5'd2, 27'h000002cf, 5'd26, 27'h00000187, 32'h00000400,
  1'd1,  5'd26, 27'h00000335, 5'd10, 27'h0000031d, 5'd7, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000235, 5'd12, 27'h000003ff, 5'd20, 27'h00000032, 32'h00000400,
  1'd1,  5'd26, 27'h0000032f, 5'd14, 27'h00000261, 5'd26, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003bd, 5'd22, 27'h000001c1, 5'd8, 27'h00000182, 32'h00000400,
  1'd1,  5'd30, 27'h0000032e, 5'd25, 27'h000001c9, 5'd18, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000050, 5'd24, 27'h0000008d, 5'd27, 27'h00000057, 32'h00000400,
  1'd1,  5'd9, 27'h0000011a, 5'd10, 27'h000000f5, 5'd0, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001d3, 5'd5, 27'h000001f7, 5'd10, 27'h000001e2, 32'h00000400,
  1'd1,  5'd5, 27'h000001e8, 5'd5, 27'h0000014b, 5'd21, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000310, 5'd15, 27'h0000036a, 5'd0, 27'h00000022, 32'h00000400,
  1'd1,  5'd7, 27'h000000fc, 5'd19, 27'h000001e2, 5'd13, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001df, 5'd17, 27'h000002e8, 5'd25, 27'h00000295, 32'h00000400,
  1'd1,  5'd10, 27'h0000000d, 5'd29, 27'h000000cc, 5'd3, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000138, 5'd30, 27'h00000117, 5'd12, 27'h000000b9, 32'h00000400,
  1'd1,  5'd7, 27'h00000368, 5'd27, 27'h0000033d, 5'd21, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a2, 5'd8, 27'h00000054, 5'd3, 27'h000002cd, 32'h00000400,
  1'd1,  5'd17, 27'h000001ef, 5'd7, 27'h00000333, 5'd10, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000027b, 5'd5, 27'h00000305, 5'd23, 27'h0000013c, 32'h00000400,
  1'd1,  5'd19, 27'h00000209, 5'd18, 27'h00000105, 5'd4, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000272, 5'd18, 27'h00000326, 5'd13, 27'h00000131, 32'h00000400,
  1'd1,  5'd18, 27'h000000e1, 5'd17, 27'h000002bc, 5'd25, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025c, 5'd26, 27'h000000a1, 5'd1, 27'h0000017a, 32'h00000400,
  1'd1,  5'd16, 27'h0000015f, 5'd27, 27'h000002ce, 5'd13, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a1, 5'd27, 27'h00000341, 5'd25, 27'h0000021a, 32'h00000400,
  1'd1,  5'd29, 27'h000003d6, 5'd9, 27'h00000265, 5'd0, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000007c, 5'd6, 27'h00000068, 5'd14, 27'h000002c3, 32'h00000400,
  1'd1,  5'd29, 27'h00000390, 5'd6, 27'h00000293, 5'd24, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c4, 5'd17, 27'h000002ce, 5'd2, 27'h0000007a, 32'h00000400,
  1'd1,  5'd26, 27'h00000104, 5'd19, 27'h000002b9, 5'd13, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f6, 5'd19, 27'h0000015b, 5'd22, 27'h0000029c, 32'h00000400,
  1'd1,  5'd30, 27'h00000162, 5'd26, 27'h0000016f, 5'd3, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000000a, 5'd30, 27'h00000115, 5'd13, 27'h000002f2, 32'h00000400,
  1'd1,  5'd26, 27'h00000221, 5'd28, 27'h000003eb, 5'd24, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e1, 5'd8, 27'h000001de, 5'd6, 27'h000000de, 32'h00000400,
  1'd1,  5'd10, 27'h00000035, 5'd9, 27'h0000030b, 5'd15, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000025b, 5'd5, 27'h0000027d, 5'd26, 27'h00000389, 32'h00000400,
  1'd1,  5'd9, 27'h0000018e, 5'd17, 27'h000002b8, 5'd9, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003d5, 5'd19, 27'h0000015e, 5'd17, 27'h000002ba, 32'h00000400,
  1'd1,  5'd5, 27'h000003e8, 5'd17, 27'h00000208, 5'd27, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031a, 5'd29, 27'h0000005a, 5'd5, 27'h000003f2, 32'h00000400,
  1'd1,  5'd8, 27'h000001d8, 5'd26, 27'h000002ac, 5'd16, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001dc, 5'd26, 27'h000001bd, 5'd30, 27'h00000086, 32'h00000400,
  1'd1,  5'd20, 27'h000000c7, 5'd5, 27'h000003e9, 5'd6, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000073, 5'd5, 27'h000000bc, 5'd19, 27'h0000005a, 32'h00000400,
  1'd1,  5'd20, 27'h00000033, 5'd6, 27'h000000a6, 5'd25, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d8, 5'd19, 27'h00000386, 5'd8, 27'h00000206, 32'h00000400,
  1'd1,  5'd19, 27'h000002c2, 5'd15, 27'h000003ca, 5'd18, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000193, 5'd18, 27'h00000380, 5'd28, 27'h000000ac, 32'h00000400,
  1'd1,  5'd16, 27'h000000ab, 5'd26, 27'h0000030b, 5'd10, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000b8, 5'd27, 27'h000002cc, 5'd18, 27'h00000145, 32'h00000400,
  1'd1,  5'd19, 27'h00000234, 5'd27, 27'h00000379, 5'd30, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000351, 5'd7, 27'h000003a9, 5'd10, 27'h000000db, 32'h00000400,
  1'd1,  5'd26, 27'h000002f4, 5'd9, 27'h000000ed, 5'd15, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ac, 5'd5, 27'h00000333, 5'd27, 27'h000002fb, 32'h00000400,
  1'd1,  5'd27, 27'h0000008c, 5'd17, 27'h000002b5, 5'd5, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000384, 5'd16, 27'h000002e5, 5'd19, 27'h000003e6, 32'h00000400,
  1'd1,  5'd28, 27'h000001fe, 5'd17, 27'h000002bb, 5'd27, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000131, 5'd29, 27'h00000381, 5'd5, 27'h00000169, 32'h00000400,
  1'd1,  5'd26, 27'h0000028e, 5'd30, 27'h0000008c, 5'd18, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000057, 5'd30, 27'h0000026b, 5'd26, 27'h00000109, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h0000004c, 5'd2, 27'h0000039b, 5'd1, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028a, 5'd4, 27'h0000038e, 5'd13, 27'h00000159, 32'h00000400,
  1'd1,  5'd4, 27'h00000333, 5'd3, 27'h0000006f, 5'd24, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000009b, 5'd11, 27'h00000159, 5'd4, 27'h000000fc, 32'h00000400,
  1'd1,  5'd0, 27'h00000220, 5'd13, 27'h000000e5, 5'd13, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000015, 5'd13, 27'h000001bf, 5'd24, 27'h00000239, 32'h00000400,
  1'd1,  5'd0, 27'h00000259, 5'd21, 27'h000001a8, 5'd4, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000039d, 5'd20, 27'h00000301, 5'd11, 27'h0000033f, 32'h00000400,
  1'd1,  5'd3, 27'h000003b5, 5'd23, 27'h0000026e, 5'd20, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000065, 5'd0, 27'h000000b5, 5'd0, 27'h00000171, 32'h00000400,
  1'd1,  5'd10, 27'h00000239, 5'd3, 27'h00000378, 5'd13, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000017a, 5'd2, 27'h000000fd, 5'd25, 27'h00000079, 32'h00000400,
  1'd1,  5'd12, 27'h0000004b, 5'd10, 27'h0000021d, 5'd3, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000311, 5'd10, 27'h0000019b, 5'd12, 27'h00000359, 32'h00000400,
  1'd1,  5'd14, 27'h00000245, 5'd15, 27'h00000044, 5'd25, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000308, 5'd25, 27'h0000027d, 5'd2, 27'h0000032a, 32'h00000400,
  1'd1,  5'd11, 27'h00000260, 5'd22, 27'h00000207, 5'd12, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000263, 5'd23, 27'h00000128, 5'd25, 27'h000001f9, 32'h00000400,
  1'd1,  5'd21, 27'h00000311, 5'd2, 27'h0000036a, 5'd3, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000321, 5'd2, 27'h000002c4, 5'd13, 27'h0000012a, 32'h00000400,
  1'd1,  5'd25, 27'h000002e5, 5'd4, 27'h000001c5, 5'd23, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d2, 5'd10, 27'h00000356, 5'd0, 27'h00000210, 32'h00000400,
  1'd1,  5'd25, 27'h000002a2, 5'd12, 27'h0000036e, 5'd14, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c9, 5'd11, 27'h00000054, 5'd25, 27'h00000283, 32'h00000400,
  1'd1,  5'd24, 27'h00000131, 5'd24, 27'h00000253, 5'd1, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000017a, 5'd24, 27'h0000032e, 5'd12, 27'h00000323, 32'h00000400,
  1'd1,  5'd21, 27'h0000011b, 5'd23, 27'h0000011c, 5'd21, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000178, 5'd0, 27'h00000196, 5'd7, 27'h0000009b, 32'h00000400,
  1'd1,  5'd1, 27'h00000139, 5'd4, 27'h000003bc, 5'd18, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000016, 5'd1, 27'h0000032b, 5'd27, 27'h0000035d, 32'h00000400,
  1'd1,  5'd0, 27'h000002e0, 5'd10, 27'h000001ef, 5'd6, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003bf, 5'd11, 27'h000001ef, 5'd19, 27'h0000018e, 32'h00000400,
  1'd1,  5'd2, 27'h0000036b, 5'd11, 27'h00000049, 5'd26, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000373, 5'd23, 27'h00000091, 5'd8, 27'h0000008c, 32'h00000400,
  1'd1,  5'd3, 27'h00000267, 5'd21, 27'h0000012a, 5'd20, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c6, 5'd21, 27'h0000022f, 5'd29, 27'h00000278, 32'h00000400,
  1'd1,  5'd15, 27'h000001f6, 5'd3, 27'h0000038d, 5'd9, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003c2, 5'd2, 27'h000001f2, 5'd17, 27'h00000092, 32'h00000400,
  1'd1,  5'd11, 27'h000001f4, 5'd2, 27'h00000380, 5'd30, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f1, 5'd11, 27'h00000209, 5'd5, 27'h00000389, 32'h00000400,
  1'd1,  5'd12, 27'h00000232, 5'd12, 27'h00000253, 5'd20, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000036b, 5'd13, 27'h00000035, 5'd29, 27'h00000316, 32'h00000400,
  1'd1,  5'd10, 27'h0000020f, 5'd22, 27'h00000272, 5'd8, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000aa, 5'd22, 27'h000000c1, 5'd16, 27'h00000077, 32'h00000400,
  1'd1,  5'd12, 27'h000000c6, 5'd22, 27'h000002be, 5'd28, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000185, 5'd1, 27'h00000378, 5'd8, 27'h00000044, 32'h00000400,
  1'd1,  5'd21, 27'h0000022a, 5'd2, 27'h000003d4, 5'd20, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002e9, 5'd1, 27'h000002d0, 5'd26, 27'h00000096, 32'h00000400,
  1'd1,  5'd24, 27'h000001d6, 5'd12, 27'h00000220, 5'd9, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000036, 5'd14, 27'h00000280, 5'd18, 27'h000002d5, 32'h00000400,
  1'd1,  5'd25, 27'h0000022a, 5'd14, 27'h00000242, 5'd28, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000235, 5'd23, 27'h000003b6, 5'd6, 27'h000002a0, 32'h00000400,
  1'd1,  5'd22, 27'h000000f0, 5'd22, 27'h000000e8, 5'd20, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003ab, 5'd25, 27'h00000306, 5'd30, 27'h000002f8, 32'h00000400,
  1'd1,  5'd0, 27'h00000013, 5'd9, 27'h0000039a, 5'd3, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003db, 5'd8, 27'h000001c9, 5'd13, 27'h00000135, 32'h00000400,
  1'd1,  5'd0, 27'h000003b7, 5'd7, 27'h00000087, 5'd24, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002df, 5'd18, 27'h00000075, 5'd0, 27'h000002d8, 32'h00000400,
  1'd1,  5'd0, 27'h0000014e, 5'd18, 27'h00000153, 5'd14, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000188, 5'd16, 27'h0000003f, 5'd22, 27'h0000012f, 32'h00000400,
  1'd1,  5'd3, 27'h000002a5, 5'd29, 27'h00000043, 5'd1, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000066, 5'd28, 27'h000003dc, 5'd12, 27'h0000030b, 32'h00000400,
  1'd1,  5'd1, 27'h00000234, 5'd29, 27'h00000275, 5'd20, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000268, 5'd6, 27'h0000009e, 5'd0, 27'h00000219, 32'h00000400,
  1'd1,  5'd11, 27'h00000272, 5'd9, 27'h00000029, 5'd11, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000f9, 5'd5, 27'h00000206, 5'd23, 27'h00000335, 32'h00000400,
  1'd1,  5'd12, 27'h0000022d, 5'd17, 27'h0000033b, 5'd0, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c8, 5'd16, 27'h00000327, 5'd10, 27'h00000232, 32'h00000400,
  1'd1,  5'd12, 27'h0000029f, 5'd17, 27'h0000001d, 5'd21, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000024f, 5'd29, 27'h0000025f, 5'd1, 27'h000000a0, 32'h00000400,
  1'd1,  5'd15, 27'h000001a1, 5'd29, 27'h000003c4, 5'd10, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000157, 5'd25, 27'h00000370, 5'd21, 27'h000002db, 32'h00000400,
  1'd1,  5'd21, 27'h0000007f, 5'd6, 27'h00000166, 5'd1, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000072, 5'd9, 27'h00000242, 5'd14, 27'h0000006f, 32'h00000400,
  1'd1,  5'd25, 27'h00000305, 5'd8, 27'h00000178, 5'd24, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003e4, 5'd19, 27'h000000df, 5'd4, 27'h0000011c, 32'h00000400,
  1'd1,  5'd21, 27'h000002ba, 5'd17, 27'h0000014d, 5'd14, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000342, 5'd16, 27'h00000083, 5'd25, 27'h000001de, 32'h00000400,
  1'd1,  5'd22, 27'h000001a8, 5'd28, 27'h00000177, 5'd3, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000328, 5'd27, 27'h000002e5, 5'd12, 27'h0000015a, 32'h00000400,
  1'd1,  5'd22, 27'h0000020d, 5'd26, 27'h000003e2, 5'd24, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000006, 5'd6, 27'h00000135, 5'd9, 27'h00000350, 32'h00000400,
  1'd1,  5'd4, 27'h00000161, 5'd6, 27'h00000361, 5'd19, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000009e, 5'd7, 27'h0000028d, 5'd30, 27'h0000020e, 32'h00000400,
  1'd1,  5'd0, 27'h000000bf, 5'd18, 27'h00000206, 5'd5, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000253, 5'd17, 27'h00000046, 5'd15, 27'h000002fd, 32'h00000400,
  1'd1,  5'd3, 27'h000000b8, 5'd16, 27'h000003cf, 5'd30, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000030d, 5'd26, 27'h0000029e, 5'd9, 27'h00000022, 32'h00000400,
  1'd1,  5'd1, 27'h00000107, 5'd26, 27'h00000034, 5'd18, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036a, 5'd28, 27'h0000010c, 5'd26, 27'h00000112, 32'h00000400,
  1'd1,  5'd14, 27'h000003d6, 5'd6, 27'h000000d7, 5'd5, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000034f, 5'd7, 27'h0000036a, 5'd20, 27'h0000028e, 32'h00000400,
  1'd1,  5'd12, 27'h000001a5, 5'd5, 27'h00000376, 5'd27, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000034a, 5'd19, 27'h0000020c, 5'd10, 27'h000000d7, 32'h00000400,
  1'd1,  5'd11, 27'h000000b3, 5'd20, 27'h000000d2, 5'd18, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000332, 5'd18, 27'h00000350, 5'd28, 27'h00000336, 32'h00000400,
  1'd1,  5'd15, 27'h000000be, 5'd28, 27'h00000352, 5'd9, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000279, 5'd26, 27'h00000283, 5'd19, 27'h0000014d, 32'h00000400,
  1'd1,  5'd15, 27'h0000005e, 5'd30, 27'h000001b0, 5'd26, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000026d, 5'd7, 27'h00000038, 5'd6, 27'h00000282, 32'h00000400,
  1'd1,  5'd25, 27'h0000028d, 5'd6, 27'h00000209, 5'd17, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000161, 5'd9, 27'h00000270, 5'd27, 27'h0000020f, 32'h00000400,
  1'd1,  5'd24, 27'h000000b2, 5'd19, 27'h00000119, 5'd7, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000013d, 5'd19, 27'h000002f7, 5'd17, 27'h00000200, 32'h00000400,
  1'd1,  5'd25, 27'h000001a4, 5'd17, 27'h00000070, 5'd28, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000003c, 5'd29, 27'h00000006, 5'd5, 27'h00000282, 32'h00000400,
  1'd1,  5'd23, 27'h00000280, 5'd27, 27'h000000b8, 5'd20, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000301, 5'd30, 27'h00000242, 5'd29, 27'h000002c3, 32'h00000400,
  1'd1,  5'd9, 27'h000002cb, 5'd0, 27'h00000095, 5'd8, 27'h0000017f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002f8, 5'd2, 27'h00000329, 5'd20, 27'h00000019, 32'h00000400,
  1'd1,  5'd8, 27'h000002dc, 5'd0, 27'h00000191, 5'd29, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000262, 5'd11, 27'h0000036f, 5'd3, 27'h00000264, 32'h00000400,
  1'd1,  5'd6, 27'h00000393, 5'd14, 27'h00000194, 5'd12, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000a1, 5'd11, 27'h000000d4, 5'd23, 27'h0000032e, 32'h00000400,
  1'd1,  5'd8, 27'h00000133, 5'd21, 27'h000003b7, 5'd4, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002fa, 5'd22, 27'h0000039b, 5'd14, 27'h0000023e, 32'h00000400,
  1'd1,  5'd8, 27'h00000259, 5'd21, 27'h0000006d, 5'd24, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000055, 5'd3, 27'h000003b3, 5'd7, 27'h000000e1, 32'h00000400,
  1'd1,  5'd18, 27'h000003de, 5'd3, 27'h000002cb, 5'd18, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f8, 5'd3, 27'h00000090, 5'd26, 27'h00000217, 32'h00000400,
  1'd1,  5'd18, 27'h000001a0, 5'd13, 27'h000001e0, 5'd2, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002fb, 5'd12, 27'h00000155, 5'd11, 27'h0000015e, 32'h00000400,
  1'd1,  5'd19, 27'h00000091, 5'd15, 27'h000001b8, 5'd25, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ca, 5'd22, 27'h000000e6, 5'd3, 27'h00000283, 32'h00000400,
  1'd1,  5'd19, 27'h00000375, 5'd25, 27'h0000007e, 5'd14, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000002f, 5'd20, 27'h00000391, 5'd20, 27'h000003c5, 32'h00000400,
  1'd1,  5'd28, 27'h000001c0, 5'd2, 27'h0000037d, 5'd4, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000362, 5'd2, 27'h00000205, 5'd15, 27'h0000005e, 32'h00000400,
  1'd1,  5'd26, 27'h00000380, 5'd4, 27'h0000020b, 5'd25, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000f7, 5'd14, 27'h000002e7, 5'd3, 27'h0000017e, 32'h00000400,
  1'd1,  5'd30, 27'h00000278, 5'd12, 27'h000000b2, 5'd12, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c1, 5'd15, 27'h00000017, 5'd25, 27'h0000025a, 32'h00000400,
  1'd1,  5'd27, 27'h00000028, 5'd21, 27'h00000095, 5'd2, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003d4, 5'd20, 27'h000002de, 5'd13, 27'h000002a5, 32'h00000400,
  1'd1,  5'd28, 27'h0000038d, 5'd22, 27'h000002e7, 5'd25, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000207, 5'd0, 27'h0000002b, 5'd2, 27'h0000002e, 32'h00000400,
  1'd1,  5'd7, 27'h0000002c, 5'd5, 27'h00000044, 5'd14, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001a7, 5'd1, 27'h000002a5, 5'd24, 27'h0000022b, 32'h00000400,
  1'd1,  5'd8, 27'h0000028c, 5'd12, 27'h00000313, 5'd7, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000190, 5'd15, 27'h000000b8, 5'd16, 27'h000002a6, 32'h00000400,
  1'd1,  5'd5, 27'h000002e8, 5'd12, 27'h000003fb, 5'd30, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000280, 5'd21, 27'h0000014d, 5'd5, 27'h000003b1, 32'h00000400,
  1'd1,  5'd7, 27'h00000059, 5'd23, 27'h000003e5, 5'd17, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000067, 5'd23, 27'h0000009e, 5'd26, 27'h000003fe, 32'h00000400,
  1'd1,  5'd18, 27'h00000219, 5'd2, 27'h0000039f, 5'd3, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003e5, 5'd0, 27'h0000025b, 5'd14, 27'h00000241, 32'h00000400,
  1'd1,  5'd16, 27'h00000028, 5'd1, 27'h000001bd, 5'd23, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000337, 5'd12, 27'h00000112, 5'd8, 27'h000002fc, 32'h00000400,
  1'd1,  5'd20, 27'h00000220, 5'd13, 27'h0000030f, 5'd19, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000dc, 5'd11, 27'h00000152, 5'd30, 27'h00000187, 32'h00000400,
  1'd1,  5'd17, 27'h000002fd, 5'd22, 27'h000000f3, 5'd9, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000079, 5'd23, 27'h0000022f, 5'd18, 27'h00000391, 32'h00000400,
  1'd1,  5'd16, 27'h00000200, 5'd21, 27'h000002da, 5'd28, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000252, 5'd4, 27'h000002bd, 5'd7, 27'h00000034, 32'h00000400,
  1'd1,  5'd30, 27'h00000064, 5'd3, 27'h000001c3, 5'd19, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000041, 5'd2, 27'h0000026c, 5'd26, 27'h0000004a, 32'h00000400,
  1'd1,  5'd29, 27'h00000262, 5'd13, 27'h00000089, 5'd5, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000348, 5'd11, 27'h0000022a, 5'd17, 27'h00000196, 32'h00000400,
  1'd1,  5'd28, 27'h000000fd, 5'd13, 27'h00000194, 5'd29, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000171, 5'd23, 27'h00000162, 5'd6, 27'h00000287, 32'h00000400,
  1'd1,  5'd27, 27'h0000010a, 5'd24, 27'h0000034d, 5'd19, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000144, 5'd24, 27'h00000170, 5'd28, 27'h00000037, 32'h00000400,
  1'd1,  5'd8, 27'h000000de, 5'd8, 27'h0000006d, 5'd2, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000014d, 5'd8, 27'h00000031, 5'd15, 27'h000000c2, 32'h00000400,
  1'd1,  5'd6, 27'h0000002c, 5'd8, 27'h000002e3, 5'd21, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fd, 5'd15, 27'h00000282, 5'd1, 27'h000003f4, 32'h00000400,
  1'd1,  5'd9, 27'h00000179, 5'd20, 27'h000001a0, 5'd15, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000176, 5'd16, 27'h000000ef, 5'd22, 27'h00000174, 32'h00000400,
  1'd1,  5'd5, 27'h00000389, 5'd30, 27'h000003cd, 5'd1, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001a6, 5'd26, 27'h00000046, 5'd10, 27'h00000165, 32'h00000400,
  1'd1,  5'd9, 27'h0000000f, 5'd26, 27'h00000249, 5'd22, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002fc, 5'd6, 27'h0000004b, 5'd0, 27'h000003e0, 32'h00000400,
  1'd1,  5'd19, 27'h00000344, 5'd9, 27'h00000112, 5'd13, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d5, 5'd10, 27'h0000006d, 5'd22, 27'h000003af, 32'h00000400,
  1'd1,  5'd19, 27'h000003e6, 5'd18, 27'h000003ec, 5'd3, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000027, 5'd15, 27'h000002a6, 5'd12, 27'h000001bc, 32'h00000400,
  1'd1,  5'd20, 27'h0000002a, 5'd20, 27'h00000018, 5'd24, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003b9, 5'd29, 27'h000001de, 5'd4, 27'h000002f6, 32'h00000400,
  1'd1,  5'd15, 27'h0000024b, 5'd26, 27'h000000f9, 5'd12, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003aa, 5'd30, 27'h00000163, 5'd23, 27'h0000018d, 32'h00000400,
  1'd1,  5'd25, 27'h000003a7, 5'd7, 27'h00000080, 5'd4, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000036f, 5'd8, 27'h000001ca, 5'd14, 27'h0000031a, 32'h00000400,
  1'd1,  5'd27, 27'h00000271, 5'd5, 27'h0000034f, 5'd22, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001df, 5'd17, 27'h00000123, 5'd2, 27'h000002ae, 32'h00000400,
  1'd1,  5'd27, 27'h0000035d, 5'd16, 27'h0000023b, 5'd15, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000378, 5'd16, 27'h00000339, 5'd22, 27'h000001dd, 32'h00000400,
  1'd1,  5'd25, 27'h000003ba, 5'd26, 27'h0000034b, 5'd2, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b7, 5'd27, 27'h00000378, 5'd11, 27'h000003e2, 32'h00000400,
  1'd1,  5'd28, 27'h0000003f, 5'd29, 27'h000003fc, 5'd23, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000173, 5'd8, 27'h000000c2, 5'd8, 27'h00000139, 32'h00000400,
  1'd1,  5'd7, 27'h000001c4, 5'd5, 27'h000000bc, 5'd20, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000379, 5'd8, 27'h000000ad, 5'd28, 27'h000003f8, 32'h00000400,
  1'd1,  5'd7, 27'h0000018c, 5'd19, 27'h00000182, 5'd8, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003c, 5'd16, 27'h00000024, 5'd17, 27'h0000016e, 32'h00000400,
  1'd1,  5'd6, 27'h000003d7, 5'd19, 27'h00000119, 5'd28, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000012e, 5'd27, 27'h000000fe, 5'd9, 27'h000002cf, 32'h00000400,
  1'd1,  5'd10, 27'h0000006b, 5'd26, 27'h00000121, 5'd17, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000002f, 5'd27, 27'h000001e2, 5'd27, 27'h0000032f, 32'h00000400,
  1'd1,  5'd16, 27'h000001cd, 5'd6, 27'h000001fa, 5'd5, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b7, 5'd8, 27'h00000293, 5'd19, 27'h00000183, 32'h00000400,
  1'd1,  5'd16, 27'h00000210, 5'd7, 27'h00000211, 5'd29, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000105, 5'd16, 27'h0000030f, 5'd9, 27'h0000011b, 32'h00000400,
  1'd1,  5'd18, 27'h000001e9, 5'd18, 27'h00000384, 5'd18, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003d0, 5'd18, 27'h0000005d, 5'd27, 27'h00000294, 32'h00000400,
  1'd1,  5'd19, 27'h000003c7, 5'd30, 27'h0000004d, 5'd6, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e5, 5'd27, 27'h000000cf, 5'd16, 27'h000001fc, 32'h00000400,
  1'd1,  5'd15, 27'h000003ad, 5'd30, 27'h000003cd, 5'd29, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e5, 5'd9, 27'h00000055, 5'd9, 27'h00000232, 32'h00000400,
  1'd1,  5'd29, 27'h000003c1, 5'd9, 27'h000000f3, 5'd18, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000029d, 5'd6, 27'h000003e3, 5'd30, 27'h0000036a, 32'h00000400,
  1'd1,  5'd28, 27'h000000bd, 5'd18, 27'h000001db, 5'd9, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000033d, 5'd19, 27'h000000f9, 5'd17, 27'h00000043, 32'h00000400,
  1'd1,  5'd30, 27'h00000309, 5'd17, 27'h00000394, 5'd29, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000025d, 5'd28, 27'h00000062, 5'd5, 27'h000003a9, 32'h00000400,
  1'd1,  5'd25, 27'h00000374, 5'd26, 27'h00000388, 5'd18, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000025a, 5'd28, 27'h00000394, 5'd25, 27'h000003fd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000271, 5'd2, 27'h000000e8, 5'd1, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000035e, 5'd2, 27'h000003c7, 5'd13, 27'h000001f5, 32'h00000400,
  1'd1,  5'd2, 27'h0000012c, 5'd2, 27'h0000015b, 5'd23, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000c2, 5'd13, 27'h0000039b, 5'd2, 27'h000000c4, 32'h00000400,
  1'd1,  5'd0, 27'h000003f1, 5'd11, 27'h000002a7, 5'd14, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000321, 5'd11, 27'h00000304, 5'd22, 27'h000000db, 32'h00000400,
  1'd1,  5'd4, 27'h0000032e, 5'd24, 27'h00000127, 5'd0, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000009e, 5'd22, 27'h000003f3, 5'd10, 27'h0000033f, 32'h00000400,
  1'd1,  5'd1, 27'h0000003e, 5'd23, 27'h000000c6, 5'd24, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003c1, 5'd1, 27'h0000007e, 5'd0, 27'h0000017a, 32'h00000400,
  1'd1,  5'd13, 27'h000002e6, 5'd1, 27'h00000329, 5'd15, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000281, 5'd2, 27'h00000353, 5'd23, 27'h000002ef, 32'h00000400,
  1'd1,  5'd13, 27'h000000ed, 5'd13, 27'h000002b2, 5'd5, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021d, 5'd12, 27'h0000027c, 5'd15, 27'h00000003, 32'h00000400,
  1'd1,  5'd11, 27'h0000028e, 5'd10, 27'h0000039d, 5'd22, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001c9, 5'd24, 27'h000003a2, 5'd1, 27'h0000008e, 32'h00000400,
  1'd1,  5'd15, 27'h000001d0, 5'd23, 27'h00000039, 5'd14, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000032, 5'd23, 27'h00000319, 5'd21, 27'h00000331, 32'h00000400,
  1'd1,  5'd22, 27'h00000258, 5'd4, 27'h000003ab, 5'd0, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d8, 5'd4, 27'h00000376, 5'd12, 27'h000000cf, 32'h00000400,
  1'd1,  5'd22, 27'h000003ae, 5'd3, 27'h00000009, 5'd21, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000385, 5'd10, 27'h00000180, 5'd1, 27'h0000018f, 32'h00000400,
  1'd1,  5'd21, 27'h000002af, 5'd12, 27'h000002bc, 5'd14, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000bb, 5'd12, 27'h000002f8, 5'd22, 27'h00000179, 32'h00000400,
  1'd1,  5'd24, 27'h00000020, 5'd21, 27'h00000282, 5'd1, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000076, 5'd25, 27'h00000056, 5'd11, 27'h000003e7, 32'h00000400,
  1'd1,  5'd22, 27'h00000034, 5'd25, 27'h00000110, 5'd20, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000035b, 5'd1, 27'h00000136, 5'd6, 27'h0000023f, 32'h00000400,
  1'd1,  5'd3, 27'h000002ec, 5'd0, 27'h00000283, 5'd16, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ab, 5'd4, 27'h00000126, 5'd28, 27'h00000300, 32'h00000400,
  1'd1,  5'd2, 27'h000001f6, 5'd10, 27'h00000287, 5'd5, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000037a, 5'd11, 27'h000002b2, 5'd17, 27'h000001d6, 32'h00000400,
  1'd1,  5'd4, 27'h000003c6, 5'd13, 27'h0000027e, 5'd28, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000023, 5'd25, 27'h00000313, 5'd9, 27'h00000280, 32'h00000400,
  1'd1,  5'd0, 27'h0000033f, 5'd22, 27'h000001f0, 5'd19, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000028e, 5'd22, 27'h0000027f, 5'd30, 27'h00000102, 32'h00000400,
  1'd1,  5'd11, 27'h0000035c, 5'd1, 27'h00000072, 5'd8, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000033b, 5'd1, 27'h000000b5, 5'd15, 27'h000003d1, 32'h00000400,
  1'd1,  5'd12, 27'h000001ba, 5'd4, 27'h000001f5, 5'd29, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000061, 5'd13, 27'h00000364, 5'd6, 27'h0000034e, 32'h00000400,
  1'd1,  5'd14, 27'h000003fb, 5'd14, 27'h000003a4, 5'd19, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000115, 5'd11, 27'h0000006e, 5'd28, 27'h0000014c, 32'h00000400,
  1'd1,  5'd14, 27'h00000112, 5'd25, 27'h000000c0, 5'd7, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001f3, 5'd21, 27'h000002f5, 5'd16, 27'h0000024c, 32'h00000400,
  1'd1,  5'd12, 27'h00000085, 5'd25, 27'h000002fc, 5'd26, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003dd, 5'd0, 27'h000002e1, 5'd10, 27'h00000088, 32'h00000400,
  1'd1,  5'd22, 27'h00000368, 5'd1, 27'h00000288, 5'd19, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000112, 5'd4, 27'h0000039a, 5'd27, 27'h00000058, 32'h00000400,
  1'd1,  5'd22, 27'h000002cd, 5'd12, 27'h00000366, 5'd9, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000008f, 5'd13, 27'h00000302, 5'd18, 27'h000002a3, 32'h00000400,
  1'd1,  5'd23, 27'h000002be, 5'd15, 27'h00000055, 5'd27, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000350, 5'd23, 27'h000003ee, 5'd8, 27'h0000009e, 32'h00000400,
  1'd1,  5'd24, 27'h0000028f, 5'd21, 27'h00000149, 5'd18, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000027b, 5'd22, 27'h000001c6, 5'd26, 27'h0000000a, 32'h00000400,
  1'd1,  5'd3, 27'h00000061, 5'd8, 27'h00000137, 5'd2, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000003e, 5'd9, 27'h000002ee, 5'd14, 27'h000002e5, 32'h00000400,
  1'd1,  5'd1, 27'h00000028, 5'd8, 27'h0000024e, 5'd24, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000006b, 5'd16, 27'h0000036b, 5'd3, 27'h000003b7, 32'h00000400,
  1'd1,  5'd2, 27'h00000170, 5'd19, 27'h000001d9, 5'd12, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002b9, 5'd15, 27'h0000034b, 5'd24, 27'h00000263, 32'h00000400,
  1'd1,  5'd2, 27'h000002d4, 5'd27, 27'h0000002a, 5'd3, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000006c, 5'd28, 27'h0000022d, 5'd15, 27'h00000138, 32'h00000400,
  1'd1,  5'd4, 27'h000001e5, 5'd26, 27'h00000222, 5'd25, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003b9, 5'd10, 27'h00000086, 5'd4, 27'h00000187, 32'h00000400,
  1'd1,  5'd14, 27'h00000074, 5'd7, 27'h00000101, 5'd12, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003bf, 5'd10, 27'h00000013, 5'd21, 27'h00000047, 32'h00000400,
  1'd1,  5'd15, 27'h000001ce, 5'd16, 27'h000000f3, 5'd4, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000101, 5'd17, 27'h00000020, 5'd12, 27'h000000d9, 32'h00000400,
  1'd1,  5'd10, 27'h0000017f, 5'd18, 27'h00000388, 5'd23, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000013e, 5'd29, 27'h0000014b, 5'd3, 27'h00000095, 32'h00000400,
  1'd1,  5'd13, 27'h00000371, 5'd28, 27'h0000035b, 5'd14, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002bc, 5'd30, 27'h0000021b, 5'd23, 27'h0000037f, 32'h00000400,
  1'd1,  5'd20, 27'h000003b1, 5'd6, 27'h00000234, 5'd5, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d6, 5'd8, 27'h0000025a, 5'd13, 27'h00000135, 32'h00000400,
  1'd1,  5'd21, 27'h00000244, 5'd8, 27'h0000008b, 5'd25, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001bc, 5'd18, 27'h0000037f, 5'd4, 27'h0000006b, 32'h00000400,
  1'd1,  5'd20, 27'h00000391, 5'd18, 27'h000002e1, 5'd11, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000008, 5'd15, 27'h00000277, 5'd22, 27'h000001a8, 32'h00000400,
  1'd1,  5'd23, 27'h000002c4, 5'd25, 27'h00000372, 5'd3, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000033e, 5'd26, 27'h000001d0, 5'd13, 27'h000000eb, 32'h00000400,
  1'd1,  5'd25, 27'h000002f5, 5'd27, 27'h0000013f, 5'd24, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001dd, 5'd7, 27'h000002be, 5'd9, 27'h00000250, 32'h00000400,
  1'd1,  5'd0, 27'h000002ae, 5'd9, 27'h00000034, 5'd17, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000242, 5'd9, 27'h0000036e, 5'd26, 27'h00000143, 32'h00000400,
  1'd1,  5'd4, 27'h000001d8, 5'd18, 27'h00000314, 5'd9, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000099, 5'd17, 27'h00000191, 5'd18, 27'h000000b1, 32'h00000400,
  1'd1,  5'd3, 27'h0000014b, 5'd15, 27'h00000284, 5'd27, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005a, 5'd26, 27'h00000088, 5'd10, 27'h0000006f, 32'h00000400,
  1'd1,  5'd2, 27'h0000013f, 5'd30, 27'h0000029f, 5'd18, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000022, 5'd26, 27'h00000359, 5'd28, 27'h000003a9, 32'h00000400,
  1'd1,  5'd14, 27'h00000031, 5'd6, 27'h000003a5, 5'd7, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002bd, 5'd7, 27'h00000137, 5'd16, 27'h0000029e, 32'h00000400,
  1'd1,  5'd11, 27'h0000014d, 5'd8, 27'h00000213, 5'd28, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002a7, 5'd20, 27'h00000296, 5'd6, 27'h00000292, 32'h00000400,
  1'd1,  5'd11, 27'h000002e4, 5'd17, 27'h00000343, 5'd17, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000039a, 5'd17, 27'h00000290, 5'd26, 27'h000001d8, 32'h00000400,
  1'd1,  5'd11, 27'h000001d2, 5'd26, 27'h00000377, 5'd6, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f9, 5'd28, 27'h000002e0, 5'd16, 27'h00000083, 32'h00000400,
  1'd1,  5'd14, 27'h00000039, 5'd29, 27'h000000d0, 5'd28, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000319, 5'd5, 27'h000000eb, 5'd6, 27'h00000340, 32'h00000400,
  1'd1,  5'd20, 27'h000003e1, 5'd6, 27'h000002c4, 5'd18, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000032b, 5'd8, 27'h00000300, 5'd27, 27'h0000039c, 32'h00000400,
  1'd1,  5'd22, 27'h000000c4, 5'd17, 27'h000002e3, 5'd7, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000035a, 5'd18, 27'h00000073, 5'd19, 27'h000003fd, 32'h00000400,
  1'd1,  5'd25, 27'h00000317, 5'd20, 27'h000001da, 5'd27, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000363, 5'd28, 27'h00000231, 5'd10, 27'h00000002, 32'h00000400,
  1'd1,  5'd21, 27'h0000037a, 5'd28, 27'h000002e6, 5'd16, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bb, 5'd27, 27'h0000010e, 5'd26, 27'h00000200, 32'h00000400,
  1'd1,  5'd8, 27'h00000191, 5'd2, 27'h0000031c, 5'd10, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000070, 5'd1, 27'h000000c1, 5'd18, 27'h000002dc, 32'h00000400,
  1'd1,  5'd7, 27'h00000359, 5'd3, 27'h000003ed, 5'd26, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000020d, 5'd13, 27'h00000288, 5'd0, 27'h000002e3, 32'h00000400,
  1'd1,  5'd6, 27'h000000ae, 5'd14, 27'h000000ee, 5'd12, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001a8, 5'd12, 27'h00000041, 5'd25, 27'h0000011a, 32'h00000400,
  1'd1,  5'd8, 27'h00000328, 5'd25, 27'h00000216, 5'd0, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002df, 5'd23, 27'h000002cf, 5'd11, 27'h00000164, 32'h00000400,
  1'd1,  5'd5, 27'h000002c1, 5'd21, 27'h000003ce, 5'd21, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e7, 5'd4, 27'h00000353, 5'd8, 27'h000002d6, 32'h00000400,
  1'd1,  5'd19, 27'h0000019b, 5'd0, 27'h00000341, 5'd16, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ef, 5'd2, 27'h00000283, 5'd27, 27'h00000348, 32'h00000400,
  1'd1,  5'd19, 27'h0000029d, 5'd15, 27'h00000072, 5'd1, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000025, 5'd15, 27'h00000082, 5'd15, 27'h000000ee, 32'h00000400,
  1'd1,  5'd19, 27'h000001bd, 5'd15, 27'h00000144, 5'd24, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000223, 5'd23, 27'h000003fd, 5'd4, 27'h000001f8, 32'h00000400,
  1'd1,  5'd19, 27'h000001b6, 5'd23, 27'h000000ed, 5'd14, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002a5, 5'd23, 27'h00000303, 5'd21, 27'h00000365, 32'h00000400,
  1'd1,  5'd26, 27'h000002ec, 5'd4, 27'h00000368, 5'd4, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b9, 5'd1, 27'h000002a9, 5'd15, 27'h000001a6, 32'h00000400,
  1'd1,  5'd30, 27'h00000241, 5'd3, 27'h00000086, 5'd25, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000231, 5'd13, 27'h000002c3, 5'd1, 27'h00000294, 32'h00000400,
  1'd1,  5'd28, 27'h000001f9, 5'd14, 27'h000001b0, 5'd13, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000071, 5'd11, 27'h0000014a, 5'd22, 27'h00000351, 32'h00000400,
  1'd1,  5'd26, 27'h000002d8, 5'd24, 27'h00000232, 5'd1, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000034e, 5'd24, 27'h000000e3, 5'd10, 27'h000002b3, 32'h00000400,
  1'd1,  5'd28, 27'h000003d7, 5'd22, 27'h000002a9, 5'd21, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000002e, 5'd0, 27'h00000205, 5'd0, 27'h00000002, 32'h00000400,
  1'd1,  5'd8, 27'h00000136, 5'd0, 27'h000001c1, 5'd14, 27'h0000002c, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000017c, 5'd5, 27'h00000094, 5'd21, 27'h0000013a, 32'h00000400,
  1'd1,  5'd7, 27'h0000014b, 5'd11, 27'h0000035c, 5'd9, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000002e, 5'd13, 27'h0000029f, 5'd19, 27'h00000393, 32'h00000400,
  1'd1,  5'd8, 27'h000000c8, 5'd14, 27'h0000023b, 5'd28, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ef, 5'd21, 27'h00000333, 5'd5, 27'h0000024c, 32'h00000400,
  1'd1,  5'd8, 27'h00000292, 5'd21, 27'h0000008b, 5'd15, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000244, 5'd24, 27'h00000297, 5'd28, 27'h00000362, 32'h00000400,
  1'd1,  5'd18, 27'h0000009b, 5'd0, 27'h00000157, 5'd2, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000299, 5'd1, 27'h00000236, 5'd11, 27'h0000012a, 32'h00000400,
  1'd1,  5'd16, 27'h00000104, 5'd2, 27'h000003e0, 5'd22, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000025d, 5'd15, 27'h000000fd, 5'd6, 27'h0000012e, 32'h00000400,
  1'd1,  5'd16, 27'h000001a1, 5'd13, 27'h000001b4, 5'd16, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000174, 5'd13, 27'h000003ef, 5'd28, 27'h0000001a, 32'h00000400,
  1'd1,  5'd17, 27'h0000012d, 5'd25, 27'h00000325, 5'd6, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003dc, 5'd25, 27'h0000030b, 5'd20, 27'h00000274, 32'h00000400,
  1'd1,  5'd17, 27'h000000d4, 5'd22, 27'h000001d5, 5'd27, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000038a, 5'd2, 27'h000001a9, 5'd8, 27'h000000bd, 32'h00000400,
  1'd1,  5'd29, 27'h000002e7, 5'd2, 27'h00000341, 5'd15, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f2, 5'd3, 27'h0000014b, 5'd26, 27'h000003eb, 32'h00000400,
  1'd1,  5'd28, 27'h000003c4, 5'd12, 27'h00000021, 5'd8, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000169, 5'd11, 27'h00000221, 5'd16, 27'h00000398, 32'h00000400,
  1'd1,  5'd28, 27'h0000036d, 5'd13, 27'h00000314, 5'd26, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000061, 5'd23, 27'h000001e1, 5'd7, 27'h00000251, 32'h00000400,
  1'd1,  5'd28, 27'h000000b1, 5'd22, 27'h000001a1, 5'd18, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000012, 5'd22, 27'h000002e0, 5'd28, 27'h0000017e, 32'h00000400,
  1'd1,  5'd6, 27'h0000016b, 5'd9, 27'h000003af, 5'd4, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000bc, 5'd7, 27'h000002fb, 5'd11, 27'h00000314, 32'h00000400,
  1'd1,  5'd7, 27'h00000187, 5'd8, 27'h00000099, 5'd22, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000171, 5'd16, 27'h000001d8, 5'd4, 27'h00000023, 32'h00000400,
  1'd1,  5'd5, 27'h00000251, 5'd18, 27'h000003c8, 5'd13, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000012b, 5'd19, 27'h00000029, 5'd25, 27'h0000019b, 32'h00000400,
  1'd1,  5'd7, 27'h00000103, 5'd30, 27'h000000fa, 5'd2, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000366, 5'd26, 27'h0000013c, 5'd10, 27'h00000228, 32'h00000400,
  1'd1,  5'd9, 27'h00000074, 5'd26, 27'h000001f4, 5'd22, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002f5, 5'd5, 27'h000002ca, 5'd3, 27'h000001bb, 32'h00000400,
  1'd1,  5'd19, 27'h0000035c, 5'd6, 27'h000001ab, 5'd13, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003dd, 5'd9, 27'h000000bd, 5'd25, 27'h00000308, 32'h00000400,
  1'd1,  5'd16, 27'h00000056, 5'd16, 27'h00000018, 5'd4, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003cd, 5'd16, 27'h000001d3, 5'd14, 27'h000001d5, 32'h00000400,
  1'd1,  5'd19, 27'h0000010c, 5'd20, 27'h000002a7, 5'd23, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000017d, 5'd29, 27'h00000097, 5'd2, 27'h000000f8, 32'h00000400,
  1'd1,  5'd19, 27'h00000300, 5'd30, 27'h0000006f, 5'd12, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000118, 5'd27, 27'h00000063, 5'd25, 27'h00000186, 32'h00000400,
  1'd1,  5'd26, 27'h00000156, 5'd9, 27'h00000045, 5'd1, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000390, 5'd9, 27'h000002b5, 5'd14, 27'h0000022c, 32'h00000400,
  1'd1,  5'd29, 27'h000001d0, 5'd10, 27'h0000003e, 5'd24, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000103, 5'd16, 27'h000000ba, 5'd1, 27'h00000367, 32'h00000400,
  1'd1,  5'd30, 27'h00000063, 5'd16, 27'h000000eb, 5'd11, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000d3, 5'd20, 27'h00000209, 5'd23, 27'h0000029d, 32'h00000400,
  1'd1,  5'd26, 27'h00000121, 5'd26, 27'h0000021b, 5'd0, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000027d, 5'd30, 27'h000003d1, 5'd15, 27'h00000038, 32'h00000400,
  1'd1,  5'd27, 27'h000000bc, 5'd30, 27'h00000346, 5'd24, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000241, 5'd6, 27'h000001d4, 5'd10, 27'h000000e9, 32'h00000400,
  1'd1,  5'd8, 27'h000001d3, 5'd7, 27'h000000f0, 5'd17, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000097, 5'd10, 27'h00000098, 5'd27, 27'h0000020c, 32'h00000400,
  1'd1,  5'd9, 27'h000003b8, 5'd19, 27'h0000036b, 5'd6, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000358, 5'd17, 27'h00000066, 5'd19, 27'h0000026d, 32'h00000400,
  1'd1,  5'd7, 27'h00000391, 5'd15, 27'h0000024b, 5'd28, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003da, 5'd29, 27'h000002f0, 5'd6, 27'h000003b3, 32'h00000400,
  1'd1,  5'd8, 27'h0000032d, 5'd26, 27'h0000005a, 5'd15, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000374, 5'd28, 27'h0000003c, 5'd26, 27'h0000029c, 32'h00000400,
  1'd1,  5'd15, 27'h00000362, 5'd10, 27'h000000f0, 5'd7, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c8, 5'd8, 27'h000001e3, 5'd19, 27'h000002f0, 32'h00000400,
  1'd1,  5'd16, 27'h0000035b, 5'd9, 27'h00000195, 5'd27, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000003, 5'd16, 27'h00000258, 5'd6, 27'h0000031a, 32'h00000400,
  1'd1,  5'd15, 27'h000002de, 5'd17, 27'h00000399, 5'd19, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011a, 5'd15, 27'h00000206, 5'd30, 27'h000000b4, 32'h00000400,
  1'd1,  5'd20, 27'h0000024f, 5'd27, 27'h00000383, 5'd9, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000241, 5'd29, 27'h000003c6, 5'd19, 27'h000002c0, 32'h00000400,
  1'd1,  5'd17, 27'h00000336, 5'd26, 27'h000001c2, 5'd26, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000f5, 5'd7, 27'h00000194, 5'd8, 27'h00000185, 32'h00000400,
  1'd1,  5'd28, 27'h000001da, 5'd6, 27'h0000030f, 5'd17, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002da, 5'd8, 27'h00000291, 5'd28, 27'h00000164, 32'h00000400,
  1'd1,  5'd27, 27'h00000308, 5'd15, 27'h000003f9, 5'd6, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d0, 5'd15, 27'h00000238, 5'd18, 27'h0000015e, 32'h00000400,
  1'd1,  5'd30, 27'h000003c9, 5'd15, 27'h0000030a, 5'd25, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001be, 5'd27, 27'h00000094, 5'd6, 27'h00000392, 32'h00000400,
  1'd1,  5'd30, 27'h000000c6, 5'd29, 27'h0000036b, 5'd19, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000389, 5'd27, 27'h00000036, 5'd29, 27'h000000f6, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000063, 5'd3, 27'h00000372, 5'd4, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000338, 5'd3, 27'h0000026b, 5'd12, 27'h000002fe, 32'h00000400,
  1'd1,  5'd1, 27'h00000025, 5'd4, 27'h00000244, 5'd20, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000001c, 5'd11, 27'h000001a3, 5'd2, 27'h00000258, 32'h00000400,
  1'd1,  5'd3, 27'h000000da, 5'd14, 27'h0000012c, 5'd15, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a4, 5'd12, 27'h0000012f, 5'd23, 27'h000000a1, 32'h00000400,
  1'd1,  5'd0, 27'h0000008e, 5'd24, 27'h00000261, 5'd2, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000e7, 5'd21, 27'h0000005d, 5'd12, 27'h0000035d, 32'h00000400,
  1'd1,  5'd3, 27'h000001c7, 5'd25, 27'h00000263, 5'd22, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001d7, 5'd2, 27'h00000061, 5'd3, 27'h000002de, 32'h00000400,
  1'd1,  5'd13, 27'h00000021, 5'd2, 27'h000002e4, 5'd11, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c5, 5'd3, 27'h00000033, 5'd23, 27'h00000225, 32'h00000400,
  1'd1,  5'd12, 27'h0000035e, 5'd15, 27'h0000016f, 5'd0, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e5, 5'd15, 27'h000001a1, 5'd10, 27'h000002d8, 32'h00000400,
  1'd1,  5'd10, 27'h0000036b, 5'd13, 27'h000002a7, 5'd23, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000224, 5'd24, 27'h00000377, 5'd3, 27'h00000352, 32'h00000400,
  1'd1,  5'd13, 27'h00000106, 5'd21, 27'h0000020c, 5'd12, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b7, 5'd22, 27'h000001fd, 5'd22, 27'h000003ed, 32'h00000400,
  1'd1,  5'd24, 27'h00000383, 5'd2, 27'h00000234, 5'd2, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000257, 5'd4, 27'h00000062, 5'd12, 27'h00000025, 32'h00000400,
  1'd1,  5'd20, 27'h000003fd, 5'd3, 27'h0000017b, 5'd24, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000213, 5'd12, 27'h000002d1, 5'd3, 27'h00000033, 32'h00000400,
  1'd1,  5'd25, 27'h00000292, 5'd12, 27'h0000039d, 5'd15, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002bd, 5'd12, 27'h00000197, 5'd23, 27'h000000fd, 32'h00000400,
  1'd1,  5'd25, 27'h000001e1, 5'd21, 27'h00000070, 5'd2, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000038b, 5'd25, 27'h00000332, 5'd15, 27'h00000157, 32'h00000400,
  1'd1,  5'd21, 27'h0000030b, 5'd21, 27'h000003ab, 5'd24, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000027, 5'd4, 27'h000000e8, 5'd6, 27'h00000092, 32'h00000400,
  1'd1,  5'd3, 27'h000002f7, 5'd4, 27'h0000011f, 5'd17, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000018e, 5'd5, 27'h0000009f, 5'd27, 27'h00000045, 32'h00000400,
  1'd1,  5'd5, 27'h00000020, 5'd10, 27'h0000032d, 5'd7, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000af, 5'd14, 27'h000001b8, 5'd17, 27'h000003b0, 32'h00000400,
  1'd1,  5'd3, 27'h0000001b, 5'd11, 27'h000001f3, 5'd28, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000160, 5'd23, 27'h0000030b, 5'd5, 27'h00000301, 32'h00000400,
  1'd1,  5'd1, 27'h0000016f, 5'd21, 27'h00000361, 5'd16, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000037f, 5'd21, 27'h00000370, 5'd29, 27'h000001c7, 32'h00000400,
  1'd1,  5'd11, 27'h000002b4, 5'd3, 27'h0000005d, 5'd8, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013b, 5'd2, 27'h000003bf, 5'd17, 27'h000000d2, 32'h00000400,
  1'd1,  5'd13, 27'h000002f5, 5'd4, 27'h000001f0, 5'd26, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000188, 5'd10, 27'h000001a5, 5'd9, 27'h0000034d, 32'h00000400,
  1'd1,  5'd12, 27'h00000240, 5'd11, 27'h000000f2, 5'd18, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000391, 5'd10, 27'h00000159, 5'd30, 27'h00000345, 32'h00000400,
  1'd1,  5'd11, 27'h0000017b, 5'd23, 27'h000002fb, 5'd8, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000db, 5'd21, 27'h00000206, 5'd17, 27'h000002e1, 32'h00000400,
  1'd1,  5'd15, 27'h000000fc, 5'd21, 27'h000002ce, 5'd28, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000023, 5'd2, 27'h00000341, 5'd8, 27'h000000b6, 32'h00000400,
  1'd1,  5'd23, 27'h0000031e, 5'd4, 27'h0000014a, 5'd18, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000099, 5'd3, 27'h00000156, 5'd29, 27'h00000387, 32'h00000400,
  1'd1,  5'd21, 27'h000001a1, 5'd14, 27'h00000190, 5'd8, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000128, 5'd11, 27'h000003a4, 5'd16, 27'h000001d8, 32'h00000400,
  1'd1,  5'd25, 27'h0000011d, 5'd13, 27'h000001bb, 5'd30, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000028e, 5'd25, 27'h00000301, 5'd10, 27'h00000107, 32'h00000400,
  1'd1,  5'd22, 27'h000001b3, 5'd21, 27'h0000035b, 5'd17, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000072, 5'd24, 27'h000002d7, 5'd29, 27'h0000031c, 32'h00000400,
  1'd1,  5'd0, 27'h000003cb, 5'd8, 27'h000001a1, 5'd3, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000007f, 5'd10, 27'h0000008f, 5'd13, 27'h00000357, 32'h00000400,
  1'd1,  5'd0, 27'h00000130, 5'd10, 27'h00000137, 5'd23, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c8, 5'd16, 27'h000003ea, 5'd2, 27'h00000342, 32'h00000400,
  1'd1,  5'd1, 27'h00000353, 5'd18, 27'h000000f1, 5'd11, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000088, 5'd16, 27'h000000c7, 5'd24, 27'h000003c3, 32'h00000400,
  1'd1,  5'd4, 27'h00000159, 5'd26, 27'h00000154, 5'd1, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000120, 5'd26, 27'h000003fd, 5'd12, 27'h00000155, 32'h00000400,
  1'd1,  5'd1, 27'h0000029c, 5'd28, 27'h0000027e, 5'd22, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000036f, 5'd5, 27'h0000026a, 5'd1, 27'h0000036f, 32'h00000400,
  1'd1,  5'd14, 27'h000002c4, 5'd8, 27'h00000389, 5'd15, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ad, 5'd7, 27'h000002ec, 5'd23, 27'h00000112, 32'h00000400,
  1'd1,  5'd13, 27'h000002cb, 5'd19, 27'h000003e3, 5'd1, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000007c, 5'd18, 27'h000001bc, 5'd12, 27'h000002c9, 32'h00000400,
  1'd1,  5'd14, 27'h000002ad, 5'd18, 27'h0000022d, 5'd21, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c2, 5'd30, 27'h0000020f, 5'd2, 27'h0000005b, 32'h00000400,
  1'd1,  5'd10, 27'h00000333, 5'd27, 27'h000000c5, 5'd13, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001c7, 5'd27, 27'h000000ec, 5'd24, 27'h000002e8, 32'h00000400,
  1'd1,  5'd23, 27'h000001dc, 5'd8, 27'h0000030d, 5'd4, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000352, 5'd8, 27'h000003db, 5'd12, 27'h00000219, 32'h00000400,
  1'd1,  5'd21, 27'h0000030e, 5'd9, 27'h000001ca, 5'd24, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000286, 5'd20, 27'h00000275, 5'd2, 27'h000000bc, 32'h00000400,
  1'd1,  5'd24, 27'h000003e0, 5'd18, 27'h00000083, 5'd11, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000240, 5'd17, 27'h00000116, 5'd20, 27'h0000030a, 32'h00000400,
  1'd1,  5'd21, 27'h000003b2, 5'd27, 27'h00000352, 5'd1, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000166, 5'd26, 27'h0000036c, 5'd15, 27'h00000048, 32'h00000400,
  1'd1,  5'd23, 27'h000003c6, 5'd26, 27'h000001ef, 5'd21, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b7, 5'd8, 27'h000002a8, 5'd7, 27'h0000022d, 32'h00000400,
  1'd1,  5'd3, 27'h000000ec, 5'd7, 27'h000003a1, 5'd19, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002b0, 5'd10, 27'h000000a0, 5'd28, 27'h00000279, 32'h00000400,
  1'd1,  5'd0, 27'h00000025, 5'd20, 27'h0000022b, 5'd6, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000037f, 5'd17, 27'h00000187, 5'd20, 27'h00000263, 32'h00000400,
  1'd1,  5'd4, 27'h000001db, 5'd15, 27'h00000268, 5'd28, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002fd, 5'd27, 27'h000002d5, 5'd5, 27'h00000299, 32'h00000400,
  1'd1,  5'd3, 27'h00000091, 5'd26, 27'h00000143, 5'd20, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a8, 5'd28, 27'h00000304, 5'd29, 27'h000003cf, 32'h00000400,
  1'd1,  5'd11, 27'h0000016a, 5'd8, 27'h0000008c, 5'd7, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000267, 5'd7, 27'h000002ee, 5'd17, 27'h00000345, 32'h00000400,
  1'd1,  5'd11, 27'h000001f4, 5'd10, 27'h0000012b, 5'd27, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001fe, 5'd17, 27'h000001b3, 5'd5, 27'h00000296, 32'h00000400,
  1'd1,  5'd15, 27'h000000e8, 5'd16, 27'h000002f3, 5'd20, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000021, 5'd18, 27'h000001ce, 5'd26, 27'h000002b6, 32'h00000400,
  1'd1,  5'd10, 27'h000003f4, 5'd26, 27'h000001d5, 5'd5, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f8, 5'd28, 27'h00000321, 5'd16, 27'h000001fb, 32'h00000400,
  1'd1,  5'd15, 27'h00000013, 5'd26, 27'h0000008d, 5'd26, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f3, 5'd8, 27'h00000150, 5'd9, 27'h000001a7, 32'h00000400,
  1'd1,  5'd21, 27'h000000d0, 5'd9, 27'h000000d3, 5'd19, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000155, 5'd6, 27'h00000262, 5'd26, 27'h0000002e, 32'h00000400,
  1'd1,  5'd20, 27'h000003fd, 5'd18, 27'h000001d4, 5'd9, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000016d, 5'd20, 27'h00000016, 5'd16, 27'h000003c5, 32'h00000400,
  1'd1,  5'd21, 27'h0000021e, 5'd16, 27'h0000033b, 5'd30, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000323, 5'd28, 27'h0000038d, 5'd9, 27'h00000220, 32'h00000400,
  1'd1,  5'd23, 27'h00000184, 5'd27, 27'h0000012e, 5'd19, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000387, 5'd26, 27'h000001c2, 5'd30, 27'h000002a6, 32'h00000400,
  1'd1,  5'd9, 27'h000001fe, 5'd3, 27'h00000048, 5'd6, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001e2, 5'd2, 27'h00000289, 5'd15, 27'h0000022b, 32'h00000400,
  1'd1,  5'd5, 27'h00000196, 5'd1, 27'h000000c1, 5'd29, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001b1, 5'd15, 27'h000001ec, 5'd2, 27'h00000169, 32'h00000400,
  1'd1,  5'd7, 27'h000002b9, 5'd15, 27'h000001c8, 5'd14, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000027, 5'd15, 27'h000001fc, 5'd21, 27'h000001f7, 32'h00000400,
  1'd1,  5'd7, 27'h00000186, 5'd20, 27'h00000368, 5'd1, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000029, 5'd20, 27'h000002fc, 5'd11, 27'h00000212, 32'h00000400,
  1'd1,  5'd5, 27'h00000212, 5'd20, 27'h000002ab, 5'd22, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000017a, 5'd4, 27'h00000048, 5'd10, 27'h000000b7, 32'h00000400,
  1'd1,  5'd19, 27'h000001a2, 5'd0, 27'h000003eb, 5'd17, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d6, 5'd2, 27'h000002d3, 5'd25, 27'h00000367, 32'h00000400,
  1'd1,  5'd17, 27'h00000054, 5'd14, 27'h00000385, 5'd3, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016b, 5'd12, 27'h00000355, 5'd11, 27'h0000034f, 32'h00000400,
  1'd1,  5'd17, 27'h00000158, 5'd11, 27'h00000347, 5'd21, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001e0, 5'd20, 27'h000002fd, 5'd2, 27'h00000163, 32'h00000400,
  1'd1,  5'd16, 27'h000003cf, 5'd24, 27'h00000222, 5'd13, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000009d, 5'd21, 27'h000003ac, 5'd23, 27'h000003c4, 32'h00000400,
  1'd1,  5'd25, 27'h000003cb, 5'd0, 27'h00000133, 5'd4, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000001, 5'd3, 27'h00000344, 5'd12, 27'h0000002b, 32'h00000400,
  1'd1,  5'd29, 27'h00000145, 5'd4, 27'h00000188, 5'd25, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003ea, 5'd13, 27'h000003c2, 5'd3, 27'h0000030b, 32'h00000400,
  1'd1,  5'd29, 27'h000003af, 5'd10, 27'h000003b2, 5'd11, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d1, 5'd12, 27'h00000321, 5'd24, 27'h00000124, 32'h00000400,
  1'd1,  5'd27, 27'h0000020e, 5'd24, 27'h000001b6, 5'd4, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000352, 5'd20, 27'h00000399, 5'd11, 27'h00000062, 32'h00000400,
  1'd1,  5'd28, 27'h0000017f, 5'd20, 27'h000002bb, 5'd21, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000102, 5'd5, 27'h00000006, 5'd4, 27'h00000013, 32'h00000400,
  1'd1,  5'd6, 27'h000000ac, 5'd2, 27'h00000397, 5'd11, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ea, 5'd1, 27'h000002f1, 5'd25, 27'h000002a7, 32'h00000400,
  1'd1,  5'd6, 27'h000002d2, 5'd11, 27'h00000330, 5'd6, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000124, 5'd12, 27'h0000037a, 5'd17, 27'h000000f3, 32'h00000400,
  1'd1,  5'd5, 27'h0000014a, 5'd13, 27'h00000275, 5'd30, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012d, 5'd21, 27'h0000013c, 5'd6, 27'h000003d1, 32'h00000400,
  1'd1,  5'd8, 27'h0000000f, 5'd23, 27'h0000039e, 5'd19, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a9, 5'd23, 27'h0000023f, 5'd29, 27'h00000170, 32'h00000400,
  1'd1,  5'd17, 27'h00000212, 5'd3, 27'h00000231, 5'd3, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000003c, 5'd2, 27'h00000068, 5'd11, 27'h00000280, 32'h00000400,
  1'd1,  5'd18, 27'h0000006b, 5'd4, 27'h000003bc, 5'd23, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000013d, 5'd10, 27'h00000181, 5'd6, 27'h0000028f, 32'h00000400,
  1'd1,  5'd18, 27'h00000215, 5'd12, 27'h0000014a, 5'd16, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a9, 5'd12, 27'h000002a8, 5'd27, 27'h00000353, 32'h00000400,
  1'd1,  5'd15, 27'h000003f8, 5'd20, 27'h00000384, 5'd5, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000003c, 5'd21, 27'h000003f0, 5'd20, 27'h0000023b, 32'h00000400,
  1'd1,  5'd18, 27'h0000020e, 5'd22, 27'h00000324, 5'd27, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000016c, 5'd1, 27'h00000051, 5'd7, 27'h000003ec, 32'h00000400,
  1'd1,  5'd26, 27'h00000069, 5'd1, 27'h000001a7, 5'd15, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000005e, 5'd0, 27'h000002b0, 5'd27, 27'h0000003c, 32'h00000400,
  1'd1,  5'd28, 27'h000002bd, 5'd10, 27'h00000350, 5'd5, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f4, 5'd14, 27'h0000008d, 5'd15, 27'h000002b9, 32'h00000400,
  1'd1,  5'd27, 27'h000002e2, 5'd13, 27'h00000370, 5'd27, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000006c, 5'd24, 27'h00000044, 5'd5, 27'h000002e4, 32'h00000400,
  1'd1,  5'd27, 27'h00000334, 5'd22, 27'h000000dc, 5'd18, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000156, 5'd24, 27'h00000319, 5'd30, 27'h0000000d, 32'h00000400,
  1'd1,  5'd8, 27'h0000021f, 5'd5, 27'h0000029f, 5'd1, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000060, 5'd7, 27'h0000016d, 5'd13, 27'h0000021f, 32'h00000400,
  1'd1,  5'd6, 27'h000002b2, 5'd5, 27'h0000020c, 5'd23, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000222, 5'd16, 27'h0000030a, 5'd3, 27'h0000009e, 32'h00000400,
  1'd1,  5'd8, 27'h000002fe, 5'd15, 27'h00000318, 5'd12, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000021e, 5'd17, 27'h00000324, 5'd25, 27'h00000138, 32'h00000400,
  1'd1,  5'd6, 27'h000003cd, 5'd30, 27'h00000215, 5'd3, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000076, 5'd30, 27'h00000304, 5'd11, 27'h000002f9, 32'h00000400,
  1'd1,  5'd10, 27'h00000033, 5'd29, 27'h000001db, 5'd22, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002da, 5'd6, 27'h00000229, 5'd3, 27'h00000370, 32'h00000400,
  1'd1,  5'd20, 27'h0000002a, 5'd5, 27'h0000035f, 5'd13, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000025a, 5'd8, 27'h00000338, 5'd22, 27'h00000105, 32'h00000400,
  1'd1,  5'd16, 27'h00000145, 5'd16, 27'h0000035c, 5'd1, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a9, 5'd17, 27'h0000023a, 5'd14, 27'h000003c7, 32'h00000400,
  1'd1,  5'd16, 27'h000000c5, 5'd15, 27'h000003b4, 5'd22, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b1, 5'd30, 27'h0000017e, 5'd1, 27'h0000007a, 32'h00000400,
  1'd1,  5'd16, 27'h0000020b, 5'd26, 27'h0000003a, 5'd14, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000308, 5'd30, 27'h000003f4, 5'd23, 27'h00000346, 32'h00000400,
  1'd1,  5'd27, 27'h00000039, 5'd9, 27'h000002b4, 5'd0, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000361, 5'd9, 27'h00000074, 5'd12, 27'h00000029, 32'h00000400,
  1'd1,  5'd27, 27'h000001b3, 5'd6, 27'h000003a1, 5'd24, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000014b, 5'd19, 27'h00000291, 5'd3, 27'h000003d6, 32'h00000400,
  1'd1,  5'd26, 27'h00000343, 5'd19, 27'h00000230, 5'd10, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003db, 5'd19, 27'h000003cf, 5'd25, 27'h000001a1, 32'h00000400,
  1'd1,  5'd29, 27'h00000349, 5'd27, 27'h00000226, 5'd4, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002de, 5'd26, 27'h00000258, 5'd13, 27'h000000aa, 32'h00000400,
  1'd1,  5'd29, 27'h000001ba, 5'd26, 27'h00000317, 5'd22, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002d0, 5'd5, 27'h000002f6, 5'd6, 27'h0000001e, 32'h00000400,
  1'd1,  5'd5, 27'h000003a3, 5'd8, 27'h00000197, 5'd19, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000c2, 5'd8, 27'h000000e8, 5'd30, 27'h000002dd, 32'h00000400,
  1'd1,  5'd10, 27'h00000091, 5'd18, 27'h00000074, 5'd5, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033d, 5'd19, 27'h000002ec, 5'd17, 27'h00000313, 32'h00000400,
  1'd1,  5'd8, 27'h000001e8, 5'd20, 27'h00000253, 5'd28, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000112, 5'd28, 27'h000003c0, 5'd5, 27'h000002f2, 32'h00000400,
  1'd1,  5'd7, 27'h00000197, 5'd29, 27'h0000003b, 5'd17, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000006f, 5'd28, 27'h0000029b, 5'd28, 27'h00000202, 32'h00000400,
  1'd1,  5'd15, 27'h00000324, 5'd9, 27'h00000357, 5'd7, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000006, 5'd9, 27'h00000172, 5'd20, 27'h0000019f, 32'h00000400,
  1'd1,  5'd19, 27'h000002f8, 5'd10, 27'h00000055, 5'd28, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000165, 5'd17, 27'h00000044, 5'd5, 27'h00000340, 32'h00000400,
  1'd1,  5'd19, 27'h0000022c, 5'd16, 27'h00000372, 5'd17, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000022, 5'd19, 27'h000001a0, 5'd28, 27'h00000162, 32'h00000400,
  1'd1,  5'd18, 27'h0000019a, 5'd28, 27'h000000bb, 5'd9, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002f0, 5'd30, 27'h0000018e, 5'd19, 27'h000000f1, 32'h00000400,
  1'd1,  5'd15, 27'h00000321, 5'd27, 27'h00000243, 5'd26, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000b6, 5'd9, 27'h0000003e, 5'd8, 27'h0000020d, 32'h00000400,
  1'd1,  5'd28, 27'h000001de, 5'd6, 27'h00000064, 5'd16, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e6, 5'd10, 27'h00000027, 5'd29, 27'h00000175, 32'h00000400,
  1'd1,  5'd27, 27'h0000003a, 5'd18, 27'h00000198, 5'd9, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000b4, 5'd17, 27'h00000067, 5'd18, 27'h0000012b, 32'h00000400,
  1'd1,  5'd29, 27'h00000148, 5'd20, 27'h0000008f, 5'd30, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000101, 5'd26, 27'h000002c9, 5'd8, 27'h00000285, 32'h00000400,
  1'd1,  5'd28, 27'h00000304, 5'd30, 27'h000000de, 5'd18, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000133, 5'd28, 27'h00000093, 5'd29, 27'h000001f6, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003bc, 5'd1, 27'h0000004e, 5'd1, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000156, 5'd0, 27'h00000067, 5'd15, 27'h000001ba, 32'h00000400,
  1'd1,  5'd0, 27'h0000026e, 5'd2, 27'h000002fc, 5'd25, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000058, 5'd14, 27'h0000015c, 5'd4, 27'h00000388, 32'h00000400,
  1'd1,  5'd3, 27'h000002ac, 5'd14, 27'h00000046, 5'd14, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000029e, 5'd14, 27'h00000351, 5'd24, 27'h00000256, 32'h00000400,
  1'd1,  5'd1, 27'h0000019e, 5'd25, 27'h000000ac, 5'd1, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000251, 5'd25, 27'h0000016a, 5'd14, 27'h000001e4, 32'h00000400,
  1'd1,  5'd0, 27'h00000177, 5'd21, 27'h00000229, 5'd22, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ec, 5'd2, 27'h000000bc, 5'd1, 27'h0000020e, 32'h00000400,
  1'd1,  5'd13, 27'h000003ea, 5'd0, 27'h000000aa, 5'd13, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000345, 5'd1, 27'h000003d3, 5'd23, 27'h000001c3, 32'h00000400,
  1'd1,  5'd13, 27'h00000076, 5'd10, 27'h000003f4, 5'd2, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000176, 5'd14, 27'h000000fe, 5'd14, 27'h00000101, 32'h00000400,
  1'd1,  5'd11, 27'h000002ae, 5'd11, 27'h0000009f, 5'd23, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000115, 5'd25, 27'h00000286, 5'd0, 27'h0000022a, 32'h00000400,
  1'd1,  5'd12, 27'h00000180, 5'd22, 27'h000002a3, 5'd14, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000040, 5'd22, 27'h00000032, 5'd24, 27'h000002d7, 32'h00000400,
  1'd1,  5'd21, 27'h0000026d, 5'd4, 27'h00000043, 5'd0, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000305, 5'd4, 27'h00000210, 5'd12, 27'h00000376, 32'h00000400,
  1'd1,  5'd24, 27'h000000bf, 5'd4, 27'h000001e0, 5'd20, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ed, 5'd13, 27'h00000228, 5'd2, 27'h000001ac, 32'h00000400,
  1'd1,  5'd24, 27'h000003d3, 5'd10, 27'h000001cf, 5'd14, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000063, 5'd12, 27'h00000273, 5'd24, 27'h000001a9, 32'h00000400,
  1'd1,  5'd21, 27'h000003ca, 5'd21, 27'h0000003e, 5'd1, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000309, 5'd24, 27'h000001cb, 5'd10, 27'h00000295, 32'h00000400,
  1'd1,  5'd22, 27'h00000372, 5'd25, 27'h00000173, 5'd22, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026a, 5'd4, 27'h00000126, 5'd7, 27'h000000e2, 32'h00000400,
  1'd1,  5'd1, 27'h000000da, 5'd2, 27'h0000015f, 5'd19, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000009c, 5'd4, 27'h000001ee, 5'd25, 27'h000003ae, 32'h00000400,
  1'd1,  5'd0, 27'h0000017b, 5'd11, 27'h000001d8, 5'd7, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001ae, 5'd10, 27'h00000395, 5'd16, 27'h000000fb, 32'h00000400,
  1'd1,  5'd0, 27'h0000027f, 5'd12, 27'h000000ce, 5'd30, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000fe, 5'd23, 27'h0000026f, 5'd7, 27'h00000216, 32'h00000400,
  1'd1,  5'd1, 27'h0000030c, 5'd25, 27'h00000172, 5'd15, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e9, 5'd21, 27'h00000361, 5'd27, 27'h00000235, 32'h00000400,
  1'd1,  5'd12, 27'h00000389, 5'd0, 27'h000001ee, 5'd9, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c0, 5'd1, 27'h0000032f, 5'd19, 27'h00000353, 32'h00000400,
  1'd1,  5'd12, 27'h000000a6, 5'd2, 27'h0000016a, 5'd30, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001e7, 5'd12, 27'h00000115, 5'd5, 27'h000001e8, 32'h00000400,
  1'd1,  5'd12, 27'h000001c6, 5'd14, 27'h000001b1, 5'd19, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001bb, 5'd10, 27'h00000388, 5'd29, 27'h000003a9, 32'h00000400,
  1'd1,  5'd13, 27'h00000197, 5'd22, 27'h0000004b, 5'd7, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000306, 5'd21, 27'h000001f2, 5'd19, 27'h000001f7, 32'h00000400,
  1'd1,  5'd14, 27'h0000038a, 5'd25, 27'h000001ff, 5'd26, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000026e, 5'd4, 27'h000001a8, 5'd9, 27'h0000016d, 32'h00000400,
  1'd1,  5'd24, 27'h000001e8, 5'd1, 27'h000002b0, 5'd20, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f1, 5'd4, 27'h0000021f, 5'd26, 27'h000003a8, 32'h00000400,
  1'd1,  5'd25, 27'h0000025f, 5'd15, 27'h00000123, 5'd6, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f3, 5'd11, 27'h00000116, 5'd17, 27'h00000074, 32'h00000400,
  1'd1,  5'd24, 27'h000000cf, 5'd12, 27'h000000f9, 5'd29, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002bf, 5'd20, 27'h00000358, 5'd10, 27'h000000de, 32'h00000400,
  1'd1,  5'd24, 27'h000000a0, 5'd23, 27'h0000002c, 5'd19, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000313, 5'd25, 27'h00000341, 5'd30, 27'h0000005b, 32'h00000400,
  1'd1,  5'd4, 27'h000001e7, 5'd6, 27'h000000f9, 5'd1, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000071, 5'd10, 27'h00000129, 5'd11, 27'h000002fc, 32'h00000400,
  1'd1,  5'd2, 27'h00000187, 5'd6, 27'h000002b2, 5'd21, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000146, 5'd15, 27'h0000039c, 5'd2, 27'h00000171, 32'h00000400,
  1'd1,  5'd1, 27'h000001a6, 5'd20, 27'h000000aa, 5'd13, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000047, 5'd19, 27'h000003ec, 5'd22, 27'h000003c5, 32'h00000400,
  1'd1,  5'd1, 27'h0000015d, 5'd30, 27'h000003c5, 5'd1, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000056, 5'd30, 27'h000000fe, 5'd12, 27'h0000000d, 32'h00000400,
  1'd1,  5'd0, 27'h0000020c, 5'd29, 27'h000000d8, 5'd21, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f4, 5'd6, 27'h00000373, 5'd4, 27'h0000020a, 32'h00000400,
  1'd1,  5'd14, 27'h00000001, 5'd8, 27'h00000320, 5'd12, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000fa, 5'd7, 27'h00000118, 5'd23, 27'h000001f2, 32'h00000400,
  1'd1,  5'd13, 27'h000002fb, 5'd15, 27'h00000225, 5'd0, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000244, 5'd17, 27'h000001d9, 5'd11, 27'h0000000e, 32'h00000400,
  1'd1,  5'd14, 27'h00000235, 5'd20, 27'h000001cb, 5'd24, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e8, 5'd29, 27'h00000281, 5'd1, 27'h00000119, 32'h00000400,
  1'd1,  5'd13, 27'h00000272, 5'd28, 27'h00000298, 5'd11, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000298, 5'd26, 27'h00000287, 5'd20, 27'h00000389, 32'h00000400,
  1'd1,  5'd22, 27'h0000013e, 5'd9, 27'h00000151, 5'd2, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000028e, 5'd5, 27'h000001a0, 5'd12, 27'h00000138, 32'h00000400,
  1'd1,  5'd21, 27'h000001fa, 5'd7, 27'h000001be, 5'd21, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000373, 5'd19, 27'h0000016f, 5'd0, 27'h0000022c, 32'h00000400,
  1'd1,  5'd23, 27'h00000331, 5'd15, 27'h000002fc, 5'd11, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000012, 5'd18, 27'h0000011d, 5'd23, 27'h000002a7, 32'h00000400,
  1'd1,  5'd21, 27'h000003e8, 5'd27, 27'h00000168, 5'd2, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000278, 5'd29, 27'h000003c7, 5'd14, 27'h00000021, 32'h00000400,
  1'd1,  5'd25, 27'h000002a9, 5'd30, 27'h000003ea, 5'd22, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002c6, 5'd10, 27'h0000001d, 5'd5, 27'h000001c8, 32'h00000400,
  1'd1,  5'd1, 27'h00000047, 5'd6, 27'h000002de, 5'd18, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000037f, 5'd9, 27'h000002eb, 5'd26, 27'h000002c3, 32'h00000400,
  1'd1,  5'd2, 27'h000002fc, 5'd16, 27'h00000039, 5'd6, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000032d, 5'd16, 27'h00000013, 5'd16, 27'h000000a9, 32'h00000400,
  1'd1,  5'd4, 27'h0000030d, 5'd19, 27'h0000025d, 5'd28, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000392, 5'd25, 27'h000003f0, 5'd9, 27'h000003a0, 32'h00000400,
  1'd1,  5'd4, 27'h000000af, 5'd27, 27'h00000151, 5'd16, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000201, 5'd27, 27'h00000349, 5'd27, 27'h0000018f, 32'h00000400,
  1'd1,  5'd14, 27'h000001ff, 5'd7, 27'h00000016, 5'd9, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fa, 5'd7, 27'h00000350, 5'd20, 27'h00000177, 32'h00000400,
  1'd1,  5'd14, 27'h000001cc, 5'd10, 27'h0000000c, 5'd26, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003b3, 5'd18, 27'h0000035e, 5'd8, 27'h0000007d, 32'h00000400,
  1'd1,  5'd15, 27'h000001a6, 5'd19, 27'h00000117, 5'd15, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001bb, 5'd16, 27'h000001f4, 5'd30, 27'h0000004b, 32'h00000400,
  1'd1,  5'd15, 27'h000000d0, 5'd26, 27'h00000248, 5'd8, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000041, 5'd29, 27'h0000011a, 5'd19, 27'h00000068, 32'h00000400,
  1'd1,  5'd12, 27'h000003c8, 5'd29, 27'h0000007d, 5'd29, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003a4, 5'd8, 27'h000003ce, 5'd6, 27'h0000038e, 32'h00000400,
  1'd1,  5'd21, 27'h00000227, 5'd10, 27'h00000103, 5'd16, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000382, 5'd6, 27'h000000bb, 5'd30, 27'h00000147, 32'h00000400,
  1'd1,  5'd21, 27'h00000169, 5'd15, 27'h0000032a, 5'd6, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000226, 5'd19, 27'h000003e8, 5'd15, 27'h0000027c, 32'h00000400,
  1'd1,  5'd24, 27'h00000341, 5'd20, 27'h000001e4, 5'd28, 27'h00000370, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000371, 5'd30, 27'h00000245, 5'd8, 27'h00000045, 32'h00000400,
  1'd1,  5'd22, 27'h0000012c, 5'd30, 27'h000001f0, 5'd15, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000017a, 5'd30, 27'h000000c8, 5'd26, 27'h0000032e, 32'h00000400,
  1'd1,  5'd5, 27'h00000387, 5'd3, 27'h000000c9, 5'd8, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002b6, 5'd2, 27'h000002dd, 5'd18, 27'h000002dd, 32'h00000400,
  1'd1,  5'd5, 27'h00000176, 5'd1, 27'h00000383, 5'd26, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000061, 5'd15, 27'h000001d3, 5'd4, 27'h00000382, 32'h00000400,
  1'd1,  5'd9, 27'h00000056, 5'd11, 27'h000003ef, 5'd11, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001d2, 5'd12, 27'h0000033e, 5'd22, 27'h00000298, 32'h00000400,
  1'd1,  5'd7, 27'h000001a6, 5'd22, 27'h000002a9, 5'd3, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003c0, 5'd22, 27'h0000025c, 5'd13, 27'h00000144, 32'h00000400,
  1'd1,  5'd9, 27'h000000e0, 5'd21, 27'h00000346, 5'd22, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001f2, 5'd3, 27'h00000000, 5'd7, 27'h000000a1, 32'h00000400,
  1'd1,  5'd19, 27'h0000034a, 5'd2, 27'h00000306, 5'd16, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000ac, 5'd0, 27'h0000008b, 5'd26, 27'h0000003e, 32'h00000400,
  1'd1,  5'd18, 27'h00000298, 5'd12, 27'h000001d1, 5'd4, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000006f, 5'd14, 27'h000000c3, 5'd12, 27'h000000d7, 32'h00000400,
  1'd1,  5'd17, 27'h00000230, 5'd10, 27'h00000297, 5'd24, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000030f, 5'd20, 27'h000002e3, 5'd1, 27'h00000124, 32'h00000400,
  1'd1,  5'd18, 27'h00000270, 5'd20, 27'h00000354, 5'd10, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000000c, 5'd24, 27'h00000094, 5'd23, 27'h000003ea, 32'h00000400,
  1'd1,  5'd26, 27'h00000391, 5'd4, 27'h000003af, 5'd3, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000ef, 5'd2, 27'h00000043, 5'd13, 27'h0000038d, 32'h00000400,
  1'd1,  5'd27, 27'h0000030a, 5'd2, 27'h00000296, 5'd25, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000328, 5'd10, 27'h00000382, 5'd3, 27'h00000050, 32'h00000400,
  1'd1,  5'd28, 27'h0000017b, 5'd14, 27'h00000067, 5'd15, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000341, 5'd13, 27'h00000381, 5'd21, 27'h0000000d, 32'h00000400,
  1'd1,  5'd27, 27'h00000387, 5'd21, 27'h00000388, 5'd2, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000039b, 5'd21, 27'h000000ed, 5'd10, 27'h00000245, 32'h00000400,
  1'd1,  5'd28, 27'h000002ff, 5'd25, 27'h00000316, 5'd25, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000247, 5'd4, 27'h00000047, 5'd5, 27'h00000028, 32'h00000400,
  1'd1,  5'd5, 27'h000003d0, 5'd2, 27'h000002f7, 5'd10, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000003e, 5'd3, 27'h00000233, 5'd23, 27'h0000002a, 32'h00000400,
  1'd1,  5'd9, 27'h00000259, 5'd12, 27'h000003fd, 5'd8, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000281, 5'd12, 27'h00000024, 5'd19, 27'h0000014d, 32'h00000400,
  1'd1,  5'd8, 27'h000000f9, 5'd12, 27'h000003ee, 5'd30, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000025, 5'd24, 27'h000000cb, 5'd9, 27'h00000075, 32'h00000400,
  1'd1,  5'd5, 27'h00000318, 5'd23, 27'h00000183, 5'd18, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000f8, 5'd22, 27'h000000fe, 5'd26, 27'h000002fc, 32'h00000400,
  1'd1,  5'd19, 27'h0000023b, 5'd1, 27'h00000299, 5'd2, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000328, 5'd2, 27'h0000005c, 5'd14, 27'h0000023a, 32'h00000400,
  1'd1,  5'd17, 27'h0000012d, 5'd0, 27'h000003d1, 5'd20, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000db, 5'd13, 27'h000001d4, 5'd9, 27'h000000b6, 32'h00000400,
  1'd1,  5'd16, 27'h00000217, 5'd11, 27'h000001e7, 5'd18, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000038a, 5'd12, 27'h00000035, 5'd29, 27'h00000358, 32'h00000400,
  1'd1,  5'd16, 27'h00000116, 5'd25, 27'h00000059, 5'd9, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000004d, 5'd23, 27'h00000377, 5'd17, 27'h0000011b, 32'h00000400,
  1'd1,  5'd16, 27'h00000013, 5'd21, 27'h000001f1, 5'd26, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001dc, 5'd3, 27'h00000183, 5'd8, 27'h0000015b, 32'h00000400,
  1'd1,  5'd30, 27'h00000173, 5'd4, 27'h000001d7, 5'd17, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000307, 5'd3, 27'h00000253, 5'd30, 27'h000000a3, 32'h00000400,
  1'd1,  5'd28, 27'h00000123, 5'd13, 27'h000001ff, 5'd5, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002cb, 5'd14, 27'h00000082, 5'd16, 27'h000003f6, 32'h00000400,
  1'd1,  5'd26, 27'h00000360, 5'd12, 27'h000002ff, 5'd29, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000012e, 5'd25, 27'h0000008e, 5'd6, 27'h000000a4, 32'h00000400,
  1'd1,  5'd27, 27'h000003ff, 5'd23, 27'h000000a8, 5'd19, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e1, 5'd24, 27'h000000a6, 5'd28, 27'h00000038, 32'h00000400,
  1'd1,  5'd5, 27'h000002e7, 5'd7, 27'h000000b8, 5'd0, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000285, 5'd9, 27'h00000027, 5'd14, 27'h000003b3, 32'h00000400,
  1'd1,  5'd5, 27'h00000333, 5'd8, 27'h000003ab, 5'd21, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000059, 5'd17, 27'h000002fe, 5'd0, 27'h000002e8, 32'h00000400,
  1'd1,  5'd6, 27'h0000003c, 5'd20, 27'h00000251, 5'd12, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000331, 5'd18, 27'h00000112, 5'd24, 27'h000000a3, 32'h00000400,
  1'd1,  5'd8, 27'h00000106, 5'd28, 27'h000002f8, 5'd1, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002f3, 5'd28, 27'h000000b9, 5'd14, 27'h00000398, 32'h00000400,
  1'd1,  5'd9, 27'h0000012f, 5'd26, 27'h0000027a, 5'd24, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000092, 5'd8, 27'h00000096, 5'd4, 27'h0000022c, 32'h00000400,
  1'd1,  5'd20, 27'h000001aa, 5'd6, 27'h00000253, 5'd13, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000018, 5'd8, 27'h00000187, 5'd21, 27'h00000016, 32'h00000400,
  1'd1,  5'd16, 27'h000003aa, 5'd19, 27'h00000098, 5'd4, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000039, 5'd19, 27'h000003ab, 5'd13, 27'h000001ee, 32'h00000400,
  1'd1,  5'd17, 27'h0000025c, 5'd17, 27'h00000005, 5'd22, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f1, 5'd29, 27'h000001b8, 5'd4, 27'h000000ce, 32'h00000400,
  1'd1,  5'd18, 27'h000003e2, 5'd29, 27'h000000eb, 5'd12, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000265, 5'd27, 27'h00000070, 5'd21, 27'h00000262, 32'h00000400,
  1'd1,  5'd27, 27'h0000024e, 5'd7, 27'h000003da, 5'd4, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002c7, 5'd9, 27'h0000030c, 5'd12, 27'h00000041, 32'h00000400,
  1'd1,  5'd27, 27'h00000154, 5'd7, 27'h00000215, 5'd22, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000037e, 5'd17, 27'h0000027f, 5'd1, 27'h000002cc, 32'h00000400,
  1'd1,  5'd30, 27'h000003cb, 5'd20, 27'h00000129, 5'd13, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000020f, 5'd17, 27'h000002b7, 5'd20, 27'h00000318, 32'h00000400,
  1'd1,  5'd27, 27'h00000124, 5'd30, 27'h00000056, 5'd0, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000240, 5'd27, 27'h00000003, 5'd14, 27'h000001d4, 32'h00000400,
  1'd1,  5'd26, 27'h000002e3, 5'd26, 27'h000003fe, 5'd25, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a7, 5'd9, 27'h000003cd, 5'd5, 27'h000000ad, 32'h00000400,
  1'd1,  5'd9, 27'h0000023e, 5'd5, 27'h0000014d, 5'd19, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002fe, 5'd6, 27'h00000269, 5'd30, 27'h00000202, 32'h00000400,
  1'd1,  5'd9, 27'h0000029c, 5'd19, 27'h0000005b, 5'd7, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000038f, 5'd17, 27'h00000110, 5'd15, 27'h0000031f, 32'h00000400,
  1'd1,  5'd5, 27'h000001ce, 5'd20, 27'h000000a3, 5'd28, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d6, 5'd30, 27'h000003d1, 5'd5, 27'h00000296, 32'h00000400,
  1'd1,  5'd6, 27'h0000036d, 5'd26, 27'h000003da, 5'd17, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003f9, 5'd30, 27'h0000028d, 5'd29, 27'h0000006b, 32'h00000400,
  1'd1,  5'd16, 27'h00000006, 5'd8, 27'h00000030, 5'd6, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000187, 5'd5, 27'h00000257, 5'd19, 27'h000001c3, 32'h00000400,
  1'd1,  5'd16, 27'h0000029a, 5'd8, 27'h000001dd, 5'd26, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000239, 5'd15, 27'h000003f1, 5'd7, 27'h000002bc, 32'h00000400,
  1'd1,  5'd16, 27'h000001e7, 5'd17, 27'h00000307, 5'd19, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000026b, 5'd16, 27'h0000030e, 5'd30, 27'h0000012b, 32'h00000400,
  1'd1,  5'd17, 27'h000000f5, 5'd26, 27'h000002cf, 5'd9, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002ce, 5'd30, 27'h0000004a, 5'd17, 27'h000000ac, 32'h00000400,
  1'd1,  5'd18, 27'h00000208, 5'd26, 27'h000000ca, 5'd27, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000039f, 5'd7, 27'h000000e1, 5'd7, 27'h000003dc, 32'h00000400,
  1'd1,  5'd30, 27'h00000135, 5'd9, 27'h00000150, 5'd16, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000009d, 5'd8, 27'h0000009e, 5'd30, 27'h0000008f, 32'h00000400,
  1'd1,  5'd28, 27'h0000006f, 5'd17, 27'h00000156, 5'd10, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000fb, 5'd17, 27'h000001bd, 5'd19, 27'h000003aa, 32'h00000400,
  1'd1,  5'd25, 27'h0000036c, 5'd19, 27'h00000005, 5'd27, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000266, 5'd28, 27'h000001ef, 5'd8, 27'h000003f9, 32'h00000400,
  1'd1,  5'd27, 27'h000001db, 5'd28, 27'h0000037c, 5'd20, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000296, 5'd29, 27'h00000197, 5'd27, 27'h0000000f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000092, 5'd0, 27'h0000031e, 5'd2, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d3, 5'd1, 27'h0000006d, 5'd15, 27'h00000084, 32'h00000400,
  1'd1,  5'd4, 27'h0000024b, 5'd0, 27'h00000106, 5'd24, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000040, 5'd14, 27'h00000397, 5'd2, 27'h000001eb, 32'h00000400,
  1'd1,  5'd2, 27'h000001d9, 5'd13, 27'h00000269, 5'd12, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000114, 5'd13, 27'h000000fc, 5'd22, 27'h00000214, 32'h00000400,
  1'd1,  5'd3, 27'h000000c4, 5'd22, 27'h0000004b, 5'd3, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000032d, 5'd22, 27'h000002b8, 5'd11, 27'h00000301, 32'h00000400,
  1'd1,  5'd4, 27'h00000049, 5'd24, 27'h0000000e, 5'd25, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000217, 5'd1, 27'h0000010d, 5'd0, 27'h000002e4, 32'h00000400,
  1'd1,  5'd15, 27'h000001ef, 5'd4, 27'h0000023c, 5'd12, 27'h00000400, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000369, 5'd1, 27'h000002de, 5'd23, 27'h000002bb, 32'h00000400,
  1'd1,  5'd12, 27'h000002f2, 5'd14, 27'h0000030a, 5'd4, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003bd, 5'd14, 27'h0000001a, 5'd11, 27'h00000075, 32'h00000400,
  1'd1,  5'd14, 27'h00000391, 5'd10, 27'h0000031e, 5'd23, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000296, 5'd23, 27'h00000179, 5'd2, 27'h00000343, 32'h00000400,
  1'd1,  5'd12, 27'h00000303, 5'd23, 27'h00000211, 5'd13, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000030c, 5'd21, 27'h000001d8, 5'd23, 27'h00000190, 32'h00000400,
  1'd1,  5'd25, 27'h000000de, 5'd4, 27'h0000033a, 5'd3, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000025b, 5'd1, 27'h000002db, 5'd13, 27'h00000362, 32'h00000400,
  1'd1,  5'd23, 27'h000002ce, 5'd1, 27'h00000134, 5'd22, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000123, 5'd15, 27'h0000016f, 5'd1, 27'h00000109, 32'h00000400,
  1'd1,  5'd23, 27'h000001b6, 5'd14, 27'h00000186, 5'd11, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000071, 5'd10, 27'h000003ad, 5'd22, 27'h00000114, 32'h00000400,
  1'd1,  5'd25, 27'h00000034, 5'd20, 27'h0000033c, 5'd4, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000246, 5'd23, 27'h000003ac, 5'd14, 27'h000001f1, 32'h00000400,
  1'd1,  5'd25, 27'h00000102, 5'd20, 27'h000002e7, 5'd24, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000061, 5'd4, 27'h00000263, 5'd8, 27'h00000187, 32'h00000400,
  1'd1,  5'd0, 27'h00000371, 5'd4, 27'h00000367, 5'd20, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000324, 5'd0, 27'h00000182, 5'd27, 27'h00000171, 32'h00000400,
  1'd1,  5'd2, 27'h0000004a, 5'd14, 27'h000002e6, 5'd8, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000205, 5'd13, 27'h00000335, 5'd20, 27'h00000249, 32'h00000400,
  1'd1,  5'd2, 27'h000002a3, 5'd11, 27'h000000ec, 5'd29, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000078, 5'd24, 27'h000001c4, 5'd8, 27'h000000d0, 32'h00000400,
  1'd1,  5'd0, 27'h000000bf, 5'd21, 27'h00000246, 5'd18, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000314, 5'd21, 27'h000002f2, 5'd30, 27'h0000013e, 32'h00000400,
  1'd1,  5'd14, 27'h00000397, 5'd4, 27'h00000125, 5'd5, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000246, 5'd3, 27'h00000116, 5'd17, 27'h00000271, 32'h00000400,
  1'd1,  5'd10, 27'h000003d4, 5'd5, 27'h00000032, 5'd28, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ea, 5'd10, 27'h00000157, 5'd6, 27'h000000cb, 32'h00000400,
  1'd1,  5'd12, 27'h000003e1, 5'd13, 27'h000002ef, 5'd17, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001dd, 5'd13, 27'h00000089, 5'd30, 27'h0000000e, 32'h00000400,
  1'd1,  5'd14, 27'h000001a9, 5'd24, 27'h000001d9, 5'd6, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000013a, 5'd22, 27'h0000015e, 5'd18, 27'h00000187, 32'h00000400,
  1'd1,  5'd12, 27'h00000043, 5'd23, 27'h0000028b, 5'd26, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000332, 5'd4, 27'h0000038f, 5'd9, 27'h000002fa, 32'h00000400,
  1'd1,  5'd25, 27'h00000102, 5'd1, 27'h0000004b, 5'd16, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000274, 5'd4, 27'h000003c5, 5'd28, 27'h000000c2, 32'h00000400,
  1'd1,  5'd23, 27'h000000c6, 5'd14, 27'h00000370, 5'd8, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000363, 5'd14, 27'h00000030, 5'd17, 27'h0000003b, 32'h00000400,
  1'd1,  5'd22, 27'h00000134, 5'd13, 27'h00000330, 5'd26, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002fe, 5'd22, 27'h00000004, 5'd9, 27'h0000033c, 32'h00000400,
  1'd1,  5'd22, 27'h000002b7, 5'd23, 27'h000003be, 5'd19, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000198, 5'd21, 27'h0000001e, 5'd27, 27'h000000bb, 32'h00000400,
  1'd1,  5'd3, 27'h0000004a, 5'd6, 27'h000000f4, 5'd4, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000010b, 5'd6, 27'h000001e7, 5'd11, 27'h00000301, 32'h00000400,
  1'd1,  5'd2, 27'h00000392, 5'd9, 27'h00000012, 5'd23, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d8, 5'd16, 27'h000003c3, 5'd5, 27'h00000035, 32'h00000400,
  1'd1,  5'd3, 27'h0000022a, 5'd17, 27'h000001a7, 5'd15, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000016, 5'd17, 27'h000002c8, 5'd23, 27'h0000027c, 32'h00000400,
  1'd1,  5'd1, 27'h000000e1, 5'd30, 27'h000002d2, 5'd2, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000038, 5'd26, 27'h00000109, 5'd11, 27'h00000244, 32'h00000400,
  1'd1,  5'd1, 27'h0000014b, 5'd28, 27'h000001ac, 5'd23, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000326, 5'd7, 27'h00000305, 5'd4, 27'h00000106, 32'h00000400,
  1'd1,  5'd11, 27'h0000015f, 5'd5, 27'h000000be, 5'd11, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000020d, 5'd7, 27'h0000032d, 5'd23, 27'h0000021c, 32'h00000400,
  1'd1,  5'd12, 27'h000002db, 5'd20, 27'h00000235, 5'd2, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023a, 5'd16, 27'h00000384, 5'd14, 27'h000003c5, 32'h00000400,
  1'd1,  5'd13, 27'h00000229, 5'd20, 27'h000000c2, 5'd21, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000250, 5'd29, 27'h0000002d, 5'd3, 27'h000000f0, 32'h00000400,
  1'd1,  5'd10, 27'h00000380, 5'd30, 27'h00000369, 5'd11, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000170, 5'd30, 27'h000001b7, 5'd25, 27'h0000003e, 32'h00000400,
  1'd1,  5'd25, 27'h000002fc, 5'd6, 27'h0000011a, 5'd1, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e2, 5'd5, 27'h00000101, 5'd11, 27'h00000191, 32'h00000400,
  1'd1,  5'd20, 27'h0000037d, 5'd10, 27'h00000104, 5'd21, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002db, 5'd17, 27'h0000029d, 5'd5, 27'h0000002c, 32'h00000400,
  1'd1,  5'd24, 27'h000000e4, 5'd20, 27'h000000ec, 5'd11, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000030a, 5'd16, 27'h000000a7, 5'd24, 27'h0000008a, 32'h00000400,
  1'd1,  5'd25, 27'h00000231, 5'd26, 27'h000000b9, 5'd4, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001f3, 5'd27, 27'h00000058, 5'd10, 27'h000002a0, 32'h00000400,
  1'd1,  5'd23, 27'h00000388, 5'd30, 27'h000003ab, 5'd23, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000287, 5'd6, 27'h0000026c, 5'd9, 27'h0000023d, 32'h00000400,
  1'd1,  5'd1, 27'h0000027c, 5'd8, 27'h0000005d, 5'd17, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000400, 5'd6, 27'h0000011c, 5'd28, 27'h00000006, 32'h00000400,
  1'd1,  5'd3, 27'h000001a2, 5'd20, 27'h00000187, 5'd9, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000032d, 5'd20, 27'h0000018a, 5'd16, 27'h0000004a, 32'h00000400,
  1'd1,  5'd4, 27'h00000221, 5'd17, 27'h000001a5, 5'd27, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000060, 5'd27, 27'h00000225, 5'd10, 27'h00000019, 32'h00000400,
  1'd1,  5'd1, 27'h000002f0, 5'd28, 27'h000001d4, 5'd18, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002de, 5'd29, 27'h000001f9, 5'd29, 27'h0000013e, 32'h00000400,
  1'd1,  5'd10, 27'h000003ac, 5'd10, 27'h00000073, 5'd6, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001f6, 5'd6, 27'h000003a8, 5'd17, 27'h00000261, 32'h00000400,
  1'd1,  5'd11, 27'h00000102, 5'd9, 27'h0000017e, 5'd29, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000034c, 5'd18, 27'h00000321, 5'd7, 27'h000000af, 32'h00000400,
  1'd1,  5'd11, 27'h0000017f, 5'd16, 27'h0000007b, 5'd15, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000025b, 5'd15, 27'h000002ed, 5'd29, 27'h00000238, 32'h00000400,
  1'd1,  5'd13, 27'h000001d3, 5'd30, 27'h0000027c, 5'd9, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000049, 5'd27, 27'h0000030b, 5'd16, 27'h000002a6, 32'h00000400,
  1'd1,  5'd15, 27'h0000018f, 5'd29, 27'h000001d6, 5'd29, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000199, 5'd7, 27'h0000002f, 5'd9, 27'h00000272, 32'h00000400,
  1'd1,  5'd20, 27'h000002b5, 5'd6, 27'h0000032c, 5'd16, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000147, 5'd5, 27'h00000119, 5'd29, 27'h000001ab, 32'h00000400,
  1'd1,  5'd21, 27'h0000029b, 5'd16, 27'h0000003f, 5'd6, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000027, 5'd17, 27'h000002c6, 5'd16, 27'h00000136, 32'h00000400,
  1'd1,  5'd21, 27'h000003e4, 5'd19, 27'h00000188, 5'd26, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000100, 5'd29, 27'h00000352, 5'd7, 27'h00000025, 32'h00000400,
  1'd1,  5'd24, 27'h000003e9, 5'd27, 27'h00000126, 5'd18, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000228, 5'd26, 27'h000002a2, 5'd30, 27'h0000027a, 32'h00000400,
  1'd1,  5'd6, 27'h000002d2, 5'd0, 27'h000000cc, 5'd5, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000a9, 5'd3, 27'h00000140, 5'd15, 27'h0000021f, 32'h00000400,
  1'd1,  5'd6, 27'h00000156, 5'd4, 27'h0000008b, 5'd27, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000004c, 5'd10, 27'h0000026d, 5'd2, 27'h00000138, 32'h00000400,
  1'd1,  5'd5, 27'h00000368, 5'd14, 27'h0000009d, 5'd13, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003dc, 5'd12, 27'h000002b0, 5'd24, 27'h0000022e, 32'h00000400,
  1'd1,  5'd8, 27'h00000190, 5'd24, 27'h000000f5, 5'd3, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cf, 5'd20, 27'h000003c7, 5'd12, 27'h000000a8, 32'h00000400,
  1'd1,  5'd7, 27'h000000b3, 5'd23, 27'h00000098, 5'd23, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001a8, 5'd1, 27'h000003ce, 5'd9, 27'h00000123, 32'h00000400,
  1'd1,  5'd16, 27'h00000030, 5'd4, 27'h000002f6, 5'd16, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000086, 5'd3, 27'h0000026b, 5'd28, 27'h000001d3, 32'h00000400,
  1'd1,  5'd16, 27'h000002cc, 5'd14, 27'h00000387, 5'd2, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000db, 5'd11, 27'h00000325, 5'd11, 27'h000003e0, 32'h00000400,
  1'd1,  5'd18, 27'h000000d0, 5'd14, 27'h0000007f, 5'd25, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ad, 5'd23, 27'h00000086, 5'd4, 27'h000002c7, 32'h00000400,
  1'd1,  5'd18, 27'h00000277, 5'd24, 27'h0000030d, 5'd10, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000010a, 5'd21, 27'h000002fe, 5'd23, 27'h00000226, 32'h00000400,
  1'd1,  5'd27, 27'h0000017a, 5'd1, 27'h000001a0, 5'd0, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003c5, 5'd2, 27'h00000030, 5'd12, 27'h000002cf, 32'h00000400,
  1'd1,  5'd26, 27'h000001a7, 5'd4, 27'h000000bf, 5'd23, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d0, 5'd14, 27'h0000013e, 5'd2, 27'h000001b3, 32'h00000400,
  1'd1,  5'd28, 27'h000001fb, 5'd11, 27'h000003f0, 5'd13, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000216, 5'd13, 27'h0000027a, 5'd25, 27'h0000009e, 32'h00000400,
  1'd1,  5'd27, 27'h000003fb, 5'd25, 27'h00000071, 5'd0, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000165, 5'd25, 27'h00000214, 5'd10, 27'h00000256, 32'h00000400,
  1'd1,  5'd28, 27'h000003d3, 5'd24, 27'h00000323, 5'd24, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002e7, 5'd4, 27'h000003ca, 5'd3, 27'h000003c3, 32'h00000400,
  1'd1,  5'd7, 27'h00000083, 5'd0, 27'h0000035c, 5'd10, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000301, 5'd5, 27'h00000029, 5'd21, 27'h00000019, 32'h00000400,
  1'd1,  5'd6, 27'h0000029b, 5'd13, 27'h0000027f, 5'd5, 27'h00000169, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000255, 5'd12, 27'h00000182, 5'd16, 27'h00000384, 32'h00000400,
  1'd1,  5'd8, 27'h00000228, 5'd11, 27'h00000148, 5'd30, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fc, 5'd24, 27'h00000326, 5'd7, 27'h000003d6, 32'h00000400,
  1'd1,  5'd10, 27'h0000005e, 5'd24, 27'h0000010c, 5'd16, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003a7, 5'd22, 27'h0000029d, 5'd27, 27'h000002fa, 32'h00000400,
  1'd1,  5'd17, 27'h00000379, 5'd0, 27'h00000065, 5'd1, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003bb, 5'd2, 27'h00000083, 5'd12, 27'h0000024c, 32'h00000400,
  1'd1,  5'd18, 27'h00000338, 5'd3, 27'h000001f2, 5'd21, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000272, 5'd14, 27'h00000326, 5'd8, 27'h00000040, 32'h00000400,
  1'd1,  5'd19, 27'h000003dc, 5'd12, 27'h00000252, 5'd18, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000036f, 5'd10, 27'h000003ed, 5'd28, 27'h00000113, 32'h00000400,
  1'd1,  5'd16, 27'h000002c3, 5'd24, 27'h00000196, 5'd6, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ce, 5'd21, 27'h000003af, 5'd17, 27'h0000029c, 32'h00000400,
  1'd1,  5'd18, 27'h000001c9, 5'd21, 27'h00000152, 5'd30, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d6, 5'd2, 27'h000001d6, 5'd5, 27'h00000372, 32'h00000400,
  1'd1,  5'd27, 27'h00000190, 5'd4, 27'h00000236, 5'd17, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002e2, 5'd2, 27'h0000033d, 5'd26, 27'h000003fe, 32'h00000400,
  1'd1,  5'd29, 27'h0000031c, 5'd14, 27'h000002b8, 5'd8, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000206, 5'd14, 27'h000003b6, 5'd19, 27'h00000236, 32'h00000400,
  1'd1,  5'd26, 27'h00000199, 5'd11, 27'h00000357, 5'd30, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000133, 5'd23, 27'h00000383, 5'd7, 27'h00000349, 32'h00000400,
  1'd1,  5'd25, 27'h000003c8, 5'd20, 27'h0000033b, 5'd18, 27'h0000001c, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001db, 5'd23, 27'h00000174, 5'd28, 27'h0000010b, 32'h00000400,
  1'd1,  5'd9, 27'h000002d1, 5'd6, 27'h00000176, 5'd5, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000029, 5'd9, 27'h00000076, 5'd14, 27'h00000217, 32'h00000400,
  1'd1,  5'd5, 27'h0000039b, 5'd8, 27'h000000f9, 5'd24, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038c, 5'd20, 27'h000000b2, 5'd0, 27'h00000198, 32'h00000400,
  1'd1,  5'd7, 27'h0000002e, 5'd15, 27'h0000026b, 5'd14, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000291, 5'd20, 27'h00000208, 5'd21, 27'h000003df, 32'h00000400,
  1'd1,  5'd7, 27'h00000005, 5'd28, 27'h00000331, 5'd3, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000210, 5'd27, 27'h00000017, 5'd11, 27'h0000038d, 32'h00000400,
  1'd1,  5'd7, 27'h00000301, 5'd29, 27'h000000d3, 5'd24, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000b0, 5'd7, 27'h000000ec, 5'd4, 27'h0000023a, 32'h00000400,
  1'd1,  5'd16, 27'h00000011, 5'd5, 27'h000001ba, 5'd12, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000293, 5'd7, 27'h00000170, 5'd23, 27'h00000328, 32'h00000400,
  1'd1,  5'd19, 27'h000000c3, 5'd20, 27'h00000066, 5'd2, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000025e, 5'd17, 27'h000002b5, 5'd12, 27'h000001a2, 32'h00000400,
  1'd1,  5'd20, 27'h000002aa, 5'd19, 27'h0000033d, 5'd21, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000018d, 5'd29, 27'h00000188, 5'd2, 27'h00000213, 32'h00000400,
  1'd1,  5'd20, 27'h0000006d, 5'd28, 27'h000003a5, 5'd14, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002dd, 5'd30, 27'h0000015e, 5'd24, 27'h0000035a, 32'h00000400,
  1'd1,  5'd26, 27'h00000329, 5'd6, 27'h00000219, 5'd1, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a0, 5'd10, 27'h00000042, 5'd11, 27'h000000e3, 32'h00000400,
  1'd1,  5'd27, 27'h00000087, 5'd6, 27'h000001b6, 5'd25, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000f7, 5'd19, 27'h000002a6, 5'd2, 27'h00000037, 32'h00000400,
  1'd1,  5'd30, 27'h0000004e, 5'd17, 27'h000001b0, 5'd13, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000029c, 5'd16, 27'h000003ae, 5'd24, 27'h0000019d, 32'h00000400,
  1'd1,  5'd26, 27'h0000000b, 5'd30, 27'h0000022b, 5'd4, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000018f, 5'd30, 27'h000003ae, 5'd10, 27'h000001fd, 32'h00000400,
  1'd1,  5'd29, 27'h0000020d, 5'd30, 27'h00000371, 5'd22, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001db, 5'd9, 27'h000002cf, 5'd6, 27'h000003ed, 32'h00000400,
  1'd1,  5'd6, 27'h000000cc, 5'd10, 27'h00000112, 5'd19, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000019c, 5'd9, 27'h000000f9, 5'd26, 27'h000002e2, 32'h00000400,
  1'd1,  5'd6, 27'h00000039, 5'd16, 27'h0000007c, 5'd9, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d5, 5'd16, 27'h0000037a, 5'd19, 27'h000003ad, 32'h00000400,
  1'd1,  5'd9, 27'h00000321, 5'd17, 27'h000002ea, 5'd30, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000283, 5'd26, 27'h0000004d, 5'd5, 27'h0000029a, 32'h00000400,
  1'd1,  5'd7, 27'h0000033a, 5'd29, 27'h00000283, 5'd17, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003f9, 5'd26, 27'h00000033, 5'd27, 27'h00000304, 32'h00000400,
  1'd1,  5'd18, 27'h0000002b, 5'd6, 27'h0000030f, 5'd7, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000258, 5'd10, 27'h00000079, 5'd19, 27'h000001bd, 32'h00000400,
  1'd1,  5'd19, 27'h00000299, 5'd8, 27'h0000026c, 5'd28, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000020, 5'd16, 27'h00000099, 5'd9, 27'h00000283, 32'h00000400,
  1'd1,  5'd16, 27'h00000140, 5'd16, 27'h00000096, 5'd16, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001bc, 5'd17, 27'h00000355, 5'd30, 27'h0000012f, 32'h00000400,
  1'd1,  5'd16, 27'h000000b3, 5'd27, 27'h000000bc, 5'd9, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000028d, 5'd30, 27'h000002c6, 5'd17, 27'h0000037b, 32'h00000400,
  1'd1,  5'd17, 27'h00000253, 5'd28, 27'h0000005b, 5'd28, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000287, 5'd9, 27'h0000019f, 5'd8, 27'h00000326, 32'h00000400,
  1'd1,  5'd28, 27'h00000199, 5'd8, 27'h00000155, 5'd17, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f9, 5'd9, 27'h00000123, 5'd29, 27'h00000037, 32'h00000400,
  1'd1,  5'd29, 27'h000001bf, 5'd16, 27'h00000188, 5'd5, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000357, 5'd20, 27'h00000279, 5'd18, 27'h00000002, 32'h00000400,
  1'd1,  5'd30, 27'h00000113, 5'd16, 27'h0000032b, 5'd27, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000069, 5'd30, 27'h0000006a, 5'd7, 27'h000001aa, 32'h00000400,
  1'd1,  5'd27, 27'h000003f2, 5'd26, 27'h00000130, 5'd19, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001fb, 5'd27, 27'h0000025a, 5'd28, 27'h00000304, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000000e1, 5'd4, 27'h0000006b, 5'd4, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000317, 5'd4, 27'h0000020d, 5'd11, 27'h00000003, 32'h00000400,
  1'd1,  5'd2, 27'h00000095, 5'd2, 27'h000002f8, 5'd24, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000005d, 5'd15, 27'h000001e7, 5'd2, 27'h000003db, 32'h00000400,
  1'd1,  5'd1, 27'h00000059, 5'd11, 27'h000001fa, 5'd14, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000028, 5'd12, 27'h000001f5, 5'd24, 27'h000001b7, 32'h00000400,
  1'd1,  5'd2, 27'h00000042, 5'd23, 27'h000001cc, 5'd4, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003b8, 5'd22, 27'h00000366, 5'd11, 27'h000001e4, 32'h00000400,
  1'd1,  5'd3, 27'h00000395, 5'd22, 27'h00000194, 5'd23, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001e8, 5'd0, 27'h000001fa, 5'd2, 27'h000000e6, 32'h00000400,
  1'd1,  5'd14, 27'h00000116, 5'd0, 27'h00000196, 5'd14, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000013b, 5'd3, 27'h0000013f, 5'd20, 27'h0000033d, 32'h00000400,
  1'd1,  5'd11, 27'h000003ad, 5'd13, 27'h00000218, 5'd0, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c5, 5'd12, 27'h000003c4, 5'd12, 27'h000002af, 32'h00000400,
  1'd1,  5'd15, 27'h000000ae, 5'd11, 27'h00000372, 5'd25, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000367, 5'd21, 27'h0000014e, 5'd0, 27'h000000f7, 32'h00000400,
  1'd1,  5'd15, 27'h000001e2, 5'd21, 27'h000003a2, 5'd14, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000031, 5'd21, 27'h00000090, 5'd24, 27'h000001c2, 32'h00000400,
  1'd1,  5'd21, 27'h00000057, 5'd2, 27'h0000035a, 5'd0, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003be, 5'd4, 27'h000001d0, 5'd11, 27'h0000038a, 32'h00000400,
  1'd1,  5'd24, 27'h000003d4, 5'd1, 27'h00000288, 5'd21, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000265, 5'd12, 27'h00000098, 5'd3, 27'h0000012b, 32'h00000400,
  1'd1,  5'd24, 27'h000000a3, 5'd13, 27'h0000025f, 5'd14, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000008e, 5'd11, 27'h00000345, 5'd21, 27'h00000164, 32'h00000400,
  1'd1,  5'd23, 27'h000001e2, 5'd24, 27'h000002df, 5'd1, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001e8, 5'd21, 27'h000001d1, 5'd10, 27'h000001f5, 32'h00000400,
  1'd1,  5'd24, 27'h000000ef, 5'd23, 27'h000003d8, 5'd24, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000009c, 5'd3, 27'h00000208, 5'd5, 27'h00000202, 32'h00000400,
  1'd1,  5'd2, 27'h0000021b, 5'd4, 27'h00000278, 5'd19, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e3, 5'd2, 27'h0000027d, 5'd30, 27'h0000037f, 32'h00000400,
  1'd1,  5'd4, 27'h0000039f, 5'd10, 27'h000003c2, 5'd6, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028a, 5'd14, 27'h000002ff, 5'd16, 27'h0000030c, 32'h00000400,
  1'd1,  5'd0, 27'h000001ff, 5'd12, 27'h00000296, 5'd28, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000028c, 5'd22, 27'h0000012d, 5'd8, 27'h0000006d, 32'h00000400,
  1'd1,  5'd4, 27'h00000226, 5'd25, 27'h000000fd, 5'd17, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029f, 5'd24, 27'h000001db, 5'd26, 27'h000000d9, 32'h00000400,
  1'd1,  5'd14, 27'h0000008e, 5'd5, 27'h00000014, 5'd6, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003e6, 5'd2, 27'h00000233, 5'd16, 27'h000001d3, 32'h00000400,
  1'd1,  5'd11, 27'h000002cd, 5'd2, 27'h00000108, 5'd29, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000007, 5'd11, 27'h000001a6, 5'd9, 27'h0000030b, 32'h00000400,
  1'd1,  5'd15, 27'h00000016, 5'd11, 27'h0000000c, 5'd15, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000359, 5'd13, 27'h00000337, 5'd28, 27'h000000dc, 32'h00000400,
  1'd1,  5'd10, 27'h000003a5, 5'd23, 27'h000003bb, 5'd10, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000377, 5'd23, 27'h0000022f, 5'd18, 27'h000003ac, 32'h00000400,
  1'd1,  5'd10, 27'h000002c7, 5'd24, 27'h0000019e, 5'd28, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000032e, 5'd1, 27'h00000253, 5'd6, 27'h000001b8, 32'h00000400,
  1'd1,  5'd21, 27'h00000355, 5'd2, 27'h000001fe, 5'd16, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022f, 5'd2, 27'h00000276, 5'd25, 27'h000003b8, 32'h00000400,
  1'd1,  5'd21, 27'h00000121, 5'd14, 27'h00000170, 5'd6, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000376, 5'd12, 27'h0000003e, 5'd17, 27'h000000d8, 32'h00000400,
  1'd1,  5'd22, 27'h00000260, 5'd14, 27'h000002a8, 5'd25, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000299, 5'd23, 27'h000002d8, 5'd6, 27'h00000323, 32'h00000400,
  1'd1,  5'd21, 27'h00000015, 5'd24, 27'h000002e4, 5'd16, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e4, 5'd22, 27'h000001bf, 5'd26, 27'h00000180, 32'h00000400,
  1'd1,  5'd0, 27'h00000312, 5'd6, 27'h000000fc, 5'd2, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ac, 5'd7, 27'h000001c1, 5'd12, 27'h000001e6, 32'h00000400,
  1'd1,  5'd2, 27'h0000004a, 5'd7, 27'h0000000e, 5'd24, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000061, 5'd17, 27'h0000023b, 5'd3, 27'h0000017f, 32'h00000400,
  1'd1,  5'd3, 27'h0000029a, 5'd19, 27'h00000383, 5'd12, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000212, 5'd17, 27'h000001f3, 5'd22, 27'h0000020b, 32'h00000400,
  1'd1,  5'd4, 27'h0000007b, 5'd29, 27'h00000396, 5'd2, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001bd, 5'd30, 27'h0000028a, 5'd15, 27'h000001a1, 32'h00000400,
  1'd1,  5'd1, 27'h000002b6, 5'd27, 27'h000000c0, 5'd20, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b4, 5'd9, 27'h000000fa, 5'd1, 27'h00000157, 32'h00000400,
  1'd1,  5'd10, 27'h000002b6, 5'd5, 27'h000000b2, 5'd14, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c9, 5'd9, 27'h0000024c, 5'd23, 27'h0000011b, 32'h00000400,
  1'd1,  5'd14, 27'h00000349, 5'd18, 27'h000001e3, 5'd3, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003bd, 5'd18, 27'h0000016f, 5'd14, 27'h000000dd, 32'h00000400,
  1'd1,  5'd13, 27'h00000059, 5'd18, 27'h000003c4, 5'd23, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000011, 5'd28, 27'h00000284, 5'd4, 27'h000003ca, 32'h00000400,
  1'd1,  5'd12, 27'h00000242, 5'd27, 27'h00000233, 5'd14, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000366, 5'd28, 27'h000000e8, 5'd23, 27'h000002ff, 32'h00000400,
  1'd1,  5'd25, 27'h0000015d, 5'd7, 27'h0000009e, 5'd3, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000394, 5'd9, 27'h00000344, 5'd10, 27'h000001ee, 32'h00000400,
  1'd1,  5'd23, 27'h0000015f, 5'd9, 27'h00000077, 5'd21, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ab, 5'd16, 27'h000001ec, 5'd0, 27'h00000024, 32'h00000400,
  1'd1,  5'd21, 27'h000000f3, 5'd16, 27'h00000195, 5'd10, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000167, 5'd18, 27'h000000d2, 5'd23, 27'h000003a2, 32'h00000400,
  1'd1,  5'd21, 27'h00000208, 5'd30, 27'h000003c6, 5'd0, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000253, 5'd30, 27'h00000174, 5'd15, 27'h00000158, 32'h00000400,
  1'd1,  5'd21, 27'h000001b5, 5'd30, 27'h000001cf, 5'd21, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000007d, 5'd9, 27'h0000035b, 5'd7, 27'h000003cf, 32'h00000400,
  1'd1,  5'd3, 27'h00000336, 5'd8, 27'h0000035c, 5'd19, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000083, 5'd9, 27'h00000046, 5'd26, 27'h000002ed, 32'h00000400,
  1'd1,  5'd2, 27'h00000120, 5'd16, 27'h00000322, 5'd8, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ea, 5'd18, 27'h000002d6, 5'd15, 27'h00000376, 32'h00000400,
  1'd1,  5'd3, 27'h00000377, 5'd16, 27'h00000215, 5'd27, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000211, 5'd30, 27'h000000d8, 5'd8, 27'h000003d4, 32'h00000400,
  1'd1,  5'd3, 27'h000001c6, 5'd29, 27'h000001e3, 5'd19, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000330, 5'd29, 27'h00000110, 5'd29, 27'h00000130, 32'h00000400,
  1'd1,  5'd13, 27'h0000001e, 5'd6, 27'h000000df, 5'd9, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002c1, 5'd9, 27'h00000016, 5'd18, 27'h00000263, 32'h00000400,
  1'd1,  5'd12, 27'h00000214, 5'd8, 27'h000000f6, 5'd30, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001b1, 5'd18, 27'h00000175, 5'd5, 27'h000003c8, 32'h00000400,
  1'd1,  5'd10, 27'h000002c1, 5'd15, 27'h0000021c, 5'd19, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c5, 5'd16, 27'h00000031, 5'd29, 27'h000003d9, 32'h00000400,
  1'd1,  5'd13, 27'h0000006a, 5'd28, 27'h0000004f, 5'd6, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000bc, 5'd28, 27'h00000050, 5'd20, 27'h00000228, 32'h00000400,
  1'd1,  5'd13, 27'h00000220, 5'd29, 27'h000000bf, 5'd29, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000069, 5'd8, 27'h000002e8, 5'd6, 27'h00000367, 32'h00000400,
  1'd1,  5'd21, 27'h00000353, 5'd7, 27'h000002ba, 5'd15, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000007c, 5'd6, 27'h00000039, 5'd26, 27'h000000e7, 32'h00000400,
  1'd1,  5'd25, 27'h00000170, 5'd19, 27'h00000299, 5'd5, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000010f, 5'd19, 27'h00000088, 5'd18, 27'h000002f4, 32'h00000400,
  1'd1,  5'd21, 27'h0000039b, 5'd20, 27'h00000053, 5'd27, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000347, 5'd30, 27'h00000112, 5'd7, 27'h000002ce, 32'h00000400,
  1'd1,  5'd24, 27'h000002b6, 5'd26, 27'h00000153, 5'd17, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000024f, 5'd30, 27'h0000010a, 5'd29, 27'h0000033b, 32'h00000400,
  1'd1,  5'd7, 27'h0000006d, 5'd1, 27'h000003e6, 5'd7, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000214, 5'd4, 27'h0000029a, 5'd19, 27'h00000023, 32'h00000400,
  1'd1,  5'd5, 27'h000000de, 5'd0, 27'h0000027d, 5'd27, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000b7, 5'd12, 27'h000000b1, 5'd2, 27'h0000017b, 32'h00000400,
  1'd1,  5'd10, 27'h0000002e, 5'd10, 27'h000001b7, 5'd13, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000037a, 5'd14, 27'h000001de, 5'd20, 27'h000003ed, 32'h00000400,
  1'd1,  5'd6, 27'h000000fb, 5'd25, 27'h000000d5, 5'd1, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000c5, 5'd24, 27'h00000122, 5'd13, 27'h000001d0, 32'h00000400,
  1'd1,  5'd5, 27'h000002aa, 5'd21, 27'h00000144, 5'd21, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000013c, 5'd2, 27'h00000251, 5'd5, 27'h00000165, 32'h00000400,
  1'd1,  5'd17, 27'h0000030d, 5'd4, 27'h000002a0, 5'd18, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000154, 5'd0, 27'h000002ff, 5'd29, 27'h00000261, 32'h00000400,
  1'd1,  5'd19, 27'h00000223, 5'd14, 27'h0000022a, 5'd0, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000024b, 5'd15, 27'h00000122, 5'd12, 27'h000002ff, 32'h00000400,
  1'd1,  5'd17, 27'h0000032d, 5'd15, 27'h00000029, 5'd20, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c7, 5'd23, 27'h000002aa, 5'd2, 27'h00000098, 32'h00000400,
  1'd1,  5'd16, 27'h000000c6, 5'd25, 27'h00000290, 5'd11, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000009b, 5'd25, 27'h00000030, 5'd21, 27'h0000035c, 32'h00000400,
  1'd1,  5'd29, 27'h000002d3, 5'd2, 27'h000001e5, 5'd3, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000294, 5'd4, 27'h0000039c, 5'd13, 27'h000003d8, 32'h00000400,
  1'd1,  5'd28, 27'h000003e5, 5'd1, 27'h0000013a, 5'd21, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000282, 5'd12, 27'h000001c4, 5'd1, 27'h000002e7, 32'h00000400,
  1'd1,  5'd27, 27'h0000034f, 5'd13, 27'h000001bc, 5'd11, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000192, 5'd10, 27'h0000018d, 5'd21, 27'h00000006, 32'h00000400,
  1'd1,  5'd27, 27'h00000323, 5'd23, 27'h000002d4, 5'd3, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002cb, 5'd21, 27'h000000c3, 5'd14, 27'h000003cf, 32'h00000400,
  1'd1,  5'd26, 27'h000000d4, 5'd22, 27'h00000226, 5'd25, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c5, 5'd4, 27'h00000246, 5'd0, 27'h00000102, 32'h00000400,
  1'd1,  5'd5, 27'h000003b4, 5'd2, 27'h00000094, 5'd13, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000016c, 5'd3, 27'h0000006d, 5'd22, 27'h00000305, 32'h00000400,
  1'd1,  5'd5, 27'h000000c4, 5'd10, 27'h000001d8, 5'd8, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000327, 5'd10, 27'h000001be, 5'd19, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h00000092, 5'd13, 27'h00000016, 5'd26, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000178, 5'd23, 27'h00000120, 5'd9, 27'h000003d0, 32'h00000400,
  1'd1,  5'd8, 27'h00000105, 5'd24, 27'h0000028e, 5'd17, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000073, 5'd21, 27'h00000037, 5'd30, 27'h00000295, 32'h00000400,
  1'd1,  5'd16, 27'h000001e4, 5'd1, 27'h0000002b, 5'd0, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000021, 5'd3, 27'h000002f3, 5'd11, 27'h00000108, 32'h00000400,
  1'd1,  5'd15, 27'h00000237, 5'd1, 27'h0000006b, 5'd22, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a1, 5'd10, 27'h00000227, 5'd9, 27'h000003d5, 32'h00000400,
  1'd1,  5'd19, 27'h00000206, 5'd12, 27'h000001d6, 5'd16, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000397, 5'd13, 27'h000003d9, 5'd27, 27'h000001c6, 32'h00000400,
  1'd1,  5'd17, 27'h0000029e, 5'd24, 27'h0000038a, 5'd6, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000191, 5'd23, 27'h000003f8, 5'd17, 27'h00000218, 32'h00000400,
  1'd1,  5'd19, 27'h000003d9, 5'd22, 27'h0000004b, 5'd28, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b7, 5'd3, 27'h000001d2, 5'd7, 27'h0000005d, 32'h00000400,
  1'd1,  5'd28, 27'h00000242, 5'd4, 27'h0000022c, 5'd19, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000091, 5'd1, 27'h000003c1, 5'd29, 27'h00000235, 32'h00000400,
  1'd1,  5'd30, 27'h000002a4, 5'd11, 27'h0000037c, 5'd10, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a0, 5'd10, 27'h0000027e, 5'd19, 27'h00000252, 32'h00000400,
  1'd1,  5'd30, 27'h000003a0, 5'd13, 27'h00000293, 5'd29, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000210, 5'd23, 27'h000001e2, 5'd9, 27'h000000a4, 32'h00000400,
  1'd1,  5'd30, 27'h000002f1, 5'd22, 27'h0000001d, 5'd15, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000041, 5'd20, 27'h00000390, 5'd28, 27'h0000020a, 32'h00000400,
  1'd1,  5'd9, 27'h0000000f, 5'd10, 27'h00000015, 5'd0, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c4, 5'd9, 27'h000001b5, 5'd10, 27'h000001a2, 32'h00000400,
  1'd1,  5'd9, 27'h000002ed, 5'd7, 27'h00000083, 5'd22, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000100, 5'd17, 27'h0000025c, 5'd2, 27'h000002ce, 32'h00000400,
  1'd1,  5'd6, 27'h0000000f, 5'd19, 27'h00000340, 5'd11, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002ae, 5'd17, 27'h00000244, 5'd22, 27'h00000128, 32'h00000400,
  1'd1,  5'd9, 27'h00000011, 5'd30, 27'h00000180, 5'd2, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000018e, 5'd27, 27'h000002c1, 5'd13, 27'h00000210, 32'h00000400,
  1'd1,  5'd10, 27'h00000057, 5'd29, 27'h000001ac, 5'd21, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000189, 5'd9, 27'h0000012a, 5'd2, 27'h00000113, 32'h00000400,
  1'd1,  5'd15, 27'h00000256, 5'd10, 27'h000000ed, 5'd12, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ae, 5'd9, 27'h0000022f, 5'd20, 27'h000002c9, 32'h00000400,
  1'd1,  5'd17, 27'h00000021, 5'd16, 27'h0000023d, 5'd1, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000065, 5'd16, 27'h000001b5, 5'd11, 27'h000003b9, 32'h00000400,
  1'd1,  5'd16, 27'h00000350, 5'd19, 27'h000002cc, 5'd20, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000004a, 5'd27, 27'h00000081, 5'd4, 27'h000003c1, 32'h00000400,
  1'd1,  5'd16, 27'h00000270, 5'd28, 27'h000001ba, 5'd12, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000008c, 5'd29, 27'h000001ae, 5'd25, 27'h000000e0, 32'h00000400,
  1'd1,  5'd27, 27'h00000113, 5'd9, 27'h0000025c, 5'd3, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000023a, 5'd8, 27'h0000010d, 5'd11, 27'h000000b7, 32'h00000400,
  1'd1,  5'd27, 27'h0000009c, 5'd9, 27'h00000092, 5'd23, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000008c, 5'd17, 27'h00000077, 5'd1, 27'h00000167, 32'h00000400,
  1'd1,  5'd30, 27'h000003d6, 5'd15, 27'h000003a5, 5'd11, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000d8, 5'd16, 27'h0000010a, 5'd25, 27'h0000023d, 32'h00000400,
  1'd1,  5'd26, 27'h000002b8, 5'd30, 27'h0000001c, 5'd3, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000358, 5'd26, 27'h000003c0, 5'd10, 27'h0000027f, 32'h00000400,
  1'd1,  5'd28, 27'h00000181, 5'd29, 27'h0000021e, 5'd22, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000035f, 5'd5, 27'h000000b2, 5'd7, 27'h00000075, 32'h00000400,
  1'd1,  5'd8, 27'h0000036e, 5'd6, 27'h0000031a, 5'd16, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000094, 5'd7, 27'h000003b6, 5'd29, 27'h00000104, 32'h00000400,
  1'd1,  5'd9, 27'h00000058, 5'd16, 27'h00000315, 5'd5, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000151, 5'd17, 27'h00000076, 5'd19, 27'h00000158, 32'h00000400,
  1'd1,  5'd6, 27'h00000333, 5'd20, 27'h00000211, 5'd30, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000000c, 5'd26, 27'h000001c2, 5'd8, 27'h00000373, 32'h00000400,
  1'd1,  5'd9, 27'h0000024b, 5'd26, 27'h000002f5, 5'd19, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000198, 5'd27, 27'h000002ae, 5'd27, 27'h0000038a, 32'h00000400,
  1'd1,  5'd15, 27'h00000379, 5'd6, 27'h000000a7, 5'd7, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000261, 5'd7, 27'h000003dd, 5'd15, 27'h00000338, 32'h00000400,
  1'd1,  5'd17, 27'h000003ae, 5'd8, 27'h0000014a, 5'd30, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002b, 5'd19, 27'h00000338, 5'd5, 27'h0000037c, 32'h00000400,
  1'd1,  5'd17, 27'h000002cd, 5'd16, 27'h00000014, 5'd19, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d5, 5'd16, 27'h00000302, 5'd29, 27'h00000197, 32'h00000400,
  1'd1,  5'd20, 27'h0000000d, 5'd29, 27'h000001f3, 5'd5, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000043, 5'd29, 27'h00000170, 5'd17, 27'h00000117, 32'h00000400,
  1'd1,  5'd15, 27'h0000020c, 5'd28, 27'h0000012f, 5'd30, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f0, 5'd9, 27'h000003c8, 5'd8, 27'h00000362, 32'h00000400,
  1'd1,  5'd30, 27'h00000360, 5'd7, 27'h00000382, 5'd17, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000020f, 5'd7, 27'h000000ed, 5'd30, 27'h000000a4, 32'h00000400,
  1'd1,  5'd30, 27'h0000003e, 5'd18, 27'h00000104, 5'd8, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000320, 5'd18, 27'h00000370, 5'd19, 27'h00000026, 32'h00000400,
  1'd1,  5'd28, 27'h00000212, 5'd19, 27'h0000032f, 5'd28, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003e4, 5'd26, 27'h000001a2, 5'd6, 27'h0000000e, 32'h00000400,
  1'd1,  5'd28, 27'h000003c9, 5'd30, 27'h00000318, 5'd17, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f6, 5'd28, 27'h000001a5, 5'd27, 27'h0000037d, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000171, 5'd1, 27'h00000313, 5'd1, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003da, 5'd0, 27'h0000023f, 5'd10, 27'h0000021e, 32'h00000400,
  1'd1,  5'd2, 27'h00000361, 5'd3, 27'h00000144, 5'd22, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e3, 5'd13, 27'h00000224, 5'd0, 27'h000000e8, 32'h00000400,
  1'd1,  5'd4, 27'h00000202, 5'd14, 27'h0000025f, 5'd15, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002ec, 5'd14, 27'h0000027f, 5'd22, 27'h000000cc, 32'h00000400,
  1'd1,  5'd4, 27'h000000d7, 5'd21, 27'h000002b1, 5'd3, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002a6, 5'd24, 27'h0000010e, 5'd12, 27'h00000090, 32'h00000400,
  1'd1,  5'd0, 27'h000000ef, 5'd23, 27'h00000017, 5'd25, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000016d, 5'd0, 27'h000001d6, 5'd5, 27'h00000007, 32'h00000400,
  1'd1,  5'd11, 27'h00000026, 5'd3, 27'h0000008a, 5'd10, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000010f, 5'd2, 27'h00000326, 5'd22, 27'h000002f2, 32'h00000400,
  1'd1,  5'd12, 27'h0000020a, 5'd11, 27'h00000237, 5'd4, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000016a, 5'd15, 27'h0000013f, 5'd11, 27'h000000cf, 32'h00000400,
  1'd1,  5'd11, 27'h00000149, 5'd13, 27'h000001a1, 5'd21, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001a3, 5'd25, 27'h000000c7, 5'd0, 27'h00000154, 32'h00000400,
  1'd1,  5'd12, 27'h0000026b, 5'd21, 27'h000003b6, 5'd12, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d7, 5'd24, 27'h000001a3, 5'd21, 27'h000001b9, 32'h00000400,
  1'd1,  5'd21, 27'h000000c3, 5'd3, 27'h0000026a, 5'd4, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003db, 5'd3, 27'h0000035c, 5'd13, 27'h00000350, 32'h00000400,
  1'd1,  5'd20, 27'h000002c0, 5'd1, 27'h0000038d, 5'd22, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003e3, 5'd13, 27'h000002a4, 5'd3, 27'h000001ba, 32'h00000400,
  1'd1,  5'd21, 27'h00000023, 5'd15, 27'h0000004a, 5'd13, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000329, 5'd15, 27'h000000c4, 5'd25, 27'h000002ed, 32'h00000400,
  1'd1,  5'd21, 27'h000000ff, 5'd25, 27'h0000005d, 5'd0, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000039d, 5'd21, 27'h00000121, 5'd11, 27'h000000ba, 32'h00000400,
  1'd1,  5'd24, 27'h00000249, 5'd25, 27'h000002dd, 5'd23, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000028f, 5'd5, 27'h0000000e, 5'd9, 27'h000003c2, 32'h00000400,
  1'd1,  5'd1, 27'h0000029b, 5'd4, 27'h0000035e, 5'd18, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000011b, 5'd0, 27'h000001f5, 5'd26, 27'h00000049, 32'h00000400,
  1'd1,  5'd2, 27'h00000175, 5'd13, 27'h00000133, 5'd6, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003df, 5'd11, 27'h00000279, 5'd17, 27'h000002da, 32'h00000400,
  1'd1,  5'd2, 27'h000002a0, 5'd12, 27'h000003f9, 5'd26, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000030a, 5'd24, 27'h000003d4, 5'd7, 27'h00000132, 32'h00000400,
  1'd1,  5'd4, 27'h000000bc, 5'd22, 27'h000002ba, 5'd20, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000026c, 5'd23, 27'h000000d1, 5'd30, 27'h00000390, 32'h00000400,
  1'd1,  5'd13, 27'h000001ea, 5'd1, 27'h000000d2, 5'd8, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002a9, 5'd0, 27'h000001c4, 5'd18, 27'h00000067, 32'h00000400,
  1'd1,  5'd11, 27'h00000029, 5'd4, 27'h00000265, 5'd30, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000038e, 5'd13, 27'h000001bb, 5'd5, 27'h0000023c, 32'h00000400,
  1'd1,  5'd12, 27'h000003eb, 5'd12, 27'h00000338, 5'd19, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001eb, 5'd11, 27'h00000154, 5'd30, 27'h0000005f, 32'h00000400,
  1'd1,  5'd12, 27'h000001a0, 5'd20, 27'h000003fe, 5'd9, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000077, 5'd25, 27'h00000060, 5'd16, 27'h000000c6, 32'h00000400,
  1'd1,  5'd11, 27'h000003ed, 5'd24, 27'h000003f0, 5'd27, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003fe, 5'd5, 27'h00000010, 5'd9, 27'h000003de, 32'h00000400,
  1'd1,  5'd24, 27'h00000163, 5'd0, 27'h00000193, 5'd17, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002bf, 5'd4, 27'h000002ff, 5'd29, 27'h000000be, 32'h00000400,
  1'd1,  5'd24, 27'h00000249, 5'd13, 27'h000003d5, 5'd8, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032a, 5'd13, 27'h000001f0, 5'd18, 27'h0000013f, 32'h00000400,
  1'd1,  5'd22, 27'h0000007d, 5'd15, 27'h000000fb, 5'd27, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b3, 5'd22, 27'h00000009, 5'd6, 27'h00000276, 32'h00000400,
  1'd1,  5'd25, 27'h0000012d, 5'd25, 27'h000000ce, 5'd18, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000001e, 5'd20, 27'h00000394, 5'd30, 27'h000000fa, 32'h00000400,
  1'd1,  5'd2, 27'h000002c8, 5'd6, 27'h000001da, 5'd3, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000351, 5'd5, 27'h00000149, 5'd14, 27'h0000036e, 32'h00000400,
  1'd1,  5'd2, 27'h000003f8, 5'd7, 27'h00000325, 5'd22, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000cd, 5'd16, 27'h000000f6, 5'd3, 27'h0000025e, 32'h00000400,
  1'd1,  5'd3, 27'h0000006c, 5'd16, 27'h00000366, 5'd11, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000155, 5'd17, 27'h000000e3, 5'd21, 27'h00000253, 32'h00000400,
  1'd1,  5'd2, 27'h0000020e, 5'd27, 27'h00000175, 5'd1, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000027, 5'd30, 27'h000001e9, 5'd10, 27'h0000039f, 32'h00000400,
  1'd1,  5'd1, 27'h0000013d, 5'd29, 27'h000001bf, 5'd21, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000210, 5'd6, 27'h00000047, 5'd0, 27'h00000057, 32'h00000400,
  1'd1,  5'd14, 27'h000001c8, 5'd8, 27'h00000021, 5'd10, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000060, 5'd7, 27'h0000014f, 5'd24, 27'h000001d7, 32'h00000400,
  1'd1,  5'd11, 27'h000003e7, 5'd18, 27'h000001fa, 5'd2, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001f7, 5'd17, 27'h0000013e, 5'd11, 27'h000002d2, 32'h00000400,
  1'd1,  5'd14, 27'h00000194, 5'd15, 27'h00000347, 5'd22, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000345, 5'd29, 27'h000001dd, 5'd1, 27'h00000136, 32'h00000400,
  1'd1,  5'd15, 27'h000001a4, 5'd26, 27'h00000386, 5'd15, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000016d, 5'd28, 27'h00000214, 5'd22, 27'h000002ad, 32'h00000400,
  1'd1,  5'd25, 27'h00000114, 5'd8, 27'h000002f6, 5'd1, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000024d, 5'd7, 27'h0000033e, 5'd13, 27'h000003e6, 32'h00000400,
  1'd1,  5'd25, 27'h00000151, 5'd5, 27'h00000366, 5'd21, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000111, 5'd19, 27'h00000181, 5'd1, 27'h000003a6, 32'h00000400,
  1'd1,  5'd21, 27'h0000023c, 5'd16, 27'h000001de, 5'd11, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000b6, 5'd18, 27'h00000361, 5'd23, 27'h000002ce, 32'h00000400,
  1'd1,  5'd21, 27'h000003e1, 5'd28, 27'h00000155, 5'd1, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000018, 5'd27, 27'h0000001f, 5'd15, 27'h000000f7, 32'h00000400,
  1'd1,  5'd25, 27'h000002db, 5'd29, 27'h00000200, 5'd25, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001fe, 5'd7, 27'h000000e1, 5'd7, 27'h0000022e, 32'h00000400,
  1'd1,  5'd4, 27'h00000024, 5'd7, 27'h000001af, 5'd19, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001b0, 5'd9, 27'h000003ba, 5'd29, 27'h00000105, 32'h00000400,
  1'd1,  5'd2, 27'h00000012, 5'd16, 27'h0000030e, 5'd9, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000313, 5'd15, 27'h0000029a, 5'd18, 27'h000000b4, 32'h00000400,
  1'd1,  5'd3, 27'h00000078, 5'd17, 27'h00000207, 5'd26, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f2, 5'd27, 27'h0000023b, 5'd10, 27'h000000fb, 32'h00000400,
  1'd1,  5'd2, 27'h0000031e, 5'd28, 27'h000000ab, 5'd16, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002fd, 5'd26, 27'h00000290, 5'd26, 27'h00000111, 32'h00000400,
  1'd1,  5'd11, 27'h000002de, 5'd8, 27'h000003b7, 5'd9, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ef, 5'd9, 27'h000002cd, 5'd17, 27'h0000008f, 32'h00000400,
  1'd1,  5'd15, 27'h0000011c, 5'd8, 27'h00000220, 5'd26, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000071, 5'd15, 27'h00000323, 5'd5, 27'h000001af, 32'h00000400,
  1'd1,  5'd14, 27'h00000042, 5'd16, 27'h00000338, 5'd15, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003b5, 5'd16, 27'h00000078, 5'd29, 27'h000000e1, 32'h00000400,
  1'd1,  5'd15, 27'h00000111, 5'd29, 27'h00000064, 5'd7, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001c6, 5'd26, 27'h00000154, 5'd17, 27'h00000054, 32'h00000400,
  1'd1,  5'd11, 27'h000001e1, 5'd30, 27'h000001a1, 5'd26, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000002d, 5'd5, 27'h000001d0, 5'd8, 27'h000001b5, 32'h00000400,
  1'd1,  5'd21, 27'h0000025d, 5'd8, 27'h000000ad, 5'd18, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002f7, 5'd5, 27'h000003ec, 5'd26, 27'h000000a0, 32'h00000400,
  1'd1,  5'd21, 27'h000001e2, 5'd17, 27'h00000089, 5'd5, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b0, 5'd18, 27'h00000155, 5'd20, 27'h0000024d, 32'h00000400,
  1'd1,  5'd25, 27'h00000198, 5'd16, 27'h00000387, 5'd28, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000086, 5'd27, 27'h00000094, 5'd7, 27'h000003f8, 32'h00000400,
  1'd1,  5'd21, 27'h00000274, 5'd30, 27'h00000016, 5'd19, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003db, 5'd29, 27'h000000c0, 5'd30, 27'h00000166, 32'h00000400,
  1'd1,  5'd8, 27'h00000052, 5'd2, 27'h0000036a, 5'd8, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ad, 5'd0, 27'h00000369, 5'd19, 27'h00000209, 32'h00000400,
  1'd1,  5'd6, 27'h000001b6, 5'd0, 27'h000001fa, 5'd28, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d9, 5'd10, 27'h00000218, 5'd2, 27'h000001c3, 32'h00000400,
  1'd1,  5'd6, 27'h00000152, 5'd10, 27'h00000381, 5'd12, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000216, 5'd15, 27'h00000025, 5'd25, 27'h000002e9, 32'h00000400,
  1'd1,  5'd9, 27'h00000114, 5'd24, 27'h000000d2, 5'd0, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000009a, 5'd21, 27'h00000351, 5'd12, 27'h0000023e, 32'h00000400,
  1'd1,  5'd6, 27'h000003c0, 5'd21, 27'h0000014d, 5'd24, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000005f, 5'd2, 27'h00000051, 5'd8, 27'h00000221, 32'h00000400,
  1'd1,  5'd17, 27'h000000ac, 5'd1, 27'h0000014d, 5'd19, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000195, 5'd3, 27'h000000eb, 5'd29, 27'h0000017a, 32'h00000400,
  1'd1,  5'd16, 27'h000003c8, 5'd11, 27'h00000042, 5'd4, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002da, 5'd14, 27'h0000023f, 5'd15, 27'h00000190, 32'h00000400,
  1'd1,  5'd15, 27'h00000265, 5'd12, 27'h000001e1, 5'd25, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000154, 5'd21, 27'h00000235, 5'd4, 27'h00000354, 32'h00000400,
  1'd1,  5'd18, 27'h000000fd, 5'd21, 27'h0000021b, 5'd11, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000027d, 5'd24, 27'h000003cb, 5'd21, 27'h00000068, 32'h00000400,
  1'd1,  5'd26, 27'h00000381, 5'd1, 27'h000002ce, 5'd2, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002f7, 5'd2, 27'h00000290, 5'd10, 27'h000001f3, 32'h00000400,
  1'd1,  5'd28, 27'h000001f8, 5'd1, 27'h000003b9, 5'd21, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000398, 5'd13, 27'h00000185, 5'd1, 27'h00000312, 32'h00000400,
  1'd1,  5'd28, 27'h00000278, 5'd13, 27'h000002aa, 5'd15, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000304, 5'd11, 27'h000000e2, 5'd22, 27'h000002b9, 32'h00000400,
  1'd1,  5'd30, 27'h000002c8, 5'd20, 27'h000003c6, 5'd3, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000031d, 5'd25, 27'h000000af, 5'd13, 27'h00000265, 32'h00000400,
  1'd1,  5'd25, 27'h000003d2, 5'd24, 27'h000002be, 5'd21, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003fb, 5'd0, 27'h0000033f, 5'd5, 27'h00000036, 32'h00000400,
  1'd1,  5'd9, 27'h0000029b, 5'd4, 27'h000002f0, 5'd13, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000197, 5'd2, 27'h00000342, 5'd25, 27'h00000253, 32'h00000400,
  1'd1,  5'd10, 27'h000000e9, 5'd11, 27'h000000b1, 5'd10, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002fb, 5'd10, 27'h00000267, 5'd20, 27'h00000172, 32'h00000400,
  1'd1,  5'd9, 27'h00000331, 5'd14, 27'h0000031c, 5'd26, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000029e, 5'd24, 27'h00000319, 5'd8, 27'h000000db, 32'h00000400,
  1'd1,  5'd8, 27'h000003f8, 5'd25, 27'h0000006e, 5'd19, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000169, 5'd23, 27'h000003a2, 5'd28, 27'h0000027d, 32'h00000400,
  1'd1,  5'd16, 27'h00000004, 5'd3, 27'h00000007, 5'd2, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000148, 5'd5, 27'h00000020, 5'd10, 27'h00000378, 32'h00000400,
  1'd1,  5'd18, 27'h0000033d, 5'd0, 27'h00000056, 5'd24, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009d, 5'd15, 27'h000000eb, 5'd7, 27'h00000201, 32'h00000400,
  1'd1,  5'd20, 27'h00000117, 5'd13, 27'h000002d7, 5'd19, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000cd, 5'd10, 27'h00000234, 5'd26, 27'h000000ca, 32'h00000400,
  1'd1,  5'd17, 27'h000001ce, 5'd22, 27'h000003ca, 5'd9, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000019f, 5'd23, 27'h00000088, 5'd17, 27'h000001c3, 32'h00000400,
  1'd1,  5'd18, 27'h00000163, 5'd22, 27'h00000281, 5'd28, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000304, 5'd1, 27'h00000215, 5'd8, 27'h00000371, 32'h00000400,
  1'd1,  5'd28, 27'h00000148, 5'd4, 27'h0000016d, 5'd16, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003a9, 5'd2, 27'h000002c6, 5'd30, 27'h0000029a, 32'h00000400,
  1'd1,  5'd27, 27'h000001da, 5'd15, 27'h000000ac, 5'd6, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003f9, 5'd13, 27'h000003fb, 5'd16, 27'h000003ff, 32'h00000400,
  1'd1,  5'd29, 27'h00000304, 5'd11, 27'h000002d4, 5'd30, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c8, 5'd22, 27'h00000170, 5'd9, 27'h000000fa, 32'h00000400,
  1'd1,  5'd27, 27'h00000109, 5'd22, 27'h0000022c, 5'd17, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a1, 5'd20, 27'h0000034c, 5'd30, 27'h00000240, 32'h00000400,
  1'd1,  5'd9, 27'h00000198, 5'd8, 27'h00000144, 5'd1, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000034d, 5'd8, 27'h00000017, 5'd15, 27'h00000134, 32'h00000400,
  1'd1,  5'd6, 27'h000001ef, 5'd8, 27'h000000d7, 5'd24, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000cf, 5'd19, 27'h00000225, 5'd0, 27'h00000377, 32'h00000400,
  1'd1,  5'd7, 27'h00000145, 5'd17, 27'h0000016d, 5'd11, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000020d, 5'd20, 27'h00000010, 5'd22, 27'h00000059, 32'h00000400,
  1'd1,  5'd9, 27'h0000031b, 5'd30, 27'h00000073, 5'd2, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d7, 5'd27, 27'h00000246, 5'd13, 27'h000003e3, 32'h00000400,
  1'd1,  5'd7, 27'h00000070, 5'd28, 27'h0000027b, 5'd24, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000123, 5'd10, 27'h00000047, 5'd3, 27'h000000f9, 32'h00000400,
  1'd1,  5'd16, 27'h0000013d, 5'd8, 27'h000001a0, 5'd10, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000036, 5'd8, 27'h00000293, 5'd24, 27'h00000095, 32'h00000400,
  1'd1,  5'd20, 27'h000001b2, 5'd18, 27'h000000e0, 5'd0, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000200, 5'd19, 27'h00000315, 5'd12, 27'h000000cf, 32'h00000400,
  1'd1,  5'd20, 27'h000000cc, 5'd18, 27'h000001bc, 5'd24, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000033e, 5'd26, 27'h00000218, 5'd2, 27'h00000115, 32'h00000400,
  1'd1,  5'd15, 27'h00000225, 5'd28, 27'h0000008e, 5'd13, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000162, 5'd29, 27'h0000012b, 5'd20, 27'h0000033e, 32'h00000400,
  1'd1,  5'd26, 27'h0000036e, 5'd7, 27'h00000261, 5'd4, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000362, 5'd5, 27'h000003c8, 5'd13, 27'h0000020a, 32'h00000400,
  1'd1,  5'd28, 27'h00000230, 5'd5, 27'h0000010b, 5'd25, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000341, 5'd18, 27'h0000027c, 5'd2, 27'h0000021f, 32'h00000400,
  1'd1,  5'd27, 27'h00000191, 5'd18, 27'h00000089, 5'd10, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000034a, 5'd18, 27'h00000379, 5'd24, 27'h00000365, 32'h00000400,
  1'd1,  5'd28, 27'h00000011, 5'd28, 27'h00000064, 5'd2, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000178, 5'd30, 27'h000001d6, 5'd12, 27'h0000005c, 32'h00000400,
  1'd1,  5'd30, 27'h0000014e, 5'd30, 27'h0000005c, 5'd24, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000eb, 5'd6, 27'h000000f8, 5'd7, 27'h00000247, 32'h00000400,
  1'd1,  5'd6, 27'h000003f7, 5'd8, 27'h000003d5, 5'd17, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002c8, 5'd8, 27'h0000030e, 5'd27, 27'h0000027a, 32'h00000400,
  1'd1,  5'd5, 27'h0000017a, 5'd18, 27'h00000180, 5'd8, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002a5, 5'd17, 27'h0000007e, 5'd17, 27'h000001b1, 32'h00000400,
  1'd1,  5'd5, 27'h00000355, 5'd16, 27'h000000fd, 5'd26, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000111, 5'd26, 27'h000000c6, 5'd5, 27'h000000b5, 32'h00000400,
  1'd1,  5'd7, 27'h000002b4, 5'd28, 27'h000001dd, 5'd15, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000173, 5'd25, 27'h00000356, 5'd28, 27'h0000019a, 32'h00000400,
  1'd1,  5'd20, 27'h0000024e, 5'd6, 27'h00000177, 5'd10, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000018f, 5'd8, 27'h00000344, 5'd16, 27'h000003b7, 32'h00000400,
  1'd1,  5'd18, 27'h000000fe, 5'd9, 27'h00000078, 5'd28, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000212, 5'd16, 27'h000002e8, 5'd10, 27'h000000c4, 32'h00000400,
  1'd1,  5'd18, 27'h000002df, 5'd16, 27'h00000370, 5'd19, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000054, 5'd20, 27'h000000f2, 5'd26, 27'h00000157, 32'h00000400,
  1'd1,  5'd16, 27'h0000021c, 5'd28, 27'h000003eb, 5'd7, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000023b, 5'd29, 27'h00000292, 5'd16, 27'h00000301, 32'h00000400,
  1'd1,  5'd17, 27'h0000014c, 5'd26, 27'h0000020d, 5'd26, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a4, 5'd5, 27'h0000021d, 5'd6, 27'h00000220, 32'h00000400,
  1'd1,  5'd30, 27'h0000021d, 5'd5, 27'h00000204, 5'd20, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b2, 5'd8, 27'h0000021d, 5'd29, 27'h0000035e, 32'h00000400,
  1'd1,  5'd29, 27'h00000372, 5'd17, 27'h000000de, 5'd7, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000255, 5'd16, 27'h00000066, 5'd16, 27'h00000284, 32'h00000400,
  1'd1,  5'd26, 27'h00000073, 5'd17, 27'h000000ac, 5'd28, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f2, 5'd30, 27'h0000031b, 5'd7, 27'h00000161, 32'h00000400,
  1'd1,  5'd29, 27'h0000037b, 5'd28, 27'h00000245, 5'd17, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000060, 5'd30, 27'h000000c0, 5'd25, 27'h000003f5, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h0000013d, 5'd1, 27'h000003c2, 5'd1, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001f0, 5'd3, 27'h000000d1, 5'd13, 27'h0000026a, 32'h00000400,
  1'd1,  5'd1, 27'h000000c4, 5'd1, 27'h00000049, 5'd23, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000267, 5'd10, 27'h0000016b, 5'd1, 27'h0000000c, 32'h00000400,
  1'd1,  5'd0, 27'h000000d8, 5'd13, 27'h00000308, 5'd12, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000025, 5'd13, 27'h000000e8, 5'd23, 27'h0000025b, 32'h00000400,
  1'd1,  5'd5, 27'h000000aa, 5'd23, 27'h000000a2, 5'd4, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b3, 5'd25, 27'h000002c5, 5'd10, 27'h0000029f, 32'h00000400,
  1'd1,  5'd0, 27'h00000174, 5'd22, 27'h00000048, 5'd23, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000025e, 5'd5, 27'h000000a1, 5'd3, 27'h00000304, 32'h00000400,
  1'd1,  5'd15, 27'h0000018a, 5'd2, 27'h00000399, 5'd10, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000327, 5'd4, 27'h000001cd, 5'd21, 27'h000001d9, 32'h00000400,
  1'd1,  5'd10, 27'h0000020d, 5'd10, 27'h00000158, 5'd3, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000133, 5'd14, 27'h000002ed, 5'd10, 27'h00000370, 32'h00000400,
  1'd1,  5'd11, 27'h000000a8, 5'd12, 27'h000003da, 5'd20, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000021, 5'd22, 27'h00000240, 5'd2, 27'h00000230, 32'h00000400,
  1'd1,  5'd12, 27'h00000350, 5'd23, 27'h000001d5, 5'd13, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000397, 5'd21, 27'h00000154, 5'd24, 27'h00000380, 32'h00000400,
  1'd1,  5'd20, 27'h00000353, 5'd2, 27'h000000b4, 5'd1, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d9, 5'd1, 27'h00000344, 5'd11, 27'h000000da, 32'h00000400,
  1'd1,  5'd24, 27'h00000087, 5'd1, 27'h000003c3, 5'd23, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001bd, 5'd11, 27'h00000326, 5'd1, 27'h00000122, 32'h00000400,
  1'd1,  5'd24, 27'h000001d5, 5'd10, 27'h000001fd, 5'd10, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e4, 5'd13, 27'h000002de, 5'd21, 27'h000003d7, 32'h00000400,
  1'd1,  5'd24, 27'h000003bc, 5'd24, 27'h000003a6, 5'd4, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000077, 5'd22, 27'h000002a0, 5'd10, 27'h000001a6, 32'h00000400,
  1'd1,  5'd23, 27'h00000125, 5'd25, 27'h0000007f, 5'd22, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000031e, 5'd1, 27'h00000164, 5'd7, 27'h00000218, 32'h00000400,
  1'd1,  5'd4, 27'h00000124, 5'd4, 27'h000003f7, 5'd16, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003df, 5'd0, 27'h00000399, 5'd30, 27'h00000105, 32'h00000400,
  1'd1,  5'd1, 27'h000002a9, 5'd11, 27'h0000001d, 5'd8, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000263, 5'd11, 27'h00000218, 5'd18, 27'h00000355, 32'h00000400,
  1'd1,  5'd4, 27'h00000298, 5'd12, 27'h000001b5, 5'd29, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000114, 5'd22, 27'h00000136, 5'd9, 27'h000002a4, 32'h00000400,
  1'd1,  5'd4, 27'h00000179, 5'd24, 27'h0000016c, 5'd15, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001eb, 5'd22, 27'h0000013b, 5'd28, 27'h000003f9, 32'h00000400,
  1'd1,  5'd11, 27'h0000008f, 5'd2, 27'h00000199, 5'd8, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000260, 5'd3, 27'h00000063, 5'd19, 27'h000000b8, 32'h00000400,
  1'd1,  5'd11, 27'h0000020e, 5'd3, 27'h000003aa, 5'd30, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f8, 5'd14, 27'h00000222, 5'd5, 27'h000002db, 32'h00000400,
  1'd1,  5'd12, 27'h00000358, 5'd12, 27'h00000378, 5'd18, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000385, 5'd14, 27'h00000110, 5'd28, 27'h00000351, 32'h00000400,
  1'd1,  5'd11, 27'h00000258, 5'd22, 27'h000003c6, 5'd8, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000046, 5'd23, 27'h0000020a, 5'd19, 27'h0000027a, 32'h00000400,
  1'd1,  5'd12, 27'h0000009d, 5'd25, 27'h000002e3, 5'd29, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000107, 5'd1, 27'h000003f3, 5'd5, 27'h000001e4, 32'h00000400,
  1'd1,  5'd22, 27'h00000108, 5'd3, 27'h000002c4, 5'd17, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ac, 5'd4, 27'h000003d2, 5'd27, 27'h000001f7, 32'h00000400,
  1'd1,  5'd24, 27'h000002c5, 5'd13, 27'h000002a0, 5'd9, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001d7, 5'd13, 27'h00000180, 5'd18, 27'h000001e1, 32'h00000400,
  1'd1,  5'd24, 27'h0000006e, 5'd13, 27'h00000176, 5'd28, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000048, 5'd20, 27'h00000336, 5'd5, 27'h00000376, 32'h00000400,
  1'd1,  5'd20, 27'h0000039d, 5'd23, 27'h0000013b, 5'd18, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000006c, 5'd22, 27'h000002ab, 5'd26, 27'h00000336, 32'h00000400,
  1'd1,  5'd4, 27'h0000008f, 5'd8, 27'h000002f2, 5'd1, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b8, 5'd6, 27'h0000017e, 5'd11, 27'h00000380, 32'h00000400,
  1'd1,  5'd4, 27'h0000033b, 5'd9, 27'h000002ad, 5'd22, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000024e, 5'd16, 27'h00000281, 5'd0, 27'h000002a6, 32'h00000400,
  1'd1,  5'd1, 27'h00000061, 5'd16, 27'h00000234, 5'd12, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000ce, 5'd18, 27'h0000032c, 5'd22, 27'h00000130, 32'h00000400,
  1'd1,  5'd0, 27'h000000a8, 5'd30, 27'h00000390, 5'd3, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e8, 5'd29, 27'h000001fc, 5'd11, 27'h0000028f, 32'h00000400,
  1'd1,  5'd2, 27'h000002c1, 5'd28, 27'h00000279, 5'd21, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000374, 5'd8, 27'h0000025f, 5'd0, 27'h000000fd, 32'h00000400,
  1'd1,  5'd13, 27'h000002e5, 5'd5, 27'h0000023b, 5'd11, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000024f, 5'd6, 27'h000000c2, 5'd24, 27'h0000034c, 32'h00000400,
  1'd1,  5'd11, 27'h000001c4, 5'd17, 27'h000000a7, 5'd3, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000310, 5'd15, 27'h000002cb, 5'd13, 27'h00000338, 32'h00000400,
  1'd1,  5'd14, 27'h00000286, 5'd16, 27'h000002ec, 5'd23, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000111, 5'd27, 27'h000000cd, 5'd5, 27'h0000008a, 32'h00000400,
  1'd1,  5'd12, 27'h000002e5, 5'd27, 27'h000003d8, 5'd11, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000035, 5'd30, 27'h000000f3, 5'd23, 27'h000000e9, 32'h00000400,
  1'd1,  5'd21, 27'h000003c3, 5'd7, 27'h00000064, 5'd1, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000bf, 5'd7, 27'h00000085, 5'd12, 27'h000001d6, 32'h00000400,
  1'd1,  5'd25, 27'h0000002e, 5'd7, 27'h0000009f, 5'd22, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000020c, 5'd20, 27'h00000244, 5'd1, 27'h000003a4, 32'h00000400,
  1'd1,  5'd20, 27'h000002f6, 5'd17, 27'h00000284, 5'd11, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000112, 5'd18, 27'h00000175, 5'd25, 27'h000002a4, 32'h00000400,
  1'd1,  5'd22, 27'h0000034d, 5'd28, 27'h00000186, 5'd4, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000022b, 5'd27, 27'h00000029, 5'd11, 27'h00000094, 32'h00000400,
  1'd1,  5'd23, 27'h000001a2, 5'd27, 27'h00000348, 5'd21, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000232, 5'd6, 27'h00000060, 5'd6, 27'h000002fa, 32'h00000400,
  1'd1,  5'd2, 27'h00000349, 5'd5, 27'h00000136, 5'd15, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000002b, 5'd10, 27'h00000025, 5'd29, 27'h000002d3, 32'h00000400,
  1'd1,  5'd4, 27'h0000032a, 5'd18, 27'h0000036b, 5'd5, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000140, 5'd18, 27'h00000234, 5'd19, 27'h0000020f, 32'h00000400,
  1'd1,  5'd3, 27'h000001ea, 5'd15, 27'h0000021b, 5'd26, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000220, 5'd28, 27'h00000209, 5'd7, 27'h0000017a, 32'h00000400,
  1'd1,  5'd5, 27'h0000009a, 5'd28, 27'h000002d1, 5'd19, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b7, 5'd29, 27'h0000036e, 5'd29, 27'h00000040, 32'h00000400,
  1'd1,  5'd11, 27'h0000008e, 5'd8, 27'h00000229, 5'd10, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000194, 5'd5, 27'h000001f2, 5'd20, 27'h00000275, 32'h00000400,
  1'd1,  5'd11, 27'h000001e6, 5'd10, 27'h00000055, 5'd27, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000012b, 5'd20, 27'h0000010d, 5'd10, 27'h0000012d, 32'h00000400,
  1'd1,  5'd12, 27'h00000325, 5'd17, 27'h0000036a, 5'd18, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000035a, 5'd18, 27'h00000319, 5'd30, 27'h00000224, 32'h00000400,
  1'd1,  5'd11, 27'h0000012a, 5'd29, 27'h00000323, 5'd6, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000295, 5'd28, 27'h00000067, 5'd20, 27'h00000213, 32'h00000400,
  1'd1,  5'd14, 27'h00000306, 5'd30, 27'h0000012d, 5'd30, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000151, 5'd9, 27'h00000100, 5'd6, 27'h00000264, 32'h00000400,
  1'd1,  5'd25, 27'h000001ed, 5'd5, 27'h00000218, 5'd16, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001c6, 5'd7, 27'h0000018a, 5'd29, 27'h000002de, 32'h00000400,
  1'd1,  5'd23, 27'h000003c3, 5'd18, 27'h00000320, 5'd8, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000c1, 5'd19, 27'h00000187, 5'd17, 27'h00000065, 32'h00000400,
  1'd1,  5'd25, 27'h0000000a, 5'd15, 27'h00000390, 5'd27, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d3, 5'd26, 27'h00000072, 5'd8, 27'h000000e3, 32'h00000400,
  1'd1,  5'd25, 27'h00000122, 5'd27, 27'h000001eb, 5'd16, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000277, 5'd28, 27'h00000018, 5'd30, 27'h000002a8, 32'h00000400,
  1'd1,  5'd6, 27'h000002e8, 5'd0, 27'h000000af, 5'd5, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003fb, 5'd1, 27'h000001f2, 5'd18, 27'h0000026a, 32'h00000400,
  1'd1,  5'd5, 27'h00000253, 5'd3, 27'h00000280, 5'd28, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000350, 5'd13, 27'h000001b9, 5'd3, 27'h0000022c, 32'h00000400,
  1'd1,  5'd8, 27'h000003e6, 5'd14, 27'h000000b7, 5'd10, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000036c, 5'd10, 27'h000003b9, 5'd25, 27'h00000045, 32'h00000400,
  1'd1,  5'd10, 27'h000000ed, 5'd21, 27'h0000032f, 5'd4, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000146, 5'd24, 27'h00000288, 5'd13, 27'h000001e5, 32'h00000400,
  1'd1,  5'd7, 27'h000003a2, 5'd25, 27'h00000262, 5'd25, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000172, 5'd4, 27'h000003ca, 5'd7, 27'h00000388, 32'h00000400,
  1'd1,  5'd18, 27'h000002db, 5'd1, 27'h000003b4, 5'd16, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000039f, 5'd0, 27'h00000166, 5'd30, 27'h0000007f, 32'h00000400,
  1'd1,  5'd17, 27'h00000301, 5'd11, 27'h00000164, 5'd1, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000016f, 5'd12, 27'h00000051, 5'd12, 27'h000000f1, 32'h00000400,
  1'd1,  5'd19, 27'h0000026a, 5'd14, 27'h000002a0, 5'd25, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000000d, 5'd24, 27'h00000170, 5'd3, 27'h000001b9, 32'h00000400,
  1'd1,  5'd16, 27'h000000a0, 5'd23, 27'h0000035c, 5'd10, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002a7, 5'd22, 27'h0000009c, 5'd24, 27'h0000011f, 32'h00000400,
  1'd1,  5'd28, 27'h00000341, 5'd4, 27'h0000013b, 5'd2, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000cc, 5'd3, 27'h000001ed, 5'd10, 27'h00000306, 32'h00000400,
  1'd1,  5'd26, 27'h00000147, 5'd4, 27'h00000364, 5'd22, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000164, 5'd13, 27'h00000076, 5'd3, 27'h0000003e, 32'h00000400,
  1'd1,  5'd27, 27'h00000385, 5'd11, 27'h000000e9, 5'd12, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c3, 5'd13, 27'h000003b7, 5'd25, 27'h000001f9, 32'h00000400,
  1'd1,  5'd30, 27'h0000009f, 5'd23, 27'h0000024d, 5'd3, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001fb, 5'd22, 27'h00000037, 5'd12, 27'h000003bd, 32'h00000400,
  1'd1,  5'd30, 27'h00000346, 5'd21, 27'h000000aa, 5'd25, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018b, 5'd1, 27'h000002a8, 5'd4, 27'h000000a8, 32'h00000400,
  1'd1,  5'd7, 27'h00000020, 5'd4, 27'h000002f1, 5'd11, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000367, 5'd3, 27'h000000f2, 5'd25, 27'h00000094, 32'h00000400,
  1'd1,  5'd8, 27'h00000305, 5'd15, 27'h00000033, 5'd6, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002b9, 5'd14, 27'h000001e8, 5'd16, 27'h00000285, 32'h00000400,
  1'd1,  5'd9, 27'h0000000d, 5'd11, 27'h00000091, 5'd29, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000258, 5'd22, 27'h00000055, 5'd9, 27'h00000274, 32'h00000400,
  1'd1,  5'd9, 27'h00000322, 5'd24, 27'h0000038d, 5'd16, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f1, 5'd24, 27'h000002a2, 5'd27, 27'h0000011c, 32'h00000400,
  1'd1,  5'd19, 27'h00000096, 5'd1, 27'h000001d1, 5'd2, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000037, 5'd2, 27'h0000007e, 5'd15, 27'h0000002d, 32'h00000400,
  1'd1,  5'd20, 27'h00000063, 5'd0, 27'h000000e7, 5'd22, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000187, 5'd12, 27'h0000019e, 5'd6, 27'h0000009d, 32'h00000400,
  1'd1,  5'd19, 27'h0000027e, 5'd11, 27'h000002ec, 5'd19, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001bd, 5'd12, 27'h000002f5, 5'd28, 27'h000002a7, 32'h00000400,
  1'd1,  5'd17, 27'h0000025f, 5'd25, 27'h000000c9, 5'd9, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001a0, 5'd21, 27'h000000d6, 5'd17, 27'h000001f9, 32'h00000400,
  1'd1,  5'd20, 27'h0000002f, 5'd22, 27'h00000186, 5'd30, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000020, 5'd3, 27'h000003b0, 5'd9, 27'h000002ae, 32'h00000400,
  1'd1,  5'd26, 27'h0000039b, 5'd4, 27'h0000027e, 5'd16, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000168, 5'd2, 27'h00000207, 5'd27, 27'h00000024, 32'h00000400,
  1'd1,  5'd29, 27'h00000249, 5'd12, 27'h000001a1, 5'd7, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002bd, 5'd14, 27'h0000030e, 5'd16, 27'h00000108, 32'h00000400,
  1'd1,  5'd28, 27'h000000f7, 5'd11, 27'h0000018e, 5'd30, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000135, 5'd23, 27'h000002b1, 5'd8, 27'h00000038, 32'h00000400,
  1'd1,  5'd28, 27'h000001c5, 5'd20, 27'h00000387, 5'd19, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000143, 5'd24, 27'h0000001e, 5'd28, 27'h000001e3, 32'h00000400,
  1'd1,  5'd6, 27'h00000207, 5'd7, 27'h0000002c, 5'd4, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000298, 5'd10, 27'h000000b6, 5'd10, 27'h0000020d, 32'h00000400,
  1'd1,  5'd8, 27'h000001e9, 5'd7, 27'h000003a4, 5'd20, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000134, 5'd16, 27'h0000018a, 5'd0, 27'h000003cf, 32'h00000400,
  1'd1,  5'd6, 27'h00000294, 5'd15, 27'h00000394, 5'd14, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000314, 5'd16, 27'h000000e4, 5'd25, 27'h000000e6, 32'h00000400,
  1'd1,  5'd8, 27'h00000069, 5'd27, 27'h0000030e, 5'd4, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ba, 5'd27, 27'h000001cf, 5'd11, 27'h0000005a, 32'h00000400,
  1'd1,  5'd6, 27'h000003ed, 5'd28, 27'h00000218, 5'd24, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000038b, 5'd8, 27'h000003f9, 5'd3, 27'h000000f1, 32'h00000400,
  1'd1,  5'd20, 27'h0000007c, 5'd8, 27'h00000374, 5'd12, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000df, 5'd6, 27'h000000c7, 5'd25, 27'h000000e0, 32'h00000400,
  1'd1,  5'd15, 27'h00000343, 5'd19, 27'h0000036f, 5'd1, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d9, 5'd20, 27'h000000ad, 5'd11, 27'h00000396, 32'h00000400,
  1'd1,  5'd19, 27'h0000010b, 5'd16, 27'h000002e8, 5'd20, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000221, 5'd30, 27'h0000003b, 5'd4, 27'h000003af, 32'h00000400,
  1'd1,  5'd18, 27'h000000b9, 5'd28, 27'h00000030, 5'd14, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001b9, 5'd25, 27'h000003b6, 5'd22, 27'h000002ef, 32'h00000400,
  1'd1,  5'd27, 27'h00000334, 5'd6, 27'h0000007e, 5'd2, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001d4, 5'd9, 27'h0000035d, 5'd11, 27'h000001e0, 32'h00000400,
  1'd1,  5'd27, 27'h00000221, 5'd9, 27'h00000384, 5'd22, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d1, 5'd17, 27'h00000128, 5'd3, 27'h0000038c, 32'h00000400,
  1'd1,  5'd26, 27'h0000024d, 5'd16, 27'h000003b8, 5'd13, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000fa, 5'd18, 27'h00000272, 5'd25, 27'h0000033c, 32'h00000400,
  1'd1,  5'd29, 27'h000002b8, 5'd26, 27'h000000c3, 5'd4, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000036d, 5'd28, 27'h00000027, 5'd12, 27'h00000300, 32'h00000400,
  1'd1,  5'd30, 27'h00000292, 5'd28, 27'h000003a2, 5'd20, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000016c, 5'd7, 27'h000000fa, 5'd7, 27'h0000030e, 32'h00000400,
  1'd1,  5'd6, 27'h00000033, 5'd6, 27'h00000359, 5'd17, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000017d, 5'd8, 27'h0000009b, 5'd30, 27'h00000303, 32'h00000400,
  1'd1,  5'd6, 27'h000000f6, 5'd16, 27'h000001ea, 5'd5, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003f2, 5'd18, 27'h000000e9, 5'd20, 27'h000001f7, 32'h00000400,
  1'd1,  5'd5, 27'h0000031b, 5'd17, 27'h000001e7, 5'd28, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000018f, 5'd26, 27'h00000226, 5'd5, 27'h000003dc, 32'h00000400,
  1'd1,  5'd7, 27'h000003cc, 5'd30, 27'h0000030f, 5'd18, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000369, 5'd29, 27'h000000cb, 5'd27, 27'h0000033e, 32'h00000400,
  1'd1,  5'd16, 27'h00000054, 5'd7, 27'h0000038a, 5'd10, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000005f, 5'd7, 27'h00000084, 5'd15, 27'h0000033d, 32'h00000400,
  1'd1,  5'd17, 27'h00000048, 5'd9, 27'h000002e6, 5'd26, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000047, 5'd15, 27'h000002f8, 5'd7, 27'h00000116, 32'h00000400,
  1'd1,  5'd16, 27'h0000036d, 5'd20, 27'h0000026b, 5'd17, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000026b, 5'd16, 27'h00000078, 5'd30, 27'h000003c5, 32'h00000400,
  1'd1,  5'd17, 27'h000003bd, 5'd28, 27'h000001ac, 5'd7, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000222, 5'd29, 27'h0000032b, 5'd20, 27'h00000218, 32'h00000400,
  1'd1,  5'd15, 27'h000003a7, 5'd29, 27'h0000026b, 5'd30, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000303, 5'd5, 27'h000001d4, 5'd7, 27'h00000264, 32'h00000400,
  1'd1,  5'd29, 27'h0000025d, 5'd6, 27'h000001f5, 5'd20, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000122, 5'd6, 27'h000002dc, 5'd28, 27'h0000019f, 32'h00000400,
  1'd1,  5'd29, 27'h00000278, 5'd19, 27'h00000157, 5'd8, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000071, 5'd17, 27'h00000302, 5'd17, 27'h000001fa, 32'h00000400,
  1'd1,  5'd27, 27'h0000010c, 5'd18, 27'h00000318, 5'd28, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000225, 5'd29, 27'h0000029a, 5'd5, 27'h00000188, 32'h00000400,
  1'd1,  5'd27, 27'h00000135, 5'd30, 27'h00000091, 5'd20, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000008c, 5'd27, 27'h000000a4, 5'd27, 27'h0000025a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000002bd, 5'd4, 27'h00000136, 5'd0, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000360, 5'd4, 27'h000000a2, 5'd14, 27'h0000019c, 32'h00000400,
  1'd1,  5'd4, 27'h000003e4, 5'd3, 27'h000000d3, 5'd23, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000354, 5'd14, 27'h0000016c, 5'd2, 27'h00000226, 32'h00000400,
  1'd1,  5'd0, 27'h000000a7, 5'd15, 27'h000000be, 5'd13, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029e, 5'd12, 27'h00000047, 5'd22, 27'h000002fe, 32'h00000400,
  1'd1,  5'd0, 27'h000002c4, 5'd22, 27'h000000aa, 5'd3, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000033f, 5'd20, 27'h00000336, 5'd10, 27'h00000156, 32'h00000400,
  1'd1,  5'd5, 27'h00000065, 5'd20, 27'h00000333, 5'd22, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000117, 5'd2, 27'h000003f6, 5'd3, 27'h00000131, 32'h00000400,
  1'd1,  5'd12, 27'h00000064, 5'd3, 27'h00000263, 5'd12, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c8, 5'd2, 27'h00000256, 5'd21, 27'h0000035e, 32'h00000400,
  1'd1,  5'd12, 27'h00000288, 5'd13, 27'h000001d7, 5'd4, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000276, 5'd11, 27'h000003cf, 5'd14, 27'h0000039c, 32'h00000400,
  1'd1,  5'd12, 27'h00000323, 5'd14, 27'h00000171, 5'd24, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000dd, 5'd23, 27'h000001f6, 5'd3, 27'h0000018c, 32'h00000400,
  1'd1,  5'd12, 27'h00000334, 5'd25, 27'h0000014f, 5'd13, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ff, 5'd21, 27'h000000fa, 5'd22, 27'h00000091, 32'h00000400,
  1'd1,  5'd25, 27'h0000009a, 5'd5, 27'h0000003e, 5'd4, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000220, 5'd2, 27'h00000111, 5'd10, 27'h000003bd, 32'h00000400,
  1'd1,  5'd20, 27'h0000031f, 5'd4, 27'h0000017a, 5'd23, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001d0, 5'd11, 27'h0000032f, 5'd2, 27'h0000001c, 32'h00000400,
  1'd1,  5'd23, 27'h000003ee, 5'd13, 27'h000000aa, 5'd11, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003d3, 5'd12, 27'h000003be, 5'd21, 27'h000001b0, 32'h00000400,
  1'd1,  5'd22, 27'h000001f0, 5'd24, 27'h00000008, 5'd1, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000312, 5'd23, 27'h000000a0, 5'd15, 27'h000000ce, 32'h00000400,
  1'd1,  5'd21, 27'h000000f3, 5'd24, 27'h00000131, 5'd21, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ba, 5'd0, 27'h000001a5, 5'd8, 27'h00000098, 32'h00000400,
  1'd1,  5'd2, 27'h00000243, 5'd3, 27'h00000209, 5'd20, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000fe, 5'd3, 27'h000001c5, 5'd28, 27'h00000224, 32'h00000400,
  1'd1,  5'd3, 27'h00000136, 5'd12, 27'h000002c3, 5'd9, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003fb, 5'd10, 27'h0000036d, 5'd15, 27'h00000240, 32'h00000400,
  1'd1,  5'd4, 27'h000003aa, 5'd13, 27'h00000225, 5'd30, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039a, 5'd24, 27'h0000014e, 5'd9, 27'h000003b9, 32'h00000400,
  1'd1,  5'd0, 27'h0000013c, 5'd20, 27'h000002ba, 5'd20, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000349, 5'd25, 27'h0000031c, 5'd26, 27'h0000004a, 32'h00000400,
  1'd1,  5'd15, 27'h00000138, 5'd4, 27'h000001a6, 5'd8, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003b0, 5'd1, 27'h000000af, 5'd19, 27'h00000238, 32'h00000400,
  1'd1,  5'd12, 27'h000000fb, 5'd2, 27'h000003d0, 5'd27, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000247, 5'd11, 27'h00000354, 5'd5, 27'h000000f5, 32'h00000400,
  1'd1,  5'd14, 27'h0000026b, 5'd12, 27'h0000024c, 5'd19, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000036, 5'd11, 27'h00000373, 5'd29, 27'h000002cc, 32'h00000400,
  1'd1,  5'd14, 27'h000002a2, 5'd25, 27'h000002d2, 5'd8, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038b, 5'd21, 27'h000002e3, 5'd19, 27'h00000322, 32'h00000400,
  1'd1,  5'd14, 27'h000000aa, 5'd22, 27'h00000141, 5'd30, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000016d, 5'd0, 27'h0000007d, 5'd8, 27'h0000005c, 32'h00000400,
  1'd1,  5'd24, 27'h0000005c, 5'd2, 27'h000002b8, 5'd17, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000145, 5'd3, 27'h00000000, 5'd25, 27'h00000382, 32'h00000400,
  1'd1,  5'd21, 27'h000002b6, 5'd15, 27'h000001f1, 5'd8, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000013, 5'd13, 27'h000001dc, 5'd17, 27'h000003f7, 32'h00000400,
  1'd1,  5'd24, 27'h00000008, 5'd13, 27'h00000322, 5'd28, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002cf, 5'd22, 27'h000001d4, 5'd8, 27'h000003b1, 32'h00000400,
  1'd1,  5'd24, 27'h000003b8, 5'd21, 27'h00000211, 5'd20, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002b0, 5'd22, 27'h00000185, 5'd30, 27'h000000f7, 32'h00000400,
  1'd1,  5'd3, 27'h00000018, 5'd6, 27'h00000181, 5'd5, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000141, 5'd6, 27'h000001b1, 5'd14, 27'h0000001c, 32'h00000400,
  1'd1,  5'd4, 27'h000002d0, 5'd6, 27'h0000039f, 5'd25, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000192, 5'd15, 27'h000003d0, 5'd3, 27'h00000014, 32'h00000400,
  1'd1,  5'd2, 27'h0000005b, 5'd18, 27'h000002fa, 5'd10, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000268, 5'd18, 27'h0000034f, 5'd20, 27'h00000384, 32'h00000400,
  1'd1,  5'd4, 27'h000003b1, 5'd28, 27'h00000020, 5'd0, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000312, 5'd29, 27'h00000363, 5'd14, 27'h00000046, 32'h00000400,
  1'd1,  5'd3, 27'h00000084, 5'd27, 27'h0000036f, 5'd23, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000064, 5'd9, 27'h00000043, 5'd2, 27'h0000003d, 32'h00000400,
  1'd1,  5'd11, 27'h00000051, 5'd8, 27'h000003a1, 5'd14, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f2, 5'd9, 27'h000000d1, 5'd21, 27'h000001ac, 32'h00000400,
  1'd1,  5'd11, 27'h000001fb, 5'd20, 27'h00000155, 5'd2, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b7, 5'd16, 27'h000002ac, 5'd13, 27'h0000001c, 32'h00000400,
  1'd1,  5'd11, 27'h0000000f, 5'd20, 27'h000001f4, 5'd25, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000020e, 5'd29, 27'h000003a8, 5'd3, 27'h000001bf, 32'h00000400,
  1'd1,  5'd13, 27'h000001c5, 5'd26, 27'h0000008c, 5'd11, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000019c, 5'd27, 27'h000000c1, 5'd24, 27'h000000a6, 32'h00000400,
  1'd1,  5'd21, 27'h0000021e, 5'd8, 27'h00000203, 5'd0, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000265, 5'd6, 27'h000002e1, 5'd14, 27'h00000351, 32'h00000400,
  1'd1,  5'd21, 27'h00000010, 5'd10, 27'h000000a9, 5'd22, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000012e, 5'd17, 27'h000001c9, 5'd4, 27'h000000c3, 32'h00000400,
  1'd1,  5'd23, 27'h0000028b, 5'd17, 27'h0000027c, 5'd12, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000e3, 5'd16, 27'h000003ad, 5'd21, 27'h000000cc, 32'h00000400,
  1'd1,  5'd20, 27'h000003f8, 5'd30, 27'h00000175, 5'd2, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003a6, 5'd30, 27'h0000012f, 5'd10, 27'h000002c6, 32'h00000400,
  1'd1,  5'd22, 27'h000003f7, 5'd30, 27'h00000064, 5'd24, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000034d, 5'd6, 27'h00000090, 5'd5, 27'h00000270, 32'h00000400,
  1'd1,  5'd2, 27'h000001fa, 5'd5, 27'h000001a3, 5'd18, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000333, 5'd6, 27'h0000035a, 5'd28, 27'h0000037d, 32'h00000400,
  1'd1,  5'd1, 27'h000000c0, 5'd19, 27'h000003c7, 5'd8, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000189, 5'd19, 27'h0000018e, 5'd16, 27'h00000043, 32'h00000400,
  1'd1,  5'd0, 27'h000002e0, 5'd18, 27'h0000039f, 5'd30, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000026f, 5'd28, 27'h0000013d, 5'd5, 27'h0000029b, 32'h00000400,
  1'd1,  5'd1, 27'h000003b3, 5'd28, 27'h000003d9, 5'd16, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002ea, 5'd29, 27'h0000012e, 5'd30, 27'h000001a5, 32'h00000400,
  1'd1,  5'd13, 27'h00000336, 5'd6, 27'h0000027c, 5'd5, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000390, 5'd6, 27'h000001ce, 5'd20, 27'h00000035, 32'h00000400,
  1'd1,  5'd12, 27'h00000371, 5'd7, 27'h000003a6, 5'd29, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000343, 5'd16, 27'h00000001, 5'd10, 27'h000000e6, 32'h00000400,
  1'd1,  5'd10, 27'h000001d5, 5'd19, 27'h0000016b, 5'd17, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000232, 5'd16, 27'h000002de, 5'd28, 27'h000002d4, 32'h00000400,
  1'd1,  5'd13, 27'h00000229, 5'd26, 27'h00000292, 5'd8, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000248, 5'd28, 27'h00000141, 5'd15, 27'h0000023a, 32'h00000400,
  1'd1,  5'd11, 27'h000002fc, 5'd26, 27'h000002d0, 5'd26, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002cc, 5'd6, 27'h00000043, 5'd7, 27'h0000020e, 32'h00000400,
  1'd1,  5'd25, 27'h00000182, 5'd7, 27'h000002a8, 5'd19, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032c, 5'd6, 27'h0000023a, 5'd28, 27'h00000296, 32'h00000400,
  1'd1,  5'd21, 27'h00000385, 5'd16, 27'h0000035e, 5'd9, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e2, 5'd15, 27'h0000023a, 5'd18, 27'h000001ac, 32'h00000400,
  1'd1,  5'd20, 27'h000003e6, 5'd18, 27'h000002c6, 5'd29, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000349, 5'd26, 27'h000003b4, 5'd9, 27'h0000006a, 32'h00000400,
  1'd1,  5'd25, 27'h00000073, 5'd25, 27'h00000383, 5'd18, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002d5, 5'd30, 27'h00000157, 5'd30, 27'h000003ec, 32'h00000400,
  1'd1,  5'd7, 27'h0000029e, 5'd4, 27'h0000033e, 5'd6, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000331, 5'd4, 27'h0000005d, 5'd20, 27'h000000ab, 32'h00000400,
  1'd1,  5'd8, 27'h0000037a, 5'd5, 27'h00000086, 5'd28, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000005a, 5'd15, 27'h0000018d, 5'd2, 27'h0000037a, 32'h00000400,
  1'd1,  5'd9, 27'h00000191, 5'd15, 27'h000001e9, 5'd10, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000258, 5'd11, 27'h0000004e, 5'd20, 27'h000003e6, 32'h00000400,
  1'd1,  5'd5, 27'h00000296, 5'd24, 27'h000002b7, 5'd0, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000027c, 5'd21, 27'h0000020c, 5'd13, 27'h0000035f, 32'h00000400,
  1'd1,  5'd7, 27'h000002e6, 5'd20, 27'h000002b8, 5'd22, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000095, 5'd0, 27'h000001dd, 5'd6, 27'h000003d0, 32'h00000400,
  1'd1,  5'd19, 27'h00000015, 5'd2, 27'h00000058, 5'd20, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002a6, 5'd1, 27'h000002e5, 5'd27, 27'h0000012d, 32'h00000400,
  1'd1,  5'd18, 27'h00000034, 5'd13, 27'h0000012d, 5'd0, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a0, 5'd13, 27'h000000c7, 5'd11, 27'h000002ac, 32'h00000400,
  1'd1,  5'd20, 27'h000001b5, 5'd11, 27'h000003bd, 5'd22, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a4, 5'd21, 27'h00000321, 5'd4, 27'h000003f4, 32'h00000400,
  1'd1,  5'd17, 27'h000000ea, 5'd23, 27'h00000165, 5'd13, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000027d, 5'd24, 27'h00000369, 5'd23, 27'h000000e8, 32'h00000400,
  1'd1,  5'd27, 27'h00000339, 5'd2, 27'h000002e5, 5'd4, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000316, 5'd0, 27'h0000011c, 5'd12, 27'h000003bd, 32'h00000400,
  1'd1,  5'd26, 27'h0000034c, 5'd2, 27'h0000017e, 5'd25, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ad, 5'd10, 27'h0000033d, 5'd2, 27'h0000022b, 32'h00000400,
  1'd1,  5'd26, 27'h00000033, 5'd11, 27'h000000c0, 5'd14, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000222, 5'd13, 27'h00000143, 5'd24, 27'h00000333, 32'h00000400,
  1'd1,  5'd29, 27'h000003f7, 5'd23, 27'h0000000b, 5'd0, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000199, 5'd21, 27'h0000019b, 5'd11, 27'h00000198, 32'h00000400,
  1'd1,  5'd27, 27'h00000222, 5'd23, 27'h00000116, 5'd25, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000037, 5'd3, 27'h00000017, 5'd2, 27'h000000d3, 32'h00000400,
  1'd1,  5'd6, 27'h000002e0, 5'd4, 27'h000000c9, 5'd10, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003bb, 5'd4, 27'h00000067, 5'd22, 27'h000000f6, 32'h00000400,
  1'd1,  5'd5, 27'h00000146, 5'd14, 27'h000001d5, 5'd7, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000027e, 5'd14, 27'h0000039f, 5'd18, 27'h000003f2, 32'h00000400,
  1'd1,  5'd9, 27'h000000f4, 5'd12, 27'h00000394, 5'd28, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002c6, 5'd23, 27'h0000003e, 5'd8, 27'h000002dc, 32'h00000400,
  1'd1,  5'd5, 27'h000001ce, 5'd20, 27'h0000039d, 5'd15, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ff, 5'd25, 27'h0000011c, 5'd30, 27'h00000365, 32'h00000400,
  1'd1,  5'd17, 27'h000000d1, 5'd2, 27'h000002fa, 5'd0, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029d, 5'd4, 27'h000003ec, 5'd12, 27'h00000108, 32'h00000400,
  1'd1,  5'd17, 27'h00000180, 5'd3, 27'h00000031, 5'd22, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000284, 5'd14, 27'h000003db, 5'd8, 27'h000003b9, 32'h00000400,
  1'd1,  5'd18, 27'h000003ac, 5'd11, 27'h000003e9, 5'd18, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003cc, 5'd13, 27'h0000018d, 5'd28, 27'h00000331, 32'h00000400,
  1'd1,  5'd18, 27'h00000282, 5'd24, 27'h000000f4, 5'd7, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000027c, 5'd21, 27'h000001e9, 5'd17, 27'h00000394, 32'h00000400,
  1'd1,  5'd15, 27'h00000372, 5'd23, 27'h00000024, 5'd29, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000276, 5'd1, 27'h000003b8, 5'd6, 27'h000000c0, 32'h00000400,
  1'd1,  5'd29, 27'h000002cc, 5'd0, 27'h00000359, 5'd20, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000221, 5'd3, 27'h000002f7, 5'd26, 27'h00000064, 32'h00000400,
  1'd1,  5'd27, 27'h0000032d, 5'd10, 27'h0000032a, 5'd7, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000035c, 5'd15, 27'h0000001d, 5'd19, 27'h000002a1, 32'h00000400,
  1'd1,  5'd30, 27'h0000011b, 5'd15, 27'h00000016, 5'd27, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000085, 5'd23, 27'h000003a8, 5'd10, 27'h00000072, 32'h00000400,
  1'd1,  5'd27, 27'h0000021e, 5'd24, 27'h0000009a, 5'd19, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000236, 5'd21, 27'h000003fe, 5'd27, 27'h0000008f, 32'h00000400,
  1'd1,  5'd6, 27'h00000341, 5'd9, 27'h000000a1, 5'd0, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000cd, 5'd7, 27'h0000023a, 5'd13, 27'h000002fe, 32'h00000400,
  1'd1,  5'd9, 27'h000001d4, 5'd5, 27'h000002f3, 5'd20, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000152, 5'd15, 27'h000002e0, 5'd2, 27'h00000318, 32'h00000400,
  1'd1,  5'd6, 27'h000000d6, 5'd15, 27'h0000026d, 5'd13, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000be, 5'd15, 27'h000003e5, 5'd23, 27'h000002e0, 32'h00000400,
  1'd1,  5'd5, 27'h00000324, 5'd29, 27'h00000275, 5'd2, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003d5, 5'd29, 27'h00000246, 5'd14, 27'h0000022c, 32'h00000400,
  1'd1,  5'd8, 27'h00000233, 5'd26, 27'h0000028d, 5'd24, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000148, 5'd7, 27'h0000038e, 5'd2, 27'h00000241, 32'h00000400,
  1'd1,  5'd16, 27'h00000102, 5'd10, 27'h00000126, 5'd15, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f2, 5'd5, 27'h000001ea, 5'd23, 27'h0000014a, 32'h00000400,
  1'd1,  5'd18, 27'h00000283, 5'd19, 27'h0000035f, 5'd0, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000cc, 5'd15, 27'h0000020c, 5'd12, 27'h00000319, 32'h00000400,
  1'd1,  5'd18, 27'h000002a7, 5'd17, 27'h00000031, 5'd22, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000c6, 5'd27, 27'h00000030, 5'd3, 27'h000002f6, 32'h00000400,
  1'd1,  5'd16, 27'h0000016c, 5'd28, 27'h000001b6, 5'd12, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002c8, 5'd27, 27'h000000cd, 5'd24, 27'h000000ae, 32'h00000400,
  1'd1,  5'd26, 27'h0000016c, 5'd6, 27'h00000371, 5'd3, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a3, 5'd7, 27'h0000015f, 5'd12, 27'h0000022d, 32'h00000400,
  1'd1,  5'd26, 27'h000003e7, 5'd8, 27'h000002ff, 5'd23, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000035, 5'd19, 27'h00000360, 5'd1, 27'h000003cd, 32'h00000400,
  1'd1,  5'd29, 27'h00000104, 5'd20, 27'h000000a6, 5'd12, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000294, 5'd20, 27'h00000211, 5'd23, 27'h000002d3, 32'h00000400,
  1'd1,  5'd27, 27'h000001b8, 5'd27, 27'h00000091, 5'd4, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000354, 5'd28, 27'h000001e4, 5'd12, 27'h00000061, 32'h00000400,
  1'd1,  5'd26, 27'h00000239, 5'd26, 27'h00000334, 5'd23, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000013d, 5'd10, 27'h00000115, 5'd8, 27'h000003eb, 32'h00000400,
  1'd1,  5'd5, 27'h0000029e, 5'd7, 27'h0000000d, 5'd15, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c8, 5'd9, 27'h000001ad, 5'd27, 27'h00000261, 32'h00000400,
  1'd1,  5'd9, 27'h000000ef, 5'd17, 27'h00000132, 5'd8, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a8, 5'd16, 27'h00000160, 5'd17, 27'h00000309, 32'h00000400,
  1'd1,  5'd10, 27'h0000012f, 5'd15, 27'h00000230, 5'd29, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000201, 5'd27, 27'h00000337, 5'd9, 27'h000000d4, 32'h00000400,
  1'd1,  5'd5, 27'h000000ce, 5'd30, 27'h0000036d, 5'd17, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000168, 5'd27, 27'h00000137, 5'd28, 27'h00000382, 32'h00000400,
  1'd1,  5'd20, 27'h000001f1, 5'd10, 27'h000000c1, 5'd6, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000038, 5'd8, 27'h00000039, 5'd18, 27'h000002ae, 32'h00000400,
  1'd1,  5'd20, 27'h000002a9, 5'd6, 27'h0000034d, 5'd30, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000339, 5'd17, 27'h00000114, 5'd7, 27'h00000358, 32'h00000400,
  1'd1,  5'd19, 27'h000000de, 5'd18, 27'h0000025f, 5'd17, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f1, 5'd20, 27'h00000165, 5'd27, 27'h0000010f, 32'h00000400,
  1'd1,  5'd18, 27'h000002af, 5'd26, 27'h00000386, 5'd6, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000375, 5'd28, 27'h00000345, 5'd20, 27'h0000007e, 32'h00000400,
  1'd1,  5'd16, 27'h000000d2, 5'd28, 27'h0000039c, 5'd29, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002dc, 5'd8, 27'h000000fa, 5'd7, 27'h00000399, 32'h00000400,
  1'd1,  5'd27, 27'h00000309, 5'd9, 27'h000001bb, 5'd18, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000aa, 5'd10, 27'h00000101, 5'd29, 27'h00000388, 32'h00000400,
  1'd1,  5'd29, 27'h000001fb, 5'd16, 27'h00000042, 5'd6, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000015c, 5'd17, 27'h000000e5, 5'd15, 27'h0000033a, 32'h00000400,
  1'd1,  5'd29, 27'h00000234, 5'd17, 27'h000003e3, 5'd26, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000024, 5'd29, 27'h00000001, 5'd8, 27'h000000ce, 32'h00000400,
  1'd1,  5'd28, 27'h000003f2, 5'd30, 27'h00000072, 5'd17, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e9, 5'd27, 27'h00000008, 5'd26, 27'h00000370, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000039d, 5'd2, 27'h000003ba, 5'd4, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000249, 5'd4, 27'h00000102, 5'd13, 27'h00000181, 32'h00000400,
  1'd1,  5'd2, 27'h00000269, 5'd3, 27'h00000070, 5'd22, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e5, 5'd12, 27'h000003ea, 5'd3, 27'h000001a3, 32'h00000400,
  1'd1,  5'd2, 27'h0000002d, 5'd12, 27'h000003e4, 5'd11, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000134, 5'd12, 27'h0000038d, 5'd21, 27'h00000272, 32'h00000400,
  1'd1,  5'd0, 27'h000002b5, 5'd22, 27'h000003b8, 5'd1, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014a, 5'd24, 27'h000000d4, 5'd11, 27'h00000146, 32'h00000400,
  1'd1,  5'd0, 27'h00000189, 5'd22, 27'h00000354, 5'd23, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ad, 5'd4, 27'h000001b3, 5'd3, 27'h0000032f, 32'h00000400,
  1'd1,  5'd15, 27'h000000a5, 5'd2, 27'h000000e7, 5'd13, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a4, 5'd2, 27'h00000323, 5'd20, 27'h000002b2, 32'h00000400,
  1'd1,  5'd11, 27'h0000033f, 5'd15, 27'h00000090, 5'd4, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000021b, 5'd14, 27'h00000006, 5'd14, 27'h00000356, 32'h00000400,
  1'd1,  5'd10, 27'h00000388, 5'd12, 27'h00000282, 5'd24, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e6, 5'd22, 27'h0000031a, 5'd5, 27'h00000001, 32'h00000400,
  1'd1,  5'd13, 27'h00000187, 5'd20, 27'h000003eb, 5'd11, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000247, 5'd21, 27'h00000089, 5'd24, 27'h0000025d, 32'h00000400,
  1'd1,  5'd21, 27'h000001bd, 5'd0, 27'h000003c8, 5'd0, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000005b, 5'd3, 27'h000003c6, 5'd13, 27'h000000c8, 32'h00000400,
  1'd1,  5'd24, 27'h000003ec, 5'd1, 27'h0000019a, 5'd22, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b9, 5'd12, 27'h000002c6, 5'd2, 27'h000002db, 32'h00000400,
  1'd1,  5'd24, 27'h00000073, 5'd14, 27'h000003e3, 5'd11, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000004c, 5'd11, 27'h000002e5, 5'd24, 27'h0000036a, 32'h00000400,
  1'd1,  5'd23, 27'h0000030a, 5'd25, 27'h000001d0, 5'd5, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000029d, 5'd21, 27'h0000032d, 5'd14, 27'h0000019c, 32'h00000400,
  1'd1,  5'd21, 27'h000002e9, 5'd21, 27'h00000043, 5'd23, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000004b, 5'd2, 27'h000001cf, 5'd6, 27'h0000001f, 32'h00000400,
  1'd1,  5'd0, 27'h00000159, 5'd0, 27'h00000192, 5'd19, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000100, 5'd3, 27'h00000190, 5'd27, 27'h0000010d, 32'h00000400,
  1'd1,  5'd3, 27'h000000c8, 5'd11, 27'h00000270, 5'd8, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000016c, 5'd10, 27'h000003a4, 5'd17, 27'h0000027e, 32'h00000400,
  1'd1,  5'd2, 27'h0000016c, 5'd12, 27'h000003d8, 5'd30, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000005d, 5'd22, 27'h000002b7, 5'd7, 27'h0000006f, 32'h00000400,
  1'd1,  5'd2, 27'h000002cc, 5'd23, 27'h00000267, 5'd17, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036f, 5'd25, 27'h00000028, 5'd29, 27'h0000016c, 32'h00000400,
  1'd1,  5'd12, 27'h00000003, 5'd2, 27'h0000012a, 5'd7, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001cf, 5'd4, 27'h000003c8, 5'd18, 27'h0000010a, 32'h00000400,
  1'd1,  5'd14, 27'h000002af, 5'd0, 27'h000001ea, 5'd29, 27'h00000071, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001a4, 5'd12, 27'h000003b1, 5'd10, 27'h00000117, 32'h00000400,
  1'd1,  5'd14, 27'h00000283, 5'd12, 27'h0000006f, 5'd18, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000000e, 5'd15, 27'h000000bd, 5'd28, 27'h00000178, 32'h00000400,
  1'd1,  5'd12, 27'h00000210, 5'd24, 27'h000003db, 5'd6, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d4, 5'd23, 27'h000000e4, 5'd18, 27'h0000015a, 32'h00000400,
  1'd1,  5'd13, 27'h0000034e, 5'd23, 27'h0000016a, 5'd30, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003d1, 5'd0, 27'h00000049, 5'd7, 27'h000003c0, 32'h00000400,
  1'd1,  5'd21, 27'h0000011a, 5'd3, 27'h00000178, 5'd16, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000123, 5'd0, 27'h0000026f, 5'd27, 27'h000000ab, 32'h00000400,
  1'd1,  5'd23, 27'h00000055, 5'd14, 27'h000000e2, 5'd5, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000025e, 5'd11, 27'h000000dd, 5'd18, 27'h00000305, 32'h00000400,
  1'd1,  5'd20, 27'h000002d1, 5'd10, 27'h00000388, 5'd29, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000148, 5'd25, 27'h00000200, 5'd9, 27'h0000012d, 32'h00000400,
  1'd1,  5'd22, 27'h000003bc, 5'd23, 27'h000002cf, 5'd19, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000201, 5'd21, 27'h000000ab, 5'd30, 27'h0000011b, 32'h00000400,
  1'd1,  5'd5, 27'h00000051, 5'd7, 27'h000000ea, 5'd4, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e1, 5'd6, 27'h00000362, 5'd12, 27'h0000018d, 32'h00000400,
  1'd1,  5'd0, 27'h00000317, 5'd6, 27'h0000004b, 5'd23, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001e9, 5'd17, 27'h00000164, 5'd4, 27'h000000c0, 32'h00000400,
  1'd1,  5'd4, 27'h000002fa, 5'd16, 27'h00000048, 5'd11, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000bf, 5'd20, 27'h00000185, 5'd24, 27'h00000029, 32'h00000400,
  1'd1,  5'd3, 27'h000002c0, 5'd27, 27'h0000012d, 5'd4, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023e, 5'd28, 27'h0000037a, 5'd12, 27'h00000394, 32'h00000400,
  1'd1,  5'd0, 27'h000003ef, 5'd26, 27'h000003c9, 5'd21, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000006f, 5'd9, 27'h0000012c, 5'd1, 27'h00000152, 32'h00000400,
  1'd1,  5'd11, 27'h000001d7, 5'd9, 27'h000001de, 5'd12, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002b3, 5'd9, 27'h00000312, 5'd23, 27'h000003cc, 32'h00000400,
  1'd1,  5'd11, 27'h00000337, 5'd15, 27'h0000025c, 5'd2, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000198, 5'd16, 27'h0000001d, 5'd12, 27'h0000039c, 32'h00000400,
  1'd1,  5'd14, 27'h00000245, 5'd18, 27'h0000006b, 5'd24, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000016c, 5'd28, 27'h00000086, 5'd2, 27'h000002ec, 32'h00000400,
  1'd1,  5'd15, 27'h00000133, 5'd26, 27'h00000103, 5'd11, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ff, 5'd30, 27'h000002b2, 5'd25, 27'h000002df, 32'h00000400,
  1'd1,  5'd21, 27'h00000212, 5'd5, 27'h0000038a, 5'd0, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002e4, 5'd10, 27'h000000b2, 5'd13, 27'h0000034d, 32'h00000400,
  1'd1,  5'd21, 27'h00000179, 5'd9, 27'h000003a4, 5'd23, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ff, 5'd16, 27'h0000026c, 5'd2, 27'h00000286, 32'h00000400,
  1'd1,  5'd23, 27'h000000f6, 5'd18, 27'h0000003d, 5'd13, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000020d, 5'd20, 27'h00000077, 5'd23, 27'h0000025b, 32'h00000400,
  1'd1,  5'd25, 27'h00000074, 5'd26, 27'h00000176, 5'd2, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000028b, 5'd28, 27'h00000247, 5'd13, 27'h00000106, 32'h00000400,
  1'd1,  5'd22, 27'h00000242, 5'd28, 27'h00000181, 5'd22, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000028e, 5'd6, 27'h00000020, 5'd5, 27'h000003d9, 32'h00000400,
  1'd1,  5'd2, 27'h000000b7, 5'd9, 27'h000002b2, 5'd20, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000292, 5'd6, 27'h00000122, 5'd30, 27'h000003e0, 32'h00000400,
  1'd1,  5'd3, 27'h00000181, 5'd20, 27'h00000139, 5'd6, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f4, 5'd17, 27'h00000088, 5'd19, 27'h0000037c, 32'h00000400,
  1'd1,  5'd3, 27'h000000cd, 5'd20, 27'h0000010e, 5'd29, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000387, 5'd30, 27'h00000247, 5'd6, 27'h00000125, 32'h00000400,
  1'd1,  5'd4, 27'h00000056, 5'd29, 27'h0000009c, 5'd15, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000039d, 5'd27, 27'h000002f1, 5'd29, 27'h00000304, 32'h00000400,
  1'd1,  5'd12, 27'h000003e0, 5'd8, 27'h000002e4, 5'd8, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003a8, 5'd8, 27'h00000286, 5'd16, 27'h00000189, 32'h00000400,
  1'd1,  5'd11, 27'h00000374, 5'd7, 27'h00000108, 5'd29, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000173, 5'd20, 27'h00000047, 5'd7, 27'h00000223, 32'h00000400,
  1'd1,  5'd15, 27'h000000a1, 5'd20, 27'h00000069, 5'd18, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000251, 5'd19, 27'h0000030f, 5'd28, 27'h0000013f, 32'h00000400,
  1'd1,  5'd13, 27'h00000009, 5'd29, 27'h0000002d, 5'd9, 27'h00000187, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003a, 5'd29, 27'h0000006d, 5'd15, 27'h0000035d, 32'h00000400,
  1'd1,  5'd13, 27'h0000008a, 5'd27, 27'h000003de, 5'd26, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000f9, 5'd8, 27'h000002ed, 5'd6, 27'h0000026f, 32'h00000400,
  1'd1,  5'd23, 27'h00000252, 5'd6, 27'h00000061, 5'd16, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000034e, 5'd8, 27'h000002c9, 5'd28, 27'h0000038c, 32'h00000400,
  1'd1,  5'd24, 27'h000003b8, 5'd16, 27'h0000009a, 5'd8, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000116, 5'd19, 27'h000002a9, 5'd20, 27'h000000b4, 32'h00000400,
  1'd1,  5'd21, 27'h000002c8, 5'd16, 27'h0000020d, 5'd28, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000025a, 5'd26, 27'h000001f9, 5'd9, 27'h000002d6, 32'h00000400,
  1'd1,  5'd25, 27'h00000125, 5'd26, 27'h000003b1, 5'd18, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002f6, 5'd29, 27'h00000083, 5'd29, 27'h000001af, 32'h00000400,
  1'd1,  5'd5, 27'h00000319, 5'd3, 27'h000001c6, 5'd5, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003dc, 5'd0, 27'h000001da, 5'd18, 27'h000002ce, 32'h00000400,
  1'd1,  5'd10, 27'h00000113, 5'd0, 27'h0000026d, 5'd25, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000170, 5'd13, 27'h000003fb, 5'd3, 27'h000000c5, 32'h00000400,
  1'd1,  5'd8, 27'h0000012d, 5'd10, 27'h00000208, 5'd12, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000117, 5'd13, 27'h00000162, 5'd21, 27'h000002c2, 32'h00000400,
  1'd1,  5'd5, 27'h000003ff, 5'd22, 27'h0000026b, 5'd4, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000044, 5'd24, 27'h0000016e, 5'd10, 27'h00000226, 32'h00000400,
  1'd1,  5'd8, 27'h00000300, 5'd24, 27'h000002f6, 5'd25, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a7, 5'd3, 27'h00000247, 5'd5, 27'h00000321, 32'h00000400,
  1'd1,  5'd20, 27'h000001da, 5'd3, 27'h00000376, 5'd16, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003bc, 5'd0, 27'h00000190, 5'd27, 27'h000001fd, 32'h00000400,
  1'd1,  5'd17, 27'h00000095, 5'd14, 27'h00000056, 5'd4, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000052, 5'd14, 27'h000002a4, 5'd15, 27'h00000191, 32'h00000400,
  1'd1,  5'd16, 27'h000002d5, 5'd15, 27'h0000001b, 5'd25, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000319, 5'd24, 27'h0000010b, 5'd0, 27'h0000032b, 32'h00000400,
  1'd1,  5'd20, 27'h000000e3, 5'd25, 27'h000001d1, 5'd13, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c0, 5'd25, 27'h00000156, 5'd24, 27'h0000035c, 32'h00000400,
  1'd1,  5'd29, 27'h0000008c, 5'd2, 27'h00000170, 5'd2, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000296, 5'd3, 27'h000000ee, 5'd12, 27'h00000194, 32'h00000400,
  1'd1,  5'd29, 27'h000000ea, 5'd2, 27'h0000015e, 5'd21, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000da, 5'd13, 27'h0000016e, 5'd2, 27'h00000177, 32'h00000400,
  1'd1,  5'd27, 27'h00000008, 5'd13, 27'h000001ab, 5'd13, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000079, 5'd14, 27'h00000252, 5'd20, 27'h00000348, 32'h00000400,
  1'd1,  5'd29, 27'h00000099, 5'd21, 27'h00000122, 5'd4, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000317, 5'd24, 27'h00000143, 5'd10, 27'h000001ef, 32'h00000400,
  1'd1,  5'd29, 27'h0000010e, 5'd23, 27'h00000019, 5'd23, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000003e, 5'd1, 27'h0000037b, 5'd2, 27'h00000026, 32'h00000400,
  1'd1,  5'd10, 27'h000000ff, 5'd2, 27'h00000157, 5'd11, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032b, 5'd4, 27'h00000215, 5'd22, 27'h00000187, 32'h00000400,
  1'd1,  5'd8, 27'h000000fb, 5'd13, 27'h0000030d, 5'd9, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000172, 5'd14, 27'h000002a2, 5'd17, 27'h0000024f, 32'h00000400,
  1'd1,  5'd7, 27'h00000187, 5'd12, 27'h00000229, 5'd30, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003a8, 5'd22, 27'h000003c4, 5'd7, 27'h0000027a, 32'h00000400,
  1'd1,  5'd9, 27'h00000129, 5'd21, 27'h0000003a, 5'd18, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000220, 5'd24, 27'h000000b6, 5'd30, 27'h00000107, 32'h00000400,
  1'd1,  5'd18, 27'h000002e1, 5'd1, 27'h000003de, 5'd1, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000219, 5'd3, 27'h000003ba, 5'd10, 27'h000001c3, 32'h00000400,
  1'd1,  5'd17, 27'h00000345, 5'd4, 27'h000001e2, 5'd25, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000022e, 5'd11, 27'h00000087, 5'd7, 27'h00000120, 32'h00000400,
  1'd1,  5'd19, 27'h000002c8, 5'd10, 27'h000003ae, 5'd15, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000212, 5'd11, 27'h000002c1, 5'd26, 27'h00000034, 32'h00000400,
  1'd1,  5'd19, 27'h000000f1, 5'd24, 27'h00000150, 5'd6, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000175, 5'd22, 27'h000000ce, 5'd15, 27'h00000245, 32'h00000400,
  1'd1,  5'd16, 27'h00000109, 5'd24, 27'h00000309, 5'd30, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b1, 5'd3, 27'h000001a7, 5'd9, 27'h0000000b, 32'h00000400,
  1'd1,  5'd26, 27'h000002f5, 5'd4, 27'h0000039e, 5'd20, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000148, 5'd4, 27'h000000a1, 5'd26, 27'h000000b5, 32'h00000400,
  1'd1,  5'd26, 27'h00000246, 5'd11, 27'h000001ce, 5'd9, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000000b, 5'd11, 27'h000001f6, 5'd16, 27'h000001b2, 32'h00000400,
  1'd1,  5'd26, 27'h000003f1, 5'd11, 27'h000003e3, 5'd29, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000012d, 5'd22, 27'h000001a0, 5'd9, 27'h00000366, 32'h00000400,
  1'd1,  5'd26, 27'h00000144, 5'd25, 27'h00000090, 5'd18, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000036, 5'd23, 27'h000003c0, 5'd29, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h0000004f, 5'd9, 27'h000002cf, 5'd1, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ef, 5'd7, 27'h000003e2, 5'd10, 27'h00000360, 32'h00000400,
  1'd1,  5'd10, 27'h0000006c, 5'd5, 27'h00000254, 5'd24, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000031, 5'd15, 27'h00000329, 5'd0, 27'h000001bd, 32'h00000400,
  1'd1,  5'd8, 27'h000003db, 5'd16, 27'h0000022c, 5'd14, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000019e, 5'd20, 27'h000001fb, 5'd20, 27'h000002f7, 32'h00000400,
  1'd1,  5'd5, 27'h000000c9, 5'd30, 27'h0000010f, 5'd4, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000136, 5'd29, 27'h00000009, 5'd11, 27'h00000291, 32'h00000400,
  1'd1,  5'd7, 27'h000003bf, 5'd30, 27'h0000008a, 5'd23, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002fb, 5'd9, 27'h00000030, 5'd4, 27'h0000025c, 32'h00000400,
  1'd1,  5'd15, 27'h000002f2, 5'd7, 27'h00000215, 5'd11, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031c, 5'd10, 27'h000000bb, 5'd23, 27'h000001c4, 32'h00000400,
  1'd1,  5'd20, 27'h000001d9, 5'd16, 27'h000003f1, 5'd3, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000371, 5'd17, 27'h00000113, 5'd12, 27'h000003cd, 32'h00000400,
  1'd1,  5'd18, 27'h0000006a, 5'd16, 27'h00000119, 5'd22, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f6, 5'd29, 27'h00000078, 5'd3, 27'h000002b5, 32'h00000400,
  1'd1,  5'd17, 27'h0000034e, 5'd27, 27'h00000231, 5'd12, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000185, 5'd30, 27'h000002cb, 5'd21, 27'h00000274, 32'h00000400,
  1'd1,  5'd30, 27'h00000064, 5'd8, 27'h000001d3, 5'd4, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000377, 5'd5, 27'h00000115, 5'd11, 27'h00000175, 32'h00000400,
  1'd1,  5'd30, 27'h000002d5, 5'd10, 27'h00000113, 5'd22, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001bb, 5'd16, 27'h00000303, 5'd0, 27'h00000212, 32'h00000400,
  1'd1,  5'd29, 27'h00000040, 5'd20, 27'h00000244, 5'd14, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e6, 5'd16, 27'h0000021a, 5'd23, 27'h0000008b, 32'h00000400,
  1'd1,  5'd26, 27'h000000ef, 5'd28, 27'h00000169, 5'd0, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d5, 5'd30, 27'h000002df, 5'd12, 27'h00000127, 32'h00000400,
  1'd1,  5'd26, 27'h0000037a, 5'd29, 27'h000003b1, 5'd23, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000197, 5'd10, 27'h0000014b, 5'd10, 27'h0000006f, 32'h00000400,
  1'd1,  5'd6, 27'h0000024e, 5'd5, 27'h000002a1, 5'd19, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002db, 5'd7, 27'h00000317, 5'd30, 27'h00000110, 32'h00000400,
  1'd1,  5'd8, 27'h0000024e, 5'd20, 27'h00000128, 5'd6, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000221, 5'd18, 27'h00000156, 5'd17, 27'h00000061, 32'h00000400,
  1'd1,  5'd8, 27'h0000002e, 5'd18, 27'h0000016e, 5'd30, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000287, 5'd29, 27'h000000cb, 5'd9, 27'h000002f3, 32'h00000400,
  1'd1,  5'd6, 27'h00000209, 5'd28, 27'h000002f9, 5'd16, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000217, 5'd30, 27'h00000168, 5'd26, 27'h0000023f, 32'h00000400,
  1'd1,  5'd18, 27'h0000005e, 5'd6, 27'h0000023a, 5'd8, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000266, 5'd7, 27'h000000cd, 5'd19, 27'h000000e3, 32'h00000400,
  1'd1,  5'd19, 27'h0000039f, 5'd8, 27'h00000275, 5'd26, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000024, 5'd19, 27'h00000126, 5'd9, 27'h00000191, 32'h00000400,
  1'd1,  5'd16, 27'h0000002d, 5'd15, 27'h000003f2, 5'd15, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000200, 5'd19, 27'h0000038d, 5'd28, 27'h00000181, 32'h00000400,
  1'd1,  5'd17, 27'h0000035b, 5'd29, 27'h0000017b, 5'd6, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003fd, 5'd26, 27'h00000214, 5'd19, 27'h00000128, 32'h00000400,
  1'd1,  5'd19, 27'h00000034, 5'd30, 27'h000001f9, 5'd26, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000290, 5'd5, 27'h0000035a, 5'd9, 27'h000002a8, 32'h00000400,
  1'd1,  5'd26, 27'h00000089, 5'd5, 27'h0000013e, 5'd18, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a7, 5'd7, 27'h000002d7, 5'd26, 27'h000003a1, 32'h00000400,
  1'd1,  5'd26, 27'h0000035a, 5'd15, 27'h00000339, 5'd7, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000213, 5'd19, 27'h00000384, 5'd19, 27'h0000019e, 32'h00000400,
  1'd1,  5'd30, 27'h0000025a, 5'd18, 27'h000000f4, 5'd26, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000026, 5'd26, 27'h000001e9, 5'd9, 27'h000001d4, 32'h00000400,
  1'd1,  5'd25, 27'h000003a9, 5'd28, 27'h0000033a, 5'd19, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c5, 5'd28, 27'h0000030b, 5'd28, 27'h000002aa, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000209, 5'd4, 27'h00000092, 5'd1, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000092, 5'd0, 27'h0000017f, 5'd11, 27'h000003dd, 32'h00000400,
  1'd1,  5'd4, 27'h000000c6, 5'd3, 27'h000001ac, 5'd22, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000024d, 5'd14, 27'h0000012a, 5'd4, 27'h0000005b, 32'h00000400,
  1'd1,  5'd0, 27'h00000331, 5'd11, 27'h000002c0, 5'd12, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ce, 5'd14, 27'h0000018c, 5'd22, 27'h000003cd, 32'h00000400,
  1'd1,  5'd3, 27'h0000014f, 5'd24, 27'h000001a4, 5'd2, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000243, 5'd21, 27'h000003f0, 5'd13, 27'h00000360, 32'h00000400,
  1'd1,  5'd2, 27'h0000009b, 5'd24, 27'h000001e1, 5'd20, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002eb, 5'd3, 27'h0000017e, 5'd3, 27'h00000392, 32'h00000400,
  1'd1,  5'd14, 27'h00000276, 5'd0, 27'h00000225, 5'd11, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000241, 5'd2, 27'h0000030f, 5'd25, 27'h00000058, 32'h00000400,
  1'd1,  5'd12, 27'h000003f2, 5'd13, 27'h000003f9, 5'd0, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000323, 5'd12, 27'h00000055, 5'd13, 27'h000001b9, 32'h00000400,
  1'd1,  5'd13, 27'h00000133, 5'd13, 27'h000002d9, 5'd25, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031c, 5'd24, 27'h00000028, 5'd0, 27'h00000348, 32'h00000400,
  1'd1,  5'd14, 27'h0000022e, 5'd22, 27'h000003fe, 5'd15, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e0, 5'd23, 27'h0000013b, 5'd22, 27'h00000216, 32'h00000400,
  1'd1,  5'd25, 27'h000002ea, 5'd2, 27'h00000016, 5'd3, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000039c, 5'd0, 27'h00000021, 5'd12, 27'h000002cd, 32'h00000400,
  1'd1,  5'd22, 27'h00000330, 5'd3, 27'h000001b3, 5'd23, 27'h000001f3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000003d, 5'd14, 27'h0000034c, 5'd3, 27'h000000d4, 32'h00000400,
  1'd1,  5'd23, 27'h00000163, 5'd11, 27'h000001d5, 5'd11, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000b8, 5'd12, 27'h0000014d, 5'd21, 27'h000002e7, 32'h00000400,
  1'd1,  5'd25, 27'h000001ad, 5'd23, 27'h00000103, 5'd0, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002dc, 5'd24, 27'h0000012a, 5'd15, 27'h000001d6, 32'h00000400,
  1'd1,  5'd24, 27'h000000e0, 5'd23, 27'h0000019c, 5'd20, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000d2, 5'd0, 27'h00000176, 5'd8, 27'h000002f8, 32'h00000400,
  1'd1,  5'd0, 27'h00000207, 5'd2, 27'h00000016, 5'd20, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000191, 5'd2, 27'h000000b1, 5'd27, 27'h0000030b, 32'h00000400,
  1'd1,  5'd1, 27'h0000002d, 5'd12, 27'h00000016, 5'd6, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f5, 5'd13, 27'h000002f6, 5'd15, 27'h000002cd, 32'h00000400,
  1'd1,  5'd4, 27'h000003ac, 5'd13, 27'h00000376, 5'd29, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000035d, 5'd20, 27'h0000033f, 5'd9, 27'h0000037f, 32'h00000400,
  1'd1,  5'd2, 27'h000003ca, 5'd25, 27'h00000046, 5'd18, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000398, 5'd23, 27'h00000253, 5'd28, 27'h000002d2, 32'h00000400,
  1'd1,  5'd14, 27'h00000216, 5'd4, 27'h000002cc, 5'd6, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000005d, 5'd3, 27'h0000001b, 5'd16, 27'h0000013f, 32'h00000400,
  1'd1,  5'd15, 27'h0000011e, 5'd1, 27'h000001a8, 5'd27, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000035c, 5'd11, 27'h00000252, 5'd6, 27'h00000359, 32'h00000400,
  1'd1,  5'd14, 27'h00000155, 5'd14, 27'h000001bb, 5'd18, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e7, 5'd14, 27'h00000118, 5'd29, 27'h0000018a, 32'h00000400,
  1'd1,  5'd10, 27'h00000171, 5'd21, 27'h000000a4, 5'd6, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000070, 5'd21, 27'h000000b4, 5'd19, 27'h0000026c, 32'h00000400,
  1'd1,  5'd13, 27'h00000324, 5'd23, 27'h00000028, 5'd27, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003fd, 5'd1, 27'h00000047, 5'd6, 27'h00000294, 32'h00000400,
  1'd1,  5'd21, 27'h000000bf, 5'd3, 27'h00000161, 5'd18, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000398, 5'd2, 27'h0000024d, 5'd27, 27'h00000061, 32'h00000400,
  1'd1,  5'd25, 27'h0000016a, 5'd14, 27'h00000119, 5'd8, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000b6, 5'd10, 27'h00000295, 5'd16, 27'h000001c0, 32'h00000400,
  1'd1,  5'd21, 27'h000003ec, 5'd11, 27'h000001e9, 5'd27, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000303, 5'd24, 27'h00000165, 5'd7, 27'h00000119, 32'h00000400,
  1'd1,  5'd20, 27'h000003c3, 5'd23, 27'h00000198, 5'd15, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001e8, 5'd20, 27'h00000354, 5'd27, 27'h00000206, 32'h00000400,
  1'd1,  5'd1, 27'h00000031, 5'd10, 27'h00000141, 5'd4, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000a1, 5'd5, 27'h000003bd, 5'd10, 27'h0000028e, 32'h00000400,
  1'd1,  5'd3, 27'h000001f9, 5'd9, 27'h00000329, 5'd25, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000d5, 5'd17, 27'h000002f4, 5'd4, 27'h00000121, 32'h00000400,
  1'd1,  5'd3, 27'h00000212, 5'd19, 27'h00000053, 5'd15, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000043, 5'd19, 27'h00000017, 5'd20, 27'h00000376, 32'h00000400,
  1'd1,  5'd1, 27'h00000329, 5'd27, 27'h000000af, 5'd1, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020a, 5'd26, 27'h00000007, 5'd11, 27'h00000334, 32'h00000400,
  1'd1,  5'd1, 27'h000003a1, 5'd26, 27'h000002f4, 5'd23, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002cf, 5'd8, 27'h000001a2, 5'd5, 27'h00000056, 32'h00000400,
  1'd1,  5'd12, 27'h000001ff, 5'd6, 27'h0000018e, 5'd11, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000151, 5'd8, 27'h000000d6, 5'd21, 27'h00000137, 32'h00000400,
  1'd1,  5'd10, 27'h00000208, 5'd19, 27'h000001dc, 5'd1, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001ba, 5'd19, 27'h000000c5, 5'd10, 27'h000001a7, 32'h00000400,
  1'd1,  5'd14, 27'h000001fa, 5'd17, 27'h000003db, 5'd22, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001f4, 5'd28, 27'h000002f5, 5'd0, 27'h00000386, 32'h00000400,
  1'd1,  5'd11, 27'h000003f0, 5'd29, 27'h000002c0, 5'd14, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000081, 5'd30, 27'h0000000b, 5'd23, 27'h000001ad, 32'h00000400,
  1'd1,  5'd25, 27'h00000036, 5'd6, 27'h0000037e, 5'd1, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000031b, 5'd10, 27'h000000fc, 5'd10, 27'h000003d9, 32'h00000400,
  1'd1,  5'd20, 27'h0000033a, 5'd7, 27'h0000002e, 5'd25, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f1, 5'd15, 27'h000002ff, 5'd4, 27'h000002e6, 32'h00000400,
  1'd1,  5'd22, 27'h0000006f, 5'd17, 27'h000000ef, 5'd10, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000147, 5'd18, 27'h000003bc, 5'd23, 27'h000002f7, 32'h00000400,
  1'd1,  5'd23, 27'h000003dd, 5'd30, 27'h0000031e, 5'd4, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002f8, 5'd26, 27'h00000039, 5'd13, 27'h00000279, 32'h00000400,
  1'd1,  5'd23, 27'h00000351, 5'd26, 27'h0000001c, 5'd21, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ef, 5'd6, 27'h000002ff, 5'd7, 27'h0000002c, 32'h00000400,
  1'd1,  5'd4, 27'h0000034c, 5'd6, 27'h0000027e, 5'd18, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000215, 5'd7, 27'h000003f3, 5'd29, 27'h000003fa, 32'h00000400,
  1'd1,  5'd5, 27'h0000004d, 5'd18, 27'h0000013c, 5'd9, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000026a, 5'd19, 27'h0000017a, 5'd18, 27'h0000002b, 32'h00000400,
  1'd1,  5'd1, 27'h00000235, 5'd20, 27'h00000121, 5'd30, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000363, 5'd30, 27'h00000324, 5'd9, 27'h00000377, 32'h00000400,
  1'd1,  5'd1, 27'h000000cf, 5'd29, 27'h0000030f, 5'd19, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000037a, 5'd27, 27'h00000274, 5'd26, 27'h0000027a, 32'h00000400,
  1'd1,  5'd11, 27'h0000023e, 5'd8, 27'h0000021d, 5'd10, 27'h000000f3, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017d, 5'd8, 27'h0000033a, 5'd17, 27'h0000008f, 32'h00000400,
  1'd1,  5'd11, 27'h000003dd, 5'd8, 27'h00000157, 5'd30, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001da, 5'd16, 27'h000002bb, 5'd8, 27'h0000036d, 32'h00000400,
  1'd1,  5'd10, 27'h000003a6, 5'd17, 27'h00000366, 5'd18, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ce, 5'd18, 27'h00000005, 5'd30, 27'h00000068, 32'h00000400,
  1'd1,  5'd15, 27'h00000006, 5'd28, 27'h0000019e, 5'd8, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d4, 5'd27, 27'h000002b1, 5'd20, 27'h000000d2, 32'h00000400,
  1'd1,  5'd15, 27'h0000005a, 5'd27, 27'h00000327, 5'd25, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001fd, 5'd8, 27'h00000307, 5'd7, 27'h00000019, 32'h00000400,
  1'd1,  5'd21, 27'h000003e0, 5'd9, 27'h000000bf, 5'd17, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000e8, 5'd6, 27'h00000089, 5'd28, 27'h0000011f, 32'h00000400,
  1'd1,  5'd24, 27'h000000d8, 5'd18, 27'h00000156, 5'd5, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000165, 5'd20, 27'h000000fa, 5'd20, 27'h00000101, 32'h00000400,
  1'd1,  5'd24, 27'h000000df, 5'd16, 27'h000000fe, 5'd29, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000170, 5'd30, 27'h000003c9, 5'd9, 27'h000002ef, 32'h00000400,
  1'd1,  5'd21, 27'h000002a0, 5'd28, 27'h0000033b, 5'd20, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001de, 5'd28, 27'h00000282, 5'd28, 27'h0000001d, 32'h00000400,
  1'd1,  5'd5, 27'h00000274, 5'd0, 27'h00000342, 5'd6, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012b, 5'd2, 27'h00000164, 5'd19, 27'h00000156, 32'h00000400,
  1'd1,  5'd6, 27'h000000ee, 5'd2, 27'h00000066, 5'd26, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000090, 5'd15, 27'h000000ac, 5'd1, 27'h00000067, 32'h00000400,
  1'd1,  5'd5, 27'h000003fd, 5'd15, 27'h000000ba, 5'd14, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000352, 5'd14, 27'h00000350, 5'd25, 27'h000000ab, 32'h00000400,
  1'd1,  5'd5, 27'h00000364, 5'd24, 27'h000000b2, 5'd2, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d7, 5'd23, 27'h000003a8, 5'd11, 27'h0000039c, 32'h00000400,
  1'd1,  5'd10, 27'h000000a3, 5'd25, 27'h000001eb, 5'd25, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c2, 5'd3, 27'h000001ec, 5'd7, 27'h000002b3, 32'h00000400,
  1'd1,  5'd19, 27'h00000399, 5'd2, 27'h00000311, 5'd20, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000290, 5'd2, 27'h0000030c, 5'd27, 27'h0000009e, 32'h00000400,
  1'd1,  5'd19, 27'h0000001b, 5'd13, 27'h000002c1, 5'd3, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c9, 5'd12, 27'h00000298, 5'd11, 27'h0000003f, 32'h00000400,
  1'd1,  5'd15, 27'h00000343, 5'd11, 27'h0000015f, 5'd22, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000110, 5'd25, 27'h000000a2, 5'd1, 27'h0000013b, 32'h00000400,
  1'd1,  5'd19, 27'h00000287, 5'd22, 27'h0000013a, 5'd12, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000062, 5'd24, 27'h000001e8, 5'd20, 27'h00000394, 32'h00000400,
  1'd1,  5'd27, 27'h000003de, 5'd1, 27'h00000116, 5'd4, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c0, 5'd2, 27'h0000021d, 5'd13, 27'h00000113, 32'h00000400,
  1'd1,  5'd26, 27'h000003f7, 5'd3, 27'h00000294, 5'd22, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000030f, 5'd12, 27'h000000b3, 5'd2, 27'h00000392, 32'h00000400,
  1'd1,  5'd29, 27'h00000216, 5'd15, 27'h000000a8, 5'd13, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003a5, 5'd11, 27'h000002b6, 5'd20, 27'h00000398, 32'h00000400,
  1'd1,  5'd28, 27'h0000016e, 5'd23, 27'h000001dc, 5'd4, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000016d, 5'd21, 27'h000003e3, 5'd14, 27'h00000152, 32'h00000400,
  1'd1,  5'd26, 27'h00000123, 5'd21, 27'h000002ca, 5'd24, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000003b, 5'd2, 27'h000000d6, 5'd1, 27'h000002b8, 32'h00000400,
  1'd1,  5'd9, 27'h000001c9, 5'd2, 27'h00000082, 5'd14, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000324, 5'd0, 27'h000000ea, 5'd24, 27'h00000018, 32'h00000400,
  1'd1,  5'd5, 27'h000002ce, 5'd13, 27'h000002df, 5'd9, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000cf, 5'd12, 27'h00000218, 5'd19, 27'h00000141, 32'h00000400,
  1'd1,  5'd9, 27'h000003ed, 5'd12, 27'h0000039e, 5'd28, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000184, 5'd21, 27'h00000339, 5'd7, 27'h0000004f, 32'h00000400,
  1'd1,  5'd9, 27'h000003a9, 5'd21, 27'h00000046, 5'd19, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000019d, 5'd23, 27'h000001eb, 5'd30, 27'h0000010a, 32'h00000400,
  1'd1,  5'd16, 27'h000003f9, 5'd5, 27'h0000003b, 5'd1, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000371, 5'd3, 27'h0000007b, 5'd12, 27'h0000029f, 32'h00000400,
  1'd1,  5'd19, 27'h000000dc, 5'd3, 27'h0000038a, 5'd21, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002cf, 5'd10, 27'h000002b8, 5'd6, 27'h000001d3, 32'h00000400,
  1'd1,  5'd17, 27'h000001f9, 5'd15, 27'h00000024, 5'd16, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000395, 5'd11, 27'h00000341, 5'd28, 27'h00000075, 32'h00000400,
  1'd1,  5'd17, 27'h0000009c, 5'd20, 27'h000003d7, 5'd6, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000371, 5'd24, 27'h0000023c, 5'd16, 27'h0000007d, 32'h00000400,
  1'd1,  5'd16, 27'h0000004a, 5'd23, 27'h00000208, 5'd30, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000094, 5'd1, 27'h00000052, 5'd5, 27'h0000021a, 32'h00000400,
  1'd1,  5'd29, 27'h000003bc, 5'd4, 27'h00000058, 5'd15, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002d9, 5'd1, 27'h000000e1, 5'd28, 27'h000002b8, 32'h00000400,
  1'd1,  5'd25, 27'h000003fb, 5'd12, 27'h000000e6, 5'd9, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002ac, 5'd15, 27'h00000164, 5'd18, 27'h000000d3, 32'h00000400,
  1'd1,  5'd28, 27'h00000085, 5'd14, 27'h00000234, 5'd27, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000010c, 5'd22, 27'h000003e7, 5'd6, 27'h0000012c, 32'h00000400,
  1'd1,  5'd26, 27'h00000254, 5'd22, 27'h0000034c, 5'd15, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000248, 5'd23, 27'h0000034c, 5'd26, 27'h00000264, 32'h00000400,
  1'd1,  5'd5, 27'h000003ee, 5'd7, 27'h0000016a, 5'd4, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003dd, 5'd8, 27'h00000061, 5'd11, 27'h000003d9, 32'h00000400,
  1'd1,  5'd6, 27'h00000065, 5'd6, 27'h00000296, 5'd21, 27'h0000002d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000294, 5'd18, 27'h00000081, 5'd5, 27'h00000019, 32'h00000400,
  1'd1,  5'd10, 27'h00000101, 5'd17, 27'h0000004c, 5'd14, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c4, 5'd16, 27'h000000ae, 5'd25, 27'h0000005d, 32'h00000400,
  1'd1,  5'd8, 27'h0000023a, 5'd25, 27'h000003f5, 5'd3, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000006a, 5'd30, 27'h000002e7, 5'd11, 27'h0000008e, 32'h00000400,
  1'd1,  5'd8, 27'h000003da, 5'd26, 27'h00000229, 5'd22, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000086, 5'd8, 27'h0000021b, 5'd1, 27'h000001da, 32'h00000400,
  1'd1,  5'd18, 27'h00000382, 5'd5, 27'h000000ea, 5'd15, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001bf, 5'd5, 27'h000003ad, 5'd21, 27'h000003ef, 32'h00000400,
  1'd1,  5'd20, 27'h000001d9, 5'd18, 27'h0000031a, 5'd3, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002f3, 5'd16, 27'h00000051, 5'd14, 27'h000000ed, 32'h00000400,
  1'd1,  5'd20, 27'h00000292, 5'd18, 27'h00000324, 5'd22, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000236, 5'd29, 27'h0000015f, 5'd0, 27'h000001a1, 32'h00000400,
  1'd1,  5'd16, 27'h0000015e, 5'd30, 27'h000000b9, 5'd15, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000000e, 5'd30, 27'h00000103, 5'd20, 27'h00000384, 32'h00000400,
  1'd1,  5'd29, 27'h00000041, 5'd6, 27'h0000008a, 5'd5, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000386, 5'd6, 27'h000002a7, 5'd10, 27'h000003a0, 32'h00000400,
  1'd1,  5'd29, 27'h000001f7, 5'd9, 27'h000001c5, 5'd20, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000151, 5'd16, 27'h00000305, 5'd3, 27'h000000c6, 32'h00000400,
  1'd1,  5'd29, 27'h000000a3, 5'd18, 27'h000003e8, 5'd10, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000165, 5'd15, 27'h000003f0, 5'd23, 27'h00000384, 32'h00000400,
  1'd1,  5'd29, 27'h000000e5, 5'd26, 27'h00000252, 5'd2, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000200, 5'd29, 27'h00000243, 5'd10, 27'h000003a1, 32'h00000400,
  1'd1,  5'd30, 27'h000000de, 5'd28, 27'h00000284, 5'd21, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000102, 5'd7, 27'h00000102, 5'd8, 27'h00000347, 32'h00000400,
  1'd1,  5'd6, 27'h000002a6, 5'd5, 27'h000002df, 5'd17, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e4, 5'd9, 27'h000001c6, 5'd29, 27'h000000d5, 32'h00000400,
  1'd1,  5'd5, 27'h00000207, 5'd17, 27'h00000077, 5'd10, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000079, 5'd16, 27'h000003be, 5'd16, 27'h0000032a, 32'h00000400,
  1'd1,  5'd7, 27'h00000293, 5'd20, 27'h000001df, 5'd30, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000013a, 5'd28, 27'h000001ba, 5'd6, 27'h000000d2, 32'h00000400,
  1'd1,  5'd8, 27'h00000239, 5'd30, 27'h00000159, 5'd18, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000cf, 5'd30, 27'h000003fe, 5'd30, 27'h000003a0, 32'h00000400,
  1'd1,  5'd16, 27'h000001d7, 5'd8, 27'h000001a1, 5'd8, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000bc, 5'd5, 27'h000003c0, 5'd15, 27'h00000277, 32'h00000400,
  1'd1,  5'd19, 27'h000001e2, 5'd5, 27'h0000018f, 5'd30, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000258, 5'd18, 27'h000001e9, 5'd5, 27'h000002b2, 32'h00000400,
  1'd1,  5'd19, 27'h000000f6, 5'd19, 27'h000001fe, 5'd16, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001b3, 5'd16, 27'h0000034b, 5'd26, 27'h000001fa, 32'h00000400,
  1'd1,  5'd18, 27'h000003b2, 5'd27, 27'h0000034a, 5'd9, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e0, 5'd27, 27'h000002b6, 5'd15, 27'h000003cb, 32'h00000400,
  1'd1,  5'd18, 27'h00000185, 5'd26, 27'h00000016, 5'd28, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000097, 5'd7, 27'h00000248, 5'd9, 27'h00000288, 32'h00000400,
  1'd1,  5'd28, 27'h00000389, 5'd5, 27'h000002f3, 5'd18, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002e7, 5'd9, 27'h00000162, 5'd29, 27'h000000bb, 32'h00000400,
  1'd1,  5'd26, 27'h00000028, 5'd19, 27'h00000111, 5'd8, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003fd, 5'd15, 27'h000002e3, 5'd17, 27'h0000028f, 32'h00000400,
  1'd1,  5'd29, 27'h00000146, 5'd16, 27'h00000006, 5'd30, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000102, 5'd25, 27'h0000038d, 5'd8, 27'h000003b2, 32'h00000400,
  1'd1,  5'd28, 27'h00000297, 5'd29, 27'h000002cd, 5'd15, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000361, 5'd30, 27'h000001b1, 5'd27, 27'h0000021f, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000001d3, 5'd0, 27'h000002ac, 5'd1, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000fb, 5'd4, 27'h0000029d, 5'd13, 27'h000002fb, 32'h00000400,
  1'd1,  5'd2, 27'h00000044, 5'd1, 27'h00000392, 5'd25, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000114, 5'd14, 27'h00000282, 5'd0, 27'h000000b8, 32'h00000400,
  1'd1,  5'd1, 27'h000003ee, 5'd11, 27'h000002d6, 5'd14, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001bb, 5'd10, 27'h000002b1, 5'd24, 27'h00000390, 32'h00000400,
  1'd1,  5'd2, 27'h000002fe, 5'd23, 27'h0000023e, 5'd3, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000293, 5'd23, 27'h000003a4, 5'd14, 27'h00000342, 32'h00000400,
  1'd1,  5'd0, 27'h000003d3, 5'd23, 27'h00000246, 5'd21, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000097, 5'd3, 27'h0000031f, 5'd2, 27'h000003e7, 32'h00000400,
  1'd1,  5'd13, 27'h0000013e, 5'd4, 27'h0000006c, 5'd11, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b0, 5'd3, 27'h00000143, 5'd25, 27'h000001c2, 32'h00000400,
  1'd1,  5'd13, 27'h000001ba, 5'd15, 27'h00000110, 5'd3, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000014c, 5'd14, 27'h0000039d, 5'd10, 27'h000002a3, 32'h00000400,
  1'd1,  5'd11, 27'h0000016f, 5'd13, 27'h00000294, 5'd22, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000109, 5'd25, 27'h00000071, 5'd2, 27'h000003eb, 32'h00000400,
  1'd1,  5'd10, 27'h000002bb, 5'd21, 27'h0000012e, 5'd11, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000027a, 5'd20, 27'h000003de, 5'd21, 27'h00000389, 32'h00000400,
  1'd1,  5'd22, 27'h000002e1, 5'd4, 27'h000001d2, 5'd3, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003b0, 5'd4, 27'h0000038e, 5'd13, 27'h0000012c, 32'h00000400,
  1'd1,  5'd24, 27'h00000182, 5'd1, 27'h0000008c, 5'd21, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000018, 5'd14, 27'h0000031f, 5'd3, 27'h000002b5, 32'h00000400,
  1'd1,  5'd23, 27'h0000007d, 5'd10, 27'h000001ed, 5'd12, 27'h0000006f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002f3, 5'd12, 27'h0000018f, 5'd23, 27'h0000009e, 32'h00000400,
  1'd1,  5'd21, 27'h0000019f, 5'd22, 27'h00000110, 5'd1, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000208, 5'd25, 27'h0000028e, 5'd12, 27'h00000400, 32'h00000400,
  1'd1,  5'd25, 27'h000000f9, 5'd22, 27'h00000254, 5'd23, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000341, 5'd1, 27'h00000301, 5'd7, 27'h00000200, 32'h00000400,
  1'd1,  5'd2, 27'h0000034d, 5'd0, 27'h00000391, 5'd18, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000016a, 5'd4, 27'h00000352, 5'd29, 27'h0000030b, 32'h00000400,
  1'd1,  5'd0, 27'h00000331, 5'd12, 27'h00000333, 5'd9, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000399, 5'd14, 27'h0000039a, 5'd19, 27'h000003bd, 32'h00000400,
  1'd1,  5'd0, 27'h0000019c, 5'd14, 27'h00000259, 5'd26, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000220, 5'd21, 27'h00000178, 5'd9, 27'h0000008e, 32'h00000400,
  1'd1,  5'd2, 27'h000001ef, 5'd24, 27'h00000269, 5'd18, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001c7, 5'd24, 27'h0000038b, 5'd27, 27'h000002b6, 32'h00000400,
  1'd1,  5'd11, 27'h00000265, 5'd5, 27'h0000008c, 5'd9, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000095, 5'd2, 27'h00000317, 5'd17, 27'h00000180, 32'h00000400,
  1'd1,  5'd15, 27'h00000075, 5'd1, 27'h000003c0, 5'd28, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000298, 5'd11, 27'h00000305, 5'd8, 27'h0000008a, 32'h00000400,
  1'd1,  5'd13, 27'h000002d1, 5'd12, 27'h0000006e, 5'd20, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f0, 5'd13, 27'h00000321, 5'd26, 27'h000002c7, 32'h00000400,
  1'd1,  5'd14, 27'h000001d8, 5'd21, 27'h00000128, 5'd6, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d5, 5'd20, 27'h000002e8, 5'd20, 27'h00000117, 32'h00000400,
  1'd1,  5'd14, 27'h0000010f, 5'd24, 27'h00000223, 5'd30, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000074, 5'd4, 27'h00000390, 5'd10, 27'h00000073, 32'h00000400,
  1'd1,  5'd25, 27'h00000169, 5'd0, 27'h00000252, 5'd19, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ac, 5'd0, 27'h0000030c, 5'd29, 27'h0000033c, 32'h00000400,
  1'd1,  5'd20, 27'h000002cc, 5'd11, 27'h00000331, 5'd6, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000182, 5'd12, 27'h0000021a, 5'd16, 27'h00000130, 32'h00000400,
  1'd1,  5'd24, 27'h00000206, 5'd14, 27'h000000f6, 5'd29, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b1, 5'd21, 27'h000003eb, 5'd5, 27'h00000393, 32'h00000400,
  1'd1,  5'd25, 27'h000001af, 5'd25, 27'h00000009, 5'd20, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000cd, 5'd25, 27'h000001d4, 5'd27, 27'h00000020, 32'h00000400,
  1'd1,  5'd1, 27'h00000286, 5'd6, 27'h00000390, 5'd0, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000250, 5'd5, 27'h000002f1, 5'd13, 27'h00000376, 32'h00000400,
  1'd1,  5'd3, 27'h0000021e, 5'd5, 27'h000001ff, 5'd25, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000378, 5'd16, 27'h0000028d, 5'd4, 27'h00000081, 32'h00000400,
  1'd1,  5'd4, 27'h000002d5, 5'd15, 27'h00000393, 5'd12, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002b3, 5'd19, 27'h000003ee, 5'd21, 27'h0000011e, 32'h00000400,
  1'd1,  5'd2, 27'h00000141, 5'd29, 27'h0000017e, 5'd1, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002fb, 5'd30, 27'h00000014, 5'd15, 27'h000001be, 32'h00000400,
  1'd1,  5'd2, 27'h000002a1, 5'd28, 27'h0000020a, 5'd25, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000181, 5'd8, 27'h00000245, 5'd2, 27'h00000276, 32'h00000400,
  1'd1,  5'd13, 27'h000003a3, 5'd9, 27'h000001f4, 5'd13, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000032d, 5'd6, 27'h0000030f, 5'd23, 27'h00000312, 32'h00000400,
  1'd1,  5'd13, 27'h00000041, 5'd18, 27'h00000096, 5'd0, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000b7, 5'd18, 27'h000000e5, 5'd11, 27'h000002ff, 32'h00000400,
  1'd1,  5'd12, 27'h00000355, 5'd16, 27'h00000122, 5'd21, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000392, 5'd27, 27'h000002cc, 5'd2, 27'h000003ea, 32'h00000400,
  1'd1,  5'd11, 27'h00000019, 5'd26, 27'h00000227, 5'd11, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001b7, 5'd30, 27'h000002c0, 5'd25, 27'h00000090, 32'h00000400,
  1'd1,  5'd21, 27'h0000006c, 5'd6, 27'h000002b7, 5'd2, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001a4, 5'd8, 27'h00000019, 5'd12, 27'h00000061, 32'h00000400,
  1'd1,  5'd24, 27'h00000313, 5'd7, 27'h00000068, 5'd21, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000036, 5'd16, 27'h000000a0, 5'd0, 27'h00000055, 32'h00000400,
  1'd1,  5'd24, 27'h0000019d, 5'd19, 27'h00000194, 5'd14, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000139, 5'd19, 27'h000003a8, 5'd20, 27'h00000371, 32'h00000400,
  1'd1,  5'd23, 27'h00000372, 5'd29, 27'h0000003b, 5'd1, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000364, 5'd28, 27'h00000389, 5'd12, 27'h000001db, 32'h00000400,
  1'd1,  5'd23, 27'h00000154, 5'd28, 27'h000002d4, 5'd23, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000286, 5'd7, 27'h000002ca, 5'd5, 27'h00000155, 32'h00000400,
  1'd1,  5'd0, 27'h0000013c, 5'd8, 27'h000000dc, 5'd19, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000039, 5'd6, 27'h0000010e, 5'd26, 27'h000003b4, 32'h00000400,
  1'd1,  5'd1, 27'h00000035, 5'd16, 27'h00000166, 5'd6, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d0, 5'd16, 27'h000003b1, 5'd19, 27'h0000033f, 32'h00000400,
  1'd1,  5'd1, 27'h00000303, 5'd19, 27'h00000212, 5'd27, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000021c, 5'd30, 27'h00000058, 5'd7, 27'h0000015e, 32'h00000400,
  1'd1,  5'd0, 27'h00000220, 5'd26, 27'h00000041, 5'd20, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a9, 5'd29, 27'h00000146, 5'd26, 27'h000001c5, 32'h00000400,
  1'd1,  5'd10, 27'h00000350, 5'd9, 27'h0000016b, 5'd5, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000038e, 5'd6, 27'h00000285, 5'd16, 27'h0000026b, 32'h00000400,
  1'd1,  5'd12, 27'h000001d4, 5'd8, 27'h000002c7, 5'd26, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000392, 5'd19, 27'h000000bb, 5'd8, 27'h000000bb, 32'h00000400,
  1'd1,  5'd14, 27'h000003fa, 5'd18, 27'h00000046, 5'd16, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000019c, 5'd19, 27'h000000ca, 5'd29, 27'h0000003d, 32'h00000400,
  1'd1,  5'd13, 27'h000001b8, 5'd26, 27'h000000d4, 5'd6, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002e4, 5'd26, 27'h0000010d, 5'd20, 27'h000000b2, 32'h00000400,
  1'd1,  5'd11, 27'h0000008e, 5'd29, 27'h000002a9, 5'd28, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000003b, 5'd9, 27'h000001a1, 5'd6, 27'h000000e6, 32'h00000400,
  1'd1,  5'd21, 27'h000000dd, 5'd6, 27'h0000024f, 5'd16, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000033d, 5'd5, 27'h0000023d, 5'd27, 27'h0000025e, 32'h00000400,
  1'd1,  5'd23, 27'h000003c8, 5'd17, 27'h00000164, 5'd6, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000203, 5'd16, 27'h000003d8, 5'd16, 27'h0000026c, 32'h00000400,
  1'd1,  5'd22, 27'h00000074, 5'd17, 27'h000003f1, 5'd27, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000291, 5'd26, 27'h00000106, 5'd6, 27'h00000123, 32'h00000400,
  1'd1,  5'd23, 27'h0000024d, 5'd26, 27'h000000b5, 5'd16, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a3, 5'd29, 27'h0000010c, 5'd30, 27'h00000363, 32'h00000400,
  1'd1,  5'd9, 27'h0000009a, 5'd4, 27'h000000d1, 5'd7, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d6, 5'd5, 27'h0000007c, 5'd19, 27'h000000f9, 32'h00000400,
  1'd1,  5'd7, 27'h000001e1, 5'd0, 27'h0000015f, 5'd26, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003f3, 5'd12, 27'h0000029d, 5'd1, 27'h0000018b, 32'h00000400,
  1'd1,  5'd7, 27'h000000c4, 5'd13, 27'h00000332, 5'd11, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000010e, 5'd13, 27'h000000a4, 5'd22, 27'h000000a7, 32'h00000400,
  1'd1,  5'd8, 27'h00000054, 5'd21, 27'h00000179, 5'd1, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000178, 5'd25, 27'h00000001, 5'd10, 27'h00000334, 32'h00000400,
  1'd1,  5'd7, 27'h000001d8, 5'd23, 27'h0000031f, 5'd22, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000095, 5'd2, 27'h00000134, 5'd9, 27'h000001d6, 32'h00000400,
  1'd1,  5'd19, 27'h000002a1, 5'd4, 27'h00000206, 5'd17, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000112, 5'd1, 27'h000000af, 5'd28, 27'h0000010c, 32'h00000400,
  1'd1,  5'd19, 27'h0000009a, 5'd11, 27'h0000023a, 5'd5, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000176, 5'd11, 27'h0000034f, 5'd13, 27'h000000e3, 32'h00000400,
  1'd1,  5'd18, 27'h0000021d, 5'd11, 27'h00000005, 5'd23, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000384, 5'd23, 27'h0000031d, 5'd4, 27'h000001b2, 32'h00000400,
  1'd1,  5'd19, 27'h000003f9, 5'd21, 27'h0000027c, 5'd11, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003bf, 5'd21, 27'h000001fd, 5'd22, 27'h00000378, 32'h00000400,
  1'd1,  5'd30, 27'h0000004a, 5'd1, 27'h00000299, 5'd3, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c4, 5'd0, 27'h000003e2, 5'd14, 27'h0000033a, 32'h00000400,
  1'd1,  5'd28, 27'h00000186, 5'd3, 27'h0000006f, 5'd24, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000010a, 5'd12, 27'h00000005, 5'd0, 27'h000003a3, 32'h00000400,
  1'd1,  5'd29, 27'h00000046, 5'd14, 27'h0000015e, 5'd13, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a8, 5'd11, 27'h00000306, 5'd24, 27'h00000283, 32'h00000400,
  1'd1,  5'd26, 27'h000002bf, 5'd23, 27'h000002ea, 5'd1, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000034d, 5'd24, 27'h000000fa, 5'd14, 27'h0000024c, 32'h00000400,
  1'd1,  5'd30, 27'h0000014d, 5'd24, 27'h00000223, 5'd22, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000197, 5'd2, 27'h000002ed, 5'd1, 27'h00000274, 32'h00000400,
  1'd1,  5'd5, 27'h000003cd, 5'd0, 27'h0000023b, 5'd12, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000303, 5'd4, 27'h000001ea, 5'd24, 27'h000001f1, 32'h00000400,
  1'd1,  5'd8, 27'h00000130, 5'd11, 27'h0000029b, 5'd5, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000122, 5'd14, 27'h000002c7, 5'd16, 27'h00000395, 32'h00000400,
  1'd1,  5'd8, 27'h00000064, 5'd13, 27'h0000020c, 5'd29, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000208, 5'd25, 27'h00000241, 5'd10, 27'h000000d2, 32'h00000400,
  1'd1,  5'd10, 27'h00000144, 5'd22, 27'h000003eb, 5'd19, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003fd, 5'd20, 27'h00000343, 5'd26, 27'h00000250, 32'h00000400,
  1'd1,  5'd19, 27'h0000034d, 5'd1, 27'h00000259, 5'd3, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000082, 5'd3, 27'h0000001f, 5'd14, 27'h0000010a, 32'h00000400,
  1'd1,  5'd15, 27'h00000394, 5'd2, 27'h00000256, 5'd23, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000314, 5'd15, 27'h0000018e, 5'd5, 27'h00000154, 32'h00000400,
  1'd1,  5'd19, 27'h0000023d, 5'd10, 27'h00000249, 5'd19, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000036e, 5'd10, 27'h00000226, 5'd29, 27'h00000300, 32'h00000400,
  1'd1,  5'd19, 27'h00000046, 5'd25, 27'h00000059, 5'd7, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000147, 5'd22, 27'h000003e9, 5'd18, 27'h00000043, 32'h00000400,
  1'd1,  5'd15, 27'h0000030f, 5'd24, 27'h000001a2, 5'd28, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e7, 5'd0, 27'h0000033b, 5'd5, 27'h000001cd, 32'h00000400,
  1'd1,  5'd28, 27'h0000003a, 5'd4, 27'h00000333, 5'd16, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000168, 5'd1, 27'h000002a9, 5'd28, 27'h0000039f, 32'h00000400,
  1'd1,  5'd27, 27'h000000c7, 5'd15, 27'h000001ad, 5'd5, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003fc, 5'd15, 27'h00000133, 5'd17, 27'h000000e3, 32'h00000400,
  1'd1,  5'd27, 27'h0000038e, 5'd12, 27'h00000107, 5'd30, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000011, 5'd24, 27'h00000261, 5'd7, 27'h0000027c, 32'h00000400,
  1'd1,  5'd28, 27'h00000066, 5'd23, 27'h0000032b, 5'd17, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000123, 5'd23, 27'h000003b6, 5'd30, 27'h000000f2, 32'h00000400,
  1'd1,  5'd8, 27'h000002ca, 5'd7, 27'h0000021a, 5'd2, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002d7, 5'd8, 27'h0000009e, 5'd14, 27'h000000d2, 32'h00000400,
  1'd1,  5'd5, 27'h00000139, 5'd6, 27'h000001f9, 5'd21, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003c3, 5'd16, 27'h00000299, 5'd1, 27'h000000ec, 32'h00000400,
  1'd1,  5'd6, 27'h0000034d, 5'd19, 27'h00000363, 5'd13, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000059, 5'd16, 27'h0000001c, 5'd21, 27'h00000192, 32'h00000400,
  1'd1,  5'd8, 27'h00000121, 5'd26, 27'h00000308, 5'd3, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021c, 5'd27, 27'h00000165, 5'd14, 27'h000001f1, 32'h00000400,
  1'd1,  5'd10, 27'h00000041, 5'd30, 27'h00000340, 5'd23, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000007f, 5'd6, 27'h00000252, 5'd2, 27'h000002f5, 32'h00000400,
  1'd1,  5'd17, 27'h0000037f, 5'd10, 27'h000000a2, 5'd10, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000030c, 5'd9, 27'h00000127, 5'd23, 27'h00000307, 32'h00000400,
  1'd1,  5'd16, 27'h00000304, 5'd16, 27'h00000016, 5'd0, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ba, 5'd20, 27'h0000000d, 5'd12, 27'h000001e1, 32'h00000400,
  1'd1,  5'd16, 27'h000002b1, 5'd17, 27'h00000202, 5'd25, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000301, 5'd28, 27'h00000246, 5'd3, 27'h0000027b, 32'h00000400,
  1'd1,  5'd20, 27'h0000017b, 5'd29, 27'h000002f0, 5'd12, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d7, 5'd27, 27'h00000308, 5'd21, 27'h000002f9, 32'h00000400,
  1'd1,  5'd28, 27'h0000034d, 5'd5, 27'h000002f6, 5'd4, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000035, 5'd8, 27'h000003b4, 5'd11, 27'h0000024d, 32'h00000400,
  1'd1,  5'd28, 27'h000000d6, 5'd10, 27'h00000050, 5'd25, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001d, 5'd17, 27'h000002ed, 5'd1, 27'h00000072, 32'h00000400,
  1'd1,  5'd29, 27'h000003d4, 5'd18, 27'h00000022, 5'd12, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000079, 5'd20, 27'h000000ac, 5'd23, 27'h000000e6, 32'h00000400,
  1'd1,  5'd28, 27'h00000252, 5'd28, 27'h00000140, 5'd3, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000133, 5'd26, 27'h000003b4, 5'd11, 27'h0000033a, 32'h00000400,
  1'd1,  5'd28, 27'h000003c0, 5'd26, 27'h0000024a, 5'd23, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000336, 5'd8, 27'h000001c1, 5'd5, 27'h000000de, 32'h00000400,
  1'd1,  5'd5, 27'h000002bb, 5'd6, 27'h000002a2, 5'd16, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000120, 5'd10, 27'h00000033, 5'd30, 27'h00000073, 32'h00000400,
  1'd1,  5'd7, 27'h000001ec, 5'd18, 27'h0000025a, 5'd7, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000397, 5'd16, 27'h000000b4, 5'd20, 27'h00000219, 32'h00000400,
  1'd1,  5'd6, 27'h00000173, 5'd15, 27'h0000033a, 5'd30, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000016e, 5'd28, 27'h000000f1, 5'd5, 27'h000001b4, 32'h00000400,
  1'd1,  5'd5, 27'h00000211, 5'd26, 27'h000000fd, 5'd18, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000f0, 5'd26, 27'h0000022a, 5'd30, 27'h00000247, 32'h00000400,
  1'd1,  5'd15, 27'h000003cf, 5'd9, 27'h00000223, 5'd8, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000305, 5'd8, 27'h00000022, 5'd16, 27'h00000096, 32'h00000400,
  1'd1,  5'd18, 27'h000003f2, 5'd6, 27'h000002df, 5'd27, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000230, 5'd20, 27'h00000165, 5'd9, 27'h0000030c, 32'h00000400,
  1'd1,  5'd20, 27'h0000028c, 5'd20, 27'h0000010a, 5'd17, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000017c, 5'd16, 27'h00000323, 5'd28, 27'h000002d3, 32'h00000400,
  1'd1,  5'd19, 27'h0000035e, 5'd29, 27'h0000011c, 5'd7, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000253, 5'd29, 27'h000001ab, 5'd17, 27'h000003f9, 32'h00000400,
  1'd1,  5'd16, 27'h000003c5, 5'd26, 27'h000001e1, 5'd26, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000331, 5'd9, 27'h00000097, 5'd8, 27'h000001bf, 32'h00000400,
  1'd1,  5'd29, 27'h000003aa, 5'd8, 27'h000002a7, 5'd18, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000021f, 5'd10, 27'h00000060, 5'd28, 27'h0000023f, 32'h00000400,
  1'd1,  5'd27, 27'h00000346, 5'd17, 27'h000003c8, 5'd10, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002ca, 5'd20, 27'h0000002e, 5'd16, 27'h000003c2, 32'h00000400,
  1'd1,  5'd30, 27'h0000008b, 5'd19, 27'h0000031a, 5'd28, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000004a, 5'd25, 27'h00000380, 5'd5, 27'h0000027d, 32'h00000400,
  1'd1,  5'd27, 27'h00000393, 5'd27, 27'h0000021e, 5'd20, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ea, 5'd28, 27'h0000035c, 5'd25, 27'h000003bf, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000000d8, 5'd0, 27'h0000016c, 5'd2, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000011a, 5'd3, 27'h000003f4, 5'd13, 27'h00000078, 32'h00000400,
  1'd1,  5'd2, 27'h00000205, 5'd0, 27'h00000243, 5'd23, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000283, 5'd11, 27'h00000225, 5'd2, 27'h00000302, 32'h00000400,
  1'd1,  5'd2, 27'h00000036, 5'd14, 27'h00000012, 5'd15, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000036a, 5'd12, 27'h00000104, 5'd24, 27'h0000023c, 32'h00000400,
  1'd1,  5'd3, 27'h000001ae, 5'd25, 27'h00000156, 5'd4, 27'h00000248, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001d8, 5'd21, 27'h000000cd, 5'd13, 27'h00000267, 32'h00000400,
  1'd1,  5'd1, 27'h000000d7, 5'd23, 27'h00000190, 5'd25, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c8, 5'd3, 27'h000001ea, 5'd2, 27'h00000244, 32'h00000400,
  1'd1,  5'd11, 27'h00000023, 5'd4, 27'h0000024e, 5'd11, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000022c, 5'd0, 27'h0000031a, 5'd22, 27'h00000166, 32'h00000400,
  1'd1,  5'd10, 27'h000003d0, 5'd10, 27'h000003a8, 5'd2, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029a, 5'd15, 27'h00000149, 5'd12, 27'h000001b1, 32'h00000400,
  1'd1,  5'd11, 27'h000000d1, 5'd11, 27'h000002f4, 5'd22, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001e6, 5'd21, 27'h000001e9, 5'd5, 27'h0000004b, 32'h00000400,
  1'd1,  5'd12, 27'h0000000c, 5'd21, 27'h000003a6, 5'd12, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a0, 5'd25, 27'h00000180, 5'd21, 27'h0000001f, 32'h00000400,
  1'd1,  5'd22, 27'h00000134, 5'd2, 27'h00000369, 5'd0, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000373, 5'd0, 27'h000000d1, 5'd10, 27'h0000034c, 32'h00000400,
  1'd1,  5'd23, 27'h0000022b, 5'd0, 27'h00000393, 5'd21, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000212, 5'd11, 27'h00000289, 5'd2, 27'h00000030, 32'h00000400,
  1'd1,  5'd23, 27'h0000009e, 5'd10, 27'h0000024d, 5'd12, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000292, 5'd13, 27'h000000ff, 5'd21, 27'h000003ee, 32'h00000400,
  1'd1,  5'd24, 27'h000003a2, 5'd22, 27'h0000027a, 5'd2, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000338, 5'd24, 27'h000000c5, 5'd14, 27'h000000f6, 32'h00000400,
  1'd1,  5'd22, 27'h0000032b, 5'd23, 27'h0000012a, 5'd22, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000202, 5'd2, 27'h0000010f, 5'd8, 27'h00000201, 32'h00000400,
  1'd1,  5'd0, 27'h00000098, 5'd5, 27'h00000023, 5'd16, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e9, 5'd2, 27'h0000020b, 5'd27, 27'h00000316, 32'h00000400,
  1'd1,  5'd2, 27'h0000001b, 5'd11, 27'h000002a9, 5'd6, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f9, 5'd10, 27'h000003f4, 5'd17, 27'h00000201, 32'h00000400,
  1'd1,  5'd0, 27'h0000004c, 5'd11, 27'h000001e0, 5'd27, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000099, 5'd25, 27'h00000074, 5'd8, 27'h000001b7, 32'h00000400,
  1'd1,  5'd2, 27'h00000113, 5'd25, 27'h000001b6, 5'd19, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000030b, 5'd23, 27'h000000a7, 5'd30, 27'h0000032e, 32'h00000400,
  1'd1,  5'd10, 27'h00000381, 5'd0, 27'h000000c2, 5'd9, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000385, 5'd1, 27'h00000239, 5'd17, 27'h00000262, 32'h00000400,
  1'd1,  5'd14, 27'h00000234, 5'd4, 27'h000000cf, 5'd29, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000018c, 5'd10, 27'h00000334, 5'd8, 27'h000001c1, 32'h00000400,
  1'd1,  5'd12, 27'h0000015e, 5'd11, 27'h000002f4, 5'd18, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000af, 5'd11, 27'h00000328, 5'd26, 27'h00000264, 32'h00000400,
  1'd1,  5'd12, 27'h00000166, 5'd23, 27'h00000076, 5'd8, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000034f, 5'd23, 27'h00000137, 5'd19, 27'h000001f9, 32'h00000400,
  1'd1,  5'd11, 27'h0000028f, 5'd23, 27'h0000012b, 5'd26, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003dc, 5'd3, 27'h0000029a, 5'd8, 27'h000002c5, 32'h00000400,
  1'd1,  5'd25, 27'h00000348, 5'd2, 27'h0000012d, 5'd16, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001fd, 5'd0, 27'h000000e7, 5'd30, 27'h00000200, 32'h00000400,
  1'd1,  5'd24, 27'h0000028a, 5'd14, 27'h00000233, 5'd6, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000004a, 5'd13, 27'h000003d2, 5'd19, 27'h0000033a, 32'h00000400,
  1'd1,  5'd23, 27'h00000221, 5'd11, 27'h0000008e, 5'd27, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000012d, 5'd24, 27'h00000340, 5'd10, 27'h00000039, 32'h00000400,
  1'd1,  5'd20, 27'h00000367, 5'd22, 27'h000001de, 5'd19, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021d, 5'd22, 27'h000003df, 5'd27, 27'h000001ac, 32'h00000400,
  1'd1,  5'd0, 27'h000002e4, 5'd7, 27'h0000018d, 5'd2, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001fd, 5'd7, 27'h000000f2, 5'd12, 27'h00000365, 32'h00000400,
  1'd1,  5'd0, 27'h00000016, 5'd5, 27'h000003ec, 5'd23, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000323, 5'd17, 27'h0000036e, 5'd0, 27'h000001dc, 32'h00000400,
  1'd1,  5'd2, 27'h0000018f, 5'd18, 27'h00000021, 5'd11, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b3, 5'd18, 27'h000001f9, 5'd23, 27'h000001ac, 32'h00000400,
  1'd1,  5'd2, 27'h0000005a, 5'd30, 27'h000002f1, 5'd5, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d3, 5'd30, 27'h00000247, 5'd14, 27'h0000027e, 32'h00000400,
  1'd1,  5'd4, 27'h0000016d, 5'd28, 27'h00000003, 5'd24, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018d, 5'd8, 27'h0000009a, 5'd3, 27'h00000035, 32'h00000400,
  1'd1,  5'd12, 27'h000002d4, 5'd9, 27'h0000030a, 5'd11, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e8, 5'd8, 27'h000001c8, 5'd23, 27'h0000001a, 32'h00000400,
  1'd1,  5'd13, 27'h0000036b, 5'd18, 27'h00000076, 5'd4, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029c, 5'd18, 27'h00000114, 5'd11, 27'h000002a9, 32'h00000400,
  1'd1,  5'd14, 27'h00000039, 5'd16, 27'h000002c1, 5'd24, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000079, 5'd30, 27'h00000223, 5'd2, 27'h000003d4, 32'h00000400,
  1'd1,  5'd12, 27'h000001e8, 5'd30, 27'h0000004d, 5'd10, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000027, 5'd26, 27'h0000014e, 5'd21, 27'h000002e7, 32'h00000400,
  1'd1,  5'd23, 27'h00000333, 5'd5, 27'h00000190, 5'd0, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000037, 5'd9, 27'h000001bf, 5'd14, 27'h00000370, 32'h00000400,
  1'd1,  5'd23, 27'h000000e2, 5'd9, 27'h00000237, 5'd23, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031c, 5'd17, 27'h00000111, 5'd3, 27'h00000001, 32'h00000400,
  1'd1,  5'd21, 27'h00000169, 5'd17, 27'h0000016f, 5'd14, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000fa, 5'd17, 27'h00000237, 5'd25, 27'h00000042, 32'h00000400,
  1'd1,  5'd21, 27'h00000032, 5'd30, 27'h000003a3, 5'd3, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c8, 5'd26, 27'h0000035c, 5'd13, 27'h00000320, 32'h00000400,
  1'd1,  5'd23, 27'h0000029d, 5'd29, 27'h000003b6, 5'd22, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000194, 5'd6, 27'h000002f0, 5'd7, 27'h00000206, 32'h00000400,
  1'd1,  5'd0, 27'h0000029d, 5'd8, 27'h00000020, 5'd16, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000047, 5'd7, 27'h000002db, 5'd27, 27'h000003f2, 32'h00000400,
  1'd1,  5'd0, 27'h0000011a, 5'd17, 27'h000002b4, 5'd7, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000033b, 5'd19, 27'h00000276, 5'd17, 27'h000000de, 32'h00000400,
  1'd1,  5'd4, 27'h0000016a, 5'd17, 27'h000003ae, 5'd28, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000240, 5'd27, 27'h00000261, 5'd8, 27'h000000d2, 32'h00000400,
  1'd1,  5'd1, 27'h00000296, 5'd26, 27'h000002ce, 5'd17, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000156, 5'd28, 27'h00000307, 5'd30, 27'h00000348, 32'h00000400,
  1'd1,  5'd12, 27'h00000141, 5'd10, 27'h00000082, 5'd9, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000006b, 5'd9, 27'h000002f0, 5'd18, 27'h000000d2, 32'h00000400,
  1'd1,  5'd12, 27'h00000313, 5'd5, 27'h0000028f, 5'd25, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001d7, 5'd15, 27'h0000024a, 5'd8, 27'h000001cb, 32'h00000400,
  1'd1,  5'd13, 27'h00000341, 5'd16, 27'h000002d1, 5'd20, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029a, 5'd18, 27'h000002ed, 5'd29, 27'h00000084, 32'h00000400,
  1'd1,  5'd12, 27'h00000047, 5'd26, 27'h00000392, 5'd7, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000003b, 5'd27, 27'h00000285, 5'd18, 27'h00000165, 32'h00000400,
  1'd1,  5'd13, 27'h000001f5, 5'd27, 27'h00000048, 5'd29, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000023, 5'd7, 27'h0000014c, 5'd10, 27'h00000126, 32'h00000400,
  1'd1,  5'd21, 27'h00000340, 5'd7, 27'h000000a6, 5'd15, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001e2, 5'd9, 27'h0000016d, 5'd29, 27'h000002d8, 32'h00000400,
  1'd1,  5'd25, 27'h000001b1, 5'd19, 27'h000001b6, 5'd6, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000180, 5'd16, 27'h0000019b, 5'd16, 27'h00000350, 32'h00000400,
  1'd1,  5'd22, 27'h000000d3, 5'd18, 27'h00000028, 5'd27, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000249, 5'd27, 27'h000000e8, 5'd6, 27'h0000006d, 32'h00000400,
  1'd1,  5'd21, 27'h000002f6, 5'd30, 27'h0000016c, 5'd20, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d4, 5'd27, 27'h000003e4, 5'd26, 27'h00000135, 32'h00000400,
  1'd1,  5'd10, 27'h000000e4, 5'd1, 27'h0000010a, 5'd10, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000030, 5'd4, 27'h00000095, 5'd16, 27'h000002c4, 32'h00000400,
  1'd1,  5'd7, 27'h0000016e, 5'd0, 27'h00000358, 5'd27, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000026d, 5'd11, 27'h000000fb, 5'd4, 27'h000003e4, 32'h00000400,
  1'd1,  5'd9, 27'h000001d8, 5'd12, 27'h00000384, 5'd12, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001c9, 5'd11, 27'h0000023a, 5'd22, 27'h00000117, 32'h00000400,
  1'd1,  5'd9, 27'h00000195, 5'd23, 27'h0000009f, 5'd1, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ed, 5'd21, 27'h0000008c, 5'd10, 27'h000001dc, 32'h00000400,
  1'd1,  5'd8, 27'h0000030a, 5'd21, 27'h000000af, 5'd25, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000012f, 5'd4, 27'h000002db, 5'd7, 27'h00000317, 32'h00000400,
  1'd1,  5'd17, 27'h00000077, 5'd1, 27'h000002d1, 5'd15, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000220, 5'd0, 27'h000003e5, 5'd28, 27'h000003c3, 32'h00000400,
  1'd1,  5'd19, 27'h00000270, 5'd10, 27'h000003f3, 5'd0, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d1, 5'd11, 27'h000003d1, 5'd13, 27'h00000218, 32'h00000400,
  1'd1,  5'd17, 27'h00000264, 5'd15, 27'h00000090, 5'd25, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000251, 5'd24, 27'h0000029d, 5'd3, 27'h000002e8, 32'h00000400,
  1'd1,  5'd18, 27'h000003b3, 5'd24, 27'h00000355, 5'd13, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000ca, 5'd23, 27'h0000003a, 5'd22, 27'h0000029d, 32'h00000400,
  1'd1,  5'd28, 27'h0000038f, 5'd4, 27'h00000004, 5'd1, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000038, 5'd1, 27'h000002d5, 5'd14, 27'h000002e4, 32'h00000400,
  1'd1,  5'd30, 27'h00000052, 5'd2, 27'h00000169, 5'd22, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001fc, 5'd12, 27'h0000002e, 5'd0, 27'h0000011b, 32'h00000400,
  1'd1,  5'd29, 27'h00000143, 5'd11, 27'h000001d3, 5'd14, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001fc, 5'd14, 27'h000001a8, 5'd23, 27'h000000a9, 32'h00000400,
  1'd1,  5'd30, 27'h00000142, 5'd25, 27'h00000056, 5'd4, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000f1, 5'd21, 27'h000000b5, 5'd11, 27'h00000265, 32'h00000400,
  1'd1,  5'd29, 27'h00000210, 5'd24, 27'h000000e9, 5'd22, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003dd, 5'd3, 27'h00000202, 5'd4, 27'h00000185, 32'h00000400,
  1'd1,  5'd6, 27'h0000005b, 5'd2, 27'h00000073, 5'd10, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ba, 5'd3, 27'h000000df, 5'd22, 27'h00000057, 32'h00000400,
  1'd1,  5'd6, 27'h0000012f, 5'd11, 27'h00000293, 5'd7, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000144, 5'd10, 27'h000002e6, 5'd17, 27'h00000242, 32'h00000400,
  1'd1,  5'd10, 27'h00000150, 5'd15, 27'h000000c1, 5'd28, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000233, 5'd24, 27'h000000fe, 5'd7, 27'h000003a3, 32'h00000400,
  1'd1,  5'd9, 27'h00000034, 5'd23, 27'h000002d5, 5'd20, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000026e, 5'd23, 27'h00000050, 5'd29, 27'h0000023d, 32'h00000400,
  1'd1,  5'd16, 27'h000001a0, 5'd0, 27'h0000029c, 5'd2, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003ce, 5'd1, 27'h000001eb, 5'd14, 27'h0000004e, 32'h00000400,
  1'd1,  5'd16, 27'h00000355, 5'd2, 27'h00000340, 5'd20, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000021e, 5'd14, 27'h0000002b, 5'd9, 27'h0000039d, 32'h00000400,
  1'd1,  5'd19, 27'h00000271, 5'd10, 27'h0000019d, 5'd19, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000304, 5'd14, 27'h000001cc, 5'd28, 27'h00000012, 32'h00000400,
  1'd1,  5'd19, 27'h00000107, 5'd20, 27'h00000320, 5'd7, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000004e, 5'd21, 27'h000003e9, 5'd19, 27'h000001bb, 32'h00000400,
  1'd1,  5'd18, 27'h00000325, 5'd22, 27'h00000093, 5'd30, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003b4, 5'd0, 27'h00000137, 5'd6, 27'h000001b6, 32'h00000400,
  1'd1,  5'd28, 27'h00000246, 5'd4, 27'h000001c7, 5'd18, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003d8, 5'd3, 27'h00000257, 5'd27, 27'h00000198, 32'h00000400,
  1'd1,  5'd28, 27'h000001d0, 5'd14, 27'h000000fe, 5'd5, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000240, 5'd12, 27'h00000367, 5'd19, 27'h00000007, 32'h00000400,
  1'd1,  5'd28, 27'h00000217, 5'd10, 27'h00000190, 5'd26, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000126, 5'd21, 27'h0000030e, 5'd6, 27'h000002a8, 32'h00000400,
  1'd1,  5'd29, 27'h000003c3, 5'd25, 27'h00000243, 5'd17, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003d6, 5'd21, 27'h000003e5, 5'd30, 27'h000000ee, 32'h00000400,
  1'd1,  5'd8, 27'h0000035d, 5'd10, 27'h00000144, 5'd3, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ac, 5'd6, 27'h000002be, 5'd13, 27'h00000124, 32'h00000400,
  1'd1,  5'd10, 27'h0000001d, 5'd9, 27'h00000027, 5'd20, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000001a, 5'd19, 27'h0000016a, 5'd0, 27'h0000021f, 32'h00000400,
  1'd1,  5'd6, 27'h00000299, 5'd19, 27'h00000230, 5'd13, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c7, 5'd16, 27'h000001a8, 5'd22, 27'h00000184, 32'h00000400,
  1'd1,  5'd8, 27'h000001a2, 5'd30, 27'h00000396, 5'd2, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000b, 5'd28, 27'h000002d0, 5'd14, 27'h000003d9, 32'h00000400,
  1'd1,  5'd10, 27'h00000072, 5'd27, 27'h00000186, 5'd23, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000137, 5'd8, 27'h000003cf, 5'd0, 27'h0000011e, 32'h00000400,
  1'd1,  5'd20, 27'h00000043, 5'd5, 27'h000000f5, 5'd10, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000019, 5'd7, 27'h0000035e, 5'd25, 27'h00000154, 32'h00000400,
  1'd1,  5'd17, 27'h0000022f, 5'd15, 27'h000003ae, 5'd2, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000023f, 5'd19, 27'h00000054, 5'd11, 27'h0000029d, 32'h00000400,
  1'd1,  5'd16, 27'h0000037b, 5'd17, 27'h00000204, 5'd21, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b7, 5'd27, 27'h000003ad, 5'd3, 27'h0000007b, 32'h00000400,
  1'd1,  5'd20, 27'h00000244, 5'd27, 27'h000002c1, 5'd12, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001d7, 5'd29, 27'h0000006d, 5'd22, 27'h00000064, 32'h00000400,
  1'd1,  5'd28, 27'h00000123, 5'd8, 27'h00000380, 5'd3, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002eb, 5'd10, 27'h000000c0, 5'd14, 27'h000000d6, 32'h00000400,
  1'd1,  5'd28, 27'h00000056, 5'd7, 27'h00000060, 5'd25, 27'h0000020c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ef, 5'd16, 27'h0000021f, 5'd4, 27'h00000022, 32'h00000400,
  1'd1,  5'd29, 27'h000002a6, 5'd17, 27'h000001b4, 5'd12, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000022b, 5'd17, 27'h0000011d, 5'd21, 27'h00000122, 32'h00000400,
  1'd1,  5'd27, 27'h0000037c, 5'd27, 27'h0000034b, 5'd2, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000028e, 5'd29, 27'h000001f1, 5'd14, 27'h0000033d, 32'h00000400,
  1'd1,  5'd29, 27'h0000012b, 5'd28, 27'h00000138, 5'd21, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002d4, 5'd9, 27'h000002f0, 5'd7, 27'h00000094, 32'h00000400,
  1'd1,  5'd6, 27'h00000106, 5'd9, 27'h00000280, 5'd17, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000018e, 5'd5, 27'h0000037b, 5'd28, 27'h00000223, 32'h00000400,
  1'd1,  5'd6, 27'h0000033e, 5'd19, 27'h00000372, 5'd7, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000308, 5'd17, 27'h000001e6, 5'd18, 27'h000001d4, 32'h00000400,
  1'd1,  5'd6, 27'h0000015d, 5'd18, 27'h00000073, 5'd30, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f3, 5'd27, 27'h000003eb, 5'd8, 27'h0000016c, 32'h00000400,
  1'd1,  5'd10, 27'h0000010e, 5'd30, 27'h000000ee, 5'd19, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b3, 5'd29, 27'h0000025e, 5'd28, 27'h00000341, 32'h00000400,
  1'd1,  5'd19, 27'h00000056, 5'd6, 27'h000001d9, 5'd9, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b0, 5'd8, 27'h00000311, 5'd18, 27'h000000a3, 32'h00000400,
  1'd1,  5'd16, 27'h00000284, 5'd9, 27'h000001d9, 5'd28, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002f0, 5'd15, 27'h000002c6, 5'd8, 27'h00000169, 32'h00000400,
  1'd1,  5'd17, 27'h00000300, 5'd15, 27'h00000349, 5'd16, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000030b, 5'd19, 27'h0000033a, 5'd28, 27'h00000369, 32'h00000400,
  1'd1,  5'd19, 27'h00000260, 5'd29, 27'h00000184, 5'd5, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002de, 5'd29, 27'h0000035b, 5'd17, 27'h00000096, 32'h00000400,
  1'd1,  5'd19, 27'h000001e5, 5'd27, 27'h0000027e, 5'd26, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000e3, 5'd6, 27'h00000213, 5'd6, 27'h000001a2, 32'h00000400,
  1'd1,  5'd30, 27'h00000335, 5'd6, 27'h00000050, 5'd20, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000370, 5'd5, 27'h000003a9, 5'd26, 27'h0000002e, 32'h00000400,
  1'd1,  5'd28, 27'h0000036c, 5'd20, 27'h000000ba, 5'd6, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000180, 5'd15, 27'h0000020c, 5'd17, 27'h00000203, 32'h00000400,
  1'd1,  5'd29, 27'h00000340, 5'd15, 27'h0000037d, 5'd27, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002fd, 5'd28, 27'h000001f7, 5'd6, 27'h00000359, 32'h00000400,
  1'd1,  5'd26, 27'h0000010e, 5'd29, 27'h0000025e, 5'd18, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000131, 5'd29, 27'h00000143, 5'd26, 27'h000000c1, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000001ae, 5'd2, 27'h000001fa, 5'd3, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d1, 5'd0, 27'h00000014, 5'd10, 27'h0000027c, 32'h00000400,
  1'd1,  5'd5, 27'h000000a8, 5'd5, 27'h00000070, 5'd25, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000178, 5'd13, 27'h00000032, 5'd4, 27'h00000310, 32'h00000400,
  1'd1,  5'd1, 27'h00000035, 5'd13, 27'h0000035c, 5'd10, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000031d, 5'd12, 27'h0000010d, 5'd24, 27'h0000006e, 32'h00000400,
  1'd1,  5'd1, 27'h00000384, 5'd21, 27'h00000226, 5'd3, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001d9, 5'd24, 27'h0000035a, 5'd14, 27'h0000011d, 32'h00000400,
  1'd1,  5'd2, 27'h000002c4, 5'd23, 27'h000002b5, 5'd24, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001db, 5'd1, 27'h00000361, 5'd1, 27'h000002b9, 32'h00000400,
  1'd1,  5'd14, 27'h000000dc, 5'd4, 27'h000001d5, 5'd13, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000074, 5'd2, 27'h0000010d, 5'd23, 27'h00000240, 32'h00000400,
  1'd1,  5'd14, 27'h0000036e, 5'd14, 27'h000002d3, 5'd4, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000326, 5'd14, 27'h000002f2, 5'd14, 27'h000000a2, 32'h00000400,
  1'd1,  5'd11, 27'h0000015c, 5'd15, 27'h000001c0, 5'd21, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000278, 5'd25, 27'h000001ab, 5'd2, 27'h000003b3, 32'h00000400,
  1'd1,  5'd10, 27'h00000223, 5'd23, 27'h00000198, 5'd12, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b3, 5'd25, 27'h00000068, 5'd22, 27'h00000241, 32'h00000400,
  1'd1,  5'd20, 27'h0000036d, 5'd1, 27'h00000160, 5'd4, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000004b, 5'd0, 27'h000002c8, 5'd13, 27'h0000033d, 32'h00000400,
  1'd1,  5'd22, 27'h000003e2, 5'd1, 27'h000000e0, 5'd24, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000187, 5'd13, 27'h0000019c, 5'd2, 27'h00000010, 32'h00000400,
  1'd1,  5'd25, 27'h000000f7, 5'd10, 27'h000003ef, 5'd15, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000b5, 5'd11, 27'h000000f7, 5'd23, 27'h000003f6, 32'h00000400,
  1'd1,  5'd22, 27'h00000172, 5'd23, 27'h000003f3, 5'd5, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000008b, 5'd23, 27'h000000ad, 5'd10, 27'h000002b7, 32'h00000400,
  1'd1,  5'd25, 27'h00000072, 5'd25, 27'h00000186, 5'd23, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000230, 5'd3, 27'h00000050, 5'd5, 27'h00000270, 32'h00000400,
  1'd1,  5'd3, 27'h000000eb, 5'd3, 27'h000003f3, 5'd17, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000126, 5'd3, 27'h00000050, 5'd26, 27'h00000133, 32'h00000400,
  1'd1,  5'd2, 27'h000000b1, 5'd12, 27'h0000023d, 5'd8, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000347, 5'd12, 27'h0000025e, 5'd19, 27'h00000331, 32'h00000400,
  1'd1,  5'd1, 27'h000003bd, 5'd14, 27'h00000006, 5'd26, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000347, 5'd23, 27'h00000359, 5'd7, 27'h0000020d, 32'h00000400,
  1'd1,  5'd0, 27'h00000298, 5'd24, 27'h0000024b, 5'd18, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000106, 5'd22, 27'h000002b0, 5'd29, 27'h0000016d, 32'h00000400,
  1'd1,  5'd12, 27'h000000f6, 5'd0, 27'h000000ef, 5'd6, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034c, 5'd3, 27'h0000005d, 5'd17, 27'h0000017b, 32'h00000400,
  1'd1,  5'd10, 27'h00000261, 5'd2, 27'h00000083, 5'd29, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000134, 5'd11, 27'h00000279, 5'd8, 27'h0000024d, 32'h00000400,
  1'd1,  5'd14, 27'h00000393, 5'd13, 27'h00000308, 5'd18, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000214, 5'd12, 27'h0000031e, 5'd28, 27'h000002e6, 32'h00000400,
  1'd1,  5'd13, 27'h0000030c, 5'd25, 27'h00000073, 5'd8, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003e, 5'd25, 27'h000002c7, 5'd17, 27'h000000ce, 32'h00000400,
  1'd1,  5'd13, 27'h00000222, 5'd25, 27'h00000141, 5'd30, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000323, 5'd2, 27'h000003aa, 5'd10, 27'h000000ea, 32'h00000400,
  1'd1,  5'd20, 27'h000002d5, 5'd1, 27'h00000342, 5'd15, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000101, 5'd3, 27'h00000313, 5'd26, 27'h000001d5, 32'h00000400,
  1'd1,  5'd24, 27'h00000316, 5'd10, 27'h00000218, 5'd8, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000032d, 5'd14, 27'h00000336, 5'd17, 27'h000003b8, 32'h00000400,
  1'd1,  5'd23, 27'h0000039c, 5'd11, 27'h0000010f, 5'd30, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000172, 5'd23, 27'h000003e7, 5'd5, 27'h0000011a, 32'h00000400,
  1'd1,  5'd21, 27'h0000008d, 5'd25, 27'h000000a8, 5'd18, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002af, 5'd24, 27'h00000104, 5'd29, 27'h00000090, 32'h00000400,
  1'd1,  5'd3, 27'h0000010c, 5'd9, 27'h00000134, 5'd2, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000006f, 5'd8, 27'h00000364, 5'd14, 27'h00000149, 32'h00000400,
  1'd1,  5'd4, 27'h000001a0, 5'd9, 27'h00000071, 5'd20, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000209, 5'd15, 27'h00000369, 5'd0, 27'h00000157, 32'h00000400,
  1'd1,  5'd4, 27'h0000021f, 5'd19, 27'h0000014a, 5'd12, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000312, 5'd16, 27'h00000361, 5'd20, 27'h000002b3, 32'h00000400,
  1'd1,  5'd0, 27'h000000db, 5'd29, 27'h0000005c, 5'd3, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f8, 5'd30, 27'h00000353, 5'd11, 27'h00000158, 32'h00000400,
  1'd1,  5'd2, 27'h00000183, 5'd26, 27'h000003a1, 5'd23, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001fb, 5'd7, 27'h00000016, 5'd1, 27'h00000038, 32'h00000400,
  1'd1,  5'd10, 27'h000002bb, 5'd10, 27'h0000001c, 5'd12, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a0, 5'd7, 27'h00000387, 5'd22, 27'h000003bf, 32'h00000400,
  1'd1,  5'd15, 27'h00000185, 5'd19, 27'h000003f9, 5'd2, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f2, 5'd16, 27'h000002f3, 5'd11, 27'h00000399, 32'h00000400,
  1'd1,  5'd11, 27'h000003c1, 5'd17, 27'h000002d6, 5'd22, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000261, 5'd28, 27'h000000ce, 5'd0, 27'h000003ab, 32'h00000400,
  1'd1,  5'd10, 27'h00000371, 5'd30, 27'h000000d5, 5'd13, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000201, 5'd26, 27'h0000033f, 5'd25, 27'h000001f6, 32'h00000400,
  1'd1,  5'd21, 27'h000001fe, 5'd10, 27'h0000013e, 5'd2, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002e0, 5'd9, 27'h00000378, 5'd10, 27'h0000019c, 32'h00000400,
  1'd1,  5'd25, 27'h0000026b, 5'd7, 27'h00000005, 5'd20, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000003f, 5'd15, 27'h000002f9, 5'd2, 27'h000002c6, 32'h00000400,
  1'd1,  5'd25, 27'h000002a9, 5'd16, 27'h00000075, 5'd11, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000249, 5'd19, 27'h00000179, 5'd23, 27'h000000c7, 32'h00000400,
  1'd1,  5'd24, 27'h0000003e, 5'd27, 27'h0000026b, 5'd4, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000050, 5'd27, 27'h000001ec, 5'd11, 27'h00000306, 32'h00000400,
  1'd1,  5'd22, 27'h0000002a, 5'd30, 27'h0000026b, 5'd23, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000266, 5'd6, 27'h000003e7, 5'd10, 27'h00000027, 32'h00000400,
  1'd1,  5'd2, 27'h0000028e, 5'd10, 27'h00000139, 5'd19, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002b1, 5'd7, 27'h000000a7, 5'd29, 27'h00000247, 32'h00000400,
  1'd1,  5'd0, 27'h000003f3, 5'd20, 27'h000000ad, 5'd7, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000365, 5'd17, 27'h00000204, 5'd18, 27'h0000023f, 32'h00000400,
  1'd1,  5'd2, 27'h0000022e, 5'd19, 27'h000001c0, 5'd30, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000004a, 5'd30, 27'h000003b2, 5'd6, 27'h0000006e, 32'h00000400,
  1'd1,  5'd0, 27'h000001ad, 5'd30, 27'h00000382, 5'd19, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000105, 5'd26, 27'h000002b0, 5'd26, 27'h0000020c, 32'h00000400,
  1'd1,  5'd13, 27'h000001e6, 5'd5, 27'h00000136, 5'd7, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000051, 5'd5, 27'h00000128, 5'd20, 27'h0000017e, 32'h00000400,
  1'd1,  5'd11, 27'h0000002a, 5'd6, 27'h00000245, 5'd28, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000322, 5'd17, 27'h000001cb, 5'd5, 27'h0000029d, 32'h00000400,
  1'd1,  5'd12, 27'h00000039, 5'd15, 27'h000003e6, 5'd17, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000000d, 5'd20, 27'h00000246, 5'd30, 27'h00000109, 32'h00000400,
  1'd1,  5'd14, 27'h00000207, 5'd28, 27'h000001e3, 5'd7, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000003a, 5'd26, 27'h0000005d, 5'd17, 27'h000003ea, 32'h00000400,
  1'd1,  5'd14, 27'h0000008e, 5'd30, 27'h0000023c, 5'd30, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a2, 5'd8, 27'h000002aa, 5'd6, 27'h000000d0, 32'h00000400,
  1'd1,  5'd21, 27'h0000033d, 5'd7, 27'h000003d0, 5'd19, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f3, 5'd8, 27'h000003b3, 5'd27, 27'h00000298, 32'h00000400,
  1'd1,  5'd21, 27'h0000005d, 5'd20, 27'h0000013d, 5'd6, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000059, 5'd16, 27'h00000287, 5'd16, 27'h00000140, 32'h00000400,
  1'd1,  5'd24, 27'h00000115, 5'd20, 27'h000000ab, 5'd30, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000dc, 5'd29, 27'h00000111, 5'd8, 27'h000002d5, 32'h00000400,
  1'd1,  5'd23, 27'h0000015e, 5'd28, 27'h000002ad, 5'd16, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000043, 5'd29, 27'h00000168, 5'd27, 27'h0000005d, 32'h00000400,
  1'd1,  5'd9, 27'h000001ca, 5'd4, 27'h000001f9, 5'd8, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000010e, 5'd4, 27'h00000279, 5'd19, 27'h000001ce, 32'h00000400,
  1'd1,  5'd7, 27'h00000332, 5'd0, 27'h0000030d, 5'd26, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ef, 5'd10, 27'h0000034a, 5'd3, 27'h00000260, 32'h00000400,
  1'd1,  5'd6, 27'h00000165, 5'd11, 27'h000003a7, 5'd12, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023a, 5'd13, 27'h000003c1, 5'd24, 27'h0000033f, 32'h00000400,
  1'd1,  5'd9, 27'h00000364, 5'd23, 27'h000000cc, 5'd3, 27'h00000364, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000008e, 5'd21, 27'h000000d6, 5'd14, 27'h00000387, 32'h00000400,
  1'd1,  5'd8, 27'h00000291, 5'd21, 27'h00000299, 5'd22, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000294, 5'd2, 27'h0000034c, 5'd8, 27'h000001fe, 32'h00000400,
  1'd1,  5'd16, 27'h000000e5, 5'd2, 27'h000002ad, 5'd19, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a6, 5'd0, 27'h00000234, 5'd28, 27'h0000003b, 32'h00000400,
  1'd1,  5'd19, 27'h000000bb, 5'd15, 27'h000001ce, 5'd3, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001d9, 5'd10, 27'h00000217, 5'd14, 27'h000002aa, 32'h00000400,
  1'd1,  5'd16, 27'h000002d7, 5'd11, 27'h00000322, 5'd20, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000024d, 5'd24, 27'h00000039, 5'd4, 27'h000002be, 32'h00000400,
  1'd1,  5'd16, 27'h000003d7, 5'd25, 27'h0000013d, 5'd14, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000042, 5'd23, 27'h00000311, 5'd25, 27'h000002e2, 32'h00000400,
  1'd1,  5'd28, 27'h000002c9, 5'd0, 27'h0000005d, 5'd0, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002ff, 5'd1, 27'h00000289, 5'd10, 27'h0000020a, 32'h00000400,
  1'd1,  5'd26, 27'h000001d7, 5'd0, 27'h000003d3, 5'd23, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000328, 5'd11, 27'h0000002c, 5'd3, 27'h00000130, 32'h00000400,
  1'd1,  5'd30, 27'h00000309, 5'd15, 27'h000000fa, 5'd15, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000012e, 5'd12, 27'h00000266, 5'd21, 27'h000003e4, 32'h00000400,
  1'd1,  5'd28, 27'h0000029f, 5'd22, 27'h000000a5, 5'd0, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021e, 5'd22, 27'h00000235, 5'd13, 27'h000003bf, 32'h00000400,
  1'd1,  5'd28, 27'h00000388, 5'd20, 27'h000002c5, 5'd23, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000037b, 5'd2, 27'h00000352, 5'd1, 27'h0000013a, 32'h00000400,
  1'd1,  5'd7, 27'h00000132, 5'd0, 27'h00000219, 5'd11, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000011b, 5'd3, 27'h00000295, 5'd25, 27'h00000205, 32'h00000400,
  1'd1,  5'd8, 27'h000002b0, 5'd12, 27'h00000094, 5'd8, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000017a, 5'd12, 27'h00000041, 5'd18, 27'h00000095, 32'h00000400,
  1'd1,  5'd6, 27'h00000015, 5'd15, 27'h00000003, 5'd27, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b5, 5'd21, 27'h00000247, 5'd6, 27'h00000256, 32'h00000400,
  1'd1,  5'd7, 27'h00000026, 5'd24, 27'h000003a0, 5'd18, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000037f, 5'd20, 27'h00000378, 5'd30, 27'h000001dd, 32'h00000400,
  1'd1,  5'd15, 27'h00000211, 5'd0, 27'h00000028, 5'd0, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000140, 5'd3, 27'h000002b9, 5'd12, 27'h00000056, 32'h00000400,
  1'd1,  5'd18, 27'h00000053, 5'd1, 27'h00000321, 5'd25, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ed, 5'd11, 27'h0000021a, 5'd6, 27'h0000002a, 32'h00000400,
  1'd1,  5'd20, 27'h00000138, 5'd13, 27'h0000005e, 5'd15, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000109, 5'd14, 27'h0000028b, 5'd28, 27'h00000371, 32'h00000400,
  1'd1,  5'd18, 27'h000000ae, 5'd22, 27'h000001cb, 5'd5, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000285, 5'd21, 27'h0000038f, 5'd15, 27'h00000262, 32'h00000400,
  1'd1,  5'd18, 27'h000003e6, 5'd23, 27'h0000014a, 5'd26, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002eb, 5'd4, 27'h00000157, 5'd6, 27'h0000036b, 32'h00000400,
  1'd1,  5'd29, 27'h000002a2, 5'd2, 27'h000000d0, 5'd19, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000336, 5'd3, 27'h000000af, 5'd26, 27'h0000005e, 32'h00000400,
  1'd1,  5'd27, 27'h00000239, 5'd14, 27'h00000358, 5'd6, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000288, 5'd13, 27'h00000183, 5'd16, 27'h00000234, 32'h00000400,
  1'd1,  5'd28, 27'h00000009, 5'd11, 27'h000001b5, 5'd26, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001be, 5'd24, 27'h00000214, 5'd6, 27'h000001cf, 32'h00000400,
  1'd1,  5'd30, 27'h00000275, 5'd20, 27'h00000348, 5'd17, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a0, 5'd25, 27'h0000021f, 5'd28, 27'h000003ff, 32'h00000400,
  1'd1,  5'd10, 27'h0000010b, 5'd7, 27'h00000098, 5'd0, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000011b, 5'd8, 27'h000001cb, 5'd11, 27'h000003c0, 32'h00000400,
  1'd1,  5'd5, 27'h00000211, 5'd5, 27'h00000263, 5'd20, 27'h000002e0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000c6, 5'd16, 27'h00000141, 5'd2, 27'h00000073, 32'h00000400,
  1'd1,  5'd10, 27'h00000022, 5'd15, 27'h00000224, 5'd11, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ba, 5'd17, 27'h000000cb, 5'd25, 27'h000002ad, 32'h00000400,
  1'd1,  5'd7, 27'h000000fe, 5'd30, 27'h0000027b, 5'd1, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c3, 5'd26, 27'h000001d7, 5'd12, 27'h00000307, 32'h00000400,
  1'd1,  5'd8, 27'h0000035b, 5'd30, 27'h00000142, 5'd25, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000188, 5'd5, 27'h000003dc, 5'd5, 27'h0000009a, 32'h00000400,
  1'd1,  5'd18, 27'h000000f9, 5'd6, 27'h000000e6, 5'd14, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000170, 5'd7, 27'h000001cf, 5'd21, 27'h000003f9, 32'h00000400,
  1'd1,  5'd17, 27'h000003d2, 5'd18, 27'h000002e2, 5'd4, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000268, 5'd20, 27'h00000078, 5'd11, 27'h000001f5, 32'h00000400,
  1'd1,  5'd17, 27'h00000371, 5'd17, 27'h0000024d, 5'd25, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000024e, 5'd30, 27'h000003e7, 5'd3, 27'h00000128, 32'h00000400,
  1'd1,  5'd19, 27'h000003f6, 5'd28, 27'h000001d5, 5'd12, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002ab, 5'd29, 27'h00000333, 5'd23, 27'h000001d7, 32'h00000400,
  1'd1,  5'd28, 27'h0000009c, 5'd7, 27'h00000344, 5'd4, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e1, 5'd9, 27'h00000091, 5'd14, 27'h000000a7, 32'h00000400,
  1'd1,  5'd28, 27'h0000012d, 5'd8, 27'h000001f2, 5'd25, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b2, 5'd15, 27'h00000273, 5'd0, 27'h000001f7, 32'h00000400,
  1'd1,  5'd30, 27'h000000b8, 5'd19, 27'h0000014b, 5'd12, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b4, 5'd19, 27'h000003d1, 5'd22, 27'h000000da, 32'h00000400,
  1'd1,  5'd29, 27'h0000032f, 5'd29, 27'h000003d0, 5'd4, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001df, 5'd26, 27'h0000024c, 5'd12, 27'h000002db, 32'h00000400,
  1'd1,  5'd26, 27'h00000385, 5'd27, 27'h00000001, 5'd22, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000001e, 5'd6, 27'h00000195, 5'd7, 27'h00000294, 32'h00000400,
  1'd1,  5'd8, 27'h00000149, 5'd10, 27'h0000001b, 5'd17, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000132, 5'd8, 27'h00000294, 5'd30, 27'h0000029b, 32'h00000400,
  1'd1,  5'd8, 27'h00000167, 5'd18, 27'h00000290, 5'd8, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000f9, 5'd19, 27'h000002af, 5'd20, 27'h000000ad, 32'h00000400,
  1'd1,  5'd6, 27'h00000169, 5'd17, 27'h000002bf, 5'd29, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000113, 5'd25, 27'h000003ce, 5'd6, 27'h00000086, 32'h00000400,
  1'd1,  5'd6, 27'h000002f7, 5'd29, 27'h0000021e, 5'd16, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000001a, 5'd30, 27'h000002b0, 5'd27, 27'h000000d8, 32'h00000400,
  1'd1,  5'd15, 27'h00000288, 5'd10, 27'h0000002f, 5'd6, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000228, 5'd5, 27'h000000e8, 5'd18, 27'h0000019c, 32'h00000400,
  1'd1,  5'd20, 27'h00000295, 5'd8, 27'h0000023f, 5'd26, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000323, 5'd16, 27'h00000275, 5'd6, 27'h000002a1, 32'h00000400,
  1'd1,  5'd19, 27'h000003e5, 5'd18, 27'h00000343, 5'd18, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003d3, 5'd15, 27'h00000297, 5'd28, 27'h000001b4, 32'h00000400,
  1'd1,  5'd20, 27'h000001ef, 5'd26, 27'h0000032f, 5'd5, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e2, 5'd26, 27'h00000274, 5'd16, 27'h000002ad, 32'h00000400,
  1'd1,  5'd18, 27'h00000265, 5'd27, 27'h00000260, 5'd30, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001dc, 5'd9, 27'h000002b6, 5'd8, 27'h00000085, 32'h00000400,
  1'd1,  5'd26, 27'h0000014e, 5'd9, 27'h0000019e, 5'd17, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f4, 5'd8, 27'h000001c5, 5'd28, 27'h0000017c, 32'h00000400,
  1'd1,  5'd27, 27'h000001f9, 5'd20, 27'h000000b6, 5'd8, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000245, 5'd17, 27'h000001be, 5'd19, 27'h00000382, 32'h00000400,
  1'd1,  5'd28, 27'h00000130, 5'd17, 27'h00000342, 5'd28, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000de, 5'd27, 27'h0000028c, 5'd6, 27'h0000022a, 32'h00000400,
  1'd1,  5'd27, 27'h00000219, 5'd29, 27'h0000034a, 5'd20, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000035e, 5'd28, 27'h000000ce, 5'd27, 27'h000000c9, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000095, 5'd0, 27'h00000384, 5'd0, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003a4, 5'd3, 27'h000001d0, 5'd14, 27'h00000077, 32'h00000400,
  1'd1,  5'd1, 27'h00000324, 5'd2, 27'h000003a0, 5'd21, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000026a, 5'd11, 27'h000000f2, 5'd2, 27'h00000169, 32'h00000400,
  1'd1,  5'd2, 27'h00000009, 5'd14, 27'h00000043, 5'd11, 27'h00000102, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001f0, 5'd11, 27'h00000299, 5'd24, 27'h00000386, 32'h00000400,
  1'd1,  5'd0, 27'h00000233, 5'd21, 27'h000001da, 5'd1, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000049, 5'd23, 27'h00000161, 5'd10, 27'h00000288, 32'h00000400,
  1'd1,  5'd3, 27'h000001ea, 5'd24, 27'h000002a4, 5'd25, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000025e, 5'd3, 27'h00000179, 5'd2, 27'h00000079, 32'h00000400,
  1'd1,  5'd11, 27'h0000009f, 5'd4, 27'h00000168, 5'd10, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000292, 5'd4, 27'h00000085, 5'd22, 27'h0000007c, 32'h00000400,
  1'd1,  5'd14, 27'h0000026f, 5'd15, 27'h0000015a, 5'd3, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000137, 5'd14, 27'h0000007d, 5'd11, 27'h00000016, 32'h00000400,
  1'd1,  5'd12, 27'h00000037, 5'd12, 27'h0000013d, 5'd22, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000018, 5'd22, 27'h00000254, 5'd2, 27'h000003aa, 32'h00000400,
  1'd1,  5'd11, 27'h0000003a, 5'd21, 27'h0000039c, 5'd14, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000022a, 5'd22, 27'h0000007e, 5'd24, 27'h0000001b, 32'h00000400,
  1'd1,  5'd22, 27'h00000003, 5'd0, 27'h00000345, 5'd1, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000019e, 5'd0, 27'h00000288, 5'd14, 27'h00000117, 32'h00000400,
  1'd1,  5'd23, 27'h00000219, 5'd3, 27'h00000232, 5'd21, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000005d, 5'd13, 27'h00000228, 5'd1, 27'h00000126, 32'h00000400,
  1'd1,  5'd22, 27'h00000153, 5'd15, 27'h0000002d, 5'd13, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000277, 5'd15, 27'h00000176, 5'd21, 27'h000003ff, 32'h00000400,
  1'd1,  5'd21, 27'h00000332, 5'd24, 27'h000003a1, 5'd2, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000087, 5'd22, 27'h00000296, 5'd11, 27'h00000376, 32'h00000400,
  1'd1,  5'd21, 27'h00000352, 5'd23, 27'h000000aa, 5'd23, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000347, 5'd0, 27'h0000005f, 5'd5, 27'h00000160, 32'h00000400,
  1'd1,  5'd3, 27'h00000152, 5'd4, 27'h0000023b, 5'd19, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000037, 5'd5, 27'h0000004d, 5'd27, 27'h000001f8, 32'h00000400,
  1'd1,  5'd1, 27'h00000167, 5'd14, 27'h0000030e, 5'd7, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000000c, 5'd11, 27'h000002bf, 5'd17, 27'h00000227, 32'h00000400,
  1'd1,  5'd4, 27'h00000324, 5'd13, 27'h0000009d, 5'd29, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000012b, 5'd24, 27'h00000096, 5'd8, 27'h000002eb, 32'h00000400,
  1'd1,  5'd1, 27'h000001fb, 5'd22, 27'h00000296, 5'd18, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000025, 5'd21, 27'h00000159, 5'd26, 27'h0000009e, 32'h00000400,
  1'd1,  5'd11, 27'h0000034d, 5'd3, 27'h0000003c, 5'd8, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000340, 5'd4, 27'h00000050, 5'd16, 27'h00000337, 32'h00000400,
  1'd1,  5'd12, 27'h000001b6, 5'd2, 27'h000001de, 5'd25, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000252, 5'd14, 27'h00000400, 5'd6, 27'h0000001c, 32'h00000400,
  1'd1,  5'd11, 27'h00000087, 5'd11, 27'h00000266, 5'd18, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000004, 5'd14, 27'h000000c2, 5'd28, 27'h00000040, 32'h00000400,
  1'd1,  5'd12, 27'h00000078, 5'd24, 27'h00000273, 5'd6, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000009, 5'd23, 27'h000003c6, 5'd16, 27'h00000091, 32'h00000400,
  1'd1,  5'd10, 27'h0000015c, 5'd25, 27'h000001dd, 5'd26, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f6, 5'd1, 27'h00000034, 5'd8, 27'h00000014, 32'h00000400,
  1'd1,  5'd23, 27'h000002a8, 5'd0, 27'h000003e6, 5'd15, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000037a, 5'd1, 27'h000000d5, 5'd29, 27'h000000c0, 32'h00000400,
  1'd1,  5'd24, 27'h0000000a, 5'd11, 27'h0000010f, 5'd8, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003ad, 5'd11, 27'h00000277, 5'd15, 27'h00000239, 32'h00000400,
  1'd1,  5'd22, 27'h000001ee, 5'd12, 27'h00000084, 5'd26, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000136, 5'd22, 27'h000003dd, 5'd9, 27'h00000224, 32'h00000400,
  1'd1,  5'd22, 27'h00000048, 5'd21, 27'h000000a1, 5'd19, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001f4, 5'd21, 27'h00000139, 5'd28, 27'h00000175, 32'h00000400,
  1'd1,  5'd2, 27'h00000294, 5'd6, 27'h000002c5, 5'd0, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003fb, 5'd10, 27'h000000ae, 5'd11, 27'h0000028e, 32'h00000400,
  1'd1,  5'd0, 27'h000001cf, 5'd9, 27'h000001c4, 5'd24, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000327, 5'd20, 27'h0000029b, 5'd4, 27'h000002e4, 32'h00000400,
  1'd1,  5'd0, 27'h0000015d, 5'd18, 27'h00000223, 5'd12, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000061, 5'd19, 27'h00000341, 5'd22, 27'h0000037f, 32'h00000400,
  1'd1,  5'd3, 27'h000003f9, 5'd29, 27'h000000a9, 5'd3, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000026d, 5'd27, 27'h000003d6, 5'd10, 27'h00000258, 32'h00000400,
  1'd1,  5'd3, 27'h000002c0, 5'd27, 27'h000000d1, 5'd25, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000029a, 5'd8, 27'h00000067, 5'd2, 27'h0000023e, 32'h00000400,
  1'd1,  5'd13, 27'h00000193, 5'd6, 27'h0000032c, 5'd14, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000345, 5'd6, 27'h00000086, 5'd20, 27'h00000390, 32'h00000400,
  1'd1,  5'd14, 27'h00000214, 5'd19, 27'h000000c6, 5'd2, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000019e, 5'd20, 27'h000000f0, 5'd11, 27'h0000006c, 32'h00000400,
  1'd1,  5'd15, 27'h00000136, 5'd20, 27'h00000296, 5'd22, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003fa, 5'd27, 27'h000001b1, 5'd4, 27'h00000271, 32'h00000400,
  1'd1,  5'd14, 27'h0000039a, 5'd26, 27'h00000367, 5'd13, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002fa, 5'd27, 27'h000001ba, 5'd23, 27'h000001b4, 32'h00000400,
  1'd1,  5'd21, 27'h0000005c, 5'd9, 27'h00000215, 5'd4, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000179, 5'd8, 27'h000003a7, 5'd14, 27'h000003a8, 32'h00000400,
  1'd1,  5'd21, 27'h00000167, 5'd6, 27'h0000031b, 5'd22, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000207, 5'd15, 27'h000002ed, 5'd5, 27'h00000067, 32'h00000400,
  1'd1,  5'd23, 27'h000003af, 5'd16, 27'h00000230, 5'd13, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003c5, 5'd16, 27'h0000006f, 5'd21, 27'h000001fa, 32'h00000400,
  1'd1,  5'd24, 27'h00000053, 5'd30, 27'h000003f1, 5'd0, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000015a, 5'd28, 27'h00000393, 5'd11, 27'h000000ab, 32'h00000400,
  1'd1,  5'd21, 27'h00000385, 5'd28, 27'h0000017c, 5'd21, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001a7, 5'd9, 27'h0000006d, 5'd10, 27'h00000100, 32'h00000400,
  1'd1,  5'd2, 27'h000001a8, 5'd9, 27'h0000032d, 5'd19, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000010, 5'd6, 27'h0000026c, 5'd26, 27'h00000105, 32'h00000400,
  1'd1,  5'd3, 27'h00000272, 5'd18, 27'h000001fb, 5'd8, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000133, 5'd19, 27'h00000014, 5'd19, 27'h0000005f, 32'h00000400,
  1'd1,  5'd1, 27'h00000287, 5'd16, 27'h000002aa, 5'd28, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002a9, 5'd29, 27'h00000244, 5'd5, 27'h000001d4, 32'h00000400,
  1'd1,  5'd4, 27'h000001b5, 5'd30, 27'h00000365, 5'd19, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ca, 5'd26, 27'h00000360, 5'd25, 27'h000003d6, 32'h00000400,
  1'd1,  5'd12, 27'h000003ac, 5'd8, 27'h0000003e, 5'd5, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e3, 5'd10, 27'h000000a3, 5'd16, 27'h000000f6, 32'h00000400,
  1'd1,  5'd10, 27'h000003cc, 5'd5, 27'h00000310, 5'd26, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ee, 5'd16, 27'h000003fc, 5'd6, 27'h00000035, 32'h00000400,
  1'd1,  5'd12, 27'h000000e0, 5'd20, 27'h000000e4, 5'd16, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000037b, 5'd15, 27'h000003a0, 5'd30, 27'h0000032a, 32'h00000400,
  1'd1,  5'd13, 27'h0000028f, 5'd27, 27'h000003e1, 5'd8, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000245, 5'd29, 27'h00000243, 5'd15, 27'h0000033c, 32'h00000400,
  1'd1,  5'd13, 27'h00000167, 5'd28, 27'h000000e6, 5'd27, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000e2, 5'd8, 27'h0000034b, 5'd6, 27'h000002a4, 32'h00000400,
  1'd1,  5'd24, 27'h00000366, 5'd9, 27'h00000308, 5'd19, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ef, 5'd5, 27'h00000395, 5'd28, 27'h000000cc, 32'h00000400,
  1'd1,  5'd23, 27'h00000272, 5'd16, 27'h000003f9, 5'd10, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000045, 5'd16, 27'h00000197, 5'd16, 27'h000000b5, 32'h00000400,
  1'd1,  5'd24, 27'h000000e1, 5'd18, 27'h000000d4, 5'd27, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000032, 5'd27, 27'h00000217, 5'd10, 27'h000000ab, 32'h00000400,
  1'd1,  5'd23, 27'h000000f7, 5'd27, 27'h00000211, 5'd16, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000103, 5'd27, 27'h00000297, 5'd26, 27'h0000009e, 32'h00000400,
  1'd1,  5'd5, 27'h000001df, 5'd4, 27'h00000120, 5'd8, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000bc, 5'd2, 27'h000002bf, 5'd16, 27'h000000f1, 32'h00000400,
  1'd1,  5'd7, 27'h00000278, 5'd4, 27'h000001d1, 5'd27, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000005, 5'd14, 27'h0000002f, 5'd3, 27'h00000143, 32'h00000400,
  1'd1,  5'd8, 27'h0000024f, 5'd15, 27'h00000070, 5'd10, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000272, 5'd14, 27'h000001ee, 5'd25, 27'h00000288, 32'h00000400,
  1'd1,  5'd9, 27'h00000087, 5'd23, 27'h00000377, 5'd3, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000247, 5'd21, 27'h00000263, 5'd12, 27'h00000186, 32'h00000400,
  1'd1,  5'd9, 27'h000000c6, 5'd24, 27'h00000045, 5'd25, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000000e, 5'd2, 27'h0000029e, 5'd9, 27'h00000038, 32'h00000400,
  1'd1,  5'd17, 27'h000002dc, 5'd0, 27'h00000400, 5'd16, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000237, 5'd1, 27'h00000099, 5'd29, 27'h00000193, 32'h00000400,
  1'd1,  5'd15, 27'h000003f5, 5'd11, 27'h00000296, 5'd2, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f5, 5'd15, 27'h00000040, 5'd14, 27'h00000220, 32'h00000400,
  1'd1,  5'd17, 27'h000001a1, 5'd15, 27'h000000fe, 5'd22, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000278, 5'd22, 27'h0000010d, 5'd4, 27'h00000310, 32'h00000400,
  1'd1,  5'd15, 27'h000002be, 5'd24, 27'h000000ee, 5'd12, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000275, 5'd22, 27'h0000001b, 5'd22, 27'h0000021f, 32'h00000400,
  1'd1,  5'd30, 27'h00000255, 5'd0, 27'h000001b6, 5'd2, 27'h00000217, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000344, 5'd5, 27'h00000076, 5'd12, 27'h000000e9, 32'h00000400,
  1'd1,  5'd25, 27'h000003d5, 5'd3, 27'h00000389, 5'd20, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b3, 5'd13, 27'h00000056, 5'd0, 27'h0000032f, 32'h00000400,
  1'd1,  5'd30, 27'h0000025a, 5'd11, 27'h0000008c, 5'd12, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000068, 5'd10, 27'h00000164, 5'd21, 27'h000000c6, 32'h00000400,
  1'd1,  5'd29, 27'h00000159, 5'd24, 27'h0000027e, 5'd4, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a1, 5'd23, 27'h00000250, 5'd13, 27'h000001dc, 32'h00000400,
  1'd1,  5'd26, 27'h0000008a, 5'd24, 27'h000003d4, 5'd25, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000039f, 5'd4, 27'h00000159, 5'd2, 27'h0000021f, 32'h00000400,
  1'd1,  5'd8, 27'h000002af, 5'd3, 27'h00000314, 5'd14, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007b, 5'd0, 27'h00000177, 5'd24, 27'h000002d9, 32'h00000400,
  1'd1,  5'd9, 27'h00000244, 5'd11, 27'h0000023a, 5'd7, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000278, 5'd10, 27'h0000024c, 5'd15, 27'h000003cf, 32'h00000400,
  1'd1,  5'd6, 27'h000001b9, 5'd13, 27'h000001f8, 5'd29, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000340, 5'd21, 27'h000003c2, 5'd6, 27'h0000027d, 32'h00000400,
  1'd1,  5'd7, 27'h000002ac, 5'd23, 27'h00000237, 5'd19, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000038a, 5'd22, 27'h0000021f, 5'd30, 27'h000003ce, 32'h00000400,
  1'd1,  5'd16, 27'h00000253, 5'd2, 27'h00000141, 5'd2, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000323, 5'd3, 27'h0000029c, 5'd10, 27'h000003f3, 32'h00000400,
  1'd1,  5'd18, 27'h00000347, 5'd4, 27'h00000140, 5'd23, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000010, 5'd14, 27'h00000326, 5'd5, 27'h00000388, 32'h00000400,
  1'd1,  5'd18, 27'h000001b5, 5'd14, 27'h0000018b, 5'd16, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000055, 5'd14, 27'h00000240, 5'd27, 27'h000002cc, 32'h00000400,
  1'd1,  5'd16, 27'h0000017f, 5'd25, 27'h00000324, 5'd8, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001d, 5'd23, 27'h000003b7, 5'd20, 27'h0000024d, 32'h00000400,
  1'd1,  5'd17, 27'h0000036e, 5'd23, 27'h000001c8, 5'd29, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000048, 5'd3, 27'h0000024d, 5'd8, 27'h000002ae, 32'h00000400,
  1'd1,  5'd26, 27'h00000380, 5'd2, 27'h000000a7, 5'd15, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000001a, 5'd1, 27'h000002cd, 5'd29, 27'h000002d1, 32'h00000400,
  1'd1,  5'd27, 27'h0000020c, 5'd13, 27'h000003c7, 5'd6, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000000, 5'd13, 27'h00000006, 5'd20, 27'h000001c0, 32'h00000400,
  1'd1,  5'd27, 27'h00000210, 5'd13, 27'h00000052, 5'd26, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000033d, 5'd20, 27'h000003f9, 5'd5, 27'h000002b5, 32'h00000400,
  1'd1,  5'd26, 27'h000001e0, 5'd21, 27'h00000366, 5'd19, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002da, 5'd21, 27'h000002d4, 5'd28, 27'h00000287, 32'h00000400,
  1'd1,  5'd8, 27'h000001db, 5'd9, 27'h00000376, 5'd0, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000359, 5'd7, 27'h000000f4, 5'd15, 27'h00000018, 32'h00000400,
  1'd1,  5'd10, 27'h000000e8, 5'd8, 27'h00000371, 5'd23, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007b, 5'd18, 27'h0000030d, 5'd0, 27'h0000015c, 32'h00000400,
  1'd1,  5'd6, 27'h000001d4, 5'd19, 27'h000001b6, 5'd14, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000154, 5'd17, 27'h000001c9, 5'd20, 27'h000002bf, 32'h00000400,
  1'd1,  5'd7, 27'h000001cf, 5'd28, 27'h00000387, 5'd0, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000020f, 5'd25, 27'h00000394, 5'd10, 27'h000002b2, 32'h00000400,
  1'd1,  5'd5, 27'h0000036b, 5'd29, 27'h0000005b, 5'd21, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001d6, 5'd7, 27'h000001d6, 5'd4, 27'h00000010, 32'h00000400,
  1'd1,  5'd17, 27'h00000339, 5'd5, 27'h000003a3, 5'd11, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ee, 5'd7, 27'h000002e6, 5'd24, 27'h0000005e, 32'h00000400,
  1'd1,  5'd17, 27'h000000e3, 5'd18, 27'h000002f0, 5'd3, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000024, 5'd16, 27'h00000162, 5'd14, 27'h00000115, 32'h00000400,
  1'd1,  5'd20, 27'h00000042, 5'd16, 27'h000000b8, 5'd22, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002de, 5'd30, 27'h00000358, 5'd0, 27'h000003c6, 32'h00000400,
  1'd1,  5'd18, 27'h00000198, 5'd29, 27'h00000193, 5'd14, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011c, 5'd27, 27'h000002ac, 5'd25, 27'h0000011f, 32'h00000400,
  1'd1,  5'd30, 27'h0000005b, 5'd7, 27'h000003cc, 5'd5, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000002e, 5'd7, 27'h0000024f, 5'd15, 27'h000000aa, 32'h00000400,
  1'd1,  5'd26, 27'h00000117, 5'd8, 27'h00000201, 5'd24, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001dd, 5'd16, 27'h000002d6, 5'd2, 27'h0000004a, 32'h00000400,
  1'd1,  5'd27, 27'h000000ca, 5'd16, 27'h00000097, 5'd14, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a1, 5'd19, 27'h00000358, 5'd22, 27'h00000217, 32'h00000400,
  1'd1,  5'd27, 27'h00000386, 5'd29, 27'h000002ba, 5'd1, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000fe, 5'd27, 27'h0000030a, 5'd13, 27'h000003b2, 32'h00000400,
  1'd1,  5'd28, 27'h000003c9, 5'd27, 27'h0000036e, 5'd22, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c0, 5'd9, 27'h00000129, 5'd7, 27'h00000178, 32'h00000400,
  1'd1,  5'd5, 27'h00000346, 5'd9, 27'h0000025f, 5'd19, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ae, 5'd5, 27'h00000189, 5'd27, 27'h00000117, 32'h00000400,
  1'd1,  5'd6, 27'h00000266, 5'd17, 27'h00000266, 5'd7, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000278, 5'd18, 27'h0000008a, 5'd20, 27'h0000020a, 32'h00000400,
  1'd1,  5'd5, 27'h000002c0, 5'd20, 27'h0000001d, 5'd28, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000235, 5'd26, 27'h00000172, 5'd8, 27'h000002c7, 32'h00000400,
  1'd1,  5'd7, 27'h000001bb, 5'd29, 27'h0000031f, 5'd19, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011e, 5'd26, 27'h000002d2, 5'd28, 27'h000000ca, 32'h00000400,
  1'd1,  5'd19, 27'h0000028f, 5'd10, 27'h00000056, 5'd5, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000008d, 5'd9, 27'h00000192, 5'd18, 27'h000000c4, 32'h00000400,
  1'd1,  5'd16, 27'h00000112, 5'd8, 27'h000001af, 5'd25, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000245, 5'd15, 27'h0000024f, 5'd10, 27'h00000000, 32'h00000400,
  1'd1,  5'd19, 27'h00000215, 5'd18, 27'h000000f5, 5'd18, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002c8, 5'd17, 27'h000000c8, 5'd30, 27'h000002fa, 32'h00000400,
  1'd1,  5'd19, 27'h000000b5, 5'd27, 27'h00000229, 5'd6, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019d, 5'd27, 27'h0000015d, 5'd16, 27'h0000032c, 32'h00000400,
  1'd1,  5'd19, 27'h00000155, 5'd28, 27'h0000013d, 5'd27, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025e, 5'd7, 27'h000003e8, 5'd6, 27'h000002e1, 32'h00000400,
  1'd1,  5'd26, 27'h0000029f, 5'd9, 27'h000001ee, 5'd16, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000238, 5'd7, 27'h000002c0, 5'd28, 27'h00000316, 32'h00000400,
  1'd1,  5'd27, 27'h00000069, 5'd20, 27'h000000e8, 5'd9, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f5, 5'd16, 27'h0000007c, 5'd15, 27'h00000310, 32'h00000400,
  1'd1,  5'd27, 27'h00000140, 5'd17, 27'h00000270, 5'd28, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000028b, 5'd30, 27'h00000382, 5'd5, 27'h00000275, 32'h00000400,
  1'd1,  5'd27, 27'h00000227, 5'd30, 27'h00000154, 5'd17, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000025d, 5'd30, 27'h000002f0, 5'd30, 27'h000000ef, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000003d4, 5'd3, 27'h0000028f, 5'd4, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002fe, 5'd1, 27'h0000017c, 5'd12, 27'h00000056, 32'h00000400,
  1'd1,  5'd2, 27'h00000229, 5'd2, 27'h00000144, 5'd21, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003f4, 5'd13, 27'h000003d5, 5'd3, 27'h000001bb, 32'h00000400,
  1'd1,  5'd1, 27'h000003d9, 5'd12, 27'h0000017c, 5'd13, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f1, 5'd14, 27'h000001b7, 5'd21, 27'h00000388, 32'h00000400,
  1'd1,  5'd2, 27'h0000012e, 5'd21, 27'h00000211, 5'd1, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000346, 5'd25, 27'h00000112, 5'd10, 27'h000003cc, 32'h00000400,
  1'd1,  5'd1, 27'h0000008b, 5'd21, 27'h00000173, 5'd25, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c0, 5'd0, 27'h000001fb, 5'd3, 27'h000001b2, 32'h00000400,
  1'd1,  5'd15, 27'h00000090, 5'd4, 27'h00000205, 5'd10, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000035, 5'd1, 27'h00000339, 5'd22, 27'h00000252, 32'h00000400,
  1'd1,  5'd14, 27'h00000286, 5'd10, 27'h0000032c, 5'd3, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ad, 5'd12, 27'h00000049, 5'd14, 27'h0000032f, 32'h00000400,
  1'd1,  5'd12, 27'h0000024b, 5'd14, 27'h0000006c, 5'd25, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003db, 5'd22, 27'h0000038b, 5'd1, 27'h0000016a, 32'h00000400,
  1'd1,  5'd14, 27'h00000037, 5'd23, 27'h0000013b, 5'd11, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000379, 5'd25, 27'h0000022b, 5'd24, 27'h00000191, 32'h00000400,
  1'd1,  5'd23, 27'h00000280, 5'd4, 27'h00000141, 5'd3, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000119, 5'd3, 27'h0000027a, 5'd14, 27'h0000019e, 32'h00000400,
  1'd1,  5'd22, 27'h00000095, 5'd3, 27'h0000000d, 5'd24, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000073, 5'd11, 27'h00000127, 5'd4, 27'h000002c8, 32'h00000400,
  1'd1,  5'd21, 27'h000002d2, 5'd11, 27'h00000259, 5'd10, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003c1, 5'd14, 27'h00000170, 5'd22, 27'h000001ab, 32'h00000400,
  1'd1,  5'd20, 27'h000002ec, 5'd21, 27'h000000ba, 5'd1, 27'h00000394, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000038a, 5'd21, 27'h0000023f, 5'd13, 27'h000003cd, 32'h00000400,
  1'd1,  5'd21, 27'h000001d0, 5'd25, 27'h0000000a, 5'd22, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d3, 5'd2, 27'h000003e1, 5'd9, 27'h00000239, 32'h00000400,
  1'd1,  5'd5, 27'h00000072, 5'd3, 27'h000003d4, 5'd17, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d8, 5'd4, 27'h000003a7, 5'd26, 27'h00000034, 32'h00000400,
  1'd1,  5'd1, 27'h00000279, 5'd10, 27'h000001b3, 5'd8, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000010e, 5'd13, 27'h0000030b, 5'd18, 27'h00000135, 32'h00000400,
  1'd1,  5'd2, 27'h00000308, 5'd14, 27'h000000b4, 5'd26, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000330, 5'd25, 27'h000001eb, 5'd10, 27'h00000119, 32'h00000400,
  1'd1,  5'd0, 27'h000002a0, 5'd24, 27'h0000025a, 5'd17, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000015f, 5'd24, 27'h0000004b, 5'd27, 27'h00000031, 32'h00000400,
  1'd1,  5'd14, 27'h000000e2, 5'd3, 27'h00000294, 5'd5, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000376, 5'd3, 27'h0000000e, 5'd20, 27'h000000ac, 32'h00000400,
  1'd1,  5'd13, 27'h000003ff, 5'd5, 27'h000000aa, 5'd26, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d1, 5'd15, 27'h000001f0, 5'd9, 27'h0000011d, 32'h00000400,
  1'd1,  5'd13, 27'h00000220, 5'd10, 27'h00000280, 5'd18, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000df, 5'd10, 27'h00000163, 5'd28, 27'h0000000b, 32'h00000400,
  1'd1,  5'd14, 27'h00000030, 5'd20, 27'h000003ff, 5'd6, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000358, 5'd25, 27'h0000023c, 5'd19, 27'h0000004c, 32'h00000400,
  1'd1,  5'd15, 27'h000001c7, 5'd20, 27'h000003f4, 5'd27, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000333, 5'd1, 27'h000001ae, 5'd9, 27'h000000c6, 32'h00000400,
  1'd1,  5'd21, 27'h000001aa, 5'd0, 27'h0000024e, 5'd18, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000004d, 5'd3, 27'h00000248, 5'd28, 27'h000000ac, 32'h00000400,
  1'd1,  5'd21, 27'h00000156, 5'd10, 27'h00000317, 5'd9, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001f4, 5'd10, 27'h00000213, 5'd18, 27'h000000bd, 32'h00000400,
  1'd1,  5'd22, 27'h000003df, 5'd15, 27'h000001ea, 5'd30, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c3, 5'd21, 27'h000002a6, 5'd6, 27'h000001d8, 32'h00000400,
  1'd1,  5'd22, 27'h000001eb, 5'd24, 27'h00000398, 5'd18, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ea, 5'd20, 27'h000002e4, 5'd28, 27'h000000de, 32'h00000400,
  1'd1,  5'd0, 27'h00000037, 5'd7, 27'h000003e9, 5'd5, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000123, 5'd5, 27'h000000f7, 5'd11, 27'h000001f6, 32'h00000400,
  1'd1,  5'd3, 27'h000003e6, 5'd8, 27'h0000005a, 5'd22, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000339, 5'd17, 27'h0000016c, 5'd3, 27'h0000009d, 32'h00000400,
  1'd1,  5'd1, 27'h0000030b, 5'd20, 27'h00000262, 5'd10, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001bb, 5'd16, 27'h000001d6, 5'd21, 27'h0000005b, 32'h00000400,
  1'd1,  5'd4, 27'h00000110, 5'd27, 27'h000001c0, 5'd2, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000004e, 5'd30, 27'h0000025a, 5'd14, 27'h0000026c, 32'h00000400,
  1'd1,  5'd1, 27'h000003f6, 5'd26, 27'h000003cb, 5'd21, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000079, 5'd7, 27'h00000206, 5'd2, 27'h000001d5, 32'h00000400,
  1'd1,  5'd14, 27'h0000032a, 5'd7, 27'h0000036c, 5'd14, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000188, 5'd7, 27'h00000066, 5'd22, 27'h00000060, 32'h00000400,
  1'd1,  5'd10, 27'h00000178, 5'd18, 27'h00000230, 5'd0, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000aa, 5'd20, 27'h0000013b, 5'd12, 27'h0000026a, 32'h00000400,
  1'd1,  5'd11, 27'h00000052, 5'd20, 27'h00000145, 5'd24, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000263, 5'd27, 27'h000000d3, 5'd3, 27'h00000148, 32'h00000400,
  1'd1,  5'd15, 27'h0000003f, 5'd30, 27'h000001e2, 5'd10, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000dc, 5'd28, 27'h0000027f, 5'd24, 27'h000000e4, 32'h00000400,
  1'd1,  5'd23, 27'h00000034, 5'd6, 27'h00000115, 5'd2, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000317, 5'd8, 27'h00000197, 5'd14, 27'h000000cb, 32'h00000400,
  1'd1,  5'd22, 27'h000002be, 5'd9, 27'h00000193, 5'd21, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b0, 5'd19, 27'h00000341, 5'd3, 27'h00000105, 32'h00000400,
  1'd1,  5'd25, 27'h0000002a, 5'd18, 27'h00000389, 5'd15, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000073, 5'd16, 27'h000003da, 5'd23, 27'h00000233, 32'h00000400,
  1'd1,  5'd25, 27'h00000184, 5'd29, 27'h000001b2, 5'd3, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002fa, 5'd27, 27'h0000002e, 5'd13, 27'h00000248, 32'h00000400,
  1'd1,  5'd23, 27'h000001dc, 5'd26, 27'h000003be, 5'd20, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000267, 5'd10, 27'h000000c6, 5'd10, 27'h00000110, 32'h00000400,
  1'd1,  5'd1, 27'h000003f9, 5'd10, 27'h0000010e, 5'd16, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000104, 5'd8, 27'h000000f6, 5'd28, 27'h00000170, 32'h00000400,
  1'd1,  5'd3, 27'h000000cf, 5'd19, 27'h0000012b, 5'd8, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000097, 5'd19, 27'h0000017c, 5'd16, 27'h000000db, 32'h00000400,
  1'd1,  5'd5, 27'h0000001e, 5'd18, 27'h00000311, 5'd28, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000001, 5'd28, 27'h00000041, 5'd6, 27'h0000014f, 32'h00000400,
  1'd1,  5'd1, 27'h000001e0, 5'd25, 27'h0000038a, 5'd19, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000294, 5'd26, 27'h00000124, 5'd27, 27'h00000180, 32'h00000400,
  1'd1,  5'd11, 27'h0000023e, 5'd5, 27'h0000033a, 5'd6, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000001d, 5'd9, 27'h00000026, 5'd18, 27'h0000024e, 32'h00000400,
  1'd1,  5'd13, 27'h000001f5, 5'd6, 27'h0000002e, 5'd28, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ae, 5'd17, 27'h00000379, 5'd7, 27'h00000185, 32'h00000400,
  1'd1,  5'd12, 27'h000000bf, 5'd19, 27'h00000234, 5'd16, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000007f, 5'd15, 27'h000002ad, 5'd26, 27'h00000315, 32'h00000400,
  1'd1,  5'd13, 27'h000003d4, 5'd30, 27'h000002ab, 5'd9, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000320, 5'd26, 27'h000003a7, 5'd20, 27'h000000b1, 32'h00000400,
  1'd1,  5'd14, 27'h0000007c, 5'd29, 27'h000001ef, 5'd26, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000032a, 5'd5, 27'h000000ed, 5'd9, 27'h000000b7, 32'h00000400,
  1'd1,  5'd24, 27'h00000063, 5'd8, 27'h000003a5, 5'd17, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f6, 5'd5, 27'h0000012b, 5'd25, 27'h0000038f, 32'h00000400,
  1'd1,  5'd22, 27'h00000108, 5'd19, 27'h00000193, 5'd7, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000a4, 5'd18, 27'h000000fd, 5'd16, 27'h0000034d, 32'h00000400,
  1'd1,  5'd24, 27'h00000286, 5'd17, 27'h000001ec, 5'd28, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000377, 5'd26, 27'h000003bb, 5'd8, 27'h000002cd, 32'h00000400,
  1'd1,  5'd25, 27'h00000088, 5'd28, 27'h0000002b, 5'd19, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ab, 5'd28, 27'h00000367, 5'd26, 27'h0000020c, 32'h00000400,
  1'd1,  5'd10, 27'h000000ce, 5'd2, 27'h00000151, 5'd5, 27'h0000035a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000378, 5'd3, 27'h000000d7, 5'd19, 27'h00000135, 32'h00000400,
  1'd1,  5'd9, 27'h0000003b, 5'd1, 27'h000001bb, 5'd27, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000003c, 5'd10, 27'h000001b1, 5'd3, 27'h00000074, 32'h00000400,
  1'd1,  5'd8, 27'h000000bd, 5'd14, 27'h0000025d, 5'd12, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000260, 5'd11, 27'h0000008f, 5'd21, 27'h00000126, 32'h00000400,
  1'd1,  5'd9, 27'h00000323, 5'd21, 27'h000002d2, 5'd2, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003f7, 5'd23, 27'h00000146, 5'd14, 27'h0000026f, 32'h00000400,
  1'd1,  5'd6, 27'h0000038f, 5'd22, 27'h000001f0, 5'd20, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031a, 5'd0, 27'h000000bf, 5'd7, 27'h000000b0, 32'h00000400,
  1'd1,  5'd18, 27'h00000256, 5'd0, 27'h000002c8, 5'd16, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000304, 5'd1, 27'h000003ea, 5'd28, 27'h0000008b, 32'h00000400,
  1'd1,  5'd19, 27'h000002cb, 5'd11, 27'h000003c7, 5'd5, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000242, 5'd11, 27'h00000287, 5'd15, 27'h00000030, 32'h00000400,
  1'd1,  5'd18, 27'h00000332, 5'd11, 27'h000001c6, 5'd22, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000320, 5'd21, 27'h000000e4, 5'd2, 27'h00000128, 32'h00000400,
  1'd1,  5'd19, 27'h0000027c, 5'd22, 27'h000002a1, 5'd13, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000111, 5'd20, 27'h00000301, 5'd25, 27'h00000335, 32'h00000400,
  1'd1,  5'd28, 27'h000000a2, 5'd2, 27'h00000001, 5'd1, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d1, 5'd2, 27'h00000116, 5'd11, 27'h0000013d, 32'h00000400,
  1'd1,  5'd26, 27'h00000037, 5'd0, 27'h0000004a, 5'd21, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000167, 5'd13, 27'h00000094, 5'd0, 27'h00000276, 32'h00000400,
  1'd1,  5'd30, 27'h0000034a, 5'd15, 27'h0000006e, 5'd13, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000036e, 5'd11, 27'h00000152, 5'd24, 27'h000000ad, 32'h00000400,
  1'd1,  5'd28, 27'h000002f8, 5'd25, 27'h000002dc, 5'd2, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000251, 5'd22, 27'h000001d7, 5'd15, 27'h0000018e, 32'h00000400,
  1'd1,  5'd26, 27'h00000206, 5'd25, 27'h00000318, 5'd21, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000b1, 5'd0, 27'h00000385, 5'd3, 27'h000000fe, 32'h00000400,
  1'd1,  5'd8, 27'h00000153, 5'd5, 27'h00000045, 5'd14, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000359, 5'd1, 27'h0000031a, 5'd24, 27'h000003dd, 32'h00000400,
  1'd1,  5'd9, 27'h000003cf, 5'd12, 27'h00000093, 5'd8, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000106, 5'd11, 27'h000002e5, 5'd15, 27'h000003a4, 32'h00000400,
  1'd1,  5'd8, 27'h00000150, 5'd12, 27'h000003a1, 5'd30, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000024a, 5'd21, 27'h0000010a, 5'd8, 27'h000003fb, 32'h00000400,
  1'd1,  5'd8, 27'h000003af, 5'd23, 27'h00000054, 5'd17, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000024f, 5'd24, 27'h00000304, 5'd28, 27'h000003b3, 32'h00000400,
  1'd1,  5'd16, 27'h00000019, 5'd0, 27'h000002a8, 5'd3, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000013, 5'd4, 27'h0000025a, 5'd11, 27'h00000400, 32'h00000400,
  1'd1,  5'd18, 27'h000001df, 5'd5, 27'h00000021, 5'd24, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000122, 5'd13, 27'h0000024a, 5'd6, 27'h00000030, 32'h00000400,
  1'd1,  5'd17, 27'h0000014f, 5'd15, 27'h00000120, 5'd17, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001cd, 5'd11, 27'h000001af, 5'd28, 27'h000001e7, 32'h00000400,
  1'd1,  5'd18, 27'h0000039b, 5'd24, 27'h0000016d, 5'd7, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000036f, 5'd25, 27'h00000048, 5'd17, 27'h000000f0, 32'h00000400,
  1'd1,  5'd20, 27'h000001aa, 5'd25, 27'h000000a4, 5'd27, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002a0, 5'd3, 27'h000003b8, 5'd8, 27'h00000299, 32'h00000400,
  1'd1,  5'd26, 27'h000002cb, 5'd0, 27'h000003e6, 5'd20, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001d5, 5'd2, 27'h000001af, 5'd29, 27'h00000067, 32'h00000400,
  1'd1,  5'd30, 27'h00000338, 5'd11, 27'h00000161, 5'd9, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003ce, 5'd11, 27'h0000033c, 5'd16, 27'h000002f5, 32'h00000400,
  1'd1,  5'd28, 27'h000000c3, 5'd12, 27'h000001f9, 5'd28, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000037, 5'd24, 27'h00000089, 5'd5, 27'h00000362, 32'h00000400,
  1'd1,  5'd27, 27'h00000306, 5'd25, 27'h00000030, 5'd15, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000133, 5'd22, 27'h000003b5, 5'd26, 27'h0000029f, 32'h00000400,
  1'd1,  5'd7, 27'h0000032c, 5'd8, 27'h00000265, 5'd1, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ce, 5'd6, 27'h00000134, 5'd12, 27'h00000339, 32'h00000400,
  1'd1,  5'd7, 27'h00000301, 5'd6, 27'h00000329, 5'd25, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000018a, 5'd19, 27'h0000024c, 5'd5, 27'h00000027, 32'h00000400,
  1'd1,  5'd9, 27'h0000025f, 5'd19, 27'h00000082, 5'd11, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000019e, 5'd18, 27'h00000122, 5'd22, 27'h00000304, 32'h00000400,
  1'd1,  5'd7, 27'h000003b0, 5'd29, 27'h000001dd, 5'd3, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000037f, 5'd25, 27'h00000396, 5'd13, 27'h0000008a, 32'h00000400,
  1'd1,  5'd6, 27'h000003dd, 5'd29, 27'h000003a4, 5'd24, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b3, 5'd6, 27'h00000330, 5'd3, 27'h000003d6, 32'h00000400,
  1'd1,  5'd18, 27'h0000037d, 5'd10, 27'h00000145, 5'd11, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000064, 5'd10, 27'h000000ff, 5'd21, 27'h000003d3, 32'h00000400,
  1'd1,  5'd19, 27'h00000152, 5'd17, 27'h000002d8, 5'd4, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000cd, 5'd17, 27'h00000351, 5'd11, 27'h000000a0, 32'h00000400,
  1'd1,  5'd17, 27'h00000256, 5'd17, 27'h00000157, 5'd20, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000005f, 5'd27, 27'h0000004b, 5'd3, 27'h000000c2, 32'h00000400,
  1'd1,  5'd18, 27'h000003db, 5'd26, 27'h000003f0, 5'd12, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000380, 5'd28, 27'h00000094, 5'd21, 27'h00000268, 32'h00000400,
  1'd1,  5'd28, 27'h00000248, 5'd6, 27'h000003f8, 5'd2, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c4, 5'd9, 27'h00000373, 5'd14, 27'h00000074, 32'h00000400,
  1'd1,  5'd30, 27'h00000220, 5'd8, 27'h0000033e, 5'd22, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003f5, 5'd18, 27'h0000026f, 5'd4, 27'h000002f0, 32'h00000400,
  1'd1,  5'd26, 27'h0000004a, 5'd17, 27'h000003a1, 5'd13, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000020c, 5'd18, 27'h000000e5, 5'd25, 27'h000001fc, 32'h00000400,
  1'd1,  5'd29, 27'h00000371, 5'd28, 27'h000002d2, 5'd1, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000312, 5'd28, 27'h000001e4, 5'd14, 27'h0000028e, 32'h00000400,
  1'd1,  5'd30, 27'h000001e7, 5'd30, 27'h0000034c, 5'd21, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000306, 5'd7, 27'h000000cf, 5'd7, 27'h0000036f, 32'h00000400,
  1'd1,  5'd8, 27'h000002c7, 5'd10, 27'h000000da, 5'd20, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000000f, 5'd10, 27'h000000e9, 5'd27, 27'h000000f8, 32'h00000400,
  1'd1,  5'd7, 27'h0000028e, 5'd18, 27'h0000028d, 5'd6, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001cd, 5'd16, 27'h00000131, 5'd17, 27'h000000a5, 32'h00000400,
  1'd1,  5'd9, 27'h0000028f, 5'd17, 27'h00000278, 5'd26, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000003a, 5'd30, 27'h00000394, 5'd6, 27'h000003fa, 32'h00000400,
  1'd1,  5'd5, 27'h00000330, 5'd29, 27'h000002bb, 5'd16, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003c1, 5'd26, 27'h00000348, 5'd27, 27'h00000284, 32'h00000400,
  1'd1,  5'd15, 27'h0000022b, 5'd6, 27'h0000006e, 5'd9, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002e8, 5'd8, 27'h00000371, 5'd18, 27'h000002c3, 32'h00000400,
  1'd1,  5'd20, 27'h00000050, 5'd9, 27'h00000274, 5'd29, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000081, 5'd16, 27'h000001a2, 5'd8, 27'h00000138, 32'h00000400,
  1'd1,  5'd20, 27'h000000fe, 5'd20, 27'h0000023f, 5'd19, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f0, 5'd19, 27'h0000015f, 5'd30, 27'h00000250, 32'h00000400,
  1'd1,  5'd19, 27'h000003bd, 5'd27, 27'h00000054, 5'd9, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002e8, 5'd28, 27'h00000139, 5'd18, 27'h00000335, 32'h00000400,
  1'd1,  5'd19, 27'h000001d9, 5'd27, 27'h000003ed, 5'd30, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000047, 5'd5, 27'h00000396, 5'd7, 27'h00000181, 32'h00000400,
  1'd1,  5'd28, 27'h0000006e, 5'd6, 27'h00000244, 5'd19, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012b, 5'd5, 27'h00000210, 5'd26, 27'h00000105, 32'h00000400,
  1'd1,  5'd28, 27'h000002a1, 5'd16, 27'h00000347, 5'd9, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000e3, 5'd15, 27'h000002dc, 5'd20, 27'h000001fa, 32'h00000400,
  1'd1,  5'd26, 27'h00000199, 5'd19, 27'h000001af, 5'd30, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024a, 5'd29, 27'h000002e6, 5'd6, 27'h00000013, 32'h00000400,
  1'd1,  5'd30, 27'h00000255, 5'd30, 27'h00000243, 5'd17, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000355, 5'd27, 27'h0000021a, 5'd29, 27'h00000199, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000379, 5'd4, 27'h00000286, 5'd5, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000fd, 5'd3, 27'h00000055, 5'd12, 27'h00000250, 32'h00000400,
  1'd1,  5'd0, 27'h00000291, 5'd4, 27'h000002b1, 5'd25, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000186, 5'd12, 27'h000002d9, 5'd0, 27'h0000012d, 32'h00000400,
  1'd1,  5'd1, 27'h000002be, 5'd10, 27'h000002fa, 5'd12, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000009e, 5'd13, 27'h00000132, 5'd21, 27'h0000003b, 32'h00000400,
  1'd1,  5'd2, 27'h00000079, 5'd20, 27'h00000336, 5'd4, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000289, 5'd25, 27'h000000b2, 5'd10, 27'h00000324, 32'h00000400,
  1'd1,  5'd3, 27'h000003ba, 5'd24, 27'h000002c8, 5'd25, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002b, 5'd0, 27'h000000b5, 5'd4, 27'h00000180, 32'h00000400,
  1'd1,  5'd11, 27'h000000c9, 5'd3, 27'h000002af, 5'd11, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000192, 5'd2, 27'h000000da, 5'd25, 27'h00000303, 32'h00000400,
  1'd1,  5'd14, 27'h00000282, 5'd13, 27'h00000288, 5'd4, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000013c, 5'd11, 27'h0000015d, 5'd13, 27'h000002a4, 32'h00000400,
  1'd1,  5'd10, 27'h00000172, 5'd10, 27'h00000399, 5'd24, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000010e, 5'd21, 27'h000002d5, 5'd1, 27'h000003b9, 32'h00000400,
  1'd1,  5'd12, 27'h000003dc, 5'd24, 27'h0000026a, 5'd13, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b0, 5'd22, 27'h00000208, 5'd21, 27'h0000019a, 32'h00000400,
  1'd1,  5'd22, 27'h0000024a, 5'd0, 27'h00000125, 5'd1, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c2, 5'd0, 27'h00000253, 5'd12, 27'h00000142, 32'h00000400,
  1'd1,  5'd22, 27'h00000309, 5'd1, 27'h000000fa, 5'd21, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000036b, 5'd11, 27'h000002ef, 5'd2, 27'h000002f1, 32'h00000400,
  1'd1,  5'd24, 27'h000002e9, 5'd13, 27'h000002c5, 5'd15, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000102, 5'd12, 27'h000003b4, 5'd25, 27'h000001b8, 32'h00000400,
  1'd1,  5'd24, 27'h00000014, 5'd21, 27'h00000026, 5'd0, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000350, 5'd22, 27'h000002a5, 5'd10, 27'h0000026c, 32'h00000400,
  1'd1,  5'd21, 27'h000003d5, 5'd23, 27'h0000019d, 5'd25, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029d, 5'd3, 27'h000000d4, 5'd9, 27'h0000007c, 32'h00000400,
  1'd1,  5'd0, 27'h00000310, 5'd2, 27'h000003f2, 5'd19, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002dd, 5'd3, 27'h00000313, 5'd26, 27'h000000b8, 32'h00000400,
  1'd1,  5'd1, 27'h00000242, 5'd13, 27'h00000177, 5'd6, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000037e, 5'd12, 27'h00000309, 5'd17, 27'h00000198, 32'h00000400,
  1'd1,  5'd2, 27'h000000c2, 5'd13, 27'h000001ea, 5'd27, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003de, 5'd21, 27'h000001d4, 5'd7, 27'h000003a8, 32'h00000400,
  1'd1,  5'd0, 27'h00000020, 5'd21, 27'h000003e6, 5'd16, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000031, 5'd24, 27'h00000189, 5'd30, 27'h000003f2, 32'h00000400,
  1'd1,  5'd15, 27'h000000e8, 5'd0, 27'h000003c1, 5'd6, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000034f, 5'd4, 27'h0000012e, 5'd17, 27'h00000035, 32'h00000400,
  1'd1,  5'd13, 27'h000000f0, 5'd4, 27'h000003f3, 5'd26, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000372, 5'd13, 27'h00000262, 5'd9, 27'h0000037b, 32'h00000400,
  1'd1,  5'd12, 27'h00000104, 5'd14, 27'h0000028c, 5'd17, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000245, 5'd14, 27'h000001c6, 5'd28, 27'h00000123, 32'h00000400,
  1'd1,  5'd12, 27'h0000025b, 5'd22, 27'h0000034a, 5'd6, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000233, 5'd22, 27'h000002ba, 5'd16, 27'h000001e2, 32'h00000400,
  1'd1,  5'd10, 27'h00000339, 5'd23, 27'h000002cb, 5'd30, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e1, 5'd4, 27'h0000010c, 5'd8, 27'h000001c5, 32'h00000400,
  1'd1,  5'd20, 27'h00000328, 5'd4, 27'h000002f4, 5'd17, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000bd, 5'd0, 27'h000001ee, 5'd29, 27'h00000277, 32'h00000400,
  1'd1,  5'd23, 27'h000002d6, 5'd11, 27'h000003f5, 5'd9, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000187, 5'd11, 27'h000002f1, 5'd18, 27'h000003fc, 32'h00000400,
  1'd1,  5'd24, 27'h0000030f, 5'd12, 27'h000000d3, 5'd29, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000100, 5'd22, 27'h0000020f, 5'd8, 27'h00000253, 32'h00000400,
  1'd1,  5'd24, 27'h000000b0, 5'd21, 27'h00000251, 5'd20, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000047, 5'd23, 27'h000001aa, 5'd28, 27'h0000023b, 32'h00000400,
  1'd1,  5'd2, 27'h00000326, 5'd7, 27'h0000025a, 5'd2, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000164, 5'd7, 27'h0000008b, 5'd11, 27'h000000ee, 32'h00000400,
  1'd1,  5'd4, 27'h000002bd, 5'd6, 27'h000003d7, 5'd20, 27'h000002f7, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000c8, 5'd16, 27'h00000245, 5'd2, 27'h00000036, 32'h00000400,
  1'd1,  5'd1, 27'h000000e1, 5'd19, 27'h00000227, 5'd13, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000038b, 5'd19, 27'h00000359, 5'd21, 27'h00000112, 32'h00000400,
  1'd1,  5'd3, 27'h00000322, 5'd28, 27'h000000d8, 5'd1, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e7, 5'd30, 27'h0000026b, 5'd14, 27'h000001c7, 32'h00000400,
  1'd1,  5'd1, 27'h0000003a, 5'd28, 27'h00000331, 5'd21, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ee, 5'd8, 27'h0000025e, 5'd2, 27'h0000031c, 32'h00000400,
  1'd1,  5'd13, 27'h00000381, 5'd6, 27'h00000055, 5'd11, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000243, 5'd8, 27'h00000222, 5'd21, 27'h000003bd, 32'h00000400,
  1'd1,  5'd10, 27'h00000282, 5'd17, 27'h00000043, 5'd1, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000320, 5'd16, 27'h00000303, 5'd10, 27'h00000298, 32'h00000400,
  1'd1,  5'd12, 27'h000000d7, 5'd18, 27'h00000154, 5'd25, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000016e, 5'd27, 27'h000003cf, 5'd4, 27'h000000db, 32'h00000400,
  1'd1,  5'd14, 27'h00000098, 5'd28, 27'h000002a6, 5'd12, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000191, 5'd25, 27'h000003d7, 5'd22, 27'h0000039c, 32'h00000400,
  1'd1,  5'd24, 27'h00000114, 5'd8, 27'h00000114, 5'd1, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000033f, 5'd5, 27'h0000019d, 5'd11, 27'h000001a6, 32'h00000400,
  1'd1,  5'd24, 27'h000003db, 5'd5, 27'h00000201, 5'd24, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c6, 5'd17, 27'h0000000b, 5'd2, 27'h00000227, 32'h00000400,
  1'd1,  5'd25, 27'h00000337, 5'd18, 27'h000001f5, 5'd11, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ae, 5'd16, 27'h000000bc, 5'd24, 27'h00000144, 32'h00000400,
  1'd1,  5'd23, 27'h0000017d, 5'd26, 27'h0000005c, 5'd0, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000304, 5'd30, 27'h000003c5, 5'd13, 27'h000000d0, 32'h00000400,
  1'd1,  5'd23, 27'h00000107, 5'd29, 27'h00000333, 5'd22, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002c5, 5'd7, 27'h0000024e, 5'd9, 27'h000003f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000315, 5'd6, 27'h0000019a, 5'd17, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000233, 5'd8, 27'h00000262, 5'd26, 27'h00000197, 32'h00000400,
  1'd1,  5'd1, 27'h00000039, 5'd16, 27'h00000089, 5'd8, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000135, 5'd16, 27'h000003fe, 5'd17, 27'h00000120, 32'h00000400,
  1'd1,  5'd4, 27'h000001e9, 5'd19, 27'h000002ff, 5'd27, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002bd, 5'd26, 27'h0000025f, 5'd8, 27'h000002ae, 32'h00000400,
  1'd1,  5'd2, 27'h000003c5, 5'd29, 27'h000001ab, 5'd17, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000096, 5'd26, 27'h00000144, 5'd29, 27'h0000012d, 32'h00000400,
  1'd1,  5'd15, 27'h000001ba, 5'd9, 27'h000001cb, 5'd7, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002e3, 5'd8, 27'h0000030f, 5'd15, 27'h000003e8, 32'h00000400,
  1'd1,  5'd11, 27'h0000039d, 5'd10, 27'h00000109, 5'd29, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001fa, 5'd17, 27'h0000038f, 5'd8, 27'h00000019, 32'h00000400,
  1'd1,  5'd14, 27'h0000025b, 5'd18, 27'h000001f7, 5'd15, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000227, 5'd15, 27'h000003e6, 5'd26, 27'h00000288, 32'h00000400,
  1'd1,  5'd12, 27'h00000120, 5'd30, 27'h00000220, 5'd9, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000338, 5'd28, 27'h00000258, 5'd17, 27'h0000015f, 32'h00000400,
  1'd1,  5'd10, 27'h00000293, 5'd29, 27'h0000014a, 5'd28, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002ab, 5'd7, 27'h00000385, 5'd9, 27'h00000185, 32'h00000400,
  1'd1,  5'd23, 27'h000003e8, 5'd9, 27'h0000018b, 5'd17, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002af, 5'd5, 27'h0000039b, 5'd27, 27'h000001b0, 32'h00000400,
  1'd1,  5'd24, 27'h00000000, 5'd17, 27'h0000014f, 5'd9, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000139, 5'd18, 27'h00000307, 5'd17, 27'h000000db, 32'h00000400,
  1'd1,  5'd21, 27'h0000009d, 5'd17, 27'h00000325, 5'd28, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031c, 5'd26, 27'h000002d5, 5'd5, 27'h0000015c, 32'h00000400,
  1'd1,  5'd24, 27'h0000021b, 5'd27, 27'h0000017e, 5'd18, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000366, 5'd27, 27'h000003b8, 5'd29, 27'h000002bc, 32'h00000400,
  1'd1,  5'd8, 27'h00000149, 5'd0, 27'h00000105, 5'd8, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000344, 5'd4, 27'h000003d9, 5'd18, 27'h0000025a, 32'h00000400,
  1'd1,  5'd8, 27'h00000198, 5'd3, 27'h00000016, 5'd26, 27'h00000009, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000326, 5'd11, 27'h00000275, 5'd0, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h00000176, 5'd12, 27'h00000308, 5'd12, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000305, 5'd15, 27'h000000f1, 5'd21, 27'h000000cd, 32'h00000400,
  1'd1,  5'd8, 27'h000003a6, 5'd22, 27'h0000010a, 5'd4, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ce, 5'd24, 27'h00000166, 5'd13, 27'h000001d7, 32'h00000400,
  1'd1,  5'd6, 27'h0000016c, 5'd24, 27'h00000313, 5'd24, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000074, 5'd1, 27'h0000010e, 5'd8, 27'h00000089, 32'h00000400,
  1'd1,  5'd19, 27'h0000012b, 5'd2, 27'h00000100, 5'd18, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003d0, 5'd2, 27'h0000004d, 5'd26, 27'h000003b4, 32'h00000400,
  1'd1,  5'd18, 27'h0000014c, 5'd12, 27'h000001df, 5'd0, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000208, 5'd11, 27'h0000018f, 5'd13, 27'h000001ce, 32'h00000400,
  1'd1,  5'd16, 27'h00000349, 5'd13, 27'h000002d8, 5'd23, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000328, 5'd24, 27'h00000372, 5'd2, 27'h00000274, 32'h00000400,
  1'd1,  5'd17, 27'h0000028a, 5'd22, 27'h000002c6, 5'd11, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000dc, 5'd22, 27'h0000016e, 5'd23, 27'h000000e2, 32'h00000400,
  1'd1,  5'd26, 27'h00000038, 5'd0, 27'h00000114, 5'd0, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000241, 5'd1, 27'h0000034f, 5'd10, 27'h00000394, 32'h00000400,
  1'd1,  5'd28, 27'h000000b3, 5'd2, 27'h000001a3, 5'd25, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000330, 5'd13, 27'h0000013b, 5'd4, 27'h00000052, 32'h00000400,
  1'd1,  5'd26, 27'h00000197, 5'd15, 27'h00000091, 5'd10, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002b5, 5'd13, 27'h000000c1, 5'd23, 27'h00000302, 32'h00000400,
  1'd1,  5'd28, 27'h00000179, 5'd20, 27'h00000361, 5'd3, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038b, 5'd20, 27'h000002e2, 5'd15, 27'h00000142, 32'h00000400,
  1'd1,  5'd30, 27'h00000008, 5'd25, 27'h000002ca, 5'd20, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000277, 5'd1, 27'h000001c4, 5'd4, 27'h0000021d, 32'h00000400,
  1'd1,  5'd6, 27'h0000024f, 5'd2, 27'h00000296, 5'd10, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000016b, 5'd4, 27'h000000c1, 5'd24, 27'h0000028c, 32'h00000400,
  1'd1,  5'd9, 27'h00000380, 5'd13, 27'h000002de, 5'd6, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000fa, 5'd15, 27'h00000116, 5'd17, 27'h00000388, 32'h00000400,
  1'd1,  5'd6, 27'h00000142, 5'd11, 27'h000000de, 5'd27, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003ad, 5'd23, 27'h000000f2, 5'd10, 27'h00000020, 32'h00000400,
  1'd1,  5'd7, 27'h000000f3, 5'd21, 27'h000002d5, 5'd18, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000089, 5'd24, 27'h0000010c, 5'd28, 27'h00000040, 32'h00000400,
  1'd1,  5'd16, 27'h000002c9, 5'd5, 27'h00000038, 5'd4, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f2, 5'd0, 27'h00000216, 5'd11, 27'h000001bd, 32'h00000400,
  1'd1,  5'd17, 27'h00000089, 5'd0, 27'h0000039e, 5'd22, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a6, 5'd11, 27'h000002d1, 5'd9, 27'h000000b0, 32'h00000400,
  1'd1,  5'd17, 27'h00000117, 5'd14, 27'h00000206, 5'd19, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002f8, 5'd15, 27'h000001d8, 5'd29, 27'h00000276, 32'h00000400,
  1'd1,  5'd17, 27'h00000156, 5'd24, 27'h000001f2, 5'd8, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000af, 5'd23, 27'h000003ea, 5'd18, 27'h000003d0, 32'h00000400,
  1'd1,  5'd18, 27'h000002d0, 5'd21, 27'h00000264, 5'd25, 27'h000003b3, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006f, 5'd1, 27'h00000273, 5'd6, 27'h0000011f, 32'h00000400,
  1'd1,  5'd25, 27'h000003ea, 5'd4, 27'h00000217, 5'd19, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000032d, 5'd3, 27'h00000018, 5'd28, 27'h0000015e, 32'h00000400,
  1'd1,  5'd29, 27'h000002c0, 5'd14, 27'h0000038b, 5'd9, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000029e, 5'd11, 27'h0000004c, 5'd15, 27'h00000245, 32'h00000400,
  1'd1,  5'd29, 27'h000002e2, 5'd14, 27'h00000185, 5'd29, 27'h000000e2, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000006a, 5'd21, 27'h0000030d, 5'd8, 27'h000002fe, 32'h00000400,
  1'd1,  5'd29, 27'h000000dd, 5'd21, 27'h00000065, 5'd20, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000034a, 5'd22, 27'h000000d6, 5'd27, 27'h00000297, 32'h00000400,
  1'd1,  5'd6, 27'h0000005c, 5'd8, 27'h0000016e, 5'd2, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000160, 5'd6, 27'h00000066, 5'd13, 27'h00000226, 32'h00000400,
  1'd1,  5'd7, 27'h00000111, 5'd8, 27'h0000034a, 5'd21, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000250, 5'd16, 27'h0000021d, 5'd0, 27'h00000014, 32'h00000400,
  1'd1,  5'd7, 27'h000000c0, 5'd19, 27'h000000af, 5'd13, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001d1, 5'd18, 27'h00000053, 5'd21, 27'h00000002, 32'h00000400,
  1'd1,  5'd9, 27'h0000002f, 5'd26, 27'h00000160, 5'd4, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000389, 5'd26, 27'h00000245, 5'd10, 27'h000002c0, 32'h00000400,
  1'd1,  5'd7, 27'h00000249, 5'd27, 27'h0000038a, 5'd22, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ea, 5'd6, 27'h00000394, 5'd5, 27'h000000a6, 32'h00000400,
  1'd1,  5'd15, 27'h00000383, 5'd6, 27'h00000071, 5'd11, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000163, 5'd8, 27'h000003a9, 5'd25, 27'h0000024e, 32'h00000400,
  1'd1,  5'd17, 27'h0000025c, 5'd17, 27'h000002e3, 5'd5, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002bd, 5'd17, 27'h00000295, 5'd14, 27'h00000262, 32'h00000400,
  1'd1,  5'd19, 27'h00000069, 5'd20, 27'h0000014f, 5'd22, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000c9, 5'd26, 27'h0000019b, 5'd1, 27'h0000011d, 32'h00000400,
  1'd1,  5'd18, 27'h00000195, 5'd26, 27'h000000f8, 5'd13, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ef, 5'd28, 27'h000000cb, 5'd23, 27'h0000023e, 32'h00000400,
  1'd1,  5'd30, 27'h000001f3, 5'd9, 27'h00000191, 5'd3, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000004c, 5'd5, 27'h0000026e, 5'd12, 27'h000002a2, 32'h00000400,
  1'd1,  5'd26, 27'h00000316, 5'd9, 27'h000000da, 5'd24, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c8, 5'd20, 27'h0000018c, 5'd0, 27'h0000014c, 32'h00000400,
  1'd1,  5'd30, 27'h00000367, 5'd18, 27'h0000011f, 5'd11, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c7, 5'd20, 27'h00000188, 5'd22, 27'h0000000c, 32'h00000400,
  1'd1,  5'd26, 27'h000002ec, 5'd26, 27'h000003cd, 5'd4, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000138, 5'd29, 27'h00000288, 5'd14, 27'h00000186, 32'h00000400,
  1'd1,  5'd29, 27'h00000276, 5'd28, 27'h00000147, 5'd24, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000130, 5'd9, 27'h000000ac, 5'd5, 27'h000003a6, 32'h00000400,
  1'd1,  5'd9, 27'h00000089, 5'd5, 27'h0000010d, 5'd20, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000136, 5'd8, 27'h000003a9, 5'd27, 27'h000002fa, 32'h00000400,
  1'd1,  5'd7, 27'h000000fc, 5'd15, 27'h00000270, 5'd6, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000137, 5'd17, 27'h00000060, 5'd16, 27'h00000154, 32'h00000400,
  1'd1,  5'd7, 27'h0000016f, 5'd17, 27'h00000356, 5'd30, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000001f, 5'd25, 27'h000003c4, 5'd7, 27'h000003b9, 32'h00000400,
  1'd1,  5'd6, 27'h00000013, 5'd27, 27'h000002f9, 5'd18, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000217, 5'd27, 27'h00000218, 5'd28, 27'h000002da, 32'h00000400,
  1'd1,  5'd16, 27'h00000283, 5'd9, 27'h000001b0, 5'd9, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000cc, 5'd6, 27'h00000374, 5'd17, 27'h000001f3, 32'h00000400,
  1'd1,  5'd16, 27'h0000016c, 5'd8, 27'h0000030f, 5'd28, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000113, 5'd17, 27'h0000000e, 5'd7, 27'h000000d8, 32'h00000400,
  1'd1,  5'd18, 27'h000003cc, 5'd19, 27'h000003f0, 5'd19, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d1, 5'd17, 27'h000000dc, 5'd30, 27'h0000038c, 32'h00000400,
  1'd1,  5'd20, 27'h00000165, 5'd29, 27'h000000ca, 5'd6, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000039e, 5'd29, 27'h000001d2, 5'd15, 27'h000002b5, 32'h00000400,
  1'd1,  5'd19, 27'h00000258, 5'd30, 27'h00000072, 5'd27, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000389, 5'd8, 27'h00000184, 5'd9, 27'h00000223, 32'h00000400,
  1'd1,  5'd26, 27'h0000033c, 5'd6, 27'h00000121, 5'd16, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a1, 5'd6, 27'h000001a4, 5'd30, 27'h000000de, 32'h00000400,
  1'd1,  5'd26, 27'h000001dd, 5'd16, 27'h00000318, 5'd8, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000fd, 5'd19, 27'h00000248, 5'd16, 27'h00000203, 32'h00000400,
  1'd1,  5'd29, 27'h000000b3, 5'd15, 27'h000003d7, 5'd29, 27'h000003da, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000325, 5'd29, 27'h00000303, 5'd9, 27'h0000034c, 32'h00000400,
  1'd1,  5'd29, 27'h00000198, 5'd27, 27'h00000353, 5'd17, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e2, 5'd30, 27'h000000bb, 5'd27, 27'h00000207, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000002c9, 5'd2, 27'h000000cd, 5'd1, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e7, 5'd4, 27'h000000c0, 5'd11, 27'h0000004c, 32'h00000400,
  1'd1,  5'd1, 27'h000003a0, 5'd4, 27'h00000308, 5'd25, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000fc, 5'd11, 27'h000000ca, 5'd3, 27'h000000bc, 32'h00000400,
  1'd1,  5'd3, 27'h000000c3, 5'd14, 27'h000000e2, 5'd10, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038c, 5'd14, 27'h00000101, 5'd24, 27'h00000146, 32'h00000400,
  1'd1,  5'd0, 27'h0000010d, 5'd24, 27'h00000135, 5'd0, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000391, 5'd21, 27'h000003e3, 5'd11, 27'h000002ad, 32'h00000400,
  1'd1,  5'd4, 27'h00000236, 5'd23, 27'h000001d1, 5'd22, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001d5, 5'd1, 27'h00000077, 5'd3, 27'h000003eb, 32'h00000400,
  1'd1,  5'd12, 27'h00000290, 5'd1, 27'h000002e9, 5'd14, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d0, 5'd1, 27'h0000008c, 5'd20, 27'h000002ef, 32'h00000400,
  1'd1,  5'd11, 27'h000003a3, 5'd14, 27'h00000120, 5'd2, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000315, 5'd10, 27'h000001ad, 5'd14, 27'h00000015, 32'h00000400,
  1'd1,  5'd12, 27'h00000223, 5'd13, 27'h000002f3, 5'd22, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001de, 5'd20, 27'h000002f3, 5'd4, 27'h00000155, 32'h00000400,
  1'd1,  5'd10, 27'h00000189, 5'd23, 27'h0000035e, 5'd14, 27'h00000189, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000349, 5'd24, 27'h000000a9, 5'd23, 27'h00000348, 32'h00000400,
  1'd1,  5'd25, 27'h000002ff, 5'd5, 27'h00000012, 5'd1, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d1, 5'd1, 27'h000002b9, 5'd11, 27'h0000006e, 32'h00000400,
  1'd1,  5'd22, 27'h000001b6, 5'd0, 27'h000001b2, 5'd24, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000266, 5'd10, 27'h00000210, 5'd4, 27'h0000007b, 32'h00000400,
  1'd1,  5'd23, 27'h00000199, 5'd10, 27'h000001d7, 5'd15, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000000c, 5'd12, 27'h000001be, 5'd22, 27'h00000361, 32'h00000400,
  1'd1,  5'd25, 27'h0000025e, 5'd21, 27'h00000164, 5'd3, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000018d, 5'd23, 27'h0000031b, 5'd12, 27'h000002ea, 32'h00000400,
  1'd1,  5'd24, 27'h00000293, 5'd21, 27'h0000028a, 5'd22, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001b3, 5'd3, 27'h00000374, 5'd5, 27'h000000ac, 32'h00000400,
  1'd1,  5'd2, 27'h0000023d, 5'd3, 27'h00000242, 5'd19, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000035f, 5'd2, 27'h0000020d, 5'd27, 27'h000000e0, 32'h00000400,
  1'd1,  5'd0, 27'h00000130, 5'd15, 27'h000001b0, 5'd8, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002b0, 5'd11, 27'h000002cb, 5'd16, 27'h0000033e, 32'h00000400,
  1'd1,  5'd2, 27'h000003c2, 5'd12, 27'h00000277, 5'd26, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000037, 5'd24, 27'h0000005e, 5'd5, 27'h00000110, 32'h00000400,
  1'd1,  5'd0, 27'h00000383, 5'd21, 27'h00000370, 5'd18, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000034b, 5'd22, 27'h000001c0, 5'd27, 27'h00000294, 32'h00000400,
  1'd1,  5'd10, 27'h00000356, 5'd3, 27'h00000180, 5'd9, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000265, 5'd4, 27'h00000214, 5'd15, 27'h0000035e, 32'h00000400,
  1'd1,  5'd14, 27'h00000125, 5'd0, 27'h0000023e, 5'd30, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000115, 5'd14, 27'h000003d5, 5'd7, 27'h00000343, 32'h00000400,
  1'd1,  5'd11, 27'h00000323, 5'd13, 27'h000002cd, 5'd16, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d1, 5'd11, 27'h0000006d, 5'd27, 27'h0000023b, 32'h00000400,
  1'd1,  5'd12, 27'h0000026e, 5'd23, 27'h00000161, 5'd8, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e2, 5'd21, 27'h0000005e, 5'd18, 27'h00000250, 32'h00000400,
  1'd1,  5'd14, 27'h000001df, 5'd22, 27'h000002f9, 5'd30, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001db, 5'd1, 27'h00000222, 5'd6, 27'h00000162, 32'h00000400,
  1'd1,  5'd24, 27'h00000073, 5'd1, 27'h0000037e, 5'd15, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000027c, 5'd3, 27'h00000291, 5'd29, 27'h00000046, 32'h00000400,
  1'd1,  5'd22, 27'h000003c9, 5'd13, 27'h000003a3, 5'd7, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003dc, 5'd11, 27'h00000088, 5'd17, 27'h00000158, 32'h00000400,
  1'd1,  5'd21, 27'h000003ec, 5'd14, 27'h00000306, 5'd26, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002ab, 5'd22, 27'h00000360, 5'd7, 27'h0000010c, 32'h00000400,
  1'd1,  5'd21, 27'h000003e2, 5'd25, 27'h00000310, 5'd19, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000023, 5'd21, 27'h00000242, 5'd30, 27'h000001ba, 32'h00000400,
  1'd1,  5'd1, 27'h000002a0, 5'd7, 27'h000002f9, 5'd0, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000034f, 5'd6, 27'h0000023e, 5'd10, 27'h00000274, 32'h00000400,
  1'd1,  5'd1, 27'h0000039d, 5'd8, 27'h0000034b, 5'd23, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000290, 5'd18, 27'h0000002a, 5'd2, 27'h000003a9, 32'h00000400,
  1'd1,  5'd4, 27'h000000ec, 5'd17, 27'h000003ad, 5'd13, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000029f, 5'd15, 27'h00000311, 5'd24, 27'h000002fe, 32'h00000400,
  1'd1,  5'd2, 27'h0000001f, 5'd30, 27'h0000001e, 5'd1, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002f, 5'd27, 27'h0000014a, 5'd13, 27'h00000042, 32'h00000400,
  1'd1,  5'd4, 27'h0000031e, 5'd28, 27'h000000bb, 5'd21, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fe, 5'd8, 27'h0000008d, 5'd2, 27'h000001a2, 32'h00000400,
  1'd1,  5'd10, 27'h000001c3, 5'd10, 27'h00000076, 5'd14, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000095, 5'd10, 27'h0000014d, 5'd25, 27'h000001cf, 32'h00000400,
  1'd1,  5'd14, 27'h000003a9, 5'd19, 27'h00000305, 5'd0, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000021c, 5'd20, 27'h000001ae, 5'd10, 27'h00000226, 32'h00000400,
  1'd1,  5'd13, 27'h000003bd, 5'd17, 27'h00000119, 5'd22, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000090, 5'd26, 27'h000003ac, 5'd4, 27'h00000273, 32'h00000400,
  1'd1,  5'd13, 27'h00000108, 5'd28, 27'h00000386, 5'd12, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000031b, 5'd30, 27'h00000352, 5'd22, 27'h000002e6, 32'h00000400,
  1'd1,  5'd23, 27'h00000251, 5'd8, 27'h000001e7, 5'd0, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000120, 5'd6, 27'h000002f1, 5'd13, 27'h000001a1, 32'h00000400,
  1'd1,  5'd21, 27'h0000001c, 5'd6, 27'h000000ba, 5'd23, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000008e, 5'd20, 27'h000001c0, 5'd1, 27'h00000062, 32'h00000400,
  1'd1,  5'd24, 27'h000001fb, 5'd18, 27'h0000030c, 5'd13, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000198, 5'd19, 27'h0000026b, 5'd24, 27'h00000156, 32'h00000400,
  1'd1,  5'd23, 27'h0000012a, 5'd26, 27'h00000199, 5'd2, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000287, 5'd30, 27'h0000000b, 5'd12, 27'h00000298, 32'h00000400,
  1'd1,  5'd20, 27'h000003db, 5'd26, 27'h00000056, 5'd21, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014e, 5'd7, 27'h00000062, 5'd5, 27'h000001e5, 32'h00000400,
  1'd1,  5'd0, 27'h00000201, 5'd7, 27'h000003c0, 5'd16, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000043, 5'd5, 27'h000003e2, 5'd28, 27'h000000a1, 32'h00000400,
  1'd1,  5'd1, 27'h00000207, 5'd19, 27'h0000003f, 5'd7, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000dc, 5'd18, 27'h000001fe, 5'd19, 27'h000003cd, 32'h00000400,
  1'd1,  5'd2, 27'h0000008a, 5'd20, 27'h000001c2, 5'd26, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000376, 5'd27, 27'h00000215, 5'd6, 27'h0000008d, 32'h00000400,
  1'd1,  5'd3, 27'h000003d9, 5'd30, 27'h0000038b, 5'd18, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000032f, 5'd30, 27'h000000b4, 5'd28, 27'h00000184, 32'h00000400,
  1'd1,  5'd14, 27'h00000275, 5'd5, 27'h0000011b, 5'd7, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003e4, 5'd7, 27'h00000189, 5'd16, 27'h0000000a, 32'h00000400,
  1'd1,  5'd11, 27'h000000d4, 5'd7, 27'h00000198, 5'd26, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000013c, 5'd17, 27'h00000223, 5'd6, 27'h00000352, 32'h00000400,
  1'd1,  5'd12, 27'h000001d3, 5'd19, 27'h00000292, 5'd20, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000119, 5'd16, 27'h0000034d, 5'd26, 27'h000001f3, 32'h00000400,
  1'd1,  5'd11, 27'h00000188, 5'd29, 27'h000000aa, 5'd9, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c2, 5'd29, 27'h000001d6, 5'd16, 27'h00000275, 32'h00000400,
  1'd1,  5'd11, 27'h00000398, 5'd30, 27'h00000306, 5'd27, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000187, 5'd6, 27'h0000026f, 5'd9, 27'h00000033, 32'h00000400,
  1'd1,  5'd20, 27'h000003c1, 5'd6, 27'h00000107, 5'd17, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000033f, 5'd7, 27'h00000085, 5'd27, 27'h000000ed, 32'h00000400,
  1'd1,  5'd22, 27'h000002e3, 5'd17, 27'h00000282, 5'd7, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000038b, 5'd18, 27'h00000371, 5'd19, 27'h000001b1, 32'h00000400,
  1'd1,  5'd20, 27'h00000314, 5'd16, 27'h00000381, 5'd28, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000170, 5'd30, 27'h00000035, 5'd8, 27'h00000025, 32'h00000400,
  1'd1,  5'd23, 27'h000000c7, 5'd28, 27'h000001cd, 5'd15, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ef, 5'd27, 27'h00000223, 5'd30, 27'h0000005a, 32'h00000400,
  1'd1,  5'd8, 27'h00000101, 5'd4, 27'h00000180, 5'd7, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000349, 5'd0, 27'h00000015, 5'd19, 27'h000000f2, 32'h00000400,
  1'd1,  5'd9, 27'h000003c4, 5'd3, 27'h000000d6, 5'd26, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000266, 5'd13, 27'h00000046, 5'd4, 27'h0000029a, 32'h00000400,
  1'd1,  5'd6, 27'h000002f5, 5'd13, 27'h00000311, 5'd12, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e7, 5'd12, 27'h000001bd, 5'd21, 27'h0000030c, 32'h00000400,
  1'd1,  5'd9, 27'h0000034e, 5'd24, 27'h000000e3, 5'd1, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000010, 5'd21, 27'h000002ea, 5'd15, 27'h000001ad, 32'h00000400,
  1'd1,  5'd9, 27'h000000ac, 5'd24, 27'h00000015, 5'd22, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000017f, 5'd4, 27'h0000027e, 5'd6, 27'h000002a8, 32'h00000400,
  1'd1,  5'd17, 27'h0000034b, 5'd2, 27'h0000005f, 5'd17, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000053, 5'd2, 27'h00000011, 5'd29, 27'h00000104, 32'h00000400,
  1'd1,  5'd18, 27'h00000284, 5'd11, 27'h00000060, 5'd3, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003e0, 5'd10, 27'h000003bb, 5'd15, 27'h00000129, 32'h00000400,
  1'd1,  5'd18, 27'h000002f8, 5'd12, 27'h000002e8, 5'd22, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000116, 5'd23, 27'h00000391, 5'd2, 27'h000001b3, 32'h00000400,
  1'd1,  5'd19, 27'h0000011b, 5'd25, 27'h00000074, 5'd13, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000262, 5'd25, 27'h00000166, 5'd23, 27'h0000009e, 32'h00000400,
  1'd1,  5'd28, 27'h000003f2, 5'd4, 27'h000000bd, 5'd4, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a4, 5'd3, 27'h00000200, 5'd12, 27'h0000028d, 32'h00000400,
  1'd1,  5'd27, 27'h00000017, 5'd3, 27'h000000a6, 5'd21, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000de, 5'd10, 27'h000001b6, 5'd1, 27'h00000354, 32'h00000400,
  1'd1,  5'd29, 27'h00000171, 5'd12, 27'h0000031d, 5'd14, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000289, 5'd12, 27'h00000100, 5'd21, 27'h0000010b, 32'h00000400,
  1'd1,  5'd27, 27'h000002b3, 5'd21, 27'h0000005e, 5'd0, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002eb, 5'd21, 27'h0000039c, 5'd13, 27'h00000224, 32'h00000400,
  1'd1,  5'd27, 27'h00000255, 5'd25, 27'h00000007, 5'd20, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000334, 5'd0, 27'h00000090, 5'd2, 27'h0000032e, 32'h00000400,
  1'd1,  5'd9, 27'h0000023d, 5'd3, 27'h0000025e, 5'd12, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ec, 5'd0, 27'h000000fa, 5'd23, 27'h000001ec, 32'h00000400,
  1'd1,  5'd5, 27'h000003b1, 5'd14, 27'h0000032d, 5'd7, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000247, 5'd12, 27'h000001ae, 5'd19, 27'h00000352, 32'h00000400,
  1'd1,  5'd7, 27'h00000182, 5'd13, 27'h000001fd, 5'd30, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b4, 5'd22, 27'h00000254, 5'd6, 27'h00000318, 32'h00000400,
  1'd1,  5'd5, 27'h000000d0, 5'd25, 27'h000002f6, 5'd17, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002c0, 5'd25, 27'h00000082, 5'd30, 27'h000002ec, 32'h00000400,
  1'd1,  5'd16, 27'h00000356, 5'd2, 27'h0000022b, 5'd1, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000c2, 5'd5, 27'h00000044, 5'd15, 27'h000001c2, 32'h00000400,
  1'd1,  5'd20, 27'h00000052, 5'd4, 27'h00000126, 5'd21, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000011c, 5'd15, 27'h00000183, 5'd5, 27'h000001da, 32'h00000400,
  1'd1,  5'd19, 27'h0000027a, 5'd11, 27'h000002c8, 5'd16, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030b, 5'd14, 27'h0000013d, 5'd27, 27'h000002b1, 32'h00000400,
  1'd1,  5'd18, 27'h000000d3, 5'd25, 27'h00000175, 5'd9, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000034e, 5'd25, 27'h0000018f, 5'd17, 27'h00000350, 32'h00000400,
  1'd1,  5'd17, 27'h0000002e, 5'd20, 27'h00000385, 5'd30, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000346, 5'd0, 27'h000000b0, 5'd5, 27'h00000319, 32'h00000400,
  1'd1,  5'd29, 27'h0000021f, 5'd4, 27'h000002dc, 5'd19, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003d0, 5'd3, 27'h0000036f, 5'd30, 27'h000000c6, 32'h00000400,
  1'd1,  5'd26, 27'h00000039, 5'd11, 27'h0000023a, 5'd7, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000042, 5'd12, 27'h000000b4, 5'd15, 27'h00000271, 32'h00000400,
  1'd1,  5'd30, 27'h00000110, 5'd14, 27'h000000c7, 5'd30, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000000, 5'd24, 27'h0000015d, 5'd7, 27'h00000100, 32'h00000400,
  1'd1,  5'd27, 27'h00000118, 5'd23, 27'h0000018c, 5'd19, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003d9, 5'd22, 27'h00000140, 5'd30, 27'h0000017e, 32'h00000400,
  1'd1,  5'd8, 27'h00000071, 5'd7, 27'h000002f8, 5'd2, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000146, 5'd6, 27'h0000038a, 5'd13, 27'h000002cc, 32'h00000400,
  1'd1,  5'd9, 27'h0000003c, 5'd9, 27'h0000023a, 5'd21, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d2, 5'd16, 27'h00000342, 5'd1, 27'h00000155, 32'h00000400,
  1'd1,  5'd6, 27'h0000023a, 5'd19, 27'h00000287, 5'd13, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002be, 5'd19, 27'h0000007f, 5'd23, 27'h000000d7, 32'h00000400,
  1'd1,  5'd9, 27'h000003db, 5'd27, 27'h0000015a, 5'd0, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000221, 5'd28, 27'h000003dd, 5'd10, 27'h0000022b, 32'h00000400,
  1'd1,  5'd7, 27'h00000076, 5'd26, 27'h00000136, 5'd21, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c4, 5'd8, 27'h00000279, 5'd4, 27'h00000234, 32'h00000400,
  1'd1,  5'd17, 27'h0000009b, 5'd6, 27'h000003a6, 5'd14, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000103, 5'd8, 27'h00000370, 5'd20, 27'h000002ee, 32'h00000400,
  1'd1,  5'd15, 27'h0000032a, 5'd18, 27'h000000bf, 5'd5, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000037b, 5'd19, 27'h000001c5, 5'd10, 27'h0000034f, 32'h00000400,
  1'd1,  5'd20, 27'h0000014f, 5'd20, 27'h00000206, 5'd24, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000f7, 5'd28, 27'h00000319, 5'd2, 27'h00000284, 32'h00000400,
  1'd1,  5'd19, 27'h0000021e, 5'd26, 27'h0000000a, 5'd10, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000375, 5'd28, 27'h000000cf, 5'd23, 27'h00000135, 32'h00000400,
  1'd1,  5'd29, 27'h00000155, 5'd9, 27'h000001bd, 5'd4, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000384, 5'd6, 27'h00000038, 5'd15, 27'h000001db, 32'h00000400,
  1'd1,  5'd28, 27'h00000312, 5'd8, 27'h00000351, 5'd23, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000d4, 5'd18, 27'h000002d8, 5'd0, 27'h00000068, 32'h00000400,
  1'd1,  5'd29, 27'h00000260, 5'd20, 27'h00000298, 5'd12, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000214, 5'd16, 27'h00000090, 5'd20, 27'h000003db, 32'h00000400,
  1'd1,  5'd29, 27'h00000322, 5'd25, 27'h000003da, 5'd0, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000fd, 5'd27, 27'h000002e1, 5'd13, 27'h000003a4, 32'h00000400,
  1'd1,  5'd27, 27'h000001e0, 5'd27, 27'h0000038d, 5'd25, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002a3, 5'd7, 27'h00000098, 5'd8, 27'h00000211, 32'h00000400,
  1'd1,  5'd7, 27'h000001d4, 5'd9, 27'h00000152, 5'd15, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000225, 5'd9, 27'h000003e9, 5'd26, 27'h0000013c, 32'h00000400,
  1'd1,  5'd8, 27'h0000037f, 5'd19, 27'h000001ac, 5'd8, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e1, 5'd19, 27'h000003a1, 5'd17, 27'h00000345, 32'h00000400,
  1'd1,  5'd8, 27'h00000300, 5'd17, 27'h0000028d, 5'd30, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000d2, 5'd27, 27'h000000ac, 5'd6, 27'h00000208, 32'h00000400,
  1'd1,  5'd9, 27'h0000014f, 5'd30, 27'h000000a6, 5'd17, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000034c, 5'd28, 27'h00000058, 5'd27, 27'h0000001c, 32'h00000400,
  1'd1,  5'd15, 27'h00000282, 5'd9, 27'h00000055, 5'd10, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002b5, 5'd6, 27'h00000138, 5'd16, 27'h000001e2, 32'h00000400,
  1'd1,  5'd18, 27'h000002f3, 5'd9, 27'h00000283, 5'd29, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001fd, 5'd17, 27'h0000016d, 5'd5, 27'h000001c1, 32'h00000400,
  1'd1,  5'd17, 27'h000003da, 5'd18, 27'h0000030b, 5'd19, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000086, 5'd19, 27'h0000024f, 5'd29, 27'h000000c9, 32'h00000400,
  1'd1,  5'd20, 27'h00000192, 5'd26, 27'h00000122, 5'd9, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000243, 5'd30, 27'h000001ec, 5'd17, 27'h0000009a, 32'h00000400,
  1'd1,  5'd18, 27'h0000023d, 5'd27, 27'h000002b9, 5'd28, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002b5, 5'd9, 27'h000000f8, 5'd6, 27'h000000a1, 32'h00000400,
  1'd1,  5'd30, 27'h0000010c, 5'd8, 27'h0000033a, 5'd16, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000255, 5'd5, 27'h000002a9, 5'd27, 27'h000003a7, 32'h00000400,
  1'd1,  5'd26, 27'h00000271, 5'd16, 27'h000003d7, 5'd10, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000017b, 5'd20, 27'h0000016d, 5'd18, 27'h000003b0, 32'h00000400,
  1'd1,  5'd26, 27'h000002cf, 5'd18, 27'h000001a2, 5'd26, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000037f, 5'd27, 27'h00000008, 5'd9, 27'h0000033f, 32'h00000400,
  1'd1,  5'd27, 27'h0000008e, 5'd26, 27'h000000da, 5'd19, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b8, 5'd26, 27'h00000103, 5'd30, 27'h000000b1, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000302, 5'd4, 27'h0000028b, 5'd4, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000001e, 5'd1, 27'h000001e8, 5'd11, 27'h000003b6, 32'h00000400,
  1'd1,  5'd2, 27'h000003fb, 5'd4, 27'h00000164, 5'd20, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000015e, 5'd12, 27'h0000025f, 5'd4, 27'h0000021e, 32'h00000400,
  1'd1,  5'd3, 27'h00000152, 5'd11, 27'h000003a0, 5'd14, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000007f, 5'd15, 27'h000001c7, 5'd23, 27'h00000028, 32'h00000400,
  1'd1,  5'd1, 27'h00000063, 5'd23, 27'h0000013f, 5'd2, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000344, 5'd20, 27'h00000396, 5'd11, 27'h000001ea, 32'h00000400,
  1'd1,  5'd4, 27'h00000289, 5'd22, 27'h0000032f, 5'd21, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035a, 5'd2, 27'h000002d1, 5'd0, 27'h0000025b, 32'h00000400,
  1'd1,  5'd12, 27'h0000035f, 5'd3, 27'h00000170, 5'd12, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000120, 5'd0, 27'h0000003c, 5'd20, 27'h0000031d, 32'h00000400,
  1'd1,  5'd10, 27'h00000207, 5'd13, 27'h00000140, 5'd0, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003aa, 5'd14, 27'h0000013b, 5'd14, 27'h00000351, 32'h00000400,
  1'd1,  5'd10, 27'h0000035a, 5'd14, 27'h00000023, 5'd21, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f1, 5'd24, 27'h0000018f, 5'd3, 27'h00000235, 32'h00000400,
  1'd1,  5'd14, 27'h00000016, 5'd21, 27'h00000269, 5'd11, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000008b, 5'd20, 27'h0000037e, 5'd21, 27'h00000135, 32'h00000400,
  1'd1,  5'd23, 27'h00000092, 5'd4, 27'h00000071, 5'd3, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000004e, 5'd3, 27'h000001a5, 5'd14, 27'h000000b4, 32'h00000400,
  1'd1,  5'd22, 27'h0000010d, 5'd3, 27'h00000342, 5'd23, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000204, 5'd14, 27'h00000214, 5'd2, 27'h0000039c, 32'h00000400,
  1'd1,  5'd24, 27'h0000000e, 5'd11, 27'h000003ef, 5'd13, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d2, 5'd14, 27'h000000e6, 5'd25, 27'h000000a9, 32'h00000400,
  1'd1,  5'd23, 27'h000000aa, 5'd21, 27'h000000d2, 5'd3, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000e8, 5'd24, 27'h000002bb, 5'd13, 27'h00000357, 32'h00000400,
  1'd1,  5'd21, 27'h00000261, 5'd22, 27'h00000011, 5'd25, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003fc, 5'd4, 27'h00000275, 5'd9, 27'h0000039f, 32'h00000400,
  1'd1,  5'd3, 27'h000001b3, 5'd1, 27'h0000022a, 5'd15, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000004f, 5'd1, 27'h00000071, 5'd28, 27'h0000015d, 32'h00000400,
  1'd1,  5'd1, 27'h000001f7, 5'd12, 27'h000002d2, 5'd7, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000008d, 5'd10, 27'h00000277, 5'd16, 27'h00000254, 32'h00000400,
  1'd1,  5'd3, 27'h000000bb, 5'd15, 27'h000000ac, 5'd25, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000009e, 5'd21, 27'h000000ab, 5'd9, 27'h00000274, 32'h00000400,
  1'd1,  5'd1, 27'h0000033a, 5'd22, 27'h00000017, 5'd19, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000379, 5'd24, 27'h00000265, 5'd30, 27'h00000112, 32'h00000400,
  1'd1,  5'd11, 27'h000003dd, 5'd4, 27'h00000003, 5'd8, 27'h000001ef, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000318, 5'd3, 27'h00000093, 5'd16, 27'h000003e5, 32'h00000400,
  1'd1,  5'd13, 27'h0000033d, 5'd1, 27'h000000e1, 5'd26, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002af, 5'd15, 27'h000000ef, 5'd7, 27'h000000fa, 32'h00000400,
  1'd1,  5'd15, 27'h00000120, 5'd15, 27'h00000185, 5'd18, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001a0, 5'd14, 27'h00000012, 5'd27, 27'h000001ec, 32'h00000400,
  1'd1,  5'd10, 27'h00000397, 5'd21, 27'h00000303, 5'd5, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e0, 5'd21, 27'h0000026d, 5'd15, 27'h000003ff, 32'h00000400,
  1'd1,  5'd10, 27'h00000269, 5'd24, 27'h00000035, 5'd26, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000137, 5'd0, 27'h00000259, 5'd7, 27'h00000210, 32'h00000400,
  1'd1,  5'd23, 27'h000000d4, 5'd4, 27'h000001e4, 5'd19, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000172, 5'd3, 27'h00000092, 5'd30, 27'h00000374, 32'h00000400,
  1'd1,  5'd24, 27'h000001c9, 5'd10, 27'h0000022d, 5'd8, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000038e, 5'd14, 27'h00000214, 5'd19, 27'h00000056, 32'h00000400,
  1'd1,  5'd21, 27'h00000201, 5'd10, 27'h00000192, 5'd29, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000026, 5'd21, 27'h0000036e, 5'd8, 27'h000001b5, 32'h00000400,
  1'd1,  5'd24, 27'h0000037f, 5'd20, 27'h000003fc, 5'd15, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c1, 5'd24, 27'h00000214, 5'd28, 27'h00000120, 32'h00000400,
  1'd1,  5'd2, 27'h00000179, 5'd8, 27'h00000353, 5'd4, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f3, 5'd5, 27'h000003e4, 5'd11, 27'h00000133, 32'h00000400,
  1'd1,  5'd3, 27'h000000f7, 5'd10, 27'h00000112, 5'd23, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000206, 5'd16, 27'h00000030, 5'd3, 27'h0000037a, 32'h00000400,
  1'd1,  5'd3, 27'h0000039f, 5'd19, 27'h00000385, 5'd12, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000007b, 5'd18, 27'h00000110, 5'd22, 27'h000002da, 32'h00000400,
  1'd1,  5'd4, 27'h0000001a, 5'd29, 27'h0000011d, 5'd4, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000355, 5'd29, 27'h00000176, 5'd12, 27'h000000f7, 32'h00000400,
  1'd1,  5'd2, 27'h000001c7, 5'd26, 27'h00000334, 5'd22, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000024c, 5'd7, 27'h000001c9, 5'd0, 27'h000001b2, 32'h00000400,
  1'd1,  5'd12, 27'h00000323, 5'd9, 27'h00000214, 5'd11, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000009e, 5'd7, 27'h000003cf, 5'd24, 27'h000002ef, 32'h00000400,
  1'd1,  5'd12, 27'h000003ab, 5'd17, 27'h0000008c, 5'd2, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000021e, 5'd16, 27'h0000035a, 5'd10, 27'h00000379, 32'h00000400,
  1'd1,  5'd11, 27'h00000341, 5'd17, 27'h00000118, 5'd22, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000366, 5'd25, 27'h00000392, 5'd4, 27'h00000036, 32'h00000400,
  1'd1,  5'd15, 27'h00000003, 5'd27, 27'h0000027b, 5'd10, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000016f, 5'd29, 27'h00000226, 5'd21, 27'h0000006c, 32'h00000400,
  1'd1,  5'd22, 27'h00000193, 5'd8, 27'h00000010, 5'd4, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000330, 5'd8, 27'h000003e6, 5'd14, 27'h000000b9, 32'h00000400,
  1'd1,  5'd21, 27'h00000047, 5'd5, 27'h000000bd, 5'd21, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000110, 5'd19, 27'h00000302, 5'd0, 27'h000000c4, 32'h00000400,
  1'd1,  5'd24, 27'h00000260, 5'd15, 27'h000003b1, 5'd12, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001bb, 5'd17, 27'h000000bf, 5'd25, 27'h000001ab, 32'h00000400,
  1'd1,  5'd22, 27'h000001b9, 5'd28, 27'h00000170, 5'd3, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000bd, 5'd30, 27'h0000023c, 5'd13, 27'h000000aa, 32'h00000400,
  1'd1,  5'd22, 27'h00000065, 5'd27, 27'h00000229, 5'd21, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000384, 5'd6, 27'h00000073, 5'd8, 27'h000003f8, 32'h00000400,
  1'd1,  5'd3, 27'h00000089, 5'd9, 27'h00000381, 5'd19, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001f4, 5'd8, 27'h000003f8, 5'd30, 27'h00000017, 32'h00000400,
  1'd1,  5'd3, 27'h00000316, 5'd17, 27'h0000037f, 5'd9, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000002, 5'd16, 27'h000003ce, 5'd19, 27'h000002ab, 32'h00000400,
  1'd1,  5'd1, 27'h000002cc, 5'd19, 27'h000002d1, 5'd28, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000343, 5'd29, 27'h0000019f, 5'd6, 27'h00000239, 32'h00000400,
  1'd1,  5'd3, 27'h00000260, 5'd27, 27'h000000de, 5'd18, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e0, 5'd28, 27'h000000b6, 5'd26, 27'h000000c1, 32'h00000400,
  1'd1,  5'd14, 27'h00000173, 5'd9, 27'h00000143, 5'd9, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000277, 5'd8, 27'h000000d7, 5'd15, 27'h000003b7, 32'h00000400,
  1'd1,  5'd11, 27'h00000205, 5'd8, 27'h000002a5, 5'd29, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000027f, 5'd15, 27'h000003b4, 5'd6, 27'h00000158, 32'h00000400,
  1'd1,  5'd12, 27'h000001dc, 5'd19, 27'h00000044, 5'd15, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000092, 5'd18, 27'h00000374, 5'd30, 27'h00000264, 32'h00000400,
  1'd1,  5'd13, 27'h00000272, 5'd30, 27'h00000301, 5'd8, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000038a, 5'd30, 27'h000000f4, 5'd17, 27'h000000da, 32'h00000400,
  1'd1,  5'd13, 27'h000002c2, 5'd26, 27'h0000024d, 5'd30, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000295, 5'd5, 27'h000002e8, 5'd6, 27'h000003ef, 32'h00000400,
  1'd1,  5'd23, 27'h00000174, 5'd6, 27'h0000027a, 5'd19, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000364, 5'd7, 27'h0000039d, 5'd28, 27'h00000373, 32'h00000400,
  1'd1,  5'd23, 27'h000003a3, 5'd17, 27'h000003a3, 5'd6, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000140, 5'd19, 27'h0000032a, 5'd19, 27'h0000001f, 32'h00000400,
  1'd1,  5'd23, 27'h000001f6, 5'd19, 27'h00000048, 5'd27, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000019e, 5'd25, 27'h000003b8, 5'd9, 27'h00000359, 32'h00000400,
  1'd1,  5'd24, 27'h00000089, 5'd26, 27'h000000fd, 5'd20, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000ae, 5'd27, 27'h000003cc, 5'd26, 27'h000000aa, 32'h00000400,
  1'd1,  5'd7, 27'h000000d6, 5'd0, 27'h00000154, 5'd7, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000040, 5'd3, 27'h000000d9, 5'd17, 27'h0000017c, 32'h00000400,
  1'd1,  5'd6, 27'h000002a2, 5'd0, 27'h00000342, 5'd26, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000201, 5'd12, 27'h00000173, 5'd0, 27'h00000175, 32'h00000400,
  1'd1,  5'd5, 27'h000001eb, 5'd12, 27'h000003d3, 5'd10, 27'h00000257, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000a6, 5'd10, 27'h00000241, 5'd23, 27'h00000257, 32'h00000400,
  1'd1,  5'd10, 27'h000000bb, 5'd25, 27'h000000e8, 5'd4, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000010, 5'd25, 27'h000002d8, 5'd12, 27'h000000a2, 32'h00000400,
  1'd1,  5'd7, 27'h0000007e, 5'd22, 27'h000003e6, 5'd23, 27'h0000009e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000024, 5'd3, 27'h00000235, 5'd10, 27'h000000e9, 32'h00000400,
  1'd1,  5'd17, 27'h00000116, 5'd1, 27'h000000ea, 5'd17, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f7, 5'd4, 27'h00000036, 5'd30, 27'h000000ef, 32'h00000400,
  1'd1,  5'd17, 27'h00000234, 5'd10, 27'h000001ba, 5'd4, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000008, 5'd15, 27'h000001e5, 5'd12, 27'h000003e2, 32'h00000400,
  1'd1,  5'd15, 27'h00000289, 5'd13, 27'h00000115, 5'd25, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003b2, 5'd23, 27'h000001f1, 5'd0, 27'h000000a7, 32'h00000400,
  1'd1,  5'd16, 27'h000003a0, 5'd24, 27'h00000190, 5'd11, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000024d, 5'd20, 27'h00000334, 5'd23, 27'h000000b3, 32'h00000400,
  1'd1,  5'd30, 27'h00000120, 5'd2, 27'h000002b8, 5'd1, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000e7, 5'd2, 27'h0000005c, 5'd11, 27'h00000382, 32'h00000400,
  1'd1,  5'd30, 27'h00000014, 5'd2, 27'h00000326, 5'd20, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ea, 5'd11, 27'h00000025, 5'd3, 27'h00000393, 32'h00000400,
  1'd1,  5'd27, 27'h00000067, 5'd12, 27'h00000291, 5'd15, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ba, 5'd14, 27'h00000381, 5'd23, 27'h000001d7, 32'h00000400,
  1'd1,  5'd26, 27'h0000017a, 5'd23, 27'h000001de, 5'd0, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003eb, 5'd23, 27'h000002da, 5'd12, 27'h00000073, 32'h00000400,
  1'd1,  5'd26, 27'h000001f3, 5'd22, 27'h0000019f, 5'd23, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000120, 5'd4, 27'h00000038, 5'd4, 27'h00000363, 32'h00000400,
  1'd1,  5'd6, 27'h000000d2, 5'd0, 27'h000002fe, 5'd12, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e6, 5'd4, 27'h000002b2, 5'd25, 27'h00000033, 32'h00000400,
  1'd1,  5'd6, 27'h00000049, 5'd12, 27'h000000d8, 5'd7, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000036c, 5'd14, 27'h0000006d, 5'd18, 27'h00000088, 32'h00000400,
  1'd1,  5'd6, 27'h00000369, 5'd15, 27'h00000151, 5'd28, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000017e, 5'd24, 27'h000002fa, 5'd7, 27'h000000c9, 32'h00000400,
  1'd1,  5'd7, 27'h000003f4, 5'd25, 27'h000002e5, 5'd19, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000024d, 5'd20, 27'h000002da, 5'd26, 27'h0000016d, 32'h00000400,
  1'd1,  5'd20, 27'h000001ec, 5'd4, 27'h00000015, 5'd4, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003cb, 5'd1, 27'h000000f8, 5'd14, 27'h000001d6, 32'h00000400,
  1'd1,  5'd19, 27'h000002f5, 5'd3, 27'h000003a8, 5'd23, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000266, 5'd15, 27'h0000008e, 5'd7, 27'h000000dc, 32'h00000400,
  1'd1,  5'd15, 27'h00000221, 5'd12, 27'h00000159, 5'd20, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c3, 5'd13, 27'h0000010f, 5'd27, 27'h000003be, 32'h00000400,
  1'd1,  5'd17, 27'h00000333, 5'd22, 27'h000000d9, 5'd9, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000253, 5'd24, 27'h00000194, 5'd15, 27'h000003f4, 32'h00000400,
  1'd1,  5'd18, 27'h0000013d, 5'd22, 27'h000002f3, 5'd27, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001dd, 5'd2, 27'h000000dc, 5'd7, 27'h0000027e, 32'h00000400,
  1'd1,  5'd27, 27'h00000332, 5'd4, 27'h00000002, 5'd19, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003bc, 5'd0, 27'h000002d6, 5'd25, 27'h000003f3, 32'h00000400,
  1'd1,  5'd28, 27'h0000014f, 5'd11, 27'h000003d3, 5'd6, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f0, 5'd10, 27'h00000188, 5'd20, 27'h00000201, 32'h00000400,
  1'd1,  5'd27, 27'h00000066, 5'd13, 27'h00000352, 5'd26, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b7, 5'd22, 27'h000002e0, 5'd8, 27'h0000010a, 32'h00000400,
  1'd1,  5'd28, 27'h00000354, 5'd21, 27'h00000242, 5'd19, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000028a, 5'd24, 27'h0000005d, 5'd30, 27'h000000b4, 32'h00000400,
  1'd1,  5'd9, 27'h0000033d, 5'd7, 27'h00000312, 5'd1, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000012, 5'd6, 27'h00000163, 5'd11, 27'h0000027c, 32'h00000400,
  1'd1,  5'd9, 27'h0000007b, 5'd9, 27'h000001ee, 5'd23, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003d7, 5'd16, 27'h00000074, 5'd3, 27'h000003c1, 32'h00000400,
  1'd1,  5'd6, 27'h00000184, 5'd16, 27'h000002b7, 5'd10, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000165, 5'd16, 27'h00000153, 5'd22, 27'h000002e7, 32'h00000400,
  1'd1,  5'd5, 27'h0000010a, 5'd27, 27'h000002be, 5'd4, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000054, 5'd27, 27'h0000013e, 5'd12, 27'h000000e7, 32'h00000400,
  1'd1,  5'd5, 27'h000000e0, 5'd26, 27'h000002e3, 5'd21, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000011, 5'd7, 27'h00000316, 5'd2, 27'h0000017f, 32'h00000400,
  1'd1,  5'd17, 27'h00000211, 5'd5, 27'h000002cf, 5'd10, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e1, 5'd10, 27'h0000013e, 5'd23, 27'h0000039b, 32'h00000400,
  1'd1,  5'd20, 27'h000000b5, 5'd17, 27'h00000268, 5'd1, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000084, 5'd19, 27'h00000400, 5'd11, 27'h0000017a, 32'h00000400,
  1'd1,  5'd16, 27'h00000135, 5'd16, 27'h00000360, 5'd23, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000264, 5'd28, 27'h0000010e, 5'd2, 27'h000000a7, 32'h00000400,
  1'd1,  5'd16, 27'h000002d8, 5'd30, 27'h00000256, 5'd12, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000050, 5'd27, 27'h00000084, 5'd24, 27'h00000301, 32'h00000400,
  1'd1,  5'd26, 27'h00000107, 5'd7, 27'h000002a4, 5'd2, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000181, 5'd5, 27'h00000107, 5'd13, 27'h000002b2, 32'h00000400,
  1'd1,  5'd29, 27'h00000130, 5'd9, 27'h00000072, 5'd22, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000303, 5'd17, 27'h00000276, 5'd2, 27'h0000019e, 32'h00000400,
  1'd1,  5'd29, 27'h00000056, 5'd16, 27'h00000242, 5'd11, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000026d, 5'd17, 27'h00000278, 5'd24, 27'h000003e3, 32'h00000400,
  1'd1,  5'd29, 27'h0000031a, 5'd29, 27'h0000027c, 5'd4, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000007c, 5'd26, 27'h00000360, 5'd12, 27'h00000253, 32'h00000400,
  1'd1,  5'd29, 27'h00000133, 5'd30, 27'h00000270, 5'd24, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000183, 5'd7, 27'h000000e9, 5'd8, 27'h00000284, 32'h00000400,
  1'd1,  5'd9, 27'h0000017d, 5'd8, 27'h00000353, 5'd18, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001c5, 5'd9, 27'h000000a8, 5'd30, 27'h00000308, 32'h00000400,
  1'd1,  5'd7, 27'h0000016d, 5'd16, 27'h000000f0, 5'd6, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000312, 5'd18, 27'h00000376, 5'd18, 27'h00000382, 32'h00000400,
  1'd1,  5'd6, 27'h000001ab, 5'd19, 27'h000001a1, 5'd25, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000034d, 5'd28, 27'h0000037f, 5'd9, 27'h000001ed, 32'h00000400,
  1'd1,  5'd7, 27'h00000310, 5'd27, 27'h000001a2, 5'd20, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000004a, 5'd30, 27'h00000151, 5'd26, 27'h00000166, 32'h00000400,
  1'd1,  5'd16, 27'h00000061, 5'd7, 27'h00000197, 5'd6, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000247, 5'd5, 27'h00000197, 5'd18, 27'h00000335, 32'h00000400,
  1'd1,  5'd15, 27'h00000290, 5'd5, 27'h00000234, 5'd26, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000263, 5'd18, 27'h00000051, 5'd8, 27'h000001a1, 32'h00000400,
  1'd1,  5'd18, 27'h00000236, 5'd17, 27'h00000226, 5'd17, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000255, 5'd20, 27'h0000024b, 5'd28, 27'h000000a3, 32'h00000400,
  1'd1,  5'd19, 27'h00000388, 5'd29, 27'h000001cf, 5'd8, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002aa, 5'd29, 27'h00000088, 5'd16, 27'h000002b7, 32'h00000400,
  1'd1,  5'd18, 27'h000001d9, 5'd30, 27'h00000135, 5'd27, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a5, 5'd7, 27'h0000019d, 5'd8, 27'h000001c6, 32'h00000400,
  1'd1,  5'd26, 27'h0000000c, 5'd9, 27'h000001b9, 5'd18, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a8, 5'd9, 27'h00000238, 5'd26, 27'h000001b9, 32'h00000400,
  1'd1,  5'd26, 27'h000000af, 5'd20, 27'h00000266, 5'd7, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000015c, 5'd19, 27'h00000396, 5'd20, 27'h0000021b, 32'h00000400,
  1'd1,  5'd30, 27'h000000d3, 5'd19, 27'h00000112, 5'd30, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000042, 5'd29, 27'h00000252, 5'd9, 27'h000002a6, 32'h00000400,
  1'd1,  5'd28, 27'h00000010, 5'd25, 27'h000003f4, 5'd19, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003ef, 5'd28, 27'h00000148, 5'd26, 27'h00000286, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000000da, 5'd1, 27'h000003ef, 5'd1, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000209, 5'd0, 27'h000002a0, 5'd10, 27'h000003ca, 32'h00000400,
  1'd1,  5'd4, 27'h000001a4, 5'd1, 27'h000002ea, 5'd25, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000176, 5'd13, 27'h000001d1, 5'd2, 27'h000003b3, 32'h00000400,
  1'd1,  5'd0, 27'h0000014a, 5'd14, 27'h000001eb, 5'd13, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000022d, 5'd12, 27'h000001d3, 5'd24, 27'h000002d0, 32'h00000400,
  1'd1,  5'd1, 27'h00000382, 5'd23, 27'h00000126, 5'd5, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000095, 5'd21, 27'h0000035d, 5'd11, 27'h000003f4, 32'h00000400,
  1'd1,  5'd5, 27'h00000053, 5'd21, 27'h000000f0, 5'd22, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000cf, 5'd4, 27'h00000389, 5'd1, 27'h0000013c, 32'h00000400,
  1'd1,  5'd11, 27'h00000226, 5'd3, 27'h000000ea, 5'd14, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d1, 5'd3, 27'h000001b9, 5'd20, 27'h000003cc, 32'h00000400,
  1'd1,  5'd14, 27'h00000385, 5'd14, 27'h00000201, 5'd4, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000012d, 5'd12, 27'h000000ee, 5'd11, 27'h00000041, 32'h00000400,
  1'd1,  5'd13, 27'h0000001f, 5'd15, 27'h0000006f, 5'd23, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000377, 5'd23, 27'h000002af, 5'd1, 27'h000001f4, 32'h00000400,
  1'd1,  5'd11, 27'h0000037e, 5'd23, 27'h00000308, 5'd13, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000007a, 5'd23, 27'h00000214, 5'd25, 27'h00000098, 32'h00000400,
  1'd1,  5'd24, 27'h000001dd, 5'd1, 27'h000003b6, 5'd1, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000036b, 5'd3, 27'h000003fd, 5'd15, 27'h00000027, 32'h00000400,
  1'd1,  5'd24, 27'h000002c3, 5'd0, 27'h000003fb, 5'd24, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000003d, 5'd11, 27'h0000024c, 5'd4, 27'h00000379, 32'h00000400,
  1'd1,  5'd21, 27'h000001dd, 5'd11, 27'h0000032c, 5'd14, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000001c, 5'd12, 27'h000000db, 5'd24, 27'h000003d3, 32'h00000400,
  1'd1,  5'd24, 27'h00000124, 5'd21, 27'h000001ef, 5'd4, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032a, 5'd23, 27'h000001ad, 5'd12, 27'h0000018c, 32'h00000400,
  1'd1,  5'd22, 27'h0000028e, 5'd25, 27'h0000013b, 5'd24, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000015, 5'd0, 27'h0000021b, 5'd7, 27'h000002b5, 32'h00000400,
  1'd1,  5'd4, 27'h00000304, 5'd2, 27'h00000141, 5'd16, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002e0, 5'd1, 27'h00000280, 5'd27, 27'h000000ec, 32'h00000400,
  1'd1,  5'd1, 27'h0000006a, 5'd13, 27'h00000194, 5'd8, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002ae, 5'd13, 27'h000003a6, 5'd18, 27'h000003df, 32'h00000400,
  1'd1,  5'd0, 27'h0000025c, 5'd11, 27'h0000027b, 5'd26, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000113, 5'd22, 27'h00000216, 5'd7, 27'h00000130, 32'h00000400,
  1'd1,  5'd1, 27'h00000038, 5'd24, 27'h000003f6, 5'd18, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f7, 5'd21, 27'h000003b4, 5'd28, 27'h00000102, 32'h00000400,
  1'd1,  5'd15, 27'h00000037, 5'd4, 27'h000001f5, 5'd7, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000334, 5'd0, 27'h000001c9, 5'd17, 27'h00000194, 32'h00000400,
  1'd1,  5'd14, 27'h00000074, 5'd2, 27'h00000250, 5'd29, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000367, 5'd12, 27'h00000257, 5'd9, 27'h000003f7, 32'h00000400,
  1'd1,  5'd11, 27'h00000378, 5'd12, 27'h000000e3, 5'd15, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011c, 5'd14, 27'h000001c0, 5'd30, 27'h000002b5, 32'h00000400,
  1'd1,  5'd13, 27'h00000005, 5'd24, 27'h00000170, 5'd6, 27'h0000021e, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003eb, 5'd25, 27'h000000d0, 5'd18, 27'h00000169, 32'h00000400,
  1'd1,  5'd13, 27'h00000392, 5'd23, 27'h0000010f, 5'd26, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000003, 5'd2, 27'h000003c2, 5'd10, 27'h000000c9, 32'h00000400,
  1'd1,  5'd25, 27'h000002bf, 5'd0, 27'h00000198, 5'd15, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000310, 5'd4, 27'h00000343, 5'd26, 27'h00000064, 32'h00000400,
  1'd1,  5'd23, 27'h0000023a, 5'd11, 27'h000001ab, 5'd6, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000001b, 5'd10, 27'h000002f2, 5'd17, 27'h00000267, 32'h00000400,
  1'd1,  5'd25, 27'h0000027c, 5'd11, 27'h000002ed, 5'd27, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000021f, 5'd25, 27'h00000328, 5'd7, 27'h000003ea, 32'h00000400,
  1'd1,  5'd22, 27'h00000175, 5'd21, 27'h000003dd, 5'd18, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000295, 5'd21, 27'h0000017a, 5'd27, 27'h00000222, 32'h00000400,
  1'd1,  5'd2, 27'h0000037b, 5'd8, 27'h00000117, 5'd1, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003be, 5'd9, 27'h0000019e, 5'd14, 27'h00000033, 32'h00000400,
  1'd1,  5'd1, 27'h000000ed, 5'd5, 27'h0000037e, 5'd25, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000c3, 5'd19, 27'h00000398, 5'd4, 27'h0000039c, 32'h00000400,
  1'd1,  5'd1, 27'h00000219, 5'd16, 27'h000002b2, 5'd13, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000008f, 5'd20, 27'h00000247, 5'd24, 27'h0000035b, 32'h00000400,
  1'd1,  5'd4, 27'h0000037d, 5'd26, 27'h000001cb, 5'd2, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000006e, 5'd29, 27'h00000168, 5'd14, 27'h000001a6, 32'h00000400,
  1'd1,  5'd3, 27'h000001f7, 5'd29, 27'h00000108, 5'd24, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003a8, 5'd9, 27'h00000046, 5'd2, 27'h000001e3, 32'h00000400,
  1'd1,  5'd14, 27'h000002c8, 5'd8, 27'h0000020a, 5'd14, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000270, 5'd7, 27'h0000033c, 5'd22, 27'h0000012c, 32'h00000400,
  1'd1,  5'd12, 27'h00000271, 5'd18, 27'h0000011b, 5'd0, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002d6, 5'd19, 27'h0000014b, 5'd10, 27'h000003b9, 32'h00000400,
  1'd1,  5'd11, 27'h000003e7, 5'd18, 27'h000003fd, 5'd23, 27'h000002a0, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000337, 5'd26, 27'h0000018c, 5'd4, 27'h00000194, 32'h00000400,
  1'd1,  5'd14, 27'h0000038d, 5'd26, 27'h0000036d, 5'd11, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000180, 5'd28, 27'h0000008d, 5'd22, 27'h000003da, 32'h00000400,
  1'd1,  5'd22, 27'h000000e4, 5'd7, 27'h00000043, 5'd0, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000184, 5'd8, 27'h000001d9, 5'd12, 27'h00000351, 32'h00000400,
  1'd1,  5'd23, 27'h00000006, 5'd7, 27'h00000220, 5'd21, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002a9, 5'd20, 27'h00000035, 5'd3, 27'h0000017c, 32'h00000400,
  1'd1,  5'd24, 27'h000001ec, 5'd15, 27'h00000258, 5'd12, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001a1, 5'd16, 27'h00000120, 5'd25, 27'h00000102, 32'h00000400,
  1'd1,  5'd23, 27'h000002df, 5'd26, 27'h000000d5, 5'd4, 27'h00000201, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000075, 5'd30, 27'h00000347, 5'd10, 27'h00000248, 32'h00000400,
  1'd1,  5'd24, 27'h000003d0, 5'd27, 27'h00000390, 5'd22, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000124, 5'd8, 27'h00000221, 5'd8, 27'h0000007f, 32'h00000400,
  1'd1,  5'd0, 27'h0000003a, 5'd7, 27'h0000029b, 5'd18, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000017c, 5'd9, 27'h0000032b, 5'd28, 27'h00000156, 32'h00000400,
  1'd1,  5'd5, 27'h00000048, 5'd16, 27'h00000215, 5'd9, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000380, 5'd20, 27'h00000006, 5'd18, 27'h00000159, 32'h00000400,
  1'd1,  5'd1, 27'h00000311, 5'd18, 27'h0000034a, 5'd28, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000208, 5'd29, 27'h0000037d, 5'd9, 27'h00000024, 32'h00000400,
  1'd1,  5'd1, 27'h000003dc, 5'd29, 27'h00000338, 5'd17, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000318, 5'd30, 27'h000000a3, 5'd28, 27'h000003e1, 32'h00000400,
  1'd1,  5'd13, 27'h000002e9, 5'd9, 27'h00000219, 5'd8, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000025b, 5'd7, 27'h000001ed, 5'd16, 27'h0000004d, 32'h00000400,
  1'd1,  5'd11, 27'h0000018f, 5'd7, 27'h000000e8, 5'd30, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f2, 5'd18, 27'h0000003f, 5'd8, 27'h00000090, 32'h00000400,
  1'd1,  5'd14, 27'h000003b9, 5'd17, 27'h0000006d, 5'd16, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000241, 5'd16, 27'h000001cf, 5'd30, 27'h0000004a, 32'h00000400,
  1'd1,  5'd14, 27'h000001fd, 5'd27, 27'h000002c6, 5'd9, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003c6, 5'd27, 27'h000003c9, 5'd19, 27'h000003ce, 32'h00000400,
  1'd1,  5'd12, 27'h00000091, 5'd29, 27'h00000225, 5'd27, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000189, 5'd8, 27'h000001e5, 5'd10, 27'h000000c9, 32'h00000400,
  1'd1,  5'd23, 27'h000003cc, 5'd9, 27'h00000120, 5'd20, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000163, 5'd6, 27'h0000007d, 5'd29, 27'h000003ff, 32'h00000400,
  1'd1,  5'd22, 27'h00000059, 5'd19, 27'h000002fd, 5'd6, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001fd, 5'd17, 27'h0000012a, 5'd16, 27'h00000210, 32'h00000400,
  1'd1,  5'd25, 27'h00000083, 5'd18, 27'h00000315, 5'd29, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000134, 5'd29, 27'h0000003e, 5'd7, 27'h0000026c, 32'h00000400,
  1'd1,  5'd22, 27'h0000038a, 5'd28, 27'h000002e6, 5'd18, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000b2, 5'd26, 27'h0000006d, 5'd28, 27'h000003f4, 32'h00000400,
  1'd1,  5'd6, 27'h00000173, 5'd1, 27'h0000030b, 5'd7, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000323, 5'd4, 27'h00000080, 5'd18, 27'h000003f5, 32'h00000400,
  1'd1,  5'd5, 27'h00000108, 5'd2, 27'h0000014f, 5'd30, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000360, 5'd13, 27'h0000032a, 5'd1, 27'h0000036c, 32'h00000400,
  1'd1,  5'd10, 27'h000000e4, 5'd11, 27'h0000024f, 5'd11, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000104, 5'd11, 27'h00000329, 5'd23, 27'h00000127, 32'h00000400,
  1'd1,  5'd9, 27'h0000006a, 5'd24, 27'h000002e9, 5'd0, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000329, 5'd24, 27'h00000352, 5'd12, 27'h00000345, 32'h00000400,
  1'd1,  5'd6, 27'h00000012, 5'd22, 27'h00000258, 5'd22, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c2, 5'd1, 27'h00000270, 5'd9, 27'h0000014f, 32'h00000400,
  1'd1,  5'd19, 27'h000003b0, 5'd3, 27'h000002bb, 5'd15, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000eb, 5'd3, 27'h0000013b, 5'd27, 27'h000001de, 32'h00000400,
  1'd1,  5'd17, 27'h00000292, 5'd15, 27'h000000a0, 5'd4, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000008d, 5'd12, 27'h00000056, 5'd10, 27'h000003fb, 32'h00000400,
  1'd1,  5'd16, 27'h00000308, 5'd13, 27'h000001ff, 5'd25, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000123, 5'd21, 27'h00000092, 5'd2, 27'h000001dd, 32'h00000400,
  1'd1,  5'd17, 27'h00000228, 5'd24, 27'h000002d4, 5'd14, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a6, 5'd23, 27'h0000039e, 5'd24, 27'h0000016e, 32'h00000400,
  1'd1,  5'd25, 27'h00000383, 5'd0, 27'h0000031f, 5'd2, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000012d, 5'd5, 27'h00000087, 5'd10, 27'h000001e0, 32'h00000400,
  1'd1,  5'd29, 27'h000002bf, 5'd3, 27'h00000252, 5'd21, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001aa, 5'd10, 27'h000001b6, 5'd2, 27'h000000aa, 32'h00000400,
  1'd1,  5'd28, 27'h0000036d, 5'd10, 27'h0000038a, 5'd13, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000138, 5'd11, 27'h00000093, 5'd24, 27'h0000007e, 32'h00000400,
  1'd1,  5'd27, 27'h000002ba, 5'd21, 27'h000002e3, 5'd1, 27'h000002d6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003c6, 5'd22, 27'h00000156, 5'd10, 27'h00000209, 32'h00000400,
  1'd1,  5'd27, 27'h00000300, 5'd23, 27'h0000017f, 5'd22, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000008b, 5'd2, 27'h000002fc, 5'd2, 27'h00000093, 32'h00000400,
  1'd1,  5'd8, 27'h00000041, 5'd3, 27'h0000024d, 5'd11, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000bc, 5'd3, 27'h00000234, 5'd23, 27'h00000365, 32'h00000400,
  1'd1,  5'd5, 27'h000000ce, 5'd12, 27'h0000032a, 5'd5, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000043, 5'd14, 27'h000003e8, 5'd17, 27'h00000258, 32'h00000400,
  1'd1,  5'd5, 27'h0000032d, 5'd12, 27'h000001db, 5'd29, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000bd, 5'd22, 27'h0000011e, 5'd8, 27'h000003c3, 32'h00000400,
  1'd1,  5'd10, 27'h0000012f, 5'd22, 27'h00000021, 5'd17, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000115, 5'd20, 27'h0000037b, 5'd30, 27'h0000026b, 32'h00000400,
  1'd1,  5'd17, 27'h00000265, 5'd2, 27'h000001ea, 5'd0, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000383, 5'd2, 27'h00000105, 5'd10, 27'h0000031e, 32'h00000400,
  1'd1,  5'd16, 27'h000000d0, 5'd3, 27'h00000076, 5'd24, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c7, 5'd11, 27'h0000022b, 5'd7, 27'h00000157, 32'h00000400,
  1'd1,  5'd18, 27'h000003cc, 5'd11, 27'h00000078, 5'd19, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a1, 5'd11, 27'h000003a2, 5'd30, 27'h000003b3, 32'h00000400,
  1'd1,  5'd20, 27'h000001f6, 5'd21, 27'h00000218, 5'd5, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000003c, 5'd22, 27'h000001fa, 5'd20, 27'h0000003e, 32'h00000400,
  1'd1,  5'd17, 27'h00000029, 5'd25, 27'h00000042, 5'd30, 27'h000002e8, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001c0, 5'd2, 27'h0000030e, 5'd7, 27'h0000007a, 32'h00000400,
  1'd1,  5'd30, 27'h000002ae, 5'd4, 27'h000002c4, 5'd17, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000152, 5'd2, 27'h00000045, 5'd29, 27'h000001f0, 32'h00000400,
  1'd1,  5'd28, 27'h000003b5, 5'd13, 27'h000001ef, 5'd6, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000056, 5'd12, 27'h000002c3, 5'd15, 27'h000002a7, 32'h00000400,
  1'd1,  5'd28, 27'h0000024b, 5'd13, 27'h00000170, 5'd29, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000373, 5'd22, 27'h00000344, 5'd5, 27'h000003af, 32'h00000400,
  1'd1,  5'd28, 27'h00000103, 5'd22, 27'h00000151, 5'd16, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000027d, 5'd25, 27'h00000176, 5'd30, 27'h000000af, 32'h00000400,
  1'd1,  5'd5, 27'h00000175, 5'd7, 27'h0000033f, 5'd2, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e3, 5'd5, 27'h00000224, 5'd10, 27'h0000035d, 32'h00000400,
  1'd1,  5'd5, 27'h0000023e, 5'd5, 27'h00000222, 5'd25, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e6, 5'd15, 27'h0000037d, 5'd2, 27'h0000028e, 32'h00000400,
  1'd1,  5'd5, 27'h000002ac, 5'd16, 27'h0000032c, 5'd11, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000003f, 5'd17, 27'h00000256, 5'd25, 27'h000002ea, 32'h00000400,
  1'd1,  5'd8, 27'h000001bf, 5'd30, 27'h0000037b, 5'd4, 27'h00000275, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e3, 5'd26, 27'h000000ed, 5'd13, 27'h0000020b, 32'h00000400,
  1'd1,  5'd9, 27'h000001f3, 5'd29, 27'h00000297, 5'd22, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029e, 5'd6, 27'h000003ad, 5'd4, 27'h00000298, 32'h00000400,
  1'd1,  5'd17, 27'h00000341, 5'd6, 27'h0000014f, 5'd10, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000179, 5'd9, 27'h000000dd, 5'd22, 27'h0000009d, 32'h00000400,
  1'd1,  5'd18, 27'h000001c1, 5'd17, 27'h000000dc, 5'd1, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000107, 5'd19, 27'h0000001c, 5'd11, 27'h00000157, 32'h00000400,
  1'd1,  5'd18, 27'h000000c3, 5'd16, 27'h00000282, 5'd22, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001b1, 5'd26, 27'h0000030a, 5'd4, 27'h0000007f, 32'h00000400,
  1'd1,  5'd17, 27'h00000188, 5'd29, 27'h00000389, 5'd10, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000295, 5'd27, 27'h00000108, 5'd22, 27'h0000003c, 32'h00000400,
  1'd1,  5'd26, 27'h00000126, 5'd10, 27'h0000011e, 5'd2, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001de, 5'd7, 27'h000000ad, 5'd13, 27'h000003e3, 32'h00000400,
  1'd1,  5'd27, 27'h0000009c, 5'd9, 27'h00000096, 5'd25, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e0, 5'd18, 27'h0000008b, 5'd3, 27'h00000179, 32'h00000400,
  1'd1,  5'd28, 27'h00000397, 5'd20, 27'h0000000e, 5'd10, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000090, 5'd19, 27'h000000f4, 5'd23, 27'h0000008e, 32'h00000400,
  1'd1,  5'd28, 27'h000001a7, 5'd27, 27'h00000208, 5'd0, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000020c, 5'd26, 27'h00000187, 5'd12, 27'h00000397, 32'h00000400,
  1'd1,  5'd27, 27'h00000190, 5'd30, 27'h000000fd, 5'd23, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002cf, 5'd5, 27'h0000018f, 5'd5, 27'h000003ee, 32'h00000400,
  1'd1,  5'd8, 27'h000000db, 5'd7, 27'h000002e4, 5'd17, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000036, 5'd8, 27'h000002bf, 5'd30, 27'h00000210, 32'h00000400,
  1'd1,  5'd5, 27'h000001aa, 5'd16, 27'h0000025a, 5'd9, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000116, 5'd16, 27'h0000005b, 5'd18, 27'h00000060, 32'h00000400,
  1'd1,  5'd5, 27'h000003c1, 5'd16, 27'h000002d3, 5'd27, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e4, 5'd28, 27'h00000301, 5'd7, 27'h00000050, 32'h00000400,
  1'd1,  5'd5, 27'h00000219, 5'd27, 27'h000000ae, 5'd19, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000f8, 5'd28, 27'h00000170, 5'd30, 27'h000001e7, 32'h00000400,
  1'd1,  5'd19, 27'h00000005, 5'd9, 27'h0000027f, 5'd7, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000003d, 5'd5, 27'h000001c6, 5'd18, 27'h0000036e, 32'h00000400,
  1'd1,  5'd19, 27'h00000188, 5'd6, 27'h000002ab, 5'd28, 27'h000000fc, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000308, 5'd18, 27'h000002bd, 5'd7, 27'h0000013b, 32'h00000400,
  1'd1,  5'd20, 27'h000000d9, 5'd16, 27'h00000258, 5'd18, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002cb, 5'd16, 27'h0000010b, 5'd28, 27'h00000337, 32'h00000400,
  1'd1,  5'd16, 27'h00000131, 5'd25, 27'h000003f7, 5'd7, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000057, 5'd27, 27'h0000022a, 5'd18, 27'h000003f8, 32'h00000400,
  1'd1,  5'd16, 27'h00000183, 5'd26, 27'h000000a5, 5'd26, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003ea, 5'd7, 27'h00000023, 5'd9, 27'h000000d7, 32'h00000400,
  1'd1,  5'd26, 27'h0000005e, 5'd7, 27'h00000018, 5'd16, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000120, 5'd9, 27'h00000123, 5'd27, 27'h0000032e, 32'h00000400,
  1'd1,  5'd29, 27'h00000051, 5'd17, 27'h00000009, 5'd7, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002e2, 5'd20, 27'h00000054, 5'd19, 27'h0000037f, 32'h00000400,
  1'd1,  5'd27, 27'h000002e8, 5'd16, 27'h0000027c, 5'd30, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002fd, 5'd26, 27'h0000033e, 5'd9, 27'h00000189, 32'h00000400,
  1'd1,  5'd29, 27'h000000d8, 5'd26, 27'h000003c4, 5'd16, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ea, 5'd27, 27'h00000162, 5'd26, 27'h00000031, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000037a, 5'd2, 27'h0000002a, 5'd3, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000a3, 5'd3, 27'h000000c7, 5'd13, 27'h000001ab, 32'h00000400,
  1'd1,  5'd0, 27'h00000361, 5'd2, 27'h0000018d, 5'd24, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000197, 5'd11, 27'h000000f4, 5'd2, 27'h000000e5, 32'h00000400,
  1'd1,  5'd3, 27'h0000006e, 5'd14, 27'h000002ca, 5'd10, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000018c, 5'd13, 27'h000001a6, 5'd23, 27'h0000020b, 32'h00000400,
  1'd1,  5'd2, 27'h000000a2, 5'd23, 27'h0000022f, 5'd2, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003aa, 5'd24, 27'h000003c8, 5'd12, 27'h00000373, 32'h00000400,
  1'd1,  5'd0, 27'h00000299, 5'd22, 27'h0000003b, 5'd24, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000067, 5'd2, 27'h000002af, 5'd1, 27'h000002a3, 32'h00000400,
  1'd1,  5'd14, 27'h000000a0, 5'd0, 27'h000003dc, 5'd11, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002d, 5'd4, 27'h0000019a, 5'd22, 27'h000002b2, 32'h00000400,
  1'd1,  5'd14, 27'h00000020, 5'd11, 27'h0000029a, 5'd4, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000200, 5'd15, 27'h000000ce, 5'd14, 27'h00000011, 32'h00000400,
  1'd1,  5'd14, 27'h00000399, 5'd12, 27'h00000334, 5'd24, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002dd, 5'd25, 27'h000000e4, 5'd1, 27'h00000347, 32'h00000400,
  1'd1,  5'd11, 27'h000003ff, 5'd22, 27'h0000017f, 5'd11, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000154, 5'd25, 27'h000002b9, 5'd22, 27'h000001a2, 32'h00000400,
  1'd1,  5'd24, 27'h0000021e, 5'd0, 27'h00000092, 5'd4, 27'h00000154, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000358, 5'd0, 27'h0000031c, 5'd11, 27'h000000b8, 32'h00000400,
  1'd1,  5'd23, 27'h000003ea, 5'd5, 27'h000000a0, 5'd21, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000262, 5'd11, 27'h00000181, 5'd4, 27'h000000af, 32'h00000400,
  1'd1,  5'd23, 27'h000003b2, 5'd12, 27'h000001e6, 5'd12, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ba, 5'd15, 27'h0000009a, 5'd21, 27'h000002c5, 32'h00000400,
  1'd1,  5'd24, 27'h00000141, 5'd23, 27'h000000cf, 5'd3, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000c0, 5'd21, 27'h00000349, 5'd12, 27'h0000032a, 32'h00000400,
  1'd1,  5'd24, 27'h00000353, 5'd22, 27'h00000239, 5'd25, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000013f, 5'd5, 27'h00000012, 5'd9, 27'h00000303, 32'h00000400,
  1'd1,  5'd1, 27'h00000055, 5'd4, 27'h000000de, 5'd18, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001a8, 5'd3, 27'h0000023c, 5'd30, 27'h000000ea, 32'h00000400,
  1'd1,  5'd0, 27'h0000010a, 5'd14, 27'h0000006b, 5'd10, 27'h00000155, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000bb, 5'd13, 27'h000000b3, 5'd19, 27'h000000e5, 32'h00000400,
  1'd1,  5'd2, 27'h00000302, 5'd12, 27'h000003a9, 5'd28, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002e5, 5'd22, 27'h0000037b, 5'd6, 27'h00000052, 32'h00000400,
  1'd1,  5'd2, 27'h000000dd, 5'd24, 27'h0000007e, 5'd16, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000376, 5'd20, 27'h0000035e, 5'd28, 27'h00000256, 32'h00000400,
  1'd1,  5'd14, 27'h00000149, 5'd1, 27'h0000014e, 5'd10, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000035, 5'd0, 27'h0000006c, 5'd18, 27'h00000146, 32'h00000400,
  1'd1,  5'd10, 27'h000002ad, 5'd1, 27'h0000017b, 5'd30, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000107, 5'd12, 27'h00000118, 5'd5, 27'h000001ff, 32'h00000400,
  1'd1,  5'd11, 27'h00000053, 5'd11, 27'h00000212, 5'd17, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001ae, 5'd14, 27'h000003de, 5'd29, 27'h000001d4, 32'h00000400,
  1'd1,  5'd10, 27'h0000022f, 5'd22, 27'h00000336, 5'd9, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000007d, 5'd24, 27'h0000009b, 5'd15, 27'h000003c3, 32'h00000400,
  1'd1,  5'd11, 27'h00000134, 5'd23, 27'h0000015e, 5'd25, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000028c, 5'd1, 27'h0000019d, 5'd9, 27'h0000006a, 32'h00000400,
  1'd1,  5'd22, 27'h000001df, 5'd0, 27'h0000002f, 5'd16, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000105, 5'd0, 27'h000000f6, 5'd26, 27'h000002a7, 32'h00000400,
  1'd1,  5'd24, 27'h000003bb, 5'd11, 27'h000003e9, 5'd6, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001c, 5'd14, 27'h0000037f, 5'd15, 27'h000002b9, 32'h00000400,
  1'd1,  5'd21, 27'h0000029b, 5'd12, 27'h0000029f, 5'd26, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000030b, 5'd22, 27'h00000296, 5'd8, 27'h000003af, 32'h00000400,
  1'd1,  5'd21, 27'h0000014c, 5'd24, 27'h000002a3, 5'd15, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000093, 5'd24, 27'h000001c4, 5'd28, 27'h000002b7, 32'h00000400,
  1'd1,  5'd2, 27'h000002d5, 5'd6, 27'h0000011c, 5'd1, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a8, 5'd8, 27'h00000337, 5'd14, 27'h00000382, 32'h00000400,
  1'd1,  5'd2, 27'h00000007, 5'd6, 27'h000002d7, 5'd20, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e7, 5'd20, 27'h000000c5, 5'd4, 27'h00000302, 32'h00000400,
  1'd1,  5'd4, 27'h00000371, 5'd15, 27'h000003a3, 5'd12, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001cd, 5'd15, 27'h000003ef, 5'd23, 27'h000002e6, 32'h00000400,
  1'd1,  5'd4, 27'h0000025a, 5'd28, 27'h000000ff, 5'd0, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ca, 5'd28, 27'h0000005c, 5'd12, 27'h00000056, 32'h00000400,
  1'd1,  5'd3, 27'h000001c7, 5'd30, 27'h000001cf, 5'd23, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000020, 5'd6, 27'h00000337, 5'd0, 27'h0000002f, 32'h00000400,
  1'd1,  5'd12, 27'h00000004, 5'd9, 27'h00000390, 5'd14, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000028f, 5'd5, 27'h00000372, 5'd21, 27'h00000087, 32'h00000400,
  1'd1,  5'd14, 27'h000001f0, 5'd17, 27'h00000197, 5'd3, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001d1, 5'd16, 27'h000002b6, 5'd10, 27'h000003d2, 32'h00000400,
  1'd1,  5'd15, 27'h00000185, 5'd20, 27'h00000158, 5'd22, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000204, 5'd29, 27'h00000060, 5'd4, 27'h000000c1, 32'h00000400,
  1'd1,  5'd10, 27'h00000322, 5'd27, 27'h0000010c, 5'd14, 27'h0000006c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ed, 5'd30, 27'h000003e4, 5'd21, 27'h000000fe, 32'h00000400,
  1'd1,  5'd24, 27'h0000021e, 5'd8, 27'h0000000e, 5'd4, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003a5, 5'd8, 27'h000000e6, 5'd14, 27'h00000227, 32'h00000400,
  1'd1,  5'd21, 27'h0000020a, 5'd7, 27'h0000029f, 5'd23, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002af, 5'd15, 27'h000002dc, 5'd4, 27'h00000037, 32'h00000400,
  1'd1,  5'd21, 27'h000002fb, 5'd17, 27'h00000162, 5'd12, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003ff, 5'd19, 27'h000003d7, 5'd22, 27'h00000163, 32'h00000400,
  1'd1,  5'd22, 27'h00000165, 5'd27, 27'h000003d3, 5'd1, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000038d, 5'd30, 27'h000003ff, 5'd11, 27'h0000016d, 32'h00000400,
  1'd1,  5'd21, 27'h0000018e, 5'd30, 27'h0000019f, 5'd24, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f3, 5'd10, 27'h000000a7, 5'd5, 27'h00000297, 32'h00000400,
  1'd1,  5'd4, 27'h00000340, 5'd8, 27'h000001ef, 5'd16, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000031f, 5'd6, 27'h000000a2, 5'd30, 27'h000000a3, 32'h00000400,
  1'd1,  5'd2, 27'h0000026b, 5'd17, 27'h00000155, 5'd7, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000134, 5'd17, 27'h0000000d, 5'd16, 27'h0000030f, 32'h00000400,
  1'd1,  5'd0, 27'h0000024b, 5'd18, 27'h000003dc, 5'd30, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000019c, 5'd26, 27'h000002fc, 5'd8, 27'h000002f2, 32'h00000400,
  1'd1,  5'd4, 27'h00000375, 5'd26, 27'h00000250, 5'd18, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000131, 5'd26, 27'h0000034b, 5'd26, 27'h0000015d, 32'h00000400,
  1'd1,  5'd10, 27'h0000022e, 5'd8, 27'h00000322, 5'd6, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000019b, 5'd8, 27'h000001d5, 5'd18, 27'h00000144, 32'h00000400,
  1'd1,  5'd14, 27'h00000361, 5'd7, 27'h0000000e, 5'd27, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c4, 5'd15, 27'h000002cd, 5'd10, 27'h0000001a, 32'h00000400,
  1'd1,  5'd10, 27'h000002a4, 5'd20, 27'h0000001b, 5'd20, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f4, 5'd20, 27'h00000083, 5'd30, 27'h00000294, 32'h00000400,
  1'd1,  5'd13, 27'h00000292, 5'd27, 27'h000001ef, 5'd6, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000158, 5'd29, 27'h00000031, 5'd16, 27'h000001e1, 32'h00000400,
  1'd1,  5'd14, 27'h00000096, 5'd27, 27'h00000366, 5'd28, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002d5, 5'd9, 27'h000000d5, 5'd5, 27'h0000025e, 32'h00000400,
  1'd1,  5'd23, 27'h00000091, 5'd10, 27'h000000fc, 5'd18, 27'h00000001, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002c2, 5'd7, 27'h000002dd, 5'd28, 27'h0000031a, 32'h00000400,
  1'd1,  5'd20, 27'h000002cf, 5'd18, 27'h0000023f, 5'd8, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003db, 5'd18, 27'h00000342, 5'd19, 27'h00000170, 32'h00000400,
  1'd1,  5'd23, 27'h000000f3, 5'd16, 27'h00000272, 5'd28, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003fe, 5'd30, 27'h000002a3, 5'd7, 27'h00000076, 32'h00000400,
  1'd1,  5'd24, 27'h000000ac, 5'd26, 27'h0000004f, 5'd15, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000102, 5'd25, 27'h000003da, 5'd30, 27'h0000036a, 32'h00000400,
  1'd1,  5'd7, 27'h000002a5, 5'd1, 27'h000002bc, 5'd5, 27'h00000222, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d7, 5'd3, 27'h000003bf, 5'd15, 27'h00000273, 32'h00000400,
  1'd1,  5'd6, 27'h000002f4, 5'd2, 27'h00000097, 5'd29, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003d1, 5'd13, 27'h000000b5, 5'd0, 27'h00000071, 32'h00000400,
  1'd1,  5'd6, 27'h00000008, 5'd12, 27'h00000398, 5'd10, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023a, 5'd10, 27'h000002e4, 5'd22, 27'h0000006c, 32'h00000400,
  1'd1,  5'd7, 27'h00000213, 5'd24, 27'h000003a3, 5'd0, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b7, 5'd24, 27'h00000371, 5'd12, 27'h0000027d, 32'h00000400,
  1'd1,  5'd6, 27'h000000fa, 5'd23, 27'h00000195, 5'd22, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000093, 5'd2, 27'h00000183, 5'd6, 27'h000001d9, 32'h00000400,
  1'd1,  5'd18, 27'h00000004, 5'd3, 27'h00000084, 5'd16, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ad, 5'd4, 27'h00000048, 5'd29, 27'h00000299, 32'h00000400,
  1'd1,  5'd16, 27'h000003ea, 5'd12, 27'h00000372, 5'd3, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030c, 5'd10, 27'h00000386, 5'd14, 27'h00000127, 32'h00000400,
  1'd1,  5'd19, 27'h00000024, 5'd11, 27'h00000256, 5'd21, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000357, 5'd20, 27'h000002d4, 5'd3, 27'h00000225, 32'h00000400,
  1'd1,  5'd16, 27'h00000166, 5'd21, 27'h000002a9, 5'd15, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000222, 5'd25, 27'h00000135, 5'd25, 27'h00000130, 32'h00000400,
  1'd1,  5'd30, 27'h000000ac, 5'd0, 27'h000001c3, 5'd0, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000de, 5'd2, 27'h000000cd, 5'd13, 27'h0000008a, 32'h00000400,
  1'd1,  5'd30, 27'h00000120, 5'd4, 27'h0000039c, 5'd21, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000264, 5'd12, 27'h00000173, 5'd2, 27'h000001fa, 32'h00000400,
  1'd1,  5'd28, 27'h000003dc, 5'd13, 27'h0000027b, 5'd15, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000002d, 5'd11, 27'h00000346, 5'd22, 27'h000002f9, 32'h00000400,
  1'd1,  5'd30, 27'h0000030f, 5'd22, 27'h00000322, 5'd4, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000b7, 5'd24, 27'h0000028d, 5'd12, 27'h00000394, 32'h00000400,
  1'd1,  5'd26, 27'h00000367, 5'd23, 27'h0000006a, 5'd23, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000199, 5'd2, 27'h00000231, 5'd3, 27'h000003e2, 32'h00000400,
  1'd1,  5'd5, 27'h000000ff, 5'd4, 27'h00000276, 5'd11, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c3, 5'd4, 27'h00000213, 5'd22, 27'h00000225, 32'h00000400,
  1'd1,  5'd7, 27'h000003b7, 5'd11, 27'h0000007c, 5'd5, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c6, 5'd14, 27'h000003bb, 5'd18, 27'h000002c3, 32'h00000400,
  1'd1,  5'd7, 27'h00000225, 5'd11, 27'h0000038f, 5'd28, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003b3, 5'd22, 27'h0000024b, 5'd7, 27'h000003f2, 32'h00000400,
  1'd1,  5'd6, 27'h00000140, 5'd25, 27'h000001de, 5'd15, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000275, 5'd23, 27'h00000038, 5'd30, 27'h0000020a, 32'h00000400,
  1'd1,  5'd17, 27'h000001a7, 5'd0, 27'h00000083, 5'd3, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000105, 5'd4, 27'h00000045, 5'd13, 27'h00000226, 32'h00000400,
  1'd1,  5'd16, 27'h0000002a, 5'd0, 27'h0000021b, 5'd20, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000396, 5'd11, 27'h000002b4, 5'd7, 27'h00000362, 32'h00000400,
  1'd1,  5'd15, 27'h00000263, 5'd10, 27'h00000358, 5'd16, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000014b, 5'd14, 27'h00000023, 5'd28, 27'h00000323, 32'h00000400,
  1'd1,  5'd16, 27'h0000024f, 5'd23, 27'h000000bc, 5'd9, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003da, 5'd25, 27'h0000008e, 5'd16, 27'h000001ef, 32'h00000400,
  1'd1,  5'd20, 27'h00000196, 5'd20, 27'h000003ae, 5'd27, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000050, 5'd2, 27'h000000de, 5'd6, 27'h0000012b, 32'h00000400,
  1'd1,  5'd28, 27'h00000206, 5'd4, 27'h000002d5, 5'd17, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000022a, 5'd5, 27'h00000013, 5'd28, 27'h00000382, 32'h00000400,
  1'd1,  5'd30, 27'h00000325, 5'd14, 27'h00000356, 5'd7, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000249, 5'd15, 27'h000001bd, 5'd19, 27'h00000330, 32'h00000400,
  1'd1,  5'd29, 27'h000000d3, 5'd14, 27'h0000014b, 5'd29, 27'h00000126, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000020e, 5'd21, 27'h000002cf, 5'd9, 27'h000001b3, 32'h00000400,
  1'd1,  5'd28, 27'h00000258, 5'd21, 27'h0000022b, 5'd18, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000191, 5'd24, 27'h0000007b, 5'd29, 27'h00000337, 32'h00000400,
  1'd1,  5'd10, 27'h00000008, 5'd7, 27'h0000021c, 5'd3, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000238, 5'd6, 27'h00000135, 5'd11, 27'h000002a3, 32'h00000400,
  1'd1,  5'd7, 27'h000001d3, 5'd5, 27'h000001fe, 5'd23, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ac, 5'd17, 27'h00000135, 5'd0, 27'h000002c9, 32'h00000400,
  1'd1,  5'd8, 27'h000001b0, 5'd17, 27'h0000032b, 5'd12, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000127, 5'd17, 27'h00000285, 5'd22, 27'h0000015b, 32'h00000400,
  1'd1,  5'd6, 27'h00000157, 5'd30, 27'h000000c0, 5'd3, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000169, 5'd27, 27'h00000241, 5'd14, 27'h000001af, 32'h00000400,
  1'd1,  5'd8, 27'h000003e5, 5'd28, 27'h0000001c, 5'd21, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000301, 5'd7, 27'h00000057, 5'd0, 27'h000003b6, 32'h00000400,
  1'd1,  5'd18, 27'h0000009c, 5'd9, 27'h00000195, 5'd13, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000033e, 5'd9, 27'h000003b0, 5'd24, 27'h000000aa, 32'h00000400,
  1'd1,  5'd17, 27'h00000027, 5'd19, 27'h000003ee, 5'd0, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000089, 5'd19, 27'h0000011b, 5'd14, 27'h00000308, 32'h00000400,
  1'd1,  5'd17, 27'h00000071, 5'd20, 27'h000000eb, 5'd23, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c1, 5'd28, 27'h00000230, 5'd2, 27'h000001d3, 32'h00000400,
  1'd1,  5'd19, 27'h00000196, 5'd26, 27'h00000168, 5'd15, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000232, 5'd29, 27'h00000150, 5'd25, 27'h00000288, 32'h00000400,
  1'd1,  5'd26, 27'h0000017e, 5'd6, 27'h000000fe, 5'd2, 27'h00000115, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000165, 5'd7, 27'h00000276, 5'd12, 27'h0000033d, 32'h00000400,
  1'd1,  5'd27, 27'h00000354, 5'd6, 27'h0000019b, 5'd25, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000bb, 5'd18, 27'h0000006b, 5'd5, 27'h0000004d, 32'h00000400,
  1'd1,  5'd27, 27'h000003ce, 5'd18, 27'h00000193, 5'd10, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034a, 5'd19, 27'h000001a2, 5'd21, 27'h00000156, 32'h00000400,
  1'd1,  5'd28, 27'h000003c0, 5'd28, 27'h000002c3, 5'd4, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001aa, 5'd27, 27'h000002a7, 5'd15, 27'h0000019c, 32'h00000400,
  1'd1,  5'd28, 27'h0000029d, 5'd27, 27'h00000364, 5'd24, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003bb, 5'd9, 27'h000001eb, 5'd7, 27'h0000016b, 32'h00000400,
  1'd1,  5'd8, 27'h0000023c, 5'd5, 27'h0000026e, 5'd16, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000eb, 5'd9, 27'h00000156, 5'd29, 27'h00000363, 32'h00000400,
  1'd1,  5'd6, 27'h000000e5, 5'd20, 27'h000001f4, 5'd8, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000015e, 5'd19, 27'h00000237, 5'd16, 27'h00000347, 32'h00000400,
  1'd1,  5'd7, 27'h00000391, 5'd15, 27'h00000377, 5'd28, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000007b, 5'd28, 27'h00000217, 5'd5, 27'h000001e3, 32'h00000400,
  1'd1,  5'd7, 27'h000001f3, 5'd27, 27'h0000006a, 5'd17, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000135, 5'd29, 27'h0000016f, 5'd28, 27'h000001d5, 32'h00000400,
  1'd1,  5'd15, 27'h00000274, 5'd9, 27'h00000206, 5'd7, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000031c, 5'd6, 27'h000000ea, 5'd17, 27'h00000031, 32'h00000400,
  1'd1,  5'd18, 27'h00000294, 5'd7, 27'h0000003a, 5'd29, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000174, 5'd19, 27'h00000128, 5'd6, 27'h000001f8, 32'h00000400,
  1'd1,  5'd18, 27'h000000b9, 5'd18, 27'h00000039, 5'd15, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c4, 5'd16, 27'h00000000, 5'd27, 27'h00000369, 32'h00000400,
  1'd1,  5'd20, 27'h00000136, 5'd30, 27'h000003a5, 5'd7, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002b4, 5'd25, 27'h000003a8, 5'd20, 27'h000001f5, 32'h00000400,
  1'd1,  5'd16, 27'h00000006, 5'd29, 27'h000001e0, 5'd28, 27'h000000eb, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d1, 5'd5, 27'h00000178, 5'd6, 27'h00000022, 32'h00000400,
  1'd1,  5'd28, 27'h000002bb, 5'd7, 27'h000001a8, 5'd18, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000a5, 5'd8, 27'h000003ad, 5'd28, 27'h00000304, 32'h00000400,
  1'd1,  5'd30, 27'h00000075, 5'd16, 27'h000003eb, 5'd8, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001f6, 5'd18, 27'h00000095, 5'd20, 27'h00000262, 32'h00000400,
  1'd1,  5'd28, 27'h000003fe, 5'd16, 27'h00000195, 5'd29, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000039d, 5'd29, 27'h000001dd, 5'd5, 27'h0000031c, 32'h00000400,
  1'd1,  5'd26, 27'h0000022a, 5'd30, 27'h00000087, 5'd19, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000136, 5'd28, 27'h000002ed, 5'd27, 27'h000001a3, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000150, 5'd3, 27'h00000167, 5'd0, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000009a, 5'd1, 27'h0000023a, 5'd10, 27'h0000015b, 32'h00000400,
  1'd1,  5'd2, 27'h00000018, 5'd4, 27'h00000306, 5'd21, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000031c, 5'd14, 27'h000003a0, 5'd0, 27'h000003e1, 32'h00000400,
  1'd1,  5'd1, 27'h0000034a, 5'd14, 27'h00000248, 5'd11, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000f4, 5'd12, 27'h00000075, 5'd20, 27'h00000368, 32'h00000400,
  1'd1,  5'd4, 27'h0000007b, 5'd24, 27'h000002cb, 5'd4, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003b8, 5'd20, 27'h00000395, 5'd13, 27'h00000373, 32'h00000400,
  1'd1,  5'd0, 27'h0000023e, 5'd23, 27'h00000119, 5'd23, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000037c, 5'd0, 27'h0000024a, 5'd1, 27'h00000039, 32'h00000400,
  1'd1,  5'd10, 27'h000001b0, 5'd2, 27'h0000015f, 5'd10, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f8, 5'd4, 27'h00000325, 5'd21, 27'h000001a8, 32'h00000400,
  1'd1,  5'd12, 27'h0000033d, 5'd13, 27'h0000019e, 5'd0, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003b9, 5'd14, 27'h00000244, 5'd15, 27'h000000af, 32'h00000400,
  1'd1,  5'd15, 27'h00000093, 5'd11, 27'h00000224, 5'd23, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009d, 5'd22, 27'h0000015f, 5'd1, 27'h0000019f, 32'h00000400,
  1'd1,  5'd13, 27'h0000016d, 5'd24, 27'h0000028f, 5'd12, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f3, 5'd21, 27'h000002f1, 5'd23, 27'h000002f7, 32'h00000400,
  1'd1,  5'd25, 27'h00000309, 5'd0, 27'h00000129, 5'd1, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022c, 5'd2, 27'h0000032d, 5'd11, 27'h00000012, 32'h00000400,
  1'd1,  5'd24, 27'h00000168, 5'd2, 27'h0000038f, 5'd22, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000011c, 5'd14, 27'h00000134, 5'd3, 27'h0000020c, 32'h00000400,
  1'd1,  5'd21, 27'h0000013c, 5'd12, 27'h00000237, 5'd11, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035e, 5'd10, 27'h000001c2, 5'd23, 27'h00000045, 32'h00000400,
  1'd1,  5'd20, 27'h000002ec, 5'd21, 27'h00000275, 5'd5, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000128, 5'd25, 27'h00000263, 5'd15, 27'h00000196, 32'h00000400,
  1'd1,  5'd24, 27'h00000302, 5'd23, 27'h00000122, 5'd24, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000007f, 5'd1, 27'h00000231, 5'd8, 27'h000001ca, 32'h00000400,
  1'd1,  5'd1, 27'h0000008e, 5'd0, 27'h0000022b, 5'd19, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001cd, 5'd3, 27'h00000141, 5'd28, 27'h00000217, 32'h00000400,
  1'd1,  5'd0, 27'h0000023c, 5'd11, 27'h0000034b, 5'd9, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000126, 5'd15, 27'h000000d1, 5'd15, 27'h0000031f, 32'h00000400,
  1'd1,  5'd2, 27'h0000031c, 5'd11, 27'h0000033d, 5'd26, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000211, 5'd25, 27'h00000314, 5'd7, 27'h00000045, 32'h00000400,
  1'd1,  5'd1, 27'h00000348, 5'd24, 27'h00000202, 5'd17, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000314, 5'd25, 27'h00000227, 5'd26, 27'h00000097, 32'h00000400,
  1'd1,  5'd12, 27'h000003de, 5'd0, 27'h0000018f, 5'd9, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000017c, 5'd2, 27'h00000308, 5'd18, 27'h000003b1, 32'h00000400,
  1'd1,  5'd12, 27'h00000325, 5'd1, 27'h00000249, 5'd28, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000121, 5'd13, 27'h0000002c, 5'd9, 27'h000000c7, 32'h00000400,
  1'd1,  5'd10, 27'h00000243, 5'd14, 27'h0000033e, 5'd17, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000382, 5'd11, 27'h00000369, 5'd29, 27'h000001d0, 32'h00000400,
  1'd1,  5'd13, 27'h00000218, 5'd22, 27'h00000268, 5'd7, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d5, 5'd22, 27'h000002d0, 5'd17, 27'h0000027c, 32'h00000400,
  1'd1,  5'd12, 27'h000001c9, 5'd21, 27'h000000d8, 5'd30, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002da, 5'd3, 27'h00000352, 5'd7, 27'h00000312, 32'h00000400,
  1'd1,  5'd22, 27'h00000380, 5'd1, 27'h000002fa, 5'd20, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000140, 5'd4, 27'h00000227, 5'd26, 27'h0000004e, 32'h00000400,
  1'd1,  5'd22, 27'h000003c3, 5'd11, 27'h0000006a, 5'd8, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000163, 5'd14, 27'h0000014c, 5'd18, 27'h000000bc, 32'h00000400,
  1'd1,  5'd25, 27'h0000006c, 5'd10, 27'h00000378, 5'd27, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002a9, 5'd23, 27'h00000110, 5'd10, 27'h000000eb, 32'h00000400,
  1'd1,  5'd21, 27'h00000085, 5'd24, 27'h00000317, 5'd18, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000350, 5'd23, 27'h000003fc, 5'd28, 27'h000001be, 32'h00000400,
  1'd1,  5'd0, 27'h00000015, 5'd9, 27'h000002eb, 5'd4, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000386, 5'd7, 27'h000000c6, 5'd13, 27'h000000e4, 32'h00000400,
  1'd1,  5'd0, 27'h000003f9, 5'd6, 27'h00000243, 5'd24, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000e9, 5'd18, 27'h00000160, 5'd0, 27'h00000298, 32'h00000400,
  1'd1,  5'd4, 27'h000002f0, 5'd19, 27'h000002c9, 5'd13, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000096, 5'd16, 27'h000001b5, 5'd23, 27'h0000039a, 32'h00000400,
  1'd1,  5'd4, 27'h00000064, 5'd30, 27'h00000158, 5'd0, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000028f, 5'd27, 27'h0000028d, 5'd14, 27'h0000012a, 32'h00000400,
  1'd1,  5'd1, 27'h00000295, 5'd27, 27'h000002ac, 5'd24, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000146, 5'd7, 27'h0000019f, 5'd0, 27'h0000016e, 32'h00000400,
  1'd1,  5'd10, 27'h00000386, 5'd7, 27'h000001f6, 5'd12, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f6, 5'd5, 27'h00000306, 5'd24, 27'h000001ba, 32'h00000400,
  1'd1,  5'd11, 27'h00000292, 5'd20, 27'h00000285, 5'd4, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000035e, 5'd15, 27'h00000346, 5'd11, 27'h00000324, 32'h00000400,
  1'd1,  5'd11, 27'h00000284, 5'd16, 27'h0000023b, 5'd22, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001f0, 5'd27, 27'h000001ff, 5'd3, 27'h000000aa, 32'h00000400,
  1'd1,  5'd13, 27'h00000027, 5'd27, 27'h000002a5, 5'd12, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000133, 5'd26, 27'h000000c8, 5'd24, 27'h000000b0, 32'h00000400,
  1'd1,  5'd23, 27'h000003b7, 5'd6, 27'h00000271, 5'd2, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000387, 5'd9, 27'h0000003f, 5'd13, 27'h00000123, 32'h00000400,
  1'd1,  5'd25, 27'h00000232, 5'd6, 27'h000001e3, 5'd21, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000008c, 5'd17, 27'h000000ec, 5'd0, 27'h000001f0, 32'h00000400,
  1'd1,  5'd21, 27'h000001e4, 5'd19, 27'h00000154, 5'd11, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000186, 5'd16, 27'h000003c1, 5'd24, 27'h000003f8, 32'h00000400,
  1'd1,  5'd22, 27'h000002cc, 5'd29, 27'h00000304, 5'd0, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000eb, 5'd30, 27'h000003e8, 5'd14, 27'h00000300, 32'h00000400,
  1'd1,  5'd23, 27'h00000281, 5'd30, 27'h0000003d, 5'd22, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b1, 5'd6, 27'h0000004d, 5'd7, 27'h0000009c, 32'h00000400,
  1'd1,  5'd0, 27'h000000b9, 5'd8, 27'h0000009b, 5'd15, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001bb, 5'd8, 27'h000002d5, 5'd28, 27'h0000011d, 32'h00000400,
  1'd1,  5'd2, 27'h00000191, 5'd17, 27'h00000136, 5'd7, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000001, 5'd15, 27'h00000222, 5'd16, 27'h0000006a, 32'h00000400,
  1'd1,  5'd2, 27'h000000e8, 5'd19, 27'h00000207, 5'd28, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f6, 5'd27, 27'h0000008e, 5'd9, 27'h00000011, 32'h00000400,
  1'd1,  5'd4, 27'h00000035, 5'd26, 27'h000003a2, 5'd18, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000d4, 5'd27, 27'h00000138, 5'd30, 27'h000003ed, 32'h00000400,
  1'd1,  5'd10, 27'h00000190, 5'd7, 27'h000000e1, 5'd6, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023d, 5'd8, 27'h00000199, 5'd19, 27'h0000000c, 32'h00000400,
  1'd1,  5'd10, 27'h0000016f, 5'd6, 27'h000003f9, 5'd28, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000195, 5'd15, 27'h000003e1, 5'd10, 27'h00000095, 32'h00000400,
  1'd1,  5'd12, 27'h00000237, 5'd16, 27'h00000028, 5'd17, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c3, 5'd20, 27'h00000064, 5'd28, 27'h0000001e, 32'h00000400,
  1'd1,  5'd11, 27'h000002d0, 5'd29, 27'h0000017a, 5'd6, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000034a, 5'd30, 27'h00000178, 5'd18, 27'h000000a0, 32'h00000400,
  1'd1,  5'd11, 27'h000002c6, 5'd27, 27'h00000378, 5'd28, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001ed, 5'd9, 27'h00000214, 5'd5, 27'h000003fe, 32'h00000400,
  1'd1,  5'd21, 27'h00000190, 5'd5, 27'h0000034b, 5'd17, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000268, 5'd7, 27'h00000205, 5'd27, 27'h0000012c, 32'h00000400,
  1'd1,  5'd24, 27'h00000076, 5'd17, 27'h000003e8, 5'd5, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000013c, 5'd19, 27'h00000007, 5'd20, 27'h000000b1, 32'h00000400,
  1'd1,  5'd24, 27'h0000035b, 5'd18, 27'h000003f3, 5'd29, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d5, 5'd27, 27'h00000256, 5'd5, 27'h000003cd, 32'h00000400,
  1'd1,  5'd22, 27'h0000034a, 5'd30, 27'h00000382, 5'd20, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003aa, 5'd27, 27'h000001c2, 5'd28, 27'h000002d1, 32'h00000400,
  1'd1,  5'd6, 27'h00000287, 5'd2, 27'h00000247, 5'd5, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000368, 5'd3, 27'h00000157, 5'd20, 27'h00000040, 32'h00000400,
  1'd1,  5'd9, 27'h00000282, 5'd4, 27'h00000356, 5'd27, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000215, 5'd15, 27'h000001ff, 5'd1, 27'h000000f2, 32'h00000400,
  1'd1,  5'd5, 27'h000000b2, 5'd11, 27'h000002ee, 5'd12, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001f8, 5'd11, 27'h0000023c, 5'd23, 27'h0000017a, 32'h00000400,
  1'd1,  5'd5, 27'h000000d1, 5'd24, 27'h00000126, 5'd1, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000027, 5'd20, 27'h0000039f, 5'd11, 27'h00000284, 32'h00000400,
  1'd1,  5'd9, 27'h000001ef, 5'd23, 27'h000000f8, 5'd20, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000234, 5'd2, 27'h00000385, 5'd9, 27'h0000021b, 32'h00000400,
  1'd1,  5'd17, 27'h000002bb, 5'd2, 27'h00000147, 5'd16, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001f8, 5'd3, 27'h000002ec, 5'd27, 27'h000001bf, 32'h00000400,
  1'd1,  5'd18, 27'h00000308, 5'd12, 27'h0000011e, 5'd0, 27'h000001b5, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002dc, 5'd13, 27'h0000007b, 5'd11, 27'h000001c1, 32'h00000400,
  1'd1,  5'd17, 27'h000001ac, 5'd11, 27'h00000130, 5'd24, 27'h000003d8, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000381, 5'd23, 27'h00000238, 5'd4, 27'h00000039, 32'h00000400,
  1'd1,  5'd16, 27'h00000178, 5'd22, 27'h00000342, 5'd11, 27'h0000006d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000068, 5'd24, 27'h0000027f, 5'd24, 27'h0000003d, 32'h00000400,
  1'd1,  5'd29, 27'h00000394, 5'd4, 27'h0000013a, 5'd0, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000287, 5'd4, 27'h000001b5, 5'd13, 27'h000000d5, 32'h00000400,
  1'd1,  5'd28, 27'h00000212, 5'd3, 27'h00000076, 5'd24, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b3, 5'd13, 27'h000001ec, 5'd3, 27'h0000022a, 32'h00000400,
  1'd1,  5'd28, 27'h00000108, 5'd11, 27'h0000008c, 5'd13, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b6, 5'd12, 27'h000002bc, 5'd22, 27'h000001d4, 32'h00000400,
  1'd1,  5'd29, 27'h000003c7, 5'd20, 27'h000003ec, 5'd1, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001e4, 5'd25, 27'h000002f0, 5'd15, 27'h00000128, 32'h00000400,
  1'd1,  5'd28, 27'h0000000b, 5'd22, 27'h00000389, 5'd21, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000361, 5'd3, 27'h00000386, 5'd2, 27'h000003a5, 32'h00000400,
  1'd1,  5'd9, 27'h0000005f, 5'd1, 27'h00000205, 5'd14, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000fe, 5'd0, 27'h00000373, 5'd22, 27'h00000185, 32'h00000400,
  1'd1,  5'd7, 27'h00000090, 5'd11, 27'h000002cd, 5'd8, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000007a, 5'd11, 27'h0000022b, 5'd19, 27'h000000ba, 32'h00000400,
  1'd1,  5'd8, 27'h000001c4, 5'd14, 27'h000003b6, 5'd26, 27'h000001be, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e2, 5'd23, 27'h0000015d, 5'd9, 27'h0000012e, 32'h00000400,
  1'd1,  5'd9, 27'h0000015a, 5'd22, 27'h000000e6, 5'd15, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000383, 5'd21, 27'h00000116, 5'd28, 27'h00000277, 32'h00000400,
  1'd1,  5'd15, 27'h000003b2, 5'd3, 27'h00000057, 5'd4, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e6, 5'd4, 27'h000001e2, 5'd13, 27'h00000285, 32'h00000400,
  1'd1,  5'd19, 27'h0000012c, 5'd1, 27'h000003ce, 5'd24, 27'h000000e3, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000202, 5'd11, 27'h000000e2, 5'd5, 27'h00000181, 32'h00000400,
  1'd1,  5'd17, 27'h00000283, 5'd14, 27'h0000020c, 5'd18, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000177, 5'd13, 27'h000000f4, 5'd26, 27'h00000111, 32'h00000400,
  1'd1,  5'd16, 27'h00000074, 5'd21, 27'h0000030c, 5'd7, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000172, 5'd20, 27'h000002e2, 5'd20, 27'h00000021, 32'h00000400,
  1'd1,  5'd20, 27'h00000294, 5'd25, 27'h000001e1, 5'd27, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000d8, 5'd3, 27'h000000d0, 5'd9, 27'h000000a4, 32'h00000400,
  1'd1,  5'd27, 27'h000002bc, 5'd1, 27'h0000026f, 5'd20, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000364, 5'd3, 27'h00000194, 5'd26, 27'h000003e0, 32'h00000400,
  1'd1,  5'd30, 27'h000002f0, 5'd15, 27'h00000179, 5'd8, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001cf, 5'd10, 27'h000001be, 5'd19, 27'h00000386, 32'h00000400,
  1'd1,  5'd27, 27'h0000018d, 5'd12, 27'h000002bd, 5'd28, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003ab, 5'd23, 27'h0000024c, 5'd7, 27'h000001e1, 32'h00000400,
  1'd1,  5'd29, 27'h000003a8, 5'd20, 27'h000003fd, 5'd18, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000056, 5'd24, 27'h0000001b, 5'd30, 27'h000002f2, 32'h00000400,
  1'd1,  5'd7, 27'h000003dd, 5'd7, 27'h00000150, 5'd3, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000102, 5'd7, 27'h000003b8, 5'd12, 27'h00000313, 32'h00000400,
  1'd1,  5'd9, 27'h00000298, 5'd8, 27'h00000248, 5'd25, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002ba, 5'd18, 27'h0000012c, 5'd1, 27'h00000178, 32'h00000400,
  1'd1,  5'd6, 27'h000000e4, 5'd17, 27'h00000169, 5'd13, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e5, 5'd19, 27'h000002de, 5'd22, 27'h00000379, 32'h00000400,
  1'd1,  5'd10, 27'h000000ba, 5'd27, 27'h000000ea, 5'd3, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000214, 5'd26, 27'h0000011c, 5'd11, 27'h000001df, 32'h00000400,
  1'd1,  5'd10, 27'h0000006b, 5'd27, 27'h00000047, 5'd22, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b3, 5'd7, 27'h0000012d, 5'd3, 27'h00000127, 32'h00000400,
  1'd1,  5'd17, 27'h000003fc, 5'd5, 27'h00000137, 5'd12, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001e1, 5'd5, 27'h000001c1, 5'd25, 27'h0000023d, 32'h00000400,
  1'd1,  5'd15, 27'h00000215, 5'd15, 27'h000003bf, 5'd0, 27'h000003a6, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000015e, 5'd17, 27'h00000188, 5'd14, 27'h00000119, 32'h00000400,
  1'd1,  5'd15, 27'h000003e2, 5'd17, 27'h000002e7, 5'd22, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000db, 5'd30, 27'h0000025e, 5'd1, 27'h00000182, 32'h00000400,
  1'd1,  5'd18, 27'h0000024b, 5'd29, 27'h0000038c, 5'd12, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e2, 5'd26, 27'h0000033c, 5'd22, 27'h000001a8, 32'h00000400,
  1'd1,  5'd26, 27'h000000b4, 5'd7, 27'h00000075, 5'd3, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038a, 5'd7, 27'h0000031f, 5'd12, 27'h0000017f, 32'h00000400,
  1'd1,  5'd27, 27'h000003d6, 5'd8, 27'h000002e2, 5'd23, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000195, 5'd18, 27'h000001cf, 5'd5, 27'h00000031, 32'h00000400,
  1'd1,  5'd28, 27'h000002ae, 5'd18, 27'h00000168, 5'd11, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000029f, 5'd18, 27'h000000c8, 5'd22, 27'h000003ed, 32'h00000400,
  1'd1,  5'd30, 27'h0000030b, 5'd30, 27'h00000038, 5'd4, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a0, 5'd26, 27'h00000034, 5'd12, 27'h000002ef, 32'h00000400,
  1'd1,  5'd28, 27'h000000a2, 5'd25, 27'h000003d6, 5'd23, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000323, 5'd10, 27'h00000125, 5'd9, 27'h0000026e, 32'h00000400,
  1'd1,  5'd8, 27'h0000034d, 5'd9, 27'h000003ca, 5'd16, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000064, 5'd8, 27'h0000021d, 5'd28, 27'h0000021c, 32'h00000400,
  1'd1,  5'd9, 27'h0000006e, 5'd15, 27'h000002e9, 5'd5, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000164, 5'd20, 27'h000000b8, 5'd17, 27'h0000020b, 32'h00000400,
  1'd1,  5'd5, 27'h00000130, 5'd19, 27'h000000ba, 5'd25, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ca, 5'd26, 27'h000000fb, 5'd6, 27'h00000004, 32'h00000400,
  1'd1,  5'd9, 27'h00000091, 5'd27, 27'h00000052, 5'd20, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002c8, 5'd27, 27'h0000012e, 5'd28, 27'h000000fa, 32'h00000400,
  1'd1,  5'd19, 27'h00000127, 5'd7, 27'h000003a2, 5'd6, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000354, 5'd5, 27'h00000196, 5'd18, 27'h00000209, 32'h00000400,
  1'd1,  5'd17, 27'h000000e8, 5'd7, 27'h00000387, 5'd27, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002e0, 5'd16, 27'h000001d4, 5'd9, 27'h00000262, 32'h00000400,
  1'd1,  5'd19, 27'h0000034d, 5'd17, 27'h00000030, 5'd15, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000029b, 5'd15, 27'h000002eb, 5'd29, 27'h000002e7, 32'h00000400,
  1'd1,  5'd20, 27'h00000058, 5'd30, 27'h00000234, 5'd8, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000109, 5'd28, 27'h000000ed, 5'd17, 27'h00000070, 32'h00000400,
  1'd1,  5'd19, 27'h000003d8, 5'd26, 27'h000001bb, 5'd25, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000230, 5'd6, 27'h0000018b, 5'd6, 27'h000002a4, 32'h00000400,
  1'd1,  5'd27, 27'h0000025f, 5'd7, 27'h000000cc, 5'd18, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000071, 5'd8, 27'h0000006c, 5'd29, 27'h00000028, 32'h00000400,
  1'd1,  5'd29, 27'h00000295, 5'd17, 27'h00000148, 5'd6, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000243, 5'd20, 27'h00000298, 5'd18, 27'h00000360, 32'h00000400,
  1'd1,  5'd27, 27'h00000112, 5'd17, 27'h00000201, 5'd29, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000132, 5'd29, 27'h000003bc, 5'd5, 27'h0000011f, 32'h00000400,
  1'd1,  5'd30, 27'h000002bb, 5'd30, 27'h00000362, 5'd18, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000017b, 5'd26, 27'h00000253, 5'd26, 27'h00000321, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000000d7, 5'd4, 27'h000001a4, 5'd4, 27'h00000103, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003a7, 5'd0, 27'h00000289, 5'd13, 27'h000001aa, 32'h00000400,
  1'd1,  5'd4, 27'h00000300, 5'd2, 27'h0000039a, 5'd22, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ef, 5'd11, 27'h000003af, 5'd0, 27'h0000038b, 32'h00000400,
  1'd1,  5'd2, 27'h00000251, 5'd10, 27'h00000173, 5'd11, 27'h00000076, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002ea, 5'd13, 27'h0000023a, 5'd21, 27'h000000c7, 32'h00000400,
  1'd1,  5'd1, 27'h000003be, 5'd24, 27'h0000027b, 5'd5, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000017f, 5'd24, 27'h000003ce, 5'd10, 27'h00000176, 32'h00000400,
  1'd1,  5'd0, 27'h000001f2, 5'd23, 27'h000002b6, 5'd23, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000022a, 5'd4, 27'h00000146, 5'd3, 27'h00000252, 32'h00000400,
  1'd1,  5'd13, 27'h0000002c, 5'd1, 27'h000003b8, 5'd11, 27'h000003e1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000b4, 5'd4, 27'h00000218, 5'd24, 27'h0000014a, 32'h00000400,
  1'd1,  5'd15, 27'h000000d4, 5'd13, 27'h00000320, 5'd3, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001b4, 5'd14, 27'h000001bf, 5'd12, 27'h00000238, 32'h00000400,
  1'd1,  5'd11, 27'h000000e9, 5'd11, 27'h000003ba, 5'd21, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000125, 5'd25, 27'h0000028b, 5'd2, 27'h00000067, 32'h00000400,
  1'd1,  5'd11, 27'h00000119, 5'd21, 27'h00000322, 5'd15, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000063, 5'd24, 27'h0000002d, 5'd20, 27'h000003de, 32'h00000400,
  1'd1,  5'd25, 27'h0000004c, 5'd1, 27'h00000173, 5'd4, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003b3, 5'd0, 27'h00000348, 5'd11, 27'h00000193, 32'h00000400,
  1'd1,  5'd22, 27'h00000354, 5'd2, 27'h0000020d, 5'd22, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000162, 5'd11, 27'h00000068, 5'd3, 27'h0000022f, 32'h00000400,
  1'd1,  5'd24, 27'h000000a1, 5'd12, 27'h00000314, 5'd12, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001e1, 5'd13, 27'h000002e1, 5'd21, 27'h0000039b, 32'h00000400,
  1'd1,  5'd21, 27'h000003b0, 5'd24, 27'h000001e5, 5'd2, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000032f, 5'd23, 27'h00000025, 5'd14, 27'h000002d9, 32'h00000400,
  1'd1,  5'd20, 27'h000003f0, 5'd25, 27'h0000003e, 5'd20, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000268, 5'd1, 27'h000002ab, 5'd8, 27'h000001e7, 32'h00000400,
  1'd1,  5'd4, 27'h0000037d, 5'd0, 27'h0000018f, 5'd16, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002c0, 5'd0, 27'h000002cf, 5'd26, 27'h0000030f, 32'h00000400,
  1'd1,  5'd2, 27'h000000db, 5'd14, 27'h000002b4, 5'd5, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000016b, 5'd11, 27'h000000d0, 5'd19, 27'h000000b3, 32'h00000400,
  1'd1,  5'd2, 27'h00000120, 5'd14, 27'h000003d7, 5'd28, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000008, 5'd24, 27'h0000000b, 5'd6, 27'h00000037, 32'h00000400,
  1'd1,  5'd2, 27'h000003f5, 5'd23, 27'h00000196, 5'd17, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000254, 5'd22, 27'h00000060, 5'd28, 27'h00000320, 32'h00000400,
  1'd1,  5'd14, 27'h0000005b, 5'd3, 27'h00000188, 5'd5, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003f6, 5'd2, 27'h0000037b, 5'd16, 27'h000001e6, 32'h00000400,
  1'd1,  5'd11, 27'h000003af, 5'd1, 27'h00000320, 5'd26, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000145, 5'd10, 27'h000002e5, 5'd5, 27'h00000131, 32'h00000400,
  1'd1,  5'd14, 27'h00000045, 5'd11, 27'h00000355, 5'd17, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000261, 5'd15, 27'h000000e5, 5'd27, 27'h0000027f, 32'h00000400,
  1'd1,  5'd15, 27'h00000065, 5'd23, 27'h00000322, 5'd7, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000335, 5'd22, 27'h0000021c, 5'd19, 27'h000002a5, 32'h00000400,
  1'd1,  5'd11, 27'h000003ed, 5'd23, 27'h000003b2, 5'd25, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000059, 5'd0, 27'h0000037a, 5'd6, 27'h00000334, 32'h00000400,
  1'd1,  5'd22, 27'h000000b8, 5'd3, 27'h00000122, 5'd17, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000381, 5'd4, 27'h000003ed, 5'd28, 27'h000000c2, 32'h00000400,
  1'd1,  5'd24, 27'h000002fd, 5'd15, 27'h00000089, 5'd6, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000221, 5'd11, 27'h00000262, 5'd19, 27'h00000094, 32'h00000400,
  1'd1,  5'd23, 27'h000002f4, 5'd12, 27'h000003ce, 5'd30, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000001e, 5'd22, 27'h000001df, 5'd6, 27'h00000364, 32'h00000400,
  1'd1,  5'd25, 27'h000001b5, 5'd24, 27'h000002fa, 5'd19, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000305, 5'd22, 27'h00000067, 5'd27, 27'h0000001b, 32'h00000400,
  1'd1,  5'd0, 27'h000001e0, 5'd10, 27'h00000101, 5'd4, 27'h000000b0, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e0, 5'd6, 27'h00000081, 5'd10, 27'h0000019e, 32'h00000400,
  1'd1,  5'd0, 27'h0000038a, 5'd8, 27'h000003dc, 5'd22, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000249, 5'd19, 27'h000002af, 5'd3, 27'h000002ab, 32'h00000400,
  1'd1,  5'd3, 27'h0000014f, 5'd17, 27'h00000328, 5'd13, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002db, 5'd19, 27'h00000043, 5'd23, 27'h00000236, 32'h00000400,
  1'd1,  5'd0, 27'h00000188, 5'd27, 27'h00000013, 5'd4, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000057, 5'd26, 27'h00000212, 5'd14, 27'h000000d1, 32'h00000400,
  1'd1,  5'd1, 27'h0000037b, 5'd30, 27'h00000295, 5'd21, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002b6, 5'd9, 27'h00000133, 5'd3, 27'h0000039f, 32'h00000400,
  1'd1,  5'd12, 27'h00000394, 5'd5, 27'h0000015f, 5'd13, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000030b, 5'd8, 27'h000003a0, 5'd22, 27'h0000029c, 32'h00000400,
  1'd1,  5'd12, 27'h00000294, 5'd18, 27'h00000106, 5'd2, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e4, 5'd17, 27'h000003f5, 5'd11, 27'h00000150, 32'h00000400,
  1'd1,  5'd12, 27'h0000022f, 5'd19, 27'h000000e7, 5'd21, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002d4, 5'd29, 27'h000002ca, 5'd3, 27'h000001a6, 32'h00000400,
  1'd1,  5'd12, 27'h000003a0, 5'd27, 27'h0000036d, 5'd12, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000000b, 5'd27, 27'h000000f2, 5'd22, 27'h00000188, 32'h00000400,
  1'd1,  5'd24, 27'h000001a9, 5'd9, 27'h000000e8, 5'd2, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000026, 5'd5, 27'h000000bd, 5'd15, 27'h000000f7, 32'h00000400,
  1'd1,  5'd24, 27'h000003cb, 5'd9, 27'h0000030a, 5'd21, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021c, 5'd18, 27'h0000037f, 5'd1, 27'h000003b5, 32'h00000400,
  1'd1,  5'd23, 27'h000000d0, 5'd15, 27'h00000301, 5'd11, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000116, 5'd17, 27'h0000003e, 5'd21, 27'h00000086, 32'h00000400,
  1'd1,  5'd25, 27'h000001df, 5'd26, 27'h00000376, 5'd3, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000203, 5'd26, 27'h0000037e, 5'd13, 27'h000003b6, 32'h00000400,
  1'd1,  5'd23, 27'h0000011e, 5'd28, 27'h000000ee, 5'd21, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000060, 5'd8, 27'h000000ff, 5'd7, 27'h00000281, 32'h00000400,
  1'd1,  5'd2, 27'h0000029c, 5'd5, 27'h00000211, 5'd17, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000299, 5'd7, 27'h000000d3, 5'd29, 27'h000001c3, 32'h00000400,
  1'd1,  5'd0, 27'h00000153, 5'd18, 27'h0000017b, 5'd6, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003a3, 5'd17, 27'h0000026b, 5'd15, 27'h0000024e, 32'h00000400,
  1'd1,  5'd0, 27'h000001cf, 5'd17, 27'h00000050, 5'd30, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000039c, 5'd27, 27'h00000375, 5'd8, 27'h0000008c, 32'h00000400,
  1'd1,  5'd4, 27'h000001e1, 5'd28, 27'h0000018a, 5'd20, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000051, 5'd29, 27'h0000022a, 5'd26, 27'h000001de, 32'h00000400,
  1'd1,  5'd12, 27'h00000047, 5'd7, 27'h0000029c, 5'd9, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001a7, 5'd7, 27'h00000317, 5'd16, 27'h00000335, 32'h00000400,
  1'd1,  5'd12, 27'h000000b3, 5'd7, 27'h00000269, 5'd30, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000024b, 5'd15, 27'h00000286, 5'd6, 27'h0000008d, 32'h00000400,
  1'd1,  5'd14, 27'h00000043, 5'd19, 27'h000000cf, 5'd17, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ea, 5'd17, 27'h00000029, 5'd27, 27'h00000067, 32'h00000400,
  1'd1,  5'd12, 27'h000002fa, 5'd27, 27'h00000187, 5'd10, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000d0, 5'd28, 27'h00000397, 5'd19, 27'h0000026e, 32'h00000400,
  1'd1,  5'd13, 27'h000003f6, 5'd28, 27'h00000257, 5'd30, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000201, 5'd6, 27'h0000005e, 5'd6, 27'h000000cc, 32'h00000400,
  1'd1,  5'd21, 27'h00000268, 5'd6, 27'h0000005e, 5'd18, 27'h0000012c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000033a, 5'd5, 27'h0000032c, 5'd27, 27'h000002ff, 32'h00000400,
  1'd1,  5'd22, 27'h0000005f, 5'd19, 27'h0000028c, 5'd6, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000197, 5'd16, 27'h0000038d, 5'd15, 27'h000003b9, 32'h00000400,
  1'd1,  5'd21, 27'h00000318, 5'd19, 27'h000001b1, 5'd28, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b7, 5'd26, 27'h000001a0, 5'd8, 27'h00000133, 32'h00000400,
  1'd1,  5'd20, 27'h000002bb, 5'd30, 27'h00000390, 5'd17, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003d1, 5'd26, 27'h00000267, 5'd25, 27'h000003b2, 32'h00000400,
  1'd1,  5'd9, 27'h0000027c, 5'd1, 27'h000001b7, 5'd10, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000250, 5'd3, 27'h000002e6, 5'd18, 27'h00000135, 32'h00000400,
  1'd1,  5'd9, 27'h000003bd, 5'd1, 27'h0000032d, 5'd25, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ae, 5'd13, 27'h0000022f, 5'd2, 27'h00000166, 32'h00000400,
  1'd1,  5'd8, 27'h00000315, 5'd14, 27'h000002a7, 5'd12, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ac, 5'd12, 27'h00000111, 5'd24, 27'h000002b7, 32'h00000400,
  1'd1,  5'd9, 27'h000000f8, 5'd21, 27'h00000183, 5'd1, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000372, 5'd25, 27'h00000301, 5'd12, 27'h0000021c, 32'h00000400,
  1'd1,  5'd10, 27'h00000117, 5'd24, 27'h00000183, 5'd24, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000180, 5'd4, 27'h00000015, 5'd5, 27'h000001d4, 32'h00000400,
  1'd1,  5'd17, 27'h000003c3, 5'd0, 27'h0000025e, 5'd16, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000160, 5'd1, 27'h000000d0, 5'd26, 27'h0000010f, 32'h00000400,
  1'd1,  5'd18, 27'h000001fe, 5'd12, 27'h000001c7, 5'd4, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011d, 5'd14, 27'h000000ba, 5'd14, 27'h00000171, 32'h00000400,
  1'd1,  5'd15, 27'h000002dc, 5'd15, 27'h00000062, 5'd22, 27'h00000234, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000115, 5'd20, 27'h00000318, 5'd2, 27'h000001dd, 32'h00000400,
  1'd1,  5'd15, 27'h00000330, 5'd24, 27'h000003cb, 5'd13, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000e9, 5'd24, 27'h00000083, 5'd21, 27'h00000276, 32'h00000400,
  1'd1,  5'd26, 27'h00000226, 5'd4, 27'h0000015d, 5'd0, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e7, 5'd4, 27'h000002d6, 5'd12, 27'h00000135, 32'h00000400,
  1'd1,  5'd29, 27'h00000028, 5'd4, 27'h000003cb, 5'd24, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000016e, 5'd13, 27'h00000380, 5'd4, 27'h0000038b, 32'h00000400,
  1'd1,  5'd30, 27'h0000004d, 5'd12, 27'h00000112, 5'd13, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000171, 5'd13, 27'h0000017e, 5'd21, 27'h00000076, 32'h00000400,
  1'd1,  5'd27, 27'h0000020b, 5'd25, 27'h000000ef, 5'd1, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a1, 5'd23, 27'h00000215, 5'd15, 27'h00000089, 32'h00000400,
  1'd1,  5'd30, 27'h000003f8, 5'd22, 27'h000000a9, 5'd24, 27'h00000114, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000008, 5'd3, 27'h00000346, 5'd4, 27'h000002c9, 32'h00000400,
  1'd1,  5'd5, 27'h000002a9, 5'd2, 27'h0000030b, 5'd11, 27'h00000119, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000196, 5'd3, 27'h0000015d, 5'd21, 27'h0000027c, 32'h00000400,
  1'd1,  5'd10, 27'h000000e5, 5'd10, 27'h000003eb, 5'd8, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000002, 5'd13, 27'h0000009b, 5'd19, 27'h00000223, 32'h00000400,
  1'd1,  5'd7, 27'h00000038, 5'd11, 27'h00000259, 5'd29, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000381, 5'd23, 27'h000002ac, 5'd8, 27'h0000018a, 32'h00000400,
  1'd1,  5'd7, 27'h000000ea, 5'd24, 27'h00000077, 5'd17, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000280, 5'd21, 27'h00000290, 5'd30, 27'h000000f3, 32'h00000400,
  1'd1,  5'd19, 27'h000000b8, 5'd3, 27'h00000130, 5'd3, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003af, 5'd0, 27'h00000068, 5'd12, 27'h0000034b, 32'h00000400,
  1'd1,  5'd16, 27'h00000333, 5'd3, 27'h0000025c, 5'd25, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000234, 5'd11, 27'h00000359, 5'd9, 27'h000000f3, 32'h00000400,
  1'd1,  5'd18, 27'h0000000a, 5'd14, 27'h0000034c, 5'd16, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003d0, 5'd12, 27'h000001a7, 5'd29, 27'h000001c2, 32'h00000400,
  1'd1,  5'd19, 27'h00000060, 5'd23, 27'h000002d5, 5'd6, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000004, 5'd25, 27'h000001b3, 5'd19, 27'h0000000b, 32'h00000400,
  1'd1,  5'd20, 27'h000000de, 5'd24, 27'h000001fe, 5'd29, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000025d, 5'd0, 27'h0000003c, 5'd5, 27'h00000395, 32'h00000400,
  1'd1,  5'd26, 27'h000000ee, 5'd1, 27'h00000390, 5'd17, 27'h00000082, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000034d, 5'd2, 27'h00000387, 5'd27, 27'h000000d1, 32'h00000400,
  1'd1,  5'd27, 27'h00000094, 5'd11, 27'h00000393, 5'd8, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000022b, 5'd12, 27'h0000011c, 5'd15, 27'h00000386, 32'h00000400,
  1'd1,  5'd26, 27'h0000038b, 5'd11, 27'h000002cb, 5'd29, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000b1, 5'd21, 27'h00000162, 5'd9, 27'h00000362, 32'h00000400,
  1'd1,  5'd29, 27'h000001c8, 5'd24, 27'h000002a9, 5'd17, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003db, 5'd25, 27'h0000021d, 5'd27, 27'h00000048, 32'h00000400,
  1'd1,  5'd9, 27'h0000007e, 5'd6, 27'h000001da, 5'd0, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c6, 5'd6, 27'h00000399, 5'd14, 27'h0000029e, 32'h00000400,
  1'd1,  5'd7, 27'h00000249, 5'd8, 27'h0000012b, 5'd22, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003a6, 5'd16, 27'h00000120, 5'd4, 27'h000003b5, 32'h00000400,
  1'd1,  5'd6, 27'h0000029b, 5'd18, 27'h000002a6, 5'd13, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000169, 5'd17, 27'h0000014d, 5'd24, 27'h000000ce, 32'h00000400,
  1'd1,  5'd8, 27'h00000031, 5'd30, 27'h00000262, 5'd3, 27'h000001f9, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000013a, 5'd27, 27'h00000101, 5'd13, 27'h000002be, 32'h00000400,
  1'd1,  5'd6, 27'h00000034, 5'd27, 27'h000003d9, 5'd22, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000272, 5'd5, 27'h000000e3, 5'd1, 27'h000003e8, 32'h00000400,
  1'd1,  5'd17, 27'h00000392, 5'd9, 27'h00000120, 5'd13, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000035b, 5'd9, 27'h0000004a, 5'd25, 27'h0000031f, 32'h00000400,
  1'd1,  5'd16, 27'h00000215, 5'd20, 27'h000001bd, 5'd0, 27'h00000284, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000308, 5'd16, 27'h0000030c, 5'd10, 27'h00000282, 32'h00000400,
  1'd1,  5'd15, 27'h0000039c, 5'd19, 27'h0000000d, 5'd22, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000037, 5'd27, 27'h00000094, 5'd4, 27'h00000197, 32'h00000400,
  1'd1,  5'd18, 27'h000001cf, 5'd27, 27'h000001c1, 5'd12, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000ac, 5'd26, 27'h000000f8, 5'd22, 27'h000001fc, 32'h00000400,
  1'd1,  5'd28, 27'h00000394, 5'd8, 27'h00000121, 5'd0, 27'h000001b8, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f9, 5'd9, 27'h00000187, 5'd13, 27'h00000110, 32'h00000400,
  1'd1,  5'd27, 27'h00000178, 5'd5, 27'h000000cb, 5'd22, 27'h000000a9, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000378, 5'd19, 27'h00000002, 5'd4, 27'h00000012, 32'h00000400,
  1'd1,  5'd29, 27'h0000027c, 5'd19, 27'h00000161, 5'd13, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000366, 5'd17, 27'h0000037f, 5'd23, 27'h000003a3, 32'h00000400,
  1'd1,  5'd27, 27'h0000025c, 5'd26, 27'h00000094, 5'd1, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036a, 5'd28, 27'h0000031e, 5'd11, 27'h000001c0, 32'h00000400,
  1'd1,  5'd26, 27'h00000345, 5'd27, 27'h00000107, 5'd22, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000273, 5'd8, 27'h00000101, 5'd10, 27'h00000043, 32'h00000400,
  1'd1,  5'd9, 27'h000000b8, 5'd9, 27'h0000016b, 5'd18, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023f, 5'd5, 27'h00000247, 5'd26, 27'h0000006b, 32'h00000400,
  1'd1,  5'd10, 27'h00000095, 5'd17, 27'h000003b5, 5'd7, 27'h000003d6, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000329, 5'd19, 27'h000003d5, 5'd20, 27'h000001af, 32'h00000400,
  1'd1,  5'd6, 27'h00000214, 5'd15, 27'h00000312, 5'd29, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033b, 5'd30, 27'h00000086, 5'd5, 27'h000000c0, 32'h00000400,
  1'd1,  5'd9, 27'h00000332, 5'd28, 27'h00000188, 5'd17, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000028, 5'd27, 27'h000002e8, 5'd26, 27'h000002ee, 32'h00000400,
  1'd1,  5'd19, 27'h00000064, 5'd6, 27'h000001ac, 5'd7, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000004f, 5'd9, 27'h00000028, 5'd18, 27'h000003b2, 32'h00000400,
  1'd1,  5'd17, 27'h0000032c, 5'd8, 27'h00000202, 5'd26, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000036d, 5'd20, 27'h0000012b, 5'd6, 27'h0000019a, 32'h00000400,
  1'd1,  5'd17, 27'h00000391, 5'd17, 27'h0000033b, 5'd17, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002c9, 5'd18, 27'h00000141, 5'd28, 27'h0000038c, 32'h00000400,
  1'd1,  5'd16, 27'h00000365, 5'd30, 27'h000001b1, 5'd5, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000249, 5'd29, 27'h000000c6, 5'd19, 27'h0000017c, 32'h00000400,
  1'd1,  5'd18, 27'h00000219, 5'd28, 27'h000002f0, 5'd30, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000400, 5'd7, 27'h000002ef, 5'd8, 27'h00000197, 32'h00000400,
  1'd1,  5'd28, 27'h00000023, 5'd9, 27'h0000030d, 5'd18, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003b7, 5'd8, 27'h000002f6, 5'd29, 27'h00000300, 32'h00000400,
  1'd1,  5'd26, 27'h0000014c, 5'd18, 27'h000003e9, 5'd9, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000297, 5'd16, 27'h000001d2, 5'd18, 27'h0000007c, 32'h00000400,
  1'd1,  5'd26, 27'h00000001, 5'd15, 27'h000002e0, 5'd27, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000319, 5'd26, 27'h0000033b, 5'd6, 27'h00000097, 32'h00000400,
  1'd1,  5'd28, 27'h000002c4, 5'd26, 27'h0000036c, 5'd18, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000309, 5'd26, 27'h00000352, 5'd26, 27'h000002a2, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000214, 5'd2, 27'h0000028e, 5'd4, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001fe, 5'd0, 27'h000002bd, 5'd10, 27'h0000030d, 32'h00000400,
  1'd1,  5'd4, 27'h0000032b, 5'd4, 27'h000003e9, 5'd24, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000005a, 5'd10, 27'h000003d3, 5'd3, 27'h00000275, 32'h00000400,
  1'd1,  5'd3, 27'h000002a3, 5'd15, 27'h000001d2, 5'd10, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000309, 5'd11, 27'h00000090, 5'd21, 27'h00000029, 32'h00000400,
  1'd1,  5'd2, 27'h000000af, 5'd22, 27'h0000003a, 5'd2, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000116, 5'd23, 27'h0000028c, 5'd13, 27'h00000291, 32'h00000400,
  1'd1,  5'd4, 27'h00000110, 5'd22, 27'h0000008e, 5'd21, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000070, 5'd2, 27'h00000274, 5'd0, 27'h000002b7, 32'h00000400,
  1'd1,  5'd14, 27'h000000f5, 5'd1, 27'h0000024c, 5'd10, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000057, 5'd2, 27'h00000008, 5'd25, 27'h0000009b, 32'h00000400,
  1'd1,  5'd11, 27'h000002bb, 5'd11, 27'h00000124, 5'd1, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001e8, 5'd13, 27'h000002c1, 5'd15, 27'h0000007d, 32'h00000400,
  1'd1,  5'd12, 27'h000000a1, 5'd14, 27'h0000035d, 5'd21, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000032a, 5'd23, 27'h00000191, 5'd4, 27'h00000044, 32'h00000400,
  1'd1,  5'd11, 27'h000000f8, 5'd25, 27'h00000232, 5'd14, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f3, 5'd23, 27'h000002b6, 5'd22, 27'h00000337, 32'h00000400,
  1'd1,  5'd20, 27'h000002ed, 5'd4, 27'h00000182, 5'd4, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000013e, 5'd1, 27'h00000216, 5'd14, 27'h0000004f, 32'h00000400,
  1'd1,  5'd22, 27'h0000018b, 5'd1, 27'h0000037d, 5'd23, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031f, 5'd14, 27'h000001df, 5'd0, 27'h00000197, 32'h00000400,
  1'd1,  5'd22, 27'h00000359, 5'd14, 27'h000001b9, 5'd13, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000180, 5'd12, 27'h00000215, 5'd23, 27'h00000148, 32'h00000400,
  1'd1,  5'd22, 27'h00000249, 5'd24, 27'h0000020a, 5'd1, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000353, 5'd24, 27'h0000000b, 5'd14, 27'h000001c2, 32'h00000400,
  1'd1,  5'd25, 27'h0000034c, 5'd20, 27'h0000035f, 5'd21, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000e5, 5'd1, 27'h000001e6, 5'd6, 27'h000003a2, 32'h00000400,
  1'd1,  5'd4, 27'h0000012e, 5'd2, 27'h0000020f, 5'd16, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001e7, 5'd4, 27'h000000b8, 5'd28, 27'h00000264, 32'h00000400,
  1'd1,  5'd1, 27'h00000230, 5'd10, 27'h00000265, 5'd8, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000303, 5'd13, 27'h00000230, 5'd17, 27'h00000310, 32'h00000400,
  1'd1,  5'd1, 27'h000003e1, 5'd11, 27'h000000f4, 5'd28, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000015c, 5'd21, 27'h00000107, 5'd10, 27'h00000068, 32'h00000400,
  1'd1,  5'd1, 27'h0000039e, 5'd24, 27'h000001cc, 5'd18, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000258, 5'd24, 27'h00000343, 5'd27, 27'h0000010d, 32'h00000400,
  1'd1,  5'd11, 27'h000001f4, 5'd4, 27'h00000324, 5'd8, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000382, 5'd2, 27'h000001db, 5'd18, 27'h00000356, 32'h00000400,
  1'd1,  5'd12, 27'h0000037e, 5'd2, 27'h000003c1, 5'd28, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ea, 5'd14, 27'h0000034d, 5'd6, 27'h000003d6, 32'h00000400,
  1'd1,  5'd12, 27'h000000e1, 5'd13, 27'h000001ec, 5'd20, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000004d, 5'd11, 27'h00000351, 5'd26, 27'h00000057, 32'h00000400,
  1'd1,  5'd12, 27'h00000232, 5'd23, 27'h000002bd, 5'd6, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a2, 5'd24, 27'h0000017e, 5'd19, 27'h000003fc, 32'h00000400,
  1'd1,  5'd11, 27'h0000031b, 5'd23, 27'h00000103, 5'd27, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000380, 5'd2, 27'h00000051, 5'd6, 27'h0000037e, 32'h00000400,
  1'd1,  5'd24, 27'h000000d2, 5'd3, 27'h000000d2, 5'd20, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000313, 5'd1, 27'h00000370, 5'd26, 27'h00000150, 32'h00000400,
  1'd1,  5'd21, 27'h000001b6, 5'd14, 27'h0000025a, 5'd6, 27'h00000173, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000032e, 5'd13, 27'h0000001b, 5'd20, 27'h0000011a, 32'h00000400,
  1'd1,  5'd25, 27'h000000ed, 5'd12, 27'h000003d3, 5'd28, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002f4, 5'd22, 27'h0000006d, 5'd7, 27'h000002da, 32'h00000400,
  1'd1,  5'd21, 27'h000002af, 5'd25, 27'h000002e8, 5'd19, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000d8, 5'd21, 27'h000002a0, 5'd30, 27'h000002b0, 32'h00000400,
  1'd1,  5'd1, 27'h000001ad, 5'd6, 27'h00000240, 5'd2, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e1, 5'd5, 27'h00000175, 5'd15, 27'h000000ed, 32'h00000400,
  1'd1,  5'd0, 27'h00000305, 5'd5, 27'h00000269, 5'd24, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b4, 5'd18, 27'h000000a5, 5'd2, 27'h00000253, 32'h00000400,
  1'd1,  5'd2, 27'h00000346, 5'd16, 27'h000003fa, 5'd11, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000236, 5'd18, 27'h000003cd, 5'd21, 27'h0000013a, 32'h00000400,
  1'd1,  5'd3, 27'h00000232, 5'd26, 27'h00000136, 5'd1, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d5, 5'd29, 27'h0000003b, 5'd14, 27'h00000271, 32'h00000400,
  1'd1,  5'd3, 27'h000001d1, 5'd28, 27'h00000172, 5'd21, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f5, 5'd6, 27'h000002de, 5'd0, 27'h00000117, 32'h00000400,
  1'd1,  5'd14, 27'h00000158, 5'd9, 27'h000003df, 5'd11, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002a1, 5'd7, 27'h00000314, 5'd23, 27'h0000021f, 32'h00000400,
  1'd1,  5'd12, 27'h0000000b, 5'd19, 27'h00000166, 5'd1, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003c2, 5'd19, 27'h00000320, 5'd14, 27'h000003ec, 32'h00000400,
  1'd1,  5'd15, 27'h000000f9, 5'd17, 27'h000002fb, 5'd25, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002da, 5'd26, 27'h0000007e, 5'd4, 27'h00000026, 32'h00000400,
  1'd1,  5'd12, 27'h00000027, 5'd27, 27'h0000005e, 5'd12, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000294, 5'd30, 27'h00000037, 5'd22, 27'h000002ab, 32'h00000400,
  1'd1,  5'd25, 27'h00000309, 5'd5, 27'h00000140, 5'd0, 27'h00000322, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000188, 5'd9, 27'h00000380, 5'd11, 27'h0000001e, 32'h00000400,
  1'd1,  5'd24, 27'h00000343, 5'd7, 27'h00000378, 5'd24, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000208, 5'd18, 27'h000002fa, 5'd4, 27'h00000182, 32'h00000400,
  1'd1,  5'd20, 27'h000003f8, 5'd19, 27'h000000a9, 5'd12, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000175, 5'd20, 27'h00000251, 5'd22, 27'h000002f9, 32'h00000400,
  1'd1,  5'd23, 27'h00000020, 5'd26, 27'h000003ed, 5'd1, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003cc, 5'd26, 27'h000003ac, 5'd14, 27'h00000325, 32'h00000400,
  1'd1,  5'd21, 27'h000002a6, 5'd30, 27'h00000232, 5'd22, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000005d, 5'd6, 27'h000000fb, 5'd5, 27'h000002dc, 32'h00000400,
  1'd1,  5'd1, 27'h000001ca, 5'd7, 27'h000002e7, 5'd20, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000025d, 5'd7, 27'h00000190, 5'd26, 27'h00000158, 32'h00000400,
  1'd1,  5'd4, 27'h000001c3, 5'd19, 27'h000002f3, 5'd5, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000128, 5'd17, 27'h000002dc, 5'd16, 27'h000003c8, 32'h00000400,
  1'd1,  5'd0, 27'h000000da, 5'd18, 27'h0000021e, 5'd28, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e7, 5'd29, 27'h00000152, 5'd8, 27'h00000145, 32'h00000400,
  1'd1,  5'd3, 27'h000003b4, 5'd26, 27'h00000109, 5'd17, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000005b, 5'd26, 27'h00000213, 5'd27, 27'h00000287, 32'h00000400,
  1'd1,  5'd13, 27'h0000012a, 5'd8, 27'h000001bf, 5'd9, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000174, 5'd5, 27'h0000032e, 5'd18, 27'h000002ab, 32'h00000400,
  1'd1,  5'd14, 27'h000001cb, 5'd7, 27'h00000356, 5'd30, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c8, 5'd18, 27'h000003db, 5'd7, 27'h0000016a, 32'h00000400,
  1'd1,  5'd14, 27'h00000216, 5'd18, 27'h00000286, 5'd19, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ca, 5'd15, 27'h0000034d, 5'd30, 27'h00000106, 32'h00000400,
  1'd1,  5'd11, 27'h000002ea, 5'd30, 27'h0000010c, 5'd9, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000031f, 5'd30, 27'h000002ff, 5'd19, 27'h0000003a, 32'h00000400,
  1'd1,  5'd11, 27'h00000017, 5'd26, 27'h00000012, 5'd27, 27'h000001db, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000007e, 5'd8, 27'h00000332, 5'd8, 27'h00000094, 32'h00000400,
  1'd1,  5'd22, 27'h000001ac, 5'd8, 27'h0000010b, 5'd20, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a6, 5'd7, 27'h000001a0, 5'd29, 27'h000000e5, 32'h00000400,
  1'd1,  5'd22, 27'h000000bb, 5'd19, 27'h00000294, 5'd6, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003da, 5'd17, 27'h0000006c, 5'd17, 27'h00000032, 32'h00000400,
  1'd1,  5'd23, 27'h000001a4, 5'd16, 27'h00000264, 5'd27, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000166, 5'd26, 27'h0000024b, 5'd9, 27'h0000013a, 32'h00000400,
  1'd1,  5'd24, 27'h0000012b, 5'd30, 27'h00000255, 5'd17, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000027f, 5'd27, 27'h00000303, 5'd27, 27'h00000271, 32'h00000400,
  1'd1,  5'd5, 27'h0000031b, 5'd2, 27'h00000208, 5'd8, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000b2, 5'd1, 27'h00000270, 5'd16, 27'h00000216, 32'h00000400,
  1'd1,  5'd10, 27'h0000000e, 5'd1, 27'h00000335, 5'd27, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a0, 5'd13, 27'h000001e9, 5'd1, 27'h000000e6, 32'h00000400,
  1'd1,  5'd5, 27'h000000c3, 5'd11, 27'h00000015, 5'd11, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b7, 5'd13, 27'h000002fe, 5'd22, 27'h00000035, 32'h00000400,
  1'd1,  5'd7, 27'h000001b5, 5'd22, 27'h000000e9, 5'd3, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001fd, 5'd24, 27'h000001b8, 5'd14, 27'h000001d0, 32'h00000400,
  1'd1,  5'd6, 27'h000000c3, 5'd24, 27'h0000030d, 5'd21, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000298, 5'd4, 27'h00000290, 5'd8, 27'h000003b6, 32'h00000400,
  1'd1,  5'd19, 27'h000002f2, 5'd4, 27'h00000326, 5'd18, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000053, 5'd0, 27'h00000348, 5'd26, 27'h000003a2, 32'h00000400,
  1'd1,  5'd16, 27'h000002ad, 5'd12, 27'h0000017f, 5'd3, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b1, 5'd14, 27'h0000018e, 5'd14, 27'h00000240, 32'h00000400,
  1'd1,  5'd20, 27'h0000003d, 5'd11, 27'h00000005, 5'd22, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019b, 5'd24, 27'h0000025c, 5'd3, 27'h00000037, 32'h00000400,
  1'd1,  5'd20, 27'h000001cc, 5'd25, 27'h00000198, 5'd15, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000311, 5'd22, 27'h00000170, 5'd22, 27'h00000178, 32'h00000400,
  1'd1,  5'd27, 27'h00000073, 5'd5, 27'h000000a8, 5'd0, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000346, 5'd3, 27'h000001be, 5'd13, 27'h00000327, 32'h00000400,
  1'd1,  5'd28, 27'h00000308, 5'd2, 27'h00000213, 5'd22, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000026e, 5'd14, 27'h000001e5, 5'd0, 27'h00000308, 32'h00000400,
  1'd1,  5'd26, 27'h00000007, 5'd14, 27'h0000004b, 5'd11, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c6, 5'd13, 27'h00000061, 5'd21, 27'h00000350, 32'h00000400,
  1'd1,  5'd27, 27'h000001a8, 5'd25, 27'h00000102, 5'd2, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003f1, 5'd22, 27'h0000021f, 5'd11, 27'h000003d7, 32'h00000400,
  1'd1,  5'd30, 27'h000000a0, 5'd23, 27'h0000012c, 5'd20, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000da, 5'd2, 27'h00000376, 5'd3, 27'h00000393, 32'h00000400,
  1'd1,  5'd7, 27'h000002c9, 5'd2, 27'h000000b2, 5'd11, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003fb, 5'd0, 27'h00000138, 5'd23, 27'h000000d3, 32'h00000400,
  1'd1,  5'd6, 27'h000001c1, 5'd13, 27'h00000052, 5'd5, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c9, 5'd15, 27'h0000005c, 5'd19, 27'h00000115, 32'h00000400,
  1'd1,  5'd7, 27'h0000015d, 5'd12, 27'h000001fb, 5'd26, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002b5, 5'd25, 27'h000001d3, 5'd9, 27'h000001e0, 32'h00000400,
  1'd1,  5'd7, 27'h0000020c, 5'd21, 27'h000000ae, 5'd20, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038c, 5'd25, 27'h000002ba, 5'd29, 27'h000003c0, 32'h00000400,
  1'd1,  5'd18, 27'h000002d3, 5'd3, 27'h000000d3, 5'd1, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f1, 5'd4, 27'h000001a8, 5'd13, 27'h000003a4, 32'h00000400,
  1'd1,  5'd19, 27'h00000087, 5'd3, 27'h00000141, 5'd25, 27'h000002ba, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016e, 5'd15, 27'h000000fc, 5'd8, 27'h0000038f, 32'h00000400,
  1'd1,  5'd18, 27'h000003d6, 5'd14, 27'h00000334, 5'd18, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d0, 5'd15, 27'h00000119, 5'd29, 27'h000003c2, 32'h00000400,
  1'd1,  5'd19, 27'h000000a2, 5'd21, 27'h00000155, 5'd8, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000267, 5'd25, 27'h0000010f, 5'd15, 27'h0000031b, 32'h00000400,
  1'd1,  5'd19, 27'h000000b6, 5'd22, 27'h0000031f, 5'd29, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ee, 5'd4, 27'h0000022e, 5'd8, 27'h000001a1, 32'h00000400,
  1'd1,  5'd30, 27'h0000006d, 5'd1, 27'h000002bd, 5'd18, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000153, 5'd3, 27'h000002b6, 5'd28, 27'h000000c5, 32'h00000400,
  1'd1,  5'd26, 27'h0000038c, 5'd10, 27'h000001ee, 5'd10, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000318, 5'd12, 27'h0000017a, 5'd15, 27'h0000024e, 32'h00000400,
  1'd1,  5'd30, 27'h00000008, 5'd11, 27'h0000027d, 5'd27, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000118, 5'd23, 27'h000001bd, 5'd6, 27'h0000011a, 32'h00000400,
  1'd1,  5'd26, 27'h00000098, 5'd20, 27'h0000035e, 5'd16, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b6, 5'd23, 27'h0000014f, 5'd30, 27'h0000001e, 32'h00000400,
  1'd1,  5'd9, 27'h00000179, 5'd8, 27'h000000f2, 5'd1, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000c9, 5'd8, 27'h00000210, 5'd11, 27'h0000003a, 32'h00000400,
  1'd1,  5'd5, 27'h00000192, 5'd5, 27'h000003f0, 5'd24, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003b4, 5'd18, 27'h000003a3, 5'd3, 27'h00000039, 32'h00000400,
  1'd1,  5'd7, 27'h000000f8, 5'd15, 27'h00000370, 5'd14, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000034b, 5'd18, 27'h00000226, 5'd24, 27'h000000ae, 32'h00000400,
  1'd1,  5'd7, 27'h0000023e, 5'd27, 27'h00000265, 5'd0, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001d3, 5'd26, 27'h0000022c, 5'd13, 27'h000002d0, 32'h00000400,
  1'd1,  5'd8, 27'h00000175, 5'd26, 27'h00000267, 5'd21, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000019f, 5'd9, 27'h00000246, 5'd2, 27'h0000031e, 32'h00000400,
  1'd1,  5'd16, 27'h00000229, 5'd6, 27'h0000027a, 5'd11, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000176, 5'd6, 27'h00000197, 5'd24, 27'h00000368, 32'h00000400,
  1'd1,  5'd17, 27'h0000008d, 5'd16, 27'h000000e1, 5'd3, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000279, 5'd19, 27'h000002d5, 5'd13, 27'h0000021d, 32'h00000400,
  1'd1,  5'd19, 27'h00000032, 5'd17, 27'h0000027f, 5'd23, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000060, 5'd29, 27'h0000008d, 5'd2, 27'h00000353, 32'h00000400,
  1'd1,  5'd17, 27'h00000307, 5'd26, 27'h000000ee, 5'd15, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002b2, 5'd26, 27'h00000238, 5'd23, 27'h0000018a, 32'h00000400,
  1'd1,  5'd28, 27'h000003ff, 5'd7, 27'h000000b0, 5'd1, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000379, 5'd8, 27'h000001de, 5'd11, 27'h000003ba, 32'h00000400,
  1'd1,  5'd26, 27'h00000188, 5'd5, 27'h000002b5, 5'd25, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000119, 5'd18, 27'h00000083, 5'd3, 27'h0000001f, 32'h00000400,
  1'd1,  5'd30, 27'h00000338, 5'd20, 27'h000000ea, 5'd12, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021b, 5'd20, 27'h00000058, 5'd24, 27'h0000001f, 32'h00000400,
  1'd1,  5'd27, 27'h000000ca, 5'd27, 27'h00000082, 5'd4, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000158, 5'd29, 27'h00000098, 5'd13, 27'h0000038e, 32'h00000400,
  1'd1,  5'd28, 27'h000001ef, 5'd26, 27'h0000023c, 5'd22, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000e8, 5'd8, 27'h0000027e, 5'd10, 27'h0000006d, 32'h00000400,
  1'd1,  5'd9, 27'h0000010a, 5'd6, 27'h00000049, 5'd16, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000034, 5'd6, 27'h00000179, 5'd27, 27'h000000a5, 32'h00000400,
  1'd1,  5'd8, 27'h000002cc, 5'd16, 27'h00000157, 5'd5, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000148, 5'd17, 27'h00000342, 5'd17, 27'h00000043, 32'h00000400,
  1'd1,  5'd8, 27'h0000028d, 5'd19, 27'h00000234, 5'd29, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000077, 5'd29, 27'h0000011d, 5'd7, 27'h0000034d, 32'h00000400,
  1'd1,  5'd7, 27'h00000221, 5'd25, 27'h000003e4, 5'd16, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b2, 5'd28, 27'h0000027f, 5'd26, 27'h00000218, 32'h00000400,
  1'd1,  5'd19, 27'h000002b2, 5'd6, 27'h000001cd, 5'd8, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000006b, 5'd10, 27'h0000004a, 5'd17, 27'h000000d3, 32'h00000400,
  1'd1,  5'd15, 27'h00000307, 5'd7, 27'h00000124, 5'd26, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b5, 5'd17, 27'h0000018f, 5'd9, 27'h00000025, 32'h00000400,
  1'd1,  5'd18, 27'h00000152, 5'd18, 27'h0000025d, 5'd17, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002a8, 5'd20, 27'h000001e9, 5'd30, 27'h00000088, 32'h00000400,
  1'd1,  5'd20, 27'h000000a9, 5'd28, 27'h000003b3, 5'd7, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000020c, 5'd27, 27'h000002c1, 5'd18, 27'h00000376, 32'h00000400,
  1'd1,  5'd17, 27'h00000047, 5'd26, 27'h000002ab, 5'd26, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003bd, 5'd10, 27'h00000013, 5'd5, 27'h000003c8, 32'h00000400,
  1'd1,  5'd25, 27'h00000399, 5'd7, 27'h0000036f, 5'd16, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000294, 5'd9, 27'h000003ef, 5'd29, 27'h000000d9, 32'h00000400,
  1'd1,  5'd30, 27'h000001df, 5'd18, 27'h000003fd, 5'd10, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c4, 5'd16, 27'h00000396, 5'd17, 27'h00000211, 32'h00000400,
  1'd1,  5'd27, 27'h0000010d, 5'd19, 27'h000000da, 5'd26, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000187, 5'd26, 27'h000003fb, 5'd10, 27'h0000002d, 32'h00000400,
  1'd1,  5'd30, 27'h00000151, 5'd28, 27'h00000252, 5'd17, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d6, 5'd29, 27'h00000320, 5'd26, 27'h0000033e, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000362, 5'd5, 27'h00000006, 5'd2, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000022c, 5'd2, 27'h0000004f, 5'd14, 27'h00000398, 32'h00000400,
  1'd1,  5'd4, 27'h000002c4, 5'd3, 27'h0000035e, 5'd21, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003fc, 5'd13, 27'h00000055, 5'd0, 27'h00000316, 32'h00000400,
  1'd1,  5'd4, 27'h00000101, 5'd13, 27'h00000023, 5'd12, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000359, 5'd10, 27'h00000330, 5'd20, 27'h000002ad, 32'h00000400,
  1'd1,  5'd3, 27'h000003f4, 5'd21, 27'h00000143, 5'd1, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d6, 5'd22, 27'h00000086, 5'd11, 27'h00000306, 32'h00000400,
  1'd1,  5'd4, 27'h00000032, 5'd25, 27'h000000bd, 5'd21, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000026d, 5'd0, 27'h00000050, 5'd5, 27'h00000060, 32'h00000400,
  1'd1,  5'd13, 27'h0000035d, 5'd4, 27'h000002b5, 5'd10, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000036d, 5'd3, 27'h0000014e, 5'd21, 27'h00000108, 32'h00000400,
  1'd1,  5'd11, 27'h00000021, 5'd13, 27'h00000050, 5'd1, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000077, 5'd14, 27'h0000011d, 5'd10, 27'h00000328, 32'h00000400,
  1'd1,  5'd13, 27'h000001df, 5'd11, 27'h000002ee, 5'd20, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f6, 5'd21, 27'h000000a8, 5'd1, 27'h000001e8, 32'h00000400,
  1'd1,  5'd15, 27'h000000d7, 5'd21, 27'h000003b4, 5'd14, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f6, 5'd21, 27'h000000a4, 5'd22, 27'h000002dc, 32'h00000400,
  1'd1,  5'd22, 27'h0000013e, 5'd4, 27'h0000039c, 5'd0, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001ff, 5'd0, 27'h00000002, 5'd14, 27'h00000208, 32'h00000400,
  1'd1,  5'd21, 27'h00000167, 5'd1, 27'h000000d7, 5'd21, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d8, 5'd12, 27'h00000037, 5'd2, 27'h00000074, 32'h00000400,
  1'd1,  5'd22, 27'h00000321, 5'd12, 27'h00000278, 5'd15, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000367, 5'd11, 27'h0000004c, 5'd21, 27'h00000082, 32'h00000400,
  1'd1,  5'd22, 27'h000002b2, 5'd25, 27'h00000245, 5'd3, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000086, 5'd24, 27'h0000033e, 5'd11, 27'h000001e9, 32'h00000400,
  1'd1,  5'd22, 27'h000000dd, 5'd24, 27'h0000007d, 5'd22, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000026f, 5'd2, 27'h00000151, 5'd6, 27'h00000002, 32'h00000400,
  1'd1,  5'd2, 27'h00000373, 5'd3, 27'h00000336, 5'd16, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f7, 5'd4, 27'h0000026c, 5'd27, 27'h00000370, 32'h00000400,
  1'd1,  5'd2, 27'h000003ef, 5'd13, 27'h000002a9, 5'd8, 27'h0000014a, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000354, 5'd14, 27'h0000025b, 5'd16, 27'h000000af, 32'h00000400,
  1'd1,  5'd2, 27'h00000141, 5'd13, 27'h00000371, 5'd30, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a5, 5'd22, 27'h000002d4, 5'd10, 27'h0000008c, 32'h00000400,
  1'd1,  5'd3, 27'h000002ad, 5'd22, 27'h000002ae, 5'd19, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000062, 5'd23, 27'h00000092, 5'd27, 27'h000000c6, 32'h00000400,
  1'd1,  5'd11, 27'h00000176, 5'd2, 27'h0000023a, 5'd6, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000180, 5'd3, 27'h00000205, 5'd18, 27'h00000060, 32'h00000400,
  1'd1,  5'd11, 27'h000003da, 5'd2, 27'h000001e9, 5'd29, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001e1, 5'd12, 27'h000003a5, 5'd7, 27'h00000281, 32'h00000400,
  1'd1,  5'd13, 27'h00000267, 5'd11, 27'h0000025e, 5'd19, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000335, 5'd10, 27'h00000314, 5'd25, 27'h000003c9, 32'h00000400,
  1'd1,  5'd14, 27'h000002ac, 5'd24, 27'h00000170, 5'd6, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d9, 5'd21, 27'h00000022, 5'd17, 27'h0000013b, 32'h00000400,
  1'd1,  5'd14, 27'h000001f9, 5'd21, 27'h00000239, 5'd29, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000326, 5'd1, 27'h00000203, 5'd7, 27'h00000389, 32'h00000400,
  1'd1,  5'd23, 27'h000001e1, 5'd4, 27'h000003cc, 5'd19, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000018b, 5'd0, 27'h00000212, 5'd26, 27'h000003b5, 32'h00000400,
  1'd1,  5'd21, 27'h000003d2, 5'd11, 27'h000001b1, 5'd5, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b4, 5'd13, 27'h000000bf, 5'd16, 27'h0000004d, 32'h00000400,
  1'd1,  5'd21, 27'h00000303, 5'd12, 27'h00000053, 5'd30, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000093, 5'd25, 27'h000002c3, 5'd6, 27'h00000389, 32'h00000400,
  1'd1,  5'd21, 27'h000001a2, 5'd22, 27'h0000008e, 5'd15, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000f3, 5'd23, 27'h0000033d, 5'd27, 27'h000000bd, 32'h00000400,
  1'd1,  5'd4, 27'h0000011b, 5'd6, 27'h000003af, 5'd1, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f7, 5'd5, 27'h00000303, 5'd12, 27'h00000326, 32'h00000400,
  1'd1,  5'd0, 27'h000001cb, 5'd9, 27'h0000026b, 5'd21, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000373, 5'd18, 27'h00000267, 5'd1, 27'h000003c4, 32'h00000400,
  1'd1,  5'd2, 27'h000002db, 5'd17, 27'h0000026f, 5'd15, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000299, 5'd17, 27'h000001d6, 5'd21, 27'h0000008c, 32'h00000400,
  1'd1,  5'd3, 27'h000003e1, 5'd29, 27'h000000ce, 5'd5, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001df, 5'd26, 27'h000001ef, 5'd10, 27'h00000177, 32'h00000400,
  1'd1,  5'd4, 27'h00000018, 5'd29, 27'h000002c8, 5'd22, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d4, 5'd5, 27'h000003c3, 5'd0, 27'h00000069, 32'h00000400,
  1'd1,  5'd11, 27'h000003f3, 5'd6, 27'h00000147, 5'd11, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000029a, 5'd5, 27'h000002d8, 5'd22, 27'h000000e1, 32'h00000400,
  1'd1,  5'd11, 27'h000000ab, 5'd18, 27'h00000123, 5'd0, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000103, 5'd15, 27'h0000020b, 5'd15, 27'h00000167, 32'h00000400,
  1'd1,  5'd10, 27'h000001ec, 5'd19, 27'h000003fa, 5'd24, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000003a, 5'd27, 27'h0000016f, 5'd3, 27'h0000024c, 32'h00000400,
  1'd1,  5'd14, 27'h00000155, 5'd29, 27'h00000396, 5'd13, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000187, 5'd29, 27'h000002b2, 5'd20, 27'h000002f7, 32'h00000400,
  1'd1,  5'd24, 27'h0000004b, 5'd6, 27'h0000026b, 5'd1, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fd, 5'd7, 27'h00000287, 5'd14, 27'h00000174, 32'h00000400,
  1'd1,  5'd25, 27'h00000330, 5'd9, 27'h0000039e, 5'd21, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000169, 5'd18, 27'h00000294, 5'd0, 27'h0000008b, 32'h00000400,
  1'd1,  5'd23, 27'h000002c2, 5'd15, 27'h00000325, 5'd15, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000201, 5'd18, 27'h00000077, 5'd24, 27'h0000001e, 32'h00000400,
  1'd1,  5'd25, 27'h0000008b, 5'd30, 27'h000001eb, 5'd3, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000334, 5'd26, 27'h0000017b, 5'd10, 27'h000003b9, 32'h00000400,
  1'd1,  5'd20, 27'h000002d8, 5'd29, 27'h0000007d, 5'd23, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d7, 5'd9, 27'h0000023d, 5'd6, 27'h000002b7, 32'h00000400,
  1'd1,  5'd4, 27'h00000210, 5'd9, 27'h00000305, 5'd17, 27'h000001e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000136, 5'd5, 27'h000002e4, 5'd29, 27'h00000363, 32'h00000400,
  1'd1,  5'd0, 27'h000002cd, 5'd16, 27'h00000236, 5'd8, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000025e, 5'd17, 27'h00000243, 5'd16, 27'h00000262, 32'h00000400,
  1'd1,  5'd0, 27'h00000243, 5'd15, 27'h000002e4, 5'd27, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000284, 5'd29, 27'h00000398, 5'd8, 27'h00000381, 32'h00000400,
  1'd1,  5'd2, 27'h000000cc, 5'd27, 27'h000003aa, 5'd16, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000da, 5'd26, 27'h000003af, 5'd26, 27'h00000086, 32'h00000400,
  1'd1,  5'd12, 27'h000002d4, 5'd9, 27'h00000154, 5'd7, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008d, 5'd7, 27'h000002d7, 5'd16, 27'h0000031b, 32'h00000400,
  1'd1,  5'd11, 27'h00000271, 5'd10, 27'h00000058, 5'd27, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000af, 5'd19, 27'h00000119, 5'd8, 27'h00000023, 32'h00000400,
  1'd1,  5'd10, 27'h0000022f, 5'd19, 27'h000002ce, 5'd20, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000157, 5'd18, 27'h000003e9, 5'd30, 27'h0000025f, 32'h00000400,
  1'd1,  5'd15, 27'h00000106, 5'd30, 27'h00000239, 5'd8, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002f4, 5'd27, 27'h0000014f, 5'd18, 27'h000000b1, 32'h00000400,
  1'd1,  5'd13, 27'h00000243, 5'd27, 27'h00000317, 5'd25, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000032c, 5'd7, 27'h000003bd, 5'd6, 27'h00000375, 32'h00000400,
  1'd1,  5'd23, 27'h000000ba, 5'd8, 27'h000001e8, 5'd19, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000323, 5'd9, 27'h00000386, 5'd28, 27'h0000006f, 32'h00000400,
  1'd1,  5'd24, 27'h00000222, 5'd20, 27'h0000010e, 5'd10, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003cd, 5'd18, 27'h0000019b, 5'd19, 27'h00000234, 32'h00000400,
  1'd1,  5'd22, 27'h00000265, 5'd18, 27'h000002b1, 5'd28, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002bb, 5'd28, 27'h00000235, 5'd10, 27'h000000aa, 32'h00000400,
  1'd1,  5'd23, 27'h000000f4, 5'd28, 27'h00000100, 5'd15, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000390, 5'd26, 27'h00000343, 5'd29, 27'h000002c4, 32'h00000400,
  1'd1,  5'd8, 27'h00000346, 5'd0, 27'h000003d1, 5'd8, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000257, 5'd4, 27'h000002ca, 5'd19, 27'h000003cc, 32'h00000400,
  1'd1,  5'd7, 27'h000003b4, 5'd2, 27'h000002dc, 5'd29, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000127, 5'd13, 27'h0000004a, 5'd2, 27'h000003ee, 32'h00000400,
  1'd1,  5'd7, 27'h0000008e, 5'd12, 27'h000003c4, 5'd13, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000008f, 5'd10, 27'h000003ac, 5'd24, 27'h00000011, 32'h00000400,
  1'd1,  5'd9, 27'h000003d3, 5'd23, 27'h000001bb, 5'd3, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002eb, 5'd23, 27'h000000ed, 5'd10, 27'h00000213, 32'h00000400,
  1'd1,  5'd7, 27'h00000136, 5'd24, 27'h000002d9, 5'd21, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003b3, 5'd3, 27'h000003e9, 5'd7, 27'h00000271, 32'h00000400,
  1'd1,  5'd20, 27'h0000023b, 5'd4, 27'h00000165, 5'd16, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000070, 5'd1, 27'h00000168, 5'd28, 27'h000003ce, 32'h00000400,
  1'd1,  5'd17, 27'h00000147, 5'd13, 27'h0000004b, 5'd4, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001fe, 5'd11, 27'h000001e8, 5'd15, 27'h000001bc, 32'h00000400,
  1'd1,  5'd16, 27'h000003c9, 5'd15, 27'h000001d7, 5'd22, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000029, 5'd24, 27'h00000107, 5'd4, 27'h0000021d, 32'h00000400,
  1'd1,  5'd18, 27'h000000ff, 5'd21, 27'h000003fa, 5'd10, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000bc, 5'd21, 27'h0000023e, 5'd23, 27'h0000005a, 32'h00000400,
  1'd1,  5'd30, 27'h00000015, 5'd3, 27'h00000370, 5'd2, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000017e, 5'd3, 27'h0000033a, 5'd11, 27'h000003eb, 32'h00000400,
  1'd1,  5'd30, 27'h0000017c, 5'd3, 27'h00000103, 5'd22, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002bd, 5'd12, 27'h000002de, 5'd4, 27'h000002ba, 32'h00000400,
  1'd1,  5'd27, 27'h000002a5, 5'd13, 27'h00000268, 5'd11, 27'h000003b7, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000d, 5'd14, 27'h00000359, 5'd22, 27'h00000338, 32'h00000400,
  1'd1,  5'd26, 27'h000003a3, 5'd24, 27'h00000295, 5'd3, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001be, 5'd21, 27'h0000035e, 5'd13, 27'h0000030d, 32'h00000400,
  1'd1,  5'd26, 27'h000002db, 5'd23, 27'h0000010a, 5'd25, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a9, 5'd4, 27'h00000320, 5'd2, 27'h00000152, 32'h00000400,
  1'd1,  5'd5, 27'h000003d8, 5'd0, 27'h000002ac, 5'd15, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ec, 5'd3, 27'h00000080, 5'd22, 27'h0000002b, 32'h00000400,
  1'd1,  5'd8, 27'h000001e8, 5'd12, 27'h00000332, 5'd8, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000185, 5'd12, 27'h00000025, 5'd17, 27'h0000017a, 32'h00000400,
  1'd1,  5'd8, 27'h00000265, 5'd10, 27'h000002c3, 5'd30, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000ec, 5'd24, 27'h00000013, 5'd5, 27'h000001a5, 32'h00000400,
  1'd1,  5'd9, 27'h0000035d, 5'd25, 27'h000002f4, 5'd16, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ac, 5'd22, 27'h000002b2, 5'd27, 27'h0000000f, 32'h00000400,
  1'd1,  5'd19, 27'h0000027d, 5'd3, 27'h000002e8, 5'd0, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000314, 5'd0, 27'h000002d8, 5'd12, 27'h00000189, 32'h00000400,
  1'd1,  5'd18, 27'h0000039f, 5'd1, 27'h00000315, 5'd23, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a6, 5'd14, 27'h000002a3, 5'd9, 27'h00000208, 32'h00000400,
  1'd1,  5'd16, 27'h000003a3, 5'd12, 27'h000001fa, 5'd17, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000019b, 5'd12, 27'h000001df, 5'd27, 27'h000000f4, 32'h00000400,
  1'd1,  5'd18, 27'h00000089, 5'd22, 27'h000001d9, 5'd9, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000030, 5'd23, 27'h000001a2, 5'd20, 27'h000001f6, 32'h00000400,
  1'd1,  5'd17, 27'h000000cc, 5'd25, 27'h00000121, 5'd25, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000041, 5'd4, 27'h000002db, 5'd9, 27'h00000060, 32'h00000400,
  1'd1,  5'd27, 27'h0000025d, 5'd0, 27'h00000028, 5'd20, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a2, 5'd5, 27'h0000003a, 5'd27, 27'h000002d7, 32'h00000400,
  1'd1,  5'd25, 27'h000003cd, 5'd11, 27'h00000397, 5'd5, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000ae, 5'd11, 27'h0000005f, 5'd16, 27'h000003c3, 32'h00000400,
  1'd1,  5'd27, 27'h000001b7, 5'd14, 27'h000002a3, 5'd29, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000362, 5'd21, 27'h000001fc, 5'd8, 27'h000001d7, 32'h00000400,
  1'd1,  5'd30, 27'h000002cf, 5'd21, 27'h000003de, 5'd16, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000307, 5'd22, 27'h000000af, 5'd26, 27'h00000119, 32'h00000400,
  1'd1,  5'd5, 27'h000002a8, 5'd8, 27'h000001c6, 5'd4, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000091, 5'd5, 27'h000001ce, 5'd13, 27'h00000100, 32'h00000400,
  1'd1,  5'd9, 27'h000000b8, 5'd8, 27'h000000a7, 5'd22, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000220, 5'd18, 27'h0000037a, 5'd1, 27'h00000288, 32'h00000400,
  1'd1,  5'd5, 27'h000003a9, 5'd16, 27'h000003c0, 5'd13, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032f, 5'd17, 27'h00000238, 5'd25, 27'h00000255, 32'h00000400,
  1'd1,  5'd5, 27'h000003b2, 5'd28, 27'h00000228, 5'd0, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000037f, 5'd29, 27'h00000267, 5'd13, 27'h00000037, 32'h00000400,
  1'd1,  5'd9, 27'h00000357, 5'd30, 27'h0000034b, 5'd23, 27'h000003e4, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000010f, 5'd7, 27'h00000338, 5'd3, 27'h00000372, 32'h00000400,
  1'd1,  5'd17, 27'h000002b2, 5'd8, 27'h00000171, 5'd10, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000dc, 5'd7, 27'h000001e1, 5'd25, 27'h0000021d, 32'h00000400,
  1'd1,  5'd17, 27'h000001f9, 5'd16, 27'h000003c5, 5'd0, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000dc, 5'd18, 27'h000002c3, 5'd12, 27'h000003d4, 32'h00000400,
  1'd1,  5'd18, 27'h00000025, 5'd19, 27'h000002e9, 5'd24, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002fe, 5'd29, 27'h000003ce, 5'd4, 27'h000003e3, 32'h00000400,
  1'd1,  5'd17, 27'h00000097, 5'd28, 27'h000000cd, 5'd11, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000101, 5'd30, 27'h0000002b, 5'd24, 27'h000003f8, 32'h00000400,
  1'd1,  5'd26, 27'h00000368, 5'd10, 27'h00000021, 5'd3, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002fb, 5'd9, 27'h00000389, 5'd13, 27'h0000007f, 32'h00000400,
  1'd1,  5'd26, 27'h00000017, 5'd9, 27'h0000003f, 5'd24, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000178, 5'd20, 27'h00000173, 5'd3, 27'h000002c8, 32'h00000400,
  1'd1,  5'd26, 27'h00000218, 5'd17, 27'h0000011e, 5'd13, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000184, 5'd19, 27'h000000cd, 5'd20, 27'h000002e9, 32'h00000400,
  1'd1,  5'd27, 27'h00000218, 5'd26, 27'h000003f6, 5'd1, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000394, 5'd26, 27'h0000018f, 5'd10, 27'h00000259, 32'h00000400,
  1'd1,  5'd27, 27'h0000037e, 5'd30, 27'h00000158, 5'd21, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001a8, 5'd8, 27'h000003e7, 5'd9, 27'h000001b8, 32'h00000400,
  1'd1,  5'd8, 27'h00000348, 5'd8, 27'h0000005d, 5'd20, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000174, 5'd6, 27'h00000343, 5'd30, 27'h0000020b, 32'h00000400,
  1'd1,  5'd10, 27'h00000104, 5'd20, 27'h000000ff, 5'd7, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003b6, 5'd16, 27'h00000187, 5'd19, 27'h00000077, 32'h00000400,
  1'd1,  5'd5, 27'h000003a9, 5'd15, 27'h0000030a, 5'd30, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001ef, 5'd27, 27'h0000022c, 5'd8, 27'h000002cf, 32'h00000400,
  1'd1,  5'd7, 27'h000003b3, 5'd29, 27'h00000039, 5'd16, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012f, 5'd27, 27'h000000bd, 5'd28, 27'h0000004d, 32'h00000400,
  1'd1,  5'd20, 27'h00000150, 5'd8, 27'h000001ba, 5'd9, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000281, 5'd7, 27'h000001ec, 5'd17, 27'h00000038, 32'h00000400,
  1'd1,  5'd16, 27'h0000014e, 5'd7, 27'h00000311, 5'd28, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000018e, 5'd18, 27'h000002bc, 5'd7, 27'h00000306, 32'h00000400,
  1'd1,  5'd15, 27'h000003c5, 5'd16, 27'h000001ba, 5'd19, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f5, 5'd19, 27'h000003b5, 5'd28, 27'h000000bf, 32'h00000400,
  1'd1,  5'd19, 27'h0000013b, 5'd29, 27'h0000001b, 5'd6, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c8, 5'd26, 27'h000000cc, 5'd19, 27'h000003f4, 32'h00000400,
  1'd1,  5'd17, 27'h0000006a, 5'd27, 27'h000003bc, 5'd28, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000383, 5'd9, 27'h00000373, 5'd6, 27'h000001f8, 32'h00000400,
  1'd1,  5'd29, 27'h000002b3, 5'd10, 27'h0000001f, 5'd17, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000311, 5'd5, 27'h0000021e, 5'd28, 27'h000003d5, 32'h00000400,
  1'd1,  5'd29, 27'h000002a2, 5'd16, 27'h00000358, 5'd9, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e9, 5'd18, 27'h0000019f, 5'd18, 27'h00000040, 32'h00000400,
  1'd1,  5'd29, 27'h00000359, 5'd20, 27'h00000165, 5'd26, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002cb, 5'd29, 27'h000000b1, 5'd8, 27'h0000012d, 32'h00000400,
  1'd1,  5'd30, 27'h000000fd, 5'd26, 27'h000000d1, 5'd17, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ad, 5'd27, 27'h000001da, 5'd29, 27'h0000002a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000361, 5'd4, 27'h000002c6, 5'd3, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000027a, 5'd4, 27'h000002ec, 5'd11, 27'h00000018, 32'h00000400,
  1'd1,  5'd0, 27'h00000279, 5'd5, 27'h00000064, 5'd23, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002ca, 5'd11, 27'h0000027f, 5'd2, 27'h0000022a, 32'h00000400,
  1'd1,  5'd2, 27'h00000269, 5'd12, 27'h00000286, 5'd15, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000255, 5'd12, 27'h00000029, 5'd23, 27'h000002b6, 32'h00000400,
  1'd1,  5'd1, 27'h000002c8, 5'd22, 27'h000003a1, 5'd0, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000340, 5'd25, 27'h0000034e, 5'd13, 27'h00000025, 32'h00000400,
  1'd1,  5'd0, 27'h00000382, 5'd24, 27'h0000013b, 5'd23, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000015c, 5'd2, 27'h00000191, 5'd2, 27'h00000043, 32'h00000400,
  1'd1,  5'd14, 27'h000002e3, 5'd0, 27'h00000240, 5'd14, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e1, 5'd3, 27'h00000102, 5'd24, 27'h0000005b, 32'h00000400,
  1'd1,  5'd15, 27'h00000061, 5'd10, 27'h000001a1, 5'd0, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000036e, 5'd13, 27'h0000028a, 5'd13, 27'h000001cd, 32'h00000400,
  1'd1,  5'd14, 27'h0000004e, 5'd11, 27'h00000313, 5'd23, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001bb, 5'd20, 27'h000002d2, 5'd4, 27'h000002b5, 32'h00000400,
  1'd1,  5'd13, 27'h00000121, 5'd22, 27'h00000103, 5'd14, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000383, 5'd25, 27'h00000120, 5'd22, 27'h00000303, 32'h00000400,
  1'd1,  5'd21, 27'h0000028d, 5'd1, 27'h000001aa, 5'd4, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003eb, 5'd4, 27'h000000e6, 5'd11, 27'h00000052, 32'h00000400,
  1'd1,  5'd24, 27'h000002ae, 5'd4, 27'h0000026c, 5'd23, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c1, 5'd12, 27'h00000137, 5'd2, 27'h00000125, 32'h00000400,
  1'd1,  5'd23, 27'h00000203, 5'd13, 27'h000000e9, 5'd11, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002eb, 5'd11, 27'h0000023f, 5'd25, 27'h000002cb, 32'h00000400,
  1'd1,  5'd20, 27'h00000305, 5'd21, 27'h0000032e, 5'd2, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000010a, 5'd21, 27'h000000b5, 5'd14, 27'h0000037d, 32'h00000400,
  1'd1,  5'd24, 27'h00000086, 5'd21, 27'h00000288, 5'd24, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003da, 5'd1, 27'h0000001a, 5'd7, 27'h00000077, 32'h00000400,
  1'd1,  5'd1, 27'h000001f3, 5'd1, 27'h00000101, 5'd18, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002c4, 5'd0, 27'h000003e5, 5'd27, 27'h000003ec, 32'h00000400,
  1'd1,  5'd1, 27'h000002e6, 5'd15, 27'h000001ee, 5'd6, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000349, 5'd11, 27'h00000399, 5'd16, 27'h000000bb, 32'h00000400,
  1'd1,  5'd3, 27'h0000007a, 5'd14, 27'h000000c9, 5'd27, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b4, 5'd24, 27'h00000138, 5'd9, 27'h000003ab, 32'h00000400,
  1'd1,  5'd2, 27'h00000062, 5'd23, 27'h00000154, 5'd20, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e8, 5'd23, 27'h0000007b, 5'd30, 27'h0000002c, 32'h00000400,
  1'd1,  5'd10, 27'h000002e2, 5'd1, 27'h00000101, 5'd9, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008b, 5'd2, 27'h0000014e, 5'd18, 27'h0000022c, 32'h00000400,
  1'd1,  5'd15, 27'h000000fb, 5'd1, 27'h000000e8, 5'd30, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000f4, 5'd10, 27'h00000224, 5'd6, 27'h00000239, 32'h00000400,
  1'd1,  5'd11, 27'h000002ba, 5'd13, 27'h000003b3, 5'd19, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ec, 5'd11, 27'h00000210, 5'd29, 27'h00000295, 32'h00000400,
  1'd1,  5'd13, 27'h0000016c, 5'd23, 27'h000000d2, 5'd8, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000b3, 5'd21, 27'h000002dd, 5'd19, 27'h0000012c, 32'h00000400,
  1'd1,  5'd15, 27'h0000014a, 5'd24, 27'h0000022c, 5'd28, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000149, 5'd2, 27'h0000005d, 5'd5, 27'h0000028a, 32'h00000400,
  1'd1,  5'd22, 27'h0000016f, 5'd4, 27'h000001e1, 5'd17, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002df, 5'd0, 27'h0000010c, 5'd30, 27'h0000037b, 32'h00000400,
  1'd1,  5'd23, 27'h000001d3, 5'd11, 27'h000002f8, 5'd9, 27'h000001c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000013a, 5'd11, 27'h000000ba, 5'd18, 27'h00000130, 32'h00000400,
  1'd1,  5'd22, 27'h00000295, 5'd11, 27'h0000038e, 5'd30, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000389, 5'd25, 27'h0000032e, 5'd9, 27'h0000016b, 32'h00000400,
  1'd1,  5'd24, 27'h0000014a, 5'd21, 27'h000002e8, 5'd16, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000e5, 5'd24, 27'h00000057, 5'd30, 27'h00000276, 32'h00000400,
  1'd1,  5'd1, 27'h0000019d, 5'd6, 27'h000003b7, 5'd1, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000001c, 5'd8, 27'h000002c0, 5'd13, 27'h00000205, 32'h00000400,
  1'd1,  5'd2, 27'h000002d9, 5'd8, 27'h000000ad, 5'd22, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003b7, 5'd19, 27'h0000024c, 5'd3, 27'h00000176, 32'h00000400,
  1'd1,  5'd2, 27'h00000312, 5'd15, 27'h0000039f, 5'd10, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000399, 5'd19, 27'h0000010d, 5'd22, 27'h00000246, 32'h00000400,
  1'd1,  5'd1, 27'h00000330, 5'd29, 27'h00000062, 5'd1, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000021a, 5'd29, 27'h0000003c, 5'd15, 27'h000001cb, 32'h00000400,
  1'd1,  5'd2, 27'h0000016b, 5'd27, 27'h00000221, 5'd23, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000002e, 5'd6, 27'h00000273, 5'd2, 27'h000001f8, 32'h00000400,
  1'd1,  5'd14, 27'h0000006b, 5'd9, 27'h00000186, 5'd12, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ab, 5'd9, 27'h000000db, 5'd23, 27'h000002c7, 32'h00000400,
  1'd1,  5'd14, 27'h000000df, 5'd20, 27'h00000198, 5'd0, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000023a, 5'd18, 27'h00000187, 5'd15, 27'h000000ff, 32'h00000400,
  1'd1,  5'd12, 27'h000003b0, 5'd16, 27'h00000053, 5'd24, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000378, 5'd26, 27'h0000000d, 5'd2, 27'h00000249, 32'h00000400,
  1'd1,  5'd11, 27'h00000141, 5'd30, 27'h0000037a, 5'd10, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002b1, 5'd27, 27'h0000009e, 5'd22, 27'h00000244, 32'h00000400,
  1'd1,  5'd24, 27'h00000106, 5'd7, 27'h000001a5, 5'd2, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000055, 5'd8, 27'h00000181, 5'd10, 27'h00000374, 32'h00000400,
  1'd1,  5'd25, 27'h0000020a, 5'd8, 27'h000001dd, 5'd24, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003d1, 5'd19, 27'h000000ad, 5'd3, 27'h0000029c, 32'h00000400,
  1'd1,  5'd23, 27'h00000292, 5'd17, 27'h00000372, 5'd13, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002aa, 5'd20, 27'h0000025c, 5'd24, 27'h0000015f, 32'h00000400,
  1'd1,  5'd21, 27'h00000394, 5'd30, 27'h000000fd, 5'd4, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b7, 5'd26, 27'h000002ef, 5'd15, 27'h000000f1, 32'h00000400,
  1'd1,  5'd21, 27'h00000037, 5'd28, 27'h0000014c, 5'd25, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000259, 5'd7, 27'h00000218, 5'd7, 27'h00000196, 32'h00000400,
  1'd1,  5'd1, 27'h000002fe, 5'd7, 27'h0000006d, 5'd16, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000106, 5'd6, 27'h00000162, 5'd28, 27'h000003c0, 32'h00000400,
  1'd1,  5'd5, 27'h0000007e, 5'd16, 27'h0000034e, 5'd6, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001c2, 5'd16, 27'h0000018f, 5'd15, 27'h00000217, 32'h00000400,
  1'd1,  5'd3, 27'h000003d7, 5'd16, 27'h00000160, 5'd27, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000aa, 5'd27, 27'h00000031, 5'd8, 27'h00000066, 32'h00000400,
  1'd1,  5'd0, 27'h000000de, 5'd30, 27'h00000238, 5'd15, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027f, 5'd26, 27'h0000007d, 5'd30, 27'h00000233, 32'h00000400,
  1'd1,  5'd11, 27'h000000a3, 5'd7, 27'h00000123, 5'd7, 27'h000003d1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000003e, 5'd7, 27'h000001a5, 5'd18, 27'h0000016a, 32'h00000400,
  1'd1,  5'd11, 27'h00000235, 5'd7, 27'h00000312, 5'd30, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001bc, 5'd20, 27'h0000027f, 5'd10, 27'h00000049, 32'h00000400,
  1'd1,  5'd13, 27'h000001e8, 5'd15, 27'h0000034d, 5'd20, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003d8, 5'd18, 27'h000003f0, 5'd29, 27'h0000030e, 32'h00000400,
  1'd1,  5'd12, 27'h000003ab, 5'd29, 27'h0000038a, 5'd9, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000cb, 5'd26, 27'h000001a6, 5'd19, 27'h000001bc, 32'h00000400,
  1'd1,  5'd11, 27'h000002d5, 5'd27, 27'h00000296, 5'd27, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000288, 5'd10, 27'h000000cc, 5'd6, 27'h00000244, 32'h00000400,
  1'd1,  5'd24, 27'h000000f9, 5'd9, 27'h000000ac, 5'd18, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000307, 5'd7, 27'h0000029e, 5'd30, 27'h00000237, 32'h00000400,
  1'd1,  5'd23, 27'h00000086, 5'd19, 27'h000001fa, 5'd7, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000333, 5'd19, 27'h000001cb, 5'd15, 27'h00000337, 32'h00000400,
  1'd1,  5'd23, 27'h000001b7, 5'd19, 27'h000000ae, 5'd30, 27'h0000036d, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035a, 5'd26, 27'h000002b7, 5'd8, 27'h0000016f, 32'h00000400,
  1'd1,  5'd22, 27'h00000235, 5'd26, 27'h000001ac, 5'd17, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000378, 5'd30, 27'h00000045, 5'd30, 27'h000003cf, 32'h00000400,
  1'd1,  5'd9, 27'h00000235, 5'd4, 27'h000001bd, 5'd8, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000000a, 5'd1, 27'h00000083, 5'd19, 27'h000003ef, 32'h00000400,
  1'd1,  5'd7, 27'h00000043, 5'd1, 27'h00000106, 5'd28, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a4, 5'd14, 27'h000002d1, 5'd3, 27'h00000098, 32'h00000400,
  1'd1,  5'd5, 27'h00000342, 5'd15, 27'h000000d3, 5'd13, 27'h000000dc, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000220, 5'd12, 27'h00000269, 5'd22, 27'h0000004b, 32'h00000400,
  1'd1,  5'd7, 27'h0000022f, 5'd22, 27'h00000111, 5'd1, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000021d, 5'd24, 27'h0000031b, 5'd11, 27'h0000029f, 32'h00000400,
  1'd1,  5'd8, 27'h000000fa, 5'd23, 27'h0000003d, 5'd23, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030b, 5'd1, 27'h000000b1, 5'd9, 27'h00000236, 32'h00000400,
  1'd1,  5'd17, 27'h000000e6, 5'd1, 27'h00000395, 5'd16, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a9, 5'd1, 27'h0000009d, 5'd28, 27'h000001c1, 32'h00000400,
  1'd1,  5'd15, 27'h0000029e, 5'd11, 27'h000003f3, 5'd2, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000000e, 5'd14, 27'h000000a0, 5'd10, 27'h00000345, 32'h00000400,
  1'd1,  5'd17, 27'h00000047, 5'd11, 27'h00000162, 5'd23, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003d3, 5'd24, 27'h000003e5, 5'd2, 27'h00000341, 32'h00000400,
  1'd1,  5'd16, 27'h0000030c, 5'd23, 27'h0000020d, 5'd14, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000005d, 5'd23, 27'h00000209, 5'd23, 27'h00000105, 32'h00000400,
  1'd1,  5'd27, 27'h000002a3, 5'd2, 27'h00000118, 5'd3, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ba, 5'd1, 27'h000001a5, 5'd13, 27'h00000034, 32'h00000400,
  1'd1,  5'd27, 27'h00000109, 5'd0, 27'h000003f7, 5'd25, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000032a, 5'd11, 27'h0000007e, 5'd0, 27'h00000391, 32'h00000400,
  1'd1,  5'd30, 27'h000000a4, 5'd11, 27'h00000287, 5'd11, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003f7, 5'd10, 27'h000002f1, 5'd23, 27'h0000035c, 32'h00000400,
  1'd1,  5'd27, 27'h0000025d, 5'd22, 27'h00000313, 5'd3, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000031a, 5'd24, 27'h0000006e, 5'd14, 27'h000002fe, 32'h00000400,
  1'd1,  5'd28, 27'h000000a6, 5'd23, 27'h000001dc, 5'd21, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000185, 5'd2, 27'h00000380, 5'd2, 27'h00000093, 32'h00000400,
  1'd1,  5'd6, 27'h000002bc, 5'd4, 27'h000000c9, 5'd13, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002b4, 5'd2, 27'h000002c3, 5'd22, 27'h00000320, 32'h00000400,
  1'd1,  5'd6, 27'h000002fe, 5'd10, 27'h000003c8, 5'd6, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000294, 5'd15, 27'h0000015c, 5'd16, 27'h00000054, 32'h00000400,
  1'd1,  5'd5, 27'h00000392, 5'd11, 27'h0000036b, 5'd30, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000035c, 5'd23, 27'h000002ea, 5'd9, 27'h000001e9, 32'h00000400,
  1'd1,  5'd8, 27'h000003f5, 5'd24, 27'h000000db, 5'd15, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002ff, 5'd20, 27'h000003cc, 5'd25, 27'h00000383, 32'h00000400,
  1'd1,  5'd16, 27'h00000255, 5'd1, 27'h00000223, 5'd4, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000060, 5'd1, 27'h000002cd, 5'd12, 27'h000003ce, 32'h00000400,
  1'd1,  5'd16, 27'h0000018f, 5'd4, 27'h000001b1, 5'd21, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001c, 5'd14, 27'h000000c5, 5'd6, 27'h000002ae, 32'h00000400,
  1'd1,  5'd18, 27'h000002b4, 5'd13, 27'h000001ca, 5'd16, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000033a, 5'd13, 27'h000000bb, 5'd26, 27'h00000184, 32'h00000400,
  1'd1,  5'd19, 27'h000003fd, 5'd22, 27'h0000029b, 5'd9, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000282, 5'd25, 27'h00000145, 5'd19, 27'h00000088, 32'h00000400,
  1'd1,  5'd15, 27'h0000037a, 5'd21, 27'h000000ff, 5'd27, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000334, 5'd1, 27'h000002ab, 5'd9, 27'h000001a0, 32'h00000400,
  1'd1,  5'd29, 27'h00000049, 5'd1, 27'h000001ab, 5'd17, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000018f, 5'd4, 27'h00000266, 5'd30, 27'h000002c0, 32'h00000400,
  1'd1,  5'd28, 27'h00000375, 5'd11, 27'h000001ba, 5'd5, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e5, 5'd13, 27'h00000209, 5'd20, 27'h0000024e, 32'h00000400,
  1'd1,  5'd30, 27'h000003a6, 5'd14, 27'h0000015c, 5'd26, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002ff, 5'd25, 27'h000001d6, 5'd8, 27'h0000039f, 32'h00000400,
  1'd1,  5'd26, 27'h000002ba, 5'd20, 27'h00000348, 5'd16, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000076, 5'd22, 27'h000002fe, 5'd28, 27'h00000028, 32'h00000400,
  1'd1,  5'd5, 27'h000003e1, 5'd5, 27'h000002e8, 5'd2, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000082, 5'd6, 27'h000001a2, 5'd10, 27'h000003a4, 32'h00000400,
  1'd1,  5'd8, 27'h000001fd, 5'd9, 27'h00000132, 5'd24, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000290, 5'd19, 27'h00000283, 5'd2, 27'h00000246, 32'h00000400,
  1'd1,  5'd9, 27'h000002f0, 5'd19, 27'h0000022f, 5'd13, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c2, 5'd18, 27'h0000013d, 5'd23, 27'h0000009f, 32'h00000400,
  1'd1,  5'd7, 27'h00000051, 5'd29, 27'h000003c3, 5'd1, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000013b, 5'd28, 27'h00000182, 5'd10, 27'h0000025e, 32'h00000400,
  1'd1,  5'd5, 27'h00000177, 5'd30, 27'h00000135, 5'd25, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002bc, 5'd7, 27'h00000330, 5'd1, 27'h00000354, 32'h00000400,
  1'd1,  5'd18, 27'h000002e0, 5'd9, 27'h000001ef, 5'd11, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ed, 5'd7, 27'h00000279, 5'd23, 27'h000002a4, 32'h00000400,
  1'd1,  5'd19, 27'h0000026a, 5'd20, 27'h000001df, 5'd0, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000177, 5'd16, 27'h00000044, 5'd13, 27'h0000023d, 32'h00000400,
  1'd1,  5'd18, 27'h00000263, 5'd19, 27'h00000256, 5'd22, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001c8, 5'd29, 27'h00000216, 5'd1, 27'h00000066, 32'h00000400,
  1'd1,  5'd19, 27'h00000026, 5'd30, 27'h00000145, 5'd11, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000386, 5'd26, 27'h00000160, 5'd21, 27'h000001bc, 32'h00000400,
  1'd1,  5'd29, 27'h000001d2, 5'd7, 27'h00000275, 5'd1, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000cc, 5'd6, 27'h000002ee, 5'd11, 27'h0000036b, 32'h00000400,
  1'd1,  5'd29, 27'h000001b8, 5'd9, 27'h00000335, 5'd22, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000333, 5'd15, 27'h00000372, 5'd4, 27'h000001f3, 32'h00000400,
  1'd1,  5'd30, 27'h00000297, 5'd16, 27'h000001ac, 5'd11, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000075, 5'd18, 27'h00000320, 5'd23, 27'h000003b8, 32'h00000400,
  1'd1,  5'd28, 27'h00000223, 5'd30, 27'h000001f6, 5'd0, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000c7, 5'd26, 27'h00000168, 5'd11, 27'h00000163, 32'h00000400,
  1'd1,  5'd30, 27'h00000039, 5'd28, 27'h00000210, 5'd21, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003e2, 5'd6, 27'h000000ba, 5'd7, 27'h000000ce, 32'h00000400,
  1'd1,  5'd7, 27'h0000037c, 5'd6, 27'h0000021e, 5'd18, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000037, 5'd10, 27'h0000007c, 5'd30, 27'h00000316, 32'h00000400,
  1'd1,  5'd7, 27'h0000013d, 5'd19, 27'h00000267, 5'd9, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f5, 5'd20, 27'h000001a0, 5'd19, 27'h0000012e, 32'h00000400,
  1'd1,  5'd8, 27'h0000022e, 5'd17, 27'h000003be, 5'd26, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000374, 5'd30, 27'h0000036f, 5'd9, 27'h000002f9, 32'h00000400,
  1'd1,  5'd8, 27'h00000366, 5'd30, 27'h000000d8, 5'd16, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000335, 5'd29, 27'h00000168, 5'd27, 27'h000001b8, 32'h00000400,
  1'd1,  5'd18, 27'h000003a0, 5'd6, 27'h000001eb, 5'd7, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000018, 5'd6, 27'h0000028d, 5'd17, 27'h000000d9, 32'h00000400,
  1'd1,  5'd19, 27'h00000147, 5'd9, 27'h00000025, 5'd28, 27'h00000084, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000f9, 5'd19, 27'h000001af, 5'd6, 27'h00000010, 32'h00000400,
  1'd1,  5'd15, 27'h00000306, 5'd18, 27'h00000063, 5'd15, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000004e, 5'd18, 27'h000003d4, 5'd27, 27'h000001c7, 32'h00000400,
  1'd1,  5'd20, 27'h00000127, 5'd26, 27'h00000066, 5'd5, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000a3, 5'd27, 27'h00000276, 5'd17, 27'h000000b0, 32'h00000400,
  1'd1,  5'd20, 27'h00000059, 5'd26, 27'h000000dc, 5'd27, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a1, 5'd8, 27'h00000042, 5'd5, 27'h00000173, 32'h00000400,
  1'd1,  5'd30, 27'h000003b7, 5'd5, 27'h000002da, 5'd19, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000331, 5'd7, 27'h00000249, 5'd25, 27'h0000039d, 32'h00000400,
  1'd1,  5'd28, 27'h0000004c, 5'd20, 27'h00000249, 5'd9, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003aa, 5'd16, 27'h00000281, 5'd20, 27'h000002aa, 32'h00000400,
  1'd1,  5'd26, 27'h000000ef, 5'd20, 27'h000001ef, 5'd30, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001d9, 5'd30, 27'h0000019e, 5'd9, 27'h00000324, 32'h00000400,
  1'd1,  5'd28, 27'h0000022a, 5'd30, 27'h000000fe, 5'd19, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000208, 5'd29, 27'h000000f1, 5'd26, 27'h00000167, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000001a1, 5'd2, 27'h000000b6, 5'd4, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f7, 5'd4, 27'h00000161, 5'd10, 27'h00000215, 32'h00000400,
  1'd1,  5'd4, 27'h00000281, 5'd2, 27'h000000ab, 5'd22, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000034b, 5'd12, 27'h0000014c, 5'd0, 27'h0000009c, 32'h00000400,
  1'd1,  5'd1, 27'h0000012c, 5'd14, 27'h000001ca, 5'd15, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003eb, 5'd14, 27'h0000020a, 5'd21, 27'h0000008c, 32'h00000400,
  1'd1,  5'd4, 27'h000003dc, 5'd24, 27'h0000038a, 5'd4, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000386, 5'd25, 27'h0000006f, 5'd11, 27'h000001b6, 32'h00000400,
  1'd1,  5'd0, 27'h000003d7, 5'd21, 27'h00000054, 5'd21, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000a6, 5'd0, 27'h00000221, 5'd0, 27'h0000002f, 32'h00000400,
  1'd1,  5'd13, 27'h00000310, 5'd1, 27'h00000379, 5'd10, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000104, 5'd4, 27'h0000000e, 5'd25, 27'h00000346, 32'h00000400,
  1'd1,  5'd14, 27'h0000031b, 5'd10, 27'h00000386, 5'd1, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e9, 5'd13, 27'h000002b2, 5'd11, 27'h0000021a, 32'h00000400,
  1'd1,  5'd12, 27'h000000ae, 5'd14, 27'h000002a0, 5'd22, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d3, 5'd22, 27'h00000268, 5'd0, 27'h00000302, 32'h00000400,
  1'd1,  5'd14, 27'h00000298, 5'd25, 27'h00000201, 5'd13, 27'h00000396, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001d3, 5'd22, 27'h000001e5, 5'd25, 27'h000002c9, 32'h00000400,
  1'd1,  5'd25, 27'h00000185, 5'd3, 27'h0000024e, 5'd1, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000033b, 5'd5, 27'h00000002, 5'd13, 27'h00000313, 32'h00000400,
  1'd1,  5'd21, 27'h000002d3, 5'd4, 27'h00000098, 5'd24, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000203, 5'd12, 27'h000002bc, 5'd4, 27'h00000350, 32'h00000400,
  1'd1,  5'd24, 27'h000002a8, 5'd14, 27'h000003be, 5'd11, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000b9, 5'd10, 27'h00000362, 5'd25, 27'h000000d4, 32'h00000400,
  1'd1,  5'd21, 27'h000000aa, 5'd22, 27'h0000027c, 5'd0, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000b8, 5'd21, 27'h0000009b, 5'd14, 27'h000001f9, 32'h00000400,
  1'd1,  5'd22, 27'h000003fd, 5'd24, 27'h000003e4, 5'd22, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f3, 5'd0, 27'h0000036e, 5'd8, 27'h0000037b, 32'h00000400,
  1'd1,  5'd5, 27'h0000004a, 5'd0, 27'h0000000c, 5'd19, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ef, 5'd4, 27'h0000009b, 5'd26, 27'h000001f0, 32'h00000400,
  1'd1,  5'd0, 27'h000001ab, 5'd10, 27'h0000027b, 5'd8, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000036, 5'd11, 27'h00000321, 5'd15, 27'h000003ae, 32'h00000400,
  1'd1,  5'd4, 27'h000003eb, 5'd14, 27'h00000025, 5'd26, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000010a, 5'd21, 27'h00000084, 5'd7, 27'h000003b2, 32'h00000400,
  1'd1,  5'd4, 27'h00000062, 5'd22, 27'h00000269, 5'd16, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000001, 5'd23, 27'h00000118, 5'd29, 27'h0000026c, 32'h00000400,
  1'd1,  5'd11, 27'h00000201, 5'd0, 27'h000003dd, 5'd9, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003ad, 5'd0, 27'h0000009d, 5'd17, 27'h00000397, 32'h00000400,
  1'd1,  5'd14, 27'h00000341, 5'd2, 27'h000000bc, 5'd27, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000022e, 5'd12, 27'h000000d2, 5'd7, 27'h000002f7, 32'h00000400,
  1'd1,  5'd13, 27'h00000326, 5'd15, 27'h000000c8, 5'd18, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000291, 5'd12, 27'h000000d6, 5'd27, 27'h00000177, 32'h00000400,
  1'd1,  5'd14, 27'h000000f0, 5'd21, 27'h0000003c, 5'd9, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000020e, 5'd21, 27'h0000023f, 5'd19, 27'h00000242, 32'h00000400,
  1'd1,  5'd14, 27'h00000048, 5'd25, 27'h00000244, 5'd26, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000330, 5'd3, 27'h000002a2, 5'd6, 27'h000001bf, 32'h00000400,
  1'd1,  5'd22, 27'h00000378, 5'd1, 27'h000003bd, 5'd18, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000074, 5'd0, 27'h00000311, 5'd29, 27'h000003ce, 32'h00000400,
  1'd1,  5'd21, 27'h00000340, 5'd15, 27'h00000064, 5'd9, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002c4, 5'd11, 27'h0000018c, 5'd20, 27'h00000187, 32'h00000400,
  1'd1,  5'd21, 27'h000000fa, 5'd12, 27'h00000246, 5'd29, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000009f, 5'd24, 27'h000000d9, 5'd7, 27'h000000bb, 32'h00000400,
  1'd1,  5'd23, 27'h000003ac, 5'd24, 27'h00000241, 5'd16, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000304, 5'd22, 27'h00000292, 5'd27, 27'h0000018c, 32'h00000400,
  1'd1,  5'd3, 27'h0000026b, 5'd6, 27'h0000014f, 5'd3, 27'h00000256, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000392, 5'd9, 27'h00000370, 5'd13, 27'h0000024c, 32'h00000400,
  1'd1,  5'd3, 27'h00000110, 5'd9, 27'h000000fe, 5'd21, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002c1, 5'd19, 27'h000000b4, 5'd3, 27'h00000140, 32'h00000400,
  1'd1,  5'd2, 27'h00000351, 5'd19, 27'h0000011a, 5'd13, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002e8, 5'd17, 27'h00000207, 5'd25, 27'h0000008a, 32'h00000400,
  1'd1,  5'd2, 27'h00000031, 5'd26, 27'h00000098, 5'd0, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002d5, 5'd26, 27'h000002ef, 5'd10, 27'h000001ad, 32'h00000400,
  1'd1,  5'd1, 27'h00000197, 5'd30, 27'h000003e1, 5'd25, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000037f, 5'd8, 27'h00000107, 5'd3, 27'h000001fb, 32'h00000400,
  1'd1,  5'd10, 27'h000002de, 5'd7, 27'h000002e4, 5'd10, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000226, 5'd9, 27'h000001aa, 5'd21, 27'h000000c4, 32'h00000400,
  1'd1,  5'd14, 27'h000003a7, 5'd15, 27'h000003d0, 5'd3, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003eb, 5'd18, 27'h00000225, 5'd10, 27'h00000326, 32'h00000400,
  1'd1,  5'd14, 27'h0000030e, 5'd17, 27'h000000b3, 5'd23, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000030f, 5'd29, 27'h0000016d, 5'd3, 27'h000000c4, 32'h00000400,
  1'd1,  5'd12, 27'h00000229, 5'd29, 27'h00000131, 5'd13, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d2, 5'd28, 27'h000002a1, 5'd24, 27'h00000286, 32'h00000400,
  1'd1,  5'd22, 27'h000002b6, 5'd9, 27'h00000323, 5'd4, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000354, 5'd6, 27'h000000b8, 5'd13, 27'h000003c6, 32'h00000400,
  1'd1,  5'd22, 27'h00000130, 5'd7, 27'h00000373, 5'd22, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ee, 5'd15, 27'h000002bc, 5'd3, 27'h000001cd, 32'h00000400,
  1'd1,  5'd22, 27'h000002ba, 5'd15, 27'h000003e3, 5'd12, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ee, 5'd17, 27'h0000008e, 5'd21, 27'h00000011, 32'h00000400,
  1'd1,  5'd22, 27'h00000315, 5'd29, 27'h00000085, 5'd3, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001d6, 5'd29, 27'h0000001f, 5'd10, 27'h0000035e, 32'h00000400,
  1'd1,  5'd25, 27'h00000087, 5'd29, 27'h00000069, 5'd23, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000035, 5'd5, 27'h000002dc, 5'd9, 27'h00000074, 32'h00000400,
  1'd1,  5'd0, 27'h00000049, 5'd8, 27'h0000005b, 5'd17, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f0, 5'd8, 27'h000002de, 5'd29, 27'h000003b6, 32'h00000400,
  1'd1,  5'd1, 27'h00000094, 5'd18, 27'h00000062, 5'd8, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000013a, 5'd18, 27'h000001ac, 5'd16, 27'h00000307, 32'h00000400,
  1'd1,  5'd1, 27'h0000003a, 5'd20, 27'h00000104, 5'd29, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001bb, 5'd29, 27'h000001f6, 5'd7, 27'h000003f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000141, 5'd30, 27'h00000397, 5'd18, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029c, 5'd30, 27'h0000037b, 5'd28, 27'h00000298, 32'h00000400,
  1'd1,  5'd13, 27'h0000036f, 5'd6, 27'h00000386, 5'd6, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000286, 5'd6, 27'h00000148, 5'd17, 27'h000001d1, 32'h00000400,
  1'd1,  5'd14, 27'h000001de, 5'd6, 27'h00000018, 5'd29, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000181, 5'd15, 27'h00000281, 5'd5, 27'h000001ad, 32'h00000400,
  1'd1,  5'd10, 27'h00000240, 5'd19, 27'h00000377, 5'd16, 27'h00000073, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000008a, 5'd18, 27'h00000049, 5'd29, 27'h000001f3, 32'h00000400,
  1'd1,  5'd14, 27'h0000012b, 5'd29, 27'h000003cf, 5'd5, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c3, 5'd30, 27'h00000105, 5'd17, 27'h00000354, 32'h00000400,
  1'd1,  5'd14, 27'h00000352, 5'd29, 27'h00000156, 5'd30, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003c5, 5'd5, 27'h0000013b, 5'd5, 27'h00000343, 32'h00000400,
  1'd1,  5'd21, 27'h000002de, 5'd7, 27'h0000008d, 5'd19, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000336, 5'd8, 27'h00000319, 5'd30, 27'h000003e5, 32'h00000400,
  1'd1,  5'd23, 27'h000003df, 5'd18, 27'h00000310, 5'd10, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001c4, 5'd18, 27'h00000358, 5'd20, 27'h0000008e, 32'h00000400,
  1'd1,  5'd23, 27'h00000381, 5'd19, 27'h00000182, 5'd30, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e9, 5'd26, 27'h0000013b, 5'd5, 27'h000001bb, 32'h00000400,
  1'd1,  5'd24, 27'h0000024b, 5'd27, 27'h00000059, 5'd18, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001c3, 5'd26, 27'h0000019f, 5'd26, 27'h00000158, 32'h00000400,
  1'd1,  5'd9, 27'h00000053, 5'd0, 27'h0000012c, 5'd8, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003c2, 5'd2, 27'h000002ba, 5'd16, 27'h0000032b, 32'h00000400,
  1'd1,  5'd7, 27'h00000321, 5'd1, 27'h000002aa, 5'd27, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001f3, 5'd11, 27'h00000098, 5'd3, 27'h00000260, 32'h00000400,
  1'd1,  5'd8, 27'h000000b1, 5'd12, 27'h00000020, 5'd15, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000210, 5'd12, 27'h00000257, 5'd24, 27'h000001a0, 32'h00000400,
  1'd1,  5'd7, 27'h00000275, 5'd25, 27'h0000007e, 5'd0, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000263, 5'd23, 27'h000000b3, 5'd13, 27'h0000015e, 32'h00000400,
  1'd1,  5'd6, 27'h000003aa, 5'd25, 27'h00000170, 5'd24, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ed, 5'd0, 27'h0000002a, 5'd10, 27'h000000c7, 32'h00000400,
  1'd1,  5'd15, 27'h0000021d, 5'd2, 27'h00000253, 5'd17, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000220, 5'd3, 27'h00000052, 5'd26, 27'h000001a7, 32'h00000400,
  1'd1,  5'd20, 27'h0000001c, 5'd13, 27'h00000334, 5'd4, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d7, 5'd12, 27'h000003a8, 5'd11, 27'h000002a3, 32'h00000400,
  1'd1,  5'd18, 27'h000000ea, 5'd11, 27'h000002a7, 5'd22, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000016, 5'd24, 27'h0000013b, 5'd4, 27'h00000362, 32'h00000400,
  1'd1,  5'd19, 27'h0000003e, 5'd21, 27'h000003d0, 5'd10, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000028d, 5'd22, 27'h000001ad, 5'd20, 27'h00000338, 32'h00000400,
  1'd1,  5'd26, 27'h00000284, 5'd3, 27'h0000014d, 5'd1, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000290, 5'd1, 27'h000003e6, 5'd10, 27'h0000015a, 32'h00000400,
  1'd1,  5'd30, 27'h00000221, 5'd3, 27'h00000328, 5'd22, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000030, 5'd13, 27'h000001b1, 5'd4, 27'h000000fc, 32'h00000400,
  1'd1,  5'd26, 27'h00000064, 5'd10, 27'h000002ed, 5'd11, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001b3, 5'd14, 27'h00000177, 5'd24, 27'h0000036e, 32'h00000400,
  1'd1,  5'd26, 27'h000000d1, 5'd25, 27'h00000085, 5'd4, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e7, 5'd24, 27'h000000e1, 5'd13, 27'h000002a4, 32'h00000400,
  1'd1,  5'd30, 27'h000001a1, 5'd22, 27'h00000018, 5'd20, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000156, 5'd2, 27'h000000e7, 5'd4, 27'h000000a2, 32'h00000400,
  1'd1,  5'd5, 27'h00000254, 5'd1, 27'h00000031, 5'd14, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003c2, 5'd3, 27'h00000068, 5'd23, 27'h000002a7, 32'h00000400,
  1'd1,  5'd9, 27'h000000d0, 5'd14, 27'h00000066, 5'd10, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d1, 5'd10, 27'h00000275, 5'd16, 27'h0000025e, 32'h00000400,
  1'd1,  5'd10, 27'h000000bb, 5'd14, 27'h000003bd, 5'd29, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001eb, 5'd23, 27'h00000340, 5'd6, 27'h00000138, 32'h00000400,
  1'd1,  5'd7, 27'h000003d1, 5'd20, 27'h00000376, 5'd16, 27'h0000034f, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000110, 5'd21, 27'h0000011c, 5'd29, 27'h000000c8, 32'h00000400,
  1'd1,  5'd16, 27'h00000036, 5'd2, 27'h000002eb, 5'd0, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000196, 5'd3, 27'h000001eb, 5'd10, 27'h0000028c, 32'h00000400,
  1'd1,  5'd18, 27'h000001d7, 5'd3, 27'h00000370, 5'd20, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000103, 5'd13, 27'h00000054, 5'd8, 27'h000002ff, 32'h00000400,
  1'd1,  5'd17, 27'h00000043, 5'd11, 27'h0000038c, 5'd18, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000091, 5'd14, 27'h000001a4, 5'd27, 27'h0000022e, 32'h00000400,
  1'd1,  5'd17, 27'h0000025d, 5'd22, 27'h00000371, 5'd10, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000357, 5'd21, 27'h000001b9, 5'd17, 27'h0000037c, 32'h00000400,
  1'd1,  5'd19, 27'h0000009f, 5'd21, 27'h000000b6, 5'd29, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000060, 5'd4, 27'h00000337, 5'd10, 27'h00000014, 32'h00000400,
  1'd1,  5'd26, 27'h000000f1, 5'd2, 27'h0000020f, 5'd19, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000033a, 5'd0, 27'h0000016f, 5'd28, 27'h000001c2, 32'h00000400,
  1'd1,  5'd26, 27'h0000010f, 5'd13, 27'h0000016f, 5'd7, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000100, 5'd14, 27'h00000195, 5'd19, 27'h000000be, 32'h00000400,
  1'd1,  5'd30, 27'h0000039a, 5'd11, 27'h0000025a, 5'd29, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000137, 5'd23, 27'h000000b3, 5'd5, 27'h000001d4, 32'h00000400,
  1'd1,  5'd26, 27'h00000233, 5'd25, 27'h0000003c, 5'd20, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000021, 5'd20, 27'h00000330, 5'd26, 27'h000001b7, 32'h00000400,
  1'd1,  5'd10, 27'h00000035, 5'd9, 27'h00000285, 5'd2, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000024f, 5'd8, 27'h000002cf, 5'd11, 27'h00000334, 32'h00000400,
  1'd1,  5'd6, 27'h000000c7, 5'd5, 27'h0000036d, 5'd21, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003d7, 5'd20, 27'h0000026b, 5'd0, 27'h0000004d, 32'h00000400,
  1'd1,  5'd7, 27'h000002d3, 5'd17, 27'h0000007e, 5'd13, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000205, 5'd19, 27'h00000361, 5'd23, 27'h000001ab, 32'h00000400,
  1'd1,  5'd8, 27'h00000099, 5'd30, 27'h000002ef, 5'd2, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000050, 5'd29, 27'h000003fc, 5'd10, 27'h0000032a, 32'h00000400,
  1'd1,  5'd10, 27'h0000001c, 5'd26, 27'h00000017, 5'd25, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000047, 5'd5, 27'h000001e9, 5'd4, 27'h0000021e, 32'h00000400,
  1'd1,  5'd19, 27'h0000039b, 5'd7, 27'h0000033c, 5'd12, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000311, 5'd9, 27'h00000244, 5'd24, 27'h000002c2, 32'h00000400,
  1'd1,  5'd19, 27'h00000069, 5'd19, 27'h000002d1, 5'd2, 27'h000001c5, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a1, 5'd18, 27'h00000161, 5'd13, 27'h0000027b, 32'h00000400,
  1'd1,  5'd18, 27'h000003eb, 5'd15, 27'h00000343, 5'd21, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000177, 5'd26, 27'h00000303, 5'd1, 27'h000001d1, 32'h00000400,
  1'd1,  5'd16, 27'h000002b9, 5'd30, 27'h00000283, 5'd15, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002cc, 5'd29, 27'h00000291, 5'd21, 27'h000002d8, 32'h00000400,
  1'd1,  5'd27, 27'h00000370, 5'd9, 27'h000002cc, 5'd4, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001b5, 5'd8, 27'h000001f4, 5'd12, 27'h0000030b, 32'h00000400,
  1'd1,  5'd30, 27'h00000305, 5'd8, 27'h00000330, 5'd24, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000007b, 5'd17, 27'h000002df, 5'd0, 27'h00000152, 32'h00000400,
  1'd1,  5'd26, 27'h0000000a, 5'd15, 27'h000003e6, 5'd15, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000021b, 5'd18, 27'h00000010, 5'd23, 27'h000000f2, 32'h00000400,
  1'd1,  5'd28, 27'h00000251, 5'd29, 27'h0000012d, 5'd0, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000265, 5'd26, 27'h00000235, 5'd11, 27'h000003c3, 32'h00000400,
  1'd1,  5'd30, 27'h00000356, 5'd28, 27'h00000216, 5'd23, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000324, 5'd5, 27'h000003d4, 5'd7, 27'h000003a5, 32'h00000400,
  1'd1,  5'd5, 27'h000000dc, 5'd8, 27'h00000126, 5'd16, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002cf, 5'd5, 27'h00000301, 5'd30, 27'h00000132, 32'h00000400,
  1'd1,  5'd9, 27'h00000090, 5'd19, 27'h0000004a, 5'd8, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002db, 5'd17, 27'h00000173, 5'd17, 27'h00000274, 32'h00000400,
  1'd1,  5'd5, 27'h00000135, 5'd17, 27'h000002d2, 5'd26, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000009f, 5'd28, 27'h0000017a, 5'd7, 27'h000003af, 32'h00000400,
  1'd1,  5'd8, 27'h000000c8, 5'd26, 27'h0000022c, 5'd16, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000099, 5'd26, 27'h0000015d, 5'd26, 27'h00000375, 32'h00000400,
  1'd1,  5'd16, 27'h00000143, 5'd5, 27'h0000031f, 5'd7, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ea, 5'd9, 27'h0000001d, 5'd16, 27'h00000149, 32'h00000400,
  1'd1,  5'd19, 27'h000001bb, 5'd7, 27'h00000390, 5'd30, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000d6, 5'd18, 27'h00000385, 5'd6, 27'h00000061, 32'h00000400,
  1'd1,  5'd19, 27'h00000069, 5'd20, 27'h00000249, 5'd19, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b7, 5'd15, 27'h00000284, 5'd27, 27'h000002f6, 32'h00000400,
  1'd1,  5'd16, 27'h00000293, 5'd30, 27'h000000a0, 5'd6, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b8, 5'd26, 27'h000000e6, 5'd17, 27'h0000010b, 32'h00000400,
  1'd1,  5'd19, 27'h000000c8, 5'd30, 27'h0000016f, 5'd30, 27'h00000214, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000234, 5'd5, 27'h00000182, 5'd5, 27'h000001e5, 32'h00000400,
  1'd1,  5'd27, 27'h000001c0, 5'd7, 27'h0000003e, 5'd17, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000f9, 5'd8, 27'h000002fd, 5'd30, 27'h000000ef, 32'h00000400,
  1'd1,  5'd30, 27'h00000129, 5'd18, 27'h0000020a, 5'd10, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000d8, 5'd18, 27'h000001df, 5'd20, 27'h000000c4, 32'h00000400,
  1'd1,  5'd26, 27'h000003c7, 5'd20, 27'h0000011b, 5'd25, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000018c, 5'd26, 27'h000000ef, 5'd10, 27'h00000009, 32'h00000400,
  1'd1,  5'd28, 27'h00000010, 5'd30, 27'h000000ab, 5'd20, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001ff, 5'd30, 27'h00000004, 5'd29, 27'h00000326, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h0000003f, 5'd2, 27'h00000347, 5'd3, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000b3, 5'd1, 27'h00000077, 5'd12, 27'h00000040, 32'h00000400,
  1'd1,  5'd1, 27'h000003a5, 5'd1, 27'h000003c4, 5'd22, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a5, 5'd13, 27'h000000c4, 5'd0, 27'h000001fe, 32'h00000400,
  1'd1,  5'd5, 27'h00000092, 5'd15, 27'h0000005d, 5'd13, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f6, 5'd14, 27'h00000254, 5'd24, 27'h00000067, 32'h00000400,
  1'd1,  5'd1, 27'h0000023d, 5'd24, 27'h00000172, 5'd4, 27'h00000011, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000315, 5'd24, 27'h000002cd, 5'd14, 27'h000002ce, 32'h00000400,
  1'd1,  5'd2, 27'h00000168, 5'd25, 27'h00000095, 5'd20, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000156, 5'd0, 27'h0000016c, 5'd2, 27'h00000263, 32'h00000400,
  1'd1,  5'd15, 27'h00000061, 5'd2, 27'h00000351, 5'd11, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000171, 5'd3, 27'h000002c6, 5'd24, 27'h000000eb, 32'h00000400,
  1'd1,  5'd13, 27'h0000028a, 5'd13, 27'h00000296, 5'd1, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000180, 5'd13, 27'h0000031a, 5'd11, 27'h000000ab, 32'h00000400,
  1'd1,  5'd11, 27'h000000fd, 5'd11, 27'h000001e0, 5'd24, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000037f, 5'd22, 27'h00000253, 5'd0, 27'h00000173, 32'h00000400,
  1'd1,  5'd10, 27'h0000022a, 5'd23, 27'h00000386, 5'd12, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000cb, 5'd22, 27'h000000ad, 5'd21, 27'h0000036c, 32'h00000400,
  1'd1,  5'd24, 27'h00000195, 5'd2, 27'h000003e5, 5'd0, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000143, 5'd4, 27'h000001ea, 5'd11, 27'h000000a0, 32'h00000400,
  1'd1,  5'd21, 27'h000003c0, 5'd1, 27'h000002fe, 5'd23, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000363, 5'd11, 27'h000003ae, 5'd0, 27'h00000039, 32'h00000400,
  1'd1,  5'd24, 27'h000002f9, 5'd13, 27'h0000034a, 5'd14, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000c9, 5'd10, 27'h00000340, 5'd24, 27'h00000166, 32'h00000400,
  1'd1,  5'd23, 27'h0000008a, 5'd25, 27'h00000298, 5'd3, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001d4, 5'd25, 27'h0000019a, 5'd12, 27'h0000019f, 32'h00000400,
  1'd1,  5'd24, 27'h00000036, 5'd22, 27'h00000247, 5'd25, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002f3, 5'd4, 27'h0000010a, 5'd6, 27'h000000d2, 32'h00000400,
  1'd1,  5'd2, 27'h0000038e, 5'd5, 27'h0000005a, 5'd15, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000d7, 5'd4, 27'h000001cc, 5'd29, 27'h0000038d, 32'h00000400,
  1'd1,  5'd5, 27'h00000017, 5'd12, 27'h0000038d, 5'd6, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003cf, 5'd13, 27'h000001d5, 5'd20, 27'h00000278, 32'h00000400,
  1'd1,  5'd3, 27'h000000a7, 5'd12, 27'h00000046, 5'd27, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003f8, 5'd20, 27'h000002e6, 5'd5, 27'h000002a7, 32'h00000400,
  1'd1,  5'd0, 27'h0000014f, 5'd25, 27'h0000033c, 5'd19, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036a, 5'd23, 27'h000003c1, 5'd28, 27'h000000b1, 32'h00000400,
  1'd1,  5'd14, 27'h0000039b, 5'd4, 27'h00000169, 5'd6, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002d1, 5'd2, 27'h0000017a, 5'd17, 27'h00000011, 32'h00000400,
  1'd1,  5'd10, 27'h00000173, 5'd3, 27'h00000154, 5'd30, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b6, 5'd11, 27'h0000020e, 5'd6, 27'h00000379, 32'h00000400,
  1'd1,  5'd13, 27'h0000032e, 5'd10, 27'h0000031c, 5'd18, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000048, 5'd12, 27'h000000c8, 5'd26, 27'h00000370, 32'h00000400,
  1'd1,  5'd12, 27'h000001d6, 5'd24, 27'h000000c3, 5'd8, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000e6, 5'd24, 27'h0000038b, 5'd19, 27'h000002eb, 32'h00000400,
  1'd1,  5'd13, 27'h00000253, 5'd23, 27'h000001ea, 5'd29, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000312, 5'd3, 27'h00000011, 5'd8, 27'h00000375, 32'h00000400,
  1'd1,  5'd22, 27'h000003dc, 5'd1, 27'h00000070, 5'd20, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000058, 5'd0, 27'h0000003a, 5'd27, 27'h00000164, 32'h00000400,
  1'd1,  5'd21, 27'h00000050, 5'd13, 27'h00000211, 5'd9, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000023, 5'd12, 27'h000003e9, 5'd15, 27'h000003bd, 32'h00000400,
  1'd1,  5'd21, 27'h000001de, 5'd13, 27'h000002c3, 5'd29, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000383, 5'd25, 27'h0000034e, 5'd8, 27'h0000037f, 32'h00000400,
  1'd1,  5'd24, 27'h000003cd, 5'd25, 27'h0000007b, 5'd15, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000005f, 5'd21, 27'h00000320, 5'd30, 27'h00000214, 32'h00000400,
  1'd1,  5'd4, 27'h0000003c, 5'd9, 27'h00000240, 5'd4, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000335, 5'd7, 27'h00000181, 5'd12, 27'h00000070, 32'h00000400,
  1'd1,  5'd0, 27'h0000012f, 5'd9, 27'h0000036e, 5'd25, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000023c, 5'd18, 27'h000000d5, 5'd3, 27'h000000f3, 32'h00000400,
  1'd1,  5'd3, 27'h0000036e, 5'd18, 27'h00000345, 5'd10, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000099, 5'd15, 27'h000003a1, 5'd25, 27'h00000303, 32'h00000400,
  1'd1,  5'd2, 27'h000000ca, 5'd26, 27'h000002da, 5'd1, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ce, 5'd27, 27'h0000017c, 5'd14, 27'h000000ea, 32'h00000400,
  1'd1,  5'd1, 27'h000002de, 5'd27, 27'h000003be, 5'd22, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000019c, 5'd5, 27'h0000035d, 5'd2, 27'h000000df, 32'h00000400,
  1'd1,  5'd11, 27'h00000056, 5'd7, 27'h000001be, 5'd12, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e5, 5'd10, 27'h0000005f, 5'd23, 27'h0000018c, 32'h00000400,
  1'd1,  5'd14, 27'h000000ec, 5'd17, 27'h00000191, 5'd2, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003aa, 5'd20, 27'h000001ea, 5'd10, 27'h0000030d, 32'h00000400,
  1'd1,  5'd13, 27'h00000396, 5'd20, 27'h000001c1, 5'd25, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000fc, 5'd26, 27'h000003a0, 5'd2, 27'h000001c4, 32'h00000400,
  1'd1,  5'd11, 27'h0000025c, 5'd28, 27'h000003d9, 5'd10, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000038b, 5'd29, 27'h000000da, 5'd22, 27'h0000000a, 32'h00000400,
  1'd1,  5'd24, 27'h000000b8, 5'd6, 27'h0000031a, 5'd2, 27'h00000094, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000018a, 5'd9, 27'h000001d4, 5'd10, 27'h0000017d, 32'h00000400,
  1'd1,  5'd24, 27'h00000217, 5'd6, 27'h0000029d, 5'd25, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000013b, 5'd20, 27'h000000b4, 5'd1, 27'h000000b7, 32'h00000400,
  1'd1,  5'd23, 27'h00000047, 5'd16, 27'h000002a9, 5'd10, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000011, 5'd20, 27'h000001d7, 5'd21, 27'h00000140, 32'h00000400,
  1'd1,  5'd22, 27'h000001d2, 5'd27, 27'h0000004b, 5'd4, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001b0, 5'd27, 27'h00000372, 5'd15, 27'h0000001b, 32'h00000400,
  1'd1,  5'd23, 27'h00000316, 5'd27, 27'h00000364, 5'd23, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000010a, 5'd8, 27'h0000032a, 5'd7, 27'h00000188, 32'h00000400,
  1'd1,  5'd1, 27'h00000162, 5'd7, 27'h000002fa, 5'd19, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d8, 5'd6, 27'h000002b8, 5'd28, 27'h00000213, 32'h00000400,
  1'd1,  5'd1, 27'h000000ae, 5'd19, 27'h00000356, 5'd8, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003c0, 5'd19, 27'h00000126, 5'd20, 27'h00000046, 32'h00000400,
  1'd1,  5'd1, 27'h00000256, 5'd17, 27'h000003a9, 5'd28, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000228, 5'd27, 27'h0000023d, 5'd9, 27'h00000143, 32'h00000400,
  1'd1,  5'd5, 27'h00000050, 5'd30, 27'h000001e2, 5'd20, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000d0, 5'd27, 27'h0000039b, 5'd29, 27'h000001fc, 32'h00000400,
  1'd1,  5'd15, 27'h0000004b, 5'd7, 27'h000002f8, 5'd6, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000013c, 5'd6, 27'h000000d3, 5'd19, 27'h00000165, 32'h00000400,
  1'd1,  5'd13, 27'h00000231, 5'd5, 27'h00000210, 5'd30, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000ec, 5'd18, 27'h0000039e, 5'd6, 27'h00000230, 32'h00000400,
  1'd1,  5'd13, 27'h00000052, 5'd18, 27'h000003b2, 5'd20, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000054, 5'd17, 27'h000001f8, 5'd28, 27'h000002ae, 32'h00000400,
  1'd1,  5'd10, 27'h000001f6, 5'd29, 27'h000001eb, 5'd5, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000178, 5'd28, 27'h000002d9, 5'd18, 27'h0000022f, 32'h00000400,
  1'd1,  5'd15, 27'h00000008, 5'd30, 27'h000001d3, 5'd27, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002d5, 5'd7, 27'h00000060, 5'd6, 27'h00000274, 32'h00000400,
  1'd1,  5'd23, 27'h00000380, 5'd9, 27'h00000192, 5'd17, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002af, 5'd6, 27'h000001c4, 5'd27, 27'h000001be, 32'h00000400,
  1'd1,  5'd25, 27'h000000bb, 5'd18, 27'h00000142, 5'd5, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000123, 5'd18, 27'h000003f6, 5'd15, 27'h000002e5, 32'h00000400,
  1'd1,  5'd23, 27'h000002ef, 5'd18, 27'h00000104, 5'd27, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000097, 5'd26, 27'h0000035a, 5'd7, 27'h000002e4, 32'h00000400,
  1'd1,  5'd24, 27'h000003c4, 5'd28, 27'h00000316, 5'd20, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000355, 5'd26, 27'h00000194, 5'd27, 27'h00000115, 32'h00000400,
  1'd1,  5'd6, 27'h0000034b, 5'd2, 27'h000001c0, 5'd8, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a5, 5'd0, 27'h000000d4, 5'd19, 27'h00000287, 32'h00000400,
  1'd1,  5'd10, 27'h000000dc, 5'd1, 27'h000001b2, 5'd28, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000172, 5'd15, 27'h0000017f, 5'd1, 27'h00000230, 32'h00000400,
  1'd1,  5'd6, 27'h000003c1, 5'd14, 27'h00000346, 5'd10, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000003f, 5'd11, 27'h00000102, 5'd21, 27'h00000283, 32'h00000400,
  1'd1,  5'd5, 27'h0000011c, 5'd21, 27'h000002d3, 5'd2, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000006d, 5'd20, 27'h000003b8, 5'd13, 27'h0000036c, 32'h00000400,
  1'd1,  5'd5, 27'h000001b9, 5'd22, 27'h0000020d, 5'd24, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032a, 5'd3, 27'h000000c8, 5'd5, 27'h00000168, 32'h00000400,
  1'd1,  5'd17, 27'h00000369, 5'd0, 27'h0000008b, 5'd16, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001cc, 5'd4, 27'h0000011f, 5'd29, 27'h0000007a, 32'h00000400,
  1'd1,  5'd15, 27'h00000295, 5'd12, 27'h000001cf, 5'd0, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000015f, 5'd15, 27'h00000102, 5'd11, 27'h000001e5, 32'h00000400,
  1'd1,  5'd20, 27'h00000164, 5'd10, 27'h000002ca, 5'd22, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000003a, 5'd25, 27'h000001a6, 5'd0, 27'h00000271, 32'h00000400,
  1'd1,  5'd19, 27'h0000037f, 5'd22, 27'h00000310, 5'd12, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000389, 5'd21, 27'h000000cc, 5'd22, 27'h0000026c, 32'h00000400,
  1'd1,  5'd25, 27'h0000038a, 5'd4, 27'h000003e7, 5'd1, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000e, 5'd2, 27'h0000011a, 5'd13, 27'h00000017, 32'h00000400,
  1'd1,  5'd28, 27'h00000351, 5'd1, 27'h0000002d, 5'd21, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000039c, 5'd11, 27'h000003bc, 5'd3, 27'h000003b7, 32'h00000400,
  1'd1,  5'd26, 27'h00000273, 5'd15, 27'h0000019c, 5'd12, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c7, 5'd11, 27'h00000055, 5'd22, 27'h000003b4, 32'h00000400,
  1'd1,  5'd26, 27'h0000009c, 5'd22, 27'h00000019, 5'd0, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000321, 5'd23, 27'h00000091, 5'd11, 27'h000000c1, 32'h00000400,
  1'd1,  5'd28, 27'h00000174, 5'd25, 27'h00000247, 5'd25, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023d, 5'd1, 27'h00000213, 5'd3, 27'h00000210, 32'h00000400,
  1'd1,  5'd9, 27'h000001f9, 5'd5, 27'h00000086, 5'd11, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000262, 5'd3, 27'h000000ba, 5'd25, 27'h0000007b, 32'h00000400,
  1'd1,  5'd10, 27'h000000d2, 5'd10, 27'h000001f1, 5'd8, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000035d, 5'd11, 27'h000001d5, 5'd20, 27'h00000272, 32'h00000400,
  1'd1,  5'd7, 27'h000000c5, 5'd14, 27'h00000101, 5'd27, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000012, 5'd24, 27'h0000016a, 5'd6, 27'h00000363, 32'h00000400,
  1'd1,  5'd7, 27'h00000055, 5'd22, 27'h00000138, 5'd17, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003d9, 5'd23, 27'h000003b7, 5'd26, 27'h000000aa, 32'h00000400,
  1'd1,  5'd17, 27'h000003cf, 5'd1, 27'h00000381, 5'd2, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002ff, 5'd4, 27'h000002b2, 5'd12, 27'h000003f9, 32'h00000400,
  1'd1,  5'd17, 27'h000000bc, 5'd1, 27'h00000071, 5'd23, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000265, 5'd15, 27'h00000074, 5'd6, 27'h0000014b, 32'h00000400,
  1'd1,  5'd17, 27'h0000002b, 5'd13, 27'h00000219, 5'd18, 27'h0000010b, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002b5, 5'd15, 27'h00000074, 5'd28, 27'h0000026d, 32'h00000400,
  1'd1,  5'd17, 27'h0000003a, 5'd25, 27'h0000025c, 5'd10, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000395, 5'd23, 27'h000002b4, 5'd19, 27'h000001ea, 32'h00000400,
  1'd1,  5'd17, 27'h000003c0, 5'd23, 27'h000000e8, 5'd30, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000d4, 5'd3, 27'h0000004c, 5'd5, 27'h00000399, 32'h00000400,
  1'd1,  5'd28, 27'h0000006b, 5'd5, 27'h0000005d, 5'd16, 27'h0000036c, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000183, 5'd2, 27'h000003c5, 5'd28, 27'h0000011c, 32'h00000400,
  1'd1,  5'd28, 27'h0000008a, 5'd14, 27'h00000356, 5'd7, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002c2, 5'd13, 27'h000003b5, 5'd20, 27'h0000004a, 32'h00000400,
  1'd1,  5'd28, 27'h00000360, 5'd13, 27'h00000011, 5'd27, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001f9, 5'd22, 27'h00000152, 5'd9, 27'h000001e3, 32'h00000400,
  1'd1,  5'd26, 27'h0000030d, 5'd20, 27'h000002ca, 5'd18, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000002c, 5'd24, 27'h000002b4, 5'd25, 27'h000003da, 32'h00000400,
  1'd1,  5'd8, 27'h00000108, 5'd8, 27'h00000122, 5'd3, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002ed, 5'd8, 27'h00000335, 5'd12, 27'h00000179, 32'h00000400,
  1'd1,  5'd6, 27'h00000193, 5'd8, 27'h00000346, 5'd23, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000023a, 5'd16, 27'h000001aa, 5'd3, 27'h0000019c, 32'h00000400,
  1'd1,  5'd5, 27'h00000311, 5'd17, 27'h00000363, 5'd13, 27'h00000055, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a1, 5'd18, 27'h000001e8, 5'd21, 27'h00000167, 32'h00000400,
  1'd1,  5'd8, 27'h00000242, 5'd27, 27'h000003c9, 5'd4, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000002f, 5'd27, 27'h000002b3, 5'd14, 27'h000001bf, 32'h00000400,
  1'd1,  5'd9, 27'h0000002d, 5'd28, 27'h000002ab, 5'd21, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000004b, 5'd6, 27'h000003a5, 5'd4, 27'h00000137, 32'h00000400,
  1'd1,  5'd18, 27'h00000389, 5'd7, 27'h0000004c, 5'd13, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002a2, 5'd10, 27'h00000029, 5'd20, 27'h00000366, 32'h00000400,
  1'd1,  5'd19, 27'h00000045, 5'd18, 27'h0000034a, 5'd5, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000020e, 5'd16, 27'h000003f9, 5'd14, 27'h000001c9, 32'h00000400,
  1'd1,  5'd15, 27'h000003d5, 5'd20, 27'h00000172, 5'd22, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000301, 5'd27, 27'h00000064, 5'd2, 27'h000001d2, 32'h00000400,
  1'd1,  5'd20, 27'h0000017a, 5'd28, 27'h0000002b, 5'd13, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000a6, 5'd29, 27'h0000027d, 5'd25, 27'h0000016a, 32'h00000400,
  1'd1,  5'd28, 27'h000002c0, 5'd5, 27'h00000324, 5'd3, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001f6, 5'd5, 27'h000002c9, 5'd11, 27'h0000021f, 32'h00000400,
  1'd1,  5'd26, 27'h000003d6, 5'd5, 27'h000001c4, 5'd22, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002ce, 5'd19, 27'h00000193, 5'd4, 27'h0000037b, 32'h00000400,
  1'd1,  5'd28, 27'h00000026, 5'd20, 27'h000000ae, 5'd14, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000213, 5'd18, 27'h0000009b, 5'd22, 27'h00000207, 32'h00000400,
  1'd1,  5'd27, 27'h0000021f, 5'd27, 27'h00000292, 5'd2, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003e6, 5'd30, 27'h00000361, 5'd12, 27'h00000259, 32'h00000400,
  1'd1,  5'd27, 27'h000003ae, 5'd26, 27'h00000242, 5'd21, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000170, 5'd6, 27'h000002fd, 5'd9, 27'h00000044, 32'h00000400,
  1'd1,  5'd5, 27'h00000383, 5'd6, 27'h0000021f, 5'd18, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003b4, 5'd7, 27'h000001ec, 5'd30, 27'h00000285, 32'h00000400,
  1'd1,  5'd5, 27'h0000028a, 5'd19, 27'h00000139, 5'd8, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000255, 5'd15, 27'h000003a8, 5'd18, 27'h00000188, 32'h00000400,
  1'd1,  5'd8, 27'h000001a8, 5'd19, 27'h00000017, 5'd27, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a0, 5'd30, 27'h00000270, 5'd8, 27'h000000ad, 32'h00000400,
  1'd1,  5'd5, 27'h00000343, 5'd27, 27'h00000046, 5'd16, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000259, 5'd26, 27'h000003ba, 5'd27, 27'h00000100, 32'h00000400,
  1'd1,  5'd16, 27'h000002ed, 5'd5, 27'h00000277, 5'd8, 27'h000000d2, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000b7, 5'd5, 27'h000001d9, 5'd16, 27'h000001e6, 32'h00000400,
  1'd1,  5'd15, 27'h000003f9, 5'd7, 27'h000001ce, 5'd27, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000277, 5'd18, 27'h0000038b, 5'd8, 27'h00000069, 32'h00000400,
  1'd1,  5'd18, 27'h00000268, 5'd15, 27'h00000262, 5'd20, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a2, 5'd17, 27'h00000294, 5'd29, 27'h0000039b, 32'h00000400,
  1'd1,  5'd16, 27'h0000027d, 5'd27, 27'h00000025, 5'd7, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000030d, 5'd29, 27'h000000c9, 5'd16, 27'h000000a8, 32'h00000400,
  1'd1,  5'd20, 27'h000000d9, 5'd28, 27'h0000019c, 5'd30, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002fd, 5'd7, 27'h00000281, 5'd5, 27'h000001f0, 32'h00000400,
  1'd1,  5'd30, 27'h0000013a, 5'd10, 27'h000000ef, 5'd20, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000dc, 5'd7, 27'h0000001e, 5'd27, 27'h000001cc, 32'h00000400,
  1'd1,  5'd30, 27'h00000293, 5'd19, 27'h00000082, 5'd9, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b8, 5'd19, 27'h000002c1, 5'd16, 27'h00000229, 32'h00000400,
  1'd1,  5'd26, 27'h00000352, 5'd19, 27'h00000210, 5'd25, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000243, 5'd29, 27'h0000002b, 5'd9, 27'h000001f5, 32'h00000400,
  1'd1,  5'd28, 27'h000003db, 5'd28, 27'h00000262, 5'd17, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f1, 5'd27, 27'h00000373, 5'd30, 27'h00000116, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h0000034e, 5'd1, 27'h00000376, 5'd1, 27'h00000349, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000030d, 5'd2, 27'h0000006f, 5'd15, 27'h00000195, 32'h00000400,
  1'd1,  5'd3, 27'h00000350, 5'd0, 27'h00000166, 5'd24, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000065, 5'd12, 27'h0000027a, 5'd3, 27'h00000364, 32'h00000400,
  1'd1,  5'd0, 27'h00000351, 5'd14, 27'h0000000e, 5'd12, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020f, 5'd13, 27'h000002b1, 5'd24, 27'h00000363, 32'h00000400,
  1'd1,  5'd2, 27'h0000005a, 5'd25, 27'h00000025, 5'd4, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003df, 5'd22, 27'h0000010e, 5'd14, 27'h000002a6, 32'h00000400,
  1'd1,  5'd3, 27'h00000199, 5'd22, 27'h0000028b, 5'd20, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f2, 5'd1, 27'h000003f5, 5'd3, 27'h00000380, 32'h00000400,
  1'd1,  5'd15, 27'h000000ee, 5'd2, 27'h00000331, 5'd14, 27'h000003bd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e3, 5'd4, 27'h0000028c, 5'd21, 27'h0000009d, 32'h00000400,
  1'd1,  5'd11, 27'h00000045, 5'd10, 27'h000003c0, 5'd1, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002bf, 5'd11, 27'h00000206, 5'd10, 27'h0000025a, 32'h00000400,
  1'd1,  5'd12, 27'h000001d4, 5'd15, 27'h00000107, 5'd22, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e2, 5'd24, 27'h0000033e, 5'd1, 27'h000001e6, 32'h00000400,
  1'd1,  5'd11, 27'h000000a6, 5'd23, 27'h00000026, 5'd13, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ae, 5'd22, 27'h00000284, 5'd22, 27'h00000101, 32'h00000400,
  1'd1,  5'd25, 27'h0000013e, 5'd1, 27'h000003d4, 5'd2, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000089, 5'd2, 27'h00000050, 5'd12, 27'h000000ab, 32'h00000400,
  1'd1,  5'd24, 27'h00000395, 5'd4, 27'h00000054, 5'd23, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f0, 5'd14, 27'h000003ae, 5'd0, 27'h000003b1, 32'h00000400,
  1'd1,  5'd23, 27'h000001f3, 5'd13, 27'h0000034c, 5'd10, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021a, 5'd10, 27'h000003cc, 5'd21, 27'h000003a2, 32'h00000400,
  1'd1,  5'd23, 27'h000001a3, 5'd22, 27'h0000012c, 5'd4, 27'h00000210, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000237, 5'd21, 27'h000001c6, 5'd12, 27'h00000282, 32'h00000400,
  1'd1,  5'd22, 27'h000003e8, 5'd22, 27'h00000145, 5'd22, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a3, 5'd4, 27'h000000c6, 5'd8, 27'h0000010f, 32'h00000400,
  1'd1,  5'd4, 27'h000001cf, 5'd5, 27'h0000001e, 5'd16, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000079, 5'd2, 27'h00000294, 5'd26, 27'h00000387, 32'h00000400,
  1'd1,  5'd4, 27'h000003f9, 5'd14, 27'h00000033, 5'd9, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000314, 5'd12, 27'h00000239, 5'd19, 27'h0000037a, 32'h00000400,
  1'd1,  5'd4, 27'h00000298, 5'd14, 27'h000002b6, 5'd26, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002f7, 5'd20, 27'h0000038e, 5'd9, 27'h0000020a, 32'h00000400,
  1'd1,  5'd0, 27'h000002aa, 5'd25, 27'h00000048, 5'd19, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002f3, 5'd21, 27'h0000030c, 5'd27, 27'h0000030a, 32'h00000400,
  1'd1,  5'd12, 27'h0000039f, 5'd4, 27'h00000230, 5'd6, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000173, 5'd1, 27'h000002ea, 5'd16, 27'h0000025c, 32'h00000400,
  1'd1,  5'd15, 27'h0000010f, 5'd3, 27'h000002ce, 5'd29, 27'h00000311, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000006f, 5'd13, 27'h00000189, 5'd8, 27'h0000033e, 32'h00000400,
  1'd1,  5'd14, 27'h00000059, 5'd13, 27'h000000ae, 5'd17, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000022c, 5'd10, 27'h00000391, 5'd28, 27'h00000114, 32'h00000400,
  1'd1,  5'd11, 27'h00000199, 5'd23, 27'h00000140, 5'd9, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000076, 5'd24, 27'h000000ae, 5'd20, 27'h000001cc, 32'h00000400,
  1'd1,  5'd15, 27'h00000083, 5'd21, 27'h00000165, 5'd30, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000012, 5'd2, 27'h0000000c, 5'd6, 27'h000002d2, 32'h00000400,
  1'd1,  5'd22, 27'h0000001b, 5'd3, 27'h00000283, 5'd19, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000064, 5'd5, 27'h00000080, 5'd30, 27'h000000fd, 32'h00000400,
  1'd1,  5'd24, 27'h000003d5, 5'd14, 27'h00000254, 5'd5, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000107, 5'd11, 27'h00000323, 5'd17, 27'h000000a2, 32'h00000400,
  1'd1,  5'd24, 27'h00000301, 5'd11, 27'h00000283, 5'd27, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001c6, 5'd25, 27'h000001a7, 5'd7, 27'h00000117, 32'h00000400,
  1'd1,  5'd23, 27'h000000e3, 5'd25, 27'h00000204, 5'd18, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000030f, 5'd22, 27'h00000333, 5'd27, 27'h00000007, 32'h00000400,
  1'd1,  5'd1, 27'h000000d2, 5'd8, 27'h00000087, 5'd5, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000179, 5'd9, 27'h000001bf, 5'd15, 27'h0000007a, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd9, 27'h00000141, 5'd24, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000389, 5'd15, 27'h0000031a, 5'd2, 27'h000001db, 32'h00000400,
  1'd1,  5'd4, 27'h00000049, 5'd17, 27'h00000068, 5'd11, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000256, 5'd16, 27'h00000103, 5'd24, 27'h0000019c, 32'h00000400,
  1'd1,  5'd4, 27'h000002d3, 5'd25, 27'h0000036f, 5'd3, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000035c, 5'd28, 27'h00000071, 5'd11, 27'h0000036a, 32'h00000400,
  1'd1,  5'd1, 27'h00000145, 5'd25, 27'h0000035c, 5'd20, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c7, 5'd9, 27'h00000197, 5'd0, 27'h00000016, 32'h00000400,
  1'd1,  5'd11, 27'h000001a6, 5'd7, 27'h0000006a, 5'd11, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d5, 5'd8, 27'h000000cd, 5'd21, 27'h00000179, 32'h00000400,
  1'd1,  5'd12, 27'h0000012d, 5'd17, 27'h00000002, 5'd0, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000015b, 5'd20, 27'h0000014a, 5'd12, 27'h00000358, 32'h00000400,
  1'd1,  5'd14, 27'h00000049, 5'd16, 27'h0000023e, 5'd23, 27'h000000c3, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000034d, 5'd26, 27'h000000ae, 5'd2, 27'h00000334, 32'h00000400,
  1'd1,  5'd10, 27'h00000320, 5'd26, 27'h00000167, 5'd14, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023c, 5'd26, 27'h00000114, 5'd25, 27'h00000234, 32'h00000400,
  1'd1,  5'd25, 27'h00000280, 5'd9, 27'h00000288, 5'd2, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003fc, 5'd6, 27'h000002df, 5'd11, 27'h0000004e, 32'h00000400,
  1'd1,  5'd21, 27'h00000016, 5'd6, 27'h0000015b, 5'd24, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d5, 5'd19, 27'h00000289, 5'd2, 27'h0000027e, 32'h00000400,
  1'd1,  5'd23, 27'h000001d1, 5'd17, 27'h00000214, 5'd11, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000046, 5'd19, 27'h000001dc, 5'd21, 27'h00000194, 32'h00000400,
  1'd1,  5'd25, 27'h00000025, 5'd26, 27'h00000157, 5'd0, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000358, 5'd28, 27'h000002c1, 5'd15, 27'h00000160, 32'h00000400,
  1'd1,  5'd21, 27'h00000233, 5'd30, 27'h00000048, 5'd23, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d9, 5'd8, 27'h00000322, 5'd5, 27'h00000244, 32'h00000400,
  1'd1,  5'd0, 27'h000003bb, 5'd5, 27'h00000262, 5'd19, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000006d, 5'd8, 27'h000000e8, 5'd29, 27'h0000000b, 32'h00000400,
  1'd1,  5'd0, 27'h000002cd, 5'd19, 27'h0000028c, 5'd9, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001a7, 5'd18, 27'h0000002f, 5'd15, 27'h00000321, 32'h00000400,
  1'd1,  5'd5, 27'h00000029, 5'd18, 27'h000000fc, 5'd27, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000002, 5'd30, 27'h000000fb, 5'd8, 27'h0000009f, 32'h00000400,
  1'd1,  5'd3, 27'h000002e2, 5'd26, 27'h000001c1, 5'd19, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000002, 5'd30, 27'h000001d0, 5'd27, 27'h0000021b, 32'h00000400,
  1'd1,  5'd13, 27'h000003c2, 5'd7, 27'h0000037c, 5'd6, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000344, 5'd6, 27'h00000312, 5'd18, 27'h00000364, 32'h00000400,
  1'd1,  5'd14, 27'h00000133, 5'd8, 27'h0000007a, 5'd26, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000b6, 5'd17, 27'h00000002, 5'd7, 27'h00000105, 32'h00000400,
  1'd1,  5'd15, 27'h00000023, 5'd16, 27'h0000012e, 5'd18, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d1, 5'd18, 27'h000001f1, 5'd30, 27'h000001db, 32'h00000400,
  1'd1,  5'd13, 27'h000002b7, 5'd30, 27'h0000023e, 5'd8, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001fa, 5'd26, 27'h00000049, 5'd20, 27'h0000015e, 32'h00000400,
  1'd1,  5'd14, 27'h0000027b, 5'd29, 27'h000001f9, 5'd30, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001ca, 5'd5, 27'h000003a5, 5'd9, 27'h000000e5, 32'h00000400,
  1'd1,  5'd25, 27'h0000026a, 5'd9, 27'h00000167, 5'd18, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000166, 5'd5, 27'h000001bc, 5'd27, 27'h0000032b, 32'h00000400,
  1'd1,  5'd25, 27'h00000003, 5'd17, 27'h0000034b, 5'd8, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c3, 5'd17, 27'h00000062, 5'd19, 27'h000002a0, 32'h00000400,
  1'd1,  5'd24, 27'h0000011a, 5'd17, 27'h000002b8, 5'd25, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032e, 5'd28, 27'h0000037a, 5'd8, 27'h00000370, 32'h00000400,
  1'd1,  5'd21, 27'h000000a3, 5'd26, 27'h00000311, 5'd17, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000036d, 5'd29, 27'h000002d2, 5'd28, 27'h00000303, 32'h00000400,
  1'd1,  5'd9, 27'h0000005e, 5'd0, 27'h000002a9, 5'd7, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038d, 5'd1, 27'h000000be, 5'd20, 27'h0000014d, 32'h00000400,
  1'd1,  5'd6, 27'h00000367, 5'd3, 27'h000003ec, 5'd28, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000002b, 5'd11, 27'h0000026c, 5'd5, 27'h00000099, 32'h00000400,
  1'd1,  5'd9, 27'h000002ab, 5'd15, 27'h000001ad, 5'd10, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002e8, 5'd11, 27'h00000096, 5'd24, 27'h00000071, 32'h00000400,
  1'd1,  5'd5, 27'h000001b4, 5'd22, 27'h000000bf, 5'd2, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002bc, 5'd21, 27'h00000312, 5'd11, 27'h00000263, 32'h00000400,
  1'd1,  5'd5, 27'h00000295, 5'd23, 27'h000001e4, 5'd20, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000006, 5'd0, 27'h00000209, 5'd5, 27'h00000155, 32'h00000400,
  1'd1,  5'd19, 27'h000003df, 5'd4, 27'h0000005a, 5'd16, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000036e, 5'd1, 27'h000000e6, 5'd26, 27'h0000026e, 32'h00000400,
  1'd1,  5'd17, 27'h00000090, 5'd14, 27'h0000003b, 5'd0, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000137, 5'd13, 27'h0000009a, 5'd14, 27'h000000cb, 32'h00000400,
  1'd1,  5'd20, 27'h00000132, 5'd13, 27'h00000122, 5'd21, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000235, 5'd20, 27'h000003de, 5'd1, 27'h000001bd, 32'h00000400,
  1'd1,  5'd20, 27'h0000001e, 5'd23, 27'h0000036c, 5'd10, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000016e, 5'd22, 27'h0000034d, 5'd21, 27'h0000035c, 32'h00000400,
  1'd1,  5'd27, 27'h0000021b, 5'd1, 27'h00000109, 5'd3, 27'h0000030c, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000190, 5'd4, 27'h0000011c, 5'd13, 27'h000002ae, 32'h00000400,
  1'd1,  5'd30, 27'h0000011e, 5'd3, 27'h0000018b, 5'd23, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000017c, 5'd12, 27'h000002ca, 5'd1, 27'h000003e9, 32'h00000400,
  1'd1,  5'd27, 27'h000002df, 5'd14, 27'h000002e4, 5'd12, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002d2, 5'd13, 27'h00000338, 5'd25, 27'h00000331, 32'h00000400,
  1'd1,  5'd27, 27'h000001d3, 5'd20, 27'h000002d9, 5'd0, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000010, 5'd24, 27'h000000d5, 5'd12, 27'h000001d9, 32'h00000400,
  1'd1,  5'd29, 27'h0000001a, 5'd25, 27'h00000211, 5'd22, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003e0, 5'd1, 27'h00000017, 5'd4, 27'h00000199, 32'h00000400,
  1'd1,  5'd9, 27'h00000068, 5'd4, 27'h00000242, 5'd14, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000039b, 5'd1, 27'h000003b0, 5'd23, 27'h0000007c, 32'h00000400,
  1'd1,  5'd8, 27'h000003a2, 5'd11, 27'h00000331, 5'd7, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a2, 5'd11, 27'h000002e4, 5'd19, 27'h00000333, 32'h00000400,
  1'd1,  5'd6, 27'h00000343, 5'd12, 27'h0000021d, 5'd30, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000078, 5'd25, 27'h000001db, 5'd8, 27'h00000308, 32'h00000400,
  1'd1,  5'd9, 27'h000002c7, 5'd23, 27'h000003f9, 5'd17, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d4, 5'd23, 27'h000001eb, 5'd29, 27'h0000015c, 32'h00000400,
  1'd1,  5'd15, 27'h0000034e, 5'd5, 27'h00000053, 5'd2, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000025c, 5'd1, 27'h000001b1, 5'd14, 27'h000000f1, 32'h00000400,
  1'd1,  5'd15, 27'h00000320, 5'd4, 27'h00000319, 5'd22, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000081, 5'd10, 27'h000001cf, 5'd7, 27'h0000002f, 32'h00000400,
  1'd1,  5'd16, 27'h000003f5, 5'd11, 27'h00000060, 5'd18, 27'h00000166, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a9, 5'd14, 27'h0000035e, 5'd29, 27'h0000004a, 32'h00000400,
  1'd1,  5'd16, 27'h000000f8, 5'd20, 27'h00000336, 5'd9, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000005b, 5'd22, 27'h00000319, 5'd15, 27'h0000027d, 32'h00000400,
  1'd1,  5'd20, 27'h000000d3, 5'd22, 27'h000000c8, 5'd26, 27'h0000009b, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000275, 5'd0, 27'h00000351, 5'd7, 27'h0000003f, 32'h00000400,
  1'd1,  5'd26, 27'h00000391, 5'd1, 27'h000001a9, 5'd20, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000005d, 5'd1, 27'h00000006, 5'd29, 27'h00000183, 32'h00000400,
  1'd1,  5'd28, 27'h0000016f, 5'd13, 27'h0000007b, 5'd9, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000006e, 5'd10, 27'h00000299, 5'd18, 27'h00000011, 32'h00000400,
  1'd1,  5'd30, 27'h000003c0, 5'd12, 27'h000002d5, 5'd26, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000092, 5'd22, 27'h0000037e, 5'd7, 27'h00000256, 32'h00000400,
  1'd1,  5'd26, 27'h000002cc, 5'd24, 27'h000001d5, 5'd18, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000047, 5'd23, 27'h00000215, 5'd26, 27'h000002e1, 32'h00000400,
  1'd1,  5'd6, 27'h0000000a, 5'd5, 27'h0000026b, 5'd3, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002e8, 5'd5, 27'h000002c9, 5'd13, 27'h000002dd, 32'h00000400,
  1'd1,  5'd8, 27'h00000202, 5'd5, 27'h000000fb, 5'd24, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000009b, 5'd20, 27'h0000027c, 5'd3, 27'h000002d9, 32'h00000400,
  1'd1,  5'd7, 27'h00000222, 5'd19, 27'h00000055, 5'd13, 27'h000000e7, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000196, 5'd16, 27'h0000021a, 5'd21, 27'h000002ae, 32'h00000400,
  1'd1,  5'd5, 27'h00000277, 5'd30, 27'h00000358, 5'd2, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000268, 5'd29, 27'h00000249, 5'd10, 27'h00000289, 32'h00000400,
  1'd1,  5'd6, 27'h00000127, 5'd30, 27'h0000017e, 5'd23, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039b, 5'd7, 27'h00000287, 5'd0, 27'h000000f1, 32'h00000400,
  1'd1,  5'd20, 27'h0000022a, 5'd9, 27'h00000034, 5'd15, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000332, 5'd5, 27'h0000033d, 5'd23, 27'h000001e4, 32'h00000400,
  1'd1,  5'd17, 27'h00000276, 5'd18, 27'h00000166, 5'd0, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000aa, 5'd17, 27'h000000c1, 5'd12, 27'h00000239, 32'h00000400,
  1'd1,  5'd18, 27'h00000217, 5'd16, 27'h00000109, 5'd24, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001b1, 5'd29, 27'h0000008d, 5'd0, 27'h00000343, 32'h00000400,
  1'd1,  5'd20, 27'h00000120, 5'd26, 27'h00000156, 5'd13, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000044, 5'd27, 27'h00000350, 5'd23, 27'h00000351, 32'h00000400,
  1'd1,  5'd26, 27'h000000f2, 5'd8, 27'h0000010d, 5'd2, 27'h00000180, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002aa, 5'd7, 27'h000000a8, 5'd11, 27'h000000f0, 32'h00000400,
  1'd1,  5'd27, 27'h0000013d, 5'd8, 27'h000003ad, 5'd25, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000392, 5'd18, 27'h0000014e, 5'd1, 27'h000003df, 32'h00000400,
  1'd1,  5'd28, 27'h000002ab, 5'd18, 27'h0000007a, 5'd15, 27'h000001f5, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000148, 5'd19, 27'h000002ef, 5'd22, 27'h00000178, 32'h00000400,
  1'd1,  5'd30, 27'h000000d5, 5'd26, 27'h000001fa, 5'd1, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002f4, 5'd26, 27'h000003d6, 5'd14, 27'h00000049, 32'h00000400,
  1'd1,  5'd28, 27'h0000034e, 5'd29, 27'h000003c9, 5'd23, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b8, 5'd5, 27'h000002b9, 5'd5, 27'h000001f5, 32'h00000400,
  1'd1,  5'd7, 27'h000003a7, 5'd8, 27'h000003cf, 5'd20, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000123, 5'd6, 27'h00000294, 5'd29, 27'h000000eb, 32'h00000400,
  1'd1,  5'd7, 27'h000002b0, 5'd17, 27'h000003ee, 5'd6, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001bb, 5'd19, 27'h00000076, 5'd18, 27'h00000105, 32'h00000400,
  1'd1,  5'd8, 27'h00000007, 5'd19, 27'h00000058, 5'd28, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003b8, 5'd26, 27'h000002f9, 5'd6, 27'h000000f6, 32'h00000400,
  1'd1,  5'd5, 27'h0000031b, 5'd29, 27'h000002a9, 5'd19, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ef, 5'd26, 27'h000003e7, 5'd28, 27'h0000033c, 32'h00000400,
  1'd1,  5'd18, 27'h0000009f, 5'd5, 27'h000001fb, 5'd8, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000382, 5'd5, 27'h00000233, 5'd16, 27'h0000009b, 32'h00000400,
  1'd1,  5'd17, 27'h00000056, 5'd8, 27'h00000155, 5'd30, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000211, 5'd15, 27'h000002ad, 5'd6, 27'h000003ed, 32'h00000400,
  1'd1,  5'd18, 27'h0000021c, 5'd16, 27'h0000036f, 5'd20, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000037a, 5'd17, 27'h00000178, 5'd26, 27'h000002f6, 32'h00000400,
  1'd1,  5'd16, 27'h000000b5, 5'd25, 27'h0000036a, 5'd9, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ed, 5'd29, 27'h000003f6, 5'd17, 27'h00000068, 32'h00000400,
  1'd1,  5'd17, 27'h00000286, 5'd26, 27'h00000157, 5'd27, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000038b, 5'd6, 27'h0000009e, 5'd8, 27'h000003ec, 32'h00000400,
  1'd1,  5'd27, 27'h00000398, 5'd8, 27'h00000051, 5'd18, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003e2, 5'd9, 27'h00000040, 5'd28, 27'h00000247, 32'h00000400,
  1'd1,  5'd29, 27'h0000030f, 5'd19, 27'h00000292, 5'd7, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000215, 5'd19, 27'h00000382, 5'd19, 27'h000000e8, 32'h00000400,
  1'd1,  5'd28, 27'h00000347, 5'd19, 27'h00000298, 5'd29, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000136, 5'd29, 27'h000001e1, 5'd5, 27'h0000019e, 32'h00000400,
  1'd1,  5'd26, 27'h00000107, 5'd30, 27'h00000214, 5'd18, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000039a, 5'd29, 27'h000003b1, 5'd29, 27'h0000032c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000340, 5'd1, 27'h000002d9, 5'd1, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000176, 5'd5, 27'h0000002e, 5'd11, 27'h0000018f, 32'h00000400,
  1'd1,  5'd3, 27'h00000343, 5'd2, 27'h0000016c, 5'd24, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000122, 5'd13, 27'h00000070, 5'd2, 27'h000002ce, 32'h00000400,
  1'd1,  5'd2, 27'h00000323, 5'd12, 27'h000001e5, 5'd11, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000099, 5'd13, 27'h0000007b, 5'd25, 27'h00000202, 32'h00000400,
  1'd1,  5'd0, 27'h00000041, 5'd21, 27'h00000233, 5'd1, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002d3, 5'd21, 27'h000001b1, 5'd11, 27'h0000003f, 32'h00000400,
  1'd1,  5'd3, 27'h0000023c, 5'd25, 27'h000001d8, 5'd23, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ed, 5'd3, 27'h000000a4, 5'd0, 27'h00000010, 32'h00000400,
  1'd1,  5'd12, 27'h00000187, 5'd3, 27'h00000198, 5'd11, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000168, 5'd5, 27'h00000084, 5'd24, 27'h000000f6, 32'h00000400,
  1'd1,  5'd11, 27'h000001e6, 5'd14, 27'h000001f2, 5'd4, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003cd, 5'd14, 27'h0000021b, 5'd12, 27'h0000011c, 32'h00000400,
  1'd1,  5'd15, 27'h000001a3, 5'd13, 27'h0000034c, 5'd21, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000325, 5'd21, 27'h000000fb, 5'd2, 27'h000003ac, 32'h00000400,
  1'd1,  5'd13, 27'h000001b8, 5'd24, 27'h0000010e, 5'd12, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d0, 5'd20, 27'h000003c7, 5'd21, 27'h00000339, 32'h00000400,
  1'd1,  5'd22, 27'h000003fc, 5'd4, 27'h0000002b, 5'd3, 27'h00000283, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001f8, 5'd1, 27'h00000003, 5'd10, 27'h0000037e, 32'h00000400,
  1'd1,  5'd24, 27'h000003f6, 5'd2, 27'h00000219, 5'd21, 27'h0000013c, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003f9, 5'd11, 27'h000001cd, 5'd2, 27'h00000174, 32'h00000400,
  1'd1,  5'd24, 27'h00000143, 5'd13, 27'h00000273, 5'd12, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f6, 5'd11, 27'h00000384, 5'd20, 27'h000002ab, 32'h00000400,
  1'd1,  5'd23, 27'h0000020b, 5'd21, 27'h000002cc, 5'd3, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a8, 5'd25, 27'h0000019f, 5'd14, 27'h000000b8, 32'h00000400,
  1'd1,  5'd22, 27'h0000037f, 5'd21, 27'h00000380, 5'd24, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a6, 5'd3, 27'h0000024e, 5'd6, 27'h000002f4, 32'h00000400,
  1'd1,  5'd0, 27'h000003d0, 5'd0, 27'h00000093, 5'd18, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d4, 5'd0, 27'h000001e6, 5'd29, 27'h0000012e, 32'h00000400,
  1'd1,  5'd2, 27'h000002e1, 5'd13, 27'h0000001b, 5'd9, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000001, 5'd11, 27'h000000d9, 5'd17, 27'h0000031f, 32'h00000400,
  1'd1,  5'd1, 27'h0000035f, 5'd14, 27'h000003d0, 5'd25, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000002e, 5'd25, 27'h00000273, 5'd5, 27'h000001e0, 32'h00000400,
  1'd1,  5'd4, 27'h00000363, 5'd22, 27'h000002b3, 5'd19, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000019f, 5'd21, 27'h000001be, 5'd26, 27'h000001f9, 32'h00000400,
  1'd1,  5'd12, 27'h0000002a, 5'd4, 27'h0000031e, 5'd9, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001a5, 5'd2, 27'h00000295, 5'd18, 27'h0000019d, 32'h00000400,
  1'd1,  5'd11, 27'h00000012, 5'd1, 27'h0000014c, 5'd27, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000347, 5'd11, 27'h00000284, 5'd7, 27'h000002e5, 32'h00000400,
  1'd1,  5'd13, 27'h00000347, 5'd13, 27'h000003c4, 5'd17, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001bc, 5'd14, 27'h000001dd, 5'd28, 27'h00000270, 32'h00000400,
  1'd1,  5'd12, 27'h00000261, 5'd25, 27'h0000034a, 5'd5, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f4, 5'd23, 27'h000002f5, 5'd15, 27'h000002b1, 32'h00000400,
  1'd1,  5'd12, 27'h00000157, 5'd23, 27'h000000d5, 5'd26, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001a8, 5'd1, 27'h0000018c, 5'd8, 27'h0000029d, 32'h00000400,
  1'd1,  5'd24, 27'h0000015a, 5'd2, 27'h00000306, 5'd16, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000031, 5'd4, 27'h00000001, 5'd26, 27'h000002a8, 32'h00000400,
  1'd1,  5'd23, 27'h00000067, 5'd13, 27'h0000033b, 5'd6, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000013d, 5'd12, 27'h000001c0, 5'd16, 27'h00000191, 32'h00000400,
  1'd1,  5'd21, 27'h000002f9, 5'd11, 27'h00000363, 5'd28, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000be, 5'd23, 27'h000000e6, 5'd6, 27'h00000059, 32'h00000400,
  1'd1,  5'd22, 27'h00000071, 5'd22, 27'h00000352, 5'd18, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000078, 5'd23, 27'h000000d1, 5'd26, 27'h000003b4, 32'h00000400,
  1'd1,  5'd0, 27'h000001a9, 5'd5, 27'h00000200, 5'd2, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000009e, 5'd7, 27'h0000036a, 5'd14, 27'h00000061, 32'h00000400,
  1'd1,  5'd3, 27'h000001d3, 5'd6, 27'h0000024b, 5'd21, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000362, 5'd20, 27'h00000090, 5'd1, 27'h000001f0, 32'h00000400,
  1'd1,  5'd4, 27'h0000027d, 5'd16, 27'h0000004f, 5'd14, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002fa, 5'd15, 27'h000003c7, 5'd23, 27'h00000023, 32'h00000400,
  1'd1,  5'd1, 27'h0000014d, 5'd26, 27'h00000247, 5'd3, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000b7, 5'd28, 27'h000002aa, 5'd12, 27'h0000038a, 32'h00000400,
  1'd1,  5'd4, 27'h0000033d, 5'd28, 27'h0000036c, 5'd21, 27'h0000021c, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000031a, 5'd9, 27'h00000153, 5'd3, 27'h00000118, 32'h00000400,
  1'd1,  5'd14, 27'h000000c5, 5'd8, 27'h00000074, 5'd11, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000307, 5'd5, 27'h000003ab, 5'd23, 27'h000000f3, 32'h00000400,
  1'd1,  5'd15, 27'h000000be, 5'd18, 27'h00000341, 5'd3, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000005c, 5'd18, 27'h00000350, 5'd14, 27'h000001fb, 32'h00000400,
  1'd1,  5'd15, 27'h00000199, 5'd16, 27'h000000c5, 5'd22, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000038e, 5'd30, 27'h000001cc, 5'd4, 27'h00000016, 32'h00000400,
  1'd1,  5'd14, 27'h0000030e, 5'd29, 27'h00000001, 5'd12, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000016, 5'd27, 27'h0000003a, 5'd22, 27'h000003c6, 32'h00000400,
  1'd1,  5'd25, 27'h00000051, 5'd10, 27'h0000002c, 5'd5, 27'h00000046, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f0, 5'd8, 27'h000003a0, 5'd11, 27'h0000015d, 32'h00000400,
  1'd1,  5'd20, 27'h00000339, 5'd9, 27'h00000231, 5'd22, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001cc, 5'd19, 27'h0000037a, 5'd0, 27'h00000137, 32'h00000400,
  1'd1,  5'd22, 27'h000002dc, 5'd17, 27'h000001c1, 5'd13, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000075, 5'd17, 27'h0000022b, 5'd23, 27'h0000018c, 32'h00000400,
  1'd1,  5'd21, 27'h0000015b, 5'd29, 27'h00000016, 5'd3, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000221, 5'd30, 27'h0000015c, 5'd13, 27'h0000035d, 32'h00000400,
  1'd1,  5'd24, 27'h0000031e, 5'd29, 27'h0000010a, 5'd22, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020c, 5'd5, 27'h0000010d, 5'd9, 27'h00000218, 32'h00000400,
  1'd1,  5'd5, 27'h0000002b, 5'd6, 27'h0000035c, 5'd17, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002eb, 5'd5, 27'h0000014b, 5'd28, 27'h0000020d, 32'h00000400,
  1'd1,  5'd2, 27'h0000035c, 5'd16, 27'h00000244, 5'd7, 27'h000003ad, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000025b, 5'd16, 27'h00000268, 5'd20, 27'h0000016e, 32'h00000400,
  1'd1,  5'd0, 27'h000000bb, 5'd15, 27'h0000026c, 5'd27, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000240, 5'd26, 27'h0000038d, 5'd9, 27'h000001a5, 32'h00000400,
  1'd1,  5'd2, 27'h00000167, 5'd26, 27'h00000083, 5'd17, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b7, 5'd30, 27'h00000076, 5'd26, 27'h00000070, 32'h00000400,
  1'd1,  5'd10, 27'h000001ec, 5'd9, 27'h00000302, 5'd9, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000015e, 5'd5, 27'h000002e1, 5'd17, 27'h00000400, 32'h00000400,
  1'd1,  5'd13, 27'h0000017e, 5'd7, 27'h0000029b, 5'd26, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000213, 5'd18, 27'h00000278, 5'd6, 27'h00000373, 32'h00000400,
  1'd1,  5'd12, 27'h00000288, 5'd19, 27'h000003dc, 5'd16, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000035c, 5'd15, 27'h00000275, 5'd29, 27'h00000392, 32'h00000400,
  1'd1,  5'd13, 27'h00000042, 5'd26, 27'h0000001c, 5'd7, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e3, 5'd27, 27'h00000252, 5'd19, 27'h00000336, 32'h00000400,
  1'd1,  5'd11, 27'h0000011d, 5'd27, 27'h00000265, 5'd30, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002da, 5'd8, 27'h000000fb, 5'd8, 27'h0000033b, 32'h00000400,
  1'd1,  5'd23, 27'h000000c6, 5'd6, 27'h00000383, 5'd16, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002f4, 5'd5, 27'h00000155, 5'd28, 27'h0000028d, 32'h00000400,
  1'd1,  5'd24, 27'h00000082, 5'd18, 27'h00000253, 5'd5, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000306, 5'd16, 27'h00000212, 5'd15, 27'h00000337, 32'h00000400,
  1'd1,  5'd24, 27'h0000017e, 5'd19, 27'h000001d1, 5'd28, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000397, 5'd26, 27'h000003a9, 5'd6, 27'h000000d3, 32'h00000400,
  1'd1,  5'd23, 27'h000003a0, 5'd28, 27'h00000024, 5'd17, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003d5, 5'd29, 27'h000002bb, 5'd26, 27'h00000233, 32'h00000400,
  1'd1,  5'd8, 27'h00000043, 5'd4, 27'h000000ea, 5'd6, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001c5, 5'd2, 27'h0000036a, 5'd16, 27'h0000038c, 32'h00000400,
  1'd1,  5'd6, 27'h00000136, 5'd5, 27'h00000038, 5'd25, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000013b, 5'd14, 27'h00000069, 5'd0, 27'h0000039e, 32'h00000400,
  1'd1,  5'd8, 27'h000001fc, 5'd13, 27'h00000191, 5'd11, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000018b, 5'd10, 27'h00000219, 5'd22, 27'h0000030e, 32'h00000400,
  1'd1,  5'd8, 27'h00000314, 5'd23, 27'h0000004f, 5'd4, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000318, 5'd21, 27'h00000251, 5'd13, 27'h00000142, 32'h00000400,
  1'd1,  5'd8, 27'h000002ae, 5'd25, 27'h00000038, 5'd21, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d0, 5'd2, 27'h00000109, 5'd6, 27'h00000163, 32'h00000400,
  1'd1,  5'd20, 27'h000000ff, 5'd0, 27'h0000009b, 5'd18, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000238, 5'd5, 27'h00000047, 5'd30, 27'h000001a5, 32'h00000400,
  1'd1,  5'd19, 27'h00000246, 5'd12, 27'h000002d6, 5'd2, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001ad, 5'd15, 27'h00000188, 5'd11, 27'h000000dd, 32'h00000400,
  1'd1,  5'd18, 27'h0000030e, 5'd12, 27'h000000ab, 5'd23, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000c3, 5'd22, 27'h000003b2, 5'd1, 27'h00000268, 32'h00000400,
  1'd1,  5'd19, 27'h000000e8, 5'd23, 27'h00000206, 5'd15, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003ba, 5'd25, 27'h000002db, 5'd21, 27'h0000020d, 32'h00000400,
  1'd1,  5'd26, 27'h000003cc, 5'd1, 27'h000001e9, 5'd3, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e3, 5'd3, 27'h00000001, 5'd11, 27'h000002f2, 32'h00000400,
  1'd1,  5'd26, 27'h0000007e, 5'd1, 27'h00000389, 5'd24, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000011f, 5'd13, 27'h000001e5, 5'd4, 27'h000002cf, 32'h00000400,
  1'd1,  5'd28, 27'h000000fb, 5'd12, 27'h00000193, 5'd10, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000008, 5'd10, 27'h000003d2, 5'd24, 27'h00000026, 32'h00000400,
  1'd1,  5'd27, 27'h00000024, 5'd22, 27'h000001f4, 5'd4, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000244, 5'd23, 27'h0000018b, 5'd10, 27'h000002af, 32'h00000400,
  1'd1,  5'd28, 27'h000001ee, 5'd21, 27'h0000028f, 5'd23, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000374, 5'd1, 27'h00000190, 5'd0, 27'h00000068, 32'h00000400,
  1'd1,  5'd7, 27'h00000191, 5'd1, 27'h000001ef, 5'd12, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000022f, 5'd2, 27'h000002b4, 5'd24, 27'h000000a6, 32'h00000400,
  1'd1,  5'd9, 27'h00000131, 5'd14, 27'h000002f6, 5'd6, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000ea, 5'd13, 27'h000003f8, 5'd17, 27'h000000f7, 32'h00000400,
  1'd1,  5'd8, 27'h000000d7, 5'd14, 27'h000001b7, 5'd26, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000015a, 5'd20, 27'h00000347, 5'd9, 27'h000001c3, 32'h00000400,
  1'd1,  5'd8, 27'h00000234, 5'd22, 27'h00000055, 5'd19, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002ac, 5'd23, 27'h00000388, 5'd28, 27'h00000249, 32'h00000400,
  1'd1,  5'd18, 27'h0000003b, 5'd1, 27'h000001c9, 5'd1, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000196, 5'd4, 27'h0000031b, 5'd12, 27'h000001e8, 32'h00000400,
  1'd1,  5'd16, 27'h00000119, 5'd3, 27'h000003a1, 5'd24, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f6, 5'd12, 27'h00000353, 5'd6, 27'h00000228, 32'h00000400,
  1'd1,  5'd19, 27'h00000234, 5'd11, 27'h000002a3, 5'd19, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000013c, 5'd15, 27'h00000134, 5'd27, 27'h00000177, 32'h00000400,
  1'd1,  5'd19, 27'h00000076, 5'd24, 27'h000001e0, 5'd8, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000039, 5'd21, 27'h0000005a, 5'd17, 27'h00000375, 32'h00000400,
  1'd1,  5'd19, 27'h00000203, 5'd25, 27'h000002bc, 5'd29, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000316, 5'd4, 27'h000000b9, 5'd9, 27'h00000300, 32'h00000400,
  1'd1,  5'd28, 27'h000003b7, 5'd0, 27'h0000024c, 5'd18, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000160, 5'd1, 27'h0000020a, 5'd29, 27'h00000044, 32'h00000400,
  1'd1,  5'd27, 27'h000000e8, 5'd11, 27'h000003ca, 5'd8, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000174, 5'd11, 27'h00000013, 5'd20, 27'h00000065, 32'h00000400,
  1'd1,  5'd28, 27'h0000035e, 5'd11, 27'h000000f0, 5'd29, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000010c, 5'd22, 27'h00000380, 5'd7, 27'h000000b0, 32'h00000400,
  1'd1,  5'd30, 27'h00000104, 5'd23, 27'h000001d3, 5'd17, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000066, 5'd24, 27'h0000016b, 5'd27, 27'h000000e0, 32'h00000400,
  1'd1,  5'd9, 27'h00000317, 5'd8, 27'h0000020b, 5'd4, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000291, 5'd9, 27'h000001c0, 5'd13, 27'h00000223, 32'h00000400,
  1'd1,  5'd9, 27'h00000202, 5'd6, 27'h00000321, 5'd24, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e9, 5'd16, 27'h000000b8, 5'd1, 27'h00000002, 32'h00000400,
  1'd1,  5'd9, 27'h0000039d, 5'd19, 27'h0000008e, 5'd15, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000032e, 5'd20, 27'h000001a2, 5'd23, 27'h00000177, 32'h00000400,
  1'd1,  5'd7, 27'h00000357, 5'd27, 27'h000003de, 5'd2, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000031b, 5'd26, 27'h00000072, 5'd11, 27'h00000391, 32'h00000400,
  1'd1,  5'd5, 27'h0000027c, 5'd27, 27'h00000009, 5'd20, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000036, 5'd7, 27'h0000023c, 5'd0, 27'h0000027a, 32'h00000400,
  1'd1,  5'd18, 27'h000002b0, 5'd9, 27'h00000184, 5'd14, 27'h0000029c, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000027c, 5'd7, 27'h00000341, 5'd24, 27'h000003f6, 32'h00000400,
  1'd1,  5'd17, 27'h000001ee, 5'd19, 27'h00000061, 5'd1, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ad, 5'd20, 27'h00000258, 5'd13, 27'h0000001c, 32'h00000400,
  1'd1,  5'd17, 27'h00000118, 5'd18, 27'h00000246, 5'd24, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000054, 5'd28, 27'h00000391, 5'd3, 27'h00000121, 32'h00000400,
  1'd1,  5'd18, 27'h000001d8, 5'd29, 27'h000002e9, 5'd12, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000017, 5'd29, 27'h0000025c, 5'd23, 27'h00000281, 32'h00000400,
  1'd1,  5'd25, 27'h00000357, 5'd6, 27'h0000000a, 5'd4, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000003b, 5'd8, 27'h0000035d, 5'd12, 27'h00000390, 32'h00000400,
  1'd1,  5'd28, 27'h00000131, 5'd6, 27'h00000005, 5'd24, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000245, 5'd19, 27'h0000035e, 5'd1, 27'h000002fb, 32'h00000400,
  1'd1,  5'd29, 27'h00000240, 5'd20, 27'h00000228, 5'd11, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000060, 5'd19, 27'h000000ad, 5'd23, 27'h000003ca, 32'h00000400,
  1'd1,  5'd30, 27'h000003f2, 5'd29, 27'h00000098, 5'd0, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002b9, 5'd26, 27'h000003ab, 5'd12, 27'h000001bb, 32'h00000400,
  1'd1,  5'd27, 27'h00000223, 5'd26, 27'h00000370, 5'd25, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000278, 5'd7, 27'h00000310, 5'd6, 27'h00000250, 32'h00000400,
  1'd1,  5'd8, 27'h000000bb, 5'd8, 27'h000003b1, 5'd17, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000312, 5'd9, 27'h000002d1, 5'd27, 27'h00000292, 32'h00000400,
  1'd1,  5'd7, 27'h000003f8, 5'd19, 27'h00000384, 5'd7, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001c5, 5'd17, 27'h000001d1, 5'd17, 27'h00000042, 32'h00000400,
  1'd1,  5'd7, 27'h00000283, 5'd20, 27'h000000bf, 5'd27, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000310, 5'd28, 27'h0000015c, 5'd6, 27'h0000003e, 32'h00000400,
  1'd1,  5'd8, 27'h00000225, 5'd29, 27'h00000380, 5'd15, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000033a, 5'd29, 27'h00000090, 5'd26, 27'h000002b0, 32'h00000400,
  1'd1,  5'd20, 27'h00000032, 5'd5, 27'h000003fa, 5'd6, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e0, 5'd10, 27'h000000c9, 5'd20, 27'h000000d8, 32'h00000400,
  1'd1,  5'd17, 27'h000000d7, 5'd5, 27'h000002cf, 5'd30, 27'h00000393, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000029d, 5'd19, 27'h000001a6, 5'd9, 27'h00000215, 32'h00000400,
  1'd1,  5'd16, 27'h00000269, 5'd18, 27'h000002fe, 5'd19, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000034, 5'd18, 27'h0000031c, 5'd27, 27'h000000d3, 32'h00000400,
  1'd1,  5'd16, 27'h0000012d, 5'd26, 27'h00000170, 5'd9, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000010e, 5'd26, 27'h0000020e, 5'd17, 27'h000001f3, 32'h00000400,
  1'd1,  5'd19, 27'h000000b3, 5'd28, 27'h000001c9, 5'd28, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d5, 5'd8, 27'h0000037d, 5'd9, 27'h0000036f, 32'h00000400,
  1'd1,  5'd29, 27'h00000127, 5'd9, 27'h0000035b, 5'd17, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002af, 5'd6, 27'h00000168, 5'd26, 27'h000001fc, 32'h00000400,
  1'd1,  5'd27, 27'h00000235, 5'd18, 27'h000002c7, 5'd8, 27'h000002b8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000101, 5'd17, 27'h00000390, 5'd15, 27'h000002cc, 32'h00000400,
  1'd1,  5'd27, 27'h00000089, 5'd15, 27'h000003bd, 5'd28, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000019c, 5'd26, 27'h000002b9, 5'd9, 27'h00000215, 32'h00000400,
  1'd1,  5'd27, 27'h000001a1, 5'd28, 27'h00000169, 5'd18, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002fc, 5'd26, 27'h0000020a, 5'd29, 27'h000000de, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001d5, 5'd4, 27'h000000bc, 5'd1, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001e5, 5'd3, 27'h000003f0, 5'd14, 27'h0000022f, 32'h00000400,
  1'd1,  5'd1, 27'h000002c4, 5'd1, 27'h00000309, 5'd20, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001b7, 5'd14, 27'h0000026e, 5'd0, 27'h00000228, 32'h00000400,
  1'd1,  5'd1, 27'h00000340, 5'd15, 27'h000001e7, 5'd14, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000260, 5'd12, 27'h00000232, 5'd22, 27'h000003c6, 32'h00000400,
  1'd1,  5'd2, 27'h00000275, 5'd20, 27'h00000366, 5'd2, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003a1, 5'd22, 27'h0000006f, 5'd11, 27'h000001a1, 32'h00000400,
  1'd1,  5'd4, 27'h00000202, 5'd22, 27'h00000302, 5'd24, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ef, 5'd4, 27'h00000272, 5'd1, 27'h00000241, 32'h00000400,
  1'd1,  5'd14, 27'h0000007c, 5'd5, 27'h0000007a, 5'd14, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000018a, 5'd0, 27'h00000381, 5'd25, 27'h0000029e, 32'h00000400,
  1'd1,  5'd14, 27'h00000162, 5'd12, 27'h000000b8, 5'd4, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000351, 5'd12, 27'h0000029a, 5'd13, 27'h000002ec, 32'h00000400,
  1'd1,  5'd12, 27'h0000023a, 5'd14, 27'h00000108, 5'd22, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018e, 5'd25, 27'h000002f9, 5'd4, 27'h00000340, 32'h00000400,
  1'd1,  5'd12, 27'h00000130, 5'd24, 27'h000000b0, 5'd13, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002bc, 5'd24, 27'h00000375, 5'd23, 27'h00000165, 32'h00000400,
  1'd1,  5'd23, 27'h0000026b, 5'd3, 27'h00000022, 5'd4, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002da, 5'd5, 27'h00000028, 5'd13, 27'h000003cd, 32'h00000400,
  1'd1,  5'd23, 27'h000001a4, 5'd0, 27'h0000026d, 5'd23, 27'h00000105, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003d1, 5'd12, 27'h0000027f, 5'd3, 27'h0000022b, 32'h00000400,
  1'd1,  5'd21, 27'h000002a7, 5'd13, 27'h00000179, 5'd14, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000b4, 5'd15, 27'h00000040, 5'd20, 27'h000003f5, 32'h00000400,
  1'd1,  5'd23, 27'h000003a9, 5'd23, 27'h000003da, 5'd5, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000020b, 5'd25, 27'h00000305, 5'd14, 27'h000000dc, 32'h00000400,
  1'd1,  5'd24, 27'h0000028b, 5'd22, 27'h0000028c, 5'd24, 27'h00000390, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000005, 5'd2, 27'h0000005c, 5'd6, 27'h000000fb, 32'h00000400,
  1'd1,  5'd4, 27'h000000d1, 5'd1, 27'h000000e1, 5'd20, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003dd, 5'd4, 27'h000001b9, 5'd26, 27'h00000325, 32'h00000400,
  1'd1,  5'd0, 27'h00000132, 5'd14, 27'h000002a2, 5'd5, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000e3, 5'd11, 27'h00000341, 5'd20, 27'h000001f8, 32'h00000400,
  1'd1,  5'd2, 27'h000000c1, 5'd13, 27'h00000041, 5'd28, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002a9, 5'd23, 27'h000000e4, 5'd9, 27'h000000ce, 32'h00000400,
  1'd1,  5'd2, 27'h000000f7, 5'd24, 27'h000001f8, 5'd20, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000135, 5'd24, 27'h00000140, 5'd29, 27'h000001d3, 32'h00000400,
  1'd1,  5'd15, 27'h0000002b, 5'd3, 27'h00000340, 5'd6, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000337, 5'd2, 27'h000001b6, 5'd19, 27'h000003d7, 32'h00000400,
  1'd1,  5'd14, 27'h00000277, 5'd1, 27'h00000376, 5'd27, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000011b, 5'd11, 27'h000001e0, 5'd10, 27'h00000081, 32'h00000400,
  1'd1,  5'd14, 27'h0000015b, 5'd15, 27'h000001e1, 5'd18, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000016b, 5'd10, 27'h00000157, 5'd26, 27'h000003fb, 32'h00000400,
  1'd1,  5'd13, 27'h000001a1, 5'd21, 27'h00000142, 5'd8, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000238, 5'd24, 27'h0000020b, 5'd16, 27'h000002c7, 32'h00000400,
  1'd1,  5'd14, 27'h00000154, 5'd20, 27'h00000349, 5'd28, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000112, 5'd3, 27'h0000000a, 5'd8, 27'h00000272, 32'h00000400,
  1'd1,  5'd24, 27'h000002c8, 5'd1, 27'h00000199, 5'd16, 27'h00000135, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002a3, 5'd4, 27'h000001c0, 5'd30, 27'h000001ee, 32'h00000400,
  1'd1,  5'd23, 27'h00000027, 5'd11, 27'h00000292, 5'd6, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000f9, 5'd11, 27'h000001b2, 5'd15, 27'h00000287, 32'h00000400,
  1'd1,  5'd23, 27'h000001c0, 5'd13, 27'h0000012f, 5'd30, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000002e, 5'd25, 27'h000002af, 5'd9, 27'h00000200, 32'h00000400,
  1'd1,  5'd22, 27'h00000354, 5'd24, 27'h000000e4, 5'd19, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000029a, 5'd22, 27'h000000b6, 5'd30, 27'h000000c4, 32'h00000400,
  1'd1,  5'd1, 27'h000002b6, 5'd7, 27'h000003d0, 5'd3, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000024c, 5'd10, 27'h00000106, 5'd11, 27'h00000220, 32'h00000400,
  1'd1,  5'd0, 27'h00000388, 5'd7, 27'h000001ad, 5'd20, 27'h000003b9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000095, 5'd18, 27'h000001f0, 5'd3, 27'h000002b6, 32'h00000400,
  1'd1,  5'd1, 27'h00000000, 5'd16, 27'h000001db, 5'd15, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000004b, 5'd17, 27'h0000037f, 5'd24, 27'h000002c9, 32'h00000400,
  1'd1,  5'd1, 27'h00000161, 5'd28, 27'h000002ee, 5'd1, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003db, 5'd29, 27'h0000010b, 5'd12, 27'h000001b3, 32'h00000400,
  1'd1,  5'd3, 27'h00000298, 5'd29, 27'h00000259, 5'd23, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000012a, 5'd5, 27'h00000335, 5'd4, 27'h00000127, 32'h00000400,
  1'd1,  5'd10, 27'h000001cc, 5'd5, 27'h00000390, 5'd12, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000023c, 5'd6, 27'h0000014d, 5'd22, 27'h00000164, 32'h00000400,
  1'd1,  5'd12, 27'h000001a7, 5'd19, 27'h000001e3, 5'd3, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000118, 5'd15, 27'h00000363, 5'd13, 27'h0000003d, 32'h00000400,
  1'd1,  5'd11, 27'h000002c7, 5'd18, 27'h000003b2, 5'd24, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000194, 5'd28, 27'h000001ed, 5'd0, 27'h000001a9, 32'h00000400,
  1'd1,  5'd12, 27'h00000376, 5'd30, 27'h000003e2, 5'd11, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001f5, 5'd28, 27'h000002b1, 5'd21, 27'h0000021b, 32'h00000400,
  1'd1,  5'd24, 27'h00000068, 5'd6, 27'h000002f8, 5'd4, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019c, 5'd6, 27'h0000031b, 5'd11, 27'h00000326, 32'h00000400,
  1'd1,  5'd21, 27'h00000184, 5'd8, 27'h0000004e, 5'd23, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000271, 5'd17, 27'h00000337, 5'd0, 27'h0000031b, 32'h00000400,
  1'd1,  5'd22, 27'h0000021e, 5'd18, 27'h00000077, 5'd14, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000046, 5'd16, 27'h000003a1, 5'd22, 27'h000000fe, 32'h00000400,
  1'd1,  5'd22, 27'h00000098, 5'd29, 27'h000002f0, 5'd4, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000009f, 5'd27, 27'h00000252, 5'd12, 27'h0000005d, 32'h00000400,
  1'd1,  5'd23, 27'h000002f4, 5'd29, 27'h0000031d, 5'd24, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003f4, 5'd6, 27'h00000002, 5'd8, 27'h0000015a, 32'h00000400,
  1'd1,  5'd2, 27'h000003db, 5'd6, 27'h000001c1, 5'd17, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000001d, 5'd5, 27'h00000181, 5'd29, 27'h000001ca, 32'h00000400,
  1'd1,  5'd0, 27'h0000026a, 5'd15, 27'h00000337, 5'd6, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002be, 5'd19, 27'h00000378, 5'd18, 27'h00000002, 32'h00000400,
  1'd1,  5'd0, 27'h000001e9, 5'd18, 27'h0000004a, 5'd28, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003d2, 5'd30, 27'h00000231, 5'd7, 27'h000002b5, 32'h00000400,
  1'd1,  5'd5, 27'h00000058, 5'd27, 27'h00000171, 5'd20, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ae, 5'd27, 27'h0000030b, 5'd27, 27'h000001a9, 32'h00000400,
  1'd1,  5'd12, 27'h0000036e, 5'd6, 27'h0000025d, 5'd8, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000bf, 5'd7, 27'h00000393, 5'd16, 27'h00000376, 32'h00000400,
  1'd1,  5'd13, 27'h00000069, 5'd7, 27'h00000166, 5'd30, 27'h00000052, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000a7, 5'd19, 27'h00000106, 5'd5, 27'h000000ff, 32'h00000400,
  1'd1,  5'd11, 27'h00000372, 5'd20, 27'h00000070, 5'd19, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000112, 5'd18, 27'h000000f1, 5'd25, 27'h000003a6, 32'h00000400,
  1'd1,  5'd14, 27'h00000331, 5'd28, 27'h000001e1, 5'd9, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002f, 5'd27, 27'h00000297, 5'd18, 27'h0000038c, 32'h00000400,
  1'd1,  5'd10, 27'h000002d1, 5'd27, 27'h000002d7, 5'd28, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000030b, 5'd8, 27'h00000303, 5'd7, 27'h000001d4, 32'h00000400,
  1'd1,  5'd21, 27'h0000022b, 5'd6, 27'h0000030f, 5'd19, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000097, 5'd8, 27'h0000023a, 5'd27, 27'h0000012d, 32'h00000400,
  1'd1,  5'd23, 27'h0000006d, 5'd18, 27'h00000127, 5'd8, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000183, 5'd20, 27'h00000103, 5'd16, 27'h00000001, 32'h00000400,
  1'd1,  5'd24, 27'h000001ad, 5'd16, 27'h000000b1, 5'd30, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000032a, 5'd28, 27'h00000191, 5'd8, 27'h0000035e, 32'h00000400,
  1'd1,  5'd24, 27'h000001b1, 5'd29, 27'h000000df, 5'd17, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002a1, 5'd27, 27'h000000cc, 5'd29, 27'h0000018d, 32'h00000400,
  1'd1,  5'd9, 27'h000002e3, 5'd2, 27'h00000080, 5'd8, 27'h00000117, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f9, 5'd4, 27'h0000033b, 5'd20, 27'h000002a5, 32'h00000400,
  1'd1,  5'd8, 27'h0000023f, 5'd0, 27'h000003fa, 5'd29, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000042, 5'd14, 27'h00000322, 5'd3, 27'h00000087, 32'h00000400,
  1'd1,  5'd6, 27'h00000191, 5'd13, 27'h00000181, 5'd11, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000ea, 5'd12, 27'h000000ae, 5'd23, 27'h00000198, 32'h00000400,
  1'd1,  5'd8, 27'h000003a6, 5'd25, 27'h000001ba, 5'd0, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000098, 5'd22, 27'h000003cb, 5'd10, 27'h000003e2, 32'h00000400,
  1'd1,  5'd8, 27'h00000389, 5'd20, 27'h000002d1, 5'd24, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002ac, 5'd4, 27'h000002a4, 5'd6, 27'h0000002b, 32'h00000400,
  1'd1,  5'd16, 27'h0000022a, 5'd1, 27'h00000162, 5'd16, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000017c, 5'd4, 27'h00000164, 5'd26, 27'h0000033d, 32'h00000400,
  1'd1,  5'd16, 27'h000003c4, 5'd11, 27'h0000031f, 5'd1, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000239, 5'd11, 27'h000003d5, 5'd14, 27'h00000308, 32'h00000400,
  1'd1,  5'd15, 27'h000003ef, 5'd14, 27'h00000315, 5'd23, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000327, 5'd21, 27'h000002aa, 5'd1, 27'h00000317, 32'h00000400,
  1'd1,  5'd19, 27'h0000019a, 5'd23, 27'h0000027b, 5'd14, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000029b, 5'd22, 27'h00000015, 5'd24, 27'h0000022e, 32'h00000400,
  1'd1,  5'd28, 27'h000002b1, 5'd0, 27'h00000142, 5'd3, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000363, 5'd0, 27'h00000324, 5'd11, 27'h00000058, 32'h00000400,
  1'd1,  5'd26, 27'h000001a3, 5'd0, 27'h00000382, 5'd21, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000340, 5'd10, 27'h00000264, 5'd4, 27'h000001a9, 32'h00000400,
  1'd1,  5'd27, 27'h0000002d, 5'd13, 27'h0000034d, 5'd11, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000150, 5'd11, 27'h000000b1, 5'd24, 27'h000003cd, 32'h00000400,
  1'd1,  5'd29, 27'h00000398, 5'd24, 27'h00000378, 5'd4, 27'h0000032d, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000095, 5'd24, 27'h000002b9, 5'd14, 27'h00000285, 32'h00000400,
  1'd1,  5'd27, 27'h000002cb, 5'd22, 27'h0000032f, 5'd25, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000163, 5'd0, 27'h0000030c, 5'd0, 27'h000001c6, 32'h00000400,
  1'd1,  5'd7, 27'h000003b8, 5'd4, 27'h000002ee, 5'd14, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000021d, 5'd0, 27'h000003e7, 5'd22, 27'h000000d9, 32'h00000400,
  1'd1,  5'd6, 27'h00000210, 5'd12, 27'h000003dd, 5'd9, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000024a, 5'd14, 27'h000003e4, 5'd18, 27'h000003cd, 32'h00000400,
  1'd1,  5'd5, 27'h0000012d, 5'd11, 27'h000001d6, 5'd30, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000356, 5'd22, 27'h00000074, 5'd6, 27'h000001d5, 32'h00000400,
  1'd1,  5'd9, 27'h0000037b, 5'd22, 27'h000003c7, 5'd17, 27'h0000007b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000035e, 5'd22, 27'h00000333, 5'd27, 27'h00000321, 32'h00000400,
  1'd1,  5'd18, 27'h0000000c, 5'd2, 27'h000000e2, 5'd3, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000198, 5'd4, 27'h0000007a, 5'd10, 27'h000002b5, 32'h00000400,
  1'd1,  5'd16, 27'h000002fd, 5'd0, 27'h00000092, 5'd21, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000cf, 5'd13, 27'h0000026d, 5'd7, 27'h0000034f, 32'h00000400,
  1'd1,  5'd16, 27'h000000e4, 5'd12, 27'h000001fb, 5'd17, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030f, 5'd13, 27'h000003e9, 5'd26, 27'h0000013c, 32'h00000400,
  1'd1,  5'd19, 27'h000003a8, 5'd24, 27'h00000027, 5'd9, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000298, 5'd22, 27'h00000329, 5'd19, 27'h000003d5, 32'h00000400,
  1'd1,  5'd19, 27'h0000005b, 5'd22, 27'h000002c6, 5'd27, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002e9, 5'd4, 27'h000002f0, 5'd5, 27'h0000035e, 32'h00000400,
  1'd1,  5'd26, 27'h000002f0, 5'd1, 27'h000000f5, 5'd18, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002d7, 5'd2, 27'h000000c3, 5'd27, 27'h000003c7, 32'h00000400,
  1'd1,  5'd28, 27'h000001dd, 5'd12, 27'h000001fd, 5'd6, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000107, 5'd15, 27'h000001e4, 5'd15, 27'h000002f1, 32'h00000400,
  1'd1,  5'd27, 27'h0000007b, 5'd10, 27'h00000205, 5'd27, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000014b, 5'd25, 27'h00000016, 5'd9, 27'h00000130, 32'h00000400,
  1'd1,  5'd27, 27'h000000c8, 5'd23, 27'h00000163, 5'd16, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002a2, 5'd25, 27'h0000008c, 5'd29, 27'h00000105, 32'h00000400,
  1'd1,  5'd6, 27'h00000198, 5'd5, 27'h000000f7, 5'd0, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000076, 5'd9, 27'h00000371, 5'd12, 27'h00000010, 32'h00000400,
  1'd1,  5'd8, 27'h000003cd, 5'd7, 27'h00000101, 5'd23, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000322, 5'd20, 27'h0000018b, 5'd3, 27'h000000ad, 32'h00000400,
  1'd1,  5'd9, 27'h000003fa, 5'd20, 27'h00000205, 5'd13, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002a3, 5'd18, 27'h000001ff, 5'd21, 27'h000001a5, 32'h00000400,
  1'd1,  5'd5, 27'h00000355, 5'd26, 27'h00000316, 5'd0, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000015d, 5'd29, 27'h0000031e, 5'd10, 27'h000002f2, 32'h00000400,
  1'd1,  5'd6, 27'h0000006a, 5'd26, 27'h00000380, 5'd25, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000000, 5'd6, 27'h000002ad, 5'd4, 27'h0000031e, 32'h00000400,
  1'd1,  5'd17, 27'h00000351, 5'd7, 27'h00000078, 5'd12, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000028c, 5'd6, 27'h0000019a, 5'd23, 27'h000000d6, 32'h00000400,
  1'd1,  5'd17, 27'h000000e9, 5'd17, 27'h000000f2, 5'd0, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000109, 5'd15, 27'h0000037f, 5'd13, 27'h000001e4, 32'h00000400,
  1'd1,  5'd15, 27'h00000242, 5'd19, 27'h000000a2, 5'd24, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000160, 5'd28, 27'h000001f4, 5'd3, 27'h000002b1, 32'h00000400,
  1'd1,  5'd18, 27'h0000012b, 5'd27, 27'h00000301, 5'd11, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000f0, 5'd30, 27'h000001a4, 5'd22, 27'h0000029a, 32'h00000400,
  1'd1,  5'd30, 27'h0000015e, 5'd7, 27'h000000fa, 5'd0, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000dc, 5'd9, 27'h00000385, 5'd14, 27'h00000115, 32'h00000400,
  1'd1,  5'd26, 27'h00000290, 5'd9, 27'h0000031c, 5'd25, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000032a, 5'd19, 27'h0000035a, 5'd3, 27'h000003da, 32'h00000400,
  1'd1,  5'd28, 27'h0000000d, 5'd16, 27'h00000200, 5'd12, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000254, 5'd16, 27'h00000296, 5'd22, 27'h000002b3, 32'h00000400,
  1'd1,  5'd28, 27'h00000341, 5'd28, 27'h0000022b, 5'd4, 27'h0000024d, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000027f, 5'd30, 27'h0000025b, 5'd11, 27'h0000022b, 32'h00000400,
  1'd1,  5'd27, 27'h00000024, 5'd28, 27'h00000279, 5'd23, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000026, 5'd6, 27'h0000033e, 5'd7, 27'h000000f5, 32'h00000400,
  1'd1,  5'd5, 27'h000003e5, 5'd7, 27'h00000183, 5'd15, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000e4, 5'd5, 27'h000002df, 5'd29, 27'h000002f5, 32'h00000400,
  1'd1,  5'd7, 27'h00000240, 5'd19, 27'h000001af, 5'd7, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003b6, 5'd16, 27'h00000027, 5'd16, 27'h0000025b, 32'h00000400,
  1'd1,  5'd7, 27'h000000d4, 5'd17, 27'h000002f0, 5'd30, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000004, 5'd27, 27'h00000267, 5'd5, 27'h000003ef, 32'h00000400,
  1'd1,  5'd6, 27'h000002b4, 5'd26, 27'h00000092, 5'd16, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003de, 5'd27, 27'h000002da, 5'd29, 27'h0000003a, 32'h00000400,
  1'd1,  5'd17, 27'h000003ff, 5'd6, 27'h00000202, 5'd7, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000215, 5'd6, 27'h0000029c, 5'd19, 27'h00000229, 32'h00000400,
  1'd1,  5'd16, 27'h00000354, 5'd6, 27'h000003e3, 5'd27, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000007c, 5'd17, 27'h00000375, 5'd8, 27'h0000012c, 32'h00000400,
  1'd1,  5'd17, 27'h00000330, 5'd19, 27'h000001b6, 5'd20, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001da, 5'd16, 27'h00000363, 5'd30, 27'h000002a8, 32'h00000400,
  1'd1,  5'd18, 27'h0000000f, 5'd30, 27'h0000007b, 5'd7, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000009c, 5'd27, 27'h000000ff, 5'd18, 27'h00000167, 32'h00000400,
  1'd1,  5'd19, 27'h000000c4, 5'd27, 27'h00000132, 5'd28, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000384, 5'd10, 27'h0000012d, 5'd9, 27'h0000023a, 32'h00000400,
  1'd1,  5'd28, 27'h00000126, 5'd6, 27'h000003eb, 5'd16, 27'h00000233, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000114, 5'd8, 27'h000002a6, 5'd26, 27'h0000017f, 32'h00000400,
  1'd1,  5'd26, 27'h000001f5, 5'd17, 27'h000003b3, 5'd10, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000026a, 5'd19, 27'h000002ee, 5'd19, 27'h00000395, 32'h00000400,
  1'd1,  5'd29, 27'h00000288, 5'd19, 27'h00000216, 5'd28, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000204, 5'd26, 27'h00000340, 5'd10, 27'h000000ea, 32'h00000400,
  1'd1,  5'd26, 27'h000000c4, 5'd29, 27'h00000379, 5'd17, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000030, 5'd28, 27'h00000315, 5'd26, 27'h0000012a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h000003c0, 5'd0, 27'h0000005c, 5'd4, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000392, 5'd0, 27'h000001f9, 5'd10, 27'h000002fe, 32'h00000400,
  1'd1,  5'd3, 27'h00000082, 5'd1, 27'h00000047, 5'd24, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000028e, 5'd14, 27'h0000014d, 5'd1, 27'h000000f4, 32'h00000400,
  1'd1,  5'd0, 27'h000003a2, 5'd13, 27'h000000f3, 5'd13, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e1, 5'd11, 27'h000001a3, 5'd24, 27'h000002e7, 32'h00000400,
  1'd1,  5'd1, 27'h00000095, 5'd25, 27'h00000213, 5'd1, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000349, 5'd20, 27'h00000322, 5'd11, 27'h00000030, 32'h00000400,
  1'd1,  5'd4, 27'h0000039e, 5'd22, 27'h0000033b, 5'd25, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001b2, 5'd3, 27'h0000004f, 5'd1, 27'h000003c9, 32'h00000400,
  1'd1,  5'd10, 27'h00000353, 5'd2, 27'h000002e6, 5'd12, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000030, 5'd3, 27'h00000241, 5'd22, 27'h00000236, 32'h00000400,
  1'd1,  5'd13, 27'h00000214, 5'd11, 27'h000001e6, 5'd0, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000cd, 5'd11, 27'h00000355, 5'd11, 27'h0000023f, 32'h00000400,
  1'd1,  5'd11, 27'h0000003e, 5'd15, 27'h00000071, 5'd21, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f3, 5'd22, 27'h00000284, 5'd2, 27'h00000115, 32'h00000400,
  1'd1,  5'd14, 27'h00000085, 5'd24, 27'h00000233, 5'd13, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002df, 5'd21, 27'h0000020a, 5'd23, 27'h00000089, 32'h00000400,
  1'd1,  5'd22, 27'h00000394, 5'd0, 27'h000000ae, 5'd4, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000023c, 5'd4, 27'h00000096, 5'd10, 27'h0000018d, 32'h00000400,
  1'd1,  5'd22, 27'h000002b4, 5'd4, 27'h000003d3, 5'd22, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002d7, 5'd11, 27'h0000031d, 5'd3, 27'h00000289, 32'h00000400,
  1'd1,  5'd21, 27'h00000143, 5'd13, 27'h000001e6, 5'd11, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000352, 5'd13, 27'h000003cc, 5'd24, 27'h000000e1, 32'h00000400,
  1'd1,  5'd21, 27'h00000343, 5'd23, 27'h0000015f, 5'd0, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000164, 5'd24, 27'h000003ad, 5'd13, 27'h00000284, 32'h00000400,
  1'd1,  5'd25, 27'h00000137, 5'd22, 27'h000002fc, 5'd22, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000bc, 5'd1, 27'h00000251, 5'd7, 27'h00000192, 32'h00000400,
  1'd1,  5'd4, 27'h000002fa, 5'd1, 27'h000003af, 5'd20, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000078, 5'd0, 27'h0000039a, 5'd25, 27'h0000037d, 32'h00000400,
  1'd1,  5'd3, 27'h00000044, 5'd13, 27'h000002a2, 5'd7, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018a, 5'd14, 27'h000001aa, 5'd19, 27'h00000219, 32'h00000400,
  1'd1,  5'd2, 27'h0000009e, 5'd14, 27'h00000113, 5'd29, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000033f, 5'd25, 27'h000000f1, 5'd9, 27'h00000196, 32'h00000400,
  1'd1,  5'd3, 27'h0000024c, 5'd20, 27'h000002c9, 5'd17, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002cf, 5'd24, 27'h000001ff, 5'd27, 27'h000002bf, 32'h00000400,
  1'd1,  5'd12, 27'h000002d0, 5'd3, 27'h00000018, 5'd7, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003c0, 5'd1, 27'h00000259, 5'd17, 27'h000000ec, 32'h00000400,
  1'd1,  5'd11, 27'h0000008d, 5'd1, 27'h000001f2, 5'd25, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000097, 5'd14, 27'h000001d5, 5'd5, 27'h000000b2, 32'h00000400,
  1'd1,  5'd12, 27'h00000301, 5'd14, 27'h000001ae, 5'd18, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000f3, 5'd10, 27'h00000190, 5'd27, 27'h00000169, 32'h00000400,
  1'd1,  5'd13, 27'h0000019e, 5'd22, 27'h000001bd, 5'd7, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000037b, 5'd23, 27'h000003a8, 5'd20, 27'h000000ff, 32'h00000400,
  1'd1,  5'd13, 27'h00000124, 5'd21, 27'h000003b5, 5'd26, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000033a, 5'd3, 27'h00000046, 5'd10, 27'h0000009a, 32'h00000400,
  1'd1,  5'd24, 27'h0000010b, 5'd1, 27'h00000060, 5'd19, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000217, 5'd1, 27'h00000211, 5'd26, 27'h00000075, 32'h00000400,
  1'd1,  5'd25, 27'h00000052, 5'd13, 27'h0000007a, 5'd6, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000019b, 5'd10, 27'h000002e0, 5'd19, 27'h0000001a, 32'h00000400,
  1'd1,  5'd20, 27'h00000393, 5'd10, 27'h000001cb, 5'd26, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000344, 5'd24, 27'h000001d6, 5'd9, 27'h000003f7, 32'h00000400,
  1'd1,  5'd23, 27'h00000042, 5'd22, 27'h000003a0, 5'd16, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000239, 5'd23, 27'h00000393, 5'd27, 27'h000002c5, 32'h00000400,
  1'd1,  5'd1, 27'h000003bb, 5'd8, 27'h000003fe, 5'd3, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000016e, 5'd8, 27'h0000015a, 5'd10, 27'h0000018a, 32'h00000400,
  1'd1,  5'd3, 27'h00000150, 5'd9, 27'h0000038c, 5'd23, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000208, 5'd18, 27'h000002e0, 5'd3, 27'h000001ba, 32'h00000400,
  1'd1,  5'd0, 27'h000001d3, 5'd20, 27'h00000284, 5'd11, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000bd, 5'd15, 27'h00000231, 5'd25, 27'h00000348, 32'h00000400,
  1'd1,  5'd0, 27'h00000273, 5'd27, 27'h000001ab, 5'd4, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c8, 5'd29, 27'h0000003a, 5'd11, 27'h000003f0, 32'h00000400,
  1'd1,  5'd1, 27'h00000072, 5'd29, 27'h0000002e, 5'd25, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000118, 5'd7, 27'h00000177, 5'd4, 27'h000000ad, 32'h00000400,
  1'd1,  5'd11, 27'h00000304, 5'd9, 27'h000002af, 5'd13, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000e5, 5'd6, 27'h000000d9, 5'd25, 27'h000002ef, 32'h00000400,
  1'd1,  5'd13, 27'h000003b3, 5'd20, 27'h000001bb, 5'd1, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000295, 5'd19, 27'h0000007a, 5'd15, 27'h00000030, 32'h00000400,
  1'd1,  5'd10, 27'h000002a1, 5'd18, 27'h000003f9, 5'd20, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000084, 5'd30, 27'h0000030d, 5'd0, 27'h000001ed, 32'h00000400,
  1'd1,  5'd15, 27'h0000002c, 5'd30, 27'h0000022d, 5'd12, 27'h0000032c, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001ba, 5'd27, 27'h0000003d, 5'd23, 27'h00000081, 32'h00000400,
  1'd1,  5'd24, 27'h000000ad, 5'd5, 27'h0000035f, 5'd0, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000005e, 5'd6, 27'h000001ef, 5'd10, 27'h00000333, 32'h00000400,
  1'd1,  5'd24, 27'h00000159, 5'd7, 27'h00000234, 5'd21, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003bd, 5'd18, 27'h0000037a, 5'd3, 27'h00000053, 32'h00000400,
  1'd1,  5'd25, 27'h0000020c, 5'd20, 27'h000001d5, 5'd12, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000cf, 5'd17, 27'h000003de, 5'd23, 27'h000003d8, 32'h00000400,
  1'd1,  5'd23, 27'h00000056, 5'd30, 27'h00000345, 5'd0, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003df, 5'd28, 27'h00000226, 5'd12, 27'h00000077, 32'h00000400,
  1'd1,  5'd25, 27'h000001bd, 5'd28, 27'h00000342, 5'd21, 27'h0000038c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000028b, 5'd8, 27'h00000202, 5'd9, 27'h000002c3, 32'h00000400,
  1'd1,  5'd5, 27'h00000004, 5'd9, 27'h000002e7, 5'd16, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000075, 5'd8, 27'h0000035d, 5'd28, 27'h0000009f, 32'h00000400,
  1'd1,  5'd1, 27'h0000028a, 5'd18, 27'h00000041, 5'd7, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000033e, 5'd19, 27'h0000034d, 5'd18, 27'h000001d0, 32'h00000400,
  1'd1,  5'd1, 27'h00000300, 5'd18, 27'h00000129, 5'd28, 27'h00000369, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a7, 5'd30, 27'h000001d7, 5'd7, 27'h000000af, 32'h00000400,
  1'd1,  5'd5, 27'h00000091, 5'd30, 27'h00000352, 5'd17, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000000a, 5'd28, 27'h000003a4, 5'd27, 27'h00000263, 32'h00000400,
  1'd1,  5'd10, 27'h000003fc, 5'd5, 27'h000000dd, 5'd6, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000392, 5'd5, 27'h000003b0, 5'd18, 27'h00000051, 32'h00000400,
  1'd1,  5'd14, 27'h00000124, 5'd5, 27'h00000207, 5'd30, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000095, 5'd20, 27'h0000008e, 5'd9, 27'h000001b8, 32'h00000400,
  1'd1,  5'd10, 27'h000001ea, 5'd17, 27'h0000004b, 5'd17, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000395, 5'd19, 27'h00000389, 5'd27, 27'h00000062, 32'h00000400,
  1'd1,  5'd11, 27'h00000193, 5'd28, 27'h0000011c, 5'd7, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002ca, 5'd30, 27'h000003e0, 5'd15, 27'h000003d8, 32'h00000400,
  1'd1,  5'd10, 27'h000001b7, 5'd26, 27'h00000177, 5'd27, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000a9, 5'd7, 27'h000000d2, 5'd5, 27'h000001d8, 32'h00000400,
  1'd1,  5'd21, 27'h00000006, 5'd6, 27'h0000012f, 5'd19, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000bb, 5'd7, 27'h00000076, 5'd26, 27'h00000040, 32'h00000400,
  1'd1,  5'd21, 27'h00000076, 5'd17, 27'h000000c9, 5'd6, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000061, 5'd20, 27'h000001e2, 5'd20, 27'h000001fe, 32'h00000400,
  1'd1,  5'd24, 27'h00000268, 5'd16, 27'h0000023e, 5'd26, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001b, 5'd30, 27'h000003d3, 5'd8, 27'h000000ab, 32'h00000400,
  1'd1,  5'd24, 27'h000000ea, 5'd28, 27'h0000039f, 5'd19, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000010d, 5'd28, 27'h00000091, 5'd27, 27'h00000219, 32'h00000400,
  1'd1,  5'd5, 27'h00000163, 5'd4, 27'h00000047, 5'd6, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001d4, 5'd4, 27'h00000386, 5'd15, 27'h000002ac, 32'h00000400,
  1'd1,  5'd5, 27'h00000364, 5'd1, 27'h00000123, 5'd30, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000038c, 5'd11, 27'h0000021f, 5'd3, 27'h0000008a, 32'h00000400,
  1'd1,  5'd9, 27'h0000038b, 5'd12, 27'h0000008d, 5'd14, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000031c, 5'd12, 27'h0000026e, 5'd22, 27'h000001d3, 32'h00000400,
  1'd1,  5'd6, 27'h00000162, 5'd21, 27'h00000289, 5'd4, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003d8, 5'd24, 27'h00000231, 5'd15, 27'h000000ef, 32'h00000400,
  1'd1,  5'd7, 27'h00000295, 5'd21, 27'h0000032e, 5'd23, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000004d, 5'd0, 27'h0000003d, 5'd7, 27'h0000021c, 32'h00000400,
  1'd1,  5'd16, 27'h00000176, 5'd2, 27'h000002a5, 5'd19, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b7, 5'd1, 27'h000003a2, 5'd29, 27'h00000040, 32'h00000400,
  1'd1,  5'd19, 27'h000001fc, 5'd13, 27'h0000005d, 5'd4, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002d, 5'd11, 27'h00000028, 5'd12, 27'h0000015f, 32'h00000400,
  1'd1,  5'd18, 27'h00000397, 5'd15, 27'h000001a1, 5'd21, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000213, 5'd25, 27'h000000d3, 5'd4, 27'h0000034e, 32'h00000400,
  1'd1,  5'd18, 27'h0000010e, 5'd24, 27'h0000010d, 5'd13, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d7, 5'd21, 27'h000001f8, 5'd23, 27'h000003d5, 32'h00000400,
  1'd1,  5'd30, 27'h000001ac, 5'd3, 27'h00000273, 5'd4, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000267, 5'd3, 27'h0000028a, 5'd15, 27'h0000002c, 32'h00000400,
  1'd1,  5'd30, 27'h0000000d, 5'd1, 27'h000000b8, 5'd25, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000076, 5'd15, 27'h00000052, 5'd4, 27'h000001cf, 32'h00000400,
  1'd1,  5'd30, 27'h00000259, 5'd13, 27'h00000210, 5'd11, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000000c, 5'd13, 27'h00000253, 5'd21, 27'h0000036b, 32'h00000400,
  1'd1,  5'd29, 27'h00000129, 5'd23, 27'h00000044, 5'd1, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000351, 5'd25, 27'h00000089, 5'd11, 27'h00000180, 32'h00000400,
  1'd1,  5'd30, 27'h00000369, 5'd24, 27'h000002fa, 5'd24, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003ce, 5'd4, 27'h0000029c, 5'd3, 27'h0000003c, 32'h00000400,
  1'd1,  5'd9, 27'h00000318, 5'd1, 27'h0000025a, 5'd12, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000029f, 5'd1, 27'h000003cf, 5'd22, 27'h00000079, 32'h00000400,
  1'd1,  5'd8, 27'h00000341, 5'd12, 27'h000002c3, 5'd6, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002a8, 5'd10, 27'h000003cb, 5'd19, 27'h0000015a, 32'h00000400,
  1'd1,  5'd8, 27'h00000156, 5'd13, 27'h0000038c, 5'd27, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000026, 5'd25, 27'h0000030f, 5'd6, 27'h00000251, 32'h00000400,
  1'd1,  5'd9, 27'h0000039c, 5'd22, 27'h000003a0, 5'd18, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000006b, 5'd23, 27'h0000035a, 5'd27, 27'h00000086, 32'h00000400,
  1'd1,  5'd18, 27'h000001e2, 5'd2, 27'h00000337, 5'd0, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000321, 5'd4, 27'h00000141, 5'd12, 27'h0000015c, 32'h00000400,
  1'd1,  5'd19, 27'h00000270, 5'd4, 27'h0000013e, 5'd22, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003f7, 5'd10, 27'h000001ba, 5'd9, 27'h0000033c, 32'h00000400,
  1'd1,  5'd19, 27'h00000328, 5'd13, 27'h00000367, 5'd16, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000249, 5'd13, 27'h0000018b, 5'd27, 27'h000000dc, 32'h00000400,
  1'd1,  5'd16, 27'h00000325, 5'd21, 27'h000000c1, 5'd5, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000276, 5'd24, 27'h000002f1, 5'd17, 27'h00000324, 32'h00000400,
  1'd1,  5'd17, 27'h000000ba, 5'd21, 27'h0000023e, 5'd29, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001de, 5'd1, 27'h00000149, 5'd9, 27'h000000a2, 32'h00000400,
  1'd1,  5'd27, 27'h000000b1, 5'd0, 27'h000003de, 5'd17, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000292, 5'd1, 27'h00000031, 5'd30, 27'h00000294, 32'h00000400,
  1'd1,  5'd27, 27'h0000022c, 5'd11, 27'h00000022, 5'd5, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000000c, 5'd15, 27'h0000005f, 5'd18, 27'h000000b1, 32'h00000400,
  1'd1,  5'd30, 27'h00000337, 5'd12, 27'h00000072, 5'd26, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000364, 5'd24, 27'h000000bb, 5'd8, 27'h000002b2, 32'h00000400,
  1'd1,  5'd25, 27'h000003e6, 5'd24, 27'h00000244, 5'd18, 27'h000003be, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000030f, 5'd21, 27'h0000030d, 5'd28, 27'h0000007b, 32'h00000400,
  1'd1,  5'd9, 27'h000000f6, 5'd9, 27'h00000157, 5'd0, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001dd, 5'd6, 27'h00000338, 5'd12, 27'h0000013c, 32'h00000400,
  1'd1,  5'd9, 27'h000003f8, 5'd10, 27'h00000128, 5'd23, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001dc, 5'd20, 27'h00000013, 5'd2, 27'h000001cb, 32'h00000400,
  1'd1,  5'd7, 27'h000001bd, 5'd18, 27'h000000e7, 5'd12, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d9, 5'd15, 27'h0000036c, 5'd23, 27'h00000287, 32'h00000400,
  1'd1,  5'd7, 27'h000000fe, 5'd28, 27'h00000115, 5'd4, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000170, 5'd30, 27'h0000021d, 5'd11, 27'h00000357, 32'h00000400,
  1'd1,  5'd7, 27'h000003ed, 5'd30, 27'h000003fb, 5'd23, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001bc, 5'd9, 27'h0000036d, 5'd0, 27'h00000004, 32'h00000400,
  1'd1,  5'd18, 27'h00000321, 5'd7, 27'h000003dd, 5'd13, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d9, 5'd7, 27'h00000356, 5'd24, 27'h000002f6, 32'h00000400,
  1'd1,  5'd18, 27'h00000127, 5'd19, 27'h000000ae, 5'd1, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000251, 5'd19, 27'h0000019d, 5'd14, 27'h00000172, 32'h00000400,
  1'd1,  5'd20, 27'h000000e7, 5'd16, 27'h000001ad, 5'd21, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001dd, 5'd28, 27'h0000005c, 5'd1, 27'h0000005e, 32'h00000400,
  1'd1,  5'd17, 27'h00000063, 5'd26, 27'h000000c4, 5'd12, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000007c, 5'd28, 27'h000000ba, 5'd23, 27'h0000006e, 32'h00000400,
  1'd1,  5'd26, 27'h00000274, 5'd6, 27'h000000ce, 5'd0, 27'h00000204, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000085, 5'd10, 27'h000000ff, 5'd13, 27'h000002e0, 32'h00000400,
  1'd1,  5'd28, 27'h0000024c, 5'd10, 27'h00000149, 5'd21, 27'h000001e8, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000af, 5'd15, 27'h0000028a, 5'd0, 27'h00000308, 32'h00000400,
  1'd1,  5'd29, 27'h000003ae, 5'd19, 27'h0000010c, 5'd12, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001d0, 5'd16, 27'h00000351, 5'd24, 27'h0000030d, 32'h00000400,
  1'd1,  5'd26, 27'h000003a7, 5'd27, 27'h000003a8, 5'd2, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000231, 5'd27, 27'h000000d2, 5'd12, 27'h0000019f, 32'h00000400,
  1'd1,  5'd30, 27'h000000c2, 5'd27, 27'h00000095, 5'd22, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d4, 5'd7, 27'h000003ed, 5'd9, 27'h000000b8, 32'h00000400,
  1'd1,  5'd7, 27'h000001fa, 5'd6, 27'h000001a1, 5'd19, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000b5, 5'd8, 27'h00000127, 5'd28, 27'h00000193, 32'h00000400,
  1'd1,  5'd7, 27'h0000027c, 5'd17, 27'h00000191, 5'd9, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c3, 5'd19, 27'h00000107, 5'd16, 27'h000001e1, 32'h00000400,
  1'd1,  5'd10, 27'h0000013c, 5'd19, 27'h00000160, 5'd26, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001bc, 5'd30, 27'h0000035d, 5'd10, 27'h00000053, 32'h00000400,
  1'd1,  5'd8, 27'h00000393, 5'd29, 27'h0000006a, 5'd19, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003ed, 5'd27, 27'h00000076, 5'd27, 27'h0000039a, 32'h00000400,
  1'd1,  5'd16, 27'h000001f7, 5'd9, 27'h0000009b, 5'd6, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000f3, 5'd7, 27'h00000140, 5'd19, 27'h000003e2, 32'h00000400,
  1'd1,  5'd15, 27'h000002ec, 5'd5, 27'h00000316, 5'd29, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002b7, 5'd17, 27'h000002c4, 5'd9, 27'h00000090, 32'h00000400,
  1'd1,  5'd19, 27'h00000160, 5'd16, 27'h000001f2, 5'd15, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000039, 5'd18, 27'h00000320, 5'd25, 27'h00000365, 32'h00000400,
  1'd1,  5'd19, 27'h0000024c, 5'd27, 27'h00000196, 5'd5, 27'h00000346, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b9, 5'd27, 27'h00000087, 5'd16, 27'h00000203, 32'h00000400,
  1'd1,  5'd17, 27'h00000380, 5'd30, 27'h00000027, 5'd30, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000b2, 5'd7, 27'h000003b2, 5'd9, 27'h000003cb, 32'h00000400,
  1'd1,  5'd28, 27'h000003c2, 5'd7, 27'h00000158, 5'd18, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002c5, 5'd5, 27'h0000026c, 5'd26, 27'h000002f6, 32'h00000400,
  1'd1,  5'd26, 27'h00000341, 5'd16, 27'h0000009b, 5'd10, 27'h0000003f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000195, 5'd18, 27'h0000026a, 5'd19, 27'h00000183, 32'h00000400,
  1'd1,  5'd26, 27'h000000d3, 5'd16, 27'h000000be, 5'd30, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000165, 5'd26, 27'h00000290, 5'd7, 27'h0000019b, 32'h00000400,
  1'd1,  5'd26, 27'h0000009c, 5'd26, 27'h000000fc, 5'd16, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b8, 5'd28, 27'h00000318, 5'd28, 27'h0000030a, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000383, 5'd0, 27'h0000026b, 5'd4, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002c7, 5'd4, 27'h000003f5, 5'd12, 27'h00000207, 32'h00000400,
  1'd1,  5'd3, 27'h0000036f, 5'd2, 27'h000000ba, 5'd20, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000326, 5'd15, 27'h00000159, 5'd2, 27'h00000096, 32'h00000400,
  1'd1,  5'd0, 27'h0000005c, 5'd14, 27'h0000022c, 5'd10, 27'h00000162, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000319, 5'd11, 27'h000002aa, 5'd22, 27'h00000289, 32'h00000400,
  1'd1,  5'd0, 27'h00000038, 5'd25, 27'h00000032, 5'd4, 27'h000001cb, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000029, 5'd20, 27'h000003c2, 5'd11, 27'h00000045, 32'h00000400,
  1'd1,  5'd4, 27'h000002b3, 5'd25, 27'h0000007f, 5'd21, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c1, 5'd0, 27'h00000383, 5'd2, 27'h0000016c, 32'h00000400,
  1'd1,  5'd13, 27'h000000ad, 5'd0, 27'h00000110, 5'd14, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001a6, 5'd2, 27'h000002d0, 5'd24, 27'h00000011, 32'h00000400,
  1'd1,  5'd13, 27'h00000242, 5'd12, 27'h000001e1, 5'd4, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000256, 5'd14, 27'h0000036d, 5'd11, 27'h00000209, 32'h00000400,
  1'd1,  5'd15, 27'h000000a7, 5'd10, 27'h0000039f, 5'd21, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000388, 5'd24, 27'h00000390, 5'd1, 27'h000003ec, 32'h00000400,
  1'd1,  5'd12, 27'h000003ed, 5'd24, 27'h0000021b, 5'd14, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000022d, 5'd21, 27'h00000123, 5'd25, 27'h000001ef, 32'h00000400,
  1'd1,  5'd25, 27'h00000144, 5'd4, 27'h000003c9, 5'd4, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ae, 5'd3, 27'h0000004b, 5'd13, 27'h000002f0, 32'h00000400,
  1'd1,  5'd25, 27'h00000102, 5'd4, 27'h000000ea, 5'd25, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e3, 5'd13, 27'h000002b2, 5'd0, 27'h000003bc, 32'h00000400,
  1'd1,  5'd25, 27'h000001c9, 5'd13, 27'h00000324, 5'd15, 27'h000000ae, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000138, 5'd12, 27'h0000016b, 5'd22, 27'h0000025c, 32'h00000400,
  1'd1,  5'd22, 27'h000003fa, 5'd21, 27'h00000221, 5'd3, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000c3, 5'd24, 27'h00000111, 5'd13, 27'h000002e4, 32'h00000400,
  1'd1,  5'd24, 27'h00000396, 5'd24, 27'h0000038e, 5'd23, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002a7, 5'd0, 27'h00000143, 5'd5, 27'h000002d5, 32'h00000400,
  1'd1,  5'd4, 27'h0000002c, 5'd3, 27'h0000032f, 5'd17, 27'h0000003c, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028c, 5'd1, 27'h000002c4, 5'd30, 27'h000002d8, 32'h00000400,
  1'd1,  5'd1, 27'h000002e6, 5'd15, 27'h00000119, 5'd9, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000033e, 5'd13, 27'h000001b9, 5'd17, 27'h000000e4, 32'h00000400,
  1'd1,  5'd2, 27'h000000d7, 5'd10, 27'h0000031f, 5'd28, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002f9, 5'd22, 27'h00000170, 5'd8, 27'h0000000d, 32'h00000400,
  1'd1,  5'd1, 27'h00000105, 5'd24, 27'h000000af, 5'd15, 27'h00000318, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ea, 5'd23, 27'h0000025c, 5'd29, 27'h00000244, 32'h00000400,
  1'd1,  5'd14, 27'h00000262, 5'd4, 27'h0000022c, 5'd7, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003e8, 5'd3, 27'h00000040, 5'd17, 27'h00000174, 32'h00000400,
  1'd1,  5'd13, 27'h00000269, 5'd0, 27'h00000008, 5'd29, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f7, 5'd12, 27'h000002a4, 5'd6, 27'h00000086, 32'h00000400,
  1'd1,  5'd13, 27'h00000048, 5'd14, 27'h000003e7, 5'd17, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000a7, 5'd10, 27'h000002a8, 5'd26, 27'h0000030e, 32'h00000400,
  1'd1,  5'd13, 27'h000002c6, 5'd24, 27'h00000315, 5'd9, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ea, 5'd20, 27'h000002ac, 5'd16, 27'h00000147, 32'h00000400,
  1'd1,  5'd11, 27'h000000c3, 5'd22, 27'h00000103, 5'd30, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001b6, 5'd0, 27'h00000326, 5'd9, 27'h00000311, 32'h00000400,
  1'd1,  5'd21, 27'h00000000, 5'd1, 27'h00000377, 5'd16, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000013f, 5'd1, 27'h000003b1, 5'd28, 27'h000002fa, 32'h00000400,
  1'd1,  5'd22, 27'h000002c8, 5'd13, 27'h0000025b, 5'd6, 27'h000001c4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000051, 5'd12, 27'h000000c1, 5'd19, 27'h00000231, 32'h00000400,
  1'd1,  5'd24, 27'h000002bf, 5'd15, 27'h000000d4, 5'd28, 27'h0000034e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000099, 5'd21, 27'h000000ca, 5'd8, 27'h0000029f, 32'h00000400,
  1'd1,  5'd22, 27'h000002e2, 5'd24, 27'h00000024, 5'd19, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000337, 5'd22, 27'h00000088, 5'd28, 27'h000002f7, 32'h00000400,
  1'd1,  5'd3, 27'h000003c9, 5'd7, 27'h00000195, 5'd1, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002cd, 5'd8, 27'h000003e4, 5'd12, 27'h00000331, 32'h00000400,
  1'd1,  5'd0, 27'h0000031e, 5'd10, 27'h0000000b, 5'd24, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e9, 5'd19, 27'h00000056, 5'd1, 27'h0000002a, 32'h00000400,
  1'd1,  5'd1, 27'h00000213, 5'd20, 27'h0000011a, 5'd14, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000007b, 5'd16, 27'h00000221, 5'd23, 27'h00000349, 32'h00000400,
  1'd1,  5'd0, 27'h000000b1, 5'd28, 27'h000002c1, 5'd3, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003bc, 5'd28, 27'h00000311, 5'd10, 27'h000002c7, 32'h00000400,
  1'd1,  5'd0, 27'h000003cb, 5'd28, 27'h000001c9, 5'd22, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003e8, 5'd9, 27'h00000023, 5'd0, 27'h000002d1, 32'h00000400,
  1'd1,  5'd11, 27'h000002d0, 5'd9, 27'h0000033b, 5'd10, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003f9, 5'd7, 27'h00000290, 5'd22, 27'h00000018, 32'h00000400,
  1'd1,  5'd11, 27'h000003f8, 5'd20, 27'h00000028, 5'd3, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000001b, 5'd19, 27'h00000307, 5'd15, 27'h000001b7, 32'h00000400,
  1'd1,  5'd10, 27'h000001e0, 5'd17, 27'h000001be, 5'd21, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000031b, 5'd26, 27'h000003fe, 5'd1, 27'h00000133, 32'h00000400,
  1'd1,  5'd14, 27'h000000de, 5'd29, 27'h00000112, 5'd14, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018b, 5'd27, 27'h000003b6, 5'd22, 27'h0000029d, 32'h00000400,
  1'd1,  5'd25, 27'h00000229, 5'd9, 27'h000001d7, 5'd2, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000001a, 5'd7, 27'h00000370, 5'd15, 27'h000000a7, 32'h00000400,
  1'd1,  5'd22, 27'h00000322, 5'd7, 27'h0000011e, 5'd22, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000021d, 5'd16, 27'h00000374, 5'd0, 27'h000003ca, 32'h00000400,
  1'd1,  5'd22, 27'h00000299, 5'd17, 27'h00000111, 5'd12, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000102, 5'd17, 27'h000000d6, 5'd25, 27'h00000115, 32'h00000400,
  1'd1,  5'd24, 27'h000002cb, 5'd26, 27'h000002a5, 5'd4, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003eb, 5'd26, 27'h000000b2, 5'd11, 27'h00000371, 32'h00000400,
  1'd1,  5'd24, 27'h000002f4, 5'd27, 27'h0000018f, 5'd22, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002bb, 5'd6, 27'h00000024, 5'd9, 27'h00000291, 32'h00000400,
  1'd1,  5'd3, 27'h000003c2, 5'd6, 27'h00000108, 5'd18, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003ce, 5'd6, 27'h0000019c, 5'd29, 27'h000002cd, 32'h00000400,
  1'd1,  5'd0, 27'h0000038c, 5'd17, 27'h00000123, 5'd10, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000365, 5'd18, 27'h000001c9, 5'd17, 27'h00000019, 32'h00000400,
  1'd1,  5'd0, 27'h0000031f, 5'd16, 27'h000001e6, 5'd26, 27'h000003de, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000397, 5'd29, 27'h0000027f, 5'd9, 27'h00000375, 32'h00000400,
  1'd1,  5'd0, 27'h00000296, 5'd29, 27'h0000017e, 5'd16, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000004e, 5'd30, 27'h000001a7, 5'd29, 27'h000000ef, 32'h00000400,
  1'd1,  5'd14, 27'h000001cc, 5'd8, 27'h0000015f, 5'd8, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000166, 5'd7, 27'h00000287, 5'd18, 27'h000000ef, 32'h00000400,
  1'd1,  5'd10, 27'h000001db, 5'd7, 27'h00000166, 5'd26, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000221, 5'd18, 27'h00000240, 5'd9, 27'h00000310, 32'h00000400,
  1'd1,  5'd14, 27'h00000226, 5'd15, 27'h000003e9, 5'd15, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000034b, 5'd16, 27'h0000008e, 5'd26, 27'h00000015, 32'h00000400,
  1'd1,  5'd11, 27'h000000ec, 5'd29, 27'h0000020e, 5'd6, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000312, 5'd29, 27'h000001d5, 5'd19, 27'h00000307, 32'h00000400,
  1'd1,  5'd13, 27'h000000c5, 5'd30, 27'h00000339, 5'd29, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000038c, 5'd9, 27'h00000038, 5'd7, 27'h000000f4, 32'h00000400,
  1'd1,  5'd22, 27'h000000a5, 5'd8, 27'h0000031f, 5'd16, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000284, 5'd6, 27'h0000020a, 5'd26, 27'h00000197, 32'h00000400,
  1'd1,  5'd25, 27'h0000003c, 5'd18, 27'h00000010, 5'd7, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a1, 5'd18, 27'h00000186, 5'd17, 27'h000002e6, 32'h00000400,
  1'd1,  5'd23, 27'h0000010b, 5'd18, 27'h000003fb, 5'd28, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f6, 5'd26, 27'h0000015d, 5'd6, 27'h0000004c, 32'h00000400,
  1'd1,  5'd22, 27'h000001b2, 5'd30, 27'h000002a9, 5'd16, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001b6, 5'd29, 27'h00000031, 5'd28, 27'h000003b4, 32'h00000400,
  1'd1,  5'd9, 27'h00000147, 5'd0, 27'h0000010f, 5'd6, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000014, 5'd4, 27'h0000020c, 5'd15, 27'h000002f4, 32'h00000400,
  1'd1,  5'd8, 27'h0000002b, 5'd4, 27'h00000386, 5'd26, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001f5, 5'd10, 27'h00000226, 5'd2, 27'h00000063, 32'h00000400,
  1'd1,  5'd9, 27'h00000265, 5'd13, 27'h00000293, 5'd12, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000034d, 5'd10, 27'h00000384, 5'd24, 27'h000001e1, 32'h00000400,
  1'd1,  5'd7, 27'h0000039b, 5'd24, 27'h00000367, 5'd3, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003dd, 5'd21, 27'h0000033c, 5'd12, 27'h00000287, 32'h00000400,
  1'd1,  5'd6, 27'h000000a8, 5'd21, 27'h00000204, 5'd24, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000199, 5'd5, 27'h0000002f, 5'd7, 27'h000003c4, 32'h00000400,
  1'd1,  5'd19, 27'h00000210, 5'd4, 27'h00000251, 5'd18, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002cb, 5'd2, 27'h000000ff, 5'd27, 27'h000002ea, 32'h00000400,
  1'd1,  5'd20, 27'h00000196, 5'd12, 27'h0000025d, 5'd1, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c3, 5'd11, 27'h000003b6, 5'd10, 27'h000002bf, 32'h00000400,
  1'd1,  5'd16, 27'h000003ec, 5'd11, 27'h00000008, 5'd25, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000f0, 5'd23, 27'h00000328, 5'd4, 27'h000001cc, 32'h00000400,
  1'd1,  5'd16, 27'h0000011a, 5'd25, 27'h00000202, 5'd12, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000037e, 5'd21, 27'h0000037c, 5'd25, 27'h00000143, 32'h00000400,
  1'd1,  5'd28, 27'h000003bf, 5'd1, 27'h00000165, 5'd0, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b5, 5'd0, 27'h0000019f, 5'd11, 27'h0000038b, 32'h00000400,
  1'd1,  5'd27, 27'h000003c7, 5'd5, 27'h0000001d, 5'd24, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002d3, 5'd10, 27'h00000307, 5'd4, 27'h00000202, 32'h00000400,
  1'd1,  5'd28, 27'h000000d2, 5'd14, 27'h00000393, 5'd13, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000037b, 5'd13, 27'h0000030a, 5'd24, 27'h00000207, 32'h00000400,
  1'd1,  5'd27, 27'h00000171, 5'd22, 27'h000001c5, 5'd3, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000100, 5'd24, 27'h000002b8, 5'd12, 27'h000000ed, 32'h00000400,
  1'd1,  5'd27, 27'h00000134, 5'd22, 27'h00000125, 5'd23, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003ef, 5'd0, 27'h000002a3, 5'd1, 27'h00000322, 32'h00000400,
  1'd1,  5'd5, 27'h00000113, 5'd2, 27'h00000161, 5'd11, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000215, 5'd1, 27'h00000075, 5'd21, 27'h00000057, 32'h00000400,
  1'd1,  5'd9, 27'h0000027b, 5'd13, 27'h00000200, 5'd9, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001e7, 5'd14, 27'h0000018f, 5'd18, 27'h00000187, 32'h00000400,
  1'd1,  5'd6, 27'h0000016f, 5'd10, 27'h00000249, 5'd27, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000197, 5'd23, 27'h00000173, 5'd9, 27'h000001cb, 32'h00000400,
  1'd1,  5'd9, 27'h00000156, 5'd21, 27'h000002e8, 5'd20, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000124, 5'd24, 27'h0000002d, 5'd26, 27'h0000015e, 32'h00000400,
  1'd1,  5'd17, 27'h0000033b, 5'd0, 27'h000003a3, 5'd1, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000010c, 5'd4, 27'h0000011d, 5'd11, 27'h000002ac, 32'h00000400,
  1'd1,  5'd15, 27'h00000388, 5'd0, 27'h0000022a, 5'd21, 27'h000001b2, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000299, 5'd13, 27'h00000081, 5'd6, 27'h00000036, 32'h00000400,
  1'd1,  5'd17, 27'h0000011b, 5'd14, 27'h0000016b, 5'd20, 27'h0000013b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000264, 5'd11, 27'h00000137, 5'd30, 27'h0000003a, 32'h00000400,
  1'd1,  5'd17, 27'h000002a1, 5'd20, 27'h000003de, 5'd5, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000305, 5'd22, 27'h00000389, 5'd17, 27'h00000300, 32'h00000400,
  1'd1,  5'd15, 27'h000002b9, 5'd22, 27'h00000251, 5'd30, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000022a, 5'd3, 27'h000000f2, 5'd6, 27'h0000008e, 32'h00000400,
  1'd1,  5'd30, 27'h000000f7, 5'd0, 27'h00000331, 5'd15, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003cc, 5'd3, 27'h00000284, 5'd30, 27'h00000149, 32'h00000400,
  1'd1,  5'd29, 27'h0000009b, 5'd13, 27'h000003b7, 5'd6, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000002f, 5'd12, 27'h000002e7, 5'd19, 27'h00000015, 32'h00000400,
  1'd1,  5'd29, 27'h000001f9, 5'd12, 27'h0000026e, 5'd26, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000d9, 5'd24, 27'h00000294, 5'd6, 27'h0000012c, 32'h00000400,
  1'd1,  5'd28, 27'h0000021a, 5'd23, 27'h0000030c, 5'd17, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f6, 5'd24, 27'h000003e3, 5'd28, 27'h000000b5, 32'h00000400,
  1'd1,  5'd8, 27'h00000049, 5'd6, 27'h0000017f, 5'd0, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000223, 5'd8, 27'h00000366, 5'd12, 27'h00000108, 32'h00000400,
  1'd1,  5'd5, 27'h000001cb, 5'd7, 27'h000001a0, 5'd21, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000014f, 5'd17, 27'h00000400, 5'd0, 27'h0000002b, 32'h00000400,
  1'd1,  5'd5, 27'h000001e9, 5'd20, 27'h0000002b, 5'd13, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003dc, 5'd20, 27'h00000266, 5'd23, 27'h0000001a, 32'h00000400,
  1'd1,  5'd9, 27'h0000035d, 5'd26, 27'h0000024a, 5'd4, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000015b, 5'd30, 27'h0000023b, 5'd15, 27'h0000014b, 32'h00000400,
  1'd1,  5'd6, 27'h000001ec, 5'd26, 27'h00000387, 5'd22, 27'h00000383, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002d2, 5'd8, 27'h000001d3, 5'd4, 27'h000000cf, 32'h00000400,
  1'd1,  5'd17, 27'h000000c8, 5'd9, 27'h00000167, 5'd14, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000279, 5'd9, 27'h000003d1, 5'd25, 27'h00000045, 32'h00000400,
  1'd1,  5'd19, 27'h00000345, 5'd18, 27'h000000cd, 5'd2, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000002, 5'd20, 27'h00000238, 5'd10, 27'h00000299, 32'h00000400,
  1'd1,  5'd17, 27'h00000072, 5'd17, 27'h00000191, 5'd22, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001fc, 5'd30, 27'h00000172, 5'd2, 27'h00000025, 32'h00000400,
  1'd1,  5'd17, 27'h00000049, 5'd28, 27'h000000dd, 5'd14, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000be, 5'd27, 27'h00000320, 5'd23, 27'h0000025b, 32'h00000400,
  1'd1,  5'd28, 27'h000002cc, 5'd5, 27'h0000012d, 5'd1, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000147, 5'd8, 27'h00000253, 5'd13, 27'h000000fc, 32'h00000400,
  1'd1,  5'd27, 27'h0000020b, 5'd5, 27'h0000022c, 5'd20, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000316, 5'd19, 27'h000002f9, 5'd1, 27'h000002aa, 32'h00000400,
  1'd1,  5'd27, 27'h000003cb, 5'd19, 27'h000002ca, 5'd13, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003d8, 5'd16, 27'h000001a6, 5'd21, 27'h00000088, 32'h00000400,
  1'd1,  5'd28, 27'h0000005d, 5'd28, 27'h00000215, 5'd1, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024a, 5'd26, 27'h00000330, 5'd13, 27'h000003c4, 32'h00000400,
  1'd1,  5'd26, 27'h00000379, 5'd28, 27'h00000277, 5'd24, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000373, 5'd6, 27'h0000002b, 5'd5, 27'h00000186, 32'h00000400,
  1'd1,  5'd9, 27'h000002b6, 5'd6, 27'h00000325, 5'd17, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000399, 5'd6, 27'h00000358, 5'd25, 27'h0000035e, 32'h00000400,
  1'd1,  5'd6, 27'h00000356, 5'd19, 27'h000000be, 5'd8, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000010d, 5'd17, 27'h000003ad, 5'd19, 27'h00000082, 32'h00000400,
  1'd1,  5'd8, 27'h000003c2, 5'd16, 27'h000001ad, 5'd30, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000005, 5'd30, 27'h00000099, 5'd9, 27'h00000359, 32'h00000400,
  1'd1,  5'd7, 27'h0000025a, 5'd26, 27'h000001ad, 5'd18, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000042, 5'd27, 27'h0000013c, 5'd29, 27'h00000083, 32'h00000400,
  1'd1,  5'd15, 27'h000002d1, 5'd9, 27'h0000014e, 5'd10, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000302, 5'd8, 27'h00000334, 5'd19, 27'h0000001e, 32'h00000400,
  1'd1,  5'd18, 27'h0000020f, 5'd7, 27'h000002b8, 5'd27, 27'h000002de, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000bd, 5'd18, 27'h00000027, 5'd8, 27'h00000305, 32'h00000400,
  1'd1,  5'd16, 27'h000003dd, 5'd20, 27'h0000025a, 5'd20, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a1, 5'd17, 27'h000002b5, 5'd29, 27'h00000036, 32'h00000400,
  1'd1,  5'd16, 27'h000003b8, 5'd26, 27'h00000238, 5'd8, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000062, 5'd27, 27'h000001c6, 5'd16, 27'h00000087, 32'h00000400,
  1'd1,  5'd19, 27'h00000210, 5'd28, 27'h0000011a, 5'd28, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000011, 5'd9, 27'h00000303, 5'd6, 27'h00000203, 32'h00000400,
  1'd1,  5'd26, 27'h00000258, 5'd7, 27'h00000122, 5'd19, 27'h00000015, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002cd, 5'd8, 27'h000003f5, 5'd25, 27'h000003b1, 32'h00000400,
  1'd1,  5'd30, 27'h000002fd, 5'd16, 27'h000003e9, 5'd9, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000315, 5'd15, 27'h000003ae, 5'd18, 27'h000001ec, 32'h00000400,
  1'd1,  5'd29, 27'h00000303, 5'd16, 27'h0000026e, 5'd29, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001be, 5'd28, 27'h000003c5, 5'd10, 27'h00000010, 32'h00000400,
  1'd1,  5'd30, 27'h0000028c, 5'd27, 27'h000000e6, 5'd17, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b0, 5'd26, 27'h000002b2, 5'd27, 27'h000003bd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001cc, 5'd2, 27'h000001be, 5'd1, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003bf, 5'd0, 27'h000002ce, 5'd11, 27'h00000281, 32'h00000400,
  1'd1,  5'd1, 27'h00000201, 5'd3, 27'h000000c7, 5'd23, 27'h00000091, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000207, 5'd13, 27'h0000014f, 5'd3, 27'h0000038c, 32'h00000400,
  1'd1,  5'd2, 27'h00000230, 5'd11, 27'h0000015d, 5'd13, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b0, 5'd10, 27'h00000198, 5'd20, 27'h000002de, 32'h00000400,
  1'd1,  5'd2, 27'h000001be, 5'd22, 27'h000000ec, 5'd5, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003fe, 5'd24, 27'h0000007c, 5'd10, 27'h0000018e, 32'h00000400,
  1'd1,  5'd2, 27'h00000394, 5'd22, 27'h00000218, 5'd20, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000016f, 5'd0, 27'h00000332, 5'd1, 27'h000003c1, 32'h00000400,
  1'd1,  5'd11, 27'h0000012d, 5'd1, 27'h000002d1, 5'd12, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000377, 5'd3, 27'h000000b2, 5'd22, 27'h00000082, 32'h00000400,
  1'd1,  5'd11, 27'h00000193, 5'd13, 27'h00000045, 5'd2, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000175, 5'd12, 27'h00000396, 5'd12, 27'h0000032f, 32'h00000400,
  1'd1,  5'd11, 27'h000003a9, 5'd15, 27'h0000017c, 5'd23, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003cd, 5'd22, 27'h00000271, 5'd4, 27'h000001ec, 32'h00000400,
  1'd1,  5'd14, 27'h0000005a, 5'd20, 27'h000002ac, 5'd10, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000023d, 5'd24, 27'h0000026a, 5'd22, 27'h00000349, 32'h00000400,
  1'd1,  5'd23, 27'h000000b7, 5'd5, 27'h000000a6, 5'd2, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002c5, 5'd2, 27'h00000350, 5'd13, 27'h000000da, 32'h00000400,
  1'd1,  5'd25, 27'h0000027b, 5'd4, 27'h00000106, 5'd21, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000005e, 5'd12, 27'h000002fe, 5'd2, 27'h00000206, 32'h00000400,
  1'd1,  5'd21, 27'h000001d3, 5'd12, 27'h00000123, 5'd12, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000325, 5'd13, 27'h0000004d, 5'd20, 27'h000002e7, 32'h00000400,
  1'd1,  5'd24, 27'h00000015, 5'd24, 27'h00000284, 5'd1, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f9, 5'd23, 27'h0000018a, 5'd12, 27'h00000385, 32'h00000400,
  1'd1,  5'd20, 27'h000003fd, 5'd21, 27'h00000239, 5'd23, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001eb, 5'd0, 27'h000002b3, 5'd7, 27'h00000021, 32'h00000400,
  1'd1,  5'd4, 27'h00000005, 5'd0, 27'h00000208, 5'd16, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003f9, 5'd0, 27'h000001e6, 5'd29, 27'h00000067, 32'h00000400,
  1'd1,  5'd0, 27'h00000318, 5'd14, 27'h000000c7, 5'd10, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003a0, 5'd15, 27'h000000ab, 5'd20, 27'h0000004c, 32'h00000400,
  1'd1,  5'd3, 27'h0000023d, 5'd15, 27'h00000136, 5'd26, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000002a, 5'd22, 27'h0000008c, 5'd8, 27'h00000292, 32'h00000400,
  1'd1,  5'd0, 27'h00000155, 5'd25, 27'h00000236, 5'd16, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000028c, 5'd21, 27'h00000031, 5'd28, 27'h00000082, 32'h00000400,
  1'd1,  5'd11, 27'h0000025b, 5'd2, 27'h00000011, 5'd10, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000264, 5'd4, 27'h00000198, 5'd15, 27'h00000224, 32'h00000400,
  1'd1,  5'd14, 27'h000003ed, 5'd0, 27'h0000000c, 5'd27, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000360, 5'd12, 27'h000003ad, 5'd8, 27'h0000000c, 32'h00000400,
  1'd1,  5'd11, 27'h00000223, 5'd11, 27'h00000329, 5'd17, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000012d, 5'd14, 27'h00000130, 5'd30, 27'h00000344, 32'h00000400,
  1'd1,  5'd15, 27'h000001a3, 5'd24, 27'h000001f4, 5'd8, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000026c, 5'd22, 27'h000003a6, 5'd20, 27'h000001bb, 32'h00000400,
  1'd1,  5'd14, 27'h00000054, 5'd24, 27'h0000029a, 5'd28, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022b, 5'd2, 27'h00000033, 5'd7, 27'h0000031d, 32'h00000400,
  1'd1,  5'd22, 27'h0000035c, 5'd0, 27'h0000029e, 5'd17, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d2, 5'd2, 27'h000002d9, 5'd27, 27'h000000b4, 32'h00000400,
  1'd1,  5'd23, 27'h000002b4, 5'd15, 27'h0000008f, 5'd10, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000020f, 5'd11, 27'h000001bf, 5'd16, 27'h00000325, 32'h00000400,
  1'd1,  5'd21, 27'h00000013, 5'd12, 27'h00000035, 5'd28, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000190, 5'd25, 27'h0000004a, 5'd5, 27'h00000272, 32'h00000400,
  1'd1,  5'd21, 27'h000000a5, 5'd22, 27'h000002b3, 5'd18, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000103, 5'd23, 27'h00000317, 5'd27, 27'h000000c5, 32'h00000400,
  1'd1,  5'd4, 27'h00000131, 5'd7, 27'h00000144, 5'd3, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000232, 5'd7, 27'h00000350, 5'd10, 27'h00000336, 32'h00000400,
  1'd1,  5'd3, 27'h0000006a, 5'd6, 27'h00000265, 5'd23, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ee, 5'd19, 27'h00000372, 5'd3, 27'h000001b9, 32'h00000400,
  1'd1,  5'd0, 27'h0000026e, 5'd16, 27'h000000da, 5'd15, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000029e, 5'd17, 27'h0000029d, 5'd24, 27'h00000074, 32'h00000400,
  1'd1,  5'd2, 27'h00000155, 5'd29, 27'h000002f4, 5'd0, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003c6, 5'd28, 27'h00000190, 5'd12, 27'h0000037f, 32'h00000400,
  1'd1,  5'd5, 27'h0000009c, 5'd29, 27'h0000030d, 5'd23, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000054, 5'd8, 27'h000001fc, 5'd1, 27'h000002b9, 32'h00000400,
  1'd1,  5'd11, 27'h000000df, 5'd8, 27'h00000273, 5'd12, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a5, 5'd5, 27'h0000017c, 5'd21, 27'h000000a9, 32'h00000400,
  1'd1,  5'd15, 27'h00000060, 5'd15, 27'h0000032b, 5'd2, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000011c, 5'd20, 27'h00000189, 5'd13, 27'h00000282, 32'h00000400,
  1'd1,  5'd10, 27'h00000389, 5'd20, 27'h000000be, 5'd23, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd10, 27'h000003b3, 5'd28, 27'h00000029, 5'd4, 27'h0000018f, 32'h00000400,
  1'd1,  5'd13, 27'h000002d1, 5'd29, 27'h000002fc, 5'd10, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001bd, 5'd27, 27'h000001bd, 5'd21, 27'h00000280, 32'h00000400,
  1'd1,  5'd23, 27'h000001a7, 5'd5, 27'h000000d0, 5'd0, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000002b, 5'd8, 27'h00000340, 5'd13, 27'h0000028d, 32'h00000400,
  1'd1,  5'd20, 27'h0000034e, 5'd8, 27'h000003d8, 5'd20, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002af, 5'd18, 27'h0000018a, 5'd0, 27'h00000375, 32'h00000400,
  1'd1,  5'd23, 27'h000003ad, 5'd19, 27'h0000037e, 5'd10, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000211, 5'd18, 27'h000000ad, 5'd23, 27'h00000360, 32'h00000400,
  1'd1,  5'd24, 27'h000003a9, 5'd27, 27'h0000001d, 5'd4, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000031f, 5'd27, 27'h00000053, 5'd11, 27'h00000004, 32'h00000400,
  1'd1,  5'd22, 27'h0000015d, 5'd25, 27'h000003a2, 5'd23, 27'h00000040, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000350, 5'd5, 27'h000000d8, 5'd7, 27'h000000c4, 32'h00000400,
  1'd1,  5'd4, 27'h00000246, 5'd9, 27'h00000323, 5'd18, 27'h000000ad, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000177, 5'd7, 27'h00000180, 5'd30, 27'h000000c5, 32'h00000400,
  1'd1,  5'd3, 27'h0000015a, 5'd18, 27'h00000049, 5'd9, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000027, 5'd18, 27'h000003f3, 5'd18, 27'h000001f1, 32'h00000400,
  1'd1,  5'd1, 27'h00000272, 5'd16, 27'h000000bb, 5'd28, 27'h00000186, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000020a, 5'd28, 27'h000000b2, 5'd8, 27'h000003bb, 32'h00000400,
  1'd1,  5'd3, 27'h0000009d, 5'd30, 27'h0000018a, 5'd19, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ae, 5'd30, 27'h00000202, 5'd26, 27'h000001b7, 32'h00000400,
  1'd1,  5'd14, 27'h00000297, 5'd8, 27'h00000051, 5'd8, 27'h0000000f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f6, 5'd10, 27'h000000a9, 5'd20, 27'h00000162, 32'h00000400,
  1'd1,  5'd13, 27'h0000020a, 5'd5, 27'h0000034f, 5'd27, 27'h0000016d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c0, 5'd18, 27'h00000368, 5'd6, 27'h00000214, 32'h00000400,
  1'd1,  5'd10, 27'h000002f8, 5'd17, 27'h0000018b, 5'd16, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003fb, 5'd16, 27'h0000023d, 5'd28, 27'h0000012f, 32'h00000400,
  1'd1,  5'd15, 27'h00000141, 5'd27, 27'h00000034, 5'd7, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ab, 5'd26, 27'h0000008e, 5'd18, 27'h000003d6, 32'h00000400,
  1'd1,  5'd10, 27'h00000314, 5'd25, 27'h000003f9, 5'd30, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000cd, 5'd8, 27'h000000ce, 5'd5, 27'h000000e2, 32'h00000400,
  1'd1,  5'd24, 27'h000002b7, 5'd6, 27'h00000067, 5'd18, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000fe, 5'd9, 27'h00000032, 5'd28, 27'h0000002e, 32'h00000400,
  1'd1,  5'd24, 27'h000001ac, 5'd19, 27'h00000389, 5'd5, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000022b, 5'd18, 27'h0000037d, 5'd16, 27'h00000076, 32'h00000400,
  1'd1,  5'd22, 27'h00000399, 5'd17, 27'h00000115, 5'd28, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bd, 5'd28, 27'h000001e0, 5'd6, 27'h0000031f, 32'h00000400,
  1'd1,  5'd20, 27'h000002fb, 5'd30, 27'h00000052, 5'd19, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a5, 5'd30, 27'h00000165, 5'd30, 27'h00000224, 32'h00000400,
  1'd1,  5'd5, 27'h0000011b, 5'd0, 27'h00000334, 5'd6, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003eb, 5'd2, 27'h000001d2, 5'd18, 27'h000000cc, 32'h00000400,
  1'd1,  5'd10, 27'h00000120, 5'd1, 27'h0000022a, 5'd27, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000234, 5'd11, 27'h0000017e, 5'd3, 27'h0000009e, 32'h00000400,
  1'd1,  5'd5, 27'h000000d0, 5'd14, 27'h0000023d, 5'd15, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002ea, 5'd11, 27'h000000c3, 5'd24, 27'h00000012, 32'h00000400,
  1'd1,  5'd6, 27'h0000010b, 5'd22, 27'h00000247, 5'd4, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003b4, 5'd23, 27'h000003de, 5'd10, 27'h0000039b, 32'h00000400,
  1'd1,  5'd7, 27'h00000293, 5'd24, 27'h00000220, 5'd23, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000e2, 5'd4, 27'h00000336, 5'd9, 27'h000001e1, 32'h00000400,
  1'd1,  5'd17, 27'h00000206, 5'd1, 27'h000003c7, 5'd16, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ed, 5'd1, 27'h000001c2, 5'd26, 27'h00000114, 32'h00000400,
  1'd1,  5'd18, 27'h00000084, 5'd11, 27'h00000182, 5'd1, 27'h00000262, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000347, 5'd12, 27'h0000018f, 5'd11, 27'h000003ce, 32'h00000400,
  1'd1,  5'd20, 27'h00000086, 5'd14, 27'h000002ab, 5'd20, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000068, 5'd21, 27'h0000036c, 5'd3, 27'h000001b6, 32'h00000400,
  1'd1,  5'd19, 27'h00000185, 5'd22, 27'h0000007d, 5'd10, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000020a, 5'd24, 27'h000000d5, 5'd21, 27'h00000346, 32'h00000400,
  1'd1,  5'd30, 27'h00000387, 5'd2, 27'h00000157, 5'd3, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002d1, 5'd0, 27'h0000021d, 5'd13, 27'h0000036a, 32'h00000400,
  1'd1,  5'd29, 27'h000003fd, 5'd2, 27'h00000366, 5'd23, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001a5, 5'd14, 27'h00000363, 5'd4, 27'h000003ce, 32'h00000400,
  1'd1,  5'd30, 27'h0000007c, 5'd15, 27'h0000018b, 5'd13, 27'h000003fa, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000c0, 5'd12, 27'h00000063, 5'd23, 27'h000000c9, 32'h00000400,
  1'd1,  5'd29, 27'h000002bb, 5'd22, 27'h00000047, 5'd3, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000114, 5'd24, 27'h000001c8, 5'd11, 27'h00000109, 32'h00000400,
  1'd1,  5'd30, 27'h0000008a, 5'd21, 27'h00000004, 5'd22, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000201, 5'd4, 27'h00000116, 5'd2, 27'h00000382, 32'h00000400,
  1'd1,  5'd7, 27'h000003a1, 5'd3, 27'h000001f3, 5'd11, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000ec, 5'd3, 27'h000003d5, 5'd20, 27'h0000035f, 32'h00000400,
  1'd1,  5'd6, 27'h0000035d, 5'd14, 27'h000003bd, 5'd8, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002b1, 5'd10, 27'h000003a8, 5'd17, 27'h00000252, 32'h00000400,
  1'd1,  5'd9, 27'h000002e0, 5'd15, 27'h000000d8, 5'd27, 27'h00000254, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e7, 5'd23, 27'h000003a0, 5'd7, 27'h00000186, 32'h00000400,
  1'd1,  5'd5, 27'h00000176, 5'd23, 27'h0000020a, 5'd20, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000d3, 5'd25, 27'h0000011d, 5'd26, 27'h000003d7, 32'h00000400,
  1'd1,  5'd18, 27'h000003a1, 5'd4, 27'h00000047, 5'd2, 27'h000003f2, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000011d, 5'd3, 27'h000000f8, 5'd11, 27'h00000333, 32'h00000400,
  1'd1,  5'd19, 27'h0000006c, 5'd1, 27'h000000d6, 5'd21, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000027e, 5'd13, 27'h000002fb, 5'd9, 27'h00000216, 32'h00000400,
  1'd1,  5'd20, 27'h00000004, 5'd13, 27'h00000087, 5'd19, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030a, 5'd13, 27'h000000e2, 5'd29, 27'h0000000a, 32'h00000400,
  1'd1,  5'd16, 27'h00000075, 5'd20, 27'h000003f5, 5'd8, 27'h0000003a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003d7, 5'd22, 27'h000002cc, 5'd17, 27'h0000014b, 32'h00000400,
  1'd1,  5'd17, 27'h000001df, 5'd24, 27'h00000386, 5'd30, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000100, 5'd3, 27'h000001db, 5'd7, 27'h0000028f, 32'h00000400,
  1'd1,  5'd26, 27'h00000227, 5'd4, 27'h000001e3, 5'd17, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000f7, 5'd3, 27'h00000068, 5'd29, 27'h000001cd, 32'h00000400,
  1'd1,  5'd30, 27'h000003d9, 5'd12, 27'h000000a4, 5'd5, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021e, 5'd12, 27'h0000027f, 5'd16, 27'h00000362, 32'h00000400,
  1'd1,  5'd30, 27'h00000215, 5'd14, 27'h0000014a, 5'd30, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000238, 5'd25, 27'h00000034, 5'd6, 27'h0000000a, 32'h00000400,
  1'd1,  5'd27, 27'h0000030d, 5'd21, 27'h00000196, 5'd17, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000177, 5'd25, 27'h000001f8, 5'd27, 27'h00000327, 32'h00000400,
  1'd1,  5'd9, 27'h0000018b, 5'd6, 27'h000001a1, 5'd2, 27'h00000392, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000004d, 5'd7, 27'h00000361, 5'd15, 27'h0000017d, 32'h00000400,
  1'd1,  5'd7, 27'h00000184, 5'd8, 27'h0000020c, 5'd22, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ab, 5'd20, 27'h000000a1, 5'd3, 27'h000001ff, 32'h00000400,
  1'd1,  5'd9, 27'h000001d3, 5'd18, 27'h000001d3, 5'd11, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b5, 5'd19, 27'h00000149, 5'd25, 27'h00000102, 32'h00000400,
  1'd1,  5'd6, 27'h000001d7, 5'd26, 27'h000002b2, 5'd2, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003fd, 5'd28, 27'h000002a5, 5'd11, 27'h0000032c, 32'h00000400,
  1'd1,  5'd8, 27'h0000030a, 5'd30, 27'h000000b6, 5'd21, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000306, 5'd6, 27'h00000104, 5'd1, 27'h000002f9, 32'h00000400,
  1'd1,  5'd18, 27'h000000d2, 5'd9, 27'h000003f9, 5'd14, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000276, 5'd5, 27'h000002f9, 5'd23, 27'h00000275, 32'h00000400,
  1'd1,  5'd16, 27'h000002cf, 5'd18, 27'h00000354, 5'd0, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000313, 5'd18, 27'h00000140, 5'd12, 27'h00000139, 32'h00000400,
  1'd1,  5'd15, 27'h00000318, 5'd19, 27'h00000221, 5'd24, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000014c, 5'd28, 27'h0000006d, 5'd1, 27'h000003a8, 32'h00000400,
  1'd1,  5'd16, 27'h0000037c, 5'd27, 27'h00000379, 5'd14, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002be, 5'd28, 27'h000000fd, 5'd21, 27'h000000b5, 32'h00000400,
  1'd1,  5'd28, 27'h00000165, 5'd7, 27'h00000019, 5'd0, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000034f, 5'd9, 27'h00000205, 5'd11, 27'h0000022c, 32'h00000400,
  1'd1,  5'd27, 27'h000001e2, 5'd7, 27'h00000213, 5'd23, 27'h0000032a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f9, 5'd20, 27'h000000e1, 5'd3, 27'h000000f4, 32'h00000400,
  1'd1,  5'd28, 27'h000001f8, 5'd19, 27'h000001b9, 5'd12, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000044, 5'd17, 27'h000000b6, 5'd24, 27'h000002c0, 32'h00000400,
  1'd1,  5'd26, 27'h0000026e, 5'd27, 27'h000001f3, 5'd1, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001dc, 5'd27, 27'h000001ad, 5'd13, 27'h000003a2, 32'h00000400,
  1'd1,  5'd29, 27'h0000038d, 5'd27, 27'h0000005b, 5'd23, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000012a, 5'd7, 27'h00000134, 5'd9, 27'h0000030a, 32'h00000400,
  1'd1,  5'd9, 27'h00000037, 5'd9, 27'h00000306, 5'd19, 27'h000001dd, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000007, 5'd6, 27'h000001ec, 5'd27, 27'h000002d9, 32'h00000400,
  1'd1,  5'd9, 27'h00000108, 5'd20, 27'h000000b8, 5'd9, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003ef, 5'd18, 27'h00000158, 5'd18, 27'h000002bf, 32'h00000400,
  1'd1,  5'd5, 27'h000001f0, 5'd20, 27'h000001a5, 5'd28, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000026d, 5'd29, 27'h0000002c, 5'd6, 27'h00000338, 32'h00000400,
  1'd1,  5'd6, 27'h000000f4, 5'd28, 27'h00000066, 5'd17, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000254, 5'd27, 27'h000002b7, 5'd29, 27'h000001a1, 32'h00000400,
  1'd1,  5'd18, 27'h0000006b, 5'd9, 27'h00000218, 5'd8, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003ed, 5'd8, 27'h0000034d, 5'd20, 27'h0000015f, 32'h00000400,
  1'd1,  5'd15, 27'h00000228, 5'd9, 27'h00000141, 5'd30, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000016b, 5'd16, 27'h000001a9, 5'd8, 27'h0000035b, 32'h00000400,
  1'd1,  5'd16, 27'h000001bb, 5'd15, 27'h00000219, 5'd19, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000036a, 5'd16, 27'h000002d6, 5'd27, 27'h0000016e, 32'h00000400,
  1'd1,  5'd19, 27'h0000032b, 5'd29, 27'h000002d6, 5'd9, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000310, 5'd29, 27'h00000051, 5'd15, 27'h00000275, 32'h00000400,
  1'd1,  5'd17, 27'h000000b1, 5'd29, 27'h0000004d, 5'd30, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000034e, 5'd8, 27'h0000002d, 5'd8, 27'h000001b2, 32'h00000400,
  1'd1,  5'd29, 27'h00000069, 5'd5, 27'h00000155, 5'd17, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000271, 5'd10, 27'h00000022, 5'd30, 27'h000002bc, 32'h00000400,
  1'd1,  5'd27, 27'h00000229, 5'd15, 27'h000003cd, 5'd8, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002d8, 5'd16, 27'h000002c8, 5'd18, 27'h00000077, 32'h00000400,
  1'd1,  5'd29, 27'h000001a9, 5'd18, 27'h00000249, 5'd29, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000010, 5'd28, 27'h00000213, 5'd7, 27'h00000011, 32'h00000400,
  1'd1,  5'd27, 27'h000000c7, 5'd30, 27'h000000f5, 5'd16, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000006f, 5'd28, 27'h0000004e, 5'd30, 27'h000001fc, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000001ab, 5'd4, 27'h00000006, 5'd3, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000dd, 5'd1, 27'h000002b2, 5'd12, 27'h000001fd, 32'h00000400,
  1'd1,  5'd2, 27'h0000025a, 5'd3, 27'h000000ee, 5'd21, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000011e, 5'd13, 27'h0000009f, 5'd1, 27'h000001b3, 32'h00000400,
  1'd1,  5'd4, 27'h00000223, 5'd11, 27'h00000284, 5'd10, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000359, 5'd12, 27'h00000089, 5'd22, 27'h00000258, 32'h00000400,
  1'd1,  5'd1, 27'h0000024a, 5'd23, 27'h000001ff, 5'd2, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000341, 5'd25, 27'h00000352, 5'd15, 27'h00000020, 32'h00000400,
  1'd1,  5'd3, 27'h00000322, 5'd22, 27'h0000014a, 5'd25, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000250, 5'd1, 27'h00000082, 5'd0, 27'h0000035f, 32'h00000400,
  1'd1,  5'd11, 27'h00000385, 5'd2, 27'h00000062, 5'd14, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000049, 5'd1, 27'h00000363, 5'd24, 27'h000001ec, 32'h00000400,
  1'd1,  5'd11, 27'h000003aa, 5'd10, 27'h00000249, 5'd0, 27'h000002ae, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000388, 5'd14, 27'h00000129, 5'd14, 27'h000001b8, 32'h00000400,
  1'd1,  5'd11, 27'h00000327, 5'd13, 27'h0000031e, 5'd25, 27'h0000016e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000356, 5'd22, 27'h00000115, 5'd2, 27'h000001bc, 32'h00000400,
  1'd1,  5'd11, 27'h000001aa, 5'd25, 27'h0000013a, 5'd12, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000002a, 5'd21, 27'h0000031c, 5'd24, 27'h000000bb, 32'h00000400,
  1'd1,  5'd22, 27'h00000112, 5'd4, 27'h0000030b, 5'd1, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000039a, 5'd1, 27'h00000301, 5'd13, 27'h00000052, 32'h00000400,
  1'd1,  5'd23, 27'h00000254, 5'd4, 27'h00000062, 5'd25, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001f, 5'd14, 27'h00000226, 5'd3, 27'h00000090, 32'h00000400,
  1'd1,  5'd21, 27'h000003a3, 5'd15, 27'h00000087, 5'd14, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000133, 5'd10, 27'h00000171, 5'd23, 27'h000002e0, 32'h00000400,
  1'd1,  5'd25, 27'h00000287, 5'd21, 27'h00000086, 5'd1, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a9, 5'd21, 27'h0000010f, 5'd11, 27'h0000030b, 32'h00000400,
  1'd1,  5'd21, 27'h0000010a, 5'd22, 27'h000001e8, 5'd20, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000190, 5'd4, 27'h00000372, 5'd9, 27'h00000227, 32'h00000400,
  1'd1,  5'd1, 27'h000003c4, 5'd4, 27'h00000310, 5'd18, 27'h000001b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000020a, 5'd2, 27'h0000027a, 5'd29, 27'h000001d3, 32'h00000400,
  1'd1,  5'd2, 27'h00000174, 5'd10, 27'h0000029a, 5'd9, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e8, 5'd14, 27'h000003c2, 5'd19, 27'h000001fe, 32'h00000400,
  1'd1,  5'd4, 27'h000002c7, 5'd13, 27'h00000283, 5'd30, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000005a, 5'd20, 27'h00000382, 5'd6, 27'h00000347, 32'h00000400,
  1'd1,  5'd1, 27'h00000197, 5'd21, 27'h000002ff, 5'd16, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002d3, 5'd24, 27'h0000014d, 5'd28, 27'h00000155, 32'h00000400,
  1'd1,  5'd15, 27'h00000031, 5'd3, 27'h000002b2, 5'd9, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000233, 5'd1, 27'h00000277, 5'd16, 27'h000002d2, 32'h00000400,
  1'd1,  5'd10, 27'h0000016a, 5'd2, 27'h00000379, 5'd29, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002ba, 5'd10, 27'h000003a4, 5'd7, 27'h00000282, 32'h00000400,
  1'd1,  5'd11, 27'h00000098, 5'd14, 27'h0000024a, 5'd17, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000167, 5'd14, 27'h00000173, 5'd27, 27'h00000360, 32'h00000400,
  1'd1,  5'd15, 27'h0000007f, 5'd23, 27'h00000097, 5'd8, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000366, 5'd24, 27'h000001b5, 5'd17, 27'h00000107, 32'h00000400,
  1'd1,  5'd13, 27'h00000090, 5'd25, 27'h00000163, 5'd29, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000023e, 5'd0, 27'h00000290, 5'd6, 27'h00000098, 32'h00000400,
  1'd1,  5'd23, 27'h0000034d, 5'd0, 27'h00000164, 5'd18, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001de, 5'd5, 27'h000000ab, 5'd28, 27'h00000368, 32'h00000400,
  1'd1,  5'd22, 27'h000000b8, 5'd12, 27'h0000035b, 5'd7, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000130, 5'd11, 27'h000002f2, 5'd16, 27'h00000216, 32'h00000400,
  1'd1,  5'd21, 27'h0000024e, 5'd13, 27'h000001f5, 5'd30, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000188, 5'd20, 27'h0000037d, 5'd6, 27'h000003b4, 32'h00000400,
  1'd1,  5'd23, 27'h0000027e, 5'd24, 27'h0000019c, 5'd15, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001df, 5'd22, 27'h00000247, 5'd29, 27'h000003a6, 32'h00000400,
  1'd1,  5'd2, 27'h000002e5, 5'd9, 27'h000002f5, 5'd4, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000010a, 5'd6, 27'h000001a6, 5'd10, 27'h00000198, 32'h00000400,
  1'd1,  5'd0, 27'h000002a5, 5'd5, 27'h00000273, 5'd23, 27'h00000146, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000260, 5'd15, 27'h0000023e, 5'd3, 27'h00000130, 32'h00000400,
  1'd1,  5'd2, 27'h000003bb, 5'd16, 27'h0000003b, 5'd11, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000316, 5'd16, 27'h000001e8, 5'd24, 27'h000000e3, 32'h00000400,
  1'd1,  5'd0, 27'h0000023a, 5'd28, 27'h00000211, 5'd0, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001f0, 5'd30, 27'h000000a8, 5'd11, 27'h0000003b, 32'h00000400,
  1'd1,  5'd2, 27'h0000001e, 5'd26, 27'h00000146, 5'd20, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000003e, 5'd6, 27'h00000361, 5'd3, 27'h000003f4, 32'h00000400,
  1'd1,  5'd11, 27'h000002ed, 5'd5, 27'h000003b5, 5'd10, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000bf, 5'd5, 27'h000002c4, 5'd25, 27'h00000247, 32'h00000400,
  1'd1,  5'd13, 27'h00000342, 5'd15, 27'h000003b8, 5'd1, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001a5, 5'd15, 27'h000003c4, 5'd13, 27'h00000060, 32'h00000400,
  1'd1,  5'd12, 27'h0000034c, 5'd18, 27'h0000030a, 5'd21, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000028, 5'd29, 27'h0000010d, 5'd1, 27'h00000265, 32'h00000400,
  1'd1,  5'd11, 27'h000003c0, 5'd30, 27'h0000027e, 5'd14, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000024b, 5'd28, 27'h000000c4, 5'd23, 27'h00000130, 32'h00000400,
  1'd1,  5'd21, 27'h000001cc, 5'd7, 27'h0000027d, 5'd4, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001ef, 5'd7, 27'h000001b9, 5'd13, 27'h000000b5, 32'h00000400,
  1'd1,  5'd23, 27'h00000314, 5'd16, 27'h000001d2, 5'd1, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b9, 5'd16, 27'h00000267, 5'd14, 27'h00000126, 32'h00000400,
  1'd1,  5'd20, 27'h000002ce, 5'd18, 27'h0000012d, 5'd20, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000232, 5'd29, 27'h0000027d, 5'd3, 27'h00000259, 32'h00000400,
  1'd1,  5'd22, 27'h0000016b, 5'd29, 27'h0000008e, 5'd13, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002f3, 5'd26, 27'h0000030b, 5'd24, 27'h000002fe, 32'h00000400,
  1'd1,  5'd0, 27'h000000d7, 5'd8, 27'h000002eb, 5'd9, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000a4, 5'd7, 27'h000000a9, 5'd18, 27'h0000012b, 32'h00000400,
  1'd1,  5'd3, 27'h00000230, 5'd6, 27'h00000271, 5'd27, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000303, 5'd19, 27'h0000038f, 5'd6, 27'h0000030b, 32'h00000400,
  1'd1,  5'd3, 27'h000003f9, 5'd15, 27'h000003e1, 5'd19, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000024c, 5'd17, 27'h00000091, 5'd26, 27'h000002c6, 32'h00000400,
  1'd1,  5'd0, 27'h000000c0, 5'd28, 27'h00000213, 5'd8, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000354, 5'd28, 27'h00000079, 5'd15, 27'h00000271, 32'h00000400,
  1'd1,  5'd1, 27'h0000001b, 5'd25, 27'h000003b4, 5'd25, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000289, 5'd10, 27'h0000014f, 5'd6, 27'h000001cf, 32'h00000400,
  1'd1,  5'd11, 27'h000002e7, 5'd8, 27'h000001ab, 5'd16, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000019e, 5'd7, 27'h0000002d, 5'd30, 27'h00000012, 32'h00000400,
  1'd1,  5'd12, 27'h000000cc, 5'd15, 27'h000003f4, 5'd9, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002d0, 5'd19, 27'h000000c0, 5'd17, 27'h000000d3, 32'h00000400,
  1'd1,  5'd14, 27'h000003aa, 5'd20, 27'h000001d4, 5'd25, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000399, 5'd27, 27'h000003ba, 5'd7, 27'h0000020e, 32'h00000400,
  1'd1,  5'd13, 27'h00000359, 5'd26, 27'h00000280, 5'd16, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000000e, 5'd30, 27'h000002fc, 5'd26, 27'h0000014f, 32'h00000400,
  1'd1,  5'd22, 27'h000001fe, 5'd5, 27'h000000f9, 5'd6, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003ef, 5'd8, 27'h00000267, 5'd20, 27'h0000016a, 32'h00000400,
  1'd1,  5'd22, 27'h0000000b, 5'd9, 27'h000000cc, 5'd29, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002b7, 5'd17, 27'h0000019f, 5'd9, 27'h0000017b, 32'h00000400,
  1'd1,  5'd21, 27'h00000103, 5'd20, 27'h0000018d, 5'd17, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000049, 5'd18, 27'h00000358, 5'd29, 27'h000001b0, 32'h00000400,
  1'd1,  5'd23, 27'h0000029c, 5'd28, 27'h00000306, 5'd7, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e3, 5'd29, 27'h0000034b, 5'd18, 27'h00000136, 32'h00000400,
  1'd1,  5'd23, 27'h00000293, 5'd29, 27'h00000081, 5'd26, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000035f, 5'd4, 27'h00000151, 5'd7, 27'h0000016e, 32'h00000400,
  1'd1,  5'd5, 27'h000003e6, 5'd3, 27'h0000036a, 5'd16, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001de, 5'd3, 27'h0000037e, 5'd29, 27'h00000360, 32'h00000400,
  1'd1,  5'd7, 27'h0000030a, 5'd14, 27'h0000031f, 5'd0, 27'h00000125, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000010e, 5'd11, 27'h00000064, 5'd13, 27'h00000321, 32'h00000400,
  1'd1,  5'd6, 27'h0000031c, 5'd11, 27'h000003a3, 5'd23, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002da, 5'd24, 27'h0000036d, 5'd0, 27'h000003ef, 32'h00000400,
  1'd1,  5'd10, 27'h0000012f, 5'd21, 27'h000003de, 5'd12, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a7, 5'd22, 27'h0000035c, 5'd22, 27'h00000267, 32'h00000400,
  1'd1,  5'd19, 27'h000000d2, 5'd3, 27'h0000005b, 5'd6, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000021b, 5'd4, 27'h00000233, 5'd19, 27'h00000284, 32'h00000400,
  1'd1,  5'd17, 27'h00000025, 5'd2, 27'h000003b3, 5'd26, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002c9, 5'd14, 27'h0000025f, 5'd2, 27'h00000327, 32'h00000400,
  1'd1,  5'd19, 27'h0000002f, 5'd13, 27'h000000bb, 5'd12, 27'h00000118, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000286, 5'd11, 27'h000002e7, 5'd25, 27'h00000160, 32'h00000400,
  1'd1,  5'd16, 27'h000001e0, 5'd24, 27'h00000021, 5'd4, 27'h00000240, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001b8, 5'd25, 27'h0000012a, 5'd12, 27'h000000d7, 32'h00000400,
  1'd1,  5'd19, 27'h0000026a, 5'd24, 27'h00000292, 5'd24, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001d8, 5'd4, 27'h00000181, 5'd4, 27'h00000101, 32'h00000400,
  1'd1,  5'd28, 27'h000003f3, 5'd2, 27'h00000300, 5'd13, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000dd, 5'd4, 27'h0000005b, 5'd20, 27'h00000335, 32'h00000400,
  1'd1,  5'd26, 27'h0000013d, 5'd15, 27'h0000014c, 5'd4, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000fa, 5'd12, 27'h0000017f, 5'd14, 27'h0000027d, 32'h00000400,
  1'd1,  5'd28, 27'h00000114, 5'd13, 27'h00000359, 5'd24, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000188, 5'd25, 27'h00000160, 5'd3, 27'h000000cc, 32'h00000400,
  1'd1,  5'd30, 27'h00000130, 5'd21, 27'h00000311, 5'd13, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001d1, 5'd21, 27'h0000022b, 5'd21, 27'h00000246, 32'h00000400,
  1'd1,  5'd8, 27'h00000015, 5'd1, 27'h000002ed, 5'd2, 27'h00000184, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000054, 5'd1, 27'h000003ad, 5'd12, 27'h00000181, 32'h00000400,
  1'd1,  5'd7, 27'h00000027, 5'd1, 27'h0000036d, 5'd22, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000105, 5'd14, 27'h0000017a, 5'd7, 27'h000003ee, 32'h00000400,
  1'd1,  5'd5, 27'h000003fe, 5'd12, 27'h000000e2, 5'd20, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000332, 5'd14, 27'h00000148, 5'd27, 27'h0000015d, 32'h00000400,
  1'd1,  5'd9, 27'h000002de, 5'd22, 27'h00000283, 5'd6, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001f0, 5'd24, 27'h000002d1, 5'd16, 27'h00000140, 32'h00000400,
  1'd1,  5'd8, 27'h0000003e, 5'd21, 27'h00000136, 5'd29, 27'h000002d9, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003de, 5'd4, 27'h00000045, 5'd3, 27'h000000d7, 32'h00000400,
  1'd1,  5'd15, 27'h000002a5, 5'd2, 27'h0000011e, 5'd10, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001c3, 5'd2, 27'h00000112, 5'd22, 27'h0000016c, 32'h00000400,
  1'd1,  5'd20, 27'h000001c2, 5'd10, 27'h00000283, 5'd9, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000fb, 5'd10, 27'h0000019c, 5'd15, 27'h0000024d, 32'h00000400,
  1'd1,  5'd19, 27'h0000027f, 5'd11, 27'h000002f5, 5'd26, 27'h000001c7, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001b3, 5'd21, 27'h000003ee, 5'd7, 27'h00000247, 32'h00000400,
  1'd1,  5'd18, 27'h00000131, 5'd24, 27'h00000091, 5'd17, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000283, 5'd24, 27'h000001b5, 5'd26, 27'h00000071, 32'h00000400,
  1'd1,  5'd29, 27'h000002c1, 5'd4, 27'h0000029c, 5'd6, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003af, 5'd3, 27'h00000147, 5'd20, 27'h0000021d, 32'h00000400,
  1'd1,  5'd28, 27'h000003cc, 5'd2, 27'h0000015d, 5'd29, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000211, 5'd13, 27'h00000261, 5'd7, 27'h00000094, 32'h00000400,
  1'd1,  5'd26, 27'h00000051, 5'd12, 27'h0000014f, 5'd19, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003cd, 5'd12, 27'h000002c8, 5'd28, 27'h00000333, 32'h00000400,
  1'd1,  5'd28, 27'h000003d3, 5'd21, 27'h00000075, 5'd9, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000118, 5'd22, 27'h000000f0, 5'd17, 27'h000002f1, 32'h00000400,
  1'd1,  5'd28, 27'h0000011e, 5'd25, 27'h00000110, 5'd30, 27'h0000024a, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003b5, 5'd9, 27'h0000021f, 5'd1, 27'h00000219, 32'h00000400,
  1'd1,  5'd9, 27'h00000193, 5'd5, 27'h0000033f, 5'd13, 27'h0000013a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000232, 5'd7, 27'h000000f6, 5'd21, 27'h0000019a, 32'h00000400,
  1'd1,  5'd8, 27'h0000010a, 5'd19, 27'h0000028c, 5'd2, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000315, 5'd20, 27'h000001c1, 5'd13, 27'h00000159, 32'h00000400,
  1'd1,  5'd10, 27'h0000004c, 5'd18, 27'h000001e1, 5'd24, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000038f, 5'd27, 27'h000003fc, 5'd1, 27'h000002ac, 32'h00000400,
  1'd1,  5'd8, 27'h0000003c, 5'd30, 27'h00000202, 5'd14, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000286, 5'd28, 27'h0000011f, 5'd23, 27'h0000038f, 32'h00000400,
  1'd1,  5'd16, 27'h000003b5, 5'd8, 27'h00000142, 5'd1, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000188, 5'd7, 27'h000000bd, 5'd10, 27'h000003db, 32'h00000400,
  1'd1,  5'd20, 27'h00000179, 5'd9, 27'h0000038f, 5'd25, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000343, 5'd17, 27'h000002ab, 5'd4, 27'h000000b6, 32'h00000400,
  1'd1,  5'd19, 27'h000002b8, 5'd16, 27'h000001f1, 5'd13, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000267, 5'd17, 27'h000003fa, 5'd24, 27'h00000098, 32'h00000400,
  1'd1,  5'd19, 27'h0000003c, 5'd28, 27'h000003eb, 5'd0, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000069, 5'd29, 27'h0000039c, 5'd12, 27'h00000090, 32'h00000400,
  1'd1,  5'd20, 27'h00000293, 5'd27, 27'h00000207, 5'd22, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001c5, 5'd9, 27'h0000020f, 5'd1, 27'h000003cc, 32'h00000400,
  1'd1,  5'd28, 27'h00000018, 5'd6, 27'h00000331, 5'd10, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000c3, 5'd9, 27'h00000260, 5'd21, 27'h0000031c, 32'h00000400,
  1'd1,  5'd26, 27'h000003ed, 5'd17, 27'h000003d6, 5'd3, 27'h000001d5, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000e7, 5'd20, 27'h00000074, 5'd11, 27'h00000057, 32'h00000400,
  1'd1,  5'd28, 27'h00000398, 5'd19, 27'h0000001b, 5'd25, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000327, 5'd27, 27'h0000023b, 5'd0, 27'h000000ea, 32'h00000400,
  1'd1,  5'd29, 27'h0000018d, 5'd26, 27'h00000277, 5'd13, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003cc, 5'd27, 27'h0000006e, 5'd25, 27'h00000210, 32'h00000400,
  1'd1,  5'd8, 27'h000002f8, 5'd9, 27'h0000035d, 5'd7, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000294, 5'd10, 27'h00000089, 5'd19, 27'h0000019f, 32'h00000400,
  1'd1,  5'd6, 27'h000003b0, 5'd8, 27'h00000202, 5'd28, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000bc, 5'd18, 27'h00000271, 5'd6, 27'h000000f7, 32'h00000400,
  1'd1,  5'd8, 27'h000002b4, 5'd17, 27'h0000018e, 5'd19, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000071, 5'd18, 27'h0000034a, 5'd26, 27'h0000024f, 32'h00000400,
  1'd1,  5'd9, 27'h00000221, 5'd26, 27'h000003e0, 5'd6, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a8, 5'd27, 27'h00000017, 5'd18, 27'h00000017, 32'h00000400,
  1'd1,  5'd7, 27'h0000001e, 5'd29, 27'h000002f8, 5'd29, 27'h000001de, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000196, 5'd6, 27'h00000237, 5'd10, 27'h0000010b, 32'h00000400,
  1'd1,  5'd19, 27'h000000bb, 5'd6, 27'h00000169, 5'd18, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003b1, 5'd9, 27'h00000345, 5'd29, 27'h00000179, 32'h00000400,
  1'd1,  5'd16, 27'h0000008d, 5'd18, 27'h000001a1, 5'd7, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000227, 5'd19, 27'h000003de, 5'd16, 27'h00000345, 32'h00000400,
  1'd1,  5'd18, 27'h00000052, 5'd17, 27'h00000350, 5'd30, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000116, 5'd28, 27'h000002af, 5'd8, 27'h0000013e, 32'h00000400,
  1'd1,  5'd18, 27'h000002ad, 5'd28, 27'h000003bd, 5'd16, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000003a, 5'd30, 27'h000001a2, 5'd27, 27'h000002a5, 32'h00000400,
  1'd1,  5'd25, 27'h000003f3, 5'd8, 27'h0000034b, 5'd7, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000398, 5'd5, 27'h0000029c, 5'd18, 27'h00000329, 32'h00000400,
  1'd1,  5'd28, 27'h000002b3, 5'd5, 27'h000000b5, 5'd29, 27'h000000f6, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000082, 5'd19, 27'h000000c7, 5'd7, 27'h000003c3, 32'h00000400,
  1'd1,  5'd27, 27'h00000009, 5'd20, 27'h000000a0, 5'd16, 27'h00000025, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000001, 5'd18, 27'h0000039b, 5'd27, 27'h000000f9, 32'h00000400,
  1'd1,  5'd27, 27'h0000024d, 5'd28, 27'h000000ad, 5'd7, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000212, 5'd29, 27'h000002e7, 5'd17, 27'h00000067, 32'h00000400,
  1'd1,  5'd26, 27'h000002a6, 5'd29, 27'h000002b2, 5'd27, 27'h00000176, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h0000004c, 5'd4, 27'h0000036b, 5'd5, 27'h00000032, 32'h00000400,
  1'd1,  5'd3, 27'h00000162, 5'd2, 27'h00000173, 5'd13, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000231, 5'd2, 27'h0000016e, 5'd25, 27'h00000208, 32'h00000400,
  1'd1,  5'd4, 27'h00000018, 5'd13, 27'h000002b2, 5'd1, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000287, 5'd13, 27'h0000023b, 5'd12, 27'h000000ff, 32'h00000400,
  1'd1,  5'd1, 27'h0000031b, 5'd13, 27'h00000343, 5'd24, 27'h000000c7, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000318, 5'd22, 27'h00000096, 5'd1, 27'h000002a8, 32'h00000400,
  1'd1,  5'd1, 27'h00000062, 5'd23, 27'h0000038b, 5'd12, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000002, 5'd21, 27'h0000011c, 5'd24, 27'h00000303, 32'h00000400,
  1'd1,  5'd13, 27'h00000345, 5'd3, 27'h00000161, 5'd3, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000053, 5'd5, 27'h00000023, 5'd15, 27'h00000007, 32'h00000400,
  1'd1,  5'd12, 27'h00000316, 5'd3, 27'h000002e1, 5'd24, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000013c, 5'd15, 27'h000000fd, 5'd3, 27'h000001dd, 32'h00000400,
  1'd1,  5'd14, 27'h00000061, 5'd10, 27'h000001f8, 5'd13, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001bd, 5'd11, 27'h00000216, 5'd21, 27'h000000b4, 32'h00000400,
  1'd1,  5'd12, 27'h000000d0, 5'd21, 27'h000001ec, 5'd4, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000be, 5'd25, 27'h00000030, 5'd14, 27'h00000166, 32'h00000400,
  1'd1,  5'd12, 27'h00000090, 5'd23, 27'h000000c0, 5'd21, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000017a, 5'd0, 27'h000000d9, 5'd0, 27'h0000031e, 32'h00000400,
  1'd1,  5'd22, 27'h00000159, 5'd2, 27'h00000350, 5'd12, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000002, 5'd4, 27'h0000036a, 5'd20, 27'h000002e3, 32'h00000400,
  1'd1,  5'd22, 27'h000002ea, 5'd11, 27'h00000080, 5'd2, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000023c, 5'd14, 27'h00000072, 5'd13, 27'h000000b1, 32'h00000400,
  1'd1,  5'd25, 27'h000002ff, 5'd13, 27'h00000390, 5'd25, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000f7, 5'd22, 27'h00000201, 5'd2, 27'h00000377, 32'h00000400,
  1'd1,  5'd25, 27'h00000147, 5'd24, 27'h0000006a, 5'd14, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003f9, 5'd24, 27'h00000225, 5'd24, 27'h0000001a, 32'h00000400,
  1'd1,  5'd1, 27'h00000303, 5'd2, 27'h00000398, 5'd5, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002c3, 5'd0, 27'h00000312, 5'd16, 27'h000000ad, 32'h00000400,
  1'd1,  5'd4, 27'h000000f9, 5'd4, 27'h00000064, 5'd29, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ec, 5'd12, 27'h000003ef, 5'd9, 27'h00000114, 32'h00000400,
  1'd1,  5'd3, 27'h000001a4, 5'd14, 27'h00000313, 5'd19, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012e, 5'd11, 27'h000003a2, 5'd25, 27'h000003a0, 32'h00000400,
  1'd1,  5'd0, 27'h00000266, 5'd25, 27'h00000093, 5'd5, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002c7, 5'd21, 27'h000001ad, 5'd16, 27'h00000150, 32'h00000400,
  1'd1,  5'd0, 27'h0000035f, 5'd23, 27'h00000135, 5'd29, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000011a, 5'd3, 27'h000001b0, 5'd10, 27'h00000059, 32'h00000400,
  1'd1,  5'd11, 27'h00000268, 5'd2, 27'h000000c1, 5'd18, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000039f, 5'd1, 27'h000002e3, 5'd28, 27'h000002aa, 32'h00000400,
  1'd1,  5'd10, 27'h000001c6, 5'd12, 27'h000000d6, 5'd9, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000029a, 5'd11, 27'h00000145, 5'd18, 27'h00000374, 32'h00000400,
  1'd1,  5'd12, 27'h0000027a, 5'd15, 27'h00000097, 5'd27, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c2, 5'd25, 27'h00000218, 5'd6, 27'h00000101, 32'h00000400,
  1'd1,  5'd13, 27'h00000037, 5'd23, 27'h00000379, 5'd19, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000035a, 5'd25, 27'h0000010d, 5'd29, 27'h0000022f, 32'h00000400,
  1'd1,  5'd25, 27'h000002b4, 5'd3, 27'h0000008f, 5'd7, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003e5, 5'd1, 27'h000002ad, 5'd17, 27'h0000003e, 32'h00000400,
  1'd1,  5'd21, 27'h0000006b, 5'd1, 27'h000000a1, 5'd26, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000cf, 5'd13, 27'h00000061, 5'd9, 27'h00000321, 32'h00000400,
  1'd1,  5'd24, 27'h000002a9, 5'd11, 27'h000001f2, 5'd18, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000303, 5'd12, 27'h00000088, 5'd25, 27'h0000035d, 32'h00000400,
  1'd1,  5'd22, 27'h00000337, 5'd20, 27'h00000322, 5'd5, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000001f, 5'd22, 27'h00000357, 5'd20, 27'h00000085, 32'h00000400,
  1'd1,  5'd23, 27'h00000246, 5'd23, 27'h0000027f, 5'd26, 27'h00000242, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000357, 5'd5, 27'h000003fe, 5'd0, 27'h000000e3, 32'h00000400,
  1'd1,  5'd0, 27'h0000000d, 5'd7, 27'h000001b7, 5'd10, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000139, 5'd8, 27'h0000004b, 5'd21, 27'h0000017b, 32'h00000400,
  1'd1,  5'd1, 27'h000001b1, 5'd16, 27'h000000fa, 5'd4, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000035f, 5'd18, 27'h00000105, 5'd13, 27'h000000f6, 32'h00000400,
  1'd1,  5'd4, 27'h0000019e, 5'd18, 27'h0000011c, 5'd25, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000006d, 5'd26, 27'h00000069, 5'd1, 27'h00000195, 32'h00000400,
  1'd1,  5'd3, 27'h00000117, 5'd29, 27'h0000000a, 5'd12, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002e3, 5'd29, 27'h00000123, 5'd22, 27'h00000111, 32'h00000400,
  1'd1,  5'd10, 27'h000001f2, 5'd5, 27'h00000221, 5'd1, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000273, 5'd9, 27'h00000050, 5'd14, 27'h00000255, 32'h00000400,
  1'd1,  5'd12, 27'h00000267, 5'd5, 27'h0000036b, 5'd24, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000013f, 5'd17, 27'h00000360, 5'd3, 27'h000001dc, 32'h00000400,
  1'd1,  5'd10, 27'h00000190, 5'd16, 27'h000000d3, 5'd10, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020f, 5'd19, 27'h0000023f, 5'd22, 27'h000002d2, 32'h00000400,
  1'd1,  5'd14, 27'h0000009f, 5'd28, 27'h00000172, 5'd3, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000058, 5'd27, 27'h000000d9, 5'd14, 27'h0000031d, 32'h00000400,
  1'd1,  5'd14, 27'h00000270, 5'd26, 27'h000002f9, 5'd22, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000287, 5'd6, 27'h0000029e, 5'd3, 27'h000003bb, 32'h00000400,
  1'd1,  5'd21, 27'h0000033d, 5'd9, 27'h00000023, 5'd10, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000014c, 5'd15, 27'h00000226, 5'd3, 27'h0000024e, 32'h00000400,
  1'd1,  5'd23, 27'h00000164, 5'd19, 27'h000001f4, 5'd15, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001e8, 5'd19, 27'h0000031a, 5'd24, 27'h0000002b, 32'h00000400,
  1'd1,  5'd21, 27'h00000031, 5'd26, 27'h000003f5, 5'd3, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035b, 5'd27, 27'h0000013f, 5'd11, 27'h00000105, 32'h00000400,
  1'd1,  5'd22, 27'h0000022f, 5'd25, 27'h000003cd, 5'd21, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000266, 5'd8, 27'h000003fc, 5'd7, 27'h000002af, 32'h00000400,
  1'd1,  5'd3, 27'h00000274, 5'd5, 27'h0000025d, 5'd20, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000056, 5'd7, 27'h00000279, 5'd27, 27'h00000196, 32'h00000400,
  1'd1,  5'd0, 27'h00000369, 5'd17, 27'h00000263, 5'd8, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000016d, 5'd15, 27'h000002d7, 5'd20, 27'h00000052, 32'h00000400,
  1'd1,  5'd3, 27'h000000ac, 5'd20, 27'h00000193, 5'd26, 27'h000002d0, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000001d, 5'd29, 27'h000003db, 5'd9, 27'h000001f4, 32'h00000400,
  1'd1,  5'd4, 27'h0000039f, 5'd30, 27'h000001de, 5'd19, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001d4, 5'd27, 27'h000003e8, 5'd30, 27'h000003c6, 32'h00000400,
  1'd1,  5'd13, 27'h00000245, 5'd6, 27'h000002b5, 5'd6, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002c9, 5'd9, 27'h0000010e, 5'd18, 27'h0000008a, 32'h00000400,
  1'd1,  5'd11, 27'h00000005, 5'd6, 27'h00000037, 5'd26, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000073, 5'd17, 27'h000000e0, 5'd6, 27'h000003a7, 32'h00000400,
  1'd1,  5'd14, 27'h000000ed, 5'd16, 27'h0000015b, 5'd19, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c4, 5'd20, 27'h000001dc, 5'd28, 27'h00000162, 32'h00000400,
  1'd1,  5'd14, 27'h000002d0, 5'd26, 27'h00000215, 5'd9, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e6, 5'd28, 27'h00000329, 5'd15, 27'h0000032a, 32'h00000400,
  1'd1,  5'd14, 27'h000000bf, 5'd28, 27'h00000379, 5'd27, 27'h0000035b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000031c, 5'd6, 27'h000002c6, 5'd8, 27'h00000145, 32'h00000400,
  1'd1,  5'd20, 27'h00000359, 5'd9, 27'h000002bb, 5'd18, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001e8, 5'd8, 27'h00000268, 5'd27, 27'h0000009e, 32'h00000400,
  1'd1,  5'd25, 27'h0000031f, 5'd16, 27'h000000e4, 5'd9, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000180, 5'd16, 27'h000002fb, 5'd16, 27'h00000355, 32'h00000400,
  1'd1,  5'd23, 27'h000001c7, 5'd16, 27'h00000120, 5'd29, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd22, 27'h000001b9, 5'd30, 27'h0000031a, 5'd9, 27'h00000366, 32'h00000400,
  1'd1,  5'd23, 27'h000000e4, 5'd28, 27'h000002e0, 5'd16, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000149, 5'd30, 27'h00000053, 5'd27, 27'h0000010e, 32'h00000400,
  1'd1,  5'd7, 27'h000001e2, 5'd2, 27'h00000371, 5'd7, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000022a, 5'd4, 27'h00000187, 5'd16, 27'h00000122, 32'h00000400,
  1'd1,  5'd10, 27'h000000b4, 5'd1, 27'h0000005e, 5'd30, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003c9, 5'd13, 27'h00000241, 5'd2, 27'h0000005a, 32'h00000400,
  1'd1,  5'd7, 27'h000003c8, 5'd11, 27'h0000037a, 5'd11, 27'h0000021a, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002cc, 5'd13, 27'h000000a1, 5'd22, 27'h0000011a, 32'h00000400,
  1'd1,  5'd9, 27'h00000100, 5'd22, 27'h0000008d, 5'd2, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000221, 5'd23, 27'h000001e9, 5'd13, 27'h000000bc, 32'h00000400,
  1'd1,  5'd10, 27'h000000ed, 5'd21, 27'h00000072, 5'd25, 27'h000001a0, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000342, 5'd1, 27'h00000151, 5'd6, 27'h000000ee, 32'h00000400,
  1'd1,  5'd17, 27'h0000008d, 5'd0, 27'h000001e3, 5'd17, 27'h0000022d, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000029, 5'd1, 27'h00000126, 5'd26, 27'h00000351, 32'h00000400,
  1'd1,  5'd20, 27'h0000012b, 5'd14, 27'h0000007b, 5'd3, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000369, 5'd12, 27'h000001d3, 5'd13, 27'h000001d0, 32'h00000400,
  1'd1,  5'd17, 27'h000002e9, 5'd12, 27'h000000b7, 5'd21, 27'h0000030b, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000306, 5'd23, 27'h000003a5, 5'd1, 27'h00000055, 32'h00000400,
  1'd1,  5'd16, 27'h0000000e, 5'd21, 27'h00000281, 5'd15, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ab, 5'd23, 27'h0000009b, 5'd23, 27'h00000172, 32'h00000400,
  1'd1,  5'd26, 27'h0000026e, 5'd3, 27'h0000016b, 5'd1, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000158, 5'd1, 27'h000002be, 5'd11, 27'h00000030, 32'h00000400,
  1'd1,  5'd27, 27'h000003f0, 5'd0, 27'h00000250, 5'd24, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000036c, 5'd12, 27'h00000086, 5'd1, 27'h00000126, 32'h00000400,
  1'd1,  5'd28, 27'h0000038f, 5'd14, 27'h00000349, 5'd13, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000008c, 5'd10, 27'h0000031e, 5'd24, 27'h000001ad, 32'h00000400,
  1'd1,  5'd26, 27'h0000021d, 5'd21, 27'h000003e0, 5'd3, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e8, 5'd22, 27'h0000021e, 5'd10, 27'h00000397, 32'h00000400,
  1'd1,  5'd26, 27'h0000025c, 5'd25, 27'h000001d5, 5'd21, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000032e, 5'd3, 27'h000002e7, 5'd1, 27'h0000004d, 32'h00000400,
  1'd1,  5'd6, 27'h000002d0, 5'd4, 27'h0000014e, 5'd10, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000be, 5'd0, 27'h00000215, 5'd25, 27'h000002f2, 32'h00000400,
  1'd1,  5'd5, 27'h00000386, 5'd10, 27'h0000037b, 5'd5, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000005f, 5'd13, 27'h00000313, 5'd15, 27'h00000203, 32'h00000400,
  1'd1,  5'd6, 27'h000002dc, 5'd12, 27'h000002f9, 5'd29, 27'h0000024c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002d3, 5'd24, 27'h000003f0, 5'd6, 27'h0000035c, 32'h00000400,
  1'd1,  5'd5, 27'h0000036f, 5'd25, 27'h00000193, 5'd19, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000140, 5'd20, 27'h000002ff, 5'd27, 27'h000003db, 32'h00000400,
  1'd1,  5'd17, 27'h00000012, 5'd2, 27'h000002c8, 5'd3, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d6, 5'd2, 27'h00000322, 5'd14, 27'h000001b1, 32'h00000400,
  1'd1,  5'd19, 27'h000002db, 5'd4, 27'h000001e0, 5'd22, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000026a, 5'd11, 27'h00000181, 5'd7, 27'h00000000, 32'h00000400,
  1'd1,  5'd16, 27'h000003b1, 5'd13, 27'h00000018, 5'd19, 27'h000003a8, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001a0, 5'd15, 27'h000001cd, 5'd28, 27'h0000003a, 32'h00000400,
  1'd1,  5'd16, 27'h00000076, 5'd23, 27'h0000015f, 5'd6, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000378, 5'd23, 27'h00000063, 5'd18, 27'h00000101, 32'h00000400,
  1'd1,  5'd19, 27'h00000261, 5'd25, 27'h0000015a, 5'd30, 27'h0000027f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003cc, 5'd0, 27'h000003f7, 5'd8, 27'h000001a2, 32'h00000400,
  1'd1,  5'd27, 27'h000001dd, 5'd2, 27'h000003ac, 5'd16, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000342, 5'd1, 27'h00000312, 5'd28, 27'h000002c4, 32'h00000400,
  1'd1,  5'd27, 27'h0000020e, 5'd11, 27'h00000072, 5'd8, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000020d, 5'd11, 27'h0000013f, 5'd19, 27'h0000024b, 32'h00000400,
  1'd1,  5'd30, 27'h00000183, 5'd14, 27'h0000010e, 5'd27, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000364, 5'd23, 27'h00000233, 5'd7, 27'h0000031b, 32'h00000400,
  1'd1,  5'd30, 27'h000001af, 5'd23, 27'h0000011c, 5'd18, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000035f, 5'd23, 27'h000001e9, 5'd25, 27'h0000036d, 32'h00000400,
  1'd1,  5'd8, 27'h00000198, 5'd5, 27'h00000323, 5'd0, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002b2, 5'd8, 27'h000003ac, 5'd15, 27'h00000188, 32'h00000400,
  1'd1,  5'd7, 27'h000002d0, 5'd6, 27'h00000237, 5'd23, 27'h00000092, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000002e, 5'd18, 27'h0000004c, 5'd4, 27'h0000015d, 32'h00000400,
  1'd1,  5'd9, 27'h000003f8, 5'd18, 27'h000001e9, 5'd13, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000332, 5'd18, 27'h000002de, 5'd24, 27'h00000020, 32'h00000400,
  1'd1,  5'd7, 27'h00000261, 5'd26, 27'h0000030c, 5'd0, 27'h000002d2, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000309, 5'd26, 27'h0000033c, 5'd11, 27'h00000262, 32'h00000400,
  1'd1,  5'd10, 27'h00000109, 5'd27, 27'h0000006e, 5'd20, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000018f, 5'd8, 27'h0000000f, 5'd4, 27'h0000027c, 32'h00000400,
  1'd1,  5'd16, 27'h0000009c, 5'd5, 27'h0000014d, 5'd14, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ba, 5'd10, 27'h00000073, 5'd23, 27'h0000019c, 32'h00000400,
  1'd1,  5'd15, 27'h00000306, 5'd15, 27'h000002df, 5'd5, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000129, 5'd17, 27'h00000239, 5'd10, 27'h00000273, 32'h00000400,
  1'd1,  5'd19, 27'h0000014e, 5'd20, 27'h00000042, 5'd21, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003e8, 5'd28, 27'h0000004e, 5'd2, 27'h0000034f, 32'h00000400,
  1'd1,  5'd15, 27'h000002fa, 5'd28, 27'h00000362, 5'd13, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000030f, 5'd28, 27'h000002ed, 5'd25, 27'h000001fc, 32'h00000400,
  1'd1,  5'd30, 27'h0000034c, 5'd7, 27'h0000014d, 5'd2, 27'h000001f4, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000309, 5'd8, 27'h000003ce, 5'd13, 27'h0000037a, 32'h00000400,
  1'd1,  5'd29, 27'h00000172, 5'd8, 27'h00000022, 5'd23, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000025e, 5'd20, 27'h0000022f, 5'd3, 27'h00000143, 32'h00000400,
  1'd1,  5'd26, 27'h000000f4, 5'd18, 27'h00000333, 5'd11, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000001e, 5'd19, 27'h000003c5, 5'd23, 27'h00000240, 32'h00000400,
  1'd1,  5'd27, 27'h0000021c, 5'd29, 27'h000003cf, 5'd1, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001e3, 5'd28, 27'h00000232, 5'd14, 27'h0000011e, 32'h00000400,
  1'd1,  5'd29, 27'h00000138, 5'd26, 27'h000001b2, 5'd20, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009e, 5'd8, 27'h000001a1, 5'd9, 27'h000003a7, 32'h00000400,
  1'd1,  5'd6, 27'h0000007e, 5'd5, 27'h000002d9, 5'd18, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b4, 5'd6, 27'h0000028a, 5'd27, 27'h0000028a, 32'h00000400,
  1'd1,  5'd10, 27'h00000050, 5'd18, 27'h000002c0, 5'd5, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003c9, 5'd20, 27'h0000002d, 5'd19, 27'h00000215, 32'h00000400,
  1'd1,  5'd6, 27'h00000086, 5'd18, 27'h00000239, 5'd26, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002e3, 5'd25, 27'h000003c2, 5'd9, 27'h00000252, 32'h00000400,
  1'd1,  5'd9, 27'h000003ac, 5'd29, 27'h00000030, 5'd19, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000343, 5'd30, 27'h000000af, 5'd28, 27'h000003b8, 32'h00000400,
  1'd1,  5'd15, 27'h00000292, 5'd8, 27'h000003a7, 5'd6, 27'h0000024b, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000183, 5'd8, 27'h00000258, 5'd18, 27'h000001a2, 32'h00000400,
  1'd1,  5'd16, 27'h000001e5, 5'd8, 27'h000002ad, 5'd30, 27'h000000ac, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000062, 5'd16, 27'h000002cc, 5'd8, 27'h00000137, 32'h00000400,
  1'd1,  5'd20, 27'h0000021a, 5'd15, 27'h00000365, 5'd20, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002b9, 5'd17, 27'h00000153, 5'd26, 27'h000001a0, 32'h00000400,
  1'd1,  5'd16, 27'h00000012, 5'd30, 27'h00000355, 5'd5, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000245, 5'd29, 27'h0000016e, 5'd18, 27'h00000293, 32'h00000400,
  1'd1,  5'd19, 27'h00000154, 5'd30, 27'h000000bd, 5'd26, 27'h0000019a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000160, 5'd7, 27'h0000003f, 5'd5, 27'h000002ea, 32'h00000400,
  1'd1,  5'd29, 27'h000002d1, 5'd6, 27'h000000c3, 5'd17, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000037f, 5'd8, 27'h00000133, 5'd30, 27'h00000147, 32'h00000400,
  1'd1,  5'd26, 27'h000002fb, 5'd17, 27'h00000076, 5'd6, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000271, 5'd17, 27'h000000f2, 5'd15, 27'h000003a9, 32'h00000400,
  1'd1,  5'd26, 27'h000002f2, 5'd18, 27'h000002ba, 5'd27, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002ef, 5'd30, 27'h0000038e, 5'd5, 27'h0000022d, 32'h00000400,
  1'd1,  5'd27, 27'h00000345, 5'd27, 27'h0000006e, 5'd20, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000002b, 5'd27, 27'h000000c8, 5'd29, 27'h00000277, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h000001de, 5'd1, 27'h00000278, 5'd4, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000241, 5'd4, 27'h000000f1, 5'd11, 27'h00000258, 32'h00000400,
  1'd1,  5'd2, 27'h000001c0, 5'd4, 27'h000001ca, 5'd24, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000331, 5'd10, 27'h000003d2, 5'd5, 27'h00000001, 32'h00000400,
  1'd1,  5'd0, 27'h0000033f, 5'd11, 27'h000003fe, 5'd10, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000031, 5'd15, 27'h00000096, 5'd24, 27'h0000027e, 32'h00000400,
  1'd1,  5'd1, 27'h00000040, 5'd25, 27'h000001a6, 5'd0, 27'h0000015a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000ac, 5'd23, 27'h00000012, 5'd12, 27'h000003b3, 32'h00000400,
  1'd1,  5'd2, 27'h000000b9, 5'd20, 27'h0000035f, 5'd22, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000e7, 5'd1, 27'h0000015f, 5'd2, 27'h000001fe, 32'h00000400,
  1'd1,  5'd13, 27'h00000020, 5'd1, 27'h00000305, 5'd10, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000020b, 5'd5, 27'h0000002f, 5'd23, 27'h0000025b, 32'h00000400,
  1'd1,  5'd11, 27'h000001c3, 5'd12, 27'h000003d2, 5'd4, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000242, 5'd11, 27'h00000034, 5'd10, 27'h00000231, 32'h00000400,
  1'd1,  5'd12, 27'h00000063, 5'd15, 27'h0000002d, 5'd24, 27'h000000c9, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000344, 5'd22, 27'h000003b0, 5'd3, 27'h000003b7, 32'h00000400,
  1'd1,  5'd12, 27'h00000224, 5'd23, 27'h000001a0, 5'd15, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000357, 5'd20, 27'h000002b0, 5'd25, 27'h000000b9, 32'h00000400,
  1'd1,  5'd23, 27'h00000162, 5'd0, 27'h000001f2, 5'd3, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e0, 5'd3, 27'h000001a5, 5'd14, 27'h00000132, 32'h00000400,
  1'd1,  5'd21, 27'h00000159, 5'd5, 27'h00000058, 5'd23, 27'h000002ad, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000025b, 5'd14, 27'h000001fe, 5'd2, 27'h0000020e, 32'h00000400,
  1'd1,  5'd24, 27'h0000026e, 5'd13, 27'h00000140, 5'd10, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000021a, 5'd14, 27'h00000184, 5'd22, 27'h0000015f, 32'h00000400,
  1'd1,  5'd21, 27'h00000192, 5'd23, 27'h000003bf, 5'd1, 27'h000000d5, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ac, 5'd23, 27'h0000021b, 5'd11, 27'h000002eb, 32'h00000400,
  1'd1,  5'd23, 27'h000002ce, 5'd25, 27'h00000204, 5'd22, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000389, 5'd3, 27'h00000142, 5'd7, 27'h0000005f, 32'h00000400,
  1'd1,  5'd1, 27'h0000010f, 5'd2, 27'h000002b5, 5'd19, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002d4, 5'd1, 27'h00000355, 5'd29, 27'h00000326, 32'h00000400,
  1'd1,  5'd2, 27'h0000005d, 5'd10, 27'h00000225, 5'd5, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000365, 5'd13, 27'h00000276, 5'd17, 27'h0000031e, 32'h00000400,
  1'd1,  5'd5, 27'h00000027, 5'd13, 27'h0000022d, 5'd29, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000e6, 5'd21, 27'h0000036a, 5'd9, 27'h00000346, 32'h00000400,
  1'd1,  5'd5, 27'h00000052, 5'd23, 27'h00000247, 5'd18, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000056, 5'd21, 27'h00000264, 5'd29, 27'h0000014c, 32'h00000400,
  1'd1,  5'd15, 27'h000001de, 5'd3, 27'h00000082, 5'd8, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017b, 5'd5, 27'h0000005c, 5'd18, 27'h00000341, 32'h00000400,
  1'd1,  5'd10, 27'h00000242, 5'd3, 27'h00000280, 5'd28, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000370, 5'd13, 27'h000001dd, 5'd8, 27'h00000265, 32'h00000400,
  1'd1,  5'd12, 27'h000003e4, 5'd14, 27'h00000098, 5'd20, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001d5, 5'd13, 27'h000000c8, 5'd27, 27'h00000169, 32'h00000400,
  1'd1,  5'd15, 27'h0000006b, 5'd24, 27'h000000b4, 5'd9, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025b, 5'd25, 27'h0000005d, 5'd18, 27'h0000018b, 32'h00000400,
  1'd1,  5'd15, 27'h00000022, 5'd25, 27'h000002c3, 5'd28, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000d4, 5'd2, 27'h0000017c, 5'd9, 27'h0000026f, 32'h00000400,
  1'd1,  5'd23, 27'h00000021, 5'd1, 27'h000003eb, 5'd19, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000025c, 5'd0, 27'h000000c3, 5'd27, 27'h000000d8, 32'h00000400,
  1'd1,  5'd20, 27'h00000399, 5'd14, 27'h0000010c, 5'd10, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000392, 5'd14, 27'h0000008c, 5'd20, 27'h0000029b, 32'h00000400,
  1'd1,  5'd25, 27'h00000128, 5'd12, 27'h000003bb, 5'd29, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000072, 5'd22, 27'h0000020e, 5'd7, 27'h000003dc, 32'h00000400,
  1'd1,  5'd21, 27'h00000285, 5'd22, 27'h0000007e, 5'd15, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000024d, 5'd24, 27'h000000d1, 5'd29, 27'h00000124, 32'h00000400,
  1'd1,  5'd0, 27'h00000332, 5'd7, 27'h000001f0, 5'd2, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002e, 5'd6, 27'h0000022c, 5'd14, 27'h000001d4, 32'h00000400,
  1'd1,  5'd3, 27'h00000320, 5'd8, 27'h00000113, 5'd22, 27'h000001bc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000127, 5'd17, 27'h000002fb, 5'd1, 27'h00000022, 32'h00000400,
  1'd1,  5'd3, 27'h00000339, 5'd19, 27'h00000071, 5'd15, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000010d, 5'd17, 27'h000000d6, 5'd21, 27'h000001ba, 32'h00000400,
  1'd1,  5'd4, 27'h00000269, 5'd28, 27'h000002ee, 5'd2, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000018a, 5'd28, 27'h0000007d, 5'd13, 27'h000002e2, 32'h00000400,
  1'd1,  5'd4, 27'h00000241, 5'd28, 27'h00000104, 5'd25, 27'h000001f6, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001e5, 5'd6, 27'h000000ec, 5'd1, 27'h0000021f, 32'h00000400,
  1'd1,  5'd15, 27'h0000004c, 5'd7, 27'h000001ae, 5'd12, 27'h00000069, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000b7, 5'd9, 27'h0000016d, 5'd25, 27'h0000000a, 32'h00000400,
  1'd1,  5'd10, 27'h0000024d, 5'd16, 27'h0000011d, 5'd3, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d2, 5'd18, 27'h0000031e, 5'd13, 27'h000001b3, 32'h00000400,
  1'd1,  5'd11, 27'h000003fb, 5'd18, 27'h000002e2, 5'd21, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000010f, 5'd30, 27'h00000284, 5'd2, 27'h0000011f, 32'h00000400,
  1'd1,  5'd12, 27'h00000055, 5'd26, 27'h000000d7, 5'd13, 27'h000002ea, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000030, 5'd26, 27'h00000040, 5'd20, 27'h0000037c, 32'h00000400,
  1'd1,  5'd20, 27'h000003ed, 5'd8, 27'h000003e5, 5'd2, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000017a, 5'd6, 27'h000001f4, 5'd15, 27'h000001a7, 32'h00000400,
  1'd1,  5'd22, 27'h000000c7, 5'd15, 27'h000003a5, 5'd3, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000f8, 5'd19, 27'h00000314, 5'd10, 27'h000003fa, 32'h00000400,
  1'd1,  5'd22, 27'h00000268, 5'd19, 27'h0000019d, 5'd23, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000035b, 5'd29, 27'h0000030b, 5'd1, 27'h0000028b, 32'h00000400,
  1'd1,  5'd22, 27'h0000024c, 5'd26, 27'h000002a1, 5'd15, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002c6, 5'd28, 27'h00000356, 5'd21, 27'h0000005c, 32'h00000400,
  1'd1,  5'd1, 27'h00000239, 5'd10, 27'h0000002f, 5'd5, 27'h0000031d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000038b, 5'd7, 27'h000003b2, 5'd20, 27'h000001ab, 32'h00000400,
  1'd1,  5'd0, 27'h00000273, 5'd6, 27'h000001d1, 5'd28, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000168, 5'd16, 27'h000002ba, 5'd8, 27'h000003ae, 32'h00000400,
  1'd1,  5'd1, 27'h00000018, 5'd20, 27'h000000a8, 5'd17, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000ae, 5'd16, 27'h000001aa, 5'd27, 27'h000001ad, 32'h00000400,
  1'd1,  5'd3, 27'h00000081, 5'd29, 27'h00000160, 5'd5, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000005, 5'd30, 27'h000003f6, 5'd18, 27'h0000026a, 32'h00000400,
  1'd1,  5'd3, 27'h000000d4, 5'd29, 27'h000000ea, 5'd26, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000162, 5'd9, 27'h0000000f, 5'd9, 27'h000001f5, 32'h00000400,
  1'd1,  5'd10, 27'h000003e7, 5'd8, 27'h00000038, 5'd16, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000270, 5'd6, 27'h000003b1, 5'd28, 27'h0000024e, 32'h00000400,
  1'd1,  5'd13, 27'h000002f9, 5'd16, 27'h0000033b, 5'd8, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000000e, 5'd15, 27'h000003eb, 5'd17, 27'h0000035d, 32'h00000400,
  1'd1,  5'd14, 27'h000003ff, 5'd17, 27'h000002b9, 5'd30, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000016, 5'd29, 27'h000002d1, 5'd7, 27'h0000026b, 32'h00000400,
  1'd1,  5'd11, 27'h00000102, 5'd30, 27'h0000033a, 5'd17, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d3, 5'd27, 27'h0000006a, 5'd29, 27'h000001ab, 32'h00000400,
  1'd1,  5'd25, 27'h000001b2, 5'd8, 27'h000002df, 5'd9, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001fb, 5'd7, 27'h0000024b, 5'd20, 27'h00000108, 32'h00000400,
  1'd1,  5'd22, 27'h000000ab, 5'd9, 27'h0000013c, 5'd27, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000021b, 5'd18, 27'h00000313, 5'd9, 27'h00000132, 32'h00000400,
  1'd1,  5'd21, 27'h0000014d, 5'd18, 27'h0000014f, 5'd19, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000030c, 5'd17, 27'h00000353, 5'd28, 27'h00000035, 32'h00000400,
  1'd1,  5'd24, 27'h0000027e, 5'd27, 27'h0000033b, 5'd9, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ca, 5'd26, 27'h000001d3, 5'd15, 27'h00000306, 32'h00000400,
  1'd1,  5'd21, 27'h000002df, 5'd27, 27'h000003c8, 5'd29, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001ac, 5'd2, 27'h00000288, 5'd5, 27'h000002f9, 32'h00000400,
  1'd1,  5'd6, 27'h00000244, 5'd2, 27'h00000102, 5'd19, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000024b, 5'd3, 27'h000000be, 5'd27, 27'h000002af, 32'h00000400,
  1'd1,  5'd7, 27'h00000351, 5'd12, 27'h000000bf, 5'd0, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003ff, 5'd12, 27'h00000225, 5'd11, 27'h000000b5, 32'h00000400,
  1'd1,  5'd5, 27'h000000e2, 5'd12, 27'h00000035, 5'd25, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000214, 5'd20, 27'h000003e3, 5'd1, 27'h00000391, 32'h00000400,
  1'd1,  5'd6, 27'h00000368, 5'd24, 27'h000002ff, 5'd14, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000036b, 5'd22, 27'h0000024c, 5'd20, 27'h000002dc, 32'h00000400,
  1'd1,  5'd18, 27'h00000351, 5'd3, 27'h0000031d, 5'd8, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000017f, 5'd2, 27'h000000c2, 5'd19, 27'h00000201, 32'h00000400,
  1'd1,  5'd19, 27'h000002b0, 5'd3, 27'h00000187, 5'd27, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000299, 5'd13, 27'h0000000d, 5'd5, 27'h0000000a, 32'h00000400,
  1'd1,  5'd18, 27'h00000224, 5'd12, 27'h0000019e, 5'd10, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000400, 5'd10, 27'h000003f8, 5'd22, 27'h00000320, 32'h00000400,
  1'd1,  5'd17, 27'h000000c4, 5'd21, 27'h00000138, 5'd0, 27'h000002a1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003fa, 5'd21, 27'h0000001e, 5'd11, 27'h000002f9, 32'h00000400,
  1'd1,  5'd16, 27'h0000028b, 5'd24, 27'h00000157, 5'd20, 27'h000003d2, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000032e, 5'd0, 27'h0000031f, 5'd2, 27'h00000129, 32'h00000400,
  1'd1,  5'd30, 27'h00000003, 5'd2, 27'h000003d1, 5'd14, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000077, 5'd4, 27'h000000f9, 5'd21, 27'h0000020b, 32'h00000400,
  1'd1,  5'd28, 27'h0000007c, 5'd11, 27'h00000355, 5'd0, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000297, 5'd12, 27'h000002b4, 5'd14, 27'h0000025e, 32'h00000400,
  1'd1,  5'd26, 27'h00000173, 5'd13, 27'h00000328, 5'd22, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002e3, 5'd21, 27'h00000220, 5'd0, 27'h00000392, 32'h00000400,
  1'd1,  5'd29, 27'h00000028, 5'd22, 27'h00000229, 5'd13, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000392, 5'd21, 27'h0000027b, 5'd21, 27'h0000011f, 32'h00000400,
  1'd1,  5'd5, 27'h000002f3, 5'd2, 27'h0000006d, 5'd4, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000b8, 5'd4, 27'h0000028f, 5'd10, 27'h000001af, 32'h00000400,
  1'd1,  5'd8, 27'h000002d9, 5'd2, 27'h000000b4, 5'd25, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000dc, 5'd11, 27'h00000123, 5'd6, 27'h00000349, 32'h00000400,
  1'd1,  5'd5, 27'h00000242, 5'd14, 27'h0000004a, 5'd16, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000157, 5'd13, 27'h000001fd, 5'd26, 27'h00000355, 32'h00000400,
  1'd1,  5'd5, 27'h000001af, 5'd22, 27'h00000303, 5'd6, 27'h00000023, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003ff, 5'd25, 27'h00000324, 5'd20, 27'h0000026a, 32'h00000400,
  1'd1,  5'd5, 27'h00000342, 5'd22, 27'h000001ac, 5'd30, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001fc, 5'd2, 27'h00000077, 5'd4, 27'h000001e5, 32'h00000400,
  1'd1,  5'd17, 27'h000002f1, 5'd5, 27'h00000048, 5'd13, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000007b, 5'd2, 27'h000002b9, 5'd21, 27'h00000307, 32'h00000400,
  1'd1,  5'd17, 27'h00000139, 5'd10, 27'h0000035a, 5'd7, 27'h000001a4, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000020a, 5'd11, 27'h00000049, 5'd16, 27'h00000356, 32'h00000400,
  1'd1,  5'd18, 27'h0000038a, 5'd15, 27'h00000170, 5'd28, 27'h000002dc, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000006a, 5'd20, 27'h000003dc, 5'd7, 27'h000002d4, 32'h00000400,
  1'd1,  5'd15, 27'h00000338, 5'd24, 27'h000003b6, 5'd15, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000266, 5'd23, 27'h000003e6, 5'd30, 27'h00000064, 32'h00000400,
  1'd1,  5'd30, 27'h000003c3, 5'd5, 27'h00000098, 5'd10, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003de, 5'd4, 27'h000001b6, 5'd17, 27'h0000013e, 32'h00000400,
  1'd1,  5'd27, 27'h00000111, 5'd1, 27'h00000047, 5'd29, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000038f, 5'd10, 27'h000001f7, 5'd8, 27'h000003e6, 32'h00000400,
  1'd1,  5'd26, 27'h000001fb, 5'd10, 27'h0000015c, 5'd16, 27'h0000025b, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003e1, 5'd12, 27'h00000302, 5'd28, 27'h000002f3, 32'h00000400,
  1'd1,  5'd26, 27'h0000026d, 5'd24, 27'h000002d2, 5'd6, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002c2, 5'd21, 27'h00000321, 5'd19, 27'h0000033a, 32'h00000400,
  1'd1,  5'd28, 27'h000003ed, 5'd21, 27'h00000050, 5'd30, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002fc, 5'd8, 27'h000001ac, 5'd3, 27'h00000245, 32'h00000400,
  1'd1,  5'd8, 27'h0000021a, 5'd9, 27'h0000020d, 5'd13, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a5, 5'd6, 27'h0000028a, 5'd22, 27'h0000003b, 32'h00000400,
  1'd1,  5'd9, 27'h00000301, 5'd16, 27'h000000eb, 5'd1, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000300, 5'd15, 27'h000002e1, 5'd13, 27'h00000248, 32'h00000400,
  1'd1,  5'd10, 27'h00000128, 5'd20, 27'h000000cc, 5'd21, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000015c, 5'd28, 27'h000003c6, 5'd4, 27'h000003a4, 32'h00000400,
  1'd1,  5'd9, 27'h000001d6, 5'd28, 27'h0000004e, 5'd12, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000057, 5'd29, 27'h00000005, 5'd22, 27'h000003f5, 32'h00000400,
  1'd1,  5'd20, 27'h00000006, 5'd5, 27'h000002e9, 5'd4, 27'h0000025f, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000036d, 5'd6, 27'h000002cf, 5'd11, 27'h00000264, 32'h00000400,
  1'd1,  5'd16, 27'h000001d6, 5'd5, 27'h000003fe, 5'd24, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000367, 5'd20, 27'h0000019b, 5'd1, 27'h000002f4, 32'h00000400,
  1'd1,  5'd18, 27'h000001f0, 5'd17, 27'h000000b0, 5'd12, 27'h0000019f, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000036a, 5'd20, 27'h0000016c, 5'd24, 27'h00000220, 32'h00000400,
  1'd1,  5'd16, 27'h000000c2, 5'd27, 27'h00000192, 5'd3, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002dc, 5'd25, 27'h00000390, 5'd13, 27'h00000249, 32'h00000400,
  1'd1,  5'd15, 27'h000003c0, 5'd28, 27'h000002e2, 5'd25, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000029f, 5'd5, 27'h0000036e, 5'd4, 27'h00000103, 32'h00000400,
  1'd1,  5'd28, 27'h000003fb, 5'd7, 27'h000002dd, 5'd12, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000130, 5'd10, 27'h0000013b, 5'd23, 27'h000001dd, 32'h00000400,
  1'd1,  5'd30, 27'h000001ae, 5'd17, 27'h000000cd, 5'd2, 27'h00000112, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000020a, 5'd18, 27'h000001de, 5'd12, 27'h000001bb, 32'h00000400,
  1'd1,  5'd28, 27'h00000114, 5'd20, 27'h00000071, 5'd24, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000f2, 5'd26, 27'h000001de, 5'd3, 27'h00000173, 32'h00000400,
  1'd1,  5'd26, 27'h00000092, 5'd29, 27'h00000370, 5'd15, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002fd, 5'd26, 27'h0000024f, 5'd22, 27'h0000023b, 32'h00000400,
  1'd1,  5'd9, 27'h00000048, 5'd8, 27'h000003a9, 5'd6, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000120, 5'd9, 27'h0000026f, 5'd20, 27'h00000167, 32'h00000400,
  1'd1,  5'd6, 27'h000001e2, 5'd5, 27'h00000318, 5'd26, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000155, 5'd18, 27'h0000011b, 5'd8, 27'h00000313, 32'h00000400,
  1'd1,  5'd7, 27'h00000026, 5'd18, 27'h00000255, 5'd20, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd9, 27'h000001dc, 5'd16, 27'h0000039c, 5'd29, 27'h0000018c, 32'h00000400,
  1'd1,  5'd6, 27'h000001b6, 5'd29, 27'h00000198, 5'd9, 27'h000003e6, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000358, 5'd27, 27'h000003ad, 5'd19, 27'h00000022, 32'h00000400,
  1'd1,  5'd6, 27'h0000039d, 5'd30, 27'h000002ab, 5'd29, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000220, 5'd9, 27'h00000179, 5'd8, 27'h00000121, 32'h00000400,
  1'd1,  5'd15, 27'h00000339, 5'd7, 27'h000003a5, 5'd15, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002d6, 5'd6, 27'h00000225, 5'd26, 27'h0000031f, 32'h00000400,
  1'd1,  5'd17, 27'h000001b1, 5'd19, 27'h0000038b, 5'd9, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000291, 5'd20, 27'h000000dc, 5'd19, 27'h0000001f, 32'h00000400,
  1'd1,  5'd15, 27'h000002f7, 5'd16, 27'h00000043, 5'd30, 27'h00000157, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031e, 5'd28, 27'h00000002, 5'd7, 27'h000000db, 32'h00000400,
  1'd1,  5'd20, 27'h00000010, 5'd28, 27'h00000166, 5'd16, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000041, 5'd28, 27'h000000f8, 5'd30, 27'h000003b8, 32'h00000400,
  1'd1,  5'd27, 27'h0000032e, 5'd7, 27'h00000302, 5'd9, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000018b, 5'd6, 27'h00000189, 5'd19, 27'h000001c8, 32'h00000400,
  1'd1,  5'd29, 27'h000001c7, 5'd8, 27'h000000cd, 5'd28, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000265, 5'd19, 27'h000002e9, 5'd10, 27'h000000fc, 32'h00000400,
  1'd1,  5'd27, 27'h00000341, 5'd20, 27'h00000008, 5'd20, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000057, 5'd16, 27'h0000024e, 5'd30, 27'h00000226, 32'h00000400,
  1'd1,  5'd29, 27'h00000022, 5'd27, 27'h000000ff, 5'd8, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000002e, 5'd27, 27'h00000234, 5'd17, 27'h00000105, 32'h00000400,
  1'd1,  5'd29, 27'h0000021b, 5'd30, 27'h00000285, 5'd27, 27'h000002b8, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd0, 27'h00000143, 5'd0, 27'h000003e2, 5'd3, 27'h00000010, 32'h00000400,
  1'd1,  5'd1, 27'h00000159, 5'd3, 27'h0000011f, 5'd13, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003d9, 5'd0, 27'h00000153, 5'd25, 27'h0000027c, 32'h00000400,
  1'd1,  5'd3, 27'h00000323, 5'd12, 27'h000003fe, 5'd0, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020d, 5'd10, 27'h000002c0, 5'd13, 27'h00000228, 32'h00000400,
  1'd1,  5'd1, 27'h000002f0, 5'd12, 27'h000003e9, 5'd22, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001f5, 5'd21, 27'h00000076, 5'd3, 27'h000002e6, 32'h00000400,
  1'd1,  5'd0, 27'h000000d0, 5'd24, 27'h0000024e, 5'd10, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000171, 5'd24, 27'h000000ff, 5'd22, 27'h000002f5, 32'h00000400,
  1'd1,  5'd12, 27'h00000287, 5'd4, 27'h000002fe, 5'd0, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000007c, 5'd0, 27'h00000287, 5'd12, 27'h0000018e, 32'h00000400,
  1'd1,  5'd11, 27'h00000022, 5'd0, 27'h0000013e, 5'd22, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ac, 5'd10, 27'h000001e6, 5'd2, 27'h00000121, 32'h00000400,
  1'd1,  5'd13, 27'h000002f7, 5'd11, 27'h0000023f, 5'd12, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000032f, 5'd11, 27'h00000223, 5'd22, 27'h0000039d, 32'h00000400,
  1'd1,  5'd14, 27'h00000179, 5'd23, 27'h000001e3, 5'd1, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000386, 5'd21, 27'h000000e9, 5'd14, 27'h000003f1, 32'h00000400,
  1'd1,  5'd10, 27'h000001c1, 5'd24, 27'h00000361, 5'd23, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000006a, 5'd1, 27'h000003b4, 5'd4, 27'h0000004e, 32'h00000400,
  1'd1,  5'd24, 27'h000001a5, 5'd2, 27'h000000e8, 5'd15, 27'h00000035, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000169, 5'd3, 27'h0000015e, 5'd24, 27'h00000304, 32'h00000400,
  1'd1,  5'd23, 27'h00000015, 5'd14, 27'h00000195, 5'd3, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000043, 5'd15, 27'h0000004d, 5'd10, 27'h00000333, 32'h00000400,
  1'd1,  5'd22, 27'h00000102, 5'd12, 27'h00000230, 5'd23, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000247, 5'd23, 27'h000003b8, 5'd3, 27'h00000206, 32'h00000400,
  1'd1,  5'd20, 27'h000002b7, 5'd23, 27'h0000026d, 5'd15, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000202, 5'd24, 27'h0000000d, 5'd21, 27'h00000357, 32'h00000400,
  1'd1,  5'd4, 27'h000002e4, 5'd1, 27'h0000036e, 5'd5, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001bf, 5'd3, 27'h00000314, 5'd18, 27'h0000008f, 32'h00000400,
  1'd1,  5'd4, 27'h00000230, 5'd5, 27'h0000001e, 5'd27, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000032b, 5'd12, 27'h000000b6, 5'd5, 27'h0000031d, 32'h00000400,
  1'd1,  5'd3, 27'h0000031c, 5'd13, 27'h000000ca, 5'd18, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f2, 5'd13, 27'h0000036c, 5'd30, 27'h0000038a, 32'h00000400,
  1'd1,  5'd1, 27'h00000309, 5'd21, 27'h000002be, 5'd8, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000097, 5'd22, 27'h00000180, 5'd18, 27'h0000018e, 32'h00000400,
  1'd1,  5'd3, 27'h000002ad, 5'd23, 27'h00000226, 5'd28, 27'h00000373, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a9, 5'd2, 27'h000003da, 5'd6, 27'h00000173, 32'h00000400,
  1'd1,  5'd12, 27'h00000166, 5'd4, 27'h00000358, 5'd19, 27'h000000e5, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000012c, 5'd1, 27'h00000329, 5'd30, 27'h00000202, 32'h00000400,
  1'd1,  5'd11, 27'h000000e0, 5'd13, 27'h000002cf, 5'd9, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003cd, 5'd13, 27'h0000003d, 5'd16, 27'h000003f6, 32'h00000400,
  1'd1,  5'd13, 27'h0000010b, 5'd15, 27'h000001b3, 5'd29, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000281, 5'd24, 27'h00000082, 5'd6, 27'h000000d4, 32'h00000400,
  1'd1,  5'd15, 27'h000000e7, 5'd24, 27'h00000179, 5'd19, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001de, 5'd23, 27'h00000111, 5'd27, 27'h000000c5, 32'h00000400,
  1'd1,  5'd23, 27'h000002a2, 5'd0, 27'h000001cf, 5'd6, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000394, 5'd3, 27'h0000037c, 5'd20, 27'h0000024d, 32'h00000400,
  1'd1,  5'd25, 27'h000000e1, 5'd3, 27'h00000337, 5'd27, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e0, 5'd11, 27'h0000028d, 5'd6, 27'h0000012e, 32'h00000400,
  1'd1,  5'd21, 27'h000003ec, 5'd13, 27'h000001d2, 5'd15, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000237, 5'd11, 27'h000003dd, 5'd27, 27'h000002c4, 32'h00000400,
  1'd1,  5'd23, 27'h00000027, 5'd25, 27'h00000292, 5'd9, 27'h00000307, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000260, 5'd22, 27'h0000018b, 5'd15, 27'h0000029d, 32'h00000400,
  1'd1,  5'd23, 27'h00000271, 5'd24, 27'h00000377, 5'd29, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000351, 5'd5, 27'h000002dc, 5'd0, 27'h00000259, 32'h00000400,
  1'd1,  5'd2, 27'h00000134, 5'd8, 27'h00000336, 5'd15, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036f, 5'd10, 27'h000000b6, 5'd24, 27'h00000114, 32'h00000400,
  1'd1,  5'd4, 27'h000001ea, 5'd15, 27'h00000340, 5'd0, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003c3, 5'd16, 27'h000003cc, 5'd10, 27'h00000365, 32'h00000400,
  1'd1,  5'd1, 27'h00000080, 5'd17, 27'h00000119, 5'd24, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002f, 5'd29, 27'h00000205, 5'd3, 27'h00000050, 32'h00000400,
  1'd1,  5'd2, 27'h000003b2, 5'd28, 27'h00000083, 5'd12, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000004d, 5'd29, 27'h000000b3, 5'd23, 27'h0000037e, 32'h00000400,
  1'd1,  5'd14, 27'h00000173, 5'd5, 27'h0000010d, 5'd0, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c6, 5'd9, 27'h000003b3, 5'd11, 27'h000003a7, 32'h00000400,
  1'd1,  5'd12, 27'h00000145, 5'd6, 27'h000002f3, 5'd22, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e5, 5'd19, 27'h00000252, 5'd2, 27'h0000035c, 32'h00000400,
  1'd1,  5'd14, 27'h00000093, 5'd18, 27'h0000009e, 5'd10, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002db, 5'd20, 27'h0000006d, 5'd22, 27'h0000026d, 32'h00000400,
  1'd1,  5'd12, 27'h000003e7, 5'd28, 27'h00000342, 5'd2, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000362, 5'd29, 27'h000003af, 5'd12, 27'h000001e9, 32'h00000400,
  1'd1,  5'd15, 27'h00000075, 5'd30, 27'h000002b0, 5'd24, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000151, 5'd6, 27'h00000046, 5'd4, 27'h000000db, 32'h00000400,
  1'd1,  5'd25, 27'h0000017a, 5'd7, 27'h00000077, 5'd12, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000350, 5'd20, 27'h000000e0, 5'd5, 27'h000000a3, 32'h00000400,
  1'd1,  5'd24, 27'h000001dc, 5'd16, 27'h0000003e, 5'd15, 27'h00000029, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000193, 5'd16, 27'h000001ac, 5'd24, 27'h000002cb, 32'h00000400,
  1'd1,  5'd21, 27'h00000111, 5'd28, 27'h000001d0, 5'd0, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000029, 5'd27, 27'h00000320, 5'd10, 27'h0000036a, 32'h00000400,
  1'd1,  5'd22, 27'h0000002a, 5'd27, 27'h000000ef, 5'd21, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000bb, 5'd9, 27'h0000010a, 5'd8, 27'h0000024d, 32'h00000400,
  1'd1,  5'd4, 27'h00000002, 5'd8, 27'h000001f9, 5'd17, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000028, 5'd8, 27'h00000220, 5'd30, 27'h00000382, 32'h00000400,
  1'd1,  5'd0, 27'h000000db, 5'd19, 27'h0000006b, 5'd9, 27'h000003c7, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003a2, 5'd18, 27'h0000021e, 5'd20, 27'h000001ec, 32'h00000400,
  1'd1,  5'd3, 27'h0000028f, 5'd19, 27'h00000030, 5'd26, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000031e, 5'd26, 27'h000002e1, 5'd9, 27'h00000189, 32'h00000400,
  1'd1,  5'd1, 27'h0000010c, 5'd26, 27'h000000ec, 5'd16, 27'h00000382, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000021a, 5'd28, 27'h0000001d, 5'd28, 27'h0000012b, 32'h00000400,
  1'd1,  5'd14, 27'h0000014a, 5'd10, 27'h000000b8, 5'd6, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d9, 5'd6, 27'h00000098, 5'd17, 27'h000001bb, 32'h00000400,
  1'd1,  5'd11, 27'h000002c6, 5'd7, 27'h000003de, 5'd26, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000027a, 5'd20, 27'h0000013c, 5'd8, 27'h000001f9, 32'h00000400,
  1'd1,  5'd12, 27'h000001dd, 5'd17, 27'h000002ec, 5'd20, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d4, 5'd16, 27'h00000269, 5'd26, 27'h00000166, 32'h00000400,
  1'd1,  5'd15, 27'h00000010, 5'd29, 27'h000003ce, 5'd6, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000127, 5'd30, 27'h0000035a, 5'd15, 27'h0000021d, 32'h00000400,
  1'd1,  5'd15, 27'h00000029, 5'd26, 27'h0000009b, 5'd27, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000133, 5'd6, 27'h000000dc, 5'd5, 27'h0000025a, 32'h00000400,
  1'd1,  5'd24, 27'h0000014c, 5'd7, 27'h00000033, 5'd18, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000c2, 5'd6, 27'h000002d2, 5'd27, 27'h00000285, 32'h00000400,
  1'd1,  5'd25, 27'h000002ba, 5'd18, 27'h000001ec, 5'd8, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000039d, 5'd18, 27'h000003cd, 5'd17, 27'h000000f6, 32'h00000400,
  1'd1,  5'd24, 27'h000000bb, 5'd19, 27'h000002cd, 5'd28, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c2, 5'd26, 27'h0000039a, 5'd6, 27'h000003a7, 32'h00000400,
  1'd1,  5'd21, 27'h000003be, 5'd30, 27'h0000036c, 5'd16, 27'h00000028, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b9, 5'd26, 27'h00000220, 5'd27, 27'h000002d4, 32'h00000400,
  1'd1,  5'd8, 27'h00000389, 5'd3, 27'h0000007c, 5'd5, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002bd, 5'd1, 27'h00000123, 5'd15, 27'h0000036e, 32'h00000400,
  1'd1,  5'd6, 27'h000000e0, 5'd4, 27'h000001b2, 5'd27, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002f5, 5'd12, 27'h00000247, 5'd1, 27'h00000058, 32'h00000400,
  1'd1,  5'd8, 27'h0000033d, 5'd11, 27'h0000017d, 5'd11, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000173, 5'd13, 27'h00000270, 5'd20, 27'h000002d9, 32'h00000400,
  1'd1,  5'd5, 27'h0000039a, 5'd21, 27'h00000292, 5'd4, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002e0, 5'd21, 27'h00000095, 5'd14, 27'h00000060, 32'h00000400,
  1'd1,  5'd9, 27'h00000021, 5'd24, 27'h00000265, 5'd23, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000242, 5'd1, 27'h000000a2, 5'd6, 27'h000001a6, 32'h00000400,
  1'd1,  5'd18, 27'h0000022b, 5'd2, 27'h00000232, 5'd16, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001a1, 5'd0, 27'h0000035e, 5'd29, 27'h00000086, 32'h00000400,
  1'd1,  5'd16, 27'h0000024c, 5'd10, 27'h00000390, 5'd0, 27'h00000260, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000400, 5'd13, 27'h000002ba, 5'd11, 27'h000002a3, 32'h00000400,
  1'd1,  5'd17, 27'h0000025c, 5'd12, 27'h00000187, 5'd23, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000317, 5'd25, 27'h0000006f, 5'd3, 27'h00000074, 32'h00000400,
  1'd1,  5'd19, 27'h00000088, 5'd25, 27'h0000026a, 5'd13, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000021a, 5'd22, 27'h00000119, 5'd25, 27'h000000dc, 32'h00000400,
  1'd1,  5'd29, 27'h0000006c, 5'd1, 27'h00000200, 5'd3, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000343, 5'd4, 27'h00000313, 5'd14, 27'h00000233, 32'h00000400,
  1'd1,  5'd30, 27'h0000019c, 5'd2, 27'h000002be, 5'd20, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002a3, 5'd11, 27'h00000156, 5'd2, 27'h00000052, 32'h00000400,
  1'd1,  5'd29, 27'h00000222, 5'd12, 27'h000001df, 5'd12, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000011e, 5'd14, 27'h0000027b, 5'd20, 27'h00000309, 32'h00000400,
  1'd1,  5'd27, 27'h000003f6, 5'd24, 27'h00000315, 5'd3, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000270, 5'd22, 27'h00000287, 5'd12, 27'h000001d7, 32'h00000400,
  1'd1,  5'd28, 27'h000002f9, 5'd23, 27'h0000032f, 5'd22, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000372, 5'd0, 27'h0000006b, 5'd1, 27'h000003f1, 32'h00000400,
  1'd1,  5'd8, 27'h00000336, 5'd2, 27'h0000020d, 5'd13, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000df, 5'd2, 27'h00000295, 5'd25, 27'h00000179, 32'h00000400,
  1'd1,  5'd9, 27'h00000053, 5'd12, 27'h000003c5, 5'd6, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000343, 5'd12, 27'h00000289, 5'd15, 27'h00000386, 32'h00000400,
  1'd1,  5'd9, 27'h000001fb, 5'd14, 27'h0000023f, 5'd28, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000278, 5'd25, 27'h000001b0, 5'd5, 27'h0000019d, 32'h00000400,
  1'd1,  5'd7, 27'h0000029b, 5'd24, 27'h0000001b, 5'd19, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000bb, 5'd21, 27'h0000004c, 5'd26, 27'h00000005, 32'h00000400,
  1'd1,  5'd18, 27'h00000352, 5'd2, 27'h0000035e, 5'd0, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000292, 5'd4, 27'h000000e2, 5'd10, 27'h00000295, 32'h00000400,
  1'd1,  5'd17, 27'h0000034b, 5'd0, 27'h000002f7, 5'd22, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000173, 5'd11, 27'h0000013f, 5'd10, 27'h000000f7, 32'h00000400,
  1'd1,  5'd18, 27'h000002d7, 5'd13, 27'h0000025b, 5'd17, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000097, 5'd11, 27'h000002e0, 5'd28, 27'h00000381, 32'h00000400,
  1'd1,  5'd16, 27'h000003b5, 5'd24, 27'h00000208, 5'd10, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003cd, 5'd22, 27'h0000017c, 5'd17, 27'h000001b5, 32'h00000400,
  1'd1,  5'd19, 27'h000002e2, 5'd23, 27'h000003f8, 5'd29, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b3, 5'd4, 27'h00000195, 5'd9, 27'h00000183, 32'h00000400,
  1'd1,  5'd30, 27'h00000052, 5'd3, 27'h000002e6, 5'd17, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000036, 5'd3, 27'h00000223, 5'd25, 27'h000003c8, 32'h00000400,
  1'd1,  5'd27, 27'h0000009f, 5'd10, 27'h0000032c, 5'd9, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000130, 5'd13, 27'h000003f8, 5'd18, 27'h000002aa, 32'h00000400,
  1'd1,  5'd28, 27'h000000f8, 5'd11, 27'h000000c8, 5'd28, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001ba, 5'd20, 27'h00000318, 5'd7, 27'h0000005a, 32'h00000400,
  1'd1,  5'd29, 27'h00000271, 5'd21, 27'h0000010e, 5'd16, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000039, 5'd21, 27'h000002f2, 5'd27, 27'h000002ca, 32'h00000400,
  1'd1,  5'd5, 27'h000000d4, 5'd6, 27'h000003c5, 5'd1, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000001d, 5'd9, 27'h000002df, 5'd15, 27'h0000016f, 32'h00000400,
  1'd1,  5'd5, 27'h00000336, 5'd9, 27'h00000305, 5'd23, 27'h000000d8, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000f3, 5'd18, 27'h0000035f, 5'd2, 27'h00000180, 32'h00000400,
  1'd1,  5'd9, 27'h000001aa, 5'd19, 27'h0000006a, 5'd10, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001a9, 5'd18, 27'h000000cc, 5'd21, 27'h000003df, 32'h00000400,
  1'd1,  5'd7, 27'h00000181, 5'd27, 27'h0000034c, 5'd4, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000239, 5'd29, 27'h000002a4, 5'd10, 27'h000003dd, 32'h00000400,
  1'd1,  5'd9, 27'h000003d1, 5'd25, 27'h000003ba, 5'd24, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000ff, 5'd5, 27'h000000da, 5'd0, 27'h000003fa, 32'h00000400,
  1'd1,  5'd17, 27'h000002f1, 5'd10, 27'h000000d9, 5'd13, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d3, 5'd6, 27'h0000011d, 5'd22, 27'h000000f6, 32'h00000400,
  1'd1,  5'd19, 27'h00000114, 5'd19, 27'h0000015a, 5'd3, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003a9, 5'd16, 27'h0000034e, 5'd13, 27'h00000187, 32'h00000400,
  1'd1,  5'd18, 27'h00000082, 5'd17, 27'h0000021e, 5'd21, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000030a, 5'd30, 27'h000003ef, 5'd0, 27'h000003a9, 32'h00000400,
  1'd1,  5'd16, 27'h00000250, 5'd27, 27'h000001ae, 5'd11, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000302, 5'd28, 27'h00000012, 5'd25, 27'h000000ca, 32'h00000400,
  1'd1,  5'd29, 27'h000003eb, 5'd9, 27'h00000256, 5'd1, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000375, 5'd5, 27'h0000026d, 5'd12, 27'h00000350, 32'h00000400,
  1'd1,  5'd29, 27'h0000038a, 5'd5, 27'h000000e5, 5'd23, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003ec, 5'd16, 27'h000001cf, 5'd0, 27'h00000306, 32'h00000400,
  1'd1,  5'd29, 27'h000002fa, 5'd17, 27'h0000037c, 5'd12, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000020d, 5'd16, 27'h000002e6, 5'd23, 27'h00000343, 32'h00000400,
  1'd1,  5'd27, 27'h000002e8, 5'd26, 27'h00000379, 5'd0, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000228, 5'd29, 27'h000002dc, 5'd14, 27'h0000022a, 32'h00000400,
  1'd1,  5'd27, 27'h0000001a, 5'd26, 27'h00000275, 5'd21, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000298, 5'd5, 27'h0000037d, 5'd8, 27'h0000006b, 32'h00000400,
  1'd1,  5'd7, 27'h0000025d, 5'd8, 27'h000002fa, 5'd16, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000006, 5'd10, 27'h00000032, 5'd28, 27'h00000123, 32'h00000400,
  1'd1,  5'd5, 27'h000003fd, 5'd20, 27'h00000121, 5'd6, 27'h00000340, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000123, 5'd16, 27'h00000079, 5'd20, 27'h000001ea, 32'h00000400,
  1'd1,  5'd8, 27'h0000016c, 5'd18, 27'h0000018b, 5'd30, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000128, 5'd30, 27'h000001b5, 5'd6, 27'h000003db, 32'h00000400,
  1'd1,  5'd8, 27'h0000003a, 5'd28, 27'h000002fc, 5'd17, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000059, 5'd28, 27'h0000026e, 5'd29, 27'h0000008e, 32'h00000400,
  1'd1,  5'd17, 27'h00000287, 5'd7, 27'h000002b3, 5'd8, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000037a, 5'd5, 27'h000003b8, 5'd16, 27'h0000011e, 32'h00000400,
  1'd1,  5'd16, 27'h00000159, 5'd8, 27'h000001bb, 5'd29, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001af, 5'd17, 27'h0000015d, 5'd5, 27'h0000029b, 32'h00000400,
  1'd1,  5'd16, 27'h00000047, 5'd16, 27'h00000374, 5'd18, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000018b, 5'd18, 27'h000001ad, 5'd28, 27'h000003d3, 32'h00000400,
  1'd1,  5'd19, 27'h0000038e, 5'd29, 27'h000000e3, 5'd8, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001c2, 5'd30, 27'h000002a4, 5'd18, 27'h0000036c, 32'h00000400,
  1'd1,  5'd16, 27'h0000002a, 5'd29, 27'h00000147, 5'd27, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000025f, 5'd6, 27'h00000350, 5'd6, 27'h000002b8, 32'h00000400,
  1'd1,  5'd28, 27'h000003b1, 5'd5, 27'h00000163, 5'd18, 27'h000001b7, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012e, 5'd7, 27'h000000ad, 5'd30, 27'h00000139, 32'h00000400,
  1'd1,  5'd29, 27'h00000209, 5'd16, 27'h000000b5, 5'd10, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000004d, 5'd16, 27'h000001dc, 5'd16, 27'h0000011a, 32'h00000400,
  1'd1,  5'd26, 27'h000003fc, 5'd16, 27'h00000179, 5'd28, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003e1, 5'd29, 27'h000001ba, 5'd8, 27'h00000178, 32'h00000400,
  1'd1,  5'd30, 27'h00000195, 5'd26, 27'h00000371, 5'd15, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000039a, 5'd29, 27'h00000026, 5'd29, 27'h0000018c, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h00000247, 5'd2, 27'h0000030b, 5'd3, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000015a, 5'd3, 27'h000002fa, 5'd15, 27'h000000c2, 32'h00000400,
  1'd1,  5'd0, 27'h0000009b, 5'd0, 27'h0000017d, 5'd21, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000376, 5'd11, 27'h000003a8, 5'd3, 27'h000002f3, 32'h00000400,
  1'd1,  5'd0, 27'h0000039a, 5'd14, 27'h00000061, 5'd13, 27'h000003fe, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000048, 5'd15, 27'h000001ce, 5'd21, 27'h00000158, 32'h00000400,
  1'd1,  5'd5, 27'h00000012, 5'd22, 27'h00000130, 5'd3, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000148, 5'd22, 27'h00000216, 5'd10, 27'h00000330, 32'h00000400,
  1'd1,  5'd2, 27'h000003da, 5'd24, 27'h000001a3, 5'd24, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002b1, 5'd3, 27'h0000024d, 5'd4, 27'h00000062, 32'h00000400,
  1'd1,  5'd11, 27'h00000235, 5'd1, 27'h00000018, 5'd15, 27'h0000015e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000283, 5'd4, 27'h00000050, 5'd21, 27'h00000029, 32'h00000400,
  1'd1,  5'd13, 27'h00000295, 5'd14, 27'h00000139, 5'd4, 27'h00000036, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000098, 5'd10, 27'h0000024c, 5'd11, 27'h000001d0, 32'h00000400,
  1'd1,  5'd13, 27'h00000231, 5'd15, 27'h000001cb, 5'd24, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000375, 5'd22, 27'h00000081, 5'd3, 27'h000002f7, 32'h00000400,
  1'd1,  5'd10, 27'h000002dc, 5'd21, 27'h000003be, 5'd11, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000015c, 5'd21, 27'h00000259, 5'd25, 27'h000002ee, 32'h00000400,
  1'd1,  5'd24, 27'h0000001c, 5'd3, 27'h00000383, 5'd0, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000255, 5'd3, 27'h0000006b, 5'd10, 27'h000003a5, 32'h00000400,
  1'd1,  5'd23, 27'h00000366, 5'd3, 27'h0000027c, 5'd23, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000013b, 5'd12, 27'h00000376, 5'd4, 27'h00000384, 32'h00000400,
  1'd1,  5'd25, 27'h00000257, 5'd14, 27'h000002d6, 5'd12, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000373, 5'd13, 27'h0000000f, 5'd23, 27'h000000cb, 32'h00000400,
  1'd1,  5'd21, 27'h00000093, 5'd24, 27'h00000002, 5'd0, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000b4, 5'd21, 27'h0000013b, 5'd14, 27'h00000216, 32'h00000400,
  1'd1,  5'd21, 27'h0000008c, 5'd24, 27'h00000270, 5'd21, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000b2, 5'd2, 27'h000000c9, 5'd5, 27'h00000373, 32'h00000400,
  1'd1,  5'd4, 27'h00000102, 5'd3, 27'h0000015a, 5'd16, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000028b, 5'd3, 27'h00000218, 5'd29, 27'h00000204, 32'h00000400,
  1'd1,  5'd4, 27'h00000011, 5'd14, 27'h00000322, 5'd9, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002cc, 5'd12, 27'h00000096, 5'd20, 27'h00000112, 32'h00000400,
  1'd1,  5'd1, 27'h00000056, 5'd11, 27'h00000325, 5'd28, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d7, 5'd23, 27'h0000038e, 5'd7, 27'h0000013f, 32'h00000400,
  1'd1,  5'd2, 27'h00000180, 5'd22, 27'h000003f8, 5'd17, 27'h000002fc, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001bf, 5'd23, 27'h0000025d, 5'd29, 27'h000000b8, 32'h00000400,
  1'd1,  5'd14, 27'h000000d4, 5'd2, 27'h00000197, 5'd10, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e5, 5'd2, 27'h00000061, 5'd16, 27'h000003a2, 32'h00000400,
  1'd1,  5'd13, 27'h000002ff, 5'd1, 27'h000002fb, 5'd27, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000108, 5'd11, 27'h00000082, 5'd7, 27'h00000079, 32'h00000400,
  1'd1,  5'd11, 27'h00000371, 5'd14, 27'h000003bd, 5'd20, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001e1, 5'd11, 27'h000001a4, 5'd27, 27'h0000033f, 32'h00000400,
  1'd1,  5'd11, 27'h00000109, 5'd21, 27'h000001ac, 5'd7, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ef, 5'd20, 27'h000002f0, 5'd16, 27'h00000197, 32'h00000400,
  1'd1,  5'd12, 27'h000000e8, 5'd24, 27'h0000009d, 5'd27, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003f6, 5'd4, 27'h000001f3, 5'd7, 27'h000000a1, 32'h00000400,
  1'd1,  5'd21, 27'h00000298, 5'd1, 27'h000001ec, 5'd19, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e9, 5'd2, 27'h0000022e, 5'd27, 27'h00000265, 32'h00000400,
  1'd1,  5'd24, 27'h00000208, 5'd15, 27'h000001ac, 5'd7, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bf, 5'd13, 27'h000002e3, 5'd16, 27'h000003c0, 32'h00000400,
  1'd1,  5'd22, 27'h00000012, 5'd15, 27'h00000153, 5'd28, 27'h00000163, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002d4, 5'd21, 27'h00000237, 5'd6, 27'h000003c6, 32'h00000400,
  1'd1,  5'd23, 27'h0000021b, 5'd21, 27'h000003c6, 5'd18, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002ef, 5'd22, 27'h000003e9, 5'd29, 27'h000000ea, 32'h00000400,
  1'd1,  5'd3, 27'h000003d6, 5'd7, 27'h0000017c, 5'd4, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000053, 5'd7, 27'h00000124, 5'd13, 27'h0000038b, 32'h00000400,
  1'd1,  5'd2, 27'h000001d6, 5'd5, 27'h000000ac, 5'd21, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000c6, 5'd20, 27'h000001ee, 5'd4, 27'h00000106, 32'h00000400,
  1'd1,  5'd0, 27'h000002f6, 5'd18, 27'h000002a1, 5'd12, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000322, 5'd19, 27'h000000ec, 5'd22, 27'h000000d7, 32'h00000400,
  1'd1,  5'd1, 27'h000001fc, 5'd26, 27'h00000060, 5'd1, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000400, 5'd28, 27'h000000ac, 5'd10, 27'h000001d6, 32'h00000400,
  1'd1,  5'd4, 27'h000001ac, 5'd27, 27'h0000022d, 5'd24, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000033f, 5'd9, 27'h000002f3, 5'd3, 27'h0000010a, 32'h00000400,
  1'd1,  5'd14, 27'h00000389, 5'd7, 27'h00000278, 5'd13, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000026c, 5'd6, 27'h00000218, 5'd20, 27'h0000031e, 32'h00000400,
  1'd1,  5'd14, 27'h000001d5, 5'd17, 27'h00000330, 5'd3, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000372, 5'd20, 27'h000001b6, 5'd13, 27'h000002ae, 32'h00000400,
  1'd1,  5'd11, 27'h000002a5, 5'd18, 27'h00000163, 5'd24, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000007c, 5'd26, 27'h0000034b, 5'd3, 27'h00000385, 32'h00000400,
  1'd1,  5'd10, 27'h00000160, 5'd27, 27'h00000189, 5'd10, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000015c, 5'd29, 27'h00000182, 5'd23, 27'h000002ba, 32'h00000400,
  1'd1,  5'd24, 27'h00000329, 5'd10, 27'h0000001b, 5'd1, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ab, 5'd9, 27'h000003a1, 5'd11, 27'h000001e5, 32'h00000400,
  1'd1,  5'd24, 27'h000000d9, 5'd20, 27'h00000147, 5'd1, 27'h000001a7, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002b1, 5'd18, 27'h00000236, 5'd10, 27'h0000032f, 32'h00000400,
  1'd1,  5'd22, 27'h0000019a, 5'd18, 27'h0000027a, 5'd23, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001f2, 5'd27, 27'h00000230, 5'd3, 27'h00000294, 32'h00000400,
  1'd1,  5'd24, 27'h000001ce, 5'd27, 27'h00000370, 5'd11, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000206, 5'd27, 27'h00000060, 5'd20, 27'h00000380, 32'h00000400,
  1'd1,  5'd0, 27'h00000112, 5'd7, 27'h0000016c, 5'd6, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000028d, 5'd9, 27'h00000248, 5'd19, 27'h00000078, 32'h00000400,
  1'd1,  5'd1, 27'h0000023e, 5'd5, 27'h000003b2, 5'd28, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000e3, 5'd19, 27'h00000203, 5'd9, 27'h000000ac, 32'h00000400,
  1'd1,  5'd3, 27'h0000031e, 5'd15, 27'h0000033f, 5'd16, 27'h00000327, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f1, 5'd17, 27'h00000375, 5'd29, 27'h0000002a, 32'h00000400,
  1'd1,  5'd1, 27'h0000020e, 5'd27, 27'h000001ba, 5'd6, 27'h00000330, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000023e, 5'd28, 27'h00000390, 5'd16, 27'h000000b7, 32'h00000400,
  1'd1,  5'd3, 27'h00000281, 5'd30, 27'h00000091, 5'd26, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000011c, 5'd8, 27'h00000342, 5'd9, 27'h00000390, 32'h00000400,
  1'd1,  5'd12, 27'h0000026c, 5'd9, 27'h000001cb, 5'd18, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000011a, 5'd9, 27'h00000196, 5'd29, 27'h00000104, 32'h00000400,
  1'd1,  5'd11, 27'h00000365, 5'd16, 27'h000001f5, 5'd7, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000228, 5'd20, 27'h000000ee, 5'd16, 27'h000000ac, 32'h00000400,
  1'd1,  5'd12, 27'h00000369, 5'd19, 27'h0000011b, 5'd27, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000057, 5'd28, 27'h000003cf, 5'd8, 27'h000000f1, 32'h00000400,
  1'd1,  5'd13, 27'h000002d3, 5'd30, 27'h00000038, 5'd17, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003cb, 5'd27, 27'h000003c5, 5'd25, 27'h000003f1, 32'h00000400,
  1'd1,  5'd25, 27'h00000075, 5'd7, 27'h0000013d, 5'd6, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a5, 5'd9, 27'h00000257, 5'd17, 27'h00000265, 32'h00000400,
  1'd1,  5'd23, 27'h000002c2, 5'd5, 27'h000001b5, 5'd26, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000023e, 5'd17, 27'h000000d7, 5'd9, 27'h000003fb, 32'h00000400,
  1'd1,  5'd25, 27'h00000011, 5'd19, 27'h00000004, 5'd17, 27'h00000268, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000375, 5'd17, 27'h000000e2, 5'd30, 27'h00000068, 32'h00000400,
  1'd1,  5'd22, 27'h000000c3, 5'd28, 27'h00000212, 5'd7, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000216, 5'd27, 27'h00000289, 5'd15, 27'h00000255, 32'h00000400,
  1'd1,  5'd25, 27'h000002bf, 5'd27, 27'h00000067, 5'd27, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000095, 5'd4, 27'h00000083, 5'd9, 27'h000000f8, 32'h00000400,
  1'd1,  5'd7, 27'h000001db, 5'd2, 27'h00000274, 5'd16, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000027b, 5'd1, 27'h000003ba, 5'd26, 27'h00000028, 32'h00000400,
  1'd1,  5'd9, 27'h00000132, 5'd12, 27'h00000057, 5'd1, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000128, 5'd14, 27'h000000bd, 5'd12, 27'h0000006c, 32'h00000400,
  1'd1,  5'd5, 27'h00000294, 5'd13, 27'h000003c1, 5'd22, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001d9, 5'd23, 27'h000001e3, 5'd2, 27'h0000004e, 32'h00000400,
  1'd1,  5'd7, 27'h00000216, 5'd24, 27'h00000155, 5'd12, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000015c, 5'd24, 27'h000003da, 5'd23, 27'h00000091, 32'h00000400,
  1'd1,  5'd19, 27'h00000056, 5'd0, 27'h000000f5, 5'd9, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000381, 5'd0, 27'h000003a3, 5'd20, 27'h00000275, 32'h00000400,
  1'd1,  5'd17, 27'h00000109, 5'd1, 27'h00000307, 5'd28, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003fe, 5'd10, 27'h000003ae, 5'd4, 27'h000002e3, 32'h00000400,
  1'd1,  5'd18, 27'h00000261, 5'd14, 27'h000000a7, 5'd13, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002f2, 5'd12, 27'h00000320, 5'd23, 27'h00000038, 32'h00000400,
  1'd1,  5'd16, 27'h0000030f, 5'd24, 27'h000001c7, 5'd0, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002cd, 5'd25, 27'h000002a4, 5'd14, 27'h0000039d, 32'h00000400,
  1'd1,  5'd16, 27'h000001d4, 5'd21, 27'h0000017c, 5'd21, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000029, 5'd1, 27'h00000052, 5'd3, 27'h000002c5, 32'h00000400,
  1'd1,  5'd28, 27'h000003c3, 5'd2, 27'h00000333, 5'd13, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b6, 5'd4, 27'h00000153, 5'd21, 27'h000000db, 32'h00000400,
  1'd1,  5'd25, 27'h000003a6, 5'd11, 27'h00000279, 5'd4, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000026a, 5'd10, 27'h00000208, 5'd12, 27'h00000134, 32'h00000400,
  1'd1,  5'd30, 27'h000001c7, 5'd13, 27'h00000320, 5'd25, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000331, 5'd21, 27'h00000115, 5'd2, 27'h00000331, 32'h00000400,
  1'd1,  5'd29, 27'h0000011a, 5'd21, 27'h0000024f, 5'd11, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000030f, 5'd23, 27'h000001b5, 5'd23, 27'h0000037a, 32'h00000400,
  1'd1,  5'd9, 27'h00000263, 5'd2, 27'h000001b1, 5'd0, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000231, 5'd4, 27'h00000308, 5'd13, 27'h000003af, 32'h00000400,
  1'd1,  5'd6, 27'h00000294, 5'd0, 27'h000001fb, 5'd25, 27'h000000f7, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003dc, 5'd13, 27'h00000118, 5'd9, 27'h000000c5, 32'h00000400,
  1'd1,  5'd7, 27'h0000016d, 5'd10, 27'h0000015f, 5'd16, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000216, 5'd12, 27'h000000ba, 5'd27, 27'h000000f6, 32'h00000400,
  1'd1,  5'd8, 27'h00000067, 5'd20, 27'h000003d9, 5'd7, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001a8, 5'd23, 27'h00000306, 5'd18, 27'h000000a0, 32'h00000400,
  1'd1,  5'd8, 27'h000001b4, 5'd21, 27'h000001bc, 5'd29, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002bd, 5'd1, 27'h000002ee, 5'd2, 27'h000001c0, 32'h00000400,
  1'd1,  5'd17, 27'h00000302, 5'd0, 27'h000003a9, 5'd15, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a6, 5'd0, 27'h000003ee, 5'd23, 27'h00000224, 32'h00000400,
  1'd1,  5'd18, 27'h00000207, 5'd13, 27'h00000008, 5'd8, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000214, 5'd14, 27'h00000302, 5'd18, 27'h00000029, 32'h00000400,
  1'd1,  5'd17, 27'h000003b9, 5'd14, 27'h0000003c, 5'd27, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002bf, 5'd25, 27'h00000338, 5'd9, 27'h00000048, 32'h00000400,
  1'd1,  5'd18, 27'h000000ea, 5'd20, 27'h0000039b, 5'd18, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000012c, 5'd25, 27'h00000184, 5'd26, 27'h000003a9, 32'h00000400,
  1'd1,  5'd29, 27'h000003db, 5'd0, 27'h0000017d, 5'd6, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000012e, 5'd0, 27'h0000015c, 5'd19, 27'h00000335, 32'h00000400,
  1'd1,  5'd27, 27'h0000035d, 5'd2, 27'h000003e6, 5'd30, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000032a, 5'd10, 27'h000002f5, 5'd10, 27'h000000b4, 32'h00000400,
  1'd1,  5'd30, 27'h0000012c, 5'd11, 27'h00000374, 5'd15, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000184, 5'd11, 27'h000000b5, 5'd28, 27'h000003e7, 32'h00000400,
  1'd1,  5'd27, 27'h0000014a, 5'd21, 27'h00000255, 5'd8, 27'h0000023f, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000036a, 5'd24, 27'h00000061, 5'd19, 27'h000002a2, 32'h00000400,
  1'd1,  5'd25, 27'h000003d8, 5'd24, 27'h0000002f, 5'd27, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000140, 5'd9, 27'h0000017a, 5'd2, 27'h000001c0, 32'h00000400,
  1'd1,  5'd8, 27'h000003a0, 5'd10, 27'h0000007f, 5'd13, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003f1, 5'd5, 27'h00000312, 5'd20, 27'h0000033d, 32'h00000400,
  1'd1,  5'd9, 27'h00000352, 5'd20, 27'h000000c5, 5'd0, 27'h00000063, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e5, 5'd16, 27'h000000d3, 5'd10, 27'h0000016c, 32'h00000400,
  1'd1,  5'd5, 27'h000000ff, 5'd16, 27'h0000030e, 5'd23, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000de, 5'd26, 27'h00000171, 5'd0, 27'h000003c5, 32'h00000400,
  1'd1,  5'd8, 27'h00000141, 5'd29, 27'h000000bd, 5'd11, 27'h0000018b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000173, 5'd27, 27'h0000013a, 5'd23, 27'h00000240, 32'h00000400,
  1'd1,  5'd16, 27'h00000286, 5'd6, 27'h0000020c, 5'd0, 27'h000001ea, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e0, 5'd7, 27'h0000018a, 5'd14, 27'h000003d5, 32'h00000400,
  1'd1,  5'd16, 27'h00000171, 5'd6, 27'h00000128, 5'd25, 27'h000002b5, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000127, 5'd18, 27'h000000e8, 5'd3, 27'h000002d7, 32'h00000400,
  1'd1,  5'd15, 27'h000002aa, 5'd20, 27'h000001d4, 5'd15, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000223, 5'd17, 27'h00000152, 5'd22, 27'h00000104, 32'h00000400,
  1'd1,  5'd17, 27'h00000139, 5'd28, 27'h000001e0, 5'd2, 27'h000003bb, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000aa, 5'd26, 27'h0000001c, 5'd13, 27'h000002ce, 32'h00000400,
  1'd1,  5'd16, 27'h00000220, 5'd28, 27'h00000147, 5'd24, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002c1, 5'd5, 27'h000001d7, 5'd0, 27'h000002e1, 32'h00000400,
  1'd1,  5'd30, 27'h00000216, 5'd7, 27'h0000018d, 5'd10, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000333, 5'd7, 27'h000001cf, 5'd23, 27'h00000336, 32'h00000400,
  1'd1,  5'd28, 27'h0000036b, 5'd17, 27'h000000c4, 5'd2, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000312, 5'd20, 27'h00000202, 5'd11, 27'h000001cb, 32'h00000400,
  1'd1,  5'd26, 27'h0000006b, 5'd19, 27'h0000013e, 5'd22, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000386, 5'd29, 27'h0000018c, 5'd0, 27'h0000038a, 32'h00000400,
  1'd1,  5'd25, 27'h00000392, 5'd29, 27'h000001ef, 5'd12, 27'h0000005f, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000020b, 5'd29, 27'h0000011f, 5'd23, 27'h0000009f, 32'h00000400,
  1'd1,  5'd7, 27'h0000027e, 5'd8, 27'h000000cd, 5'd10, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000023e, 5'd6, 27'h000002af, 5'd20, 27'h000000ad, 32'h00000400,
  1'd1,  5'd5, 27'h000003b4, 5'd9, 27'h000001ff, 5'd26, 27'h00000054, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002a4, 5'd16, 27'h00000261, 5'd7, 27'h000000f3, 32'h00000400,
  1'd1,  5'd5, 27'h000002f4, 5'd16, 27'h00000178, 5'd16, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000278, 5'd20, 27'h000001df, 5'd27, 27'h000000c1, 32'h00000400,
  1'd1,  5'd5, 27'h000003d8, 5'd30, 27'h00000001, 5'd9, 27'h0000019d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000199, 5'd26, 27'h00000236, 5'd20, 27'h00000156, 32'h00000400,
  1'd1,  5'd5, 27'h00000124, 5'd30, 27'h000003e0, 5'd28, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000170, 5'd5, 27'h00000231, 5'd8, 27'h0000017f, 32'h00000400,
  1'd1,  5'd16, 27'h0000003a, 5'd7, 27'h000002c0, 5'd18, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000364, 5'd7, 27'h00000290, 5'd28, 27'h000003d6, 32'h00000400,
  1'd1,  5'd17, 27'h000002d9, 5'd18, 27'h00000173, 5'd9, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000031a, 5'd17, 27'h000001c7, 5'd19, 27'h0000020e, 32'h00000400,
  1'd1,  5'd19, 27'h000001a3, 5'd17, 27'h000003fc, 5'd26, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000314, 5'd28, 27'h00000145, 5'd8, 27'h000001bf, 32'h00000400,
  1'd1,  5'd16, 27'h0000004d, 5'd30, 27'h000001c8, 5'd17, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000283, 5'd27, 27'h00000069, 5'd27, 27'h00000294, 32'h00000400,
  1'd1,  5'd29, 27'h00000045, 5'd10, 27'h000000a5, 5'd5, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000060, 5'd5, 27'h000003c7, 5'd17, 27'h00000256, 32'h00000400,
  1'd1,  5'd30, 27'h0000037b, 5'd9, 27'h000000f4, 5'd29, 27'h0000015f, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000000c, 5'd20, 27'h0000029a, 5'd6, 27'h000003fe, 32'h00000400,
  1'd1,  5'd28, 27'h00000252, 5'd19, 27'h000003d7, 5'd18, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000065, 5'd18, 27'h000000ae, 5'd27, 27'h0000028e, 32'h00000400,
  1'd1,  5'd30, 27'h000000fc, 5'd30, 27'h00000165, 5'd7, 27'h00000021, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000030b, 5'd29, 27'h0000006c, 5'd18, 27'h00000111, 32'h00000400,
  1'd1,  5'd28, 27'h0000031b, 5'd27, 27'h00000178, 5'd26, 27'h000000bf, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000000fa, 5'd2, 27'h000001d7, 5'd2, 27'h000001ec, 32'h00000400,
  1'd1,  5'd1, 27'h00000040, 5'd0, 27'h0000017e, 5'd13, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003c6, 5'd4, 27'h000002eb, 5'd20, 27'h000002d6, 32'h00000400,
  1'd1,  5'd1, 27'h00000230, 5'd10, 27'h0000015a, 5'd2, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000007e, 5'd11, 27'h00000101, 5'd11, 27'h00000016, 32'h00000400,
  1'd1,  5'd0, 27'h0000002c, 5'd11, 27'h000000cf, 5'd21, 27'h00000300, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b4, 5'd23, 27'h00000115, 5'd0, 27'h000001e5, 32'h00000400,
  1'd1,  5'd3, 27'h0000013c, 5'd22, 27'h00000201, 5'd14, 27'h000000b3, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002de, 5'd22, 27'h000003e8, 5'd24, 27'h0000007a, 32'h00000400,
  1'd1,  5'd15, 27'h00000140, 5'd5, 27'h000000a7, 5'd4, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000308, 5'd4, 27'h00000195, 5'd10, 27'h00000311, 32'h00000400,
  1'd1,  5'd15, 27'h000001fe, 5'd0, 27'h0000037f, 5'd21, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000041, 5'd10, 27'h0000024f, 5'd0, 27'h0000030f, 32'h00000400,
  1'd1,  5'd12, 27'h00000334, 5'd12, 27'h00000132, 5'd13, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003d0, 5'd12, 27'h00000234, 5'd24, 27'h0000030e, 32'h00000400,
  1'd1,  5'd12, 27'h0000007d, 5'd22, 27'h000003d7, 5'd3, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000007f, 5'd23, 27'h00000193, 5'd11, 27'h00000261, 32'h00000400,
  1'd1,  5'd12, 27'h000000c8, 5'd25, 27'h00000241, 5'd23, 27'h0000000a, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000000e, 5'd3, 27'h000002fe, 5'd2, 27'h000000a7, 32'h00000400,
  1'd1,  5'd21, 27'h00000182, 5'd1, 27'h00000309, 5'd12, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000213, 5'd4, 27'h00000358, 5'd23, 27'h0000002f, 32'h00000400,
  1'd1,  5'd25, 27'h00000317, 5'd12, 27'h0000016c, 5'd3, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000015e, 5'd14, 27'h000002fb, 5'd13, 27'h00000178, 32'h00000400,
  1'd1,  5'd25, 27'h000002ec, 5'd12, 27'h00000265, 5'd24, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000202, 5'd22, 27'h0000032e, 5'd2, 27'h000001ea, 32'h00000400,
  1'd1,  5'd21, 27'h000003d6, 5'd24, 27'h000000b5, 5'd10, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000001d, 5'd24, 27'h000000f0, 5'd21, 27'h0000006e, 32'h00000400,
  1'd1,  5'd4, 27'h0000006d, 5'd0, 27'h0000017d, 5'd7, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000015f, 5'd0, 27'h000001d8, 5'd19, 27'h00000203, 32'h00000400,
  1'd1,  5'd2, 27'h000000ab, 5'd2, 27'h00000203, 5'd28, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000c6, 5'd14, 27'h00000350, 5'd9, 27'h00000137, 32'h00000400,
  1'd1,  5'd3, 27'h000000c2, 5'd13, 27'h000001c7, 5'd20, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002af, 5'd13, 27'h00000063, 5'd30, 27'h00000069, 32'h00000400,
  1'd1,  5'd1, 27'h000000ca, 5'd22, 27'h000001ef, 5'd5, 27'h000002f2, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001e7, 5'd22, 27'h00000357, 5'd15, 27'h00000246, 32'h00000400,
  1'd1,  5'd5, 27'h00000072, 5'd20, 27'h00000368, 5'd27, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ee, 5'd3, 27'h000000c7, 5'd10, 27'h00000089, 32'h00000400,
  1'd1,  5'd10, 27'h000002a1, 5'd3, 27'h000001a6, 5'd18, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000028d, 5'd2, 27'h000003c4, 5'd28, 27'h000002e7, 32'h00000400,
  1'd1,  5'd12, 27'h0000017c, 5'd11, 27'h0000013b, 5'd7, 27'h000002fb, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000020c, 5'd11, 27'h000001b8, 5'd17, 27'h00000200, 32'h00000400,
  1'd1,  5'd15, 27'h00000078, 5'd13, 27'h00000022, 5'd27, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000293, 5'd22, 27'h00000231, 5'd7, 27'h000002f9, 32'h00000400,
  1'd1,  5'd13, 27'h0000011f, 5'd22, 27'h0000020c, 5'd18, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000037c, 5'd24, 27'h000001fd, 5'd30, 27'h00000218, 32'h00000400,
  1'd1,  5'd25, 27'h0000007b, 5'd2, 27'h00000327, 5'd10, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002b8, 5'd0, 27'h0000012e, 5'd17, 27'h00000002, 32'h00000400,
  1'd1,  5'd21, 27'h00000051, 5'd0, 27'h00000002, 5'd26, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000013a, 5'd11, 27'h00000180, 5'd6, 27'h000000c7, 32'h00000400,
  1'd1,  5'd25, 27'h00000094, 5'd13, 27'h00000365, 5'd19, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000028e, 5'd15, 27'h00000013, 5'd28, 27'h000003f1, 32'h00000400,
  1'd1,  5'd24, 27'h0000024e, 5'd25, 27'h000002ab, 5'd8, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000031f, 5'd24, 27'h00000350, 5'd17, 27'h000000d5, 32'h00000400,
  1'd1,  5'd21, 27'h0000038e, 5'd20, 27'h000003df, 5'd29, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000083, 5'd6, 27'h00000280, 5'd3, 27'h000001c8, 32'h00000400,
  1'd1,  5'd3, 27'h00000165, 5'd7, 27'h0000025b, 5'd11, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000178, 5'd5, 27'h000002b1, 5'd24, 27'h00000167, 32'h00000400,
  1'd1,  5'd2, 27'h000000a6, 5'd16, 27'h00000168, 5'd5, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003c1, 5'd18, 27'h000002f2, 5'd12, 27'h00000256, 32'h00000400,
  1'd1,  5'd4, 27'h00000256, 5'd19, 27'h00000087, 5'd20, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000208, 5'd29, 27'h000001d9, 5'd2, 27'h00000245, 32'h00000400,
  1'd1,  5'd0, 27'h000002f5, 5'd27, 27'h00000252, 5'd14, 27'h0000031b, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000261, 5'd30, 27'h0000036c, 5'd22, 27'h00000117, 32'h00000400,
  1'd1,  5'd13, 27'h00000267, 5'd6, 27'h000000a1, 5'd0, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d2, 5'd9, 27'h000003fa, 5'd12, 27'h000003b3, 32'h00000400,
  1'd1,  5'd11, 27'h000003f5, 5'd6, 27'h000003ea, 5'd25, 27'h0000020a, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f1, 5'd15, 27'h000003ec, 5'd4, 27'h000002a7, 32'h00000400,
  1'd1,  5'd13, 27'h00000208, 5'd19, 27'h000000e7, 5'd10, 27'h00000304, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001c6, 5'd18, 27'h000002b3, 5'd24, 27'h00000163, 32'h00000400,
  1'd1,  5'd13, 27'h0000008a, 5'd29, 27'h000002de, 5'd3, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000135, 5'd26, 27'h000001c8, 5'd12, 27'h000002e4, 32'h00000400,
  1'd1,  5'd10, 27'h0000015d, 5'd26, 27'h00000333, 5'd24, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000c4, 5'd9, 27'h0000028d, 5'd2, 27'h000003b6, 32'h00000400,
  1'd1,  5'd22, 27'h000001d7, 5'd6, 27'h000001aa, 5'd12, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001c6, 5'd16, 27'h0000018b, 5'd3, 27'h0000038d, 32'h00000400,
  1'd1,  5'd22, 27'h00000231, 5'd20, 27'h00000253, 5'd10, 27'h0000022a, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f8, 5'd16, 27'h000002c3, 5'd24, 27'h000001bf, 32'h00000400,
  1'd1,  5'd22, 27'h0000006f, 5'd26, 27'h00000293, 5'd3, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000283, 5'd28, 27'h000000aa, 5'd10, 27'h0000029e, 32'h00000400,
  1'd1,  5'd23, 27'h00000289, 5'd29, 27'h0000026b, 5'd22, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000113, 5'd8, 27'h000001c1, 5'd7, 27'h0000013a, 32'h00000400,
  1'd1,  5'd2, 27'h00000153, 5'd7, 27'h0000039f, 5'd17, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000034c, 5'd6, 27'h0000008e, 5'd26, 27'h00000250, 32'h00000400,
  1'd1,  5'd4, 27'h00000250, 5'd16, 27'h00000170, 5'd6, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000010f, 5'd18, 27'h00000303, 5'd17, 27'h00000323, 32'h00000400,
  1'd1,  5'd0, 27'h000001f9, 5'd19, 27'h00000028, 5'd28, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000d5, 5'd29, 27'h000001a9, 5'd7, 27'h00000179, 32'h00000400,
  1'd1,  5'd2, 27'h00000366, 5'd28, 27'h0000015b, 5'd15, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000229, 5'd27, 27'h0000021e, 5'd29, 27'h000003f7, 32'h00000400,
  1'd1,  5'd15, 27'h0000002e, 5'd6, 27'h000002b9, 5'd5, 27'h0000034d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000347, 5'd8, 27'h0000029b, 5'd19, 27'h00000103, 32'h00000400,
  1'd1,  5'd11, 27'h000001de, 5'd5, 27'h0000025e, 5'd29, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001fd, 5'd17, 27'h000003f1, 5'd8, 27'h000000be, 32'h00000400,
  1'd1,  5'd13, 27'h00000006, 5'd18, 27'h0000035b, 5'd20, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f5, 5'd20, 27'h00000240, 5'd28, 27'h00000158, 32'h00000400,
  1'd1,  5'd15, 27'h0000018b, 5'd28, 27'h000002df, 5'd8, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000037d, 5'd28, 27'h000000db, 5'd16, 27'h000002bb, 32'h00000400,
  1'd1,  5'd13, 27'h000002ff, 5'd27, 27'h000002b3, 5'd29, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000354, 5'd5, 27'h00000274, 5'd7, 27'h0000004a, 32'h00000400,
  1'd1,  5'd24, 27'h000003ce, 5'd7, 27'h0000008a, 5'd20, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000302, 5'd5, 27'h0000028e, 5'd29, 27'h000002de, 32'h00000400,
  1'd1,  5'd24, 27'h000000ee, 5'd18, 27'h00000273, 5'd9, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000001e, 5'd20, 27'h00000077, 5'd19, 27'h0000037b, 32'h00000400,
  1'd1,  5'd20, 27'h0000033a, 5'd16, 27'h00000236, 5'd29, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000382, 5'd29, 27'h0000020f, 5'd5, 27'h000003aa, 32'h00000400,
  1'd1,  5'd24, 27'h000000a5, 5'd27, 27'h000002b4, 5'd15, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000005e, 5'd26, 27'h00000074, 5'd26, 27'h0000010b, 32'h00000400,
  1'd1,  5'd5, 27'h00000195, 5'd3, 27'h00000293, 5'd5, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000328, 5'd0, 27'h00000016, 5'd17, 27'h00000175, 32'h00000400,
  1'd1,  5'd6, 27'h000000f4, 5'd5, 27'h00000032, 5'd27, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032a, 5'd14, 27'h00000240, 5'd3, 27'h000000ed, 32'h00000400,
  1'd1,  5'd8, 27'h000001f3, 5'd12, 27'h00000276, 5'd13, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000013a, 5'd13, 27'h000000d5, 5'd25, 27'h00000141, 32'h00000400,
  1'd1,  5'd5, 27'h00000243, 5'd25, 27'h000001ce, 5'd1, 27'h00000345, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003f2, 5'd25, 27'h0000011d, 5'd14, 27'h000001a8, 32'h00000400,
  1'd1,  5'd8, 27'h000001cc, 5'd24, 27'h000002a7, 5'd20, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000012d, 5'd1, 27'h000003cb, 5'd6, 27'h0000015b, 32'h00000400,
  1'd1,  5'd18, 27'h00000030, 5'd1, 27'h0000016f, 5'd17, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000040, 5'd0, 27'h000001d8, 5'd26, 27'h000000f7, 32'h00000400,
  1'd1,  5'd17, 27'h000001cf, 5'd14, 27'h0000004a, 5'd1, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000020f, 5'd14, 27'h00000373, 5'd12, 27'h00000142, 32'h00000400,
  1'd1,  5'd19, 27'h00000279, 5'd10, 27'h00000168, 5'd23, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000218, 5'd23, 27'h0000033a, 5'd3, 27'h000000af, 32'h00000400,
  1'd1,  5'd18, 27'h000001cf, 5'd20, 27'h00000392, 5'd14, 27'h00000140, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000b0, 5'd23, 27'h00000227, 5'd20, 27'h000003db, 32'h00000400,
  1'd1,  5'd27, 27'h0000038b, 5'd4, 27'h000002ea, 5'd0, 27'h0000020b, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003a8, 5'd2, 27'h0000024b, 5'd11, 27'h00000213, 32'h00000400,
  1'd1,  5'd28, 27'h00000374, 5'd4, 27'h0000021c, 5'd23, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000315, 5'd14, 27'h00000022, 5'd3, 27'h00000377, 32'h00000400,
  1'd1,  5'd28, 27'h000000b0, 5'd13, 27'h0000025c, 5'd11, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000234, 5'd14, 27'h000001ab, 5'd21, 27'h00000027, 32'h00000400,
  1'd1,  5'd27, 27'h00000139, 5'd21, 27'h00000088, 5'd0, 27'h0000022f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000063, 5'd22, 27'h0000003a, 5'd12, 27'h0000037b, 32'h00000400,
  1'd1,  5'd29, 27'h0000008a, 5'd20, 27'h00000337, 5'd23, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000ce, 5'd0, 27'h000000de, 5'd0, 27'h00000029, 32'h00000400,
  1'd1,  5'd9, 27'h0000006f, 5'd1, 27'h00000117, 5'd12, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000c2, 5'd1, 27'h00000258, 5'd24, 27'h00000210, 32'h00000400,
  1'd1,  5'd5, 27'h0000014f, 5'd13, 27'h00000011, 5'd7, 27'h00000338, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000027, 5'd14, 27'h0000029b, 5'd16, 27'h0000022e, 32'h00000400,
  1'd1,  5'd8, 27'h000003ee, 5'd13, 27'h000001b7, 5'd28, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000121, 5'd24, 27'h0000013b, 5'd8, 27'h00000325, 32'h00000400,
  1'd1,  5'd8, 27'h00000218, 5'd21, 27'h000002af, 5'd19, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000143, 5'd21, 27'h00000170, 5'd26, 27'h00000372, 32'h00000400,
  1'd1,  5'd20, 27'h00000209, 5'd1, 27'h00000371, 5'd2, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001ba, 5'd2, 27'h000001ae, 5'd15, 27'h00000098, 32'h00000400,
  1'd1,  5'd16, 27'h00000248, 5'd13, 27'h000003b1, 5'd6, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000036, 5'd11, 27'h000003c2, 5'd17, 27'h0000013a, 32'h00000400,
  1'd1,  5'd20, 27'h000000eb, 5'd13, 27'h000003a7, 5'd26, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000295, 5'd24, 27'h000000bc, 5'd9, 27'h00000199, 32'h00000400,
  1'd1,  5'd16, 27'h0000006b, 5'd23, 27'h00000183, 5'd17, 27'h00000237, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000002b, 5'd23, 27'h00000135, 5'd30, 27'h00000223, 32'h00000400,
  1'd1,  5'd28, 27'h000003a8, 5'd0, 27'h000000e8, 5'd9, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003f2, 5'd4, 27'h000002ac, 5'd19, 27'h0000005d, 32'h00000400,
  1'd1,  5'd29, 27'h00000274, 5'd3, 27'h000002c7, 5'd26, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000005a, 5'd15, 27'h00000087, 5'd8, 27'h0000035b, 32'h00000400,
  1'd1,  5'd26, 27'h000002da, 5'd15, 27'h0000003d, 5'd15, 27'h000002e6, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003c1, 5'd14, 27'h000001f2, 5'd26, 27'h000001cf, 32'h00000400,
  1'd1,  5'd27, 27'h000003e6, 5'd20, 27'h000003f6, 5'd5, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000278, 5'd21, 27'h00000002, 5'd18, 27'h00000328, 32'h00000400,
  1'd1,  5'd28, 27'h000003bc, 5'd24, 27'h00000294, 5'd30, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000101, 5'd6, 27'h00000033, 5'd1, 27'h000000bf, 32'h00000400,
  1'd1,  5'd8, 27'h000000a5, 5'd7, 27'h000001cc, 5'd13, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000007f, 5'd8, 27'h000000e0, 5'd21, 27'h00000214, 32'h00000400,
  1'd1,  5'd8, 27'h00000204, 5'd17, 27'h0000022a, 5'd3, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001ba, 5'd15, 27'h000003f2, 5'd14, 27'h00000115, 32'h00000400,
  1'd1,  5'd10, 27'h00000114, 5'd16, 27'h00000121, 5'd24, 27'h00000151, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000090, 5'd30, 27'h0000016a, 5'd2, 27'h0000001e, 32'h00000400,
  1'd1,  5'd7, 27'h00000173, 5'd27, 27'h0000038b, 5'd10, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000350, 5'd30, 27'h0000011a, 5'd20, 27'h0000031b, 32'h00000400,
  1'd1,  5'd17, 27'h0000039e, 5'd5, 27'h00000363, 5'd1, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001cd, 5'd8, 27'h0000037c, 5'd14, 27'h000003ab, 32'h00000400,
  1'd1,  5'd17, 27'h000002e0, 5'd9, 27'h000000cd, 5'd21, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a9, 5'd15, 27'h000003a2, 5'd0, 27'h00000003, 32'h00000400,
  1'd1,  5'd16, 27'h00000366, 5'd19, 27'h000001e3, 5'd12, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000d8, 5'd15, 27'h00000228, 5'd24, 27'h000001de, 32'h00000400,
  1'd1,  5'd20, 27'h00000100, 5'd30, 27'h0000017f, 5'd2, 27'h000003a7, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000025f, 5'd27, 27'h00000071, 5'd11, 27'h00000105, 32'h00000400,
  1'd1,  5'd20, 27'h000001d9, 5'd28, 27'h000001f3, 5'd21, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000018a, 5'd8, 27'h00000150, 5'd0, 27'h0000031c, 32'h00000400,
  1'd1,  5'd28, 27'h000003ca, 5'd5, 27'h00000288, 5'd15, 27'h0000018f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000037e, 5'd6, 27'h00000172, 5'd21, 27'h00000056, 32'h00000400,
  1'd1,  5'd28, 27'h00000230, 5'd18, 27'h00000062, 5'd0, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000334, 5'd19, 27'h00000243, 5'd11, 27'h0000000a, 32'h00000400,
  1'd1,  5'd27, 27'h0000003f, 5'd18, 27'h00000115, 5'd23, 27'h0000038d, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000031a, 5'd28, 27'h00000072, 5'd4, 27'h000002c9, 32'h00000400,
  1'd1,  5'd28, 27'h00000338, 5'd26, 27'h0000018b, 5'd14, 27'h000002bf, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003d8, 5'd26, 27'h000000ec, 5'd23, 27'h000002fd, 32'h00000400,
  1'd1,  5'd6, 27'h00000179, 5'd7, 27'h0000014c, 5'd5, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000190, 5'd10, 27'h0000012b, 5'd15, 27'h0000021e, 32'h00000400,
  1'd1,  5'd9, 27'h00000365, 5'd6, 27'h0000030a, 5'd27, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000022, 5'd19, 27'h00000168, 5'd5, 27'h000002b9, 32'h00000400,
  1'd1,  5'd9, 27'h000000ac, 5'd19, 27'h00000161, 5'd19, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003fd, 5'd19, 27'h00000084, 5'd28, 27'h00000166, 32'h00000400,
  1'd1,  5'd8, 27'h00000377, 5'd30, 27'h00000097, 5'd5, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000100, 5'd29, 27'h000002bb, 5'd18, 27'h00000348, 32'h00000400,
  1'd1,  5'd9, 27'h00000253, 5'd26, 27'h000001c3, 5'd30, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002a7, 5'd9, 27'h0000029f, 5'd8, 27'h0000023a, 32'h00000400,
  1'd1,  5'd20, 27'h00000170, 5'd6, 27'h0000009d, 5'd18, 27'h000002a2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000173, 5'd8, 27'h00000371, 5'd27, 27'h00000036, 32'h00000400,
  1'd1,  5'd19, 27'h000001cb, 5'd16, 27'h000001bd, 5'd6, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001fc, 5'd19, 27'h00000369, 5'd17, 27'h00000085, 32'h00000400,
  1'd1,  5'd20, 27'h00000130, 5'd18, 27'h00000209, 5'd26, 27'h0000029e, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000339, 5'd27, 27'h00000395, 5'd9, 27'h000003dd, 32'h00000400,
  1'd1,  5'd16, 27'h00000008, 5'd29, 27'h00000196, 5'd19, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000e0, 5'd28, 27'h0000030a, 5'd28, 27'h000003fb, 32'h00000400,
  1'd1,  5'd29, 27'h00000178, 5'd5, 27'h0000031c, 5'd8, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000029a, 5'd5, 27'h0000022d, 5'd17, 27'h000000ac, 32'h00000400,
  1'd1,  5'd27, 27'h000002d0, 5'd8, 27'h00000181, 5'd29, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000016e, 5'd20, 27'h0000021f, 5'd6, 27'h00000153, 32'h00000400,
  1'd1,  5'd27, 27'h00000180, 5'd18, 27'h0000030a, 5'd15, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000025, 5'd17, 27'h0000010e, 5'd26, 27'h0000006f, 32'h00000400,
  1'd1,  5'd26, 27'h000003c1, 5'd28, 27'h00000074, 5'd7, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000008a, 5'd29, 27'h0000021c, 5'd15, 27'h000003d4, 32'h00000400,
  1'd1,  5'd29, 27'h0000018a, 5'd26, 27'h000003d1, 5'd30, 27'h00000374, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000002ed, 5'd1, 27'h000001d9, 5'd1, 27'h000002a8, 32'h00000400,
  1'd1,  5'd5, 27'h00000076, 5'd4, 27'h00000319, 5'd11, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001cb, 5'd0, 27'h000000da, 5'd20, 27'h000003b5, 32'h00000400,
  1'd1,  5'd1, 27'h00000131, 5'd13, 27'h00000115, 5'd5, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000039d, 5'd11, 27'h000003b7, 5'd15, 27'h00000069, 32'h00000400,
  1'd1,  5'd1, 27'h00000198, 5'd12, 27'h00000198, 5'd24, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ee, 5'd21, 27'h00000262, 5'd3, 27'h000003f6, 32'h00000400,
  1'd1,  5'd3, 27'h0000033c, 5'd25, 27'h000001c8, 5'd11, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000014b, 5'd20, 27'h00000387, 5'd25, 27'h000002fa, 32'h00000400,
  1'd1,  5'd13, 27'h00000254, 5'd5, 27'h0000004b, 5'd1, 27'h000000fe, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000298, 5'd2, 27'h00000104, 5'd11, 27'h00000328, 32'h00000400,
  1'd1,  5'd11, 27'h00000211, 5'd0, 27'h00000307, 5'd24, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000007c, 5'd12, 27'h00000168, 5'd0, 27'h00000104, 32'h00000400,
  1'd1,  5'd13, 27'h000000ca, 5'd15, 27'h00000148, 5'd14, 27'h000000a6, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002df, 5'd11, 27'h000002ee, 5'd23, 27'h00000031, 32'h00000400,
  1'd1,  5'd13, 27'h000000f8, 5'd25, 27'h0000021f, 5'd3, 27'h000000c8, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000ab, 5'd23, 27'h000001e3, 5'd10, 27'h000002f9, 32'h00000400,
  1'd1,  5'd11, 27'h00000254, 5'd24, 27'h000001bb, 5'd24, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000227, 5'd1, 27'h00000129, 5'd2, 27'h00000390, 32'h00000400,
  1'd1,  5'd22, 27'h000001ec, 5'd2, 27'h000003a2, 5'd14, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e2, 5'd4, 27'h00000259, 5'd25, 27'h0000028e, 32'h00000400,
  1'd1,  5'd22, 27'h0000010f, 5'd11, 27'h00000160, 5'd5, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e5, 5'd11, 27'h000000ea, 5'd12, 27'h0000031f, 32'h00000400,
  1'd1,  5'd25, 27'h000001c0, 5'd14, 27'h000003ae, 5'd21, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000391, 5'd22, 27'h00000014, 5'd2, 27'h000000ce, 32'h00000400,
  1'd1,  5'd22, 27'h000000dc, 5'd21, 27'h000001e4, 5'd10, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000a8, 5'd23, 27'h000003e4, 5'd21, 27'h000001ff, 32'h00000400,
  1'd1,  5'd1, 27'h00000381, 5'd3, 27'h0000013d, 5'd8, 27'h000001af, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b1, 5'd2, 27'h000000ae, 5'd19, 27'h000000a6, 32'h00000400,
  1'd1,  5'd3, 27'h00000263, 5'd0, 27'h000003e4, 5'd27, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003f2, 5'd14, 27'h000002a5, 5'd8, 27'h00000127, 32'h00000400,
  1'd1,  5'd4, 27'h0000000d, 5'd14, 27'h00000164, 5'd19, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001f7, 5'd11, 27'h000003da, 5'd25, 27'h000003a1, 32'h00000400,
  1'd1,  5'd4, 27'h0000038c, 5'd22, 27'h000002c9, 5'd9, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000189, 5'd25, 27'h000002a8, 5'd19, 27'h00000374, 32'h00000400,
  1'd1,  5'd5, 27'h0000007e, 5'd23, 27'h0000027b, 5'd26, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000087, 5'd5, 27'h00000076, 5'd8, 27'h000003c0, 32'h00000400,
  1'd1,  5'd14, 27'h0000021a, 5'd1, 27'h00000308, 5'd16, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001e6, 5'd4, 27'h00000286, 5'd27, 27'h000001e1, 32'h00000400,
  1'd1,  5'd11, 27'h000002ec, 5'd14, 27'h0000022b, 5'd6, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003ad, 5'd11, 27'h00000173, 5'd20, 27'h0000010b, 32'h00000400,
  1'd1,  5'd14, 27'h000000cd, 5'd12, 27'h000000bf, 5'd27, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000b3, 5'd22, 27'h0000007f, 5'd9, 27'h0000010f, 32'h00000400,
  1'd1,  5'd11, 27'h000002f1, 5'd25, 27'h000001d9, 5'd19, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d2, 5'd20, 27'h0000039c, 5'd29, 27'h000000e7, 32'h00000400,
  1'd1,  5'd21, 27'h000002fc, 5'd0, 27'h0000024b, 5'd8, 27'h000003e7, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001f2, 5'd1, 27'h00000158, 5'd17, 27'h00000161, 32'h00000400,
  1'd1,  5'd24, 27'h000001f0, 5'd3, 27'h000001c6, 5'd28, 27'h00000088, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000327, 5'd13, 27'h00000256, 5'd7, 27'h00000248, 32'h00000400,
  1'd1,  5'd22, 27'h00000100, 5'd10, 27'h0000031b, 5'd18, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000c7, 5'd15, 27'h00000110, 5'd29, 27'h0000015e, 32'h00000400,
  1'd1,  5'd22, 27'h000001af, 5'd25, 27'h00000081, 5'd5, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000175, 5'd22, 27'h000003e7, 5'd17, 27'h0000034d, 32'h00000400,
  1'd1,  5'd22, 27'h00000199, 5'd23, 27'h000001c2, 5'd30, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000008c, 5'd7, 27'h00000333, 5'd2, 27'h00000170, 32'h00000400,
  1'd1,  5'd2, 27'h0000034a, 5'd5, 27'h000003f5, 5'd11, 27'h0000001f, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000377, 5'd8, 27'h0000021a, 5'd21, 27'h000000b3, 32'h00000400,
  1'd1,  5'd0, 27'h000003b8, 5'd17, 27'h000002fc, 5'd0, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003ab, 5'd16, 27'h00000033, 5'd12, 27'h0000019b, 32'h00000400,
  1'd1,  5'd0, 27'h0000023a, 5'd18, 27'h0000038b, 5'd24, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000007b, 5'd27, 27'h00000138, 5'd2, 27'h0000037f, 32'h00000400,
  1'd1,  5'd0, 27'h0000011a, 5'd26, 27'h000002a3, 5'd13, 27'h0000023d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000258, 5'd25, 27'h00000376, 5'd22, 27'h000001ed, 32'h00000400,
  1'd1,  5'd13, 27'h000001cd, 5'd8, 27'h00000155, 5'd4, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000071, 5'd9, 27'h000000d7, 5'd14, 27'h0000003a, 32'h00000400,
  1'd1,  5'd10, 27'h000001e9, 5'd9, 27'h0000014d, 5'd22, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001b1, 5'd19, 27'h00000379, 5'd3, 27'h000003d8, 32'h00000400,
  1'd1,  5'd13, 27'h0000015c, 5'd16, 27'h00000220, 5'd13, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002cd, 5'd17, 27'h00000237, 5'd24, 27'h000001f1, 32'h00000400,
  1'd1,  5'd13, 27'h0000029e, 5'd27, 27'h000002cc, 5'd5, 27'h00000013, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003ec, 5'd28, 27'h00000036, 5'd14, 27'h0000013b, 32'h00000400,
  1'd1,  5'd14, 27'h00000205, 5'd26, 27'h000001dd, 5'd21, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d0, 5'd5, 27'h0000034e, 5'd2, 27'h000003bb, 32'h00000400,
  1'd1,  5'd22, 27'h00000096, 5'd5, 27'h000003b1, 5'd11, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000380, 5'd19, 27'h000002c3, 5'd4, 27'h000001df, 32'h00000400,
  1'd1,  5'd21, 27'h000002ad, 5'd16, 27'h00000379, 5'd12, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000015f, 5'd16, 27'h000002a8, 5'd25, 27'h0000023f, 32'h00000400,
  1'd1,  5'd24, 27'h00000244, 5'd29, 27'h0000011f, 5'd0, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003d1, 5'd27, 27'h000000cd, 5'd12, 27'h00000207, 32'h00000400,
  1'd1,  5'd25, 27'h000001cd, 5'd28, 27'h00000155, 5'd20, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000346, 5'd9, 27'h000003eb, 5'd8, 27'h0000039d, 32'h00000400,
  1'd1,  5'd2, 27'h00000189, 5'd6, 27'h000002f5, 5'd19, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000102, 5'd10, 27'h00000079, 5'd30, 27'h0000032f, 32'h00000400,
  1'd1,  5'd3, 27'h000003b7, 5'd16, 27'h00000124, 5'd6, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000078, 5'd18, 27'h000000d0, 5'd15, 27'h000002c7, 32'h00000400,
  1'd1,  5'd0, 27'h0000001a, 5'd18, 27'h00000157, 5'd29, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003d0, 5'd29, 27'h0000026f, 5'd7, 27'h0000003a, 32'h00000400,
  1'd1,  5'd3, 27'h00000141, 5'd28, 27'h00000398, 5'd17, 27'h0000039f, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000fc, 5'd26, 27'h00000162, 5'd29, 27'h0000035b, 32'h00000400,
  1'd1,  5'd10, 27'h0000032e, 5'd6, 27'h0000011f, 5'd7, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000341, 5'd7, 27'h000000b5, 5'd19, 27'h00000215, 32'h00000400,
  1'd1,  5'd12, 27'h0000010e, 5'd6, 27'h000003a3, 5'd29, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002f7, 5'd18, 27'h00000350, 5'd9, 27'h000002d4, 32'h00000400,
  1'd1,  5'd14, 27'h00000223, 5'd18, 27'h00000350, 5'd18, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a6, 5'd15, 27'h00000379, 5'd27, 27'h0000017a, 32'h00000400,
  1'd1,  5'd15, 27'h0000011e, 5'd28, 27'h0000007a, 5'd9, 27'h000000a0, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002a7, 5'd28, 27'h00000101, 5'd17, 27'h000003a5, 32'h00000400,
  1'd1,  5'd14, 27'h00000155, 5'd29, 27'h000001e4, 5'd27, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000050, 5'd9, 27'h000001a4, 5'd5, 27'h00000142, 32'h00000400,
  1'd1,  5'd21, 27'h000000cc, 5'd7, 27'h0000001e, 5'd18, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000285, 5'd6, 27'h0000029f, 5'd28, 27'h000000fd, 32'h00000400,
  1'd1,  5'd25, 27'h0000028c, 5'd17, 27'h00000262, 5'd10, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000046, 5'd15, 27'h000002c2, 5'd18, 27'h000001d1, 32'h00000400,
  1'd1,  5'd22, 27'h00000135, 5'd18, 27'h00000044, 5'd26, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000012c, 5'd29, 27'h00000338, 5'd9, 27'h0000017d, 32'h00000400,
  1'd1,  5'd23, 27'h000003e4, 5'd29, 27'h000003e6, 5'd18, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000210, 5'd27, 27'h000003d9, 5'd27, 27'h000001e9, 32'h00000400,
  1'd1,  5'd9, 27'h000000c6, 5'd1, 27'h000000e6, 5'd8, 27'h00000123, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000c7, 5'd1, 27'h000001c6, 5'd19, 27'h000002c7, 32'h00000400,
  1'd1,  5'd10, 27'h000000e5, 5'd2, 27'h00000279, 5'd30, 27'h000002d3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000cf, 5'd11, 27'h000002c5, 5'd0, 27'h00000195, 32'h00000400,
  1'd1,  5'd6, 27'h000002e3, 5'd15, 27'h0000009c, 5'd13, 27'h0000026f, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000370, 5'd11, 27'h000003d9, 5'd24, 27'h00000232, 32'h00000400,
  1'd1,  5'd7, 27'h00000029, 5'd25, 27'h000001c2, 5'd3, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000014d, 5'd23, 27'h000002d2, 5'd15, 27'h0000014d, 32'h00000400,
  1'd1,  5'd9, 27'h00000329, 5'd25, 27'h000000e3, 5'd21, 27'h000003ac, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000176, 5'd1, 27'h00000136, 5'd9, 27'h00000148, 32'h00000400,
  1'd1,  5'd17, 27'h00000381, 5'd2, 27'h000001d0, 5'd18, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000180, 5'd3, 27'h00000299, 5'd26, 27'h000001a5, 32'h00000400,
  1'd1,  5'd17, 27'h000000c1, 5'd12, 27'h000003b8, 5'd4, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000014c, 5'd11, 27'h000001ac, 5'd14, 27'h00000302, 32'h00000400,
  1'd1,  5'd18, 27'h00000142, 5'd15, 27'h0000013b, 5'd25, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002c3, 5'd22, 27'h00000038, 5'd0, 27'h000003a6, 32'h00000400,
  1'd1,  5'd16, 27'h000002d4, 5'd24, 27'h000003ef, 5'd11, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000309, 5'd21, 27'h00000310, 5'd23, 27'h0000015e, 32'h00000400,
  1'd1,  5'd29, 27'h00000191, 5'd2, 27'h000003ee, 5'd1, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a7, 5'd3, 27'h000001a9, 5'd15, 27'h00000030, 32'h00000400,
  1'd1,  5'd26, 27'h0000017e, 5'd0, 27'h0000008e, 5'd22, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000001c, 5'd11, 27'h000002b2, 5'd4, 27'h00000225, 32'h00000400,
  1'd1,  5'd30, 27'h0000009d, 5'd13, 27'h0000006c, 5'd11, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000106, 5'd13, 27'h00000066, 5'd24, 27'h00000196, 32'h00000400,
  1'd1,  5'd26, 27'h00000281, 5'd23, 27'h0000022e, 5'd1, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000277, 5'd22, 27'h00000026, 5'd15, 27'h00000119, 32'h00000400,
  1'd1,  5'd28, 27'h00000137, 5'd20, 27'h00000386, 5'd25, 27'h000002d1, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003bb, 5'd4, 27'h000001b0, 5'd0, 27'h00000287, 32'h00000400,
  1'd1,  5'd9, 27'h0000012a, 5'd4, 27'h000000f1, 5'd13, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000076, 5'd4, 27'h0000021c, 5'd23, 27'h0000022c, 32'h00000400,
  1'd1,  5'd10, 27'h0000009b, 5'd10, 27'h0000022f, 5'd6, 27'h000001a9, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000137, 5'd10, 27'h000001c4, 5'd16, 27'h000000eb, 32'h00000400,
  1'd1,  5'd9, 27'h000000de, 5'd10, 27'h000002fd, 5'd29, 27'h00000200, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003bd, 5'd22, 27'h00000240, 5'd7, 27'h00000282, 32'h00000400,
  1'd1,  5'd7, 27'h00000112, 5'd21, 27'h0000018c, 5'd19, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a6, 5'd23, 27'h0000033b, 5'd27, 27'h000002f0, 32'h00000400,
  1'd1,  5'd15, 27'h00000361, 5'd5, 27'h00000087, 5'd1, 27'h00000159, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000008a, 5'd3, 27'h000001b2, 5'd12, 27'h000003ca, 32'h00000400,
  1'd1,  5'd17, 27'h00000162, 5'd15, 27'h00000122, 5'd5, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001f5, 5'd13, 27'h00000028, 5'd20, 27'h00000088, 32'h00000400,
  1'd1,  5'd20, 27'h000001fd, 5'd12, 27'h0000035d, 5'd26, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000351, 5'd22, 27'h000001bb, 5'd6, 27'h00000173, 32'h00000400,
  1'd1,  5'd19, 27'h000002fe, 5'd25, 27'h000001ed, 5'd16, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000026d, 5'd22, 27'h000003f5, 5'd27, 27'h00000320, 32'h00000400,
  1'd1,  5'd25, 27'h000003f3, 5'd0, 27'h0000012a, 5'd5, 27'h0000034c, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000014d, 5'd2, 27'h00000330, 5'd18, 27'h00000255, 32'h00000400,
  1'd1,  5'd26, 27'h0000000a, 5'd1, 27'h00000024, 5'd27, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000339, 5'd11, 27'h000002e9, 5'd7, 27'h000003b6, 32'h00000400,
  1'd1,  5'd29, 27'h000003df, 5'd14, 27'h0000005f, 5'd16, 27'h000000b4, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000367, 5'd13, 27'h0000036c, 5'd28, 27'h0000035e, 32'h00000400,
  1'd1,  5'd29, 27'h0000002c, 5'd24, 27'h00000234, 5'd8, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003af, 5'd24, 27'h00000241, 5'd18, 27'h0000032c, 32'h00000400,
  1'd1,  5'd30, 27'h0000005b, 5'd21, 27'h000001e5, 5'd28, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000140, 5'd9, 27'h0000030f, 5'd4, 27'h00000249, 32'h00000400,
  1'd1,  5'd6, 27'h000002bc, 5'd8, 27'h00000185, 5'd11, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001af, 5'd7, 27'h000000c5, 5'd22, 27'h00000147, 32'h00000400,
  1'd1,  5'd10, 27'h00000069, 5'd17, 27'h000002cd, 5'd3, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000148, 5'd18, 27'h000001c1, 5'd11, 27'h00000328, 32'h00000400,
  1'd1,  5'd9, 27'h00000263, 5'd18, 27'h000001ae, 5'd24, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000391, 5'd30, 27'h00000030, 5'd2, 27'h00000391, 32'h00000400,
  1'd1,  5'd8, 27'h0000003e, 5'd26, 27'h00000293, 5'd10, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ef, 5'd28, 27'h00000391, 5'd23, 27'h000003dd, 32'h00000400,
  1'd1,  5'd19, 27'h000003f9, 5'd8, 27'h00000291, 5'd4, 27'h000003c5, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000139, 5'd8, 27'h0000028a, 5'd14, 27'h0000039b, 32'h00000400,
  1'd1,  5'd19, 27'h0000035c, 5'd9, 27'h0000009b, 5'd23, 27'h000001a3, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000037, 5'd18, 27'h000000f3, 5'd3, 27'h00000091, 32'h00000400,
  1'd1,  5'd16, 27'h00000308, 5'd15, 27'h00000212, 5'd14, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000386, 5'd16, 27'h000003ea, 5'd20, 27'h000002f8, 32'h00000400,
  1'd1,  5'd16, 27'h000003a0, 5'd25, 27'h000003f7, 5'd4, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001a4, 5'd26, 27'h00000081, 5'd13, 27'h000001bc, 32'h00000400,
  1'd1,  5'd18, 27'h00000380, 5'd30, 27'h00000058, 5'd22, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002c7, 5'd8, 27'h00000067, 5'd3, 27'h00000295, 32'h00000400,
  1'd1,  5'd29, 27'h00000279, 5'd7, 27'h000002ff, 5'd13, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002fa, 5'd7, 27'h000001b9, 5'd21, 27'h00000311, 32'h00000400,
  1'd1,  5'd28, 27'h0000035b, 5'd16, 27'h000001be, 5'd4, 27'h0000019c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002dd, 5'd16, 27'h0000026f, 5'd10, 27'h00000400, 32'h00000400,
  1'd1,  5'd27, 27'h00000376, 5'd16, 27'h0000039c, 5'd20, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000d6, 5'd29, 27'h00000058, 5'd2, 27'h000001ee, 32'h00000400,
  1'd1,  5'd27, 27'h00000344, 5'd28, 27'h00000137, 5'd13, 27'h000000f2, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003b9, 5'd28, 27'h00000179, 5'd23, 27'h00000255, 32'h00000400,
  1'd1,  5'd9, 27'h000000ce, 5'd9, 27'h0000003a, 5'd9, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000398, 5'd7, 27'h000002d9, 5'd17, 27'h00000297, 32'h00000400,
  1'd1,  5'd8, 27'h000000f3, 5'd8, 27'h0000016d, 5'd29, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000093, 5'd18, 27'h000002c2, 5'd5, 27'h000003f3, 32'h00000400,
  1'd1,  5'd7, 27'h0000029a, 5'd15, 27'h00000321, 5'd16, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a6, 5'd20, 27'h00000209, 5'd29, 27'h000000b1, 32'h00000400,
  1'd1,  5'd9, 27'h00000103, 5'd28, 27'h0000029f, 5'd8, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000101, 5'd28, 27'h0000025a, 5'd20, 27'h00000083, 32'h00000400,
  1'd1,  5'd5, 27'h0000026e, 5'd29, 27'h00000237, 5'd27, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000019f, 5'd6, 27'h000001f6, 5'd5, 27'h0000027a, 32'h00000400,
  1'd1,  5'd18, 27'h000000d2, 5'd5, 27'h000001bd, 5'd17, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001f, 5'd8, 27'h000002ee, 5'd28, 27'h00000036, 32'h00000400,
  1'd1,  5'd18, 27'h000003d9, 5'd17, 27'h000002e6, 5'd9, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003a1, 5'd17, 27'h00000275, 5'd15, 27'h00000294, 32'h00000400,
  1'd1,  5'd16, 27'h000002ef, 5'd20, 27'h0000005a, 5'd30, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000005b, 5'd27, 27'h00000167, 5'd5, 27'h000001f3, 32'h00000400,
  1'd1,  5'd19, 27'h000003b2, 5'd26, 27'h00000222, 5'd16, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002e9, 5'd28, 27'h00000001, 5'd29, 27'h00000115, 32'h00000400,
  1'd1,  5'd27, 27'h00000012, 5'd6, 27'h000000b1, 5'd8, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000048, 5'd6, 27'h0000038c, 5'd16, 27'h00000332, 32'h00000400,
  1'd1,  5'd29, 27'h0000038f, 5'd6, 27'h000001e4, 5'd27, 27'h00000319, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000368, 5'd19, 27'h000002ac, 5'd5, 27'h00000235, 32'h00000400,
  1'd1,  5'd29, 27'h00000139, 5'd20, 27'h0000015b, 5'd17, 27'h000000c0, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000cb, 5'd16, 27'h000000c5, 5'd30, 27'h00000100, 32'h00000400,
  1'd1,  5'd28, 27'h0000008d, 5'd29, 27'h000001f1, 5'd8, 27'h000001e3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000393, 5'd26, 27'h00000245, 5'd19, 27'h00000219, 32'h00000400,
  1'd1,  5'd30, 27'h000002c1, 5'd29, 27'h000002f4, 5'd29, 27'h000001b7, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h00000224, 5'd4, 27'h000003a6, 5'd2, 27'h000000d3, 32'h00000400,
  1'd1,  5'd2, 27'h00000340, 5'd2, 27'h00000150, 5'd14, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000ef, 5'd0, 27'h00000309, 5'd24, 27'h000002a1, 32'h00000400,
  1'd1,  5'd0, 27'h000003ca, 5'd14, 27'h0000018c, 5'd2, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000305, 5'd11, 27'h0000008d, 5'd12, 27'h000000de, 32'h00000400,
  1'd1,  5'd1, 27'h000002e7, 5'd12, 27'h000002e9, 5'd23, 27'h00000363, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003e8, 5'd21, 27'h00000208, 5'd3, 27'h00000023, 32'h00000400,
  1'd1,  5'd0, 27'h0000003d, 5'd24, 27'h000001d2, 5'd14, 27'h00000019, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000f6, 5'd23, 27'h0000001d, 5'd24, 27'h000001d7, 32'h00000400,
  1'd1,  5'd14, 27'h000003de, 5'd4, 27'h0000018f, 5'd0, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000aa, 5'd2, 27'h0000001a, 5'd15, 27'h00000094, 32'h00000400,
  1'd1,  5'd12, 27'h00000377, 5'd1, 27'h0000000b, 5'd25, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001ee, 5'd14, 27'h00000122, 5'd2, 27'h0000013e, 32'h00000400,
  1'd1,  5'd13, 27'h0000026a, 5'd12, 27'h0000024e, 5'd11, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000018e, 5'd13, 27'h0000020e, 5'd22, 27'h000002f0, 32'h00000400,
  1'd1,  5'd14, 27'h000003cb, 5'd20, 27'h00000362, 5'd2, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000377, 5'd24, 27'h000001c0, 5'd11, 27'h00000239, 32'h00000400,
  1'd1,  5'd15, 27'h000001bf, 5'd25, 27'h0000008a, 5'd24, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000038e, 5'd2, 27'h000000b8, 5'd4, 27'h0000007d, 32'h00000400,
  1'd1,  5'd25, 27'h0000019c, 5'd1, 27'h000002de, 5'd10, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ce, 5'd0, 27'h000001f4, 5'd21, 27'h000002fd, 32'h00000400,
  1'd1,  5'd23, 27'h00000314, 5'd13, 27'h0000030e, 5'd5, 27'h0000001d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000025e, 5'd12, 27'h0000039c, 5'd13, 27'h00000160, 32'h00000400,
  1'd1,  5'd20, 27'h00000304, 5'd10, 27'h00000314, 5'd20, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003a9, 5'd25, 27'h000002cc, 5'd4, 27'h000002fb, 32'h00000400,
  1'd1,  5'd25, 27'h00000245, 5'd24, 27'h000003f5, 5'd14, 27'h000000da, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000032e, 5'd21, 27'h00000246, 5'd21, 27'h000000f9, 32'h00000400,
  1'd1,  5'd4, 27'h0000009d, 5'd3, 27'h00000260, 5'd6, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003be, 5'd0, 27'h000001ed, 5'd17, 27'h0000000b, 32'h00000400,
  1'd1,  5'd2, 27'h0000006d, 5'd1, 27'h000002be, 5'd28, 27'h0000027c, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000022a, 5'd11, 27'h000002b3, 5'd8, 27'h000003b9, 32'h00000400,
  1'd1,  5'd5, 27'h00000032, 5'd11, 27'h0000022f, 5'd19, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000061, 5'd14, 27'h0000010f, 5'd27, 27'h0000007b, 32'h00000400,
  1'd1,  5'd2, 27'h00000167, 5'd24, 27'h00000149, 5'd9, 27'h00000065, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001a3, 5'd23, 27'h000001b1, 5'd15, 27'h00000308, 32'h00000400,
  1'd1,  5'd4, 27'h0000005c, 5'd21, 27'h000003ef, 5'd27, 27'h000003cd, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000221, 5'd0, 27'h00000343, 5'd5, 27'h000003f9, 32'h00000400,
  1'd1,  5'd12, 27'h00000260, 5'd2, 27'h0000016f, 5'd16, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000011d, 5'd3, 27'h000001cf, 5'd30, 27'h0000015b, 32'h00000400,
  1'd1,  5'd11, 27'h00000180, 5'd10, 27'h0000015b, 5'd8, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000312, 5'd12, 27'h00000311, 5'd20, 27'h00000135, 32'h00000400,
  1'd1,  5'd11, 27'h00000370, 5'd12, 27'h00000018, 5'd27, 27'h00000195, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000152, 5'd25, 27'h00000061, 5'd9, 27'h00000336, 32'h00000400,
  1'd1,  5'd12, 27'h0000029b, 5'd22, 27'h000001b5, 5'd18, 27'h000001f1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001c1, 5'd24, 27'h00000162, 5'd26, 27'h00000300, 32'h00000400,
  1'd1,  5'd23, 27'h00000310, 5'd0, 27'h000000db, 5'd7, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000393, 5'd1, 27'h00000387, 5'd19, 27'h0000020e, 32'h00000400,
  1'd1,  5'd22, 27'h0000039c, 5'd2, 27'h00000392, 5'd28, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003f4, 5'd15, 27'h000000a2, 5'd7, 27'h00000174, 32'h00000400,
  1'd1,  5'd23, 27'h00000104, 5'd12, 27'h00000213, 5'd17, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000009c, 5'd14, 27'h000002be, 5'd30, 27'h0000028c, 32'h00000400,
  1'd1,  5'd23, 27'h0000008c, 5'd23, 27'h00000081, 5'd10, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000a3, 5'd24, 27'h0000012b, 5'd17, 27'h000003c5, 32'h00000400,
  1'd1,  5'd21, 27'h0000031b, 5'd21, 27'h000001f0, 5'd30, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000019f, 5'd9, 27'h00000352, 5'd5, 27'h000000a9, 32'h00000400,
  1'd1,  5'd3, 27'h0000038a, 5'd8, 27'h000001bd, 5'd11, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000003f, 5'd10, 27'h00000025, 5'd23, 27'h00000132, 32'h00000400,
  1'd1,  5'd0, 27'h0000024f, 5'd20, 27'h000001f9, 5'd1, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000148, 5'd17, 27'h000003a7, 5'd13, 27'h000003dc, 32'h00000400,
  1'd1,  5'd0, 27'h00000313, 5'd17, 27'h00000196, 5'd24, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000330, 5'd29, 27'h000002bb, 5'd0, 27'h000001f9, 32'h00000400,
  1'd1,  5'd1, 27'h00000120, 5'd25, 27'h000003c9, 5'd11, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003e5, 5'd30, 27'h000002fa, 5'd22, 27'h000003ca, 32'h00000400,
  1'd1,  5'd10, 27'h0000038c, 5'd7, 27'h000001f4, 5'd2, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a4, 5'd7, 27'h00000400, 5'd11, 27'h000000bc, 32'h00000400,
  1'd1,  5'd10, 27'h0000027f, 5'd7, 27'h00000221, 5'd21, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d5, 5'd20, 27'h000001e1, 5'd2, 27'h0000037d, 32'h00000400,
  1'd1,  5'd11, 27'h00000143, 5'd18, 27'h00000234, 5'd15, 27'h000000d6, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000d0, 5'd16, 27'h000000c5, 5'd23, 27'h0000012b, 32'h00000400,
  1'd1,  5'd11, 27'h00000245, 5'd28, 27'h00000261, 5'd1, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003bf, 5'd28, 27'h00000049, 5'd13, 27'h0000009d, 32'h00000400,
  1'd1,  5'd11, 27'h000003f6, 5'd30, 27'h00000040, 5'd23, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003ab, 5'd7, 27'h00000114, 5'd0, 27'h00000163, 32'h00000400,
  1'd1,  5'd23, 27'h000001e8, 5'd9, 27'h0000017a, 5'd12, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000324, 5'd17, 27'h000002f2, 5'd2, 27'h000001e3, 32'h00000400,
  1'd1,  5'd22, 27'h000000fe, 5'd18, 27'h0000032e, 5'd15, 27'h000000b5, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000011c, 5'd17, 27'h000001c5, 5'd24, 27'h000003b5, 32'h00000400,
  1'd1,  5'd22, 27'h00000238, 5'd30, 27'h000003de, 5'd2, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003b3, 5'd27, 27'h00000009, 5'd13, 27'h00000159, 32'h00000400,
  1'd1,  5'd24, 27'h000001be, 5'd30, 27'h00000279, 5'd24, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000023c, 5'd9, 27'h000001e4, 5'd10, 27'h000000c3, 32'h00000400,
  1'd1,  5'd3, 27'h000002c6, 5'd6, 27'h00000312, 5'd20, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000017a, 5'd9, 27'h000002d1, 5'd29, 27'h000003db, 32'h00000400,
  1'd1,  5'd2, 27'h00000261, 5'd18, 27'h0000022d, 5'd6, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003b4, 5'd20, 27'h0000002d, 5'd19, 27'h000001d4, 32'h00000400,
  1'd1,  5'd0, 27'h000000fb, 5'd15, 27'h00000293, 5'd26, 27'h00000122, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003bd, 5'd26, 27'h00000389, 5'd8, 27'h0000033b, 32'h00000400,
  1'd1,  5'd1, 27'h0000026d, 5'd27, 27'h000003bd, 5'd16, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002dd, 5'd30, 27'h000000d9, 5'd28, 27'h00000091, 32'h00000400,
  1'd1,  5'd11, 27'h000001b5, 5'd5, 27'h000001ac, 5'd8, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001b6, 5'd8, 27'h00000214, 5'd19, 27'h00000088, 32'h00000400,
  1'd1,  5'd11, 27'h00000360, 5'd6, 27'h000001bf, 5'd28, 27'h000000ba, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e5, 5'd17, 27'h0000011b, 5'd9, 27'h00000270, 32'h00000400,
  1'd1,  5'd11, 27'h00000068, 5'd15, 27'h00000283, 5'd19, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000265, 5'd19, 27'h0000023d, 5'd29, 27'h00000174, 32'h00000400,
  1'd1,  5'd11, 27'h00000359, 5'd30, 27'h0000011b, 5'd6, 27'h000002cd, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003d5, 5'd27, 27'h000002ea, 5'd15, 27'h00000296, 32'h00000400,
  1'd1,  5'd15, 27'h00000143, 5'd26, 27'h000001d2, 5'd26, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000031e, 5'd7, 27'h00000144, 5'd9, 27'h00000155, 32'h00000400,
  1'd1,  5'd25, 27'h00000083, 5'd7, 27'h00000112, 5'd17, 27'h000003b5, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000058, 5'd9, 27'h000002fe, 5'd30, 27'h0000038d, 32'h00000400,
  1'd1,  5'd21, 27'h0000017b, 5'd18, 27'h00000021, 5'd9, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000265, 5'd16, 27'h00000183, 5'd20, 27'h0000017e, 32'h00000400,
  1'd1,  5'd20, 27'h0000037f, 5'd15, 27'h000003e3, 5'd28, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000008, 5'd26, 27'h00000156, 5'd8, 27'h000002ad, 32'h00000400,
  1'd1,  5'd21, 27'h00000188, 5'd30, 27'h00000247, 5'd17, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000022a, 5'd27, 27'h00000371, 5'd29, 27'h00000056, 32'h00000400,
  1'd1,  5'd6, 27'h000000ff, 5'd3, 27'h0000008d, 5'd5, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d4, 5'd1, 27'h00000081, 5'd17, 27'h000002bd, 32'h00000400,
  1'd1,  5'd6, 27'h0000011f, 5'd0, 27'h0000011e, 5'd26, 27'h00000202, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000098, 5'd11, 27'h000002d0, 5'd3, 27'h000000dc, 32'h00000400,
  1'd1,  5'd8, 27'h0000012e, 5'd10, 27'h00000164, 5'd12, 27'h000001cf, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001e0, 5'd12, 27'h000003c1, 5'd22, 27'h000001ee, 32'h00000400,
  1'd1,  5'd7, 27'h000002ea, 5'd25, 27'h00000143, 5'd3, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000069, 5'd21, 27'h000001b5, 5'd13, 27'h000002ac, 32'h00000400,
  1'd1,  5'd8, 27'h00000316, 5'd24, 27'h000001fb, 5'd25, 27'h00000006, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e7, 5'd1, 27'h00000002, 5'd7, 27'h000000f6, 32'h00000400,
  1'd1,  5'd20, 27'h0000002d, 5'd4, 27'h0000029d, 5'd16, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000079, 5'd2, 27'h000002b7, 5'd28, 27'h00000118, 32'h00000400,
  1'd1,  5'd16, 27'h000002aa, 5'd13, 27'h0000033c, 5'd4, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000321, 5'd10, 27'h0000024b, 5'd13, 27'h00000096, 32'h00000400,
  1'd1,  5'd19, 27'h000000d4, 5'd10, 27'h00000199, 5'd24, 27'h000000a8, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001c6, 5'd24, 27'h000003ec, 5'd3, 27'h0000005a, 32'h00000400,
  1'd1,  5'd16, 27'h000000eb, 5'd22, 27'h0000004e, 5'd11, 27'h00000314, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000175, 5'd21, 27'h000003c7, 5'd21, 27'h0000017d, 32'h00000400,
  1'd1,  5'd30, 27'h000002a2, 5'd0, 27'h000000f0, 5'd0, 27'h000002e3, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003c7, 5'd2, 27'h0000004d, 5'd11, 27'h00000092, 32'h00000400,
  1'd1,  5'd30, 27'h000000d1, 5'd4, 27'h00000325, 5'd21, 27'h000000c6, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000244, 5'd15, 27'h000001d5, 5'd2, 27'h000000e6, 32'h00000400,
  1'd1,  5'd28, 27'h000000a9, 5'd14, 27'h00000219, 5'd14, 27'h000003b0, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000009a, 5'd11, 27'h000002d1, 5'd25, 27'h00000154, 32'h00000400,
  1'd1,  5'd27, 27'h000000b0, 5'd23, 27'h000001fc, 5'd4, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000390, 5'd23, 27'h000002d9, 5'd13, 27'h00000171, 32'h00000400,
  1'd1,  5'd29, 27'h000000d0, 5'd24, 27'h00000107, 5'd22, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002aa, 5'd1, 27'h00000177, 5'd1, 27'h00000338, 32'h00000400,
  1'd1,  5'd6, 27'h0000000a, 5'd3, 27'h000000f8, 5'd12, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000016b, 5'd1, 27'h00000061, 5'd23, 27'h00000269, 32'h00000400,
  1'd1,  5'd8, 27'h00000082, 5'd15, 27'h0000002b, 5'd9, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000398, 5'd13, 27'h000003d4, 5'd17, 27'h00000309, 32'h00000400,
  1'd1,  5'd5, 27'h000003ef, 5'd10, 27'h00000371, 5'd29, 27'h0000011a, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002e5, 5'd22, 27'h000000f1, 5'd8, 27'h00000335, 32'h00000400,
  1'd1,  5'd9, 27'h00000128, 5'd21, 27'h000000f5, 5'd17, 27'h00000087, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001ff, 5'd24, 27'h000000ed, 5'd28, 27'h0000023c, 32'h00000400,
  1'd1,  5'd19, 27'h00000236, 5'd3, 27'h0000034b, 5'd1, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003f2, 5'd1, 27'h000003dd, 5'd10, 27'h0000028d, 32'h00000400,
  1'd1,  5'd19, 27'h00000146, 5'd14, 27'h00000118, 5'd8, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000ab, 5'd14, 27'h000000f6, 5'd19, 27'h0000030b, 32'h00000400,
  1'd1,  5'd15, 27'h0000026e, 5'd15, 27'h000000d5, 5'd30, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000225, 5'd25, 27'h000001e7, 5'd9, 27'h000001a7, 32'h00000400,
  1'd1,  5'd17, 27'h00000363, 5'd23, 27'h00000298, 5'd20, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000066, 5'd23, 27'h000000ce, 5'd25, 27'h000003db, 32'h00000400,
  1'd1,  5'd30, 27'h000002bb, 5'd3, 27'h00000283, 5'd7, 27'h00000086, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000387, 5'd0, 27'h000002db, 5'd18, 27'h00000225, 32'h00000400,
  1'd1,  5'd29, 27'h00000261, 5'd4, 27'h0000005a, 5'd30, 27'h000003c6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003f7, 5'd10, 27'h000002e1, 5'd8, 27'h0000002c, 32'h00000400,
  1'd1,  5'd30, 27'h00000159, 5'd12, 27'h0000000d, 5'd15, 27'h000003bf, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000154, 5'd12, 27'h00000046, 5'd30, 27'h0000033e, 32'h00000400,
  1'd1,  5'd26, 27'h000002ae, 5'd21, 27'h000003f6, 5'd10, 27'h000000d7, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002c1, 5'd25, 27'h000002fd, 5'd17, 27'h000001c1, 32'h00000400,
  1'd1,  5'd30, 27'h00000187, 5'd22, 27'h000000f3, 5'd30, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000130, 5'd8, 27'h00000106, 5'd2, 27'h000000be, 32'h00000400,
  1'd1,  5'd7, 27'h000001a3, 5'd6, 27'h000000a2, 5'd14, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000306, 5'd8, 27'h000000ce, 5'd24, 27'h00000100, 32'h00000400,
  1'd1,  5'd5, 27'h000003d0, 5'd19, 27'h000001d6, 5'd2, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000037, 5'd15, 27'h000002da, 5'd12, 27'h000003fc, 32'h00000400,
  1'd1,  5'd8, 27'h0000005d, 5'd15, 27'h00000277, 5'd24, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000196, 5'd26, 27'h000001c7, 5'd4, 27'h0000026d, 32'h00000400,
  1'd1,  5'd8, 27'h0000013c, 5'd27, 27'h00000021, 5'd10, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000022e, 5'd29, 27'h00000283, 5'd21, 27'h0000011f, 32'h00000400,
  1'd1,  5'd16, 27'h000000b2, 5'd9, 27'h00000152, 5'd1, 27'h0000031c, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000005d, 5'd9, 27'h000001d1, 5'd10, 27'h000001eb, 32'h00000400,
  1'd1,  5'd16, 27'h00000072, 5'd5, 27'h000000d8, 5'd23, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000028f, 5'd17, 27'h000001fe, 5'd1, 27'h00000191, 32'h00000400,
  1'd1,  5'd19, 27'h0000028c, 5'd20, 27'h000001c2, 5'd13, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000bd, 5'd15, 27'h000003db, 5'd21, 27'h00000053, 32'h00000400,
  1'd1,  5'd20, 27'h000001f8, 5'd30, 27'h000003d3, 5'd2, 27'h00000020, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000022a, 5'd27, 27'h000003d5, 5'd13, 27'h000001fe, 32'h00000400,
  1'd1,  5'd17, 27'h000002fb, 5'd28, 27'h00000032, 5'd20, 27'h00000347, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003e6, 5'd7, 27'h0000027d, 5'd2, 27'h000003d0, 32'h00000400,
  1'd1,  5'd26, 27'h000003d3, 5'd6, 27'h00000122, 5'd14, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000033a, 5'd5, 27'h00000390, 5'd24, 27'h0000017a, 32'h00000400,
  1'd1,  5'd25, 27'h000003ef, 5'd19, 27'h000003a4, 5'd0, 27'h000003bc, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002a0, 5'd16, 27'h000000de, 5'd11, 27'h000003a3, 32'h00000400,
  1'd1,  5'd26, 27'h0000016a, 5'd16, 27'h0000013d, 5'd23, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002a5, 5'd27, 27'h0000002a, 5'd1, 27'h00000218, 32'h00000400,
  1'd1,  5'd28, 27'h00000398, 5'd29, 27'h0000020e, 5'd11, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000064, 5'd27, 27'h000002f8, 5'd23, 27'h0000014a, 32'h00000400,
  1'd1,  5'd8, 27'h00000038, 5'd9, 27'h00000085, 5'd9, 27'h00000178, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000331, 5'd6, 27'h000001c2, 5'd16, 27'h00000312, 32'h00000400,
  1'd1,  5'd8, 27'h00000382, 5'd7, 27'h00000370, 5'd27, 27'h00000285, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000194, 5'd19, 27'h00000109, 5'd6, 27'h0000016a, 32'h00000400,
  1'd1,  5'd9, 27'h00000030, 5'd17, 27'h000001ce, 5'd20, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ff, 5'd17, 27'h00000286, 5'd28, 27'h000000c8, 32'h00000400,
  1'd1,  5'd7, 27'h00000069, 5'd28, 27'h0000014f, 5'd8, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000009, 5'd30, 27'h000001cb, 5'd20, 27'h000000b4, 32'h00000400,
  1'd1,  5'd9, 27'h00000233, 5'd28, 27'h000002eb, 5'd30, 27'h000000e8, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000001e, 5'd5, 27'h000001a1, 5'd6, 27'h0000022a, 32'h00000400,
  1'd1,  5'd15, 27'h0000026d, 5'd5, 27'h000003a7, 5'd18, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000004e, 5'd8, 27'h000003cc, 5'd28, 27'h00000207, 32'h00000400,
  1'd1,  5'd18, 27'h00000292, 5'd18, 27'h0000000c, 5'd6, 27'h000003ed, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000032e, 5'd16, 27'h000001eb, 5'd15, 27'h00000264, 32'h00000400,
  1'd1,  5'd19, 27'h000001af, 5'd16, 27'h000001a3, 5'd28, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000117, 5'd27, 27'h000002c8, 5'd6, 27'h000002f6, 32'h00000400,
  1'd1,  5'd18, 27'h0000020f, 5'd29, 27'h00000051, 5'd17, 27'h00000277, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000049, 5'd26, 27'h0000036d, 5'd30, 27'h000003ce, 32'h00000400,
  1'd1,  5'd27, 27'h000001a9, 5'd7, 27'h0000017a, 5'd6, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000016f, 5'd8, 27'h00000087, 5'd16, 27'h0000039b, 32'h00000400,
  1'd1,  5'd29, 27'h00000156, 5'd9, 27'h00000257, 5'd30, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000b2, 5'd20, 27'h00000290, 5'd6, 27'h000001db, 32'h00000400,
  1'd1,  5'd26, 27'h00000195, 5'd17, 27'h000002b7, 5'd15, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000011f, 5'd20, 27'h000002a4, 5'd27, 27'h0000018c, 32'h00000400,
  1'd1,  5'd27, 27'h0000005c, 5'd27, 27'h000000d5, 5'd8, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000028e, 5'd29, 27'h00000116, 5'd16, 27'h00000112, 32'h00000400,
  1'd1,  5'd25, 27'h000003e2, 5'd27, 27'h000003c4, 5'd26, 27'h000001e5, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000003f0, 5'd4, 27'h0000006a, 5'd3, 27'h00000203, 32'h00000400,
  1'd1,  5'd3, 27'h00000231, 5'd1, 27'h0000004e, 5'd15, 27'h00000034, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001a3, 5'd0, 27'h000001d9, 5'd23, 27'h00000103, 32'h00000400,
  1'd1,  5'd1, 27'h0000009f, 5'd13, 27'h0000014a, 5'd1, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003d3, 5'd15, 27'h00000092, 5'd12, 27'h000003da, 32'h00000400,
  1'd1,  5'd2, 27'h000003fc, 5'd12, 27'h000000ea, 5'd25, 27'h00000326, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000001f, 5'd22, 27'h000002f3, 5'd2, 27'h000003da, 32'h00000400,
  1'd1,  5'd4, 27'h00000254, 5'd23, 27'h000003ff, 5'd15, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000396, 5'd24, 27'h00000143, 5'd23, 27'h0000034a, 32'h00000400,
  1'd1,  5'd12, 27'h0000001f, 5'd4, 27'h00000065, 5'd0, 27'h00000193, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002fd, 5'd1, 27'h000003f3, 5'd11, 27'h0000020b, 32'h00000400,
  1'd1,  5'd11, 27'h000003a6, 5'd1, 27'h0000036c, 5'd20, 27'h00000309, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000da, 5'd11, 27'h000003c9, 5'd1, 27'h000001f5, 32'h00000400,
  1'd1,  5'd14, 27'h00000335, 5'd12, 27'h00000169, 5'd15, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000035, 5'd11, 27'h00000235, 5'd22, 27'h0000039a, 32'h00000400,
  1'd1,  5'd13, 27'h000000e8, 5'd24, 27'h00000079, 5'd1, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000193, 5'd24, 27'h00000332, 5'd12, 27'h0000004d, 32'h00000400,
  1'd1,  5'd10, 27'h000002af, 5'd22, 27'h000001d7, 5'd22, 27'h00000080, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000100, 5'd1, 27'h0000003a, 5'd4, 27'h00000280, 32'h00000400,
  1'd1,  5'd23, 27'h00000268, 5'd1, 27'h000003eb, 5'd10, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000036, 5'd0, 27'h000001b8, 5'd22, 27'h0000039a, 32'h00000400,
  1'd1,  5'd23, 27'h000002ce, 5'd13, 27'h00000096, 5'd4, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000305, 5'd15, 27'h0000012b, 5'd10, 27'h0000027f, 32'h00000400,
  1'd1,  5'd21, 27'h000001e4, 5'd10, 27'h0000015a, 5'd24, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002c5, 5'd25, 27'h00000300, 5'd0, 27'h00000350, 32'h00000400,
  1'd1,  5'd20, 27'h000003f5, 5'd24, 27'h0000012a, 5'd15, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000143, 5'd25, 27'h00000121, 5'd24, 27'h00000256, 32'h00000400,
  1'd1,  5'd2, 27'h000003ad, 5'd0, 27'h000001d9, 5'd8, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a9, 5'd3, 27'h00000060, 5'd18, 27'h00000023, 32'h00000400,
  1'd1,  5'd1, 27'h00000330, 5'd3, 27'h00000133, 5'd29, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002c8, 5'd10, 27'h000001d3, 5'd8, 27'h0000012a, 32'h00000400,
  1'd1,  5'd3, 27'h00000225, 5'd11, 27'h0000008d, 5'd19, 27'h0000029f, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001a0, 5'd14, 27'h000000c7, 5'd26, 27'h00000387, 32'h00000400,
  1'd1,  5'd0, 27'h00000349, 5'd24, 27'h0000007a, 5'd6, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003ea, 5'd24, 27'h00000302, 5'd18, 27'h000002d2, 32'h00000400,
  1'd1,  5'd0, 27'h0000020e, 5'd25, 27'h00000214, 5'd26, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c5, 5'd2, 27'h000003d0, 5'd10, 27'h00000099, 32'h00000400,
  1'd1,  5'd12, 27'h00000323, 5'd3, 27'h00000082, 5'd18, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002e4, 5'd3, 27'h000002a7, 5'd26, 27'h00000022, 32'h00000400,
  1'd1,  5'd10, 27'h00000348, 5'd11, 27'h00000166, 5'd9, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d6, 5'd11, 27'h000002bf, 5'd18, 27'h00000147, 32'h00000400,
  1'd1,  5'd11, 27'h00000385, 5'd11, 27'h000001e7, 5'd26, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000231, 5'd24, 27'h000001ac, 5'd9, 27'h0000012c, 32'h00000400,
  1'd1,  5'd13, 27'h00000153, 5'd24, 27'h0000004e, 5'd19, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000266, 5'd22, 27'h00000307, 5'd27, 27'h00000154, 32'h00000400,
  1'd1,  5'd21, 27'h00000316, 5'd0, 27'h000003a1, 5'd7, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000010a, 5'd0, 27'h0000019d, 5'd20, 27'h000001c7, 32'h00000400,
  1'd1,  5'd22, 27'h00000250, 5'd0, 27'h00000250, 5'd26, 27'h0000026e, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002be, 5'd13, 27'h00000204, 5'd7, 27'h00000242, 32'h00000400,
  1'd1,  5'd20, 27'h00000323, 5'd12, 27'h00000168, 5'd16, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000d5, 5'd13, 27'h000003d7, 5'd28, 27'h000000bb, 32'h00000400,
  1'd1,  5'd21, 27'h000002f9, 5'd24, 27'h000000b7, 5'd8, 27'h00000367, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003c7, 5'd21, 27'h000002f3, 5'd18, 27'h00000008, 32'h00000400,
  1'd1,  5'd25, 27'h00000261, 5'd22, 27'h00000064, 5'd30, 27'h00000192, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001df, 5'd9, 27'h0000033e, 5'd0, 27'h000001c4, 32'h00000400,
  1'd1,  5'd2, 27'h00000110, 5'd8, 27'h000003dd, 5'd12, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002c9, 5'd5, 27'h000000ef, 5'd24, 27'h000000a7, 32'h00000400,
  1'd1,  5'd3, 27'h00000171, 5'd20, 27'h00000022, 5'd3, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000007f, 5'd18, 27'h00000183, 5'd11, 27'h0000030c, 32'h00000400,
  1'd1,  5'd3, 27'h0000000d, 5'd18, 27'h0000019d, 5'd24, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000058, 5'd28, 27'h000000a6, 5'd3, 27'h00000010, 32'h00000400,
  1'd1,  5'd4, 27'h000003e3, 5'd26, 27'h00000136, 5'd10, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000335, 5'd27, 27'h000002ba, 5'd22, 27'h000003bc, 32'h00000400,
  1'd1,  5'd12, 27'h000003a0, 5'd5, 27'h000001cc, 5'd1, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e8, 5'd7, 27'h0000015c, 5'd10, 27'h000001ec, 32'h00000400,
  1'd1,  5'd12, 27'h000003a4, 5'd6, 27'h0000037a, 5'd23, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000015f, 5'd16, 27'h00000194, 5'd4, 27'h000003e9, 32'h00000400,
  1'd1,  5'd12, 27'h000000e1, 5'd20, 27'h000001c6, 5'd11, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f1, 5'd17, 27'h000000d1, 5'd24, 27'h00000352, 32'h00000400,
  1'd1,  5'd13, 27'h000000a6, 5'd28, 27'h00000330, 5'd4, 27'h00000358, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000030b, 5'd29, 27'h000003fe, 5'd15, 27'h00000112, 32'h00000400,
  1'd1,  5'd14, 27'h000001d6, 5'd29, 27'h00000330, 5'd23, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001e2, 5'd8, 27'h00000146, 5'd4, 27'h000003b4, 32'h00000400,
  1'd1,  5'd21, 27'h0000020b, 5'd9, 27'h000002bf, 5'd12, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000256, 5'd16, 27'h000000ab, 5'd2, 27'h00000310, 32'h00000400,
  1'd1,  5'd21, 27'h00000225, 5'd15, 27'h0000034c, 5'd10, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000025a, 5'd19, 27'h0000015e, 5'd24, 27'h00000124, 32'h00000400,
  1'd1,  5'd24, 27'h0000003a, 5'd30, 27'h00000319, 5'd2, 27'h0000011e, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000004d, 5'd27, 27'h00000136, 5'd11, 27'h000000b9, 32'h00000400,
  1'd1,  5'd23, 27'h000001e3, 5'd27, 27'h00000093, 5'd20, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002a, 5'd7, 27'h00000017, 5'd8, 27'h000000ff, 32'h00000400,
  1'd1,  5'd0, 27'h00000275, 5'd10, 27'h00000070, 5'd20, 27'h000001c6, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000011a, 5'd9, 27'h00000135, 5'd28, 27'h00000216, 32'h00000400,
  1'd1,  5'd1, 27'h00000374, 5'd20, 27'h00000123, 5'd7, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000023, 5'd17, 27'h0000018a, 5'd18, 27'h0000003a, 32'h00000400,
  1'd1,  5'd1, 27'h000000ff, 5'd20, 27'h000000fc, 5'd27, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd1, 27'h000003f7, 5'd28, 27'h00000321, 5'd8, 27'h000000e5, 32'h00000400,
  1'd1,  5'd3, 27'h0000015d, 5'd29, 27'h0000003e, 5'd18, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000168, 5'd28, 27'h000000c4, 5'd26, 27'h000000e4, 32'h00000400,
  1'd1,  5'd12, 27'h00000315, 5'd7, 27'h00000006, 5'd5, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000026b, 5'd9, 27'h00000055, 5'd17, 27'h000003ff, 32'h00000400,
  1'd1,  5'd13, 27'h000000bb, 5'd5, 27'h000000b5, 5'd27, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002d3, 5'd18, 27'h00000161, 5'd9, 27'h000002aa, 32'h00000400,
  1'd1,  5'd11, 27'h00000153, 5'd17, 27'h00000217, 5'd19, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000002f, 5'd18, 27'h00000329, 5'd28, 27'h0000010b, 32'h00000400,
  1'd1,  5'd15, 27'h00000113, 5'd26, 27'h00000029, 5'd10, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000255, 5'd27, 27'h00000117, 5'd19, 27'h00000367, 32'h00000400,
  1'd1,  5'd12, 27'h00000086, 5'd30, 27'h00000032, 5'd27, 27'h000003a4, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000027, 5'd5, 27'h00000338, 5'd9, 27'h0000003f, 32'h00000400,
  1'd1,  5'd24, 27'h0000014a, 5'd6, 27'h000001c6, 5'd17, 27'h00000002, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d7, 5'd9, 27'h000002e7, 5'd29, 27'h00000357, 32'h00000400,
  1'd1,  5'd22, 27'h00000001, 5'd18, 27'h00000346, 5'd6, 27'h000000b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c6, 5'd18, 27'h00000366, 5'd18, 27'h00000194, 32'h00000400,
  1'd1,  5'd23, 27'h0000015c, 5'd20, 27'h0000013f, 5'd29, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000025a, 5'd28, 27'h0000038d, 5'd8, 27'h00000172, 32'h00000400,
  1'd1,  5'd23, 27'h000002af, 5'd26, 27'h00000237, 5'd19, 27'h0000032f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000ba, 5'd26, 27'h00000049, 5'd27, 27'h000002d6, 32'h00000400,
  1'd1,  5'd9, 27'h00000135, 5'd2, 27'h000000b7, 5'd7, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000fb, 5'd1, 27'h0000035f, 5'd19, 27'h00000300, 32'h00000400,
  1'd1,  5'd7, 27'h000003f4, 5'd2, 27'h0000032b, 5'd28, 27'h000001ff, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000148, 5'd10, 27'h000001e0, 5'd2, 27'h00000265, 32'h00000400,
  1'd1,  5'd10, 27'h00000083, 5'd13, 27'h000002b2, 5'd13, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003da, 5'd12, 27'h000001ca, 5'd24, 27'h000003fe, 32'h00000400,
  1'd1,  5'd7, 27'h0000035b, 5'd25, 27'h0000008c, 5'd4, 27'h00000156, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011e, 5'd25, 27'h000000e1, 5'd15, 27'h000001ea, 32'h00000400,
  1'd1,  5'd8, 27'h00000126, 5'd21, 27'h0000010f, 5'd25, 27'h000002c3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000d9, 5'd0, 27'h000001ee, 5'd9, 27'h000001ec, 32'h00000400,
  1'd1,  5'd17, 27'h000003d5, 5'd1, 27'h000000b7, 5'd16, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000cf, 5'd3, 27'h00000181, 5'd28, 27'h00000388, 32'h00000400,
  1'd1,  5'd16, 27'h000000ad, 5'd13, 27'h000000b0, 5'd1, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000255, 5'd12, 27'h0000017c, 5'd14, 27'h000002ff, 32'h00000400,
  1'd1,  5'd18, 27'h0000008d, 5'd11, 27'h0000014f, 5'd24, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003d7, 5'd23, 27'h0000025c, 5'd3, 27'h00000323, 32'h00000400,
  1'd1,  5'd17, 27'h00000139, 5'd22, 27'h000002ea, 5'd14, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002f7, 5'd22, 27'h00000344, 5'd25, 27'h00000031, 32'h00000400,
  1'd1,  5'd30, 27'h000001b7, 5'd4, 27'h00000013, 5'd2, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000224, 5'd4, 27'h00000107, 5'd12, 27'h00000163, 32'h00000400,
  1'd1,  5'd29, 27'h00000309, 5'd1, 27'h0000018f, 5'd24, 27'h00000334, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ba, 5'd11, 27'h0000024d, 5'd4, 27'h00000306, 32'h00000400,
  1'd1,  5'd26, 27'h000002c8, 5'd15, 27'h00000087, 5'd13, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd29, 27'h000000f8, 5'd15, 27'h000001f0, 5'd22, 27'h0000030e, 32'h00000400,
  1'd1,  5'd26, 27'h00000066, 5'd23, 27'h000002b9, 5'd3, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000024e, 5'd25, 27'h00000286, 5'd12, 27'h0000005f, 32'h00000400,
  1'd1,  5'd29, 27'h000002d0, 5'd22, 27'h000002bb, 5'd22, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021b, 5'd0, 27'h000000c1, 5'd3, 27'h00000126, 32'h00000400,
  1'd1,  5'd8, 27'h00000034, 5'd1, 27'h000002b9, 5'd12, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000049, 5'd2, 27'h00000044, 5'd25, 27'h00000047, 32'h00000400,
  1'd1,  5'd7, 27'h000000ef, 5'd10, 27'h000002f1, 5'd7, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000356, 5'd15, 27'h000000c0, 5'd19, 27'h00000106, 32'h00000400,
  1'd1,  5'd7, 27'h0000014a, 5'd11, 27'h00000184, 5'd27, 27'h00000032, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000251, 5'd24, 27'h0000011f, 5'd9, 27'h000003cb, 32'h00000400,
  1'd1,  5'd5, 27'h0000010e, 5'd23, 27'h0000018e, 5'd16, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000002c, 5'd25, 27'h0000011d, 5'd25, 27'h00000362, 32'h00000400,
  1'd1,  5'd20, 27'h000001bf, 5'd2, 27'h00000215, 5'd3, 27'h000003e5, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000301, 5'd3, 27'h000003f0, 5'd10, 27'h000002aa, 32'h00000400,
  1'd1,  5'd17, 27'h00000067, 5'd10, 27'h000001d6, 5'd7, 27'h00000083, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001c9, 5'd13, 27'h00000282, 5'd20, 27'h000001f9, 32'h00000400,
  1'd1,  5'd16, 27'h0000039c, 5'd14, 27'h00000222, 5'd26, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000008b, 5'd24, 27'h0000002d, 5'd9, 27'h00000128, 32'h00000400,
  1'd1,  5'd17, 27'h00000227, 5'd21, 27'h00000021, 5'd15, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000367, 5'd20, 27'h000003ae, 5'd26, 27'h00000243, 32'h00000400,
  1'd1,  5'd25, 27'h0000039a, 5'd1, 27'h00000154, 5'd9, 27'h0000019b, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000027, 5'd3, 27'h000001d9, 5'd16, 27'h000003b4, 32'h00000400,
  1'd1,  5'd29, 27'h0000023d, 5'd2, 27'h00000370, 5'd28, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000237, 5'd10, 27'h000001ae, 5'd10, 27'h00000125, 32'h00000400,
  1'd1,  5'd26, 27'h0000031b, 5'd14, 27'h0000012e, 5'd20, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000275, 5'd13, 27'h000000e4, 5'd27, 27'h00000208, 32'h00000400,
  1'd1,  5'd30, 27'h000003c5, 5'd23, 27'h000000de, 5'd9, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000302, 5'd21, 27'h0000021f, 5'd17, 27'h0000004d, 32'h00000400,
  1'd1,  5'd27, 27'h000003a2, 5'd24, 27'h00000285, 5'd26, 27'h000000fa, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000050, 5'd6, 27'h000002a4, 5'd3, 27'h000003fe, 32'h00000400,
  1'd1,  5'd6, 27'h00000030, 5'd7, 27'h00000153, 5'd12, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000039a, 5'd9, 27'h000001ce, 5'd25, 27'h000001e0, 32'h00000400,
  1'd1,  5'd10, 27'h00000030, 5'd20, 27'h00000034, 5'd2, 27'h0000005c, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000012c, 5'd17, 27'h00000121, 5'd10, 27'h000002f6, 32'h00000400,
  1'd1,  5'd8, 27'h0000024d, 5'd15, 27'h0000023b, 5'd24, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000352, 5'd27, 27'h000003ca, 5'd4, 27'h00000030, 32'h00000400,
  1'd1,  5'd10, 27'h000000ab, 5'd28, 27'h000000e6, 5'd14, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000311, 5'd30, 27'h0000007a, 5'd25, 27'h0000032e, 32'h00000400,
  1'd1,  5'd16, 27'h0000013f, 5'd10, 27'h00000138, 5'd2, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000231, 5'd8, 27'h00000302, 5'd12, 27'h000002b1, 32'h00000400,
  1'd1,  5'd17, 27'h000000c0, 5'd7, 27'h000002bd, 5'd24, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c4, 5'd17, 27'h000001b0, 5'd0, 27'h00000030, 32'h00000400,
  1'd1,  5'd16, 27'h0000014e, 5'd16, 27'h00000223, 5'd14, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000d2, 5'd17, 27'h00000268, 5'd21, 27'h00000044, 32'h00000400,
  1'd1,  5'd18, 27'h000001bd, 5'd26, 27'h0000009c, 5'd1, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001ea, 5'd29, 27'h000000e0, 5'd14, 27'h0000011a, 32'h00000400,
  1'd1,  5'd20, 27'h00000168, 5'd25, 27'h0000038f, 5'd20, 27'h000003a5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003b7, 5'd9, 27'h00000221, 5'd1, 27'h00000261, 32'h00000400,
  1'd1,  5'd28, 27'h00000302, 5'd10, 27'h000000c0, 5'd10, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003f5, 5'd8, 27'h0000020f, 5'd24, 27'h000000d4, 32'h00000400,
  1'd1,  5'd28, 27'h00000366, 5'd18, 27'h00000368, 5'd4, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000038a, 5'd17, 27'h000003a3, 5'd13, 27'h000000f4, 32'h00000400,
  1'd1,  5'd29, 27'h0000033d, 5'd18, 27'h000000cc, 5'd25, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000363, 5'd30, 27'h000000e1, 5'd4, 27'h000001f5, 32'h00000400,
  1'd1,  5'd30, 27'h00000302, 5'd30, 27'h000001e0, 5'd10, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000205, 5'd28, 27'h0000023f, 5'd22, 27'h000000d2, 32'h00000400,
  1'd1,  5'd7, 27'h000001b5, 5'd7, 27'h000002a1, 5'd7, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000292, 5'd5, 27'h00000108, 5'd20, 27'h0000020f, 32'h00000400,
  1'd1,  5'd6, 27'h000001ee, 5'd7, 27'h000001e6, 5'd29, 27'h0000001e, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a2, 5'd16, 27'h000003a9, 5'd5, 27'h0000033a, 32'h00000400,
  1'd1,  5'd5, 27'h000001e8, 5'd17, 27'h000001cc, 5'd17, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001fd, 5'd16, 27'h000002b8, 5'd26, 27'h00000087, 32'h00000400,
  1'd1,  5'd6, 27'h000000c1, 5'd29, 27'h000001b5, 5'd5, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000146, 5'd29, 27'h00000247, 5'd17, 27'h00000307, 32'h00000400,
  1'd1,  5'd8, 27'h00000327, 5'd28, 27'h000001e9, 5'd30, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001bf, 5'd7, 27'h000001ec, 5'd5, 27'h00000213, 32'h00000400,
  1'd1,  5'd19, 27'h00000122, 5'd9, 27'h000000a2, 5'd19, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000330, 5'd7, 27'h000002cb, 5'd30, 27'h000001f4, 32'h00000400,
  1'd1,  5'd18, 27'h000002ae, 5'd20, 27'h00000240, 5'd8, 27'h00000351, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002b5, 5'd20, 27'h0000011f, 5'd17, 27'h0000025f, 32'h00000400,
  1'd1,  5'd19, 27'h000001d2, 5'd15, 27'h000002a8, 5'd28, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000027b, 5'd28, 27'h000001f4, 5'd6, 27'h00000262, 32'h00000400,
  1'd1,  5'd19, 27'h00000230, 5'd28, 27'h00000045, 5'd19, 27'h00000287, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e6, 5'd26, 27'h0000028e, 5'd25, 27'h000003bf, 32'h00000400,
  1'd1,  5'd28, 27'h00000052, 5'd6, 27'h0000028f, 5'd6, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003f5, 5'd9, 27'h00000091, 5'd16, 27'h00000273, 32'h00000400,
  1'd1,  5'd30, 27'h000001ec, 5'd6, 27'h000001a3, 5'd30, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000288, 5'd20, 27'h000000a9, 5'd9, 27'h000000e4, 32'h00000400,
  1'd1,  5'd26, 27'h000003c0, 5'd19, 27'h00000361, 5'd16, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000030f, 5'd20, 27'h0000027d, 5'd26, 27'h00000061, 32'h00000400,
  1'd1,  5'd26, 27'h00000154, 5'd29, 27'h000000d7, 5'd5, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000037c, 5'd28, 27'h000002ca, 5'd16, 27'h00000209, 32'h00000400,
  1'd1,  5'd25, 27'h00000363, 5'd29, 27'h0000008b, 5'd29, 27'h000002c1, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd3, 27'h0000013e, 5'd3, 27'h00000132, 5'd0, 27'h000000e9, 32'h00000400,
  1'd1,  5'd0, 27'h000003d6, 5'd2, 27'h000001c6, 5'd11, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000013e, 5'd2, 27'h000003b3, 5'd23, 27'h0000014c, 32'h00000400,
  1'd1,  5'd4, 27'h000001bb, 5'd12, 27'h000002f2, 5'd2, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000354, 5'd10, 27'h00000158, 5'd14, 27'h00000008, 32'h00000400,
  1'd1,  5'd4, 27'h0000038d, 5'd14, 27'h00000100, 5'd21, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001d9, 5'd25, 27'h00000047, 5'd0, 27'h000003cd, 32'h00000400,
  1'd1,  5'd4, 27'h000003f2, 5'd21, 27'h00000353, 5'd10, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000023b, 5'd24, 27'h000003cb, 5'd24, 27'h000002b5, 32'h00000400,
  1'd1,  5'd11, 27'h000002b6, 5'd2, 27'h00000187, 5'd0, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002fe, 5'd1, 27'h00000027, 5'd11, 27'h000003e9, 32'h00000400,
  1'd1,  5'd15, 27'h00000095, 5'd3, 27'h00000269, 5'd25, 27'h00000144, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003f1, 5'd14, 27'h000003fb, 5'd3, 27'h000000bd, 32'h00000400,
  1'd1,  5'd11, 27'h0000019c, 5'd14, 27'h0000015d, 5'd10, 27'h0000028f, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000012b, 5'd14, 27'h00000126, 5'd21, 27'h00000350, 32'h00000400,
  1'd1,  5'd12, 27'h00000319, 5'd25, 27'h000000ce, 5'd1, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000a1, 5'd25, 27'h00000333, 5'd13, 27'h000001e5, 32'h00000400,
  1'd1,  5'd14, 27'h00000103, 5'd22, 27'h0000009a, 5'd21, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000346, 5'd4, 27'h00000222, 5'd3, 27'h000000a9, 32'h00000400,
  1'd1,  5'd21, 27'h000002e9, 5'd3, 27'h0000020c, 5'd14, 27'h000001a5, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000044, 5'd4, 27'h00000292, 5'd25, 27'h00000335, 32'h00000400,
  1'd1,  5'd24, 27'h00000267, 5'd11, 27'h00000293, 5'd4, 27'h000001a2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000335, 5'd14, 27'h000002f9, 5'd11, 27'h0000002d, 32'h00000400,
  1'd1,  5'd22, 27'h0000003c, 5'd11, 27'h0000039c, 5'd24, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000344, 5'd24, 27'h00000379, 5'd1, 27'h0000011d, 32'h00000400,
  1'd1,  5'd25, 27'h00000315, 5'd20, 27'h000002f1, 5'd14, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003d0, 5'd25, 27'h00000164, 5'd23, 27'h0000036d, 32'h00000400,
  1'd1,  5'd3, 27'h00000040, 5'd3, 27'h000002b1, 5'd7, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001d5, 5'd4, 27'h00000186, 5'd19, 27'h000002a4, 32'h00000400,
  1'd1,  5'd2, 27'h0000030f, 5'd4, 27'h000003d6, 5'd27, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd4, 27'h000000a9, 5'd11, 27'h00000076, 5'd7, 27'h00000089, 32'h00000400,
  1'd1,  5'd0, 27'h000000f3, 5'd12, 27'h000000c7, 5'd19, 27'h00000188, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000001c, 5'd13, 27'h000000f1, 5'd29, 27'h00000102, 32'h00000400,
  1'd1,  5'd0, 27'h000001e4, 5'd21, 27'h0000024d, 5'd7, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000012a, 5'd21, 27'h00000051, 5'd20, 27'h0000018e, 32'h00000400,
  1'd1,  5'd3, 27'h0000021c, 5'd20, 27'h00000358, 5'd28, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000026d, 5'd1, 27'h000003b5, 5'd5, 27'h00000195, 32'h00000400,
  1'd1,  5'd11, 27'h00000290, 5'd2, 27'h000002c6, 5'd19, 27'h000000bd, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001fa, 5'd2, 27'h00000197, 5'd28, 27'h0000005a, 32'h00000400,
  1'd1,  5'd12, 27'h00000361, 5'd12, 27'h00000343, 5'd10, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001c9, 5'd12, 27'h00000371, 5'd20, 27'h0000026a, 32'h00000400,
  1'd1,  5'd13, 27'h000002e6, 5'd14, 27'h000003d5, 5'd27, 27'h0000030e, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000d4, 5'd21, 27'h00000060, 5'd9, 27'h0000009e, 32'h00000400,
  1'd1,  5'd13, 27'h00000380, 5'd25, 27'h00000039, 5'd16, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000001, 5'd23, 27'h00000125, 5'd26, 27'h000003b2, 32'h00000400,
  1'd1,  5'd23, 27'h00000178, 5'd1, 27'h000002dc, 5'd9, 27'h000002a8, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000170, 5'd0, 27'h0000033e, 5'd20, 27'h0000012e, 32'h00000400,
  1'd1,  5'd24, 27'h00000277, 5'd4, 27'h00000122, 5'd27, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000031e, 5'd13, 27'h0000008f, 5'd8, 27'h00000131, 32'h00000400,
  1'd1,  5'd23, 27'h000003de, 5'd10, 27'h000003fa, 5'd16, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001e7, 5'd12, 27'h0000011c, 5'd27, 27'h000003ca, 32'h00000400,
  1'd1,  5'd23, 27'h000003c0, 5'd23, 27'h0000029c, 5'd8, 27'h0000016a, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000021b, 5'd21, 27'h000003aa, 5'd15, 27'h00000332, 32'h00000400,
  1'd1,  5'd23, 27'h000001d6, 5'd23, 27'h000000e1, 5'd29, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000119, 5'd7, 27'h000001d7, 5'd1, 27'h00000199, 32'h00000400,
  1'd1,  5'd4, 27'h00000399, 5'd8, 27'h00000289, 5'd14, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036b, 5'd8, 27'h000003d4, 5'd23, 27'h00000067, 32'h00000400,
  1'd1,  5'd0, 27'h0000030f, 5'd19, 27'h0000019a, 5'd2, 27'h000000cc, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000268, 5'd17, 27'h00000384, 5'd12, 27'h0000012d, 32'h00000400,
  1'd1,  5'd0, 27'h000000c0, 5'd17, 27'h000000c4, 5'd21, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f6, 5'd29, 27'h000002ee, 5'd3, 27'h000000b3, 32'h00000400,
  1'd1,  5'd2, 27'h00000012, 5'd27, 27'h00000258, 5'd14, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002d4, 5'd27, 27'h000002ed, 5'd20, 27'h000002e4, 32'h00000400,
  1'd1,  5'd14, 27'h00000182, 5'd9, 27'h000003fe, 5'd0, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002d1, 5'd6, 27'h0000034d, 5'd10, 27'h0000017e, 32'h00000400,
  1'd1,  5'd12, 27'h00000300, 5'd6, 27'h00000060, 5'd24, 27'h0000036a, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001d7, 5'd20, 27'h000000e9, 5'd0, 27'h00000088, 32'h00000400,
  1'd1,  5'd14, 27'h00000109, 5'd17, 27'h00000342, 5'd11, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002f1, 5'd18, 27'h00000287, 5'd20, 27'h000003b9, 32'h00000400,
  1'd1,  5'd13, 27'h000001a3, 5'd26, 27'h00000333, 5'd0, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000026, 5'd27, 27'h000001f5, 5'd11, 27'h00000348, 32'h00000400,
  1'd1,  5'd15, 27'h000001cf, 5'd26, 27'h00000228, 5'd20, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000170, 5'd5, 27'h00000152, 5'd2, 27'h000001b4, 32'h00000400,
  1'd1,  5'd23, 27'h00000050, 5'd9, 27'h00000235, 5'd14, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000068, 5'd18, 27'h000000e1, 5'd0, 27'h00000099, 32'h00000400,
  1'd1,  5'd23, 27'h000000b6, 5'd15, 27'h00000230, 5'd11, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000117, 5'd19, 27'h00000019, 5'd22, 27'h000001cc, 32'h00000400,
  1'd1,  5'd25, 27'h00000351, 5'd27, 27'h000002ab, 5'd0, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000381, 5'd30, 27'h00000292, 5'd15, 27'h0000017d, 32'h00000400,
  1'd1,  5'd20, 27'h0000036b, 5'd28, 27'h0000032e, 5'd25, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000008f, 5'd6, 27'h000000cf, 5'd7, 27'h0000034c, 32'h00000400,
  1'd1,  5'd3, 27'h000000b7, 5'd7, 27'h00000317, 5'd19, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000355, 5'd9, 27'h00000073, 5'd26, 27'h0000008e, 32'h00000400,
  1'd1,  5'd3, 27'h00000098, 5'd19, 27'h00000059, 5'd8, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000049, 5'd17, 27'h0000013f, 5'd17, 27'h00000074, 32'h00000400,
  1'd1,  5'd2, 27'h0000033c, 5'd19, 27'h00000321, 5'd29, 27'h000000e0, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000021c, 5'd30, 27'h0000025f, 5'd5, 27'h0000020e, 32'h00000400,
  1'd1,  5'd1, 27'h000002c3, 5'd27, 27'h00000047, 5'd16, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003fa, 5'd29, 27'h000000ed, 5'd27, 27'h00000033, 32'h00000400,
  1'd1,  5'd12, 27'h000003e3, 5'd8, 27'h0000017c, 5'd6, 27'h000003d7, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000010e, 5'd6, 27'h0000010f, 5'd17, 27'h0000017a, 32'h00000400,
  1'd1,  5'd13, 27'h0000011e, 5'd7, 27'h0000005e, 5'd26, 27'h000000bc, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000012c, 5'd18, 27'h000000b8, 5'd8, 27'h00000209, 32'h00000400,
  1'd1,  5'd10, 27'h00000345, 5'd20, 27'h0000018b, 5'd18, 27'h00000185, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000174, 5'd17, 27'h000001f5, 5'd28, 27'h00000388, 32'h00000400,
  1'd1,  5'd13, 27'h000001d0, 5'd29, 27'h000003e9, 5'd6, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001ea, 5'd28, 27'h00000047, 5'd16, 27'h0000008b, 32'h00000400,
  1'd1,  5'd10, 27'h000001c4, 5'd29, 27'h000002b5, 5'd30, 27'h000002cc, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000384, 5'd6, 27'h00000376, 5'd6, 27'h0000001a, 32'h00000400,
  1'd1,  5'd23, 27'h0000031b, 5'd9, 27'h000001d1, 5'd19, 27'h0000005a, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000016, 5'd8, 27'h000002e2, 5'd30, 27'h0000039d, 32'h00000400,
  1'd1,  5'd24, 27'h00000237, 5'd17, 27'h0000009c, 5'd9, 27'h000002e2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002f6, 5'd19, 27'h000000fb, 5'd15, 27'h0000032c, 32'h00000400,
  1'd1,  5'd24, 27'h0000039a, 5'd15, 27'h0000024f, 5'd28, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002aa, 5'd30, 27'h00000080, 5'd7, 27'h00000148, 32'h00000400,
  1'd1,  5'd20, 27'h00000380, 5'd27, 27'h0000029b, 5'd19, 27'h0000023b, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002e2, 5'd29, 27'h00000232, 5'd29, 27'h000001b1, 32'h00000400,
  1'd1,  5'd6, 27'h00000337, 5'd1, 27'h00000392, 5'd9, 27'h00000213, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000c8, 5'd3, 27'h000001c3, 5'd18, 27'h00000148, 32'h00000400,
  1'd1,  5'd9, 27'h0000038f, 5'd2, 27'h0000038c, 5'd27, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000010c, 5'd11, 27'h00000077, 5'd2, 27'h0000000d, 32'h00000400,
  1'd1,  5'd5, 27'h000001d4, 5'd13, 27'h00000094, 5'd14, 27'h00000388, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000284, 5'd12, 27'h000001b3, 5'd22, 27'h0000022b, 32'h00000400,
  1'd1,  5'd5, 27'h000001a0, 5'd24, 27'h000001a6, 5'd2, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000f7, 5'd25, 27'h0000034c, 5'd10, 27'h00000175, 32'h00000400,
  1'd1,  5'd9, 27'h000003cc, 5'd21, 27'h00000165, 5'd22, 27'h00000018, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001a6, 5'd0, 27'h00000371, 5'd7, 27'h00000140, 32'h00000400,
  1'd1,  5'd18, 27'h00000350, 5'd3, 27'h000001c6, 5'd19, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000019d, 5'd0, 27'h000003f4, 5'd29, 27'h0000002c, 32'h00000400,
  1'd1,  5'd16, 27'h0000022d, 5'd10, 27'h000002a9, 5'd0, 27'h000001c9, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039e, 5'd11, 27'h000003e3, 5'd12, 27'h00000264, 32'h00000400,
  1'd1,  5'd20, 27'h00000107, 5'd14, 27'h0000032a, 5'd23, 27'h00000067, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000193, 5'd21, 27'h0000020d, 5'd4, 27'h0000021d, 32'h00000400,
  1'd1,  5'd18, 27'h00000117, 5'd23, 27'h00000221, 5'd10, 27'h000003f4, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000027c, 5'd25, 27'h00000012, 5'd23, 27'h00000292, 32'h00000400,
  1'd1,  5'd29, 27'h0000008b, 5'd1, 27'h000003ec, 5'd1, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000041, 5'd0, 27'h00000361, 5'd10, 27'h000002bf, 32'h00000400,
  1'd1,  5'd30, 27'h00000075, 5'd3, 27'h000000cd, 5'd22, 27'h0000039e, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000089, 5'd13, 27'h00000248, 5'd4, 27'h00000127, 32'h00000400,
  1'd1,  5'd29, 27'h000000da, 5'd13, 27'h000002b5, 5'd14, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000364, 5'd12, 27'h0000017b, 5'd24, 27'h0000006b, 32'h00000400,
  1'd1,  5'd30, 27'h0000024a, 5'd24, 27'h000002f1, 5'd1, 27'h0000016c, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000001d, 5'd25, 27'h0000022f, 5'd14, 27'h000001a7, 32'h00000400,
  1'd1,  5'd30, 27'h000001e0, 5'd20, 27'h00000330, 5'd24, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001d1, 5'd1, 27'h00000093, 5'd5, 27'h00000035, 32'h00000400,
  1'd1,  5'd5, 27'h000003dd, 5'd0, 27'h00000126, 5'd10, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003d3, 5'd2, 27'h000002b0, 5'd25, 27'h000000d7, 32'h00000400,
  1'd1,  5'd8, 27'h000001ed, 5'd13, 27'h00000084, 5'd7, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000340, 5'd14, 27'h0000023d, 5'd20, 27'h00000203, 32'h00000400,
  1'd1,  5'd8, 27'h000003fe, 5'd10, 27'h000002e7, 5'd29, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000118, 5'd24, 27'h00000034, 5'd8, 27'h000001c9, 32'h00000400,
  1'd1,  5'd6, 27'h000001db, 5'd24, 27'h0000032a, 5'd19, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002a6, 5'd22, 27'h00000044, 5'd25, 27'h000003ac, 32'h00000400,
  1'd1,  5'd19, 27'h0000030e, 5'd1, 27'h000002d0, 5'd2, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000020a, 5'd1, 27'h000000f2, 5'd15, 27'h00000199, 32'h00000400,
  1'd1,  5'd16, 27'h00000186, 5'd13, 27'h00000086, 5'd9, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002ef, 5'd11, 27'h0000013b, 5'd19, 27'h000001e8, 32'h00000400,
  1'd1,  5'd18, 27'h00000297, 5'd13, 27'h0000028d, 5'd29, 27'h000002af, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003bb, 5'd24, 27'h000003a8, 5'd5, 27'h00000251, 32'h00000400,
  1'd1,  5'd19, 27'h0000034f, 5'd21, 27'h0000015d, 5'd19, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001c5, 5'd23, 27'h00000325, 5'd28, 27'h0000002f, 32'h00000400,
  1'd1,  5'd28, 27'h0000006b, 5'd0, 27'h00000020, 5'd6, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002cf, 5'd0, 27'h00000371, 5'd15, 27'h0000035f, 32'h00000400,
  1'd1,  5'd26, 27'h000000aa, 5'd0, 27'h000002a2, 5'd27, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000220, 5'd15, 27'h00000124, 5'd8, 27'h00000058, 32'h00000400,
  1'd1,  5'd27, 27'h00000125, 5'd11, 27'h0000000b, 5'd17, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000019d, 5'd14, 27'h0000032c, 5'd28, 27'h0000016e, 32'h00000400,
  1'd1,  5'd28, 27'h00000164, 5'd21, 27'h000001c3, 5'd5, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000316, 5'd21, 27'h000003f9, 5'd19, 27'h0000031b, 32'h00000400,
  1'd1,  5'd28, 27'h000000b2, 5'd24, 27'h0000002a, 5'd27, 27'h00000301, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000297, 5'd7, 27'h000000ef, 5'd4, 27'h00000219, 32'h00000400,
  1'd1,  5'd9, 27'h00000025, 5'd8, 27'h00000104, 5'd10, 27'h000003e8, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001d8, 5'd8, 27'h00000127, 5'd25, 27'h000002cf, 32'h00000400,
  1'd1,  5'd8, 27'h000001f8, 5'd17, 27'h0000010f, 5'd2, 27'h00000174, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000008d, 5'd20, 27'h000001c9, 5'd13, 27'h000002e0, 32'h00000400,
  1'd1,  5'd10, 27'h000000af, 5'd15, 27'h000002d7, 5'd22, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000214, 5'd27, 27'h000001ab, 5'd0, 27'h00000205, 32'h00000400,
  1'd1,  5'd9, 27'h0000013e, 5'd27, 27'h0000004f, 5'd11, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000376, 5'd25, 27'h000003aa, 5'd23, 27'h00000170, 32'h00000400,
  1'd1,  5'd20, 27'h0000002b, 5'd5, 27'h00000318, 5'd3, 27'h0000035c, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000020a, 5'd9, 27'h00000154, 5'd15, 27'h00000107, 32'h00000400,
  1'd1,  5'd18, 27'h0000032b, 5'd8, 27'h000003be, 5'd23, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002cf, 5'd15, 27'h00000313, 5'd4, 27'h00000393, 32'h00000400,
  1'd1,  5'd17, 27'h0000024a, 5'd20, 27'h00000142, 5'd12, 27'h0000018c, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000284, 5'd18, 27'h000001cc, 5'd25, 27'h0000017c, 32'h00000400,
  1'd1,  5'd17, 27'h000001be, 5'd27, 27'h0000021d, 5'd2, 27'h0000015d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000034e, 5'd30, 27'h00000174, 5'd12, 27'h00000173, 32'h00000400,
  1'd1,  5'd19, 27'h000001be, 5'd26, 27'h0000029f, 5'd22, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001de, 5'd10, 27'h00000026, 5'd4, 27'h000000b5, 32'h00000400,
  1'd1,  5'd26, 27'h00000276, 5'd6, 27'h00000302, 5'd12, 27'h0000033e, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001a6, 5'd9, 27'h0000026e, 5'd23, 27'h000000a1, 32'h00000400,
  1'd1,  5'd30, 27'h00000085, 5'd15, 27'h0000038f, 5'd4, 27'h000001b0, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000035a, 5'd19, 27'h00000252, 5'd13, 27'h000000ed, 32'h00000400,
  1'd1,  5'd25, 27'h00000376, 5'd17, 27'h000000f6, 5'd22, 27'h0000032b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000051, 5'd27, 27'h000001f0, 5'd3, 27'h000002d7, 32'h00000400,
  1'd1,  5'd30, 27'h00000386, 5'd25, 27'h0000036e, 5'd14, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000208, 5'd29, 27'h00000267, 5'd24, 27'h000000a8, 32'h00000400,
  1'd1,  5'd8, 27'h000000bc, 5'd10, 27'h00000035, 5'd5, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001f2, 5'd8, 27'h00000214, 5'd17, 27'h0000008a, 32'h00000400,
  1'd1,  5'd9, 27'h0000031e, 5'd7, 27'h00000323, 5'd30, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000295, 5'd18, 27'h00000353, 5'd9, 27'h000001a1, 32'h00000400,
  1'd1,  5'd7, 27'h0000032a, 5'd16, 27'h000003c3, 5'd20, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000196, 5'd18, 27'h0000013f, 5'd27, 27'h000000ba, 32'h00000400,
  1'd1,  5'd9, 27'h000000a6, 5'd27, 27'h000001d4, 5'd9, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001e8, 5'd29, 27'h00000246, 5'd16, 27'h000002fd, 32'h00000400,
  1'd1,  5'd10, 27'h00000112, 5'd30, 27'h00000111, 5'd28, 27'h00000380, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000002a, 5'd9, 27'h000002b6, 5'd9, 27'h000000c5, 32'h00000400,
  1'd1,  5'd17, 27'h00000255, 5'd6, 27'h000003f8, 5'd16, 27'h0000008a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002a6, 5'd8, 27'h00000080, 5'd29, 27'h0000002c, 32'h00000400,
  1'd1,  5'd16, 27'h0000031e, 5'd16, 27'h000003d7, 5'd8, 27'h0000002b, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000292, 5'd18, 27'h000001af, 5'd19, 27'h0000009b, 32'h00000400,
  1'd1,  5'd18, 27'h00000275, 5'd19, 27'h000002a7, 5'd30, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000010, 5'd29, 27'h00000112, 5'd8, 27'h0000019e, 32'h00000400,
  1'd1,  5'd15, 27'h00000340, 5'd26, 27'h00000065, 5'd19, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003dc, 5'd27, 27'h000001ea, 5'd29, 27'h0000014c, 32'h00000400,
  1'd1,  5'd30, 27'h000000bd, 5'd8, 27'h00000017, 5'd10, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000012d, 5'd7, 27'h000001f4, 5'd17, 27'h000001ac, 32'h00000400,
  1'd1,  5'd29, 27'h00000234, 5'd5, 27'h0000010a, 5'd25, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000185, 5'd17, 27'h000003be, 5'd7, 27'h0000032d, 32'h00000400,
  1'd1,  5'd29, 27'h00000076, 5'd20, 27'h0000020d, 5'd17, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000012b, 5'd18, 27'h000002f5, 5'd30, 27'h0000033e, 32'h00000400,
  1'd1,  5'd28, 27'h000002da, 5'd28, 27'h00000230, 5'd7, 27'h00000255, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003e5, 5'd27, 27'h000000e6, 5'd20, 27'h00000137, 32'h00000400,
  1'd1,  5'd30, 27'h000000f0, 5'd30, 27'h00000245, 5'd28, 27'h00000298, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd1, 27'h000003b5, 5'd4, 27'h0000039d, 5'd4, 27'h0000005f, 32'h00000400,
  1'd1,  5'd0, 27'h00000106, 5'd2, 27'h00000337, 5'd11, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000002, 5'd3, 27'h0000017f, 5'd22, 27'h0000020b, 32'h00000400,
  1'd1,  5'd4, 27'h0000029d, 5'd14, 27'h00000233, 5'd1, 27'h000000e9, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000034f, 5'd12, 27'h000003e9, 5'd10, 27'h000002f0, 32'h00000400,
  1'd1,  5'd0, 27'h000001c9, 5'd12, 27'h000001c0, 5'd21, 27'h000003b4, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000ec, 5'd22, 27'h000002e5, 5'd4, 27'h000002d4, 32'h00000400,
  1'd1,  5'd3, 27'h0000018b, 5'd21, 27'h000002ec, 5'd11, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000022, 5'd23, 27'h0000014c, 5'd22, 27'h0000031d, 32'h00000400,
  1'd1,  5'd10, 27'h00000191, 5'd1, 27'h000002f5, 5'd1, 27'h00000250, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000161, 5'd4, 27'h000002a7, 5'd12, 27'h00000054, 32'h00000400,
  1'd1,  5'd12, 27'h0000036d, 5'd1, 27'h00000201, 5'd25, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000200, 5'd13, 27'h00000065, 5'd1, 27'h000001c5, 32'h00000400,
  1'd1,  5'd10, 27'h00000276, 5'd14, 27'h00000391, 5'd11, 27'h0000028b, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000156, 5'd12, 27'h000001c9, 5'd22, 27'h000000cd, 32'h00000400,
  1'd1,  5'd13, 27'h000003bb, 5'd22, 27'h00000111, 5'd0, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000005b, 5'd24, 27'h00000138, 5'd10, 27'h000001a9, 32'h00000400,
  1'd1,  5'd12, 27'h0000023f, 5'd23, 27'h000001e2, 5'd24, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000004, 5'd4, 27'h000000fb, 5'd4, 27'h000002ed, 32'h00000400,
  1'd1,  5'd23, 27'h0000004e, 5'd2, 27'h00000335, 5'd13, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000021b, 5'd1, 27'h000000cc, 5'd24, 27'h0000028e, 32'h00000400,
  1'd1,  5'd22, 27'h00000193, 5'd11, 27'h0000033f, 5'd1, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003cf, 5'd13, 27'h0000024e, 5'd15, 27'h000000d1, 32'h00000400,
  1'd1,  5'd25, 27'h000002c5, 5'd14, 27'h000002a8, 5'd24, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003b0, 5'd22, 27'h000000ff, 5'd4, 27'h000003e6, 32'h00000400,
  1'd1,  5'd21, 27'h00000388, 5'd22, 27'h000003f6, 5'd11, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000e6, 5'd25, 27'h0000028e, 5'd23, 27'h00000147, 32'h00000400,
  1'd1,  5'd3, 27'h000003cc, 5'd0, 27'h00000398, 5'd5, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000033f, 5'd0, 27'h00000341, 5'd18, 27'h0000024b, 32'h00000400,
  1'd1,  5'd4, 27'h000000d8, 5'd3, 27'h00000086, 5'd28, 27'h0000018d, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000002c, 5'd13, 27'h000000db, 5'd5, 27'h00000279, 32'h00000400,
  1'd1,  5'd2, 27'h000002d2, 5'd14, 27'h00000226, 5'd18, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000027c, 5'd13, 27'h000001a2, 5'd29, 27'h000003a4, 32'h00000400,
  1'd1,  5'd3, 27'h00000026, 5'd23, 27'h00000075, 5'd5, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000e4, 5'd24, 27'h000003c4, 5'd19, 27'h0000012f, 32'h00000400,
  1'd1,  5'd4, 27'h000000c2, 5'd24, 27'h0000020f, 5'd28, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002e6, 5'd1, 27'h00000202, 5'd9, 27'h000000a1, 32'h00000400,
  1'd1,  5'd15, 27'h000000d1, 5'd3, 27'h0000021a, 5'd15, 27'h000002e7, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001b6, 5'd2, 27'h00000241, 5'd27, 27'h00000047, 32'h00000400,
  1'd1,  5'd13, 27'h00000035, 5'd11, 27'h000003ff, 5'd7, 27'h000002f4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000163, 5'd12, 27'h000000ff, 5'd16, 27'h000003e8, 32'h00000400,
  1'd1,  5'd13, 27'h000000d4, 5'd14, 27'h00000086, 5'd30, 27'h00000315, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003de, 5'd25, 27'h00000146, 5'd8, 27'h000003a9, 32'h00000400,
  1'd1,  5'd12, 27'h00000080, 5'd21, 27'h00000184, 5'd18, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000241, 5'd24, 27'h0000025e, 5'd27, 27'h000003d1, 32'h00000400,
  1'd1,  5'd25, 27'h0000026b, 5'd2, 27'h0000031d, 5'd9, 27'h00000171, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000273, 5'd5, 27'h00000081, 5'd19, 27'h000000c7, 32'h00000400,
  1'd1,  5'd24, 27'h000002ec, 5'd2, 27'h0000030c, 5'd29, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000350, 5'd13, 27'h000003b7, 5'd5, 27'h000003a4, 32'h00000400,
  1'd1,  5'd24, 27'h0000026a, 5'd14, 27'h00000379, 5'd16, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000295, 5'd11, 27'h00000243, 5'd28, 27'h000002c8, 32'h00000400,
  1'd1,  5'd25, 27'h0000017a, 5'd25, 27'h000002fd, 5'd8, 27'h00000348, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003ca, 5'd23, 27'h00000166, 5'd20, 27'h000001cb, 32'h00000400,
  1'd1,  5'd25, 27'h00000270, 5'd22, 27'h000003d1, 5'd26, 27'h000000a7, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003ee, 5'd5, 27'h000002a0, 5'd2, 27'h00000144, 32'h00000400,
  1'd1,  5'd1, 27'h000000b1, 5'd6, 27'h000002fc, 5'd10, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000226, 5'd7, 27'h00000295, 5'd22, 27'h000002ae, 32'h00000400,
  1'd1,  5'd3, 27'h000001a8, 5'd15, 27'h0000035e, 5'd3, 27'h00000049, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000253, 5'd18, 27'h0000005b, 5'd15, 27'h000000c2, 32'h00000400,
  1'd1,  5'd0, 27'h000000d9, 5'd19, 27'h000000b7, 5'd20, 27'h0000036b, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000003f, 5'd30, 27'h0000001a, 5'd2, 27'h0000006f, 32'h00000400,
  1'd1,  5'd3, 27'h00000224, 5'd27, 27'h000001e8, 5'd14, 27'h00000253, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038f, 5'd30, 27'h0000011f, 5'd21, 27'h0000003f, 32'h00000400,
  1'd1,  5'd11, 27'h00000206, 5'd5, 27'h00000116, 5'd3, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000023b, 5'd9, 27'h00000244, 5'd13, 27'h00000337, 32'h00000400,
  1'd1,  5'd13, 27'h000001cf, 5'd5, 27'h0000036c, 5'd22, 27'h00000109, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000301, 5'd19, 27'h000001be, 5'd2, 27'h000001d5, 32'h00000400,
  1'd1,  5'd10, 27'h00000350, 5'd18, 27'h0000034b, 5'd15, 27'h000001a6, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000382, 5'd18, 27'h0000037e, 5'd25, 27'h0000005d, 32'h00000400,
  1'd1,  5'd13, 27'h00000331, 5'd27, 27'h00000197, 5'd3, 27'h0000012d, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000094, 5'd28, 27'h000001f2, 5'd10, 27'h0000022d, 32'h00000400,
  1'd1,  5'd14, 27'h000001f0, 5'd26, 27'h000001ac, 5'd25, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000215, 5'd5, 27'h000003e1, 5'd4, 27'h000002e0, 32'h00000400,
  1'd1,  5'd24, 27'h0000039f, 5'd7, 27'h00000244, 5'd13, 27'h00000398, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000036b, 5'd16, 27'h000002c2, 5'd1, 27'h0000008e, 32'h00000400,
  1'd1,  5'd22, 27'h00000373, 5'd18, 27'h000003f7, 5'd13, 27'h0000023a, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002ce, 5'd16, 27'h000001b0, 5'd22, 27'h0000021a, 32'h00000400,
  1'd1,  5'd23, 27'h00000384, 5'd26, 27'h0000009c, 5'd1, 27'h00000010, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003a0, 5'd27, 27'h0000004f, 5'd12, 27'h00000184, 32'h00000400,
  1'd1,  5'd24, 27'h000001a8, 5'd26, 27'h000003d5, 5'd24, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000345, 5'd6, 27'h00000006, 5'd7, 27'h00000272, 32'h00000400,
  1'd1,  5'd2, 27'h000002d8, 5'd5, 27'h000002d1, 5'd18, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000003b, 5'd6, 27'h0000020b, 5'd27, 27'h000001f3, 32'h00000400,
  1'd1,  5'd3, 27'h000003aa, 5'd15, 27'h00000219, 5'd5, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000025, 5'd15, 27'h00000247, 5'd16, 27'h0000010d, 32'h00000400,
  1'd1,  5'd2, 27'h00000130, 5'd16, 27'h000001c7, 5'd29, 27'h000002da, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000c6, 5'd26, 27'h0000002e, 5'd8, 27'h0000020d, 32'h00000400,
  1'd1,  5'd3, 27'h0000008a, 5'd28, 27'h0000011d, 5'd18, 27'h00000142, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000029c, 5'd30, 27'h00000272, 5'd30, 27'h000003ce, 32'h00000400,
  1'd1,  5'd12, 27'h0000019f, 5'd10, 27'h00000052, 5'd10, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000333, 5'd7, 27'h0000016e, 5'd20, 27'h000000b2, 32'h00000400,
  1'd1,  5'd11, 27'h00000034, 5'd7, 27'h00000336, 5'd27, 27'h000000af, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000149, 5'd18, 27'h00000353, 5'd9, 27'h00000169, 32'h00000400,
  1'd1,  5'd14, 27'h0000023d, 5'd19, 27'h00000038, 5'd20, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000018d, 5'd16, 27'h00000082, 5'd28, 27'h0000031b, 32'h00000400,
  1'd1,  5'd13, 27'h0000008b, 5'd26, 27'h00000097, 5'd6, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001f7, 5'd26, 27'h00000073, 5'd17, 27'h00000364, 32'h00000400,
  1'd1,  5'd10, 27'h00000300, 5'd30, 27'h00000344, 5'd30, 27'h00000089, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000356, 5'd10, 27'h00000024, 5'd5, 27'h0000016c, 32'h00000400,
  1'd1,  5'd21, 27'h000003fa, 5'd7, 27'h00000030, 5'd16, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002d3, 5'd6, 27'h000003fe, 5'd26, 27'h0000017b, 32'h00000400,
  1'd1,  5'd24, 27'h000000ee, 5'd16, 27'h00000396, 5'd9, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000041, 5'd16, 27'h00000348, 5'd15, 27'h000003f2, 32'h00000400,
  1'd1,  5'd24, 27'h00000033, 5'd17, 27'h000003bf, 5'd28, 27'h000000ce, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000322, 5'd28, 27'h00000031, 5'd8, 27'h000002ec, 32'h00000400,
  1'd1,  5'd21, 27'h00000174, 5'd30, 27'h0000002a, 5'd17, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000058, 5'd29, 27'h00000073, 5'd26, 27'h000002b6, 32'h00000400,
  1'd1,  5'd6, 27'h0000032d, 5'd1, 27'h000001f9, 5'd8, 27'h00000332, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000277, 5'd3, 27'h00000027, 5'd19, 27'h00000237, 32'h00000400,
  1'd1,  5'd9, 27'h000002d5, 5'd2, 27'h000003f5, 5'd30, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000e8, 5'd11, 27'h00000287, 5'd3, 27'h000001bf, 32'h00000400,
  1'd1,  5'd5, 27'h0000031d, 5'd13, 27'h00000256, 5'd15, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000127, 5'd14, 27'h00000122, 5'd21, 27'h000002c4, 32'h00000400,
  1'd1,  5'd8, 27'h000000c5, 5'd25, 27'h0000029f, 5'd0, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003f1, 5'd22, 27'h00000127, 5'd11, 27'h000002f9, 32'h00000400,
  1'd1,  5'd9, 27'h00000067, 5'd24, 27'h000002b8, 5'd23, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003af, 5'd2, 27'h0000001d, 5'd5, 27'h00000298, 32'h00000400,
  1'd1,  5'd17, 27'h0000007a, 5'd4, 27'h00000017, 5'd16, 27'h00000361, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000000d, 5'd3, 27'h00000395, 5'd26, 27'h000002e3, 32'h00000400,
  1'd1,  5'd18, 27'h00000123, 5'd14, 27'h00000180, 5'd3, 27'h0000000d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000013b, 5'd11, 27'h00000097, 5'd13, 27'h00000068, 32'h00000400,
  1'd1,  5'd19, 27'h00000095, 5'd15, 27'h00000080, 5'd22, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000387, 5'd21, 27'h000003f2, 5'd1, 27'h000000ee, 32'h00000400,
  1'd1,  5'd17, 27'h000002d1, 5'd24, 27'h00000336, 5'd10, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000011c, 5'd23, 27'h0000017a, 5'd25, 27'h0000032d, 32'h00000400,
  1'd1,  5'd28, 27'h00000029, 5'd2, 27'h000000e9, 5'd3, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000158, 5'd4, 27'h0000029a, 5'd11, 27'h00000166, 32'h00000400,
  1'd1,  5'd26, 27'h000001c9, 5'd4, 27'h000000a6, 5'd22, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000237, 5'd14, 27'h00000378, 5'd4, 27'h000002dc, 32'h00000400,
  1'd1,  5'd27, 27'h00000087, 5'd13, 27'h00000167, 5'd13, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000347, 5'd15, 27'h00000198, 5'd23, 27'h0000015b, 32'h00000400,
  1'd1,  5'd28, 27'h0000003d, 5'd21, 27'h000003fb, 5'd0, 27'h0000037e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000019c, 5'd22, 27'h00000105, 5'd13, 27'h00000185, 32'h00000400,
  1'd1,  5'd29, 27'h0000026f, 5'd25, 27'h000000dd, 5'd25, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000000a, 5'd1, 27'h000003e6, 5'd1, 27'h00000086, 32'h00000400,
  1'd1,  5'd8, 27'h00000022, 5'd2, 27'h0000038f, 5'd11, 27'h00000310, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002db, 5'd3, 27'h00000088, 5'd24, 27'h00000100, 32'h00000400,
  1'd1,  5'd10, 27'h00000082, 5'd13, 27'h0000037d, 5'd5, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000001d, 5'd12, 27'h000000f0, 5'd20, 27'h000001f5, 32'h00000400,
  1'd1,  5'd5, 27'h000000fc, 5'd12, 27'h00000111, 5'd26, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000187, 5'd25, 27'h0000015e, 5'd10, 27'h00000094, 32'h00000400,
  1'd1,  5'd9, 27'h000001fe, 5'd22, 27'h00000086, 5'd19, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021b, 5'd23, 27'h000001ef, 5'd30, 27'h0000032a, 32'h00000400,
  1'd1,  5'd19, 27'h000001d0, 5'd1, 27'h0000025e, 5'd4, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003e1, 5'd1, 27'h00000365, 5'd15, 27'h000001c4, 32'h00000400,
  1'd1,  5'd20, 27'h0000029f, 5'd10, 27'h000002c7, 5'd9, 27'h0000029a, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000087, 5'd13, 27'h00000121, 5'd16, 27'h000002d6, 32'h00000400,
  1'd1,  5'd18, 27'h0000034d, 5'd13, 27'h000000a3, 5'd27, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003ca, 5'd23, 27'h000001e7, 5'd6, 27'h000001d3, 32'h00000400,
  1'd1,  5'd17, 27'h00000385, 5'd25, 27'h0000009b, 5'd17, 27'h00000243, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001fb, 5'd23, 27'h00000310, 5'd26, 27'h00000337, 32'h00000400,
  1'd1,  5'd27, 27'h00000131, 5'd0, 27'h0000007b, 5'd6, 27'h0000028e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e9, 5'd1, 27'h000002ad, 5'd16, 27'h00000078, 32'h00000400,
  1'd1,  5'd28, 27'h000000a5, 5'd2, 27'h0000035a, 5'd29, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000017e, 5'd12, 27'h000002ae, 5'd7, 27'h000003bf, 32'h00000400,
  1'd1,  5'd28, 27'h00000312, 5'd10, 27'h000001f1, 5'd18, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000309, 5'd10, 27'h00000221, 5'd29, 27'h0000029e, 32'h00000400,
  1'd1,  5'd27, 27'h0000023c, 5'd22, 27'h000003bd, 5'd7, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000282, 5'd23, 27'h000002bf, 5'd20, 27'h00000093, 32'h00000400,
  1'd1,  5'd27, 27'h00000200, 5'd23, 27'h0000000f, 5'd29, 27'h000001fe, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011c, 5'd9, 27'h0000006b, 5'd2, 27'h00000143, 32'h00000400,
  1'd1,  5'd10, 27'h0000001a, 5'd6, 27'h000001b0, 5'd13, 27'h0000014f, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003f2, 5'd8, 27'h00000317, 5'd23, 27'h00000347, 32'h00000400,
  1'd1,  5'd10, 27'h000000bd, 5'd17, 27'h000003eb, 5'd3, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000105, 5'd20, 27'h000000c1, 5'd13, 27'h0000038a, 32'h00000400,
  1'd1,  5'd7, 27'h0000036a, 5'd16, 27'h00000204, 5'd24, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000025a, 5'd29, 27'h0000014e, 5'd2, 27'h00000013, 32'h00000400,
  1'd1,  5'd7, 27'h0000039f, 5'd27, 27'h000001ac, 5'd11, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000003b, 5'd30, 27'h000003a5, 5'd23, 27'h00000326, 32'h00000400,
  1'd1,  5'd18, 27'h0000010d, 5'd8, 27'h0000003e, 5'd1, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000015e, 5'd8, 27'h00000033, 5'd15, 27'h00000192, 32'h00000400,
  1'd1,  5'd16, 27'h000000c5, 5'd5, 27'h00000263, 5'd21, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000266, 5'd15, 27'h0000024b, 5'd4, 27'h00000347, 32'h00000400,
  1'd1,  5'd16, 27'h0000024c, 5'd19, 27'h000001d0, 5'd13, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002fe, 5'd18, 27'h00000008, 5'd22, 27'h000001ce, 32'h00000400,
  1'd1,  5'd18, 27'h000002d7, 5'd26, 27'h00000257, 5'd0, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001f2, 5'd26, 27'h000002c3, 5'd14, 27'h000000ea, 32'h00000400,
  1'd1,  5'd16, 27'h00000011, 5'd26, 27'h0000006e, 5'd23, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000017b, 5'd5, 27'h000000ae, 5'd2, 27'h0000008e, 32'h00000400,
  1'd1,  5'd30, 27'h000002ba, 5'd8, 27'h00000175, 5'd15, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000317, 5'd5, 27'h00000176, 5'd25, 27'h0000023a, 32'h00000400,
  1'd1,  5'd26, 27'h000000a6, 5'd19, 27'h000002cc, 5'd5, 27'h00000003, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000e8, 5'd15, 27'h0000026c, 5'd14, 27'h00000215, 32'h00000400,
  1'd1,  5'd30, 27'h00000242, 5'd16, 27'h000003d1, 5'd21, 27'h000000ca, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000285, 5'd27, 27'h0000015b, 5'd4, 27'h00000132, 32'h00000400,
  1'd1,  5'd29, 27'h00000264, 5'd30, 27'h000000c8, 5'd10, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e3, 5'd30, 27'h000001aa, 5'd25, 27'h00000165, 32'h00000400,
  1'd1,  5'd8, 27'h00000228, 5'd5, 27'h000003e7, 5'd9, 27'h0000029d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000091, 5'd8, 27'h000002e8, 5'd20, 27'h0000022b, 32'h00000400,
  1'd1,  5'd5, 27'h000000f1, 5'd8, 27'h000002f7, 5'd28, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000d9, 5'd20, 27'h000001ee, 5'd7, 27'h00000290, 32'h00000400,
  1'd1,  5'd9, 27'h0000014d, 5'd18, 27'h000003fa, 5'd17, 27'h0000017b, 32'hfffffc00,
  1'd1,  5'd7, 27'h000003a5, 5'd19, 27'h00000181, 5'd26, 27'h00000034, 32'h00000400,
  1'd1,  5'd7, 27'h00000376, 5'd30, 27'h00000157, 5'd5, 27'h00000374, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000030e, 5'd27, 27'h000003fb, 5'd16, 27'h00000024, 32'h00000400,
  1'd1,  5'd5, 27'h000001b4, 5'd29, 27'h000002aa, 5'd29, 27'h000000b1, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001dc, 5'd7, 27'h0000016a, 5'd9, 27'h000000c8, 32'h00000400,
  1'd1,  5'd18, 27'h000002ac, 5'd10, 27'h00000085, 5'd16, 27'h00000218, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003c4, 5'd8, 27'h0000008b, 5'd26, 27'h00000014, 32'h00000400,
  1'd1,  5'd16, 27'h00000272, 5'd20, 27'h00000257, 5'd5, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000139, 5'd19, 27'h0000008e, 5'd16, 27'h000000c9, 32'h00000400,
  1'd1,  5'd18, 27'h000000b0, 5'd18, 27'h00000044, 5'd26, 27'h0000011f, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000397, 5'd29, 27'h000000ff, 5'd6, 27'h0000017e, 32'h00000400,
  1'd1,  5'd19, 27'h000002dd, 5'd28, 27'h000000d6, 5'd17, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000098, 5'd30, 27'h000000c4, 5'd28, 27'h0000015a, 32'h00000400,
  1'd1,  5'd30, 27'h00000328, 5'd8, 27'h000000e8, 5'd6, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000030a, 5'd6, 27'h000000ce, 5'd20, 27'h00000212, 32'h00000400,
  1'd1,  5'd28, 27'h000003f8, 5'd6, 27'h00000272, 5'd26, 27'h0000003d, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001bc, 5'd17, 27'h000002db, 5'd7, 27'h0000022a, 32'h00000400,
  1'd1,  5'd26, 27'h000000e2, 5'd17, 27'h0000017b, 5'd18, 27'h000002c6, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000008d, 5'd20, 27'h00000222, 5'd27, 27'h000000d8, 32'h00000400,
  1'd1,  5'd29, 27'h000000d1, 5'd27, 27'h00000152, 5'd6, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000bc, 5'd26, 27'h000002cf, 5'd16, 27'h00000349, 32'h00000400,
  1'd1,  5'd30, 27'h000003a6, 5'd27, 27'h000002be, 5'd28, 27'h00000239, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000031b, 5'd4, 27'h0000034a, 5'd4, 27'h000002ea, 32'h00000400,
  1'd1,  5'd0, 27'h0000009e, 5'd0, 27'h000001bd, 5'd14, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000006a, 5'd1, 27'h0000009d, 5'd20, 27'h00000300, 32'h00000400,
  1'd1,  5'd0, 27'h000001b6, 5'd13, 27'h000003f0, 5'd1, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002ba, 5'd13, 27'h0000034f, 5'd10, 27'h00000323, 32'h00000400,
  1'd1,  5'd1, 27'h000002ea, 5'd12, 27'h0000034a, 5'd23, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001d6, 5'd20, 27'h000003c0, 5'd0, 27'h0000039b, 32'h00000400,
  1'd1,  5'd1, 27'h0000027e, 5'd20, 27'h00000338, 5'd10, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000036a, 5'd24, 27'h000001ab, 5'd25, 27'h000000de, 32'h00000400,
  1'd1,  5'd10, 27'h00000220, 5'd1, 27'h00000335, 5'd4, 27'h0000036e, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000276, 5'd4, 27'h0000007a, 5'd13, 27'h000002a0, 32'h00000400,
  1'd1,  5'd15, 27'h0000011b, 5'd1, 27'h000003dd, 5'd22, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000223, 5'd13, 27'h000000c3, 5'd1, 27'h000003e7, 32'h00000400,
  1'd1,  5'd11, 27'h000001b8, 5'd12, 27'h0000028b, 5'd11, 27'h0000010a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000206, 5'd13, 27'h000002f2, 5'd21, 27'h000000e7, 32'h00000400,
  1'd1,  5'd12, 27'h000002aa, 5'd24, 27'h00000388, 5'd4, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000282, 5'd23, 27'h000002fd, 5'd10, 27'h00000261, 32'h00000400,
  1'd1,  5'd15, 27'h000000a4, 5'd25, 27'h000002ed, 5'd25, 27'h00000145, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003f0, 5'd4, 27'h000000b0, 5'd4, 27'h0000009f, 32'h00000400,
  1'd1,  5'd24, 27'h000002cc, 5'd5, 27'h0000002b, 5'd11, 27'h000003b8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000082, 5'd3, 27'h0000027a, 5'd22, 27'h000002e0, 32'h00000400,
  1'd1,  5'd21, 27'h00000020, 5'd14, 27'h00000292, 5'd0, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000001c, 5'd10, 27'h000003f9, 5'd15, 27'h00000117, 32'h00000400,
  1'd1,  5'd25, 27'h0000009a, 5'd13, 27'h00000021, 5'd23, 27'h000000b6, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000010a, 5'd23, 27'h00000393, 5'd0, 27'h00000244, 32'h00000400,
  1'd1,  5'd25, 27'h00000163, 5'd22, 27'h000003c3, 5'd12, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002f1, 5'd22, 27'h00000266, 5'd24, 27'h000000cf, 32'h00000400,
  1'd1,  5'd1, 27'h0000030c, 5'd0, 27'h0000032f, 5'd5, 27'h0000039d, 32'hfffffc00,
  1'd1,  5'd1, 27'h000000df, 5'd3, 27'h0000009b, 5'd16, 27'h000002fd, 32'h00000400,
  1'd1,  5'd1, 27'h0000013b, 5'd4, 27'h0000007e, 5'd28, 27'h00000107, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001cb, 5'd13, 27'h00000127, 5'd5, 27'h000003ab, 32'h00000400,
  1'd1,  5'd4, 27'h0000038e, 5'd13, 27'h000001f6, 5'd16, 27'h00000245, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000287, 5'd12, 27'h00000045, 5'd29, 27'h00000010, 32'h00000400,
  1'd1,  5'd4, 27'h000000b1, 5'd24, 27'h00000237, 5'd8, 27'h000000dd, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000037c, 5'd23, 27'h000000e9, 5'd16, 27'h000003a2, 32'h00000400,
  1'd1,  5'd2, 27'h0000013c, 5'd24, 27'h000001f7, 5'd27, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000322, 5'd2, 27'h00000173, 5'd8, 27'h000002c1, 32'h00000400,
  1'd1,  5'd14, 27'h000003da, 5'd0, 27'h000002a7, 5'd17, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003da, 5'd2, 27'h00000213, 5'd28, 27'h000002a5, 32'h00000400,
  1'd1,  5'd13, 27'h0000002c, 5'd12, 27'h00000128, 5'd9, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000121, 5'd11, 27'h0000017c, 5'd16, 27'h0000023c, 32'h00000400,
  1'd1,  5'd14, 27'h0000014a, 5'd12, 27'h0000029a, 5'd26, 27'h000000f1, 32'hfffffc00,
  1'd1,  5'd14, 27'h000002f8, 5'd23, 27'h0000009d, 5'd6, 27'h0000001c, 32'h00000400,
  1'd1,  5'd10, 27'h000001b1, 5'd23, 27'h00000306, 5'd16, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003b3, 5'd21, 27'h00000059, 5'd26, 27'h0000000f, 32'h00000400,
  1'd1,  5'd23, 27'h000000b2, 5'd2, 27'h000003e6, 5'd10, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002bc, 5'd3, 27'h00000224, 5'd18, 27'h0000023b, 32'h00000400,
  1'd1,  5'd23, 27'h00000029, 5'd3, 27'h000001f2, 5'd30, 27'h00000074, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000028f, 5'd11, 27'h00000196, 5'd10, 27'h00000051, 32'h00000400,
  1'd1,  5'd23, 27'h000002f2, 5'd11, 27'h000003bc, 5'd19, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000028a, 5'd15, 27'h000001a0, 5'd26, 27'h00000075, 32'h00000400,
  1'd1,  5'd24, 27'h000003e2, 5'd23, 27'h000002b7, 5'd8, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003ee, 5'd22, 27'h0000029a, 5'd17, 27'h000000c8, 32'h00000400,
  1'd1,  5'd25, 27'h000002b9, 5'd20, 27'h000003d7, 5'd27, 27'h00000335, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000030d, 5'd5, 27'h00000375, 5'd4, 27'h0000003a, 32'h00000400,
  1'd1,  5'd2, 27'h000001fe, 5'd7, 27'h00000149, 5'd12, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000239, 5'd8, 27'h00000039, 5'd22, 27'h00000064, 32'h00000400,
  1'd1,  5'd5, 27'h00000072, 5'd16, 27'h00000269, 5'd3, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000214, 5'd18, 27'h000000d7, 5'd14, 27'h00000355, 32'h00000400,
  1'd1,  5'd4, 27'h000001df, 5'd19, 27'h0000008c, 5'd24, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000039e, 5'd29, 27'h000001ce, 5'd2, 27'h000000ad, 32'h00000400,
  1'd1,  5'd2, 27'h0000026a, 5'd30, 27'h00000261, 5'd11, 27'h00000068, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000096, 5'd28, 27'h0000035a, 5'd24, 27'h00000311, 32'h00000400,
  1'd1,  5'd13, 27'h0000037f, 5'd7, 27'h0000031b, 5'd2, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000014d, 5'd6, 27'h00000176, 5'd10, 27'h00000166, 32'h00000400,
  1'd1,  5'd13, 27'h0000039b, 5'd7, 27'h00000004, 5'd23, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000034e, 5'd18, 27'h0000014b, 5'd2, 27'h00000141, 32'h00000400,
  1'd1,  5'd11, 27'h00000124, 5'd18, 27'h00000327, 5'd14, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000347, 5'd15, 27'h000002d6, 5'd21, 27'h00000325, 32'h00000400,
  1'd1,  5'd14, 27'h000002ad, 5'd25, 27'h0000035f, 5'd0, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000006a, 5'd26, 27'h0000014d, 5'd14, 27'h00000012, 32'h00000400,
  1'd1,  5'd12, 27'h0000015e, 5'd26, 27'h000001d1, 5'd25, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000330, 5'd8, 27'h000002a0, 5'd3, 27'h000001a7, 32'h00000400,
  1'd1,  5'd24, 27'h000002a0, 5'd5, 27'h00000143, 5'd11, 27'h00000130, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000d7, 5'd20, 27'h0000027e, 5'd4, 27'h000003ba, 32'h00000400,
  1'd1,  5'd23, 27'h000002ac, 5'd15, 27'h00000289, 5'd11, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ea, 5'd18, 27'h00000293, 5'd25, 27'h00000000, 32'h00000400,
  1'd1,  5'd24, 27'h000002f9, 5'd27, 27'h0000011e, 5'd0, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000341, 5'd28, 27'h00000304, 5'd15, 27'h0000019e, 32'h00000400,
  1'd1,  5'd23, 27'h00000380, 5'd26, 27'h00000091, 5'd23, 27'h000001d1, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000a1, 5'd5, 27'h00000299, 5'd7, 27'h0000006f, 32'h00000400,
  1'd1,  5'd3, 27'h000000f6, 5'd7, 27'h00000001, 5'd17, 27'h0000014d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000365, 5'd5, 27'h000003ad, 5'd26, 27'h00000161, 32'h00000400,
  1'd1,  5'd2, 27'h00000151, 5'd19, 27'h0000011f, 5'd7, 27'h000000c1, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000025e, 5'd18, 27'h000000cc, 5'd20, 27'h000001f1, 32'h00000400,
  1'd1,  5'd4, 27'h0000005f, 5'd19, 27'h000001e8, 5'd29, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000277, 5'd27, 27'h0000016b, 5'd6, 27'h0000032c, 32'h00000400,
  1'd1,  5'd1, 27'h0000032c, 5'd28, 27'h000000c6, 5'd15, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001bd, 5'd26, 27'h00000050, 5'd30, 27'h0000005e, 32'h00000400,
  1'd1,  5'd13, 27'h000001da, 5'd7, 27'h00000175, 5'd5, 27'h0000014e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001d2, 5'd6, 27'h0000016c, 5'd16, 27'h000002a1, 32'h00000400,
  1'd1,  5'd13, 27'h0000038d, 5'd6, 27'h00000007, 5'd28, 27'h000000bf, 32'hfffffc00,
  1'd1,  5'd12, 27'h000002ec, 5'd16, 27'h00000371, 5'd6, 27'h0000027f, 32'h00000400,
  1'd1,  5'd13, 27'h00000055, 5'd17, 27'h000002cf, 5'd16, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000018, 5'd15, 27'h000003ad, 5'd30, 27'h000003d3, 32'h00000400,
  1'd1,  5'd12, 27'h00000190, 5'd28, 27'h0000038a, 5'd8, 27'h000002b2, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000011d, 5'd30, 27'h0000011a, 5'd17, 27'h000002b6, 32'h00000400,
  1'd1,  5'd11, 27'h0000015a, 5'd28, 27'h00000359, 5'd29, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000ca, 5'd10, 27'h00000033, 5'd5, 27'h00000358, 32'h00000400,
  1'd1,  5'd21, 27'h0000034b, 5'd9, 27'h0000010e, 5'd16, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e5, 5'd6, 27'h0000002b, 5'd25, 27'h00000368, 32'h00000400,
  1'd1,  5'd24, 27'h000001ae, 5'd15, 27'h00000336, 5'd6, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000001d, 5'd17, 27'h0000037b, 5'd18, 27'h00000310, 32'h00000400,
  1'd1,  5'd22, 27'h0000020b, 5'd20, 27'h0000029e, 5'd29, 27'h0000039b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002d1, 5'd30, 27'h000000c1, 5'd9, 27'h00000019, 32'h00000400,
  1'd1,  5'd22, 27'h000002f7, 5'd28, 27'h000001f2, 5'd18, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000087, 5'd27, 27'h000000fb, 5'd26, 27'h000000d3, 32'h00000400,
  1'd1,  5'd8, 27'h000000a1, 5'd1, 27'h000003f3, 5'd7, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000030a, 5'd2, 27'h00000080, 5'd18, 27'h000001de, 32'h00000400,
  1'd1,  5'd5, 27'h00000339, 5'd0, 27'h000003de, 5'd26, 27'h0000007c, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000200, 5'd10, 27'h000003f7, 5'd3, 27'h0000020c, 32'h00000400,
  1'd1,  5'd9, 27'h000002fe, 5'd14, 27'h00000150, 5'd13, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000302, 5'd10, 27'h0000033b, 5'd24, 27'h00000242, 32'h00000400,
  1'd1,  5'd5, 27'h000000ff, 5'd22, 27'h00000007, 5'd1, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000360, 5'd23, 27'h000003f6, 5'd10, 27'h00000315, 32'h00000400,
  1'd1,  5'd6, 27'h00000262, 5'd21, 27'h0000002b, 5'd22, 27'h00000150, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000283, 5'd1, 27'h00000266, 5'd9, 27'h0000005e, 32'h00000400,
  1'd1,  5'd18, 27'h00000248, 5'd3, 27'h000003c0, 5'd18, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000167, 5'd3, 27'h00000309, 5'd28, 27'h000001fe, 32'h00000400,
  1'd1,  5'd15, 27'h000002a1, 5'd13, 27'h0000019d, 5'd4, 27'h000003f7, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000039f, 5'd14, 27'h00000004, 5'd13, 27'h00000144, 32'h00000400,
  1'd1,  5'd19, 27'h0000025d, 5'd11, 27'h000002f9, 5'd21, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000025a, 5'd24, 27'h000000b3, 5'd0, 27'h0000039e, 32'h00000400,
  1'd1,  5'd18, 27'h000001d2, 5'd25, 27'h000001f5, 5'd11, 27'h000003f3, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001d2, 5'd21, 27'h0000038e, 5'd25, 27'h000002de, 32'h00000400,
  1'd1,  5'd30, 27'h000000bc, 5'd0, 27'h000001f2, 5'd2, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001ea, 5'd4, 27'h00000184, 5'd14, 27'h000002c5, 32'h00000400,
  1'd1,  5'd28, 27'h00000237, 5'd5, 27'h00000035, 5'd22, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000227, 5'd12, 27'h00000172, 5'd5, 27'h0000008c, 32'h00000400,
  1'd1,  5'd29, 27'h0000033d, 5'd12, 27'h000000f3, 5'd14, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002be, 5'd14, 27'h00000205, 5'd23, 27'h00000087, 32'h00000400,
  1'd1,  5'd26, 27'h0000029d, 5'd24, 27'h000003bd, 5'd1, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000017b, 5'd21, 27'h000003a3, 5'd11, 27'h0000025b, 32'h00000400,
  1'd1,  5'd27, 27'h00000148, 5'd23, 27'h000001df, 5'd22, 27'h00000381, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000002, 5'd1, 27'h00000356, 5'd0, 27'h0000013d, 32'h00000400,
  1'd1,  5'd6, 27'h0000031b, 5'd0, 27'h00000324, 5'd11, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003e9, 5'd2, 27'h0000021a, 5'd20, 27'h000002cf, 32'h00000400,
  1'd1,  5'd8, 27'h00000003, 5'd15, 27'h00000174, 5'd9, 27'h00000158, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000284, 5'd11, 27'h000003c4, 5'd15, 27'h00000352, 32'h00000400,
  1'd1,  5'd8, 27'h000003ab, 5'd14, 27'h0000011f, 5'd29, 27'h000001df, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000cb, 5'd25, 27'h0000022c, 5'd8, 27'h00000097, 32'h00000400,
  1'd1,  5'd6, 27'h00000356, 5'd24, 27'h000002f6, 5'd20, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000297, 5'd23, 27'h00000234, 5'd29, 27'h000003b9, 32'h00000400,
  1'd1,  5'd18, 27'h000001f6, 5'd0, 27'h00000120, 5'd0, 27'h00000395, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000088, 5'd3, 27'h0000037d, 5'd11, 27'h0000009c, 32'h00000400,
  1'd1,  5'd17, 27'h000000ba, 5'd12, 27'h000001b3, 5'd8, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000023a, 5'd11, 27'h0000014a, 5'd18, 27'h000002da, 32'h00000400,
  1'd1,  5'd17, 27'h000002bf, 5'd14, 27'h00000186, 5'd26, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000370, 5'd24, 27'h00000192, 5'd8, 27'h0000003d, 32'h00000400,
  1'd1,  5'd20, 27'h0000005b, 5'd20, 27'h000002cb, 5'd18, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000283, 5'd23, 27'h00000078, 5'd27, 27'h00000323, 32'h00000400,
  1'd1,  5'd28, 27'h000003b3, 5'd2, 27'h000001c4, 5'd6, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000025f, 5'd2, 27'h0000028a, 5'd18, 27'h00000271, 32'h00000400,
  1'd1,  5'd30, 27'h00000274, 5'd2, 27'h000000b5, 5'd27, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002bb, 5'd14, 27'h00000163, 5'd9, 27'h000000ba, 32'h00000400,
  1'd1,  5'd28, 27'h00000022, 5'd13, 27'h000001aa, 5'd15, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000021f, 5'd11, 27'h00000288, 5'd30, 27'h00000041, 32'h00000400,
  1'd1,  5'd30, 27'h00000094, 5'd24, 27'h00000125, 5'd9, 27'h00000339, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000032d, 5'd22, 27'h00000172, 5'd15, 27'h00000380, 32'h00000400,
  1'd1,  5'd29, 27'h000001d8, 5'd23, 27'h000001c7, 5'd29, 27'h00000331, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000b2, 5'd7, 27'h00000066, 5'd0, 27'h00000193, 32'h00000400,
  1'd1,  5'd9, 27'h00000011, 5'd9, 27'h000001bc, 5'd13, 27'h0000022e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000026a, 5'd8, 27'h0000002a, 5'd25, 27'h00000341, 32'h00000400,
  1'd1,  5'd5, 27'h000000ef, 5'd15, 27'h0000031e, 5'd3, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000a7, 5'd16, 27'h0000025b, 5'd15, 27'h0000013e, 32'h00000400,
  1'd1,  5'd6, 27'h0000033d, 5'd18, 27'h00000376, 5'd21, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000162, 5'd28, 27'h00000300, 5'd2, 27'h000001cc, 32'h00000400,
  1'd1,  5'd8, 27'h000002ce, 5'd27, 27'h00000139, 5'd14, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000104, 5'd28, 27'h00000313, 5'd25, 27'h0000030f, 32'h00000400,
  1'd1,  5'd19, 27'h0000019b, 5'd5, 27'h00000142, 5'd4, 27'h000001b9, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000022a, 5'd8, 27'h000002c2, 5'd12, 27'h000003ae, 32'h00000400,
  1'd1,  5'd18, 27'h00000369, 5'd6, 27'h000001d3, 5'd21, 27'h000000ec, 32'hfffffc00,
  1'd1,  5'd20, 27'h000001bd, 5'd18, 27'h00000211, 5'd0, 27'h000000d2, 32'h00000400,
  1'd1,  5'd19, 27'h00000335, 5'd17, 27'h0000012d, 5'd13, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000018f, 5'd20, 27'h00000116, 5'd23, 27'h000003f9, 32'h00000400,
  1'd1,  5'd16, 27'h000002e1, 5'd30, 27'h0000022a, 5'd0, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003c3, 5'd28, 27'h0000026a, 5'd11, 27'h00000262, 32'h00000400,
  1'd1,  5'd16, 27'h000003be, 5'd29, 27'h00000327, 5'd21, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000026a, 5'd6, 27'h00000124, 5'd4, 27'h0000028d, 32'h00000400,
  1'd1,  5'd30, 27'h00000245, 5'd9, 27'h00000390, 5'd11, 27'h00000312, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000011a, 5'd5, 27'h000001b7, 5'd25, 27'h0000033a, 32'h00000400,
  1'd1,  5'd29, 27'h00000033, 5'd16, 27'h000002f6, 5'd4, 27'h0000031a, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b2, 5'd19, 27'h0000012d, 5'd11, 27'h000001f1, 32'h00000400,
  1'd1,  5'd26, 27'h000003d8, 5'd17, 27'h00000011, 5'd22, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000ab, 5'd28, 27'h0000003d, 5'd3, 27'h00000190, 32'h00000400,
  1'd1,  5'd27, 27'h00000215, 5'd27, 27'h00000312, 5'd12, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000052, 5'd29, 27'h0000014e, 5'd21, 27'h0000016e, 32'h00000400,
  1'd1,  5'd7, 27'h00000271, 5'd9, 27'h0000002b, 5'd9, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000131, 5'd5, 27'h000002ca, 5'd30, 27'h00000037, 32'h00000400,
  1'd1,  5'd5, 27'h00000262, 5'd17, 27'h0000003b, 5'd8, 27'h00000141, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000331, 5'd19, 27'h0000003f, 5'd15, 27'h0000033c, 32'h00000400,
  1'd1,  5'd6, 27'h000001a9, 5'd19, 27'h00000176, 5'd29, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000009b, 5'd29, 27'h0000036e, 5'd8, 27'h00000381, 32'h00000400,
  1'd1,  5'd6, 27'h00000345, 5'd30, 27'h00000285, 5'd19, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000185, 5'd26, 27'h000001f5, 5'd29, 27'h0000014d, 32'h00000400,
  1'd1,  5'd16, 27'h00000042, 5'd6, 27'h0000033c, 5'd10, 27'h00000081, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000008b, 5'd6, 27'h0000028c, 5'd19, 27'h000003b8, 32'h00000400,
  1'd1,  5'd16, 27'h0000011c, 5'd9, 27'h000000e7, 5'd30, 27'h0000006b, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000289, 5'd17, 27'h0000019b, 5'd9, 27'h00000008, 32'h00000400,
  1'd1,  5'd16, 27'h000001d6, 5'd15, 27'h0000027c, 5'd20, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000385, 5'd15, 27'h000003e8, 5'd27, 27'h00000319, 32'h00000400,
  1'd1,  5'd17, 27'h00000383, 5'd28, 27'h0000014c, 5'd10, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000012d, 5'd27, 27'h00000108, 5'd17, 27'h000000ca, 32'h00000400,
  1'd1,  5'd15, 27'h000002f1, 5'd27, 27'h0000000f, 5'd29, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000a6, 5'd8, 27'h0000009c, 5'd7, 27'h00000318, 32'h00000400,
  1'd1,  5'd30, 27'h000002a1, 5'd10, 27'h00000056, 5'd18, 27'h0000016b, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002af, 5'd7, 27'h00000245, 5'd29, 27'h000000b9, 32'h00000400,
  1'd1,  5'd29, 27'h00000127, 5'd17, 27'h00000166, 5'd8, 27'h0000015b, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000018, 5'd18, 27'h000000b3, 5'd18, 27'h00000200, 32'h00000400,
  1'd1,  5'd27, 27'h000003d2, 5'd17, 27'h00000143, 5'd26, 27'h0000017c, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001f0, 5'd30, 27'h000002e5, 5'd6, 27'h00000348, 32'h00000400,
  1'd1,  5'd30, 27'h000000fd, 5'd29, 27'h000000b6, 5'd20, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003b5, 5'd29, 27'h00000094, 5'd30, 27'h0000007b, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h00000178, 5'd1, 27'h000002ad, 5'd0, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000012d, 5'd1, 27'h00000332, 5'd14, 27'h0000002a, 32'h00000400,
  1'd1,  5'd2, 27'h000003e2, 5'd3, 27'h000001d7, 5'd21, 27'h000002fe, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001da, 5'd11, 27'h0000003e, 5'd4, 27'h00000309, 32'h00000400,
  1'd1,  5'd5, 27'h00000085, 5'd10, 27'h0000032e, 5'd25, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036c, 5'd22, 27'h00000340, 5'd3, 27'h00000348, 32'h00000400,
  1'd1,  5'd0, 27'h00000195, 5'd22, 27'h00000396, 5'd15, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000020d, 5'd24, 27'h00000079, 5'd22, 27'h00000114, 32'h00000400,
  1'd1,  5'd13, 27'h000003e0, 5'd4, 27'h00000012, 5'd1, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000259, 5'd1, 27'h00000028, 5'd12, 27'h00000080, 32'h00000400,
  1'd1,  5'd13, 27'h000000a4, 5'd1, 27'h00000105, 5'd22, 27'h000002c0, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000117, 5'd11, 27'h00000022, 5'd4, 27'h0000005d, 32'h00000400,
  1'd1,  5'd15, 27'h00000071, 5'd15, 27'h000001c4, 5'd14, 27'h000001d9, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000034, 5'd12, 27'h0000001f, 5'd23, 27'h00000354, 32'h00000400,
  1'd1,  5'd15, 27'h00000041, 5'd21, 27'h000002c2, 5'd4, 27'h00000060, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000209, 5'd22, 27'h0000018e, 5'd14, 27'h000000c3, 32'h00000400,
  1'd1,  5'd10, 27'h000001ce, 5'd23, 27'h00000069, 5'd25, 27'h0000006a, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000220, 5'd4, 27'h000000e3, 5'd0, 27'h0000039b, 32'h00000400,
  1'd1,  5'd21, 27'h000003e1, 5'd1, 27'h000002bc, 5'd10, 27'h00000389, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000025e, 5'd2, 27'h00000289, 5'd23, 27'h00000328, 32'h00000400,
  1'd1,  5'd20, 27'h000003da, 5'd11, 27'h00000132, 5'd3, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000308, 5'd13, 27'h0000017f, 5'd11, 27'h000003eb, 32'h00000400,
  1'd1,  5'd20, 27'h000002dd, 5'd14, 27'h0000009c, 5'd22, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000329, 5'd23, 27'h0000008e, 5'd0, 27'h000000db, 32'h00000400,
  1'd1,  5'd23, 27'h0000000f, 5'd23, 27'h000001a3, 5'd15, 27'h000001b3, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000037a, 5'd25, 27'h00000084, 5'd25, 27'h00000224, 32'h00000400,
  1'd1,  5'd4, 27'h0000013c, 5'd0, 27'h000002b6, 5'd7, 27'h00000085, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000035a, 5'd3, 27'h00000335, 5'd19, 27'h0000004d, 32'h00000400,
  1'd1,  5'd0, 27'h0000005d, 5'd4, 27'h0000038f, 5'd30, 27'h00000297, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000021b, 5'd11, 27'h000002b2, 5'd8, 27'h000003ef, 32'h00000400,
  1'd1,  5'd0, 27'h00000143, 5'd14, 27'h0000002d, 5'd19, 27'h000000bb, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002e7, 5'd10, 27'h000003da, 5'd27, 27'h00000378, 32'h00000400,
  1'd1,  5'd1, 27'h00000216, 5'd21, 27'h00000129, 5'd7, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000375, 5'd21, 27'h000000ea, 5'd17, 27'h000001c1, 32'h00000400,
  1'd1,  5'd3, 27'h00000393, 5'd23, 27'h00000306, 5'd25, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003dd, 5'd4, 27'h000000b4, 5'd10, 27'h00000056, 32'h00000400,
  1'd1,  5'd13, 27'h0000021c, 5'd4, 27'h000002d4, 5'd18, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009b, 5'd1, 27'h0000002e, 5'd30, 27'h000002cf, 32'h00000400,
  1'd1,  5'd10, 27'h000001e4, 5'd14, 27'h000003ee, 5'd9, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000369, 5'd12, 27'h00000146, 5'd16, 27'h000000c4, 32'h00000400,
  1'd1,  5'd13, 27'h0000023d, 5'd14, 27'h0000022b, 5'd27, 27'h000000d4, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000253, 5'd25, 27'h00000161, 5'd7, 27'h00000176, 32'h00000400,
  1'd1,  5'd13, 27'h0000000c, 5'd24, 27'h00000236, 5'd17, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000037e, 5'd22, 27'h000001ba, 5'd28, 27'h0000002c, 32'h00000400,
  1'd1,  5'd20, 27'h00000343, 5'd4, 27'h00000098, 5'd9, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000291, 5'd0, 27'h000003fa, 5'd16, 27'h00000175, 32'h00000400,
  1'd1,  5'd22, 27'h000002cb, 5'd4, 27'h0000017e, 5'd25, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000275, 5'd12, 27'h0000030d, 5'd10, 27'h00000107, 32'h00000400,
  1'd1,  5'd24, 27'h000003dc, 5'd14, 27'h000002ee, 5'd17, 27'h000003ff, 32'hfffffc00,
  1'd1,  5'd22, 27'h000002d0, 5'd12, 27'h000002ed, 5'd28, 27'h000001f7, 32'h00000400,
  1'd1,  5'd23, 27'h00000184, 5'd21, 27'h0000032c, 5'd7, 27'h0000001b, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000304, 5'd25, 27'h0000015b, 5'd20, 27'h000000b1, 32'h00000400,
  1'd1,  5'd24, 27'h000003ed, 5'd21, 27'h0000000a, 5'd26, 27'h0000029b, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000279, 5'd7, 27'h000000ae, 5'd5, 27'h0000009d, 32'h00000400,
  1'd1,  5'd4, 27'h00000095, 5'd8, 27'h00000031, 5'd13, 27'h000001ae, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000032d, 5'd9, 27'h000002e9, 5'd23, 27'h0000039a, 32'h00000400,
  1'd1,  5'd4, 27'h000002fb, 5'd18, 27'h00000031, 5'd2, 27'h0000027e, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000038e, 5'd15, 27'h00000257, 5'd12, 27'h0000034f, 32'h00000400,
  1'd1,  5'd2, 27'h00000128, 5'd19, 27'h00000307, 5'd22, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001ec, 5'd26, 27'h0000017a, 5'd2, 27'h0000019c, 32'h00000400,
  1'd1,  5'd2, 27'h0000025b, 5'd29, 27'h000001c3, 5'd14, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd4, 27'h000002f4, 5'd28, 27'h0000027a, 5'd21, 27'h0000006c, 32'h00000400,
  1'd1,  5'd13, 27'h00000379, 5'd7, 27'h000002b2, 5'd4, 27'h000002e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000108, 5'd9, 27'h00000374, 5'd10, 27'h00000306, 32'h00000400,
  1'd1,  5'd14, 27'h000000eb, 5'd9, 27'h0000018b, 5'd22, 27'h0000013d, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000029a, 5'd18, 27'h000003c1, 5'd0, 27'h000000f2, 32'h00000400,
  1'd1,  5'd12, 27'h00000017, 5'd19, 27'h00000315, 5'd13, 27'h000002b4, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000167, 5'd15, 27'h000002ec, 5'd25, 27'h000002af, 32'h00000400,
  1'd1,  5'd13, 27'h000003d4, 5'd30, 27'h00000344, 5'd4, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000013, 5'd26, 27'h00000338, 5'd11, 27'h0000030b, 32'h00000400,
  1'd1,  5'd14, 27'h0000028e, 5'd27, 27'h000001e8, 5'd23, 27'h000001e1, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000091, 5'd6, 27'h000002dd, 5'd3, 27'h000001b1, 32'h00000400,
  1'd1,  5'd23, 27'h00000177, 5'd8, 27'h00000122, 5'd13, 27'h0000010c, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002ad, 5'd19, 27'h00000185, 5'd4, 27'h0000037b, 32'h00000400,
  1'd1,  5'd23, 27'h00000038, 5'd20, 27'h000000c5, 5'd15, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003c3, 5'd16, 27'h00000111, 5'd22, 27'h000003b2, 32'h00000400,
  1'd1,  5'd21, 27'h0000005b, 5'd29, 27'h00000277, 5'd0, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd24, 27'h000002ed, 5'd29, 27'h00000192, 5'd15, 27'h00000153, 32'h00000400,
  1'd1,  5'd24, 27'h000000db, 5'd26, 27'h00000290, 5'd21, 27'h000003ce, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000ff, 5'd7, 27'h00000236, 5'd7, 27'h0000017f, 32'h00000400,
  1'd1,  5'd4, 27'h000003c2, 5'd9, 27'h0000030f, 5'd16, 27'h00000329, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003a4, 5'd9, 27'h000000fa, 5'd29, 27'h0000021d, 32'h00000400,
  1'd1,  5'd2, 27'h0000005e, 5'd17, 27'h0000013b, 5'd9, 27'h000000c2, 32'hfffffc00,
  1'd1,  5'd4, 27'h000003e4, 5'd17, 27'h0000003d, 5'd17, 27'h000000a8, 32'h00000400,
  1'd1,  5'd3, 27'h0000010f, 5'd19, 27'h0000039c, 5'd28, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039c, 5'd30, 27'h0000032d, 5'd6, 27'h00000145, 32'h00000400,
  1'd1,  5'd2, 27'h00000045, 5'd29, 27'h00000288, 5'd16, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000039b, 5'd30, 27'h0000013e, 5'd28, 27'h0000036b, 32'h00000400,
  1'd1,  5'd11, 27'h00000048, 5'd7, 27'h00000040, 5'd7, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002eb, 5'd6, 27'h000002ac, 5'd15, 27'h00000369, 32'h00000400,
  1'd1,  5'd14, 27'h00000376, 5'd6, 27'h000002f3, 5'd27, 27'h000003eb, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001d7, 5'd20, 27'h000000c6, 5'd5, 27'h0000018c, 32'h00000400,
  1'd1,  5'd11, 27'h000003c2, 5'd20, 27'h000000a5, 5'd16, 27'h000000f0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000395, 5'd18, 27'h000003a3, 5'd29, 27'h000003e1, 32'h00000400,
  1'd1,  5'd14, 27'h00000258, 5'd28, 27'h000001b9, 5'd9, 27'h000000f8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000339, 5'd27, 27'h00000081, 5'd17, 27'h00000292, 32'h00000400,
  1'd1,  5'd11, 27'h00000231, 5'd30, 27'h000000b4, 5'd28, 27'h000003f1, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000346, 5'd9, 27'h000000f7, 5'd6, 27'h00000282, 32'h00000400,
  1'd1,  5'd22, 27'h00000259, 5'd5, 27'h00000198, 5'd18, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd24, 27'h000003b4, 5'd10, 27'h0000008d, 5'd28, 27'h0000025f, 32'h00000400,
  1'd1,  5'd23, 27'h000003dc, 5'd15, 27'h0000034b, 5'd9, 27'h0000037b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000000fd, 5'd15, 27'h000003ad, 5'd20, 27'h00000009, 32'h00000400,
  1'd1,  5'd21, 27'h000000e1, 5'd20, 27'h00000186, 5'd27, 27'h000001fc, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000044, 5'd29, 27'h000002e1, 5'd6, 27'h00000146, 32'h00000400,
  1'd1,  5'd20, 27'h00000339, 5'd29, 27'h00000391, 5'd20, 27'h00000280, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000011b, 5'd28, 27'h00000224, 5'd26, 27'h0000027a, 32'h00000400,
  1'd1,  5'd5, 27'h000000fc, 5'd1, 27'h00000207, 5'd7, 27'h00000031, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001c8, 5'd2, 27'h0000006d, 5'd19, 27'h000003e2, 32'h00000400,
  1'd1,  5'd9, 27'h00000120, 5'd2, 27'h00000081, 5'd28, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000281, 5'd15, 27'h000000e7, 5'd0, 27'h000002fb, 32'h00000400,
  1'd1,  5'd6, 27'h00000326, 5'd13, 27'h00000075, 5'd13, 27'h0000011c, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001d0, 5'd10, 27'h00000217, 5'd22, 27'h00000202, 32'h00000400,
  1'd1,  5'd9, 27'h00000382, 5'd23, 27'h000002eb, 5'd4, 27'h000000cb, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000003f, 5'd21, 27'h00000302, 5'd13, 27'h000002c2, 32'h00000400,
  1'd1,  5'd6, 27'h00000044, 5'd23, 27'h000003aa, 5'd25, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000036b, 5'd3, 27'h0000030c, 5'd6, 27'h00000057, 32'h00000400,
  1'd1,  5'd18, 27'h00000395, 5'd2, 27'h0000021a, 5'd19, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000024a, 5'd2, 27'h000003f6, 5'd28, 27'h000003ae, 32'h00000400,
  1'd1,  5'd19, 27'h000003fd, 5'd14, 27'h0000028b, 5'd1, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000215, 5'd14, 27'h000000e2, 5'd13, 27'h000003d1, 32'h00000400,
  1'd1,  5'd19, 27'h0000033d, 5'd15, 27'h00000005, 5'd22, 27'h00000153, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000217, 5'd23, 27'h0000020e, 5'd4, 27'h00000079, 32'h00000400,
  1'd1,  5'd17, 27'h00000055, 5'd20, 27'h0000039d, 5'd12, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000031c, 5'd25, 27'h0000027b, 5'd23, 27'h000002a5, 32'h00000400,
  1'd1,  5'd28, 27'h000002f5, 5'd2, 27'h0000004a, 5'd0, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001ea, 5'd4, 27'h00000046, 5'd14, 27'h000001a3, 32'h00000400,
  1'd1,  5'd26, 27'h00000297, 5'd3, 27'h00000032, 5'd25, 27'h0000012f, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000002b, 5'd12, 27'h000002f8, 5'd2, 27'h00000042, 32'h00000400,
  1'd1,  5'd29, 27'h000001f0, 5'd14, 27'h000000e0, 5'd10, 27'h0000036f, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000291, 5'd12, 27'h00000214, 5'd25, 27'h00000085, 32'h00000400,
  1'd1,  5'd28, 27'h000000ca, 5'd25, 27'h00000117, 5'd4, 27'h000002bd, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000119, 5'd21, 27'h000003ff, 5'd13, 27'h00000389, 32'h00000400,
  1'd1,  5'd29, 27'h0000024f, 5'd24, 27'h000002ba, 5'd24, 27'h00000325, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d0, 5'd0, 27'h0000018a, 5'd3, 27'h00000238, 32'h00000400,
  1'd1,  5'd9, 27'h00000273, 5'd0, 27'h00000148, 5'd12, 27'h000002e9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000325, 5'd3, 27'h00000337, 5'd25, 27'h00000303, 32'h00000400,
  1'd1,  5'd10, 27'h0000003f, 5'd11, 27'h000000c4, 5'd7, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000134, 5'd11, 27'h0000034e, 5'd20, 27'h000000f6, 32'h00000400,
  1'd1,  5'd9, 27'h00000159, 5'd12, 27'h00000225, 5'd27, 27'h00000197, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000be, 5'd20, 27'h000002f6, 5'd10, 27'h00000032, 32'h00000400,
  1'd1,  5'd8, 27'h0000017b, 5'd24, 27'h000001a8, 5'd19, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000022c, 5'd21, 27'h00000375, 5'd28, 27'h000000a9, 32'h00000400,
  1'd1,  5'd16, 27'h0000023c, 5'd4, 27'h000002f7, 5'd0, 27'h00000059, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000049, 5'd1, 27'h000000f8, 5'd11, 27'h000003b3, 32'h00000400,
  1'd1,  5'd19, 27'h0000027e, 5'd13, 27'h000002e8, 5'd5, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001f, 5'd12, 27'h000003a3, 5'd16, 27'h00000310, 32'h00000400,
  1'd1,  5'd18, 27'h00000079, 5'd12, 27'h000000ee, 5'd29, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000025e, 5'd21, 27'h00000391, 5'd8, 27'h00000391, 32'h00000400,
  1'd1,  5'd18, 27'h00000352, 5'd22, 27'h000001e6, 5'd16, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000173, 5'd21, 27'h000000da, 5'd27, 27'h000002ff, 32'h00000400,
  1'd1,  5'd27, 27'h000003ac, 5'd2, 27'h00000199, 5'd8, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000002e, 5'd2, 27'h0000032e, 5'd16, 27'h000000ad, 32'h00000400,
  1'd1,  5'd26, 27'h00000230, 5'd3, 27'h00000301, 5'd27, 27'h0000007e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000011, 5'd13, 27'h000001fb, 5'd8, 27'h00000341, 32'h00000400,
  1'd1,  5'd30, 27'h000002e8, 5'd11, 27'h0000037f, 5'd19, 27'h000000ab, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000059, 5'd15, 27'h00000037, 5'd26, 27'h000001c3, 32'h00000400,
  1'd1,  5'd27, 27'h00000194, 5'd25, 27'h00000261, 5'd9, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003ca, 5'd25, 27'h000002a6, 5'd16, 27'h00000395, 32'h00000400,
  1'd1,  5'd26, 27'h000003fe, 5'd21, 27'h00000098, 5'd30, 27'h000001da, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003d9, 5'd7, 27'h00000146, 5'd3, 27'h0000023c, 32'h00000400,
  1'd1,  5'd5, 27'h00000131, 5'd8, 27'h000003a2, 5'd10, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002a7, 5'd5, 27'h00000328, 5'd25, 27'h0000006e, 32'h00000400,
  1'd1,  5'd8, 27'h00000397, 5'd17, 27'h000003fd, 5'd2, 27'h00000110, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d8, 5'd16, 27'h000000f3, 5'd11, 27'h000002a0, 32'h00000400,
  1'd1,  5'd9, 27'h00000112, 5'd17, 27'h0000026a, 5'd23, 27'h000000d0, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a4, 5'd30, 27'h00000355, 5'd1, 27'h000001e5, 32'h00000400,
  1'd1,  5'd9, 27'h00000035, 5'd26, 27'h00000312, 5'd11, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000f5, 5'd30, 27'h000001a5, 5'd23, 27'h00000108, 32'h00000400,
  1'd1,  5'd17, 27'h00000365, 5'd5, 27'h00000284, 5'd2, 27'h00000058, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000de, 5'd10, 27'h0000005a, 5'd12, 27'h0000018e, 32'h00000400,
  1'd1,  5'd18, 27'h000000d5, 5'd7, 27'h000000e7, 5'd23, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001b, 5'd19, 27'h000003aa, 5'd0, 27'h0000016b, 32'h00000400,
  1'd1,  5'd19, 27'h00000298, 5'd17, 27'h000001c4, 5'd11, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001f5, 5'd17, 27'h000002d9, 5'd21, 27'h000002b5, 32'h00000400,
  1'd1,  5'd17, 27'h000002b4, 5'd30, 27'h000001ad, 5'd0, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000e0, 5'd30, 27'h00000101, 5'd10, 27'h00000157, 32'h00000400,
  1'd1,  5'd15, 27'h000002b7, 5'd29, 27'h000002cd, 5'd21, 27'h000003dd, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000393, 5'd8, 27'h00000209, 5'd2, 27'h0000021f, 32'h00000400,
  1'd1,  5'd30, 27'h0000022c, 5'd8, 27'h000002c0, 5'd13, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000da, 5'd7, 27'h00000384, 5'd22, 27'h000003cd, 32'h00000400,
  1'd1,  5'd27, 27'h0000022f, 5'd16, 27'h000001de, 5'd2, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002e3, 5'd16, 27'h00000158, 5'd12, 27'h000001c0, 32'h00000400,
  1'd1,  5'd29, 27'h0000039c, 5'd19, 27'h0000028b, 5'd21, 27'h000002a6, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000398, 5'd27, 27'h0000037f, 5'd0, 27'h0000036d, 32'h00000400,
  1'd1,  5'd26, 27'h00000341, 5'd27, 27'h00000098, 5'd13, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000050, 5'd27, 27'h0000003b, 5'd22, 27'h00000041, 32'h00000400,
  1'd1,  5'd8, 27'h00000228, 5'd7, 27'h00000126, 5'd5, 27'h0000011d, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000229, 5'd5, 27'h0000010f, 5'd26, 27'h0000031b, 32'h00000400,
  1'd1,  5'd9, 27'h000003b7, 5'd20, 27'h000000e8, 5'd7, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000273, 5'd17, 27'h00000071, 5'd15, 27'h00000379, 32'h00000400,
  1'd1,  5'd6, 27'h000002fe, 5'd17, 27'h0000020c, 5'd30, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001e4, 5'd29, 27'h000003e7, 5'd9, 27'h0000022f, 32'h00000400,
  1'd1,  5'd6, 27'h000001b0, 5'd30, 27'h00000247, 5'd19, 27'h0000028c, 32'hfffffc00,
  1'd1,  5'd9, 27'h000002d9, 5'd26, 27'h000002e3, 5'd26, 27'h0000025d, 32'h00000400,
  1'd1,  5'd19, 27'h00000163, 5'd6, 27'h0000014a, 5'd6, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000236, 5'd8, 27'h00000259, 5'd15, 27'h0000022d, 32'h00000400,
  1'd1,  5'd19, 27'h0000004f, 5'd8, 27'h00000335, 5'd26, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000d8, 5'd19, 27'h0000013e, 5'd7, 27'h000001eb, 32'h00000400,
  1'd1,  5'd17, 27'h00000262, 5'd16, 27'h000000c1, 5'd16, 27'h000001ee, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000043, 5'd18, 27'h0000003b, 5'd27, 27'h00000308, 32'h00000400,
  1'd1,  5'd18, 27'h00000364, 5'd27, 27'h00000317, 5'd8, 27'h000000de, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000091, 5'd30, 27'h000001e6, 5'd19, 27'h00000225, 32'h00000400,
  1'd1,  5'd15, 27'h000003af, 5'd30, 27'h000001c4, 5'd29, 27'h000001e7, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002c8, 5'd5, 27'h000000e3, 5'd7, 27'h0000020e, 32'h00000400,
  1'd1,  5'd26, 27'h00000024, 5'd8, 27'h0000027f, 5'd19, 27'h0000025c, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000016e, 5'd5, 27'h0000016d, 5'd27, 27'h00000008, 32'h00000400,
  1'd1,  5'd26, 27'h00000250, 5'd20, 27'h000000a8, 5'd7, 27'h000001fb, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000339, 5'd17, 27'h00000202, 5'd15, 27'h00000358, 32'h00000400,
  1'd1,  5'd28, 27'h000003c4, 5'd17, 27'h00000160, 5'd30, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003bf, 5'd26, 27'h00000028, 5'd7, 27'h0000029b, 32'h00000400,
  1'd1,  5'd30, 27'h0000028c, 5'd26, 27'h0000024a, 5'd18, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003a4, 5'd30, 27'h000002a1, 5'd28, 27'h000001fd, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h0000017f, 5'd4, 27'h000001a6, 5'd1, 27'h00000133, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000382, 5'd4, 27'h0000027c, 5'd13, 27'h00000270, 32'h00000400,
  1'd1,  5'd1, 27'h00000039, 5'd1, 27'h000002e8, 5'd21, 27'h00000022, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000008a, 5'd10, 27'h000001a7, 5'd2, 27'h00000017, 32'h00000400,
  1'd1,  5'd1, 27'h00000292, 5'd13, 27'h000002ec, 5'd23, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003ff, 5'd21, 27'h00000261, 5'd4, 27'h00000294, 32'h00000400,
  1'd1,  5'd1, 27'h0000037c, 5'd23, 27'h000003a4, 5'd15, 27'h000001a8, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000015c, 5'd21, 27'h000003d8, 5'd25, 27'h0000016a, 32'h00000400,
  1'd1,  5'd10, 27'h00000380, 5'd4, 27'h0000028d, 5'd4, 27'h000002c5, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000009d, 5'd3, 27'h000001e1, 5'd12, 27'h000001a3, 32'h00000400,
  1'd1,  5'd10, 27'h000003f4, 5'd2, 27'h00000183, 5'd25, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000372, 5'd13, 27'h0000024d, 5'd4, 27'h00000191, 32'h00000400,
  1'd1,  5'd15, 27'h000000a2, 5'd11, 27'h00000068, 5'd13, 27'h00000005, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000331, 5'd14, 27'h0000002c, 5'd25, 27'h00000242, 32'h00000400,
  1'd1,  5'd11, 27'h0000033e, 5'd21, 27'h00000366, 5'd4, 27'h00000257, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000225, 5'd24, 27'h000000c6, 5'd10, 27'h000003e9, 32'h00000400,
  1'd1,  5'd14, 27'h0000029a, 5'd22, 27'h00000060, 5'd24, 27'h000001fd, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003aa, 5'd0, 27'h000000b3, 5'd5, 27'h00000021, 32'h00000400,
  1'd1,  5'd22, 27'h0000038b, 5'd1, 27'h000001ef, 5'd14, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000248, 5'd3, 27'h000000ec, 5'd22, 27'h0000030a, 32'h00000400,
  1'd1,  5'd25, 27'h000002c8, 5'd11, 27'h00000283, 5'd3, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001ea, 5'd11, 27'h00000373, 5'd13, 27'h000003f8, 32'h00000400,
  1'd1,  5'd21, 27'h0000006e, 5'd14, 27'h000002f2, 5'd23, 27'h000003c1, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000037, 5'd24, 27'h000002f0, 5'd2, 27'h00000392, 32'h00000400,
  1'd1,  5'd22, 27'h0000030d, 5'd24, 27'h0000002b, 5'd11, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000db, 5'd24, 27'h000002a9, 5'd24, 27'h000002f8, 32'h00000400,
  1'd1,  5'd2, 27'h00000124, 5'd2, 27'h0000025e, 5'd6, 27'h0000038e, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000027a, 5'd4, 27'h000001b4, 5'd18, 27'h000000e4, 32'h00000400,
  1'd1,  5'd3, 27'h000002df, 5'd4, 27'h000000b4, 5'd27, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000361, 5'd13, 27'h00000274, 5'd6, 27'h00000171, 32'h00000400,
  1'd1,  5'd2, 27'h00000174, 5'd13, 27'h000000e3, 5'd17, 27'h0000026a, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000120, 5'd10, 27'h00000238, 5'd26, 27'h00000293, 32'h00000400,
  1'd1,  5'd4, 27'h00000118, 5'd21, 27'h00000095, 5'd7, 27'h00000238, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000248, 5'd21, 27'h00000169, 5'd16, 27'h0000039d, 32'h00000400,
  1'd1,  5'd4, 27'h000000bc, 5'd23, 27'h00000304, 5'd26, 27'h0000038b, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000222, 5'd1, 27'h00000039, 5'd6, 27'h000002cb, 32'h00000400,
  1'd1,  5'd11, 27'h0000032a, 5'd4, 27'h000001a5, 5'd17, 27'h00000090, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ab, 5'd1, 27'h0000038f, 5'd27, 27'h000000ea, 32'h00000400,
  1'd1,  5'd12, 27'h000000c8, 5'd13, 27'h000002e0, 5'd5, 27'h000003af, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000015b, 5'd14, 27'h0000019d, 5'd17, 27'h0000015c, 32'h00000400,
  1'd1,  5'd13, 27'h00000295, 5'd12, 27'h0000017a, 5'd30, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000301, 5'd22, 27'h0000033b, 5'd8, 27'h00000346, 32'h00000400,
  1'd1,  5'd15, 27'h000001c6, 5'd22, 27'h0000024d, 5'd19, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd11, 27'h000002e4, 5'd22, 27'h0000005e, 5'd27, 27'h000001ab, 32'h00000400,
  1'd1,  5'd23, 27'h00000326, 5'd1, 27'h000003f6, 5'd7, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd23, 27'h000001da, 5'd1, 27'h00000261, 5'd16, 27'h0000018b, 32'h00000400,
  1'd1,  5'd25, 27'h00000241, 5'd0, 27'h00000107, 5'd28, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000370, 5'd14, 27'h00000034, 5'd10, 27'h00000114, 32'h00000400,
  1'd1,  5'd25, 27'h000001c6, 5'd14, 27'h00000173, 5'd16, 27'h000002be, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000df, 5'd11, 27'h00000335, 5'd26, 27'h00000307, 32'h00000400,
  1'd1,  5'd21, 27'h00000265, 5'd22, 27'h00000366, 5'd5, 27'h000002c2, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000102, 5'd25, 27'h000000b8, 5'd18, 27'h00000222, 32'h00000400,
  1'd1,  5'd22, 27'h00000377, 5'd22, 27'h000003dd, 5'd28, 27'h000002cf, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000020, 5'd5, 27'h000000fb, 5'd3, 27'h000003d2, 32'h00000400,
  1'd1,  5'd1, 27'h00000095, 5'd8, 27'h00000001, 5'd15, 27'h00000104, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000381, 5'd6, 27'h000000b1, 5'd22, 27'h000001d4, 32'h00000400,
  1'd1,  5'd3, 27'h000002bd, 5'd16, 27'h0000015a, 5'd1, 27'h000002a5, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000367, 5'd16, 27'h00000355, 5'd14, 27'h00000279, 32'h00000400,
  1'd1,  5'd0, 27'h00000200, 5'd19, 27'h00000319, 5'd25, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003e7, 5'd30, 27'h0000008a, 5'd2, 27'h00000276, 32'h00000400,
  1'd1,  5'd0, 27'h00000221, 5'd29, 27'h000000c9, 5'd11, 27'h000001ad, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000088, 5'd27, 27'h000001fe, 5'd23, 27'h00000204, 32'h00000400,
  1'd1,  5'd15, 27'h0000002b, 5'd5, 27'h00000324, 5'd0, 27'h00000198, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000ee, 5'd8, 27'h00000103, 5'd13, 27'h0000034f, 32'h00000400,
  1'd1,  5'd11, 27'h0000039a, 5'd9, 27'h00000152, 5'd25, 27'h00000288, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000017d, 5'd15, 27'h00000361, 5'd2, 27'h00000255, 32'h00000400,
  1'd1,  5'd14, 27'h00000339, 5'd18, 27'h000000ce, 5'd14, 27'h00000138, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003d9, 5'd19, 27'h000001dc, 5'd21, 27'h00000244, 32'h00000400,
  1'd1,  5'd13, 27'h00000148, 5'd28, 27'h000001cf, 5'd2, 27'h00000317, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000234, 5'd25, 27'h0000038b, 5'd14, 27'h000002cd, 32'h00000400,
  1'd1,  5'd12, 27'h0000017c, 5'd28, 27'h000003f4, 5'd25, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000093, 5'd5, 27'h0000022f, 5'd3, 27'h00000162, 32'h00000400,
  1'd1,  5'd23, 27'h00000136, 5'd5, 27'h000000eb, 5'd13, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000398, 5'd19, 27'h00000363, 5'd0, 27'h0000004b, 32'h00000400,
  1'd1,  5'd24, 27'h000002c8, 5'd19, 27'h0000013a, 5'd10, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000120, 5'd18, 27'h000002cf, 5'd23, 27'h000001bc, 32'h00000400,
  1'd1,  5'd23, 27'h00000305, 5'd29, 27'h000001f0, 5'd0, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000020a, 5'd29, 27'h00000333, 5'd13, 27'h0000027d, 32'h00000400,
  1'd1,  5'd21, 27'h00000145, 5'd28, 27'h0000039b, 5'd21, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003bc, 5'd5, 27'h00000353, 5'd5, 27'h000000b2, 32'h00000400,
  1'd1,  5'd1, 27'h00000258, 5'd8, 27'h00000031, 5'd16, 27'h0000012b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000018c, 5'd6, 27'h00000304, 5'd27, 27'h00000392, 32'h00000400,
  1'd1,  5'd4, 27'h00000091, 5'd20, 27'h000000bc, 5'd8, 27'h0000008b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000008c, 5'd16, 27'h00000315, 5'd17, 27'h000001ff, 32'h00000400,
  1'd1,  5'd0, 27'h0000013d, 5'd17, 27'h0000034f, 5'd28, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000008a, 5'd27, 27'h0000013a, 5'd10, 27'h00000072, 32'h00000400,
  1'd1,  5'd3, 27'h00000198, 5'd27, 27'h00000251, 5'd20, 27'h00000199, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000008b, 5'd30, 27'h000003a2, 5'd26, 27'h00000163, 32'h00000400,
  1'd1,  5'd14, 27'h0000013f, 5'd9, 27'h00000024, 5'd5, 27'h0000030d, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000239, 5'd7, 27'h000002b7, 5'd16, 27'h000001fc, 32'h00000400,
  1'd1,  5'd14, 27'h000002e3, 5'd5, 27'h000001f1, 5'd29, 27'h00000247, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000036, 5'd17, 27'h0000002f, 5'd10, 27'h0000007a, 32'h00000400,
  1'd1,  5'd14, 27'h000002c1, 5'd18, 27'h000002be, 5'd20, 27'h0000020e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000fe, 5'd17, 27'h00000042, 5'd27, 27'h00000399, 32'h00000400,
  1'd1,  5'd10, 27'h00000360, 5'd30, 27'h000002be, 5'd7, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003cc, 5'd27, 27'h00000328, 5'd19, 27'h000003f4, 32'h00000400,
  1'd1,  5'd14, 27'h0000002c, 5'd29, 27'h0000018b, 5'd29, 27'h00000101, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000322, 5'd6, 27'h00000153, 5'd10, 27'h000000e5, 32'h00000400,
  1'd1,  5'd25, 27'h00000326, 5'd10, 27'h00000056, 5'd16, 27'h000000db, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000a0, 5'd8, 27'h00000326, 5'd26, 27'h0000015c, 32'h00000400,
  1'd1,  5'd24, 27'h000000d4, 5'd16, 27'h00000352, 5'd7, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd20, 27'h000003be, 5'd20, 27'h000001b0, 5'd19, 27'h0000036e, 32'h00000400,
  1'd1,  5'd21, 27'h00000311, 5'd18, 27'h000002b7, 5'd28, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd22, 27'h000003f2, 5'd26, 27'h0000039e, 5'd8, 27'h000001a9, 32'h00000400,
  1'd1,  5'd22, 27'h000001a2, 5'd26, 27'h000003fe, 5'd16, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000287, 5'd27, 27'h000001c4, 5'd28, 27'h000000f1, 32'h00000400,
  1'd1,  5'd5, 27'h00000291, 5'd2, 27'h000000d5, 5'd9, 27'h00000294, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000388, 5'd0, 27'h00000343, 5'd19, 27'h00000146, 32'h00000400,
  1'd1,  5'd10, 27'h0000012f, 5'd4, 27'h000000cd, 5'd28, 27'h0000018e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000062, 5'd14, 27'h000001cf, 5'd1, 27'h00000248, 32'h00000400,
  1'd1,  5'd7, 27'h00000021, 5'd11, 27'h00000207, 5'd12, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000005b, 5'd10, 27'h00000187, 5'd25, 27'h00000044, 32'h00000400,
  1'd1,  5'd9, 27'h000000c1, 5'd20, 27'h000002bb, 5'd2, 27'h000003cb, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000308, 5'd23, 27'h00000358, 5'd11, 27'h00000303, 32'h00000400,
  1'd1,  5'd8, 27'h00000293, 5'd22, 27'h000001aa, 5'd24, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f3, 5'd0, 27'h00000173, 5'd9, 27'h0000016a, 32'h00000400,
  1'd1,  5'd17, 27'h00000035, 5'd0, 27'h00000302, 5'd15, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000369, 5'd0, 27'h0000000a, 5'd29, 27'h00000055, 32'h00000400,
  1'd1,  5'd15, 27'h00000209, 5'd11, 27'h000003b0, 5'd2, 27'h000003ef, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000025, 5'd13, 27'h00000341, 5'd15, 27'h000000bb, 32'h00000400,
  1'd1,  5'd18, 27'h0000001e, 5'd11, 27'h0000025b, 5'd22, 27'h00000223, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000032a, 5'd25, 27'h00000117, 5'd0, 27'h00000071, 32'h00000400,
  1'd1,  5'd16, 27'h000000ec, 5'd22, 27'h00000132, 5'd11, 27'h00000099, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000009b, 5'd22, 27'h00000136, 5'd21, 27'h00000125, 32'h00000400,
  1'd1,  5'd28, 27'h000003f9, 5'd3, 27'h000003e9, 5'd4, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000353, 5'd2, 27'h00000040, 5'd14, 27'h0000039f, 32'h00000400,
  1'd1,  5'd27, 27'h0000011a, 5'd4, 27'h0000016c, 5'd25, 27'h0000010d, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000025, 5'd11, 27'h00000316, 5'd0, 27'h00000047, 32'h00000400,
  1'd1,  5'd27, 27'h000001fa, 5'd15, 27'h000000c7, 5'd12, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003b3, 5'd13, 27'h000000e1, 5'd21, 27'h00000228, 32'h00000400,
  1'd1,  5'd28, 27'h00000079, 5'd22, 27'h00000093, 5'd5, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000042, 5'd22, 27'h0000026b, 5'd14, 27'h000003a3, 32'h00000400,
  1'd1,  5'd30, 27'h0000004f, 5'd22, 27'h00000019, 5'd25, 27'h00000093, 32'hfffffc00,
  1'd1,  5'd8, 27'h000001f5, 5'd4, 27'h00000289, 5'd0, 27'h00000007, 32'h00000400,
  1'd1,  5'd9, 27'h000002ea, 5'd2, 27'h00000161, 5'd13, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002c5, 5'd5, 27'h0000005f, 5'd22, 27'h000002c3, 32'h00000400,
  1'd1,  5'd6, 27'h0000037c, 5'd15, 27'h00000120, 5'd9, 27'h000003b6, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000025b, 5'd11, 27'h000002ad, 5'd17, 27'h0000024b, 32'h00000400,
  1'd1,  5'd8, 27'h00000220, 5'd10, 27'h000001e5, 5'd26, 27'h0000017a, 32'hfffffc00,
  1'd1,  5'd6, 27'h000000b1, 5'd23, 27'h00000138, 5'd7, 27'h00000232, 32'h00000400,
  1'd1,  5'd8, 27'h000002d0, 5'd22, 27'h000000c6, 5'd19, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000304, 5'd23, 27'h00000288, 5'd30, 27'h00000282, 32'h00000400,
  1'd1,  5'd18, 27'h0000022d, 5'd1, 27'h000000d7, 5'd3, 27'h000002ac, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000241, 5'd2, 27'h00000145, 5'd14, 27'h00000033, 32'h00000400,
  1'd1,  5'd19, 27'h000000ce, 5'd14, 27'h0000019f, 5'd7, 27'h0000010e, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000274, 5'd11, 27'h000002cf, 5'd18, 27'h000002c2, 32'h00000400,
  1'd1,  5'd16, 27'h000002f6, 5'd14, 27'h000003ce, 5'd29, 27'h00000078, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000053, 5'd23, 27'h00000343, 5'd6, 27'h0000018c, 32'h00000400,
  1'd1,  5'd16, 27'h000001f4, 5'd25, 27'h0000019c, 5'd18, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001fe, 5'd25, 27'h000000e3, 5'd25, 27'h00000373, 32'h00000400,
  1'd1,  5'd27, 27'h000001bf, 5'd1, 27'h000001a9, 5'd5, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000391, 5'd4, 27'h00000276, 5'd18, 27'h00000242, 32'h00000400,
  1'd1,  5'd25, 27'h00000362, 5'd4, 27'h0000003e, 5'd28, 27'h0000002f, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000020d, 5'd12, 27'h00000180, 5'd5, 27'h00000128, 32'h00000400,
  1'd1,  5'd28, 27'h00000048, 5'd11, 27'h0000036f, 5'd15, 27'h0000033a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000389, 5'd13, 27'h0000023e, 5'd27, 27'h00000172, 32'h00000400,
  1'd1,  5'd27, 27'h0000012d, 5'd21, 27'h000001c6, 5'd9, 27'h000000f4, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000210, 5'd23, 27'h0000024b, 5'd18, 27'h00000333, 32'h00000400,
  1'd1,  5'd29, 27'h000002ce, 5'd21, 27'h00000122, 5'd26, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002da, 5'd6, 27'h00000298, 5'd2, 27'h00000287, 32'h00000400,
  1'd1,  5'd9, 27'h00000201, 5'd9, 27'h0000009a, 5'd12, 27'h000001dc, 32'hfffffc00,
  1'd1,  5'd6, 27'h000002d1, 5'd6, 27'h00000120, 5'd22, 27'h00000267, 32'h00000400,
  1'd1,  5'd7, 27'h000000a8, 5'd19, 27'h0000013d, 5'd0, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000152, 5'd19, 27'h00000157, 5'd14, 27'h00000336, 32'h00000400,
  1'd1,  5'd6, 27'h000000ca, 5'd15, 27'h000002d8, 5'd22, 27'h000003df, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023b, 5'd26, 27'h000002f0, 5'd4, 27'h000001aa, 32'h00000400,
  1'd1,  5'd8, 27'h0000005d, 5'd30, 27'h00000361, 5'd12, 27'h000001b6, 32'hfffffc00,
  1'd1,  5'd5, 27'h000000b2, 5'd26, 27'h00000064, 5'd23, 27'h000000e8, 32'h00000400,
  1'd1,  5'd19, 27'h00000330, 5'd8, 27'h00000314, 5'd0, 27'h00000072, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000006, 5'd9, 27'h000001e3, 5'd14, 27'h00000334, 32'h00000400,
  1'd1,  5'd17, 27'h00000043, 5'd5, 27'h0000022d, 5'd20, 27'h000002d8, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000029d, 5'd20, 27'h0000019b, 5'd4, 27'h0000026e, 32'h00000400,
  1'd1,  5'd17, 27'h00000211, 5'd17, 27'h000002f6, 5'd13, 27'h00000228, 32'hfffffc00,
  1'd1,  5'd20, 27'h000000b3, 5'd15, 27'h00000236, 5'd24, 27'h000002ff, 32'h00000400,
  1'd1,  5'd18, 27'h00000207, 5'd30, 27'h00000056, 5'd5, 27'h00000030, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000081, 5'd29, 27'h00000168, 5'd10, 27'h000002d1, 32'h00000400,
  1'd1,  5'd20, 27'h00000092, 5'd30, 27'h0000036d, 5'd25, 27'h0000033b, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000019c, 5'd7, 27'h0000035c, 5'd3, 27'h000003e8, 32'h00000400,
  1'd1,  5'd26, 27'h0000022d, 5'd5, 27'h0000028c, 5'd12, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003f9, 5'd6, 27'h0000038d, 5'd24, 27'h000003fb, 32'h00000400,
  1'd1,  5'd26, 27'h00000322, 5'd20, 27'h0000012c, 5'd3, 27'h000003c3, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000218, 5'd17, 27'h00000265, 5'd11, 27'h00000352, 32'h00000400,
  1'd1,  5'd27, 27'h000002c0, 5'd19, 27'h0000033b, 5'd23, 27'h0000035d, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000054, 5'd29, 27'h00000392, 5'd0, 27'h00000273, 32'h00000400,
  1'd1,  5'd28, 27'h00000116, 5'd29, 27'h00000206, 5'd12, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000a8, 5'd28, 27'h0000000e, 5'd20, 27'h000003bf, 32'h00000400,
  1'd1,  5'd6, 27'h000000eb, 5'd7, 27'h00000105, 5'd9, 27'h00000037, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000286, 5'd7, 27'h000002a2, 5'd27, 27'h000002eb, 32'h00000400,
  1'd1,  5'd7, 27'h00000276, 5'd16, 27'h00000037, 5'd8, 27'h00000298, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000297, 5'd18, 27'h0000032c, 5'd17, 27'h00000353, 32'h00000400,
  1'd1,  5'd5, 27'h0000027a, 5'd19, 27'h000001ae, 5'd30, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000245, 5'd26, 27'h00000400, 5'd6, 27'h00000319, 32'h00000400,
  1'd1,  5'd6, 27'h0000009f, 5'd26, 27'h00000321, 5'd17, 27'h00000341, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000036, 5'd28, 27'h00000030, 5'd26, 27'h00000261, 32'h00000400,
  1'd1,  5'd19, 27'h00000379, 5'd7, 27'h0000025d, 5'd7, 27'h00000128, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002d9, 5'd6, 27'h00000136, 5'd18, 27'h0000015b, 32'h00000400,
  1'd1,  5'd18, 27'h0000020a, 5'd9, 27'h0000037a, 5'd27, 27'h000003c9, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000356, 5'd18, 27'h0000034f, 5'd6, 27'h000000c8, 32'h00000400,
  1'd1,  5'd20, 27'h00000087, 5'd18, 27'h00000298, 5'd18, 27'h00000249, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002f9, 5'd16, 27'h0000034f, 5'd29, 27'h0000024f, 32'h00000400,
  1'd1,  5'd19, 27'h00000044, 5'd28, 27'h00000196, 5'd8, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000255, 5'd28, 27'h0000013c, 5'd19, 27'h000001c0, 32'h00000400,
  1'd1,  5'd20, 27'h000000fe, 5'd30, 27'h0000036d, 5'd27, 27'h000003c4, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000300, 5'd6, 27'h00000076, 5'd10, 27'h0000004d, 32'h00000400,
  1'd1,  5'd29, 27'h000002ee, 5'd9, 27'h0000033b, 5'd19, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000365, 5'd5, 27'h00000261, 5'd30, 27'h00000036, 32'h00000400,
  1'd1,  5'd30, 27'h0000009c, 5'd16, 27'h0000010e, 5'd8, 27'h00000177, 32'hfffffc00,
  1'd1,  5'd26, 27'h000003c1, 5'd16, 27'h0000031f, 5'd20, 27'h00000279, 32'h00000400,
  1'd1,  5'd26, 27'h0000015e, 5'd17, 27'h0000030c, 5'd29, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000376, 5'd30, 27'h000003bd, 5'd8, 27'h000001fd, 32'h00000400,
  1'd1,  5'd25, 27'h0000038d, 5'd28, 27'h00000397, 5'd19, 27'h000000a5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003dc, 5'd29, 27'h0000016b, 5'd29, 27'h00000249, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h00000079, 5'd2, 27'h00000289, 5'd2, 27'h0000007a, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000073, 5'd4, 27'h00000187, 5'd14, 27'h000001f9, 32'h00000400,
  1'd1,  5'd3, 27'h000002d7, 5'd0, 27'h00000239, 5'd20, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000128, 5'd14, 27'h00000179, 5'd2, 27'h00000388, 32'h00000400,
  1'd1,  5'd2, 27'h000001b3, 5'd11, 27'h0000020d, 5'd21, 27'h0000005e, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000375, 5'd24, 27'h000001d3, 5'd4, 27'h000000dd, 32'h00000400,
  1'd1,  5'd3, 27'h000001a5, 5'd23, 27'h0000015b, 5'd11, 27'h0000003b, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000008c, 5'd22, 27'h000000f7, 5'd22, 27'h00000271, 32'h00000400,
  1'd1,  5'd11, 27'h000000b3, 5'd2, 27'h000001f4, 5'd3, 27'h00000252, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002ef, 5'd3, 27'h0000034d, 5'd12, 27'h000002d1, 32'h00000400,
  1'd1,  5'd15, 27'h0000009e, 5'd1, 27'h00000047, 5'd21, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003e9, 5'd14, 27'h00000106, 5'd3, 27'h00000166, 32'h00000400,
  1'd1,  5'd11, 27'h000000b2, 5'd12, 27'h00000062, 5'd12, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000031a, 5'd13, 27'h00000236, 5'd22, 27'h000002fd, 32'h00000400,
  1'd1,  5'd12, 27'h00000114, 5'd21, 27'h000002d4, 5'd3, 27'h000000f5, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000035, 5'd25, 27'h00000051, 5'd15, 27'h000001cc, 32'h00000400,
  1'd1,  5'd12, 27'h00000282, 5'd23, 27'h000000fb, 5'd22, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000081, 5'd0, 27'h0000028e, 5'd1, 27'h000002b1, 32'h00000400,
  1'd1,  5'd23, 27'h0000013d, 5'd4, 27'h00000155, 5'd13, 27'h000001bd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000108, 5'd0, 27'h000000a0, 5'd21, 27'h0000037a, 32'h00000400,
  1'd1,  5'd25, 27'h00000046, 5'd15, 27'h00000198, 5'd4, 27'h000002c4, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000228, 5'd15, 27'h000001bd, 5'd12, 27'h0000005d, 32'h00000400,
  1'd1,  5'd23, 27'h0000005d, 5'd11, 27'h0000018b, 5'd24, 27'h000000e4, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002f7, 5'd22, 27'h00000204, 5'd1, 27'h0000020f, 32'h00000400,
  1'd1,  5'd24, 27'h0000028a, 5'd22, 27'h00000343, 5'd10, 27'h00000274, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000230, 5'd21, 27'h000001e9, 5'd22, 27'h000003ce, 32'h00000400,
  1'd1,  5'd4, 27'h0000030e, 5'd2, 27'h0000018a, 5'd5, 27'h000002bc, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000254, 5'd3, 27'h00000294, 5'd20, 27'h0000020f, 32'h00000400,
  1'd1,  5'd3, 27'h00000032, 5'd1, 27'h000002d4, 5'd27, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd2, 27'h000002da, 5'd11, 27'h00000252, 5'd6, 27'h000003bf, 32'h00000400,
  1'd1,  5'd3, 27'h00000146, 5'd12, 27'h000001f8, 5'd16, 27'h000003d3, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000000b, 5'd12, 27'h000002c8, 5'd28, 27'h00000342, 32'h00000400,
  1'd1,  5'd1, 27'h00000242, 5'd21, 27'h0000017d, 5'd5, 27'h000003f5, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002ea, 5'd24, 27'h00000004, 5'd16, 27'h0000009e, 32'h00000400,
  1'd1,  5'd2, 27'h00000128, 5'd21, 27'h000000ae, 5'd27, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ba, 5'd0, 27'h000002d6, 5'd5, 27'h0000035c, 32'h00000400,
  1'd1,  5'd11, 27'h00000251, 5'd1, 27'h000003e1, 5'd19, 27'h00000137, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000141, 5'd2, 27'h00000250, 5'd27, 27'h0000000b, 32'h00000400,
  1'd1,  5'd13, 27'h00000110, 5'd14, 27'h00000048, 5'd6, 27'h0000010f, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000017e, 5'd10, 27'h000002fc, 5'd19, 27'h0000018e, 32'h00000400,
  1'd1,  5'd13, 27'h00000154, 5'd10, 27'h000003f5, 5'd26, 27'h0000004b, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000c9, 5'd25, 27'h000000e9, 5'd6, 27'h0000013c, 32'h00000400,
  1'd1,  5'd12, 27'h000001ca, 5'd22, 27'h0000009e, 5'd18, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000272, 5'd22, 27'h00000254, 5'd27, 27'h00000366, 32'h00000400,
  1'd1,  5'd20, 27'h0000037d, 5'd1, 27'h0000009e, 5'd8, 27'h000001d8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000312, 5'd0, 27'h00000091, 5'd17, 27'h0000015d, 32'h00000400,
  1'd1,  5'd23, 27'h00000064, 5'd3, 27'h00000109, 5'd27, 27'h000003fc, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000227, 5'd11, 27'h00000360, 5'd9, 27'h00000303, 32'h00000400,
  1'd1,  5'd22, 27'h0000029c, 5'd13, 27'h00000165, 5'd18, 27'h00000209, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035d, 5'd12, 27'h00000075, 5'd29, 27'h0000013a, 32'h00000400,
  1'd1,  5'd25, 27'h000001f3, 5'd25, 27'h000002de, 5'd9, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000023c, 5'd24, 27'h0000007a, 5'd18, 27'h000000b9, 32'h00000400,
  1'd1,  5'd22, 27'h000002fc, 5'd21, 27'h00000294, 5'd26, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002d4, 5'd8, 27'h00000055, 5'd2, 27'h000002d9, 32'h00000400,
  1'd1,  5'd4, 27'h000002f6, 5'd8, 27'h00000141, 5'd11, 27'h000002f8, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001b1, 5'd8, 27'h0000001d, 5'd25, 27'h0000028d, 32'h00000400,
  1'd1,  5'd2, 27'h00000119, 5'd18, 27'h0000008c, 5'd4, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000020b, 5'd17, 27'h00000006, 5'd12, 27'h00000214, 32'h00000400,
  1'd1,  5'd1, 27'h00000352, 5'd16, 27'h00000072, 5'd21, 27'h00000258, 32'hfffffc00,
  1'd1,  5'd2, 27'h000001ae, 5'd26, 27'h0000031a, 5'd0, 27'h000001f1, 32'h00000400,
  1'd1,  5'd1, 27'h0000001d, 5'd28, 27'h00000024, 5'd13, 27'h000002db, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000107, 5'd28, 27'h000001d1, 5'd24, 27'h00000342, 32'h00000400,
  1'd1,  5'd11, 27'h000000c7, 5'd7, 27'h000000f0, 5'd1, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd10, 27'h000002ec, 5'd7, 27'h000001b6, 5'd11, 27'h00000186, 32'h00000400,
  1'd1,  5'd15, 27'h000001bc, 5'd8, 27'h000003db, 5'd24, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000028f, 5'd15, 27'h000003b7, 5'd1, 27'h00000064, 32'h00000400,
  1'd1,  5'd14, 27'h0000011c, 5'd17, 27'h00000009, 5'd10, 27'h0000025e, 32'hfffffc00,
  1'd1,  5'd13, 27'h000000c3, 5'd15, 27'h0000023c, 5'd24, 27'h00000059, 32'h00000400,
  1'd1,  5'd14, 27'h00000240, 5'd28, 27'h00000216, 5'd0, 27'h000003ea, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000bd, 5'd27, 27'h000001a5, 5'd13, 27'h000001bb, 32'h00000400,
  1'd1,  5'd11, 27'h0000039b, 5'd30, 27'h0000012e, 5'd23, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001bd, 5'd5, 27'h00000285, 5'd5, 27'h00000082, 32'h00000400,
  1'd1,  5'd22, 27'h000000de, 5'd8, 27'h00000223, 5'd12, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000141, 5'd17, 27'h00000114, 5'd1, 27'h00000002, 32'h00000400,
  1'd1,  5'd22, 27'h00000057, 5'd16, 27'h0000034a, 5'd13, 27'h00000191, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000395, 5'd19, 27'h0000017e, 5'd25, 27'h0000018e, 32'h00000400,
  1'd1,  5'd21, 27'h00000116, 5'd30, 27'h00000295, 5'd1, 27'h000000ee, 32'hfffffc00,
  1'd1,  5'd24, 27'h000000a2, 5'd27, 27'h0000016f, 5'd14, 27'h0000037e, 32'h00000400,
  1'd1,  5'd23, 27'h00000379, 5'd30, 27'h0000025f, 5'd21, 27'h00000143, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000197, 5'd6, 27'h0000024b, 5'd5, 27'h000002df, 32'h00000400,
  1'd1,  5'd2, 27'h00000285, 5'd8, 27'h0000004f, 5'd18, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000011b, 5'd7, 27'h0000029f, 5'd27, 27'h000001e5, 32'h00000400,
  1'd1,  5'd1, 27'h00000271, 5'd18, 27'h000003ce, 5'd5, 27'h00000336, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001bf, 5'd19, 27'h00000297, 5'd16, 27'h000001e6, 32'h00000400,
  1'd1,  5'd5, 27'h00000034, 5'd19, 27'h00000362, 5'd28, 27'h00000043, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000000c, 5'd26, 27'h000002d8, 5'd5, 27'h000002c7, 32'h00000400,
  1'd1,  5'd1, 27'h0000013d, 5'd26, 27'h000003fe, 5'd17, 27'h0000004d, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003d5, 5'd30, 27'h00000102, 5'd29, 27'h00000210, 32'h00000400,
  1'd1,  5'd14, 27'h000003a5, 5'd8, 27'h00000001, 5'd8, 27'h00000149, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003a2, 5'd8, 27'h000002ed, 5'd16, 27'h00000326, 32'h00000400,
  1'd1,  5'd14, 27'h00000390, 5'd6, 27'h000001ff, 5'd27, 27'h000001c1, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000333, 5'd20, 27'h00000010, 5'd6, 27'h00000282, 32'h00000400,
  1'd1,  5'd15, 27'h000001d4, 5'd18, 27'h000001ae, 5'd19, 27'h0000032e, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000198, 5'd17, 27'h000002c9, 5'd28, 27'h000000bd, 32'h00000400,
  1'd1,  5'd13, 27'h00000367, 5'd27, 27'h000001ef, 5'd7, 27'h000003c2, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003a8, 5'd26, 27'h0000023a, 5'd15, 27'h000002f8, 32'h00000400,
  1'd1,  5'd11, 27'h000002bf, 5'd29, 27'h00000130, 5'd26, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000323, 5'd7, 27'h0000035b, 5'd7, 27'h000002de, 32'h00000400,
  1'd1,  5'd25, 27'h000002a4, 5'd8, 27'h0000035a, 5'd18, 27'h0000007f, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000248, 5'd6, 27'h000002ae, 5'd30, 27'h0000004c, 32'h00000400,
  1'd1,  5'd24, 27'h0000014e, 5'd16, 27'h000003d6, 5'd6, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000345, 5'd18, 27'h000003ba, 5'd15, 27'h00000290, 32'h00000400,
  1'd1,  5'd25, 27'h00000137, 5'd20, 27'h00000234, 5'd26, 27'h00000075, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000140, 5'd26, 27'h000000c2, 5'd7, 27'h0000015d, 32'h00000400,
  1'd1,  5'd24, 27'h0000011b, 5'd28, 27'h00000385, 5'd17, 27'h0000022c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000016b, 5'd28, 27'h000003e7, 5'd27, 27'h0000036b, 32'h00000400,
  1'd1,  5'd7, 27'h000003a7, 5'd2, 27'h00000334, 5'd5, 27'h00000167, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000020c, 5'd3, 27'h000002e8, 5'd16, 27'h000000fd, 32'h00000400,
  1'd1,  5'd6, 27'h000001ac, 5'd2, 27'h00000120, 5'd29, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000018f, 5'd13, 27'h0000021b, 5'd2, 27'h0000007a, 32'h00000400,
  1'd1,  5'd7, 27'h00000376, 5'd10, 27'h0000030d, 5'd10, 27'h000003e2, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000330, 5'd11, 27'h000003c1, 5'd23, 27'h00000037, 32'h00000400,
  1'd1,  5'd6, 27'h0000011f, 5'd20, 27'h00000369, 5'd4, 27'h0000008d, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000346, 5'd20, 27'h000003c2, 5'd12, 27'h000000cf, 32'h00000400,
  1'd1,  5'd7, 27'h000002df, 5'd20, 27'h000003cf, 5'd25, 27'h00000293, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000131, 5'd5, 27'h0000009c, 5'd9, 27'h000002dd, 32'h00000400,
  1'd1,  5'd16, 27'h00000314, 5'd4, 27'h000000a0, 5'd16, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000063, 5'd3, 27'h000001fa, 5'd29, 27'h000000f2, 32'h00000400,
  1'd1,  5'd18, 27'h00000196, 5'd10, 27'h000003b8, 5'd2, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001b, 5'd10, 27'h00000304, 5'd22, 27'h0000014d, 32'h00000400,
  1'd1,  5'd20, 27'h0000014b, 5'd24, 27'h000002f3, 5'd2, 27'h000002e4, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002a8, 5'd21, 27'h000001ec, 5'd11, 27'h00000367, 32'h00000400,
  1'd1,  5'd19, 27'h000003ff, 5'd21, 27'h0000038a, 5'd21, 27'h00000053, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000292, 5'd2, 27'h00000012, 5'd0, 27'h000002ce, 32'h00000400,
  1'd1,  5'd28, 27'h00000150, 5'd4, 27'h000000bb, 5'd11, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000271, 5'd4, 27'h000000f2, 5'd21, 27'h0000004e, 32'h00000400,
  1'd1,  5'd30, 27'h00000197, 5'd12, 27'h000000d8, 5'd4, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000316, 5'd10, 27'h0000020a, 5'd10, 27'h000003fc, 32'h00000400,
  1'd1,  5'd30, 27'h00000080, 5'd12, 27'h000003b7, 5'd23, 27'h000001d6, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000014, 5'd22, 27'h000002ae, 5'd2, 27'h00000317, 32'h00000400,
  1'd1,  5'd26, 27'h0000026e, 5'd22, 27'h000001e1, 5'd11, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000390, 5'd23, 27'h00000029, 5'd21, 27'h000003e8, 32'h00000400,
  1'd1,  5'd8, 27'h0000032a, 5'd0, 27'h00000015, 5'd4, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000025d, 5'd4, 27'h000001f6, 5'd10, 27'h000001a9, 32'h00000400,
  1'd1,  5'd9, 27'h00000137, 5'd3, 27'h000003a3, 5'd25, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000013f, 5'd12, 27'h00000177, 5'd7, 27'h00000122, 32'h00000400,
  1'd1,  5'd6, 27'h000002d8, 5'd10, 27'h00000288, 5'd19, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000026c, 5'd15, 27'h000001c8, 5'd28, 27'h0000022e, 32'h00000400,
  1'd1,  5'd7, 27'h00000150, 5'd24, 27'h000001f0, 5'd9, 27'h000001d4, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000373, 5'd21, 27'h00000023, 5'd20, 27'h0000009b, 32'h00000400,
  1'd1,  5'd6, 27'h000000cb, 5'd23, 27'h0000007f, 5'd30, 27'h0000008f, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000a5, 5'd1, 27'h0000007a, 5'd3, 27'h00000172, 32'h00000400,
  1'd1,  5'd15, 27'h0000020d, 5'd0, 27'h00000354, 5'd11, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000331, 5'd10, 27'h000001fd, 5'd6, 27'h00000199, 32'h00000400,
  1'd1,  5'd19, 27'h000002b0, 5'd11, 27'h0000033a, 5'd17, 27'h0000027a, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000018c, 5'd14, 27'h000001c3, 5'd27, 27'h000002ca, 32'h00000400,
  1'd1,  5'd19, 27'h000003e7, 5'd23, 27'h000000d8, 5'd10, 27'h0000012a, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000385, 5'd22, 27'h00000252, 5'd17, 27'h00000018, 32'h00000400,
  1'd1,  5'd17, 27'h0000025c, 5'd22, 27'h000003a4, 5'd28, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000124, 5'd4, 27'h000002d4, 5'd9, 27'h000000a5, 32'h00000400,
  1'd1,  5'd28, 27'h000003c9, 5'd3, 27'h0000019c, 5'd20, 27'h00000148, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001cb, 5'd1, 27'h00000053, 5'd26, 27'h00000203, 32'h00000400,
  1'd1,  5'd27, 27'h00000259, 5'd15, 27'h00000192, 5'd9, 27'h000000fd, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000a2, 5'd15, 27'h000000b8, 5'd20, 27'h00000107, 32'h00000400,
  1'd1,  5'd29, 27'h00000277, 5'd13, 27'h000000f5, 5'd30, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000032d, 5'd23, 27'h0000021d, 5'd8, 27'h0000003c, 32'h00000400,
  1'd1,  5'd29, 27'h00000299, 5'd21, 27'h0000031d, 5'd16, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000003, 5'd24, 27'h000000e9, 5'd30, 27'h0000010b, 32'h00000400,
  1'd1,  5'd9, 27'h000002f2, 5'd10, 27'h0000006e, 5'd4, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000d, 5'd6, 27'h00000352, 5'd15, 27'h000000a0, 32'h00000400,
  1'd1,  5'd7, 27'h00000040, 5'd8, 27'h00000195, 5'd24, 27'h00000152, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000030f, 5'd18, 27'h000001a2, 5'd3, 27'h00000117, 32'h00000400,
  1'd1,  5'd7, 27'h00000247, 5'd20, 27'h00000223, 5'd10, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000009c, 5'd17, 27'h00000111, 5'd25, 27'h0000007a, 32'h00000400,
  1'd1,  5'd8, 27'h000003ea, 5'd27, 27'h000003db, 5'd4, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd7, 27'h000002df, 5'd29, 27'h000001f3, 5'd14, 27'h000002bd, 32'h00000400,
  1'd1,  5'd6, 27'h000000b2, 5'd27, 27'h000003d4, 5'd20, 27'h00000362, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000390, 5'd9, 27'h000002ea, 5'd1, 27'h0000020d, 32'h00000400,
  1'd1,  5'd20, 27'h0000002b, 5'd5, 27'h0000038b, 5'd11, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd18, 27'h00000281, 5'd7, 27'h000000f0, 5'd24, 27'h000002b3, 32'h00000400,
  1'd1,  5'd16, 27'h000002e0, 5'd17, 27'h000001d7, 5'd2, 27'h00000273, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001c8, 5'd15, 27'h00000317, 5'd13, 27'h00000347, 32'h00000400,
  1'd1,  5'd16, 27'h000002ce, 5'd19, 27'h000001b3, 5'd25, 27'h000002ce, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039e, 5'd28, 27'h000002ac, 5'd2, 27'h000000c6, 32'h00000400,
  1'd1,  5'd16, 27'h000003f8, 5'd27, 27'h000001a0, 5'd12, 27'h00000286, 32'hfffffc00,
  1'd1,  5'd16, 27'h000000e4, 5'd30, 27'h00000114, 5'd22, 27'h0000038f, 32'h00000400,
  1'd1,  5'd30, 27'h00000259, 5'd8, 27'h00000152, 5'd1, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000014, 5'd7, 27'h00000079, 5'd10, 27'h00000160, 32'h00000400,
  1'd1,  5'd28, 27'h000003a0, 5'd7, 27'h000000e4, 5'd24, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd29, 27'h000001b9, 5'd17, 27'h000002f1, 5'd3, 27'h000002e9, 32'h00000400,
  1'd1,  5'd27, 27'h00000260, 5'd20, 27'h00000135, 5'd15, 27'h00000116, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000193, 5'd17, 27'h0000033e, 5'd23, 27'h000002e5, 32'h00000400,
  1'd1,  5'd26, 27'h0000013a, 5'd30, 27'h00000158, 5'd3, 27'h00000221, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003a9, 5'd29, 27'h000001fe, 5'd14, 27'h000001d3, 32'h00000400,
  1'd1,  5'd29, 27'h00000357, 5'd30, 27'h00000371, 5'd23, 27'h000001d2, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000087, 5'd6, 27'h00000030, 5'd6, 27'h00000094, 32'h00000400,
  1'd1,  5'd7, 27'h00000303, 5'd8, 27'h00000133, 5'd29, 27'h00000264, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000032a, 5'd16, 27'h00000096, 5'd7, 27'h000001b2, 32'h00000400,
  1'd1,  5'd10, 27'h00000079, 5'd16, 27'h00000004, 5'd20, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003d4, 5'd18, 27'h0000028e, 5'd27, 27'h0000002e, 32'h00000400,
  1'd1,  5'd5, 27'h00000358, 5'd27, 27'h000000e1, 5'd8, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000017, 5'd30, 27'h000002d3, 5'd16, 27'h00000027, 32'h00000400,
  1'd1,  5'd7, 27'h000003d8, 5'd26, 27'h0000017d, 5'd27, 27'h00000368, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000037a, 5'd7, 27'h00000254, 5'd5, 27'h00000197, 32'h00000400,
  1'd1,  5'd17, 27'h000003e8, 5'd7, 27'h0000008f, 5'd19, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000002d, 5'd5, 27'h0000022d, 5'd28, 27'h000002cd, 32'h00000400,
  1'd1,  5'd18, 27'h000000f5, 5'd19, 27'h0000012b, 5'd8, 27'h00000244, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000231, 5'd17, 27'h000000a2, 5'd16, 27'h000003dd, 32'h00000400,
  1'd1,  5'd18, 27'h0000026f, 5'd19, 27'h000000ea, 5'd29, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000321, 5'd29, 27'h000000e4, 5'd8, 27'h000001e1, 32'h00000400,
  1'd1,  5'd15, 27'h0000035d, 5'd30, 27'h000003b4, 5'd16, 27'h0000038a, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003d2, 5'd30, 27'h00000091, 5'd30, 27'h000000bd, 32'h00000400,
  1'd1,  5'd29, 27'h0000022a, 5'd7, 27'h0000006a, 5'd8, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd28, 27'h000001b7, 5'd7, 27'h00000361, 5'd16, 27'h00000241, 32'h00000400,
  1'd1,  5'd27, 27'h000001d1, 5'd7, 27'h000003d4, 5'd28, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000034f, 5'd18, 27'h000001c7, 5'd8, 27'h00000351, 32'h00000400,
  1'd1,  5'd30, 27'h00000305, 5'd20, 27'h00000264, 5'd19, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001e9, 5'd17, 27'h00000152, 5'd26, 27'h0000006f, 32'h00000400,
  1'd1,  5'd30, 27'h00000201, 5'd30, 27'h00000342, 5'd9, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000200, 5'd30, 27'h00000349, 5'd16, 27'h00000036, 32'h00000400,
  1'd1,  5'd26, 27'h00000359, 5'd27, 27'h00000324, 5'd30, 27'h000001f2, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h0000019d, 5'd3, 27'h0000003a, 5'd4, 27'h000000a7, 32'h00000400,
  1'd1,  5'd1, 27'h0000031c, 5'd2, 27'h00000297, 5'd13, 27'h00000320, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000062, 5'd0, 27'h0000002b, 5'd25, 27'h0000011d, 32'h00000400,
  1'd1,  5'd2, 27'h00000359, 5'd13, 27'h000001f2, 5'd4, 27'h00000042, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000003b, 5'd12, 27'h0000033c, 5'd22, 27'h0000010e, 32'h00000400,
  1'd1,  5'd4, 27'h000001ac, 5'd24, 27'h00000350, 5'd0, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000004, 5'd21, 27'h00000260, 5'd12, 27'h0000015a, 32'h00000400,
  1'd1,  5'd1, 27'h00000052, 5'd25, 27'h00000317, 5'd21, 27'h0000038f, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a7, 5'd2, 27'h000000d7, 5'd1, 27'h00000222, 32'h00000400,
  1'd1,  5'd14, 27'h00000291, 5'd0, 27'h000003ae, 5'd11, 27'h0000037c, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000a7, 5'd4, 27'h00000209, 5'd24, 27'h0000023a, 32'h00000400,
  1'd1,  5'd11, 27'h00000277, 5'd12, 27'h0000013e, 5'd4, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000367, 5'd13, 27'h0000020c, 5'd15, 27'h0000005d, 32'h00000400,
  1'd1,  5'd13, 27'h0000013c, 5'd12, 27'h00000041, 5'd23, 27'h000001fa, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000316, 5'd25, 27'h0000008e, 5'd4, 27'h000003b5, 32'h00000400,
  1'd1,  5'd12, 27'h000000ec, 5'd25, 27'h00000281, 5'd13, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd13, 27'h000002c2, 5'd24, 27'h000002bc, 5'd21, 27'h000002b1, 32'h00000400,
  1'd1,  5'd22, 27'h00000228, 5'd0, 27'h00000113, 5'd3, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000300, 5'd2, 27'h0000027f, 5'd11, 27'h0000037a, 32'h00000400,
  1'd1,  5'd25, 27'h000001dc, 5'd3, 27'h00000107, 5'd24, 27'h00000344, 32'hfffffc00,
  1'd1,  5'd25, 27'h000001ce, 5'd11, 27'h00000334, 5'd4, 27'h000002d5, 32'h00000400,
  1'd1,  5'd25, 27'h00000134, 5'd12, 27'h00000074, 5'd12, 27'h000003f6, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000322, 5'd11, 27'h000002ce, 5'd21, 27'h0000030e, 32'h00000400,
  1'd1,  5'd25, 27'h00000311, 5'd23, 27'h00000127, 5'd2, 27'h00000108, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000276, 5'd21, 27'h00000357, 5'd11, 27'h000002e5, 32'h00000400,
  1'd1,  5'd20, 27'h000002e5, 5'd24, 27'h000000c2, 5'd24, 27'h000001ba, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000376, 5'd2, 27'h000003e6, 5'd6, 27'h00000369, 32'h00000400,
  1'd1,  5'd2, 27'h00000097, 5'd2, 27'h000000b5, 5'd19, 27'h0000009d, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000215, 5'd5, 27'h00000026, 5'd30, 27'h00000320, 32'h00000400,
  1'd1,  5'd1, 27'h00000308, 5'd11, 27'h00000098, 5'd5, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001d5, 5'd12, 27'h00000330, 5'd17, 27'h00000335, 32'h00000400,
  1'd1,  5'd0, 27'h00000315, 5'd12, 27'h000000b1, 5'd28, 27'h00000066, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001b4, 5'd24, 27'h000002ce, 5'd8, 27'h0000036a, 32'h00000400,
  1'd1,  5'd0, 27'h000003a3, 5'd21, 27'h00000295, 5'd18, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000259, 5'd22, 27'h00000214, 5'd30, 27'h000000d3, 32'h00000400,
  1'd1,  5'd12, 27'h00000028, 5'd3, 27'h00000380, 5'd9, 27'h000000ed, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000026, 5'd4, 27'h0000005f, 5'd19, 27'h0000035f, 32'h00000400,
  1'd1,  5'd14, 27'h00000260, 5'd3, 27'h00000361, 5'd29, 27'h00000291, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000fc, 5'd13, 27'h00000152, 5'd10, 27'h00000101, 32'h00000400,
  1'd1,  5'd15, 27'h000001bb, 5'd15, 27'h00000083, 5'd15, 27'h00000299, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000218, 5'd14, 27'h0000026b, 5'd27, 27'h00000129, 32'h00000400,
  1'd1,  5'd10, 27'h000002f7, 5'd24, 27'h00000361, 5'd9, 27'h00000050, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000319, 5'd23, 27'h00000280, 5'd16, 27'h00000290, 32'h00000400,
  1'd1,  5'd14, 27'h000001a8, 5'd24, 27'h00000152, 5'd27, 27'h000000c5, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003b8, 5'd2, 27'h000002bf, 5'd6, 27'h0000018c, 32'h00000400,
  1'd1,  5'd20, 27'h0000033a, 5'd3, 27'h00000327, 5'd17, 27'h000002e1, 32'hfffffc00,
  1'd1,  5'd21, 27'h000003e0, 5'd2, 27'h00000175, 5'd29, 27'h00000209, 32'h00000400,
  1'd1,  5'd21, 27'h0000031d, 5'd13, 27'h00000179, 5'd7, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000000a, 5'd11, 27'h00000167, 5'd18, 27'h000000f0, 32'h00000400,
  1'd1,  5'd24, 27'h000003ec, 5'd15, 27'h000000d8, 5'd27, 27'h00000272, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000017f, 5'd22, 27'h0000014d, 5'd6, 27'h0000003d, 32'h00000400,
  1'd1,  5'd22, 27'h0000039d, 5'd24, 27'h00000347, 5'd16, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000024e, 5'd25, 27'h00000185, 5'd29, 27'h00000006, 32'h00000400,
  1'd1,  5'd2, 27'h000002c4, 5'd8, 27'h00000042, 5'd4, 27'h00000164, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002fe, 5'd9, 27'h00000256, 5'd11, 27'h00000144, 32'h00000400,
  1'd1,  5'd4, 27'h0000000f, 5'd5, 27'h000001e3, 5'd25, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd3, 27'h000001be, 5'd18, 27'h00000352, 5'd0, 27'h000002ee, 32'h00000400,
  1'd1,  5'd0, 27'h000002af, 5'd19, 27'h000001ca, 5'd11, 27'h0000039a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000033b, 5'd20, 27'h0000025f, 5'd20, 27'h0000037b, 32'h00000400,
  1'd1,  5'd2, 27'h00000004, 5'd27, 27'h00000214, 5'd2, 27'h000000cf, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000379, 5'd29, 27'h00000011, 5'd10, 27'h00000291, 32'h00000400,
  1'd1,  5'd4, 27'h000003b9, 5'd30, 27'h00000273, 5'd24, 27'h00000303, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000155, 5'd6, 27'h0000027e, 5'd1, 27'h000001d6, 32'h00000400,
  1'd1,  5'd13, 27'h000002ad, 5'd6, 27'h000001d6, 5'd11, 27'h000001c2, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000099, 5'd7, 27'h000000f9, 5'd21, 27'h00000064, 32'h00000400,
  1'd1,  5'd15, 27'h0000002b, 5'd17, 27'h00000025, 5'd3, 27'h000003dc, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000020c, 5'd18, 27'h00000034, 5'd14, 27'h000000e7, 32'h00000400,
  1'd1,  5'd10, 27'h000001ee, 5'd16, 27'h0000035e, 5'd23, 27'h000000d1, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003a7, 5'd26, 27'h000001fc, 5'd1, 27'h000002fa, 32'h00000400,
  1'd1,  5'd14, 27'h00000062, 5'd27, 27'h000001ee, 5'd10, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000284, 5'd29, 27'h000002af, 5'd23, 27'h000001f9, 32'h00000400,
  1'd1,  5'd21, 27'h000002c1, 5'd9, 27'h0000033c, 5'd0, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000145, 5'd7, 27'h00000297, 5'd14, 27'h00000063, 32'h00000400,
  1'd1,  5'd25, 27'h00000346, 5'd15, 27'h00000392, 5'd2, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000003f, 5'd16, 27'h00000203, 5'd11, 27'h0000012c, 32'h00000400,
  1'd1,  5'd23, 27'h000000b6, 5'd17, 27'h0000036e, 5'd23, 27'h0000028a, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000000e, 5'd29, 27'h00000254, 5'd1, 27'h000000b6, 32'h00000400,
  1'd1,  5'd21, 27'h000000e9, 5'd26, 27'h000002ec, 5'd11, 27'h000001f0, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000109, 5'd28, 27'h0000015c, 5'd24, 27'h0000001a, 32'h00000400,
  1'd1,  5'd1, 27'h000003b2, 5'd9, 27'h000000df, 5'd10, 27'h0000012e, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000072, 5'd7, 27'h00000377, 5'd18, 27'h0000037c, 32'h00000400,
  1'd1,  5'd3, 27'h000001c9, 5'd6, 27'h00000076, 5'd30, 27'h000000cd, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000048, 5'd17, 27'h00000317, 5'd5, 27'h00000265, 32'h00000400,
  1'd1,  5'd3, 27'h000003ce, 5'd19, 27'h0000037f, 5'd18, 27'h000002eb, 32'hfffffc00,
  1'd1,  5'd0, 27'h000003c1, 5'd16, 27'h000002fc, 5'd29, 27'h0000034a, 32'h00000400,
  1'd1,  5'd1, 27'h00000335, 5'd26, 27'h0000033c, 5'd8, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd1, 27'h000001ed, 5'd29, 27'h00000046, 5'd18, 27'h0000001b, 32'h00000400,
  1'd1,  5'd1, 27'h00000093, 5'd26, 27'h0000032b, 5'd30, 27'h000003f9, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000008f, 5'd7, 27'h0000030b, 5'd8, 27'h000003b9, 32'h00000400,
  1'd1,  5'd15, 27'h000001bf, 5'd5, 27'h000002cc, 5'd17, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000017d, 5'd6, 27'h00000208, 5'd26, 27'h000002c7, 32'h00000400,
  1'd1,  5'd11, 27'h00000006, 5'd16, 27'h000001ee, 5'd5, 27'h0000033c, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000039b, 5'd18, 27'h00000263, 5'd18, 27'h000002cb, 32'h00000400,
  1'd1,  5'd13, 27'h00000180, 5'd17, 27'h000001f8, 5'd28, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd14, 27'h000001e1, 5'd28, 27'h00000338, 5'd7, 27'h000003bd, 32'h00000400,
  1'd1,  5'd15, 27'h000000c0, 5'd30, 27'h000002a9, 5'd16, 27'h00000079, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000016b, 5'd27, 27'h000002ed, 5'd28, 27'h000000b9, 32'h00000400,
  1'd1,  5'd25, 27'h00000343, 5'd5, 27'h000003f7, 5'd6, 27'h00000270, 32'hfffffc00,
  1'd1,  5'd23, 27'h000003c6, 5'd6, 27'h0000030c, 5'd17, 27'h0000007d, 32'h00000400,
  1'd1,  5'd23, 27'h0000018c, 5'd5, 27'h000003fc, 5'd27, 27'h00000399, 32'hfffffc00,
  1'd1,  5'd25, 27'h000002e9, 5'd18, 27'h0000007b, 5'd9, 27'h000002bc, 32'h00000400,
  1'd1,  5'd23, 27'h0000011f, 5'd17, 27'h00000351, 5'd19, 27'h00000194, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000231, 5'd15, 27'h00000341, 5'd29, 27'h0000016b, 32'h00000400,
  1'd1,  5'd24, 27'h000003f5, 5'd27, 27'h000000ce, 5'd8, 27'h00000044, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000032e, 5'd26, 27'h0000021e, 5'd18, 27'h000003cb, 32'h00000400,
  1'd1,  5'd21, 27'h000002c1, 5'd28, 27'h000000f9, 5'd26, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000375, 5'd0, 27'h00000029, 5'd6, 27'h0000035d, 32'h00000400,
  1'd1,  5'd8, 27'h00000227, 5'd2, 27'h00000034, 5'd20, 27'h000000d9, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000007e, 5'd0, 27'h000001c8, 5'd27, 27'h000000d2, 32'h00000400,
  1'd1,  5'd5, 27'h000003f6, 5'd15, 27'h000000bb, 5'd3, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000250, 5'd15, 27'h00000192, 5'd14, 27'h000002c3, 32'h00000400,
  1'd1,  5'd9, 27'h00000262, 5'd14, 27'h0000022b, 5'd24, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000239, 5'd25, 27'h0000003a, 5'd0, 27'h000002b8, 32'h00000400,
  1'd1,  5'd7, 27'h00000245, 5'd25, 27'h000000cb, 5'd11, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001be, 5'd20, 27'h000003ef, 5'd25, 27'h0000027f, 32'h00000400,
  1'd1,  5'd15, 27'h000002ac, 5'd1, 27'h000001bf, 5'd9, 27'h000000fb, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000010c, 5'd1, 27'h0000027c, 5'd20, 27'h000001dc, 32'h00000400,
  1'd1,  5'd15, 27'h00000210, 5'd2, 27'h000002a7, 5'd29, 27'h00000378, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000016e, 5'd14, 27'h000001f5, 5'd3, 27'h0000035c, 32'h00000400,
  1'd1,  5'd19, 27'h0000008b, 5'd11, 27'h00000388, 5'd25, 27'h000000d3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000ea, 5'd21, 27'h000000fa, 5'd1, 27'h0000022f, 32'h00000400,
  1'd1,  5'd16, 27'h000001ee, 5'd25, 27'h00000153, 5'd10, 27'h0000026c, 32'hfffffc00,
  1'd1,  5'd19, 27'h0000039e, 5'd22, 27'h000000b0, 5'd20, 27'h0000033b, 32'h00000400,
  1'd1,  5'd26, 27'h00000305, 5'd4, 27'h00000124, 5'd1, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000034f, 5'd2, 27'h00000068, 5'd15, 27'h00000150, 32'h00000400,
  1'd1,  5'd26, 27'h00000112, 5'd2, 27'h000000bc, 5'd22, 27'h000003ec, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002fe, 5'd12, 27'h0000005c, 5'd4, 27'h0000010e, 32'h00000400,
  1'd1,  5'd26, 27'h0000000e, 5'd10, 27'h0000024f, 5'd13, 27'h00000366, 32'hfffffc00,
  1'd1,  5'd27, 27'h000002e9, 5'd15, 27'h00000039, 5'd25, 27'h000000a4, 32'h00000400,
  1'd1,  5'd28, 27'h000002cb, 5'd23, 27'h00000237, 5'd4, 27'h0000004a, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000206, 5'd22, 27'h0000025b, 5'd11, 27'h00000389, 32'h00000400,
  1'd1,  5'd29, 27'h000002f7, 5'd21, 27'h00000039, 5'd22, 27'h00000098, 32'hfffffc00,
  1'd1,  5'd5, 27'h000003ac, 5'd3, 27'h00000350, 5'd4, 27'h00000059, 32'h00000400,
  1'd1,  5'd7, 27'h000001eb, 5'd2, 27'h000000c4, 5'd14, 27'h00000014, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000292, 5'd2, 27'h0000009a, 5'd24, 27'h00000084, 32'h00000400,
  1'd1,  5'd8, 27'h00000399, 5'd10, 27'h00000367, 5'd6, 27'h000003e9, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000247, 5'd13, 27'h000001bf, 5'd18, 27'h000000f5, 32'h00000400,
  1'd1,  5'd7, 27'h000000be, 5'd14, 27'h00000375, 5'd28, 27'h000003f0, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000013, 5'd23, 27'h00000238, 5'd7, 27'h000001fe, 32'h00000400,
  1'd1,  5'd9, 27'h00000234, 5'd25, 27'h0000028c, 5'd20, 27'h000000df, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000037c, 5'd23, 27'h00000146, 5'd28, 27'h0000007f, 32'h00000400,
  1'd1,  5'd18, 27'h00000324, 5'd4, 27'h000001d8, 5'd4, 27'h00000333, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002bc, 5'd0, 27'h000000f7, 5'd11, 27'h000001b0, 32'h00000400,
  1'd1,  5'd18, 27'h000000dc, 5'd13, 27'h0000036e, 5'd8, 27'h000002b3, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000033f, 5'd12, 27'h000001f7, 5'd18, 27'h0000006e, 32'h00000400,
  1'd1,  5'd19, 27'h0000004c, 5'd15, 27'h000001f5, 5'd27, 27'h0000034a, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003f5, 5'd22, 27'h0000021e, 5'd9, 27'h00000308, 32'h00000400,
  1'd1,  5'd18, 27'h00000217, 5'd25, 27'h00000338, 5'd16, 27'h000001cc, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000ad, 5'd22, 27'h0000007c, 5'd28, 27'h000001c5, 32'h00000400,
  1'd1,  5'd25, 27'h000003f2, 5'd2, 27'h000002ff, 5'd7, 27'h000003aa, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c7, 5'd4, 27'h000001f9, 5'd17, 27'h0000002f, 32'h00000400,
  1'd1,  5'd28, 27'h00000099, 5'd3, 27'h0000001d, 5'd26, 27'h0000031f, 32'hfffffc00,
  1'd1,  5'd26, 27'h000002e5, 5'd12, 27'h000001eb, 5'd9, 27'h00000004, 32'h00000400,
  1'd1,  5'd29, 27'h00000034, 5'd11, 27'h0000022b, 5'd16, 27'h000000a1, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000036b, 5'd15, 27'h0000010c, 5'd28, 27'h00000266, 32'h00000400,
  1'd1,  5'd26, 27'h00000011, 5'd21, 27'h000000ee, 5'd7, 27'h000001d0, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000027c, 5'd25, 27'h000002eb, 5'd16, 27'h000001a4, 32'h00000400,
  1'd1,  5'd27, 27'h00000080, 5'd23, 27'h00000381, 5'd29, 27'h000002fd, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000053, 5'd9, 27'h0000028e, 5'd3, 27'h00000221, 32'h00000400,
  1'd1,  5'd8, 27'h000000b7, 5'd9, 27'h00000255, 5'd12, 27'h00000352, 32'hfffffc00,
  1'd1,  5'd6, 27'h000003b6, 5'd10, 27'h000000cd, 5'd24, 27'h00000248, 32'h00000400,
  1'd1,  5'd8, 27'h00000051, 5'd19, 27'h000000db, 5'd4, 27'h00000269, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000339, 5'd18, 27'h0000004a, 5'd11, 27'h000003b1, 32'h00000400,
  1'd1,  5'd6, 27'h00000308, 5'd15, 27'h00000207, 5'd20, 27'h000002f6, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000395, 5'd28, 27'h0000011d, 5'd5, 27'h0000007f, 32'h00000400,
  1'd1,  5'd7, 27'h0000021e, 5'd26, 27'h000002fa, 5'd15, 27'h0000013e, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000011d, 5'd30, 27'h00000194, 5'd23, 27'h000001a6, 32'h00000400,
  1'd1,  5'd17, 27'h000003f2, 5'd9, 27'h000001bd, 5'd1, 27'h00000261, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003be, 5'd9, 27'h00000280, 5'd15, 27'h00000187, 32'h00000400,
  1'd1,  5'd17, 27'h0000036e, 5'd7, 27'h00000082, 5'd22, 27'h000001ec, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000001b, 5'd20, 27'h0000020a, 5'd2, 27'h0000024a, 32'h00000400,
  1'd1,  5'd17, 27'h0000024a, 5'd16, 27'h000003f4, 5'd13, 27'h000002ed, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000007f, 5'd19, 27'h0000008e, 5'd25, 27'h00000332, 32'h00000400,
  1'd1,  5'd18, 27'h0000019a, 5'd28, 27'h000002e4, 5'd3, 27'h000002c1, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000078, 5'd28, 27'h0000009b, 5'd14, 27'h00000309, 32'h00000400,
  1'd1,  5'd16, 27'h000000f8, 5'd30, 27'h000002e9, 5'd25, 27'h00000276, 32'hfffffc00,
  1'd1,  5'd30, 27'h000000a7, 5'd10, 27'h00000074, 5'd1, 27'h00000084, 32'h00000400,
  1'd1,  5'd27, 27'h0000038f, 5'd6, 27'h00000181, 5'd13, 27'h000003d9, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000030d, 5'd6, 27'h00000047, 5'd24, 27'h000000dd, 32'h00000400,
  1'd1,  5'd25, 27'h000003e4, 5'd15, 27'h000003f4, 5'd3, 27'h000001f2, 32'hfffffc00,
  1'd1,  5'd30, 27'h000002f9, 5'd16, 27'h000002c9, 5'd11, 27'h000003b0, 32'h00000400,
  1'd1,  5'd29, 27'h0000018d, 5'd18, 27'h0000035c, 5'd24, 27'h00000024, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003de, 5'd26, 27'h000002b2, 5'd1, 27'h000003dd, 32'h00000400,
  1'd1,  5'd29, 27'h0000023e, 5'd29, 27'h00000342, 5'd10, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000077, 5'd25, 27'h000003cf, 5'd20, 27'h00000342, 32'h00000400,
  1'd1,  5'd7, 27'h00000321, 5'd6, 27'h000002fa, 5'd9, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000007c, 5'd10, 27'h000000f2, 5'd27, 27'h0000025d, 32'h00000400,
  1'd1,  5'd8, 27'h000003e5, 5'd16, 27'h00000252, 5'd7, 27'h0000001a, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000377, 5'd17, 27'h000002e8, 5'd17, 27'h000002c4, 32'h00000400,
  1'd1,  5'd9, 27'h000001bf, 5'd18, 27'h00000190, 5'd30, 27'h00000111, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000280, 5'd30, 27'h0000010b, 5'd9, 27'h000003fd, 32'h00000400,
  1'd1,  5'd9, 27'h000003dd, 5'd29, 27'h000000f4, 5'd16, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000305, 5'd30, 27'h0000017e, 5'd30, 27'h00000201, 32'h00000400,
  1'd1,  5'd18, 27'h0000031b, 5'd6, 27'h0000008a, 5'd8, 27'h0000000c, 32'hfffffc00,
  1'd1,  5'd19, 27'h000000d1, 5'd10, 27'h000000f9, 5'd17, 27'h0000001d, 32'h00000400,
  1'd1,  5'd16, 27'h00000382, 5'd6, 27'h00000143, 5'd25, 27'h00000356, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000160, 5'd19, 27'h00000289, 5'd5, 27'h00000231, 32'h00000400,
  1'd1,  5'd20, 27'h000000c2, 5'd19, 27'h00000302, 5'd18, 27'h0000000e, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000027a, 5'd18, 27'h00000194, 5'd27, 27'h00000356, 32'h00000400,
  1'd1,  5'd16, 27'h0000018c, 5'd26, 27'h000003b9, 5'd7, 27'h00000236, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000338, 5'd28, 27'h000001bf, 5'd20, 27'h000000ea, 32'h00000400,
  1'd1,  5'd19, 27'h00000345, 5'd28, 27'h0000010b, 5'd26, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000262, 5'd8, 27'h00000117, 5'd8, 27'h000003b3, 32'h00000400,
  1'd1,  5'd30, 27'h00000105, 5'd8, 27'h000002fe, 5'd16, 27'h000002c7, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000256, 5'd9, 27'h000003b8, 5'd28, 27'h0000026a, 32'h00000400,
  1'd1,  5'd26, 27'h0000037e, 5'd17, 27'h000003c9, 5'd7, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000069, 5'd20, 27'h0000026a, 5'd20, 27'h000000b9, 32'h00000400,
  1'd1,  5'd30, 27'h000002c1, 5'd18, 27'h000003f5, 5'd26, 27'h00000350, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000ae, 5'd27, 27'h0000038b, 5'd7, 27'h000000b7, 32'h00000400,
  1'd1,  5'd28, 27'h000000ba, 5'd28, 27'h000000dd, 5'd18, 27'h00000379, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000033f, 5'd28, 27'h000000c4, 5'd26, 27'h0000026e, 32'h00000400,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd2, 27'h000002fa, 5'd2, 27'h0000010a, 5'd1, 27'h0000025d, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000228, 5'd1, 27'h0000021a, 5'd13, 27'h00000222, 32'h00000400,
  1'd1,  5'd3, 27'h0000019c, 5'd3, 27'h0000019f, 5'd23, 27'h00000147, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000006c, 5'd12, 27'h000000d7, 5'd2, 27'h00000130, 32'h00000400,
  1'd1,  5'd1, 27'h0000030b, 5'd13, 27'h00000036, 5'd23, 27'h000002d5, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000007a, 5'd24, 27'h000000f6, 5'd4, 27'h000002d4, 32'h00000400,
  1'd1,  5'd0, 27'h000001b1, 5'd22, 27'h0000015f, 5'd10, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000018f, 5'd21, 27'h0000037e, 5'd24, 27'h0000013f, 32'h00000400,
  1'd1,  5'd11, 27'h0000001f, 5'd4, 27'h000003b2, 5'd3, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000163, 5'd3, 27'h000002c8, 5'd13, 27'h000000af, 32'h00000400,
  1'd1,  5'd10, 27'h00000351, 5'd4, 27'h00000138, 5'd23, 27'h00000129, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000f2, 5'd14, 27'h000002f9, 5'd4, 27'h00000134, 32'h00000400,
  1'd1,  5'd14, 27'h00000053, 5'd11, 27'h000000a5, 5'd22, 27'h000002b1, 32'hfffffc00,
  1'd1,  5'd15, 27'h000001ae, 5'd24, 27'h00000370, 5'd0, 27'h000000bf, 32'h00000400,
  1'd1,  5'd12, 27'h00000353, 5'd23, 27'h000001cf, 5'd11, 27'h000000b8, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001a6, 5'd23, 27'h00000201, 5'd21, 27'h00000226, 32'h00000400,
  1'd1,  5'd24, 27'h000003d4, 5'd1, 27'h000002ae, 5'd1, 27'h00000016, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000086, 5'd1, 27'h00000083, 5'd12, 27'h0000028f, 32'h00000400,
  1'd1,  5'd25, 27'h000001fa, 5'd3, 27'h00000391, 5'd23, 27'h0000007d, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000019, 5'd11, 27'h00000282, 5'd1, 27'h000002a5, 32'h00000400,
  1'd1,  5'd21, 27'h000000f2, 5'd11, 27'h000001c8, 5'd11, 27'h00000170, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000261, 5'd13, 27'h0000009b, 5'd24, 27'h0000037b, 32'h00000400,
  1'd1,  5'd21, 27'h00000024, 5'd24, 27'h00000358, 5'd1, 27'h00000282, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000025f, 5'd23, 27'h000000d7, 5'd12, 27'h00000276, 32'h00000400,
  1'd1,  5'd22, 27'h000003d7, 5'd23, 27'h00000228, 5'd23, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000005b, 5'd2, 27'h0000029c, 5'd7, 27'h00000074, 32'h00000400,
  1'd1,  5'd1, 27'h000002fd, 5'd1, 27'h000002f1, 5'd18, 27'h00000259, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000036e, 5'd0, 27'h000001d8, 5'd28, 27'h00000113, 32'h00000400,
  1'd1,  5'd2, 27'h000003af, 5'd13, 27'h00000070, 5'd5, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd2, 27'h0000036b, 5'd13, 27'h00000034, 5'd18, 27'h00000039, 32'h00000400,
  1'd1,  5'd1, 27'h000001e1, 5'd12, 27'h0000017a, 5'd28, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000181, 5'd21, 27'h00000134, 5'd8, 27'h00000385, 32'h00000400,
  1'd1,  5'd2, 27'h000003b7, 5'd22, 27'h0000021a, 5'd20, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd0, 27'h000000e9, 5'd23, 27'h0000028a, 5'd29, 27'h0000033c, 32'h00000400,
  1'd1,  5'd11, 27'h00000277, 5'd0, 27'h000000c2, 5'd8, 27'h00000267, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000018a, 5'd1, 27'h0000039d, 5'd17, 27'h0000029a, 32'h00000400,
  1'd1,  5'd11, 27'h00000040, 5'd0, 27'h000003f5, 5'd29, 27'h00000251, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000296, 5'd10, 27'h0000027f, 5'd7, 27'h00000288, 32'h00000400,
  1'd1,  5'd14, 27'h00000318, 5'd11, 27'h00000311, 5'd20, 27'h00000026, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000025c, 5'd13, 27'h000001b9, 5'd26, 27'h00000008, 32'h00000400,
  1'd1,  5'd11, 27'h0000028f, 5'd21, 27'h00000314, 5'd7, 27'h00000160, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000188, 5'd21, 27'h00000054, 5'd17, 27'h000000af, 32'h00000400,
  1'd1,  5'd12, 27'h00000209, 5'd21, 27'h00000030, 5'd29, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000019d, 5'd1, 27'h00000183, 5'd8, 27'h00000082, 32'h00000400,
  1'd1,  5'd22, 27'h0000013a, 5'd2, 27'h0000023e, 5'd15, 27'h00000377, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000127, 5'd1, 27'h00000177, 5'd27, 27'h0000011b, 32'h00000400,
  1'd1,  5'd23, 27'h000000e5, 5'd13, 27'h0000019d, 5'd6, 27'h00000007, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000035e, 5'd14, 27'h00000376, 5'd16, 27'h0000016f, 32'h00000400,
  1'd1,  5'd24, 27'h000000ef, 5'd13, 27'h0000026f, 5'd27, 27'h000001aa, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000319, 5'd25, 27'h000002e0, 5'd5, 27'h000001f7, 32'h00000400,
  1'd1,  5'd21, 27'h000001b5, 5'd24, 27'h000002ba, 5'd19, 27'h0000020d, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000007c, 5'd24, 27'h00000345, 5'd28, 27'h000000e9, 32'h00000400,
  1'd1,  5'd1, 27'h000001ba, 5'd9, 27'h000001a7, 5'd1, 27'h000002cb, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000395, 5'd6, 27'h00000300, 5'd12, 27'h00000344, 32'h00000400,
  1'd1,  5'd3, 27'h00000357, 5'd5, 27'h0000037f, 5'd25, 27'h0000014c, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001c0, 5'd16, 27'h0000001c, 5'd3, 27'h00000165, 32'h00000400,
  1'd1,  5'd0, 27'h00000321, 5'd20, 27'h00000060, 5'd14, 27'h000001eb, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000326, 5'd19, 27'h00000241, 5'd23, 27'h0000026b, 32'h00000400,
  1'd1,  5'd2, 27'h000003b1, 5'd27, 27'h000001a3, 5'd3, 27'h00000316, 32'hfffffc00,
  1'd1,  5'd3, 27'h000000e6, 5'd28, 27'h0000011b, 5'd14, 27'h00000217, 32'h00000400,
  1'd1,  5'd0, 27'h000003b8, 5'd30, 27'h00000247, 5'd24, 27'h000003c0, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000006a, 5'd6, 27'h000001da, 5'd0, 27'h000003c5, 32'h00000400,
  1'd1,  5'd11, 27'h000001c4, 5'd7, 27'h000003d9, 5'd14, 27'h00000355, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000013, 5'd9, 27'h00000369, 5'd24, 27'h000001d7, 32'h00000400,
  1'd1,  5'd11, 27'h000000f0, 5'd19, 27'h00000039, 5'd0, 27'h000003f8, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000f7, 5'd18, 27'h00000146, 5'd12, 27'h0000005a, 32'h00000400,
  1'd1,  5'd12, 27'h0000012b, 5'd17, 27'h00000107, 5'd21, 27'h000001e0, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000083, 5'd30, 27'h0000039d, 5'd3, 27'h000000c3, 32'h00000400,
  1'd1,  5'd12, 27'h000001df, 5'd30, 27'h000001df, 5'd12, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000024f, 5'd29, 27'h0000034d, 5'd21, 27'h000000b7, 32'h00000400,
  1'd1,  5'd23, 27'h000003d1, 5'd9, 27'h00000329, 5'd1, 27'h0000035e, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000aa, 5'd7, 27'h000001df, 5'd13, 27'h000003f7, 32'h00000400,
  1'd1,  5'd23, 27'h000000b6, 5'd17, 27'h000002d4, 5'd1, 27'h00000279, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000095, 5'd19, 27'h000000ea, 5'd11, 27'h000000c4, 32'h00000400,
  1'd1,  5'd20, 27'h000003b7, 5'd18, 27'h000000b8, 5'd20, 27'h000002b9, 32'hfffffc00,
  1'd1,  5'd23, 27'h000002b2, 5'd29, 27'h00000158, 5'd1, 27'h000000dc, 32'h00000400,
  1'd1,  5'd21, 27'h000002df, 5'd27, 27'h000001a5, 5'd12, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000316, 5'd30, 27'h0000028d, 5'd20, 27'h000003e7, 32'h00000400,
  1'd1,  5'd4, 27'h0000020c, 5'd8, 27'h000000b6, 5'd5, 27'h0000028d, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000024f, 5'd5, 27'h0000010d, 5'd17, 27'h000002ce, 32'h00000400,
  1'd1,  5'd4, 27'h00000012, 5'd7, 27'h00000215, 5'd27, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002e, 5'd16, 27'h000001dc, 5'd9, 27'h00000119, 32'h00000400,
  1'd1,  5'd5, 27'h0000007f, 5'd17, 27'h00000003, 5'd15, 27'h000003b2, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000002d, 5'd19, 27'h000003b3, 5'd28, 27'h00000177, 32'h00000400,
  1'd1,  5'd2, 27'h00000074, 5'd28, 27'h000002dc, 5'd5, 27'h0000024f, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000256, 5'd29, 27'h00000385, 5'd16, 27'h00000259, 32'h00000400,
  1'd1,  5'd1, 27'h0000022f, 5'd25, 27'h000003a1, 5'd25, 27'h00000397, 32'hfffffc00,
  1'd1,  5'd12, 27'h000001d2, 5'd10, 27'h00000032, 5'd7, 27'h0000038e, 32'h00000400,
  1'd1,  5'd12, 27'h00000208, 5'd7, 27'h000000ac, 5'd20, 27'h000000c4, 32'hfffffc00,
  1'd1,  5'd10, 27'h000001ec, 5'd9, 27'h00000104, 5'd28, 27'h000002d8, 32'h00000400,
  1'd1,  5'd14, 27'h00000372, 5'd18, 27'h0000021c, 5'd7, 27'h000001bf, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000271, 5'd16, 27'h00000357, 5'd19, 27'h00000188, 32'h00000400,
  1'd1,  5'd11, 27'h000002b3, 5'd19, 27'h0000004d, 5'd26, 27'h000000b7, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000218, 5'd26, 27'h00000021, 5'd10, 27'h0000012b, 32'h00000400,
  1'd1,  5'd11, 27'h00000012, 5'd30, 27'h000003eb, 5'd15, 27'h00000246, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000006e, 5'd28, 27'h000002b3, 5'd28, 27'h00000340, 32'h00000400,
  1'd1,  5'd20, 27'h00000375, 5'd8, 27'h0000015d, 5'd6, 27'h000003cf, 32'hfffffc00,
  1'd1,  5'd23, 27'h000000e1, 5'd8, 27'h0000015e, 5'd17, 27'h00000187, 32'h00000400,
  1'd1,  5'd22, 27'h000002a6, 5'd8, 27'h000002e8, 5'd26, 27'h0000022b, 32'hfffffc00,
  1'd1,  5'd23, 27'h0000026f, 5'd15, 27'h00000235, 5'd8, 27'h000003a4, 32'h00000400,
  1'd1,  5'd22, 27'h000000ac, 5'd16, 27'h000001da, 5'd20, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000043, 5'd18, 27'h000001e8, 5'd29, 27'h00000306, 32'h00000400,
  1'd1,  5'd25, 27'h0000027f, 5'd27, 27'h00000321, 5'd8, 27'h00000324, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000084, 5'd29, 27'h00000349, 5'd17, 27'h00000253, 32'h00000400,
  1'd1,  5'd24, 27'h00000169, 5'd26, 27'h00000282, 5'd30, 27'h00000211, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000021d, 5'd2, 27'h00000394, 5'd6, 27'h00000063, 32'h00000400,
  1'd1,  5'd6, 27'h00000302, 5'd4, 27'h00000119, 5'd19, 27'h0000019e, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000033e, 5'd1, 27'h00000279, 5'd27, 27'h00000028, 32'h00000400,
  1'd1,  5'd5, 27'h000002d4, 5'd13, 27'h00000038, 5'd0, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000272, 5'd11, 27'h00000323, 5'd12, 27'h000003b3, 32'h00000400,
  1'd1,  5'd8, 27'h00000048, 5'd14, 27'h000001d0, 5'd21, 27'h00000106, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000048, 5'd25, 27'h00000105, 5'd3, 27'h00000283, 32'h00000400,
  1'd1,  5'd5, 27'h0000023e, 5'd24, 27'h00000023, 5'd12, 27'h0000004f, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003b6, 5'd24, 27'h000000e4, 5'd21, 27'h000003b3, 32'h00000400,
  1'd1,  5'd19, 27'h000002c4, 5'd1, 27'h0000014a, 5'd5, 27'h00000372, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000316, 5'd0, 27'h0000015d, 5'd19, 27'h00000037, 32'h00000400,
  1'd1,  5'd18, 27'h000003ae, 5'd0, 27'h000000b9, 5'd29, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000003a, 5'd13, 27'h000003d7, 5'd1, 27'h0000030f, 32'h00000400,
  1'd1,  5'd20, 27'h000001eb, 5'd10, 27'h00000315, 5'd22, 27'h000001ac, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003a4, 5'd22, 27'h000000bd, 5'd5, 27'h00000009, 32'h00000400,
  1'd1,  5'd17, 27'h00000143, 5'd21, 27'h0000036e, 5'd12, 27'h00000124, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001ac, 5'd22, 27'h0000034c, 5'd23, 27'h00000073, 32'h00000400,
  1'd1,  5'd30, 27'h0000017e, 5'd1, 27'h00000326, 5'd3, 27'h00000266, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000036e, 5'd3, 27'h0000009b, 5'd14, 27'h0000008d, 32'h00000400,
  1'd1,  5'd29, 27'h000001e6, 5'd2, 27'h00000056, 5'd24, 27'h000003d5, 32'hfffffc00,
  1'd1,  5'd26, 27'h000001c6, 5'd15, 27'h000000ce, 5'd3, 27'h0000035e, 32'h00000400,
  1'd1,  5'd29, 27'h00000137, 5'd14, 27'h00000052, 5'd13, 27'h000002df, 32'hfffffc00,
  1'd1,  5'd26, 27'h0000005a, 5'd11, 27'h000001ed, 5'd22, 27'h000001ff, 32'h00000400,
  1'd1,  5'd26, 27'h00000399, 5'd22, 27'h00000042, 5'd0, 27'h00000039, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000135, 5'd21, 27'h00000206, 5'd13, 27'h0000015b, 32'h00000400,
  1'd1,  5'd28, 27'h000002ce, 5'd22, 27'h000001a4, 5'd25, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000034, 5'd5, 27'h00000053, 5'd2, 27'h00000272, 32'h00000400,
  1'd1,  5'd7, 27'h0000009e, 5'd4, 27'h000002e5, 5'd15, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000031e, 5'd1, 27'h00000225, 5'd24, 27'h00000319, 32'h00000400,
  1'd1,  5'd5, 27'h00000369, 5'd11, 27'h000000b0, 5'd5, 27'h000001cd, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000037d, 5'd11, 27'h00000253, 5'd18, 27'h00000071, 32'h00000400,
  1'd1,  5'd8, 27'h000001e1, 5'd12, 27'h00000071, 5'd28, 27'h000003ae, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000108, 5'd23, 27'h0000036e, 5'd10, 27'h00000013, 32'h00000400,
  1'd1,  5'd6, 27'h00000257, 5'd21, 27'h00000219, 5'd16, 27'h00000196, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001a5, 5'd21, 27'h00000217, 5'd29, 27'h000001d8, 32'h00000400,
  1'd1,  5'd19, 27'h00000243, 5'd4, 27'h0000022b, 5'd2, 27'h000003d4, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001f8, 5'd2, 27'h00000347, 5'd14, 27'h0000012e, 32'h00000400,
  1'd1,  5'd17, 27'h0000006c, 5'd12, 27'h00000025, 5'd6, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000346, 5'd14, 27'h00000374, 5'd20, 27'h0000000c, 32'h00000400,
  1'd1,  5'd20, 27'h000001b3, 5'd12, 27'h000001e4, 5'd30, 27'h00000308, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000011b, 5'd21, 27'h0000004f, 5'd6, 27'h00000299, 32'h00000400,
  1'd1,  5'd16, 27'h000001df, 5'd22, 27'h000001a4, 5'd20, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000399, 5'd24, 27'h0000028a, 5'd28, 27'h00000237, 32'h00000400,
  1'd1,  5'd29, 27'h00000298, 5'd4, 27'h0000031e, 5'd7, 27'h00000226, 32'hfffffc00,
  1'd1,  5'd29, 27'h0000007c, 5'd2, 27'h0000004d, 5'd30, 27'h000002a7, 32'h00000400,
  1'd1,  5'd27, 27'h0000027a, 5'd11, 27'h000001fd, 5'd7, 27'h00000047, 32'hfffffc00,
  1'd1,  5'd27, 27'h000000c1, 5'd15, 27'h000000b6, 5'd15, 27'h00000278, 32'h00000400,
  1'd1,  5'd26, 27'h000001a0, 5'd14, 27'h000003ba, 5'd28, 27'h00000132, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003ef, 5'd24, 27'h00000391, 5'd10, 27'h000000aa, 32'h00000400,
  1'd1,  5'd27, 27'h000001e5, 5'd25, 27'h00000183, 5'd19, 27'h00000012, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000009b, 5'd23, 27'h00000276, 5'd26, 27'h000002c6, 32'h00000400,
  1'd1,  5'd5, 27'h000001b0, 5'd8, 27'h0000013e, 5'd4, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd9, 27'h000003eb, 5'd5, 27'h00000347, 5'd10, 27'h000001bb, 32'h00000400,
  1'd1,  5'd9, 27'h0000025d, 5'd9, 27'h00000061, 5'd25, 27'h000002ab, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001e5, 5'd18, 27'h000001a9, 5'd2, 27'h0000034c, 32'h00000400,
  1'd1,  5'd7, 27'h0000016c, 5'd17, 27'h000003bd, 5'd15, 27'h00000096, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001ee, 5'd17, 27'h000002cf, 5'd22, 27'h0000030b, 32'h00000400,
  1'd1,  5'd5, 27'h000000c7, 5'd25, 27'h000003f6, 5'd5, 27'h00000033, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000283, 5'd26, 27'h000000fe, 5'd10, 27'h00000229, 32'h00000400,
  1'd1,  5'd5, 27'h00000323, 5'd30, 27'h00000368, 5'd23, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000036a, 5'd9, 27'h000003cc, 5'd2, 27'h00000329, 32'h00000400,
  1'd1,  5'd18, 27'h00000299, 5'd9, 27'h000003be, 5'd14, 27'h00000354, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000114, 5'd6, 27'h000001a4, 5'd20, 27'h000002e4, 32'h00000400,
  1'd1,  5'd20, 27'h000001f5, 5'd19, 27'h0000019e, 5'd2, 27'h0000025a, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000dc, 5'd19, 27'h0000021c, 5'd12, 27'h00000261, 32'h00000400,
  1'd1,  5'd18, 27'h0000013c, 5'd19, 27'h00000172, 5'd22, 27'h0000002e, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002c3, 5'd27, 27'h00000097, 5'd3, 27'h0000026b, 32'h00000400,
  1'd1,  5'd16, 27'h0000020c, 5'd26, 27'h0000001f, 5'd14, 27'h0000000b, 32'hfffffc00,
  1'd1,  5'd18, 27'h000003bf, 5'd28, 27'h000000c6, 5'd21, 27'h000000fa, 32'h00000400,
  1'd1,  5'd25, 27'h00000370, 5'd7, 27'h0000005b, 5'd1, 27'h0000023e, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000015b, 5'd5, 27'h000000d3, 5'd15, 27'h000000bf, 32'h00000400,
  1'd1,  5'd26, 27'h000002e3, 5'd5, 27'h000000bd, 5'd23, 27'h00000357, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000dd, 5'd18, 27'h00000148, 5'd2, 27'h00000115, 32'h00000400,
  1'd1,  5'd28, 27'h000001c0, 5'd19, 27'h00000347, 5'd14, 27'h00000131, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002bc, 5'd17, 27'h00000085, 5'd25, 27'h00000336, 32'h00000400,
  1'd1,  5'd29, 27'h00000290, 5'd29, 27'h000000d0, 5'd4, 27'h0000005d, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000140, 5'd30, 27'h0000020f, 5'd12, 27'h000002eb, 32'h00000400,
  1'd1,  5'd30, 27'h000001ce, 5'd27, 27'h00000274, 5'd22, 27'h0000027d, 32'hfffffc00,
  1'd1,  5'd9, 27'h0000035e, 5'd6, 27'h00000056, 5'd5, 27'h000000dd, 32'h00000400,
  1'd1,  5'd8, 27'h00000010, 5'd5, 27'h000003a8, 5'd28, 27'h00000375, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000131, 5'd18, 27'h0000020e, 5'd5, 27'h000002d7, 32'h00000400,
  1'd1,  5'd8, 27'h0000003a, 5'd16, 27'h000000e4, 5'd20, 27'h00000227, 32'hfffffc00,
  1'd1,  5'd7, 27'h000001df, 5'd15, 27'h000003a8, 5'd29, 27'h0000003e, 32'h00000400,
  1'd1,  5'd8, 27'h0000015d, 5'd28, 27'h000001c3, 5'd7, 27'h0000021d, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000142, 5'd30, 27'h000002e8, 5'd19, 27'h0000003a, 32'h00000400,
  1'd1,  5'd5, 27'h00000370, 5'd27, 27'h00000327, 5'd26, 27'h000002ee, 32'hfffffc00,
  1'd1,  5'd18, 27'h000001ae, 5'd8, 27'h0000015d, 5'd8, 27'h000003c8, 32'h00000400,
  1'd1,  5'd16, 27'h000003c2, 5'd10, 27'h00000067, 5'd16, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000021d, 5'd7, 27'h000003ac, 5'd29, 27'h0000005a, 32'h00000400,
  1'd1,  5'd19, 27'h0000021b, 5'd17, 27'h0000007c, 5'd6, 27'h000001f7, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000005d, 5'd17, 27'h0000006c, 5'd18, 27'h0000005c, 32'h00000400,
  1'd1,  5'd15, 27'h000003eb, 5'd17, 27'h000000a4, 5'd30, 27'h0000039c, 32'hfffffc00,
  1'd1,  5'd16, 27'h000003fc, 5'd30, 27'h00000212, 5'd9, 27'h00000368, 32'h00000400,
  1'd1,  5'd16, 27'h00000307, 5'd27, 27'h000003c0, 5'd16, 27'h000001d7, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002be, 5'd26, 27'h000000f3, 5'd30, 27'h0000006a, 32'h00000400,
  1'd1,  5'd28, 27'h000000bd, 5'd7, 27'h000000a1, 5'd9, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd25, 27'h000003cc, 5'd6, 27'h00000370, 5'd19, 27'h000003a6, 32'h00000400,
  1'd1,  5'd29, 27'h000003e2, 5'd7, 27'h000003cf, 5'd27, 27'h00000219, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000169, 5'd17, 27'h0000007b, 5'd9, 27'h000003fc, 32'h00000400,
  1'd1,  5'd27, 27'h000002eb, 5'd17, 27'h00000262, 5'd19, 27'h00000181, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000346, 5'd17, 27'h00000182, 5'd26, 27'h0000017d, 32'h00000400,
  1'd1,  5'd25, 27'h00000383, 5'd27, 27'h00000300, 5'd9, 27'h000002aa, 32'hfffffc00,
  1'd1,  5'd28, 27'h000003c1, 5'd27, 27'h00000032, 5'd18, 27'h0000018e, 32'h00000400,
  1'd1,  5'd29, 27'h00000070, 5'd27, 27'h00000373, 5'd26, 27'h00000087, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd5, 27'h000000a4, 5'd4, 27'h0000019d, 5'd3, 27'h0000011c, 32'h00000400,
  1'd1,  5'd4, 27'h00000255, 5'd2, 27'h0000036d, 5'd10, 27'h0000030f, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000037f, 5'd4, 27'h000000a8, 5'd25, 27'h00000327, 32'h00000400,
  1'd1,  5'd1, 27'h000002c6, 5'd12, 27'h00000077, 5'd3, 27'h00000097, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000050, 5'd12, 27'h00000304, 5'd21, 27'h0000022a, 32'h00000400,
  1'd1,  5'd3, 27'h000001af, 5'd22, 27'h0000019e, 5'd4, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd4, 27'h000001d0, 5'd21, 27'h000003cb, 5'd12, 27'h000002b3, 32'h00000400,
  1'd1,  5'd3, 27'h000002e7, 5'd23, 27'h000000d4, 5'd25, 27'h00000057, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001f6, 5'd0, 27'h0000026f, 5'd4, 27'h000002e9, 32'h00000400,
  1'd1,  5'd13, 27'h00000309, 5'd3, 27'h000001f7, 5'd12, 27'h00000271, 32'hfffffc00,
  1'd1,  5'd11, 27'h0000026b, 5'd0, 27'h000000c6, 5'd21, 27'h000002e9, 32'h00000400,
  1'd1,  5'd13, 27'h00000399, 5'd12, 27'h0000022b, 5'd1, 27'h000003e3, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000024a, 5'd13, 27'h00000260, 5'd20, 27'h000003ac, 32'h00000400,
  1'd1,  5'd10, 27'h000001dc, 5'd24, 27'h000000be, 5'd1, 27'h000003a3, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000011b, 5'd23, 27'h0000035a, 5'd15, 27'h00000076, 32'h00000400,
  1'd1,  5'd13, 27'h000002d9, 5'd21, 27'h0000034d, 5'd21, 27'h000000be, 32'hfffffc00,
  1'd1,  5'd20, 27'h000002d2, 5'd1, 27'h00000202, 5'd0, 27'h00000148, 32'h00000400,
  1'd1,  5'd21, 27'h000000d4, 5'd2, 27'h0000012d, 5'd12, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000083, 5'd3, 27'h00000122, 5'd23, 27'h00000038, 32'h00000400,
  1'd1,  5'd22, 27'h000002b2, 5'd12, 27'h00000364, 5'd0, 27'h0000031e, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000380, 5'd14, 27'h00000127, 5'd13, 27'h0000009f, 32'h00000400,
  1'd1,  5'd25, 27'h00000041, 5'd12, 27'h00000134, 5'd23, 27'h0000035f, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002ce, 5'd23, 27'h00000166, 5'd0, 27'h000003c5, 32'h00000400,
  1'd1,  5'd20, 27'h000003be, 5'd24, 27'h000000c9, 5'd10, 27'h000002b7, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000195, 5'd25, 27'h00000160, 5'd25, 27'h00000173, 32'h00000400,
  1'd1,  5'd3, 27'h00000143, 5'd1, 27'h00000130, 5'd5, 27'h00000296, 32'hfffffc00,
  1'd1,  5'd3, 27'h000002fd, 5'd0, 27'h0000021b, 5'd17, 27'h000003ee, 32'h00000400,
  1'd1,  5'd1, 27'h0000006a, 5'd2, 27'h000003d6, 5'd29, 27'h000002ca, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001ec, 5'd13, 27'h00000186, 5'd9, 27'h00000035, 32'h00000400,
  1'd1,  5'd4, 27'h000001a2, 5'd12, 27'h00000005, 5'd18, 27'h00000305, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000371, 5'd13, 27'h0000030d, 5'd29, 27'h000001e9, 32'h00000400,
  1'd1,  5'd2, 27'h00000278, 5'd25, 27'h0000009b, 5'd7, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000089, 5'd21, 27'h00000049, 5'd16, 27'h00000312, 32'h00000400,
  1'd1,  5'd0, 27'h0000024f, 5'd22, 27'h00000163, 5'd27, 27'h000001ab, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003eb, 5'd2, 27'h000003c2, 5'd8, 27'h00000063, 32'h00000400,
  1'd1,  5'd10, 27'h00000340, 5'd1, 27'h000001e6, 5'd20, 27'h000001e5, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000158, 5'd0, 27'h00000025, 5'd28, 27'h00000195, 32'h00000400,
  1'd1,  5'd14, 27'h000001a4, 5'd12, 27'h00000367, 5'd8, 27'h000003b1, 32'hfffffc00,
  1'd1,  5'd13, 27'h000001bb, 5'd13, 27'h000002f1, 5'd20, 27'h000002a0, 32'h00000400,
  1'd1,  5'd12, 27'h000000ca, 5'd15, 27'h0000001f, 5'd26, 27'h000002c8, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000182, 5'd20, 27'h0000035d, 5'd6, 27'h00000093, 32'h00000400,
  1'd1,  5'd11, 27'h00000197, 5'd24, 27'h000001e2, 5'd18, 27'h00000225, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000019c, 5'd22, 27'h00000192, 5'd29, 27'h000001ea, 32'h00000400,
  1'd1,  5'd21, 27'h00000256, 5'd4, 27'h00000138, 5'd5, 27'h000003d0, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000376, 5'd2, 27'h000002cc, 5'd16, 27'h0000026c, 32'h00000400,
  1'd1,  5'd25, 27'h0000014a, 5'd1, 27'h000002f0, 5'd26, 27'h00000337, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000083, 5'd14, 27'h00000099, 5'd10, 27'h0000006e, 32'h00000400,
  1'd1,  5'd25, 27'h000001ad, 5'd12, 27'h0000028b, 5'd20, 27'h00000127, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002a5, 5'd10, 27'h00000170, 5'd27, 27'h00000279, 32'h00000400,
  1'd1,  5'd24, 27'h00000113, 5'd22, 27'h00000209, 5'd9, 27'h0000024e, 32'hfffffc00,
  1'd1,  5'd21, 27'h000002e8, 5'd24, 27'h000003df, 5'd17, 27'h00000057, 32'h00000400,
  1'd1,  5'd22, 27'h0000030f, 5'd24, 27'h00000312, 5'd27, 27'h0000026b, 32'hfffffc00,
  1'd1,  5'd1, 27'h000002aa, 5'd7, 27'h00000211, 5'd2, 27'h000000dc, 32'h00000400,
  1'd1,  5'd3, 27'h00000037, 5'd6, 27'h0000024f, 5'd14, 27'h00000172, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000136, 5'd7, 27'h000003d7, 5'd21, 27'h0000021b, 32'h00000400,
  1'd1,  5'd3, 27'h000003b0, 5'd19, 27'h00000257, 5'd3, 27'h0000017e, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000015d, 5'd18, 27'h0000006d, 5'd10, 27'h000002a4, 32'h00000400,
  1'd1,  5'd1, 27'h0000002b, 5'd19, 27'h0000032e, 5'd21, 27'h000002c9, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000130, 5'd25, 27'h000003c1, 5'd4, 27'h00000115, 32'h00000400,
  1'd1,  5'd4, 27'h00000365, 5'd30, 27'h000001b9, 5'd14, 27'h00000121, 32'hfffffc00,
  1'd1,  5'd4, 27'h0000001c, 5'd28, 27'h000003d1, 5'd24, 27'h0000009e, 32'h00000400,
  1'd1,  5'd13, 27'h0000009d, 5'd10, 27'h00000107, 5'd0, 27'h0000026d, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000001f, 5'd9, 27'h0000011b, 5'd10, 27'h00000194, 32'h00000400,
  1'd1,  5'd13, 27'h0000038e, 5'd7, 27'h0000012f, 5'd24, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd11, 27'h000003f6, 5'd18, 27'h000002ab, 5'd0, 27'h000000d5, 32'h00000400,
  1'd1,  5'd13, 27'h00000334, 5'd16, 27'h00000270, 5'd15, 27'h000001e4, 32'hfffffc00,
  1'd1,  5'd14, 27'h0000026a, 5'd15, 27'h0000020f, 5'd22, 27'h00000060, 32'h00000400,
  1'd1,  5'd15, 27'h0000019a, 5'd30, 27'h000001b8, 5'd3, 27'h000002f1, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000082, 5'd27, 27'h00000215, 5'd13, 27'h0000014f, 32'h00000400,
  1'd1,  5'd13, 27'h0000013a, 5'd27, 27'h00000368, 5'd25, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000017f, 5'd5, 27'h000001cf, 5'd1, 27'h0000006f, 32'h00000400,
  1'd1,  5'd23, 27'h0000013e, 5'd7, 27'h000003f2, 5'd13, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000060, 5'd18, 27'h00000383, 5'd1, 27'h000002b8, 32'h00000400,
  1'd1,  5'd23, 27'h00000111, 5'd18, 27'h000002ba, 5'd12, 27'h0000030a, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000350, 5'd20, 27'h0000002a, 5'd22, 27'h00000298, 32'h00000400,
  1'd1,  5'd22, 27'h00000290, 5'd28, 27'h0000032e, 5'd0, 27'h000003a0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001f7, 5'd29, 27'h000002dc, 5'd14, 27'h000000ff, 32'h00000400,
  1'd1,  5'd21, 27'h000000c8, 5'd29, 27'h000000ef, 5'd24, 27'h000002ff, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000007e, 5'd8, 27'h000001a8, 5'd15, 27'h000002a3, 32'h00000400,
  1'd1,  5'd4, 27'h00000097, 5'd8, 27'h00000320, 5'd30, 27'h00000165, 32'hfffffc00,
  1'd1,  5'd0, 27'h000002cb, 5'd18, 27'h000001b3, 5'd8, 27'h00000055, 32'h00000400,
  1'd1,  5'd0, 27'h000000ee, 5'd16, 27'h0000000a, 5'd18, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd2, 27'h000000c4, 5'd18, 27'h00000039, 5'd27, 27'h000000d9, 32'h00000400,
  1'd1,  5'd2, 27'h0000022d, 5'd29, 27'h0000018b, 5'd6, 27'h0000018a, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000391, 5'd29, 27'h00000191, 5'd18, 27'h00000081, 32'h00000400,
  1'd1,  5'd2, 27'h000002b1, 5'd26, 27'h00000380, 5'd30, 27'h0000005b, 32'hfffffc00,
  1'd1,  5'd10, 27'h0000025d, 5'd5, 27'h000003f0, 5'd5, 27'h00000309, 32'h00000400,
  1'd1,  5'd12, 27'h0000016d, 5'd5, 27'h00000206, 5'd15, 27'h000003a9, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000107, 5'd6, 27'h000000a5, 5'd27, 27'h00000211, 32'h00000400,
  1'd1,  5'd13, 27'h000001bf, 5'd16, 27'h000000c2, 5'd6, 27'h00000328, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000115, 5'd17, 27'h000001ae, 5'd16, 27'h000003c6, 32'h00000400,
  1'd1,  5'd11, 27'h00000007, 5'd19, 27'h00000244, 5'd26, 27'h0000037a, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000319, 5'd27, 27'h00000121, 5'd8, 27'h000002f2, 32'h00000400,
  1'd1,  5'd10, 27'h000003f4, 5'd29, 27'h00000085, 5'd19, 27'h00000070, 32'hfffffc00,
  1'd1,  5'd11, 27'h000000c1, 5'd30, 27'h0000007a, 5'd28, 27'h000003b8, 32'h00000400,
  1'd1,  5'd24, 27'h000002ee, 5'd8, 27'h00000102, 5'd5, 27'h0000033f, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000391, 5'd5, 27'h000003c7, 5'd18, 27'h00000351, 32'h00000400,
  1'd1,  5'd21, 27'h000003f3, 5'd6, 27'h000001e8, 5'd29, 27'h00000134, 32'hfffffc00,
  1'd1,  5'd21, 27'h00000233, 5'd16, 27'h000002c9, 5'd8, 27'h000002f4, 32'h00000400,
  1'd1,  5'd23, 27'h00000299, 5'd18, 27'h0000009e, 5'd15, 27'h000002f9, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000023a, 5'd19, 27'h000000e3, 5'd29, 27'h000003ca, 32'h00000400,
  1'd1,  5'd22, 27'h000003a5, 5'd25, 27'h000003e3, 5'd10, 27'h000000a4, 32'hfffffc00,
  1'd1,  5'd22, 27'h000000be, 5'd30, 27'h0000021d, 5'd16, 27'h0000036a, 32'h00000400,
  1'd1,  5'd25, 27'h00000167, 5'd27, 27'h00000114, 5'd28, 27'h00000062, 32'hfffffc00,
  1'd1,  5'd8, 27'h000002d8, 5'd4, 27'h0000030e, 5'd8, 27'h0000010b, 32'h00000400,
  1'd1,  5'd6, 27'h000000c8, 5'd4, 27'h00000330, 5'd18, 27'h000000ea, 32'hfffffc00,
  1'd1,  5'd7, 27'h000000cc, 5'd3, 27'h000003c1, 5'd30, 27'h000001a4, 32'h00000400,
  1'd1,  5'd5, 27'h000003df, 5'd15, 27'h000000b5, 5'd1, 27'h00000224, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000029a, 5'd14, 27'h000001be, 5'd13, 27'h00000355, 32'h00000400,
  1'd1,  5'd5, 27'h00000386, 5'd15, 27'h00000167, 5'd21, 27'h00000027, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000028, 5'd24, 27'h00000145, 5'd3, 27'h000001ec, 32'h00000400,
  1'd1,  5'd6, 27'h00000142, 5'd21, 27'h00000282, 5'd12, 27'h00000182, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000023a, 5'd23, 27'h00000195, 5'd21, 27'h000003f6, 32'h00000400,
  1'd1,  5'd18, 27'h0000034e, 5'd3, 27'h000002ce, 5'd7, 27'h0000014b, 32'hfffffc00,
  1'd1,  5'd15, 27'h0000028c, 5'd3, 27'h00000347, 5'd20, 27'h0000000c, 32'h00000400,
  1'd1,  5'd18, 27'h0000017e, 5'd1, 27'h0000025d, 5'd28, 27'h00000302, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000024, 5'd13, 27'h0000035f, 5'd0, 27'h00000335, 32'h00000400,
  1'd1,  5'd20, 27'h00000217, 5'd10, 27'h0000036d, 5'd23, 27'h00000384, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000103, 5'd22, 27'h000001fc, 5'd1, 27'h00000384, 32'h00000400,
  1'd1,  5'd19, 27'h000001dc, 5'd23, 27'h000002ad, 5'd11, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000007d, 5'd22, 27'h000003ea, 5'd20, 27'h00000342, 32'h00000400,
  1'd1,  5'd30, 27'h000000e0, 5'd2, 27'h00000266, 5'd0, 27'h00000263, 32'hfffffc00,
  1'd1,  5'd27, 27'h00000340, 5'd0, 27'h000001a6, 5'd13, 27'h000002c6, 32'h00000400,
  1'd1,  5'd26, 27'h0000008f, 5'd0, 27'h00000137, 5'd21, 27'h00000208, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000302, 5'd15, 27'h000001cc, 5'd3, 27'h000002c1, 32'h00000400,
  1'd1,  5'd29, 27'h000002ef, 5'd12, 27'h00000301, 5'd13, 27'h0000004c, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000035b, 5'd13, 27'h00000264, 5'd20, 27'h0000033d, 32'h00000400,
  1'd1,  5'd27, 27'h00000005, 5'd23, 27'h00000202, 5'd4, 27'h000003fb, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000009e, 5'd21, 27'h00000226, 5'd15, 27'h0000010d, 32'h00000400,
  1'd1,  5'd28, 27'h00000010, 5'd22, 27'h000000aa, 5'd24, 27'h0000009a, 32'hfffffc00,
  1'd1,  5'd8, 27'h000003fc, 5'd0, 27'h00000308, 5'd3, 27'h0000037c, 32'h00000400,
  1'd1,  5'd10, 27'h0000006c, 5'd5, 27'h00000096, 5'd15, 27'h0000016f, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000398, 5'd2, 27'h0000006e, 5'd21, 27'h00000233, 32'h00000400,
  1'd1,  5'd6, 27'h0000020f, 5'd10, 27'h00000208, 5'd5, 27'h00000232, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000186, 5'd12, 27'h00000237, 5'd15, 27'h00000296, 32'h00000400,
  1'd1,  5'd9, 27'h0000036f, 5'd12, 27'h000001e7, 5'd26, 27'h00000231, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000161, 5'd23, 27'h00000095, 5'd8, 27'h00000295, 32'h00000400,
  1'd1,  5'd5, 27'h0000023c, 5'd22, 27'h000000d8, 5'd16, 27'h00000205, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001c1, 5'd21, 27'h000003ff, 5'd30, 27'h000001e2, 32'h00000400,
  1'd1,  5'd17, 27'h0000016c, 5'd0, 27'h000002ac, 5'd4, 27'h0000008e, 32'hfffffc00,
  1'd1,  5'd18, 27'h0000037e, 5'd0, 27'h00000143, 5'd13, 27'h00000131, 32'h00000400,
  1'd1,  5'd15, 27'h000002f9, 5'd13, 27'h00000099, 5'd9, 27'h00000387, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e9, 5'd13, 27'h000000ca, 5'd16, 27'h000003c7, 32'h00000400,
  1'd1,  5'd19, 27'h0000025c, 5'd12, 27'h000001d5, 5'd26, 27'h000002a7, 32'hfffffc00,
  1'd1,  5'd17, 27'h00000135, 5'd23, 27'h00000190, 5'd8, 27'h000003fc, 32'h00000400,
  1'd1,  5'd18, 27'h00000051, 5'd23, 27'h000000e4, 5'd20, 27'h00000113, 32'hfffffc00,
  1'd1,  5'd17, 27'h0000012a, 5'd21, 27'h000003a2, 5'd28, 27'h00000150, 32'h00000400,
  1'd1,  5'd28, 27'h00000289, 5'd0, 27'h0000028c, 5'd7, 27'h000003ab, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000290, 5'd3, 27'h000002a7, 5'd27, 27'h0000036a, 32'h00000400,
  1'd1,  5'd25, 27'h00000356, 5'd12, 27'h000001c6, 5'd9, 27'h00000139, 32'hfffffc00,
  1'd1,  5'd30, 27'h000003b3, 5'd13, 27'h00000189, 5'd15, 27'h00000229, 32'h00000400,
  1'd1,  5'd30, 27'h00000070, 5'd10, 27'h000003f6, 5'd30, 27'h00000386, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000031e, 5'd24, 27'h0000034d, 5'd8, 27'h0000038a, 32'h00000400,
  1'd1,  5'd27, 27'h000002cf, 5'd21, 27'h00000117, 5'd16, 27'h00000391, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000165, 5'd21, 27'h000000a2, 5'd28, 27'h0000013b, 32'h00000400,
  1'd1,  5'd7, 27'h000003f9, 5'd8, 27'h00000149, 5'd3, 27'h00000321, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000e6, 5'd7, 27'h000003e7, 5'd13, 27'h0000013f, 32'h00000400,
  1'd1,  5'd9, 27'h00000024, 5'd9, 27'h000002ac, 5'd22, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd10, 27'h000000c6, 5'd19, 27'h00000373, 5'd3, 27'h00000292, 32'h00000400,
  1'd1,  5'd6, 27'h000003c1, 5'd18, 27'h00000093, 5'd10, 27'h00000235, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000217, 5'd20, 27'h000002a6, 5'd21, 27'h00000291, 32'h00000400,
  1'd1,  5'd5, 27'h00000376, 5'd30, 27'h000000a6, 5'd1, 27'h0000013f, 32'hfffffc00,
  1'd1,  5'd6, 27'h00000054, 5'd26, 27'h000000a8, 5'd13, 27'h00000343, 32'h00000400,
  1'd1,  5'd8, 27'h00000355, 5'd27, 27'h0000016e, 5'd23, 27'h00000290, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001d4, 5'd9, 27'h000003a1, 5'd2, 27'h00000088, 32'h00000400,
  1'd1,  5'd15, 27'h000002d9, 5'd6, 27'h00000089, 5'd10, 27'h0000021f, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000239, 5'd9, 27'h0000037f, 5'd24, 27'h000001f5, 32'h00000400,
  1'd1,  5'd16, 27'h000001c3, 5'd16, 27'h00000126, 5'd2, 27'h000003a2, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000189, 5'd15, 27'h000003e8, 5'd12, 27'h0000015e, 32'h00000400,
  1'd1,  5'd16, 27'h000002da, 5'd20, 27'h000002a0, 5'd21, 27'h000002f0, 32'hfffffc00,
  1'd1,  5'd18, 27'h000002c4, 5'd26, 27'h000003f0, 5'd4, 27'h00000067, 32'h00000400,
  1'd1,  5'd20, 27'h00000155, 5'd29, 27'h000000cc, 5'd13, 27'h000002a4, 32'hfffffc00,
  1'd1,  5'd16, 27'h000001e3, 5'd30, 27'h0000001d, 5'd22, 27'h00000114, 32'h00000400,
  1'd1,  5'd27, 27'h000002f9, 5'd6, 27'h0000025d, 5'd4, 27'h000000a2, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000035, 5'd5, 27'h000002eb, 5'd13, 27'h00000159, 32'h00000400,
  1'd1,  5'd28, 27'h0000033b, 5'd7, 27'h00000232, 5'd25, 27'h000000f9, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003bb, 5'd18, 27'h00000243, 5'd4, 27'h00000131, 32'h00000400,
  1'd1,  5'd27, 27'h000003d9, 5'd18, 27'h000001fc, 5'd10, 27'h00000175, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000031c, 5'd18, 27'h00000019, 5'd23, 27'h0000035c, 32'h00000400,
  1'd1,  5'd28, 27'h000003d1, 5'd26, 27'h0000014b, 5'd1, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000021f, 5'd29, 27'h00000201, 5'd10, 27'h00000219, 32'h00000400,
  1'd1,  5'd30, 27'h0000009f, 5'd28, 27'h000003ad, 5'd23, 27'h000003ba, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000149, 5'd9, 27'h000000a5, 5'd9, 27'h0000015d, 32'h00000400,
  1'd1,  5'd7, 27'h000003f7, 5'd5, 27'h00000122, 5'd30, 27'h00000281, 32'hfffffc00,
  1'd1,  5'd10, 27'h00000106, 5'd20, 27'h00000230, 5'd5, 27'h000001f6, 32'h00000400,
  1'd1,  5'd9, 27'h00000229, 5'd20, 27'h00000034, 5'd15, 27'h0000027b, 32'hfffffc00,
  1'd1,  5'd6, 27'h0000013f, 5'd18, 27'h000003a7, 5'd27, 27'h000000a6, 32'h00000400,
  1'd1,  5'd6, 27'h00000027, 5'd26, 27'h000000b2, 5'd7, 27'h00000095, 32'hfffffc00,
  1'd1,  5'd8, 27'h000000d5, 5'd26, 27'h000003df, 5'd16, 27'h0000030d, 32'h00000400,
  1'd1,  5'd6, 27'h00000284, 5'd27, 27'h000001db, 5'd30, 27'h00000215, 32'hfffffc00,
  1'd1,  5'd19, 27'h00000070, 5'd5, 27'h000003f5, 5'd5, 27'h000001bb, 32'h00000400,
  1'd1,  5'd20, 27'h000002a3, 5'd7, 27'h00000298, 5'd18, 27'h000000aa, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000009d, 5'd10, 27'h000000c2, 5'd27, 27'h00000010, 32'h00000400,
  1'd1,  5'd18, 27'h00000033, 5'd19, 27'h00000012, 5'd7, 27'h000003cc, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000371, 5'd20, 27'h00000044, 5'd16, 27'h0000038b, 32'h00000400,
  1'd1,  5'd17, 27'h00000344, 5'd18, 27'h00000398, 5'd25, 27'h00000376, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000035e, 5'd29, 27'h00000213, 5'd5, 27'h000000fc, 32'h00000400,
  1'd1,  5'd19, 27'h000001fd, 5'd28, 27'h00000064, 5'd15, 27'h00000342, 32'hfffffc00,
  1'd1,  5'd17, 27'h000002c9, 5'd30, 27'h000000ce, 5'd26, 27'h0000028e, 32'h00000400,
  1'd1,  5'd26, 27'h0000001e, 5'd7, 27'h0000011d, 5'd8, 27'h000000b2, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000155, 5'd8, 27'h000002a5, 5'd16, 27'h00000201, 32'h00000400,
  1'd1,  5'd26, 27'h000002d6, 5'd7, 27'h000000ea, 5'd27, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002a9, 5'd20, 27'h0000010f, 5'd9, 27'h0000035f, 32'h00000400,
  1'd1,  5'd28, 27'h000002f6, 5'd17, 27'h000002ca, 5'd19, 27'h000002ef, 32'hfffffc00,
  1'd1,  5'd27, 27'h000001a7, 5'd15, 27'h000003ca, 5'd30, 27'h000002bf, 32'h00000400,
  1'd1,  5'd26, 27'h000002aa, 5'd29, 27'h00000026, 5'd7, 27'h00000212, 32'hfffffc00,
  1'd1,  5'd29, 27'h00000106, 5'd27, 27'h0000019e, 5'd18, 27'h00000218, 32'h00000400,
  1'd1,  5'd29, 27'h0000037d, 5'd26, 27'h0000024b, 5'd26, 27'h00000054, 32'hfffffc00,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd0,  5'd0, 27'h00000000, 5'd0, 27'h00000000, 5'd0, 27'h00000000, 32'h00000000,
  1'd1,  5'd4, 27'h000000e6, 5'd3, 27'h000001da, 5'd2, 27'h00000327, 32'h00000400,
  1'd1,  5'd1, 27'h000002d1, 5'd4, 27'h0000024e, 5'd15, 27'h00000161, 32'hfffffc00,
  1'd1,  5'd4, 27'h00000024, 5'd3, 27'h0000038b, 5'd21, 27'h0000025c, 32'h00000400,
  1'd1,  5'd3, 27'h00000100, 5'd12, 27'h00000242, 5'd2, 27'h00000359, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000343, 5'd13, 27'h00000082, 5'd24, 27'h00000092, 32'h00000400,
  1'd1,  5'd1, 27'h00000143, 5'd21, 27'h00000091, 5'd1, 27'h00000365, 32'hfffffc00,
  1'd1,  5'd0, 27'h000001e9, 5'd25, 27'h000001d4, 5'd10, 27'h000003cb, 32'h00000400,
  1'd1,  5'd3, 27'h0000006d, 5'd25, 27'h00000175, 5'd23, 27'h000002bb, 32'hfffffc00,
  1'd1,  5'd13, 27'h00000077, 5'd0, 27'h000000f8, 5'd2, 27'h00000374, 32'h00000400,
  1'd1,  5'd10, 27'h0000024d, 5'd4, 27'h000002f0, 5'd14, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd14, 27'h000000b5, 5'd4, 27'h00000368, 5'd25, 27'h0000030f, 32'h00000400,
  1'd1,  5'd11, 27'h00000350, 5'd13, 27'h00000268, 5'd1, 27'h00000045, 32'hfffffc00,
  1'd1,  5'd13, 27'h0000013d, 5'd13, 27'h0000009e, 5'd23, 27'h00000013, 32'h00000400,
  1'd1,  5'd12, 27'h00000054, 5'd24, 27'h000000c0, 5'd3, 27'h000001ca, 32'hfffffc00,
  1'd1,  5'd12, 27'h000000f2, 5'd22, 27'h0000034e, 5'd11, 27'h0000008b, 32'h00000400,
  1'd1,  5'd13, 27'h000003de, 5'd23, 27'h000000c5, 5'd21, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000021c, 5'd3, 27'h0000000b, 5'd1, 27'h000001ba, 32'h00000400,
  1'd1,  5'd24, 27'h0000027e, 5'd5, 27'h0000001c, 5'd10, 27'h000001ce, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000016f, 5'd4, 27'h000000ef, 5'd21, 27'h00000049, 32'h00000400,
  1'd1,  5'd20, 27'h000002b3, 5'd12, 27'h0000026f, 5'd2, 27'h000000ef, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000257, 5'd13, 27'h0000019e, 5'd14, 27'h00000045, 32'h00000400,
  1'd1,  5'd24, 27'h0000012f, 5'd21, 27'h000000cc, 5'd0, 27'h00000241, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000039e, 5'd25, 27'h00000317, 5'd12, 27'h0000007a, 32'h00000400,
  1'd1,  5'd23, 27'h00000026, 5'd23, 27'h000001f6, 5'd21, 27'h0000002a, 32'hfffffc00,
  1'd1,  5'd3, 27'h0000019a, 5'd3, 27'h0000011e, 5'd6, 27'h0000031e, 32'h00000400,
  1'd1,  5'd4, 27'h00000283, 5'd4, 27'h00000130, 5'd16, 27'h000003db, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000017a, 5'd3, 27'h0000004a, 5'd27, 27'h00000317, 32'h00000400,
  1'd1,  5'd2, 27'h000003f6, 5'd12, 27'h00000216, 5'd7, 27'h000001f8, 32'hfffffc00,
  1'd1,  5'd0, 27'h0000017a, 5'd14, 27'h00000234, 5'd17, 27'h00000289, 32'h00000400,
  1'd1,  5'd3, 27'h000001c7, 5'd13, 27'h0000026b, 5'd30, 27'h0000017d, 32'hfffffc00,
  1'd1,  5'd2, 27'h00000364, 5'd21, 27'h00000209, 5'd9, 27'h0000029f, 32'h00000400,
  1'd1,  5'd3, 27'h000000ff, 5'd22, 27'h000003ea, 5'd18, 27'h00000360, 32'hfffffc00,
  1'd1,  5'd1, 27'h0000014a, 5'd23, 27'h00000399, 5'd28, 27'h0000025f, 32'h00000400,
  1'd1,  5'd10, 27'h00000327, 5'd4, 27'h000002e1, 5'd10, 27'h00000120, 32'hfffffc00,
  1'd1,  5'd11, 27'h00000349, 5'd4, 27'h00000324, 5'd19, 27'h000000f7, 32'h00000400,
  1'd1,  5'd13, 27'h000002e4, 5'd2, 27'h000001b2, 5'd30, 27'h00000385, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003c5, 5'd13, 27'h0000011a, 5'd5, 27'h000003ad, 32'h00000400,
  1'd1,  5'd10, 27'h0000039b, 5'd14, 27'h000002b0, 5'd19, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000ab, 5'd15, 27'h000000de, 5'd29, 27'h00000127, 32'h00000400,
  1'd1,  5'd14, 27'h00000273, 5'd24, 27'h0000014f, 5'd9, 27'h000003fd, 32'hfffffc00,
  1'd1,  5'd12, 27'h0000010b, 5'd21, 27'h00000036, 5'd19, 27'h00000162, 32'h00000400,
  1'd1,  5'd15, 27'h00000016, 5'd25, 27'h0000008f, 5'd28, 27'h000003c8, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000044, 5'd0, 27'h000003c9, 5'd6, 27'h00000087, 32'h00000400,
  1'd1,  5'd25, 27'h00000266, 5'd3, 27'h00000189, 5'd16, 27'h00000230, 32'hfffffc00,
  1'd1,  5'd21, 27'h000001c3, 5'd1, 27'h00000161, 5'd26, 27'h00000241, 32'h00000400,
  1'd1,  5'd21, 27'h00000149, 5'd13, 27'h000002dc, 5'd7, 27'h0000021b, 32'hfffffc00,
  1'd1,  5'd21, 27'h0000024c, 5'd14, 27'h00000265, 5'd18, 27'h00000238, 32'h00000400,
  1'd1,  5'd24, 27'h0000033c, 5'd15, 27'h00000030, 5'd29, 27'h000002b0, 32'hfffffc00,
  1'd1,  5'd24, 27'h000001d8, 5'd25, 27'h00000101, 5'd9, 27'h0000035c, 32'h00000400,
  1'd1,  5'd23, 27'h00000011, 5'd21, 27'h000002e7, 5'd17, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd22, 27'h0000037e, 5'd22, 27'h0000025b, 5'd28, 27'h00000378, 32'h00000400,
  1'd1,  5'd4, 27'h0000022b, 5'd6, 27'h0000017b, 5'd3, 27'h00000343, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000006, 5'd9, 27'h000002c7, 5'd13, 27'h000000bb, 32'h00000400,
  1'd1,  5'd5, 27'h00000048, 5'd5, 27'h000001b4, 5'd25, 27'h00000220, 32'hfffffc00,
  1'd1,  5'd2, 27'h000003ff, 5'd16, 27'h000000af, 5'd2, 27'h000000dc, 32'h00000400,
  1'd1,  5'd5, 27'h0000002a, 5'd20, 27'h0000013b, 5'd21, 27'h00000048, 32'hfffffc00,
  1'd1,  5'd0, 27'h00000093, 5'd29, 27'h00000346, 5'd3, 27'h0000013a, 32'h00000400,
  1'd1,  5'd1, 27'h000000ae, 5'd30, 27'h00000283, 5'd11, 27'h00000190, 32'hfffffc00,
  1'd1,  5'd3, 27'h000003bf, 5'd28, 27'h00000051, 5'd25, 27'h00000107, 32'h00000400,
  1'd1,  5'd10, 27'h00000196, 5'd8, 27'h00000079, 5'd3, 27'h0000003e, 32'hfffffc00,
  1'd1,  5'd15, 27'h000000b9, 5'd6, 27'h00000091, 5'd11, 27'h0000022e, 32'h00000400,
  1'd1,  5'd11, 27'h000001bf, 5'd5, 27'h0000039d, 5'd20, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000147, 5'd20, 27'h00000111, 5'd3, 27'h0000013d, 32'h00000400,
  1'd1,  5'd14, 27'h000000b8, 5'd16, 27'h0000015e, 5'd13, 27'h00000292, 32'hfffffc00,
  1'd1,  5'd13, 27'h000003ea, 5'd20, 27'h00000052, 5'd22, 27'h000002bc, 32'h00000400,
  1'd1,  5'd13, 27'h00000165, 5'd29, 27'h00000261, 5'd0, 27'h0000033d, 32'hfffffc00,
  1'd1,  5'd11, 27'h000001c9, 5'd27, 27'h0000039b, 5'd10, 27'h000001e1, 32'h00000400,
  1'd1,  5'd11, 27'h00000232, 5'd26, 27'h00000149, 5'd25, 27'h000002dd, 32'hfffffc00,
  1'd1,  5'd24, 27'h00000353, 5'd8, 27'h0000008c, 5'd2, 27'h0000029b, 32'h00000400,
  1'd1,  5'd23, 27'h0000008b, 5'd9, 27'h00000074, 5'd10, 27'h000001ed, 32'hfffffc00,
  1'd1,  5'd21, 27'h000000bd, 5'd17, 27'h00000373, 5'd2, 27'h0000034c, 32'h00000400,
  1'd1,  5'd24, 27'h000000c0, 5'd19, 27'h00000194, 5'd11, 27'h000001b1, 32'hfffffc00,
  1'd1,  5'd25, 27'h0000011c, 5'd18, 27'h00000044, 5'd21, 27'h00000263, 32'h00000400,
  1'd1,  5'd24, 27'h00000030, 5'd28, 27'h0000033e, 5'd2, 27'h0000020f, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000348, 5'd26, 27'h00000066, 5'd12, 27'h0000039b, 32'h00000400,
  1'd1,  5'd22, 27'h0000028d, 5'd30, 27'h000001da, 5'd25, 27'h00000239, 32'hfffffc00,
  1'd1,  5'd1, 27'h00000196, 5'd5, 27'h00000266, 5'd19, 27'h00000360, 32'h00000400,
  1'd1,  5'd3, 27'h0000012c, 5'd5, 27'h000000bb, 5'd30, 27'h00000206, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000008a, 5'd16, 27'h0000018a, 5'd9, 27'h00000297, 32'h00000400,
  1'd1,  5'd1, 27'h00000275, 5'd17, 27'h00000324, 5'd19, 27'h00000100, 32'hfffffc00,
  1'd1,  5'd3, 27'h00000018, 5'd19, 27'h0000026a, 5'd28, 27'h00000142, 32'h00000400,
  1'd1,  5'd0, 27'h0000038e, 5'd27, 27'h000001ed, 5'd7, 27'h000001c0, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000047, 5'd28, 27'h000003a5, 5'd20, 27'h0000010f, 32'h00000400,
  1'd1,  5'd0, 27'h00000011, 5'd30, 27'h000002a0, 5'd27, 27'h000000ff, 32'hfffffc00,
  1'd1,  5'd14, 27'h00000265, 5'd9, 27'h0000015b, 5'd6, 27'h000001c3, 32'h00000400,
  1'd1,  5'd15, 27'h000000a0, 5'd7, 27'h000000b8, 5'd16, 27'h0000009f, 32'hfffffc00,
  1'd1,  5'd14, 27'h000003da, 5'd6, 27'h0000036d, 5'd29, 27'h0000007c, 32'h00000400,
  1'd1,  5'd15, 27'h00000013, 5'd19, 27'h0000039a, 5'd7, 27'h00000064, 32'hfffffc00,
  1'd1,  5'd12, 27'h000003b6, 5'd19, 27'h00000366, 5'd17, 27'h0000020f, 32'h00000400,
  1'd1,  5'd11, 27'h000002a8, 5'd19, 27'h000003f3, 5'd26, 27'h00000216, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000286, 5'd30, 27'h00000026, 5'd5, 27'h0000023a, 32'h00000400,
  1'd1,  5'd13, 27'h000001a1, 5'd29, 27'h00000397, 5'd18, 27'h000002d7, 32'hfffffc00,
  1'd1,  5'd12, 27'h00000039, 5'd26, 27'h00000327, 5'd30, 27'h00000282, 32'h00000400,
  1'd1,  5'd25, 27'h000001e5, 5'd6, 27'h0000006f, 5'd8, 27'h00000183, 32'hfffffc00,
  1'd1,  5'd23, 27'h00000058, 5'd9, 27'h000000be, 5'd16, 27'h000003d4, 32'h00000400,
  1'd1,  5'd23, 27'h000001e5, 5'd8, 27'h00000372, 5'd28, 27'h000001bb, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000031, 5'd18, 27'h000002c1, 5'd8, 27'h00000084, 32'h00000400,
  1'd1,  5'd22, 27'h0000027c, 5'd16, 27'h0000013d, 5'd18, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd24, 27'h0000033e, 5'd20, 27'h0000007a, 5'd30, 27'h000000a6, 32'h00000400,
  1'd1,  5'd20, 27'h000003c0, 5'd28, 27'h0000003d, 5'd6, 27'h000001e9, 32'hfffffc00,
  1'd1,  5'd22, 27'h00000397, 5'd26, 27'h000000cd, 5'd17, 27'h00000342, 32'h00000400,
  1'd1,  5'd24, 27'h000002ba, 5'd28, 27'h0000013f, 5'd27, 27'h000001c3, 32'hfffffc00,
  1'd1,  5'd9, 27'h000000ca, 5'd3, 27'h0000028f, 5'd6, 27'h0000037f, 32'h00000400,
  1'd1,  5'd7, 27'h0000011d, 5'd1, 27'h0000036a, 5'd17, 27'h00000353, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000299, 5'd3, 27'h00000161, 5'd28, 27'h000003e0, 32'h00000400,
  1'd1,  5'd8, 27'h00000039, 5'd12, 27'h00000193, 5'd2, 27'h00000278, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000269, 5'd12, 27'h00000379, 5'd12, 27'h00000176, 32'h00000400,
  1'd1,  5'd6, 27'h000002c9, 5'd11, 27'h000002cc, 5'd23, 27'h000001a1, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000015f, 5'd22, 27'h0000037f, 5'd1, 27'h00000288, 32'h00000400,
  1'd1,  5'd9, 27'h00000079, 5'd21, 27'h00000102, 5'd10, 27'h0000037f, 32'hfffffc00,
  1'd1,  5'd5, 27'h0000032c, 5'd24, 27'h0000029b, 5'd23, 27'h000002ed, 32'h00000400,
  1'd1,  5'd18, 27'h000003c2, 5'd3, 27'h00000119, 5'd10, 27'h00000051, 32'hfffffc00,
  1'd1,  5'd17, 27'h000001b2, 5'd4, 27'h00000368, 5'd17, 27'h00000108, 32'h00000400,
  1'd1,  5'd18, 27'h000000ca, 5'd2, 27'h0000016c, 5'd30, 27'h000000e1, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000155, 5'd12, 27'h00000182, 5'd1, 27'h00000380, 32'h00000400,
  1'd1,  5'd17, 27'h00000269, 5'd11, 27'h0000032d, 5'd23, 27'h00000176, 32'hfffffc00,
  1'd1,  5'd16, 27'h000002c1, 5'd25, 27'h00000267, 5'd4, 27'h000002e5, 32'h00000400,
  1'd1,  5'd16, 27'h00000212, 5'd25, 27'h000000a3, 5'd11, 27'h000002f3, 32'hfffffc00,
  1'd1,  5'd19, 27'h000003e5, 5'd24, 27'h0000028f, 5'd25, 27'h00000163, 32'h00000400,
  1'd1,  5'd29, 27'h00000074, 5'd0, 27'h000003d5, 5'd4, 27'h0000009c, 32'hfffffc00,
  1'd1,  5'd27, 27'h000003f0, 5'd1, 27'h00000228, 5'd12, 27'h000003be, 32'h00000400,
  1'd1,  5'd29, 27'h0000023b, 5'd4, 27'h0000030c, 5'd21, 27'h00000323, 32'hfffffc00,
  1'd1,  5'd28, 27'h0000018d, 5'd13, 27'h0000004c, 5'd4, 27'h00000198, 32'h00000400,
  1'd1,  5'd29, 27'h0000037a, 5'd13, 27'h000003bb, 5'd10, 27'h000003ca, 32'hfffffc00,
  1'd1,  5'd28, 27'h000000ec, 5'd13, 27'h0000017f, 5'd24, 27'h00000335, 32'h00000400,
  1'd1,  5'd28, 27'h0000003d, 5'd24, 27'h00000061, 5'd2, 27'h00000207, 32'hfffffc00,
  1'd1,  5'd25, 27'h00000391, 5'd23, 27'h000000fa, 5'd12, 27'h00000163, 32'h00000400,
  1'd1,  5'd26, 27'h000003b8, 5'd25, 27'h00000158, 5'd24, 27'h00000017, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000180, 5'd4, 27'h00000083, 5'd2, 27'h0000025a, 32'h00000400,
  1'd1,  5'd7, 27'h000001c0, 5'd2, 27'h0000016b, 5'd12, 27'h000001d3, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000257, 5'd0, 27'h000003f3, 5'd21, 27'h0000038d, 32'h00000400,
  1'd1,  5'd7, 27'h0000003d, 5'd14, 27'h00000001, 5'd7, 27'h000002d4, 32'hfffffc00,
  1'd1,  5'd5, 27'h000001c8, 5'd10, 27'h000001a5, 5'd16, 27'h000000b7, 32'h00000400,
  1'd1,  5'd7, 27'h000001d2, 5'd14, 27'h000000c7, 5'd29, 27'h00000008, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002c1, 5'd21, 27'h00000129, 5'd5, 27'h0000036e, 32'h00000400,
  1'd1,  5'd9, 27'h000002ae, 5'd23, 27'h000003ca, 5'd17, 27'h0000011b, 32'hfffffc00,
  1'd1,  5'd8, 27'h00000375, 5'd24, 27'h0000033f, 5'd28, 27'h0000026c, 32'h00000400,
  1'd1,  5'd16, 27'h000001d2, 5'd1, 27'h000002b1, 5'd2, 27'h00000168, 32'hfffffc00,
  1'd1,  5'd18, 27'h000000ad, 5'd4, 27'h0000029a, 5'd10, 27'h0000031e, 32'h00000400,
  1'd1,  5'd18, 27'h000001c4, 5'd12, 27'h000002ae, 5'd8, 27'h00000000, 32'hfffffc00,
  1'd1,  5'd15, 27'h000003a5, 5'd10, 27'h00000385, 5'd19, 27'h00000123, 32'h00000400,
  1'd1,  5'd16, 27'h000003c1, 5'd11, 27'h00000035, 5'd27, 27'h000002b6, 32'hfffffc00,
  1'd1,  5'd16, 27'h00000174, 5'd21, 27'h00000058, 5'd9, 27'h000000a5, 32'h00000400,
  1'd1,  5'd19, 27'h000002d6, 5'd21, 27'h00000033, 5'd20, 27'h0000004e, 32'hfffffc00,
  1'd1,  5'd17, 27'h000000e9, 5'd21, 27'h00000333, 5'd27, 27'h000002b9, 32'h00000400,
  1'd1,  5'd29, 27'h0000008a, 5'd3, 27'h000002c8, 5'd9, 27'h00000371, 32'hfffffc00,
  1'd1,  5'd30, 27'h0000005a, 5'd4, 27'h0000038b, 5'd29, 27'h000003a5, 32'h00000400,
  1'd1,  5'd27, 27'h000003b5, 5'd15, 27'h000001c4, 5'd7, 27'h00000041, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000030, 5'd14, 27'h00000383, 5'd15, 27'h00000201, 32'h00000400,
  1'd1,  5'd26, 27'h000000c3, 5'd15, 27'h0000000e, 5'd26, 27'h000002fa, 32'hfffffc00,
  1'd1,  5'd26, 27'h000000b4, 5'd20, 27'h000002d0, 5'd6, 27'h000003c8, 32'h00000400,
  1'd1,  5'd30, 27'h000003f0, 5'd21, 27'h000003a8, 5'd16, 27'h000002f5, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002fe, 5'd25, 27'h0000023d, 5'd30, 27'h00000021, 32'h00000400,
  1'd1,  5'd7, 27'h000001c1, 5'd5, 27'h000002ce, 5'd3, 27'h0000034b, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000322, 5'd6, 27'h00000061, 5'd10, 27'h00000366, 32'h00000400,
  1'd1,  5'd8, 27'h000003a6, 5'd5, 27'h00000365, 5'd23, 27'h000002ec, 32'hfffffc00,
  1'd1,  5'd7, 27'h0000000c, 5'd18, 27'h00000119, 5'd3, 27'h000002f5, 32'h00000400,
  1'd1,  5'd5, 27'h0000013a, 5'd20, 27'h00000147, 5'd12, 27'h000000a3, 32'hfffffc00,
  1'd1,  5'd5, 27'h000002af, 5'd17, 27'h00000383, 5'd24, 27'h000003e1, 32'h00000400,
  1'd1,  5'd5, 27'h00000138, 5'd30, 27'h000003e3, 5'd3, 27'h000003e0, 32'hfffffc00,
  1'd1,  5'd9, 27'h00000161, 5'd30, 27'h000001e6, 5'd12, 27'h000003cd, 32'h00000400,
  1'd1,  5'd10, 27'h0000009e, 5'd29, 27'h000001b7, 5'd24, 27'h00000203, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000007e, 5'd5, 27'h000000f4, 5'd1, 27'h00000156, 32'h00000400,
  1'd1,  5'd17, 27'h000003df, 5'd8, 27'h00000084, 5'd15, 27'h00000061, 32'hfffffc00,
  1'd1,  5'd15, 27'h000002bd, 5'd7, 27'h000003a2, 5'd23, 27'h00000128, 32'h00000400,
  1'd1,  5'd16, 27'h0000004e, 5'd20, 27'h000001cb, 5'd4, 27'h00000295, 32'hfffffc00,
  1'd1,  5'd19, 27'h000001de, 5'd20, 27'h00000173, 5'd12, 27'h000003af, 32'h00000400,
  1'd1,  5'd17, 27'h0000002a, 5'd18, 27'h00000093, 5'd25, 27'h00000306, 32'hfffffc00,
  1'd1,  5'd17, 27'h000003e2, 5'd26, 27'h000003cb, 5'd4, 27'h000000df, 32'h00000400,
  1'd1,  5'd16, 27'h000003ce, 5'd29, 27'h0000036c, 5'd14, 27'h000000e6, 32'hfffffc00,
  1'd1,  5'd20, 27'h00000150, 5'd29, 27'h000002fa, 5'd24, 27'h0000023c, 32'h00000400,
  1'd1,  5'd28, 27'h00000141, 5'd7, 27'h00000065, 5'd2, 27'h00000265, 32'hfffffc00,
  1'd1,  5'd28, 27'h00000280, 5'd9, 27'h00000294, 5'd13, 27'h00000207, 32'h00000400,
  1'd1,  5'd29, 27'h000001d4, 5'd9, 27'h00000352, 5'd21, 27'h00000229, 32'hfffffc00,
  1'd1,  5'd27, 27'h0000015a, 5'd17, 27'h00000197, 5'd1, 27'h0000000b, 32'h00000400,
  1'd1,  5'd29, 27'h000000e6, 5'd16, 27'h000003f0, 5'd13, 27'h0000006e, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000338, 5'd16, 27'h000000ca, 5'd22, 27'h00000169, 32'h00000400,
  1'd1,  5'd27, 27'h0000009e, 5'd29, 27'h00000070, 5'd10, 27'h0000037d, 32'hfffffc00,
  1'd1,  5'd29, 27'h000002f4, 5'd27, 27'h00000279, 5'd21, 27'h000002af, 32'h00000400,
  1'd1,  5'd7, 27'h0000003b, 5'd5, 27'h0000012b, 5'd7, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd6, 27'h000001d9, 5'd8, 27'h00000184, 5'd27, 27'h0000005e, 32'h00000400,
  1'd1,  5'd8, 27'h000000e5, 5'd19, 27'h00000085, 5'd9, 27'h00000004, 32'hfffffc00,
  1'd1,  5'd8, 27'h0000021c, 5'd16, 27'h000001ba, 5'd17, 27'h0000035d, 32'h00000400,
  1'd1,  5'd8, 27'h00000312, 5'd19, 27'h000000ef, 5'd29, 27'h00000056, 32'hfffffc00,
  1'd1,  5'd7, 27'h00000388, 5'd26, 27'h00000040, 5'd7, 27'h000003ee, 32'h00000400,
  1'd1,  5'd7, 27'h000001d9, 5'd29, 27'h000002c1, 5'd19, 27'h00000313, 32'hfffffc00,
  1'd1,  5'd5, 27'h00000390, 5'd27, 27'h0000031a, 5'd29, 27'h000003ff, 32'h00000400,
  1'd1,  5'd16, 27'h000001d4, 5'd7, 27'h0000016f, 5'd9, 27'h00000077, 32'hfffffc00,
  1'd1,  5'd20, 27'h0000011b, 5'd8, 27'h0000009c, 5'd18, 27'h000002a5, 32'h00000400,
  1'd1,  5'd20, 27'h000000e7, 5'd6, 27'h000003cc, 5'd30, 27'h000003a1, 32'hfffffc00,
  1'd1,  5'd15, 27'h00000356, 5'd15, 27'h0000030e, 5'd9, 27'h000001fd, 32'h00000400,
  1'd1,  5'd18, 27'h000000cb, 5'd19, 27'h00000130, 5'd17, 27'h00000038, 32'hfffffc00,
  1'd1,  5'd19, 27'h000002d2, 5'd15, 27'h000002b3, 5'd26, 27'h000001ae, 32'h00000400,
  1'd1,  5'd18, 27'h00000138, 5'd29, 27'h00000062, 5'd5, 27'h00000136, 32'hfffffc00,
  1'd1,  5'd16, 27'h0000000e, 5'd27, 27'h000002e7, 5'd20, 27'h00000295, 32'h00000400,
  1'd1,  5'd17, 27'h0000013a, 5'd28, 27'h0000014d, 5'd27, 27'h00000179, 32'hfffffc00,
  1'd1,  5'd29, 27'h000003d8, 5'd10, 27'h000000eb, 5'd5, 27'h00000140, 32'h00000400,
  1'd1,  5'd26, 27'h000001c8, 5'd10, 27'h0000013d, 5'd18, 27'h0000015c, 32'hfffffc00,
  1'd1,  5'd28, 27'h000002a6, 5'd8, 27'h000000e6, 5'd29, 27'h000002b7, 32'h00000400,
  1'd1,  5'd29, 27'h000002bb, 5'd16, 27'h000003d0, 5'd8, 27'h00000289, 32'hfffffc00,
  1'd1,  5'd26, 27'h00000292, 5'd19, 27'h00000097, 5'd18, 27'h000003a0, 32'h00000400,
  1'd1,  5'd29, 27'h00000102, 5'd16, 27'h0000003d, 5'd27, 27'h0000008c, 32'hfffffc00,
  1'd1,  5'd30, 27'h000001a2, 5'd29, 27'h0000007d, 5'd9, 27'h0000014d, 32'h00000400,
  1'd1,  5'd27, 27'h0000037a, 5'd27, 27'h000001c9, 5'd16, 27'h0000023c, 32'hfffffc00,
  1'd1,  5'd30, 27'h00000262, 5'd28, 27'h000001b0, 5'd26, 27'h0000013d, 32'h00000400};
