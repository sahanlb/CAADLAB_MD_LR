-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
0U/op8AfrDbNdFggUUot6syEcZdwCnbnvKHMTW0TAKHIdnWaV5vk/uX8SobLgg4X
0XZlluvEzyUnQBVMA/xmx4zfmfrfnPKz9xnClsS9VTVpiPHfwVj0pa0YIZL3osxq
wvlU6pSc3ZTQxWW7LCXZ7ohfTtmtmtqagv6pCbWciw8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13232)
`protect data_block
O6xvFFJBvT/4t+s51b1kTT+ybYjyxMgSfnqdOX4eel/rwwVpgGFpXsJdJiEBSDWa
82S4fpO1Zjr27EefHuSPjYNKIPjxmP2g6BIT3QE2E0ifYj0BPh3S1+raPq99BWhs
2y/v91zsgB8UixD1sAcMPnSjNtRc1uUgFexK+tAHSXx3QNVlRIA/Rt2nwzead0BG
7qe400fHLxOuKw+AB2v83jm2QtgeyxoERbI/0AvxFnbgCvuXEG83wYmhMYJSPyWr
gHyQ4jyomya81CVNFKmLs3dYpodRkA5vsD05VdfiOFca2HDBr5VjF7gXiKX1tq56
jg9lJqIo/H/9E8Ftsmu9Tc6C9rEZwNXVoZ6fnp9P5GF3Z559B92pnRxE3c1nH8+X
e3cVNqx5VTrd66/SHUSjhGOpOQgSDFw+1tTkQnsM+Ix51TnZSIFuoesuT9hrl5r2
jdpExWjblZ5GjD69IBkLb6soSA0oN7jwQJ3PFQQxzm5p7DgeYvxUx1/XRqeUhBJG
xRd0faNwz72pq+im2qNUlEklzmSm/XjwDF5LmPaPSLcAxCGWoHwT8Fbaahqt3+az
zp617fRsmm9EHZXpkjHXYSZ26rtWwm7TcnZnQJg/K/7AtBBrTbi/3bA46xGXsmxZ
HtG4UcyJHD0p6AcWC6pP75LGh/aNmo3zrNBmol20/rVEzPRICcWvrwuTF6sqB98Q
4iIEsn6x7Mmech/iYTCCpHM2kq6tPdaUrUqFSadL8GGxcpRwViN0J5ntji6HHK10
bQWauxFtWFXBcCMXw9RZucu7eK78BV0uBkvONv0piLjQGKXBrK5UH/uGzcOP6A4b
3T3rwb+VSJuOoNkfRtewFXKjedZ9GO+DiO35htR/ok/Sbj37mmib9KDb3KUJ7HA9
a9QWkdoxjUAISQecXbL2NDxrGSmAc7xyhdeB95wQ6x9an192RXBUaCQFThTIl/Hd
YQfnaHfTWgQbDrUH0j935DsOs9LKWIuR2momLaNsGNzaObEq7+mn5I4vm4CiC4EH
lKUqgbmF4hF7KRHG71tNX8F2dA/t/ql/yuLxj0asNq5UOSDOEs7rnDJofNw8+wxk
fWpCfFzySozPE0LLisBhLfotC4gwa3D2lX7afxHe5th5otwRYI8Tm5DqUMj826AG
4alGxBxOtHwHUbPy4NaWNiWZuk7L1kosDYQ3RR/5GhBB8ZoO5S89J4Ou9c82kkjB
SnnT1oCHm/m020TS6f+pEsiimuKn7HPvBHnooLGxun6wHt5+t0xbUlPQeGzt1Y7Q
xu9+Z8L0h/qbbDVzxkitlwHPBAQ1koSK2FpE9eKEuc3L12mBMZrHUPPNFjFdJt8q
iYyNOiHfyKzvn4usms+x+q1u7Suakoderhj0vUeZzdk7N/ySKTOgEkHAQdLvFJx5
CZ7mmU5f1txhT+YxOzzupp0P3IlJulUMvQnNGsl0V6OGnBGWmMrL5eiMZCqylVZW
TA2B2ZdjaoqQqGwe4zx5PpWoyMSkwZYoEzdVqQ6ryIsgAM0TOewOEsTEEh59oycn
7dD9cvmL8uqA6At2GJ5bPTGCzik05kGb9otRCrv53mk8O3DxlN12MlvdHCn3r4Bx
dDi9nGfhIL6vxhZ5i8Phsw22oApgAFtVNazyFgEC2Y8pfJBZzMb17i/UdC5msj5y
SuWSB8g8ZnRfwSVZXyHzaux9ISzS3WJDFBPkEP9WcMGHiz3SoVJ7mt0hyh9x29OD
xsrKn9LEZCyhcq8OFinBnIdtNu8leKDWZIAeRPvKHCUR9CUEAT5EkvbPfYjRm5yd
GmHbNi2X9drDJ6o3TiWDvuhoDajVAZyoKz33775iifAG5CaUJLXbdknhtThz8Qqp
Hb4gUpVd+XpZZFFfTbit8jdHakj+9RbQ7mRfQjJnVsjECDgel1l4eO6iF0bVk9pH
x05GoP9jkpWakC7dVy4eaFOkdIyG2QaG8OZdYsYh/rDhtpPURCQElLw4qZyvhdL/
mkAu3iKm0cC1D0iLKKa3kUiWpz2v/wfEUgRLrzmuqxdZ+Sx+Sl/lNxLTIqgjCGj4
lqN3l00trZadBJrh0MEq17EucbKjfpVT78a/1fx4A40ISLUmaMmqsf/DIQebdvGw
g5sShe9YKQZcZGl08u/A6uz6lIX1jZPOfOGQCiyHKVsQtTbocawkd5+sGPsnH6b/
6H8V7T5s5x/3QqHcjzeViHId1ChaRVOuzBGM/MwwpHPu+tAlKY/cJa8JAD/X82jf
/vHiPZOjjs6SpMQ/5TzYqmwHAG0/9955E8ESv63h/kCdLUbSaZ3YcStwAnBRETih
3m6XsXPGL91P5l4TMR10cRe6ucnBRm0Tkgrn4usAEYlRVGVgryFA35Cv+0zJORGz
DfXucgh9+ttTrV2L1HQBFzZABV2wmFUwfRzraN3D/3W31dXm6MudQ28fh44S1FFx
IsSBnsOxli380AXa0JAcXqZi6yzGWxLmhmYhuwaRh3Xg/aU3jh9cLJXbs6EXBtro
kbPR+PCC/Nx/KVxqzK20OxyPHklRxqbIlaSCw4/QiVNSSYqh42cVuzQs4LYeg4A6
LMWMQ8NB2pKWZYOIzX35iN07GyncCX8GB90S6r/zKgHfAG5x38Xu4Htjmg2A7dAK
zDJChi4tq5idssRolU9yIfNoMB6B30jWRizAtvZ1nJh3IbMT7AR669n7KaTiyq/h
ipO06PcpcMrnRLhGKLVv9vZ6U5RtFMALQ64ZnAFkdduHS91TkN3o/ou+7fcx3tKH
nbIJKMA7lEPc/Occpx/GaneUj/Ijk+ElwNdGOzaAyQZFXpNFTteQA21BCvNvWU0J
0UsMKOVx6r4No5XZ6fox/WOaKJ85OvHYGZAc/c4O5WWOMOMbhcvUHg+sgye9UWDo
GurNS5XFyuqZYJUprvCpG/0Ryl96y/6zaE/0psGEmR5vd+s5O/ieZwuCbNu/z1g9
DYDST+2cGu42QznHzbTWMsNj6XFyKUDzdMS4MBGfejNmncSNlhbKkWvtqNTIZCKP
xKNHKV0RdXRRAenJ01EuXc1QvDodPG/409HRLT4TB80rwxTAk7hBFL6EarFXJNEL
7L9r3Axim9eWLnmwonSfMfSawnXWCgSng6dFUv6k6St3jPEkHTi4yTNVVqIhYQxf
GKClzqD91gAxZGx8RcvWEFOCKtRo+DKgY1eF+pzZTeUH7dLn0oaBw9GTuIW47sf2
7pXksu9PiyK8Az5G5UftGCUNqAj+8sh2mdBMOBTxsh3xxwaUWokRo1HQFryvRSf+
UZCz73JW+NbQ0osxP55OTtOsOa/X8F5+/m9wcnEepWccODyEecrzgMGBrFTJQ6cR
uHSqyS+iKmQPuv0FWFUm7fOCKnKqRn9TC/RiXlOWgmlRgiQRQlVNu65m+ufZit/K
gdab1TwcdVs47gcVMMwo+po0Y01xclER5a4oSFILzDbDoRPc6BEw3kQtu5VrJbkV
ALoVRgpXUNqmS8pta0KlCjHpcxcsT4A/3+/JAT7A0xDNMPwgTOIBRm00IxcpbSVg
AwG/SR1IroRBvj/gJ6ToVVV4MtNy7t1PGFUCsX1JhUiUQ53Zf3sao7HCDPdgAsCg
GKwl9g2L+sJBsZwEbFqZObUJCfIwvztvF4eYdLUWXURV4cMryg6XtVFVfVa4PevW
wy8tuJkq5CmrlD/HfCd2GZkUDja0cjsz0Jd6OhcLpAvjjIucpVc6Dr4bgk728yds
0jBx75riN2XqteeVtlGi8hMZWZwZtvosnkOh7NX9Sh9w3dL3YK1T2e0DdfrorcmC
xZSnAsqPyjkPVUnfNAKH0/GPhxamUJG/2X3GLjBpvvg23YUe6aYkp7FkKwVg9hd5
S3tbOXxcjkn1ILVDIBwymcSf15PMn+lIP3D9yELAlCiy2UA4sGRc5NANNq8SNZZj
af8Ybaa4CTwhW6dRpHutUnwEzj1a+Xd/HTQ5cxllfVe6s0rAyl4MFtJRv03Ni3VP
S5GCs5dEalm9CaSUtlrQr9p+VchzoePtVL7YN6eaIBUqXGea4NIAR21Qs228NIlR
sCg8yFGwj4EGJVyz7dotvmwDIBozFdEyYGO/oZRlDU9GSZftMAkYvDgrXYvwb7pa
U8Nlxalvop40dSSoU2Dsk+DwUuNWh2yg3JUqWrqiLmq6Zen4Anz3bQ9WktON28Bz
r3ISK1QTPutbZtYRkVEetIzHpHwn6zCt6qwUaIZG0LK2KHYg58jJ8nqL+Gr4ieDD
PfDsyRLuFeSxaPvjKIzXCmUT+pnYIIeITbNi0BnbVScC6CJyJUIO1exg5sPs/bTJ
fm2tDCFQXXQqe/igLROZ4PB07Tlu6pBw+R3+OekjthpPbPydctOHqgDHubGC6iEV
RcQnO4J6rQ07Ipdgue1QPG+VVd9yPW9Q0khIwAfcUM0X+2JmNrm16BD36ak/PWga
9rIDTOrGdaMcR5PkyhpyvqbbrNhR07yL0dcRNBded7ufoK2AsGOKs6A4WaMlE1vX
fj0IjX1jjuqAWik4c2ciAVBVZ64Hg/+7rQtOAIxt6SPwnxBUA5HuIfzW8h4bIN1o
JWT/sr+uoURzTEUbMqaz9pa0j+f78USyEFJ90VI3Eh+HdXiViqpVRhyIQ4RYVQbN
IScNf9lFXIq48ioHYgawEO1phWp/99Gv4fo9Am2vqa/fcsfSg4ETiJbyBk2brGIw
JSCgltRnqa0Ep0ZHzRPt5pYYat4TZ+izRYMbJqjAyyWL1L8iWL1RnDctgr2XVR2G
3cSZbs+PwnENXCHE+6tKESFh3h08EZwpd4h+acfzfNHRAbM2erelZG/MibsGMNa3
PZrWwML6cvBc53v8gPyAmYoJUgtFlssu4GBr6Uv1HWkMmzB+rNSH4GGPxlNAiAt+
oPkqhc1w0u/xf1xFam/6P5aY4qkj/iVVjMpI/TtmH/C8YhKZSgTeqrVerW2+KSJf
eOZ3Hlx68qR2I01lK2J4YtCvTqfH3FNCYDwHId5sc3Sywezuw2qCyjxQ3AgdQsU0
WD2yBd6GKy82Yyvf7fKYQ7Z/hwZ12fVMh8iPZhXnRW/FYvG7QqvpKHewL+k5CcpI
STU2A6bPEQj39fCmOWzxrv+m0zArxRRuc3OSKFZaNhu4OMptOtZcqKuLkvxSZEE7
tTHNF6YJmJCZWQYky7VmoQyAzSjyJXjU8jutqZnKbdk5SGs6PG07cW9ahjdBLDXw
ADkhTTpMdfsPXZWNPlfk7UO4k3TwlNMGp4iu1eW0GHw3mSWNpKubNUv3H9UTtu9k
ic3MWzIH/MG4DHsF4Jin21CNjmdv0ycElbglB6Ap6sMExXxBVbQ7PuZ/Fpkcz60h
1asuPXYpbbCTmH+EfyWTBNJ+VsuWkDfcuVhDmAL36yyQYJ1vzUzesVIHZ7+nPD2e
7/cQFD3WijfjCow1F4ricg61lX8+Ne6vYPGMpjwgw1OLdIaAuTTmH1dxoXgOLDq4
PplU6Zp6I6AxmZsVOLaf3uJGTzKWKZ3L4gDKOZV7Zm92Rp2D4koSz9tHukKcOHtO
HiyfqHlkrZRCmQQM82vEHL6gckqQKos+pCs2cRtbXdo4VANSecoc7ARxc0K6M5DK
L/XtDWXsEpYiLqy6X4f1HicE+OBP7+ljbUTJB8h9ZVqWW/yzqKlRRHmy6ReIsmyt
JrR4ve52TentFvAs6rvuPOGzcy2FqBYJ6cAzY2T+auY+zm3KUv9IR61XUQ5Otsnj
EFbIML9X37BjududNeXZIBCsvJ8iYubXqz6g0BT7hjpfHV7bxjQ9EcWcCaK4Tuou
wp6R0av4WSvvDUXC823Inoo2Om0ys9DP0n5Z88S3MebiW4F781MIGwGjHJVK/7m5
RCYLoarTSSV0Nn9B9mIWymjZmrEakeQYu0EycKhrsIXf8YaX9lVb7UCw5aSo05J6
6ctXYHIKeNV/bXejCcIt4GrliQi1vmcoBPftsFeC4Oeyh10tc1bVFaruQmcxdCkh
j0Nxkl0pX7mfWwnnVrMIr+Lh4wWzonM7ocLcmHliro6/xUqQf6yoIzAHUuV4XUAb
30Oo8EIZYALUM+DXZHN403T0WBH7nlMpG10caSphKH720EzTpD/SCBVzj2gsRZ7o
IFuFNUZ+U/i7jQ54sfDhx9pP6L0uanF3jLKUqZQqwFEiyIAfnJUegK9Eb+GrHPcK
69o89IguBKBy8eRuoH/8J3SvOa9YZwvPxvjzL1qD6hyJVL6HwYPWCAQ0iMp9n/4g
3Q31iC2dhTUjTXuffVeqzPXih4z0tReYzmEdGFyQNyFQfa7EOXDMcv6QuTIxSTY2
mBJ31pJW4Qc2PTrcJFjJTYoMSnHtAbZvCp+ARBoLk3peB8vHaN7gAWl8nBRWU7N9
tD7Ewibe/+lA0nl5ajeEvQ+/D6KOtS7AMRNWa1xLQiJVZQ7HqUu62jkNntcBMisi
y8Vz3qwDKiWakKFIRypIo4Kn7EIX2E1AHpUQfrw3ZDsWtXhaz8RvwUzo+QeILXB6
920HiiiI1wlXciChWEOuLwnJpDHw8Mmm8dthyWEpeYTN1ZgyEvdiNGUfD6Lhph2S
WRgS02NkLtVNmO4g8HAyybjgJZGI48NberK9mtxNuf3d2LZe0VrUXaYW+V5DLIb5
wS8aCW5W+wh9zUQNOWXyimrWvYkKAYbLh1qPgKlh6iY9Nv+0NSWOjUedC7imk0oA
vWf6yKSLjrDs1/oJvhnj/T6KyKL1tjy4AF5zEvQarFx0efzRD4xU83CLpinKlpPb
3rQZFsVceeTd7VZQnZ/hPbRxroq4/imtuxXagC1nDQav85L2P+/Rv4ATCdFdcBpu
XdIm0NaMoZD73mRjoncjZSBStmDgUDlUklmlV7dyIXdDHDXqzbHMvja+yss4zNa7
t0eq7XbiDTILehXm1Ng//D6wwYcLU3ukeM9JGhn8wu70hS8u58F7Aky8sRPyJWrB
zwbpa2QkkP8HmDJbdK9jQTdLJVzVELzqi6IcRqoOGWDR+gIz7Ukpixc42AbJFdPQ
Y9McjPEG0w+Qpk4AQdrtrwsJwJNJ3JbabiFZoFdBzqE4Lm4Jsab2FtVDJ8Wpg/Ia
2p2sJnBx60EHnYg/bCFHJYQxb27NsbDIIYptV8jRnWQ0+wc1QNaPFo07iwZbR8AY
58sidwd7BUcKE7HKimm9bbnzZ5JYpxELVPrD07rNUDZ0UtVW9WdRqtQjMS0EVcxU
0M/K4B2j0CPY6FycfNiwXNLe/v+h2K6t/pKp8HLSidAGXdsIfGO9aaYuU7xFUzlp
H1xNEQ5UDruehj+n9FUc/MdPf/3nZI/LlsIwyDcIrGSYfi8BK8UuEKTn7r7bmlZt
05AOlXnCyTYbZK80nhmn1xFqe2VDSHpkyvz95fDcdA6d7tb7FU5wLxLnvwMS7uQs
guN5fWOA1PfL46XxpTW0V5Kftb0xTmOH9qRdLTycF/gPZlOl0h4Jm9sB8JJEcOJw
7gcLJdO7hsBH2HrB/3fSNhf4LHz1Xw6JWNjdY8ab4q15aHL22iZmq/RdGMRint0S
mrrQN/KFPE/C3scRdX+tTca4BXQYrVrO/MA2Qq9F0cE83BgGwGznxvtqM0v3VrxK
hajEzY2TfCDwAYXW3XYHFBuAkH9OTFY/BkG5lNtQbiTqOJYTP/BgRBHfx7h/j6jp
+4FTOUGQtbFWrWqoDN97GPz/k+t7f7iisy4or/LyjurXEWbCLewIp9yVVbr9Y1T9
BQbtZWIOPOS7ATa1pcF4mSG31X72eeF6huKEoC1yv13lUbLemTBeABMChMElbgeE
s8SBrXH0HRV8f4Wztga9gGO2wecq0fJsOXZ9Pdhko6AIAbnkg6Ok63IqjClLPmRC
S+9BhwBVasmV04VK1P/Pji11DaXclKCeCd3GchazYm82plDaP6WjX5H/pIXGy4y6
nbmuBS/SuP+9mQuHaGai3szeIWh6MW1pvTxp6mb5chDRiucEyHgAvgbLcLVWGh6+
TgD4sJltvFJFjpr2vufunkuwpm+GS9uRJ9Mp6g5rcg6ZxOC43qutfvReSSCbsiu8
wkJHPtxasRYNxdToZNZqlXGm/W56zQTlbq656SDszPXqwDhA0c8PZ9B5+9ZJb4Ov
gcEpxHs8C7XrxRTn4lUR3Ras5s55dui+3TCuOAPSn4fiTxep69sl3QzOLtYdcN/a
VFGZfdZC0He4GTqLP4kcGGnz1BpFUfcLN8x5Y2QyrooJ9nZzDlkEK1uPxPYhi0X0
GYffVBaQvGeQf0LoM2J1yxB+aRPHdx0zfmHdSrd/OpvKb4uirmU0snG3duuC9qFk
2/4Xr+l2mX1r1mcjtqMHui9Cq7IbxF2bjQV7HWRz+U9BUr63nvVkAhX54GPIqFXo
OAMo4AxfVT4ITJZI+unqdUPpcWYE+tFurokxr/8aex4eoGOoeKnZt1K69j7YZUiT
rhGeQP1soWbmOkHfP5IcRcCdtQhngVg/0dAG4flLCJgE20bRhwezSIpLZBWfBbaO
UbKFRcIRbKbLFH9jMNwTCBP81yHl81XQrKaM5LP0a9hcaMDi8r7NP9huZRhyAwIY
Kv8EsFmQVZpuh2qAr+QLTRC6HWfH/ciOri70isQKVhxHsQbHFLDF/opQlkIUVG8i
imBynUAKnIrXlJtcBHF4eJWo1H/X4PBlqX0IVT0OgTqhksmPPg3fZNr/+XddnWbv
Sw+vIQIR4EPLieX/UP4kIoSPFMqj98MSvWPa5rtuo7sQ0oUCFbHHMNxnNwbVS3hf
n5zp+L65zFxUwv0w3FIqXgdOSpIjOXQNfAFHUgUY6pzWzVNFlOcYiiYIQP4W3mmM
8qFJbv4IThrP1OJinDU1AjIYJ7hH1Kyi/84KYl43NAG2TyjTQvSNZzY5NeewcAi9
OPcThL4x1rvUeB0mEmhfnXApgRS/35F4GGGlix30BpJy2P0r0XagdbLWZbDe0l8r
osZAtd1Urb/JXF32gZuMMt5bRF1sEbqIVjzJ7i+xkDBR0x/VflysO2byKEazh3p1
N9xBcIu6Aq+/pNRT94EFWpv4j9g2I7oeH4FWT4BD+h2NyrIxiQ91g3gsuSvoOcTJ
cTiIxHkxpXGpOvLbFLd7q7pk8uWav0FFZ92aXdPSy2ABGECXX8GPELoo4tvkUDf1
fJKSBrwTd/ehhgjPuUlgrKx9u3yEC2Txx3GohsU5VZ2Jqr7PGp8kfeQijTPXt4dA
SA4VxzY/pTx91o2thTWYvgOPD08iaoHECjvTW9Xi4T1ErWzHEXi9/FvvpyENFxdu
tVMjKC/Nu+aTCwDx2Q2CTiaj2qLYJLE51U4ZWHWP28Ol+Bas/tK2V2iDvJJ9rnCY
gm8E8jZh1vH1Xso2rHF7ScgFZXY6OtCcgjrC1ion2CjahcReXReK1/PSp2BDCHPY
1RlHBGR1EjUpKwpZo+PFLpzhPqcIRpoJvFvGshpQAE6Vku47QuN59f6YDplRoIob
Dmk8NHABnff4nWuIh7pUMBFvumiDCgpzZXTKw+rAFDxpvljfM/RmNsAu6vkmzgbh
j5yUj8PburgG+gYXLyH+oTuOMEZ/s72otp4pms7K2HmyzHTwSsogS+whaK9Nio5V
sn8UhZCc4M38zmbFkB4eHyarTx01pSBKCD5zIFMqPwwzZ4+9T6Il9/alj32rSdaP
0WT8ln44EEooY4gBpyiGgyamGPUxP8H7D7JjikJR9LxCZvToPX/s6Hy+xp8SHkJQ
qmA5WtzRlNQt9mZHu6lHWfHzoU7r8mlWWxx1LjQrTQ00Hjysn+4mGIcLQ5f9DaGV
E91dpC8+c572RvhVGXyC1/TYg4hZZS32A9VBWD9uo4cz+gG4CPOfHvnlwT5bDMs3
OYcRiqrSkNjibfwTSGsM5QEnchFrh18B+hTZg+04yiIDubaerVZeKoPco2mKmoAF
Hgyd/w8+PnUPN6qTeVoO01jfPHloDEx80NT7cJBHQ0lRSyyb8ToXuYTe/omm1V0j
4YTvDaEjquuFFfblfalzt/6kVQngcQ5wOvuF3IgBNaL4/UTh9SlY7R1Q6M5gC6aw
2fwbu+3S788b5O+HDzvjQAYSRsXwp09Hl7l8vTcwO5kfp8r7LXUc+ZkIP69pgXiy
EW9zZjBLlRHPD+EhWWN93P5H7BkK1P0TIEsijq+mldDE3IErX2K+I2VAMk0prg8V
n0jJJSF0udAoNpEv7GDa1rkv5yQWT9HzxghhAUHsLr2ZPwuTU54HrU5d4DngBIEW
kH/6Blqmn9rp/ri9ovf1na/+ksSYKoqsgN6YWHI6zP6/N/N8IdyvP8iF4TgImWuY
m69YY1Ag2xAdwneHKWdfuUH8Ycr/x/pAWSBdvUr+gu8igsb7lxJi8NcLJ3phaeY0
VIxXsH+RD1FSUI1sgXfqlxQAoN5fsN22PW0cVe0OmQq6aqGpFmsIyKP3jCgjYqpJ
Jxo2kypuS7+agesgVA3Ep5PoWLJWLcrx3M+5PBaNzHjYiIAG+fqg/5g9U/0g8Qmv
9x1MpAXE+KFNMkfgr2x42xYGH30fzX4lNihSf5DxDBi5DXLPExsurHPkbtv1qO9j
zL8qyi2mYh+27TeOtou7FKboz5TRLZUDAfPGrGtGw/eYfQBj+tZ84AfXlNJfLbZ8
nm+lSCWuyRT3TdPzTVEFwLVWICAj0jSb4wE1ihlnca0lBsmHsHwq7VIOjkgyBs/h
4lLTJ4UjKqxzSp/PFMLZC3/jiKaxCLEZoYjZitLbZ/jw+MxbbI9X7rztZtSEH0Sr
vyuY0ihw9TLcjUyPG1qlqrmqemrwf0jI7OX9w3JcKHjP4DNLGeTlMQHNr1HLDthr
tVFurEj2u8vsX95H/047OrOiyXnyZECGO3D+MsmepBfeU26uRq7fmkmNUGuOhR0P
q7OdvlCIi9M/5yDjTiNLx5zlW/5UXapxKnq3YIaC90qHOj6Xrusl5QHdjA+8Fnp7
fBPwEvlOP1qFWBU0zF7fdS9doUtaBMHVaXpYPsmuQDAAiVxcB4OnfW5fi/jPkmDF
n1KJFYaJHJR+JmPY+OLlXbAPpU/6buLhtKjvJS3zKngNEflknIYadgURYU8TXnFr
3ix2fNBNUbWa088KOFYIt1yAkZRKEs1lVYnfPBdCRfxa2XcxoDONW39zC71Epl8m
Z2F23P1bHy7z6wIRcncOsbjqzky+CHRdfKFzieJG3H3bW4WgvcjU392sf3u1JnZo
ZmSCVb82YVcXrffdWTfKGzHUUhHyOCElKFfBZwRF0xfy6zgbKjcRWD7c0kMpE/Am
ULKJ0fY3WAubqCoPQCu2NqFJH2ZC1PXJz7OAgW/5ZULAzvXwuuO4Q3uRlHvrq0Qf
BlTGlp2Wb0zp6qxBXtTn6XKU+ldrDq5US2a3ttEgGZApOoUY+eymklX3mlLNdR53
M0hLyz4qtTzfDMnHJ/y7cd773nFfWnkMsOV3aTiRkAoJTi3g9KFTqYgX+rfOZoiS
gvZ44kbMXFOrBJn7N7hp5rdEMnDXf9C8E0mA/K8gcmzZLykboHK1A881PxkQGjQj
navXBwupawMp2CdQfc1ccZ97AOo//ICkW3OLkHkwRvXuwZ4RJkgfz+82XZnX3omi
mEkYe8KU8LNb0/DMxPyYdxLD5e3dIbjLEGTRGPUFq3jv4+WujMO+55pC0EnpOCH+
6r7FKgH/JRzxovhBDF933D+4qLffASXPnkEa5Jjw8p+zqVlndl7TlsUXX7U5aOuX
Me9bjTa2TIhmwFHsiUS5oSIeWz4eAqe74yKGQsrKLa5Lb7QCvpI+1BRt0px8EeqN
gNPWVJ47CIbEuA52darWZjH4moN/Q1GOoD/1dMbmDcbHkjg8RP0lcBTdd4QukSy1
DTwN+nqYzXFZO0Xte6/w/z01gHtGh1tdNlXLBY2sVw4MIjVFx4uP9xiyRtS3JyMR
J4zd1C8eTDdxHQBdKOVIzcB4AInwjEmyiGd40v/wfQXvrSWe0tCAALXZ6unSGyLJ
DlxJCH9eN9LK8TusTWgQd74mkvnKiCMWuVMB94rP7LQhtHux6HzywdU4XGtcUpSQ
Vsr5m8r518J2561LvLPfISKvePzwhnp5Axhu7UrPIScWNuou5lcaZwhGZ26+Qy5J
CdnEU4nmOyQqp23W1m2JileDnLFKMUOOmDyhijbu8vp17HFfegrbh/8vPkKHvYBk
iW/rs81AIG0spvHxUsQVrUsmf6jaQ8u/AgKrdrHqsW7YMkPmBJpU64oy4irvPdg0
kt3ASL429FrAcbztTgbqlmmVKKvf2jTgspXHi42FVB1x8hdFaj8vZWp3MCGKmMzI
YuomcFt5mgQb5PThYI5jQ05tqxLFHJmQo8iGIMh2PEyU6nJqUlNuxb3Ra/GnQ6Bu
2VDHyo7rEstrlXRxwc5BfEKR7lUQS4FcSZ3HXt2M4Z4VkLKBpzLZI4poUAkN2rnS
xXL4RuJ9WXD5pUXAMIBYwFwZsn7dUSI9Mxw2jecw7kKh3yBQ+OF87593GKnPEESm
8hqvNJMBuAXNp8WNaUPQW3kDbzlRDKqXkFKmvHCENkxzpdhx/N/eW6kodJ7DZGpi
NatyHD0rL848adWY2FA6RuHLo/cOuOfgh2mVfTKsEamkIdD35+GdkJy0wRF+iJsa
eOa2zp59IM4KoacucekES7QfLOG0t3SBEiu7mzHY8jxIXRDntmyFR+e2qNPNKRku
B1WeqmntQZ98R4agMGsSLMSmc5sFw9f2iMqcpAKcXs8vm49N3+3r4H7WTvq0Ftxp
X4pbUDppuE7V5je9X7TVfTZbzr2ieFqS/oKod4ZLQIT1GO2SU1kfsN0ppwgwQ17o
BKWTICWiHX8/yjkQeyWoKseIGK6yjhLCJHkPp0BvaNoNMbdkn1ABH5KFptzrWXZS
UeP0J0fgnMXPy8wVj0bpWGbSf2PXN94piI5uqQegGJqNUSrU+OR5tnCykbpg/JI3
oB8c9XKnUzng0VBic3VqEkwJTNQTGKMDJ5pBFKSmrZi+i/0GymLOcAUhHwSdf6Cx
epyiOE7tnHQeI37FGmihM2IegcxdxeDPW0DdMRgLdbK9nypXdSKAmyrorMiuJqot
JR6BksBdcr6gapFLOsit0glHkmbybnIwN8OTORQe3Cvllkon+7ZxtYtYPzJWmI3A
IyVNOQLbvwv52+ohj4OPD+4r6IsdHqsIusLDsUlWevJ4r5kvoF/Wn3KcLUbsK46/
MYG5l5A8y9sgeu6052UOkeZdAS+CqJ4Fd7QR5WNpRvAzv1AhKAfF2AWzX2C5wHy9
TLAglN5mB2xYrWI2LsqlQCMbdnRUsvKrTCAkNAgGr8Kn6mAOW9kOegNlLXskHaNx
ExcJu90kXu6CUWN32/Q+LPpkXYuSzn4QlfwnEs+9CwNm/37nsibDiURJAz3KK/L5
jbBL4msMPogUknMfEF1tgBz7aQdxA4n5uXkTCaXH8IEKN0Lesu8rOvhf7iblEQL2
MDcZzDKw1K8wYnK0ccRQCfDhCu8f2CQeqjJr1Xp5J52NDiAkImccf4moJ0WuaUcX
bn1MMofis1sm5AN6/Hb6FSPLjsQWKl3Va6POuI23ocfoiZTV3Fuzp1x6CG5Zyt2i
W/de16QhqlCtpPfPfknwsp16Mecd1ik2UHolQa3Vz0kYvYGl6WgxtFabcG0xyVo3
UeT75O8/mG9PyABsKp2FzKE1qRg0mrE7Fm/zeBX9aaPVmCEHxWDCHFh5DKwbhPRj
m/gH2J6rKKLB+PG7ZEBJxNWbXi5nBRpvRkDaA7H7xkh7uHOlALdsCx6d9wOQXEjL
sAANZk2n/Iimtgw4PtYrYnTEU+g90QcY+5YEeGN/Rj0QLyC5z/3do5/MWO/VzBLQ
zDUkgtYJCS0qoKmGngABANUfowxTvLT1poc213BxjQvamMeaDCxyTRK4KyjKQrrQ
CkqYht/2veR2nqXd8cngu9bN38JA7P91Rs72/2NQ+iubDaWL0ZHWV3wBlZ29COvy
mBoAsDoyDtMJhvwTEIfo3YD2ITF834toGXhABsBoB+AYheR0QyOck1XpKno5hrp1
3NXpqS0IRU5RRpG7HVTAbcjYIbniJlG/ff0RS8T9LIXgLWFOGIWNtlbufQNDL4fo
RnPHYmUpP7K0KNGsJ9pfBayV93uTYR/1b2Q7ZBWtl21RkCL4dlCpmfKsGJXOXZAv
TqrJDDLNZtFtlljzTCXL5UKzOaqxEMz8sCzOY6TmU/BQqw5eWo7HI+XqMWqbUMlO
HcNDBmF+3q93053PiEUOppRfXt6Dv50Z+1IHqIdEhLyzhZRKtaDx//ypBo3kD8iP
uBjO4iAmD3J6LAamkdhZzslrAuXdnDNtMcVBgr0tQqjdDilvQZ+4az2JaZ+XGz2A
rcZfUvtnqzZs7NHVquCMzLoB2MZX8HZOz2qG5QEXojdSMi7f1LZxyGJ8t1Tj0eyK
zj1rQP7n1i6p8KgUjQJUbLjlqjCnpRc+zxIfMO3acMGOaseupE/h8Pg8yrL3Jt0I
WximzJ7JuYRTfOmW077ez+CmJiEILUcSEW1GUvVJ1Ef+F8/i9OYiRo5uuUF2DKEK
XSxI6cV0SfKaqnMpANkpCHerE52D+nvaKOeUwmYBEqftskyZjSdKxbDTuPLaJKXG
kvNoeXWh8OfGY+ny7TtTv9EFCVnEI6OBAQ3KA84WF4fd2MvtFdLr2A5hRr8r6dyP
s8KzRQM5ic64WZNDH3WQ/sGDjAX5FpkkJ/I9BNQ7KzVZyOYr/IUPuJtwTXyOkhDj
dkr6DWSz+4P5mPK/COzrOfBXn62Wbw3cm5+/a7d5kQZutET2CtnmnVW7MBl4mpgz
cfJIev7lsO02eBAyRDksqt3JxaxdrfDEjuTPr1lRYCWFfD1AQvWWy07QwPffdju5
oxpGpIpx2MwgBXnp4TWAqtmWaPSftWa+Sb5Js+a/d1fpmcm2PxOTVa125Bx8EXcZ
1xWoYar0gOmMqaB2KhV/iClLTEI8fudQxx5MxE7Fv2Zn1bk+rWq2tcgVpIdL2Xjf
ZOH2z6qvu18Za+LU/le8pw86DJOGSpEafUxeAWpqS+euCOyjqjD135JSOqNK2hfx
9Uk2iCvYEhl04LGVyzJ9tk8N75fSwP47L3OHib2fBBNmgIe21DRC1lor1ZTezyVt
HT2dMlAzDMiXKrvReBVy0UdHUPhmgQqc9jTREpX3oNTxoOC1k+djY8/HsmBxsRao
o29/y3xGP57ZKhZizghfDBg71I3fpaMpemW9GR8HWJHfIOhZt6+GmJ7S7knfEcAC
M2VArPR+6xO9x9j4wQXfw2E+aocvVB+aJV5CkhM0ktgXXdsVDjd4Xo1qWDy+BTkS
Zt9gLVmqz/b5lpv+j2p3opeHQGrgPrwV0VdPUOIYU2h7TQVvA5M4w2p9Nv55WOX0
iAdIWgtgSYBXFoEkawD8TpmBu67cnMCOdj3d8+eFril6oAwtAqk9YGZTs22GWVkn
rCsv+Qd77GYoHq3IacMUay3WmFy1SwvUNtIJshC6EdbLYYn9umA7/XOuzPWbYbMw
Csewdb96cimxQehu+xr9m2uQFwSfBgDZzhYAA+174E5B0/GrUwD1SWw2LTOeG/4/
MsYBNl1i1Elq4WVR/272Cr2B+dfvtYrzefoTqJbb7xjkW5Ars0dyc7g7+46Ri1z7
FGl91l4Ffkr3X7WNJOoK2vJeIHiE6oSasb290He9QKROf2raTZU2xYSrcU8CbdYL
cmuxZ/wAPBpW+0BOePGXkkmR1QEWh3p1J+EdchLwuogyEQZ65pbo2ykCVypnPIWy
n9UPtrNx1p67PHx1Gbc2T0pM1qGxI/QUkCMprhwiDY7Hpn4NtrfR1+UaJ4U/LvKJ
Yqwi3WfwNUjwbEwNqVYlezxXPomaZG58M7UQzv91KKxgX43vkQJMgggp0ik+rDY6
nAvO8yKBPsQCod11zI/fwOpD4ZQR26N3bUs5GtFcmMtSgmzT27jZKJjsJhon4lHu
bmmo/e1RnpKXN6xJZ0nkeTm7vCravoK37G10V2ARPbItyGx5YBlIwY+/2X0Trxt9
1GOmoj/JekWLJneJJa+Zkg6fqXoTbrMyuNBPoAQNP/0Xg1V1GpAkAl3IRWpkNyRH
XunuWBSp4oGuhMsxuc5RCxla5MluRnRVQJzm2kGjJNiYmyboeXMxXYH+IJKk2v7G
FrcyfXeMQor2wpRUN7Ry8ZXEvthdYMs2U5GD5TeLgVLgJkz2L8DcFHwVlH21SXpv
n0giFoZdB6MTdNlKPuGtMW3o7WqSAghnDSpyHxXlr71FaV2CE51rj7jOPvwPp7Qy
k1i1IfBaOeet8j1D0OMlPvO6UhaItA5Uqi9rKUZTzDHBeqRkh6HALbTNZ04QHxX4
ERnWR1ZKNxY+jygXGkkGhSzCCxyaH57gbRxnXOzKNl+eQQPQbcRMc23C73hXfD60
ueU7kmjOtQfn5s7JJSFaCheMZJhijLFcC3oTPhCZhkvR0Sr2UnzeafQpuatA9MaU
ZV2AF95EdSvcNmBCoE79n/XABveocOJTuHTs75WCD+DCSSf5GgaFJwvmhC05/B+f
LYH+ZjZC26+FuVgvp+wnPjcCHWSJiK/QNrUKL99ess1Zs5UCqvtCRBflaYrPxrbu
HBlA/USS09DE3mqiaCxaKc2vmS2FEKHISBjy7ZJ4KauiB8W5UDnhbgxHpfp3TNWm
72PtF6FS2d1YCc2oDKTfzmCMFAI0MpndNbeG2Yq8dyZTzv1jDCOGzxQRu+W+Z5U3
u8nQ04D/hEoOoKxYoPltejFP4hZ4RNqSmUx+XMqW4CKB4s9+l3N8fNklguQeMqja
99gNpKby2thiRntGtZPpoNa87VEjGDWr2RMmWvnddp0e1w6fSZP4Vpn9dJXyMPlB
NLYq4AxRhA7yOoG4HYdOKcMY1oISHwIambmII/eZFM8JyJjelQ3wG8B9Gx/Ow6HX
oD8sp3Mmw425onPZ1k7GL9kmYKuqy9F05tIrVeX08pQ/JvVRkOZMuVObzmtJhfPc
GyW74IPVvJroldjbEcvYKEwZG33vvyoQcPOatA5unqIn6buEHzMxOo+WTF5JIV+3
EynM1dcuDoseHbuDfg5Z7najC5wPrT3vxOD5TZx0sCPrO14SooutM3DD6blwjmiG
ymol8CxsM/+VWcxuIejbkpDSNPdQfxNDChxFDZVyBsdyOS5DJa7ARkMwitE73+DQ
c1ZUdK56ybwyPm9cZdyX8otuhhDg9RVv48yguuVKEo0XJ/Yorlmb05EDNSOmFXib
NAchQNcT6dByClnfY0W6CELYGsgLb0FxuoJNidiISsyU8yo8SWGNnfKp5KNqYR3C
cU+U7enyic3dGtscMqvv7cP45lQqAT6hW+nJRBqrjygMMldmibprijzQFI9NSfvQ
gDq8S9fOdW9+DVefgynpuxn2LIaJe2GKo9aDeNIm11dea0ksSYTvUFJbPObck6Xv
C1YtbgS5dzAaBGGpgCGgCZ+GOlYHYb5cSKCFnh9649Kd0qNO3I9+i2ZwAtYn5ndM
lF7C+82jVEQeCCpOwM08aBbF3nPkhqkzr0WSnP36MlzgQo4O/d5GpcbmKIEWBnsJ
wafQBULX7Z73HTDAvh0qimm1VhfJ1iQ5PQ0cfwn8xxXWktavNAfsaiJGOJyGmyRu
NN2CSt0HyhyQiHVzldIiWahLQV3haAeT9O+J7jKDweoMar5LsZrNl9/ZJcDQMcCR
kAUn+Ctak6JfkW5e7S5pp1uCgb9ZPS+PEDrcra+fxNw=
`protect end_protected
