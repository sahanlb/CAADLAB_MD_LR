-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gV/iQkMIEtzAUNi82lGbSR22eoeiENK0zIALIf/kf0ls/q7pmed0r1knYRb70WAd
4+DPI7acCOyZNoDpEvm/ijdCwfketHPjIn1ac+1gfmF7+/Gx5s6k21Ewmj/TQT0W
+LhPXfcT6yBKVotwi6L/y9NoOJdItSNwZKkvqlFNKOw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 19708)

`protect DATA_BLOCK
oKtD7F+aNE9vbKa+10nM8wiKXmLMgFE8Uq3O+prvoYZ82+7xNq57Vj+Mqm4ePneV
cftk9cYkkjyq5LmyNIONNf4OL/dqub/3EQ4dWnYWHkomxQQ802xXco+65pNWBYlg
4nGFpocBMWeh6KWrsdMR6T9t+KWaXaWnoQYN4mg45nNwesbYV+NlNCuBRiBTrY8g
ZO2gtNfidnJ9OyVhrR6SPvsLyYbxAa6KnN94M8v93U6gTgSCZGwjWNyXQaLMRena
TmFXu+B4HTH01q//ErLSfZM+V5hj+snzvQzYsDOe8vSHKd9NuXB+Qw0SOQQIsbhW
L+bPfXsXTBavWtEzwA2Mplorx6Jp8bg4z56ZMUKq8oOdfLya7qICv+GjWfvObBjg
UikEk7EAgrY0wA4+WFEfSsyoZVu1CtQ2y3ChfeaprHCoKnjNPbcifCDw3OpnGmnO
XXT7lhKN62WymJQ5pyr9QFxbUDg8gwR8cXFcVq8DDNbe0wrNTl2XBG11/lhL8G7P
RKIsHUl14fr5EdFNUQhj96OhTlsWrY3DKnai/JR8rriJlU/eDnTIir/qrxduBa9N
xNYtJFGPI4QM0aAgqpd7WVePAwdqYyddOmJ05oH2BfDtj7svn9W2a+bRFt00k5YE
C4Iaic5KAPAUWwFO2IzuBFxW4xIFJHgquPipF6Ia/jhvRjklUb15xwNwt8YEjJFL
PVEe0BA4XCi13RSoynIxwzj4+bxnKdg3g+5Nbxm2Ax4jVjGFZWELqthRPf4OvmsS
YrqABXKi/M1KZnPHekncy7zuJD7apuk2nPc62Mx/sIqNfoXGzDfjCxAPz3+0chIF
jTNxTORl8dZV+59S2g1nG0D5DhG07fZ3R8Liy8J+nlfMVp7uILQyRshTpzqNaRv3
Ee2RkX+27ZT3YX5j4N7WlwDvzP3vDF3sIrS4N3YJYBKXkc9Q1XRmasc+M5kXQW/u
K4FQ9Gk39vsNpHDIvZcl51shy9L/48P/3v5EIvvW6P0XUCj9a2/oNoQszdtPZpcn
zG+cB1HTnsimBn/DIzkh2EuuzSOvbJUCqQlkyDPEw4c5TBXQrvBkhtSqTSrTlHv0
CiDFRP2PuaMyy3Ekughww6wzmP54VPD6tHR3AeOzfjevH2KfVce4Ymz5WFU5Ccjq
Z+6UyBHLd5nCwZ4IP9fuzLHjhU2jyDwRl3VssHIHx+DhuW9uRVILwHfR5n7TUokd
keCt5zvRD72wUajsrQ+7DScMmM1nYXJ7mxU70aaO9L3ZOHTPupB7PdSQjfFjzXqP
Iho5O28u5DzONVK/C/WfURcGObeMQpkC5lvbrHWCMTsmQ5qVSAjrz2j8HbTZRDlv
xCfhYt7+Y4T01IIUlH5qKpsj/jC8YrOCCu6Vf/WpIHvtyiDFtNxeGwCUSmm4Z8Pa
cSi9x2lQXUhbFLR4A8LcsQ8CA8jhpScsGTZA71ExoeDTrwTETFvjD3PS4hcaRGqI
YZk2jU6TQD6ZZHRjxRUVtNth7rLEZnpArLHAFmUn+BqJNOINMmw23MPhIxzzt7va
ZSuKTSkTmZb4p5Ip58YY1Y7r7J7Pc1CyG0TKz8hsmNHXImflD8CQAm2/PVPeygA7
7+5i/9YDvhnjUySI18E/bzKBB89U9Kr4nl7liImAKXGl5dMP0+Zy1up3rHr9cS4U
Fh7ABMWajd/JlbP1uE4zhtFs2OSiPsUHhGrU6VRpAfze9k+5dYCZ/SZONzIcO63E
3aMO3e1VPmXGl/5lvdBYT8xakvtKOSWimwN0t0h03MTMtTBMgljHi7cpXHk4RUgO
iKxfMv56CrT984kw/565dge6zk9rkoywsY0QvbcxRVWSL5st5b4anDxocjxPc92q
d3V/XtMtbJ/KKJQCewCsn9LW3R8gDHKVQpLeSRZspid6Tg4mv3/b3977Z29FwUqB
kFb+jhDstUq19GtlbCS0Y11pnx95DggOfhqFtZm9FvPj8G+AyDNQEkh9FWwYNuaX
SAYonFKdQdQVz3eh8OIXWaQf/6zDEMsgLivFmGic/ZZpJUK09upD4OCSLB2tMAQc
MDNjD5AVHy/SXKcjA73d4+45faajP2t+xR/eq0o1nR1haSKJtBSBnJrphYFgly3m
Cc549iunNw16S9HH7rrtWoU9nhGSWCYeBEJiZRypx2EB9I4Xb5zdJC4HZHrSK9Zn
NuxzkkXHKRxCPldpN8wcH1+BIRz6ApG3VMcPdzyc4yTm7qacLyfVFw2eeNEVjj2+
05W/kCXhxIKXA1nyuSjxTonYfIkuQRqCtOCOL3DXeV3mc3aRx+XTeMIReptmd3jS
uT2952T9rDR4tUAmLIBcNQwPn3p8AK4WZ7X8WLX50dcAluq6CGwi60H6gMGupfHK
K4HS3LpUoCedl5DingJnwwZU7Q16wvv/bqvdnWSTDCog+XptpgWN7RaWhvUs8XfJ
w24sysZHrM7ijtc65et1UXDl+VERmXueDaHhM/+mcZvCy/YYiHG+LWUON4dqglSk
oqhjM06KjdlLMNlSFY6+QCnUt5tjABg5ymeWPBHwgL5WLX5aQQx2TSrHO9CVHF42
3EIKIC7OLgWfeDG2HlyUgbu+X/fHHI+XLIPL5qyx6Tv7aLn1Zpb1TA4bkPJ/Gdjc
diI3My6IZLFgJqnpEIpBOmRMOW9i00514gxBDvdC2MOV9cPH+DH+d0ktgClJkCEv
yvwS2yRwAWcg/71vRWUMilSSC6ktnjiUGGy0Ln6dQHTEv9Sq6Y5wt15NPgzNtQe0
eyhxhfF/noXVJc/oVt/u5NuuuYpn0rhm9Bl3viNtP7ZO6DqDw9/nByVkBO83Nzmx
Nf6cuQWEZSipDmJ7A1bUh/y5WoLcY0n4sOgJlLWn29XrFutz7qrBu08VayIcTiB0
YuCqG+jg+chi3d6UsMqV8XZR6qnRMDgm8ZX4eOSjO2D3e4iW+J1QKgZHHsVxZIF8
PCdEp4HXlc24WLIoNF40pG/AE7bNzB9+E/ZqsKh4FWxDrKsUy++ltBAo9+ThKtBI
sA1TiCbIlegfBIA0Zswe7XavCTGr3RZpJtNnmDaxF4wF1Fa7U6v8T+/Kz2kGUyHi
dPJUG3W1H6Qpqo6Dug8GZmfVP4jDpJCTqhWJX3saaJWZCmUlpKPY3SJXxBuupW2E
VtdA4EEfMZbPk7pvwc+Uy8kozZzw75+l1b+N/2OWPkb6qLG+bpTlBkAfMXTgHlv6
7NESVueMyIdgpCbzE5FR0v/jr0NV6tUTJ2uZchbhSV993ig+o/olGHAvdudvdN5j
icudUDxcrCjBf9YU0ttmgX0b5knnQbEBsXYenlVWqwqLghtLT9wPOhkdAioASGcU
4ulOK1KeMTQKasuYKKd3sWxpUgeAdBiKlqZ7xhd0rYwcDIvkqxbcTVGTJC6M/hDK
4RCYpUW4M6dMWws9DiQyQSB3GKQGUNeazSC7QBjGTQtmA2b0u8VVrFmtOoJeJYqf
lnseRtKjiZKZTfoJUdvH46wgenjpW/O5Ndby2/pJNfhA7w+47aI48IRWZG5aOX9w
vKU3umKIheqec5n4RCHWmR2LHS69cHQByFRbrEM6kiJmo88JyGIqdU6qqmXwOu2b
97/hOUE/23rGbzNcb4uwAEGz5s0WnAKhlHsMmN1sqQJgHJ3IM7AJZVRptkv7gd/k
+xuCfESt0D5k2Yx8SspXgsYzMMV0KJ+LGWrkFREai13WNMCEKHdBwz1mWWZE+SH+
LYrWfoJAsAj45KtgrkjsU6L/Pzoy6FyaT/Qb372O6lXeUkkR66BspcQKFuNPP3nN
TIKBvjfl+X3h+SjA2re12/T81ad+5fxbis9gcEL8wGrJOZsvWfHG8xB2w9OQ3bmA
cDxdtO3IHnmMYi62pCF2yz9WTJ7di8E8AyUIkfaIbqv19oIJ7VZa5SIaazi2Llje
4r/dTgMYI0CWZxxrpzzr4N9vewSl1XktJgbLFqFpM7JNhzj4+fUXLKCYae93+kkM
MhorwBf9JAylX0iHIUn2/uuKdnjMTJfntX7IOQ9JCa7+w5Im+4/WH3kwznkqEdW7
thX7xcZ11Z4b0HBLzf/UH4zuAZKHCh+fmwPdeegSuZxfT5t9WL+WJGB2CdcuI7yn
ewBlGHI2oPZ/Ypa/YGyPaKgAY3u92p18/uLpRJwvvpxr3/fnzor/9G+ffMrQV/hD
GPNNmIGwkO4d2H9xjh3uE84i556RkGPxbHmbYxWBIijdIEi+4rpnmib1BLkrrk26
BUxNjNp0ZbOJmz5UsGUEjApSXo7wvB1RiQiZ9yuI01MuXLYVEYy8y3lG/z0Nz022
N11T8zEF5nHPXss1QF1aPDWqmGPeclBTWHivefTE2zeOIQkfwQtB5qlDKbvGwybM
By0s08fsd/eN7YA51NJ1nxYFaYClG0MgC8KymxwifBcJTIuYv0ewTzItiymRB45R
Xd86e7HUpSn4dmPsBMcF6qAEDgGpvKE2pEKsr8ls/kEgEMTN1yISoSTCUuOu6Vno
gi5j25xTEXp8qfLZQUZ2H6SkODkY2QTodcnqaEcL4VchFcEaG9gCzbqPowiW57nI
SiG6BCAbuRk0j9YG4AY8nGfNsAuuq1r36nbDUggLMTMMJuEOisKDQI0C4hT7QG5s
Amf0LDtDUPXbRtyM7URpGbsOaeh/4NB5UIW4NE3Bw3PA2kWMkUdWoG9Xcgx1Bz/A
Nxlcppo8JKnAu+7OgGMnjSjrzLyuwZ1el/dAhPPov0cUJEtc14OT3vsjNVoRTVVq
+fwblbGGjL/PQDb0aqUJ7tdLKFyHm8P0B1ZMWOf1KhPeX4s8fCeDTbjwN7fXEWVQ
s8iJXNWAEhNebisYsE3AKV7OtXHvJqwQeKMCBlJbRW1Uh72262BbS72Z4Z4txaKr
iIX8/omAtjmYhTVNx8UfKVyqwahOWhg6Iw83m6A+goZxsf3Q2q5PFFYEAWMuKBj1
N0qnvhhAAhlppPKcWoL0gxNQvxEdZCQe1VX9DUWvp7TJP7R9Ag3V99MA5g2QZlIO
z1lDW1rhJdi047akpFe6kK91tNJQuMus5yR2xID3KZ1dKhwbQjDTlGdo3iB+0Ow7
vgeB1U0dJ6Xfds0BWuofJNvVNyTDiu6g9BrerODgwrdaUG0HxmmulnBrq6K7oYpH
9Kwq0ztGUn1HZqz6dftokjkXajjAUSiXIMt8x/rdqGSSBkhbhSNN3gWwub/6wA3s
8+RZP7ksKkw25/Nh+wp9FOmTOXJLsi7ah1QqoQtOBE9UuR0gkksCo8CzW+9DJlJt
DZlZBffe5u71fMpt+pFrEY7RnTiFd7/af7BDzbQJ4buUVqobuc9gAZ1Xt1WVkJnm
u8FLvn2ZpaEyfzehMyvCsLKptwkGjB89iMjEfMruTXrXbqysLjuImbCwsbRnBumK
s6uvQBTVe0ppHXQ2yEhNTIDJTPsPTiZXdyPKcvHIWmqyPIrJJQXfHYxkYPpqUKG0
0agacUZd76Y6gPLCIcEXYlmlaLP2E8frflrzofE8uwqjWYT8o1R9fc3RlK5D4xKC
jtM3UxzOWRw9YGCnOUO0tDYRQ9IO6dkBjVx0b4Eg4zrNNqPKQFeIMDjjssMoSK3J
zAzSyXNultsQdn7d0Cbnqb8SFCpw+laPvsg1nWf0B6lUm26CXfSLmKLQr2xY9M+b
jj8aLSzN2So/iFf34USilpMYQ2/YmMRSVT2ItC/5MAVNsXjKePDjcY8n1TqJz7ef
aeyPPzjWhTEnOqO2uj38G64pj9tGmPDLVi2HB79Y/AoU9Z4qvYkpW0pOVRrd3YDi
5aLTp778+xl8CqFN6I0coTxKIV9OZwxCXrf++Lo9fD3B2MpEKcnG3/GGoT593avT
7PkK+J6NI546fMMCxglT8DEI2OZH4RU2SqxfieQDJYuVNDq2LhNTieY8/1VWkUR9
PQ2SQDpo44BT1Xu70hHNkzKIRR7hC8mAbSN1xAN79euh4h7AXuZjrjpcKIBmCqws
o+iw0Oo3x4Fu0QOwRu+xYOY/rfHqu3jz+7IAy8/uxGNsVBTAXYDFRPAfA62BI4JT
cPokN0GLB4ZbDXvUtL6Nn/e8Uij701per4g9A/Z0a/HT4VjJqeM30ccUhdPFmh7y
5RrPqnxOhgsU7JA9T+pJ0PVsbI4OcgLOZGm2M4VHS63/OakXFUl6VI7vOhvdGM4T
Xb3L2U5k7spxXVwpDA9VNgAUJ1U9JUCdNYS3olj+7PpR7JVeHmI4raEuJ58En1Cw
4udiyOfoMCzQ+MkjSzF6h4OamcD6yz1wB7VNv9dyn6K1QEEuRu2BH7w1fpPLSvrA
1xhVOMANDwIx2YRmewiuXl+9py9r3FKcfdw3zwUDgvRYcyHyZb/3q++B2xdMOn80
/6EFuyaUpFVMznOWlnWxkjw9vfBx4pbJaO0BP00+wSYYHPkOcmvzJRaenagyRIkx
HL5xIaSGroeQ6u3FeIA3+x/N2GFZNztO/8cZ3CyuW5ZbLkLRRUL7e47oU4qqmG24
409mPjTNxpbt4p5OD+5iT6i5zvfAfMY68l8GvDje9/yKYZfK+SEagjBqa57zHmk7
/Bu8Ocoqdi0W/K/do/kfUZ0AbniHJTdVLE3FlgfWDfuheqlFW2SYSl5p7lqVnmU7
4R60CfL49TbFhC8vfU/LKIknWOvYtWrj6qSEORaxFs588tikhk1SPFgYGEtHIoDi
3J0vzAuOFUltkvcBN74p62ATcUlOPMApgPz5BE1d/W/sceGa1nz/XYJg/Db7/lqa
6CkMqP7CMVAQ3hr4ciUL4LjPvklfc7lIjdjekK/UFh4f88IgKzRzb6v3Wsc29xKT
0RnxgeTVkcAWi7Mf4c5ASC2J34K9BShko0Ho7QQtxb2K+bp9cTjwIAEybMYTOmfr
OJPkKq6NfsQII3DzWo3d/+oIUUO5F2cobJgUbdYbXeEtOATr/itmeiu7RhAzyG/t
xcSbP+7ta/+d9jvxfcqU0VzGDEIajo80EN6Y1VJEQpf1Bfia2S0EDSPhLD+bon6d
A8+1DLYg6nMANoVU68BZomjIYaR52bYdQWyOqBuyakqmcqdDIO/jvstK0z0Ax3bb
9PuFzKBIkWrCrJpb32VthGMWsG4wEoI4B/2DeBCc98eNwua/+d2HTlsPgeRcLAux
HZkE5jHwBVW/DHYyT8eMyhH4Wup4qsc8ze9RYMY1cSbuLg8egFE3aayxJkCcagRa
MVLOJUBPSKZGbwlf2107krB0kWLBoCzimWstNaFRfmxGK+JKWyMB8w1XXtwsc7kN
mczt7Q67Sx2AUvysNTfBu22aaPzwwnDoAAVLXlX8+OBinauo4q/GfP2S86I2hD69
x1IPbvHA9J6COreOE812GxK0/rsRR8c0PFLLmDRws600usFYlIYW3++9Wi8XoiLX
YT7+bFEbHus4WKsqKHlQMZ64jfRTW4oGvDFQi3qyS9amqG/3gkxCduphPUHvF3sy
P5BT66Cc4xAQ0iY6rJ3ZzkAu/SjEwKeb2Hv1lt56aZ/N5N/HQ9VZB/qgAqt8KoBe
m8yXDNZGPxbQDA5Ma+nfwejgs5HqsCwVqNqh3CK5tsZ34wYZiRUvTAJocLxDoZJ1
EeuNctPzMF1yQWNMlQ+3z2WzOh10si6ghPczMkfrcUeHtTCUF1uSDAj/BlXUFabK
ynS/2vUg5Brg27dlPFb0ej2ZtWxDnjBIsLwvq5WzTQclZ7Z6R0VZIVoPkeVpDgLP
YlP0ZsvsN7xmzn1ZuyHwQXHLuFpILjFbzbj722giz5EeOJeQ7e9iMRgo6rynT4yq
wwm9w1gp1GJEZXGWLVmLEDYjbViyAySarNP9PBH7sGTbugNhewLbEU/asIkrHI1n
p3wdkKbgbPWFpKEtwocUeXZfNwXYQIHEb5RcYDZDmJ6DBuZLrFMKyXuXGYBL5Jqo
Mqq2NyKPJEE+HBKMBxNT887dabeEzRnhRX+3tdebxFwijK1S/PYz5tSKuV5qH/CP
oymePknGs1ACFXqEIKjyDDtj7BmJ2cyIEhR0Qn5CNbdjaF7Q29XCaSe97RJhdn+t
bG0WalB8xun044/W/kw+LpChYzMRZzMy3P/vb8Z5/hlNRJlGV2L+1r/iGEOrLiRp
9LzdXOHP+8RXAaGs2L3rcuZWkni0lZFoBNQbFPRn4dTh9bK0oxvErRySjRB9PzNA
vOYzHFhyOqpWjsS6Y0nsriwQLVb37zqlNgrX6J9dFzWvplx6tok0VFt5J3FhINW8
C/+Sc4RUtDLnmzT2Ku0rYm2f/FXOjMPJI2nOZmvls2Q0JTic6JgnaeUDdzjaDqTl
Cu+fdpSyhPBjDx7xSs2gMRvGFVQWtxYzqUU4ZIQx/It7JxBZA1e8Kn9n5e/Yuc1m
QpjTalhGrMFElLOhXYzVZWtswq6JdgQaLnj2pN/FDCOojaM0l0hdvBjG5laFUaRj
HFDIIxC0YmG7oniWAAluqfGy5J1zYxTd2KbQcpDrZIOPx5rFG3dQskyffPAisb1y
5o1CEg09ZLg73+H8GEqHNa1p75Rap9ZNJrrVuG5OyaAYrwXyYP1sBDQF5Gnw97X0
kQ69cJ/J+XYptTuADyE5ASojI9lsH27GkJR3SJRYn/BrQBRDLDRFftws0l9zfFQs
zvZsVFlpv1U84t9wE/vvbdipbygq6u1dIZLY/cKAQPP9GaRN5bZYqAr07nJwJxW3
yhZvCwc3SkMO2qgCtYZQRqlcUAX0RBzi63ouEAadUwQNVt1hrP7bLQG98AtIIcaA
yTq+RmuKyyWz0FuWx/ctIIp5/S+R/Uced+MXatHZF0C0w30YJN/QNltNPcKIYWre
jBD35eDYL6/3duLsqOgdtlLjBb5RffEsE9QE/hNMrJARpFhJkhzUjFWyun4PXm8k
auBq5o3nLYt2LTFQboZ5hQP104Sij+r/MPogk+wdNeKHIeHvXAZYQrVEiODJgeFF
iBC6SDB60xE4wFCXZLhIYgDpnvKTEeLxbZqrgfTDfXhnlxB/uWDlZ5NwS3uZo5gQ
K66nLftxBNmkH5YCG3QlMYK6SjLyAHe7UTl9CavcCCbDyob/ubx6IrRjJu/k1+F/
MKJRn4idBRT6qn0qBM2Ir+7afC09SdhAXiGT2KZaSK8IRqXllbkfMmuU43N03G+r
YYyCaignaEhKd5bOoguVI1vIHIrfIG/cAXHXdPWn2Aa0DENuOvTWLVYKuz6ZCjHy
NKd/7W8pQZVOHle2uOxCe1tNlOWEX3MGV8PbSo8RDIZpv6bmIa41tawanglR984L
WYY+7BVG7KRwia5C2NSB5u+ckNsd+0KoYJijV7nGxJKZCdNKQnZS75d8Mf5r8odo
3WId2cT0py4hjNB3RUZvyCYtvxvLltrzaAodlOG4KIz5R2GngaY509hNx74RKw3o
58pG5J8SMaCN+7FD367ybX/mN4tck3Rqtz7qKXheNLRjW+8HWGMbBy5jNBm6zFQO
8sgFazyn8bPsOX2nHqJIYyuvVQgc2ukks/s/HQPTdbewpfqRBj1g/KnCgwiP88QA
x3CpL/1gcuNMoD5aI2cchYU1Ps9mycZgs8xLWT0CqC9Rw+4fa5uWpi3k2m1oBHpK
eT5k2ctBuWU4jiuCYT2ptdKI9z44QxL4T7m+2OVxbBR2vbT4WWo4I46d4UzbJU2k
XpWHyZ3ABsA/SrLyPpibANBskChzJibr2QdL9wE/1JO9XxKm3GyIPu+lR1jE+tvC
bAwf0dbdHtDcRHL2xUoJ+0mscarS9GTn/KaTgSleqcUtbU2sAZTSETgWKTyJlBfr
csgHjj0jDBEjoWGnOWb1tuUs5wuq6ednMCBKKE08pD7PFyMqNvW5owhwRrf1GEPd
tBy/+8ZppXvKqM9XIZZWo6laMxZIQBcVomCHJWZJd1lnAubjBlSgRX3KwHCz0h+a
BnjlIy9QJsW7clBtF3FNV9aHs8kaPztBXI7VetX9KU/49GAjWb8TQO2ALBp/zlUd
Gpww1vgEh9NJFoVZ1CoMWChdNU26LOJ2kZsBqbcCEKaqoYAdgdJLRttjSAVQiZgC
hU5KwW+psunQQ7ZS/NtibrWsTpS3hdZSnYChKQTrP4Z1VnYvaQCT6XCBIe5z8xcy
WrZHx5e7jyNkyHOsh5i5SULEktuAVT22OrNmZA77t7b9ur3kiAcqym7USqeP8ol7
17aufIXeNipzWXUcYW+7DEbcvzaRs7TCPenerdnrantFwr0tQlKz04cpqdxW18YT
t9OLge+tflp/XF+QzWExPCvVbCevuRf8rWXc4fw233J/cMzZRaPku6QtL96ebUt0
/QotTkqbs+QVcPB0yYYrxOYSsTXsT38Tc8EuG+B/QAbLp11hw0tRggjn4YPwmP1c
n3Ml2Hkhr3qL23lILz5vUzcVPs/M73maqbbSLb87cPrBkabp9oxNrYs259IoY9/K
ATiFD+NsZQvK9zExoOHDehIFeeRYOgc4be4xNRKc+o0RA3VowJYL7iBitf1+h2a7
Ilp6WC6erb3efGaepHX7btwjEC7MSS9dfi6CCn+EcgEhjuwK6QcZ9kIkFlMDQU+0
fSrWgb7DqGBBMlQutTRDP25HiEK5ivkr7FRhxmOdMpGpnXgOJH0Cd+27+U0+QJ2X
Fje8vi0cmsHHhmQ5nnfdjKC0mdLpDR00mHBKsm8w/LCDE86y0WNisjgo9LMWQwxK
j9XWe+HID6VCm3Q0PdYmiDDshnCscQsc9W26nbAsvA3kFPWmuNhg9TpGsknADM13
N9qCF20kY0CjgsqmiDAS17OssuwROid4NqFAAbc5jylUhFtW7LDSeDhEh7ggiKA8
0CNFCiUwalBfArOMYeqN7pvU9C/0jHdj2h9uuUQcbVsD+LLBDtePdkIF5drmj3vm
xxWYDphtCYt2TjI4AdL6gj1lMRWm0VkQdw4T/fZWOD7PFb/3texKQeJ5tiwtVzev
9AtnUZc/DbACOftBckNZJr1rSaEEXRQaR2KsdfjDShFfUqlBRJYxvZFUoPb+gQCV
hX/WDnP8MDYZdlvAoIUr4NlkntRCxrfaA5hkvNBl0+6JHAz2jeEciq3RqgWWe5dL
DeAL9XvbOxEUTfWTmpP8SrnWZZ8hCSu8inuglQKl5MGL0lz8hRN/kfwvyIUxrqG1
4vJrMeoMOKBxxJBXVOTfEOKIcD+WOR3L6HlyekwMolRBpgNFStCubTfdPMXLISz2
tbxGBZsFAFxeQQGIUchb31h8qbZEQdB+Gnc18QHW8DVYfuZR4rki7iTxKgw4KvEJ
GYMOFg+dFVPvWLT4hzz4xZRsO5JFtMl00O7I+ZKoXaXjaoFOR4nQUhf1OSMNCN56
TQTacu9qipymtc8s9fA3cg9r4ioXxWaZ2mPCGfOH9E5F+qJmtAhvgcbTgnF+ROH0
mSKYNNCX7pZT5F506341c6OcARYIreFI6JqE1m5u96rVNhF2B5hqVy8jCI9+tLkE
InqiBkk2VlX/Y6EcprEbzwnC9yye4Nr4NfMfLsiavVRJTBB6QdRrTl6B9f6Sd0Qa
2Y+gtrGU5kvXyqK8vEXZnNK8CoWfgi9Dzc07Nn8hZSkGN0MQi3vOeu19runy6f9u
obfy75GnQZiI9DiQyUwmvNPQpmhV5ZFJMd/AFoEAVhFpS/fmvYNDxv5H0oyPWyx/
bvDNKYE4zbpS2O6mWDqzqgz3iewZcJqCbv2sWg74A7BzK9CY/JDHeX8YeBXme2aj
jK0AN3aomt3ihhVsh0g3o4pR2LeRq6XingEQ5Om2AS/fVTBc3De/3plE7mZa57fx
yMh1T/I9z7lKkftelHTGh8CnPAnF+/QXYAcu5WjyqnPvRfLEV5nLkyVnMFC7N/vY
VziWIyBt3/riDaFSuObAUEeeO9/xoObn3nsIw6QBXdpfmIsjVMg5EJ42ouEPd/uR
IJQOCJrBxlzNW/vNTJddjsyctbPa2J55Ku1qiaEvQORm/b7KJYdburcV9o/9Kg7j
i0vy4b6y9tKKwKeUZRuXgcHmx+WcjBWiDmTQqzlQsb5w4GTFTotZZX6tCQglXTAs
vwDcvUHYt0OhIepLtats3e75CtJkz2FxuL3LTvFu1Ow+OVd2lrdo7JlwfgGzGYPx
nn3X0f/slVrQed14zAp0BsamGimCE5OXhJcKlPhrxfF4wBudUCQ58rkZmZIfK6p0
nLxlPYDM9ebn2Ak1GDBGZQoJmWIOeBSXEJ8kkdQQ69UWeyRhs4pQeLwoUSlWmtzQ
hT6Jp2zWpHniLic5jPdLCuM+p8KQhRcgZ8T/C4JK2Dp8uit527dcF1NDdZS04yl9
7Aq64UWI8H/INVlAEnexQInRb+h4Ae5dVlDM379jOh1rXtuGrttiDC4o8B7/zn20
3gjEJ2wsRxe9aHz2RYSHAGozj7Ddh9m4wruliOd8aVelONi6ba9WrDYOBKtecCQd
ruK68oM6AwF83F0+qGt26ISrO/b9vXTVIg2kC1EE/GVreed97CzQxhjJeAjgvSC9
EBBKxp7kGz0yI89xoUlS6PPYQT9nS18SqbMRX/nCT/F7DMLtQXtAHmmRED2NCWsq
Jpl5oaBLLBG0WnRlxX6DZY+B9myQ5ZZNTU0psr48kWuCTh4dPphA8gk6oTmPrrEf
Gej+dEjk9ruiXnk7x/fu7O2Kup8hVlFypl2nUevU2/ILvoG6yjvj/clJX82u8z3c
J3qoKQxdSa0tP/mitMfDVJZKq3gSsYN9rx3Yaj6w5HKKQhw1ISI+828JhIpXirGQ
AfRVaAvJZkCI9G6E8u/HT8sWZ4G9FNmGavLBNodfpKbuY3aKPWemhWofjNxn/FG0
xF85ezUw9M2orwDYvRo3Hcxdxlz+3TLTWrlaC+1UcIgnANOIa5MBDhIV5wq2O0G2
UmHB0seM+fnhZW/5ToufA8TTzFHrKnXs2KvYWA4+9/YMs8q5GlFQH2Lccx2VtDff
vpNGJszlo8RvUYkyQCaCIb7jB2TiD0HPDSJYgFPMLIm+fANi/mdtJRXQxWd44H82
8Oj4IA+JGVMeh3C7SXZA0EzNYAK8bvu2+eSr+u46mLoHEL2m/HMCXuwflzGnsKI+
xUZa9SLd+Ff5euSK61ttRdmtjPWjr9szBcd7/HTsqO9XfAN3Sygm9pX238AlrLex
IIKkkzJ7wG3llvwQnIBxdEJ7n267Emvmbw+fPDgINTYD3i/KrUFI7ZthrfXLcNF3
r7uXPndv9dp3+vRkvLOtBXHNAjEpFseAsFCarPXPN0tFlBc6uG4Zm1MBtlX1d2/I
es0HOWXqtodvfOXzXzhUEuTQ0FRvI69tjn1VeD45X4in6oXAOjJrIo2V7ESZB/na
8FzCK4J2EFNUAfVDMsrRNgWk1bEmrpCw3f90+u4RvU9jS/zykCByYFfpaZxbFkiR
nPp3aKIP0MANCiwDIzlYwz7YYnZgD8yd3y/HNluo5Nl3VYJmWI38kA+6+Eim9O+Z
9zyxbIg+OyhkvlgD16CVJPnkN8YzryNYjLTxMZWqthoX1gvPm5z97LO2GeoP3I7X
0Mgu9Nftgr2xkOC4UHoODg8wm3OnqV6gUhAdOVErxSv4BlzFEV660Hol+nJXvjxi
oL+FShFgdhNKuMNEF5vS4KKYLF/Go1HZfsia0VtSY1xm/wKO7m+YsI5/5q1kuiRE
/pGAj+B/UQboXbmKpfbSYfRpSvRn8MzF0sszqUUDIy1mqa3GLDrS2TnYBY0HwqTh
6OOti/b/8jzhNvSOUb/AoPWXicPfOdHT4hpmX7a2FPm4askKKQeIfVx+WiG80VRR
0XPEIRyb1cJnhXQikiG/QV+mY4cMOV8JsuO1eSqo76xB8oYY24eesalvUrsKMXTV
DOE/R7mdSV1V6TLyhryKKd86BFxeQLQHAj/6iW/5gIkWr8HUYjj+UrjQdixd4CnF
z/Ze+5USnV466wAPN5aWd/7HLlqJN+k+RDNQn+g0W02v7ntWBWG0qi6GL2oFp+25
H4RJmygTor95xFhO//AccxfS54kL6zWhiz2PJM0fwmaaYTY3ChVS0atbewXogTF9
1HOQG8Iq9SY1Oshdix/1DSA4V4VUYCthHZRNS3Sen5B4zmIlNspGuSmf7vCTmQNJ
xjzPWqv5rq7r4C8YnFbH305e5GG6hi8hLELs3Ba8+uFGLyc8dwPw4KViLWd5JuMZ
wwhKq0UcF3sxsJ6f5GKKXwoFZEPqEZgrQke9RhNl9YfgEXMlSavzZsPC5/DM8Vhd
d/29aB/L8xKme9eTrAbPyF3F2k1WlQcONmuix+F5fss2Iz7Afh7E+eszWKOQnOKY
v+Moj5aMgZXWiMn64MeYp3vWPQusoLM0OSwIME8+j2AGg9qjeZa+7F/EBdSCggMG
C39RK/nM7kNd/QVyV0CqSJF74xgz26ZY0RQ7FIPWKikucN6UuQLDLUWWeQdMbxpo
IvdUSFkEhAfaVTqFvv3EB1o+JsRmTHLliUHw/DrtYLX0jBQleYxRJs0ZKJNs1o/g
e1K1s6WRg9rGE3zhnmvWNapK1BW9LfUSyf+T4Oe2OhqhHAnU6s41p1QnlAzvs/3m
dx//yG6ct6F/7gucuNwAu8brygZYiYjjH0R+qmwn41Vav3L4AMVjUviW13JlPM9D
lFzrKw3rUkeqbhxa9r0xJz/EwJjeMVR9Vc0hOW1dXBa/yvsEDfprhLAF1cMpYqfw
Wu9g3Zb/MYPvy9Eou56tI4bx84/QvESvVoGKl0tCBvoma3ruIt/QwhMTGr1XVfcq
Yw1LfYd3m/p81BprXgdGpWLdw8heYiko+LSNHWjeheakYuks3h0LXwx4yzILWz3c
8H1PQvVCKZy+4ioMxw30tJRN0Rr3vS1o/bneIIN0GC3xfNW5iMmUtB0KApyv3eWv
YyS/IX+T+xXxFKG33dqZpIDzx67sa8/njBSZFjRFPLErt7JSQi42kcWqVHfDIxuj
/dS/c9hZwqhA4F7yKl9FwiNv3YdgBq+afKjsTYg9cNfwwAwNDNavhT6Mzl4SNVBC
QH9qZ6/vLhiBeEYZysU1cNs/ETZCwkr4ja2jBXhZuXR6tg0WOZuZ4olTXRGQm8rc
uwLtQ2EmURKNZR1+6LafqcM7ZhOAFLbKzmAH+cxMOyAzC+emir/9/2fKg6oaKMZz
RvNTBAeVQI70D+zt4fYHeKK+2gmJ06NUsH+cT21Kyx4W4dz96aKugsonpqXQ0BGB
FDHmSslUFJ5WOklzmeulhGwlj3NOdxmjPW97/7DvE8WeY+QJ2N/rnYafbk8ipeEP
ESoV3W/KAp262JiNbgwZdGc+YYm6mqzoZf95X4EryMsl8KjGPzBgi2c4AIaH+Mf3
o20FqZzdkqyF0/gv3EBK80vuewHMZB8UkaoqUtpPNr7BhqdaJCJaIskmyhB3hCaA
TmPg/RXEDMU8bPTBl4kNYR9zazqmHqDtRxIqqhUDIMOQOyuAdG1UGB1euslwzD79
cNrv/R8L9hGkt4PgH6nY0JxN09G0ijnbB3/NCxNlEsNhx3B6fo01E8uhs1oHFxhn
dOh/Rqj+dUs2145ZpSaO32tZtcy3tarOVo7Uru9/WVra96R4oJ6nSFly9uy4CrnW
GU5+P/qNfooS0n2UCyyf551IKMpF/HrVECX6gct7dMJblpoEzL2LXp9hEz+p07a1
67UKQTL5Gk8cjRefGYVfvIDuI2BxY8OTZYLv4h0yTUSm0hPCzlagzmpoynAmGITr
R9ml7MAX8qOl+RMtMaAbtVR6a/O6g/eJpgMf0NlhUGngSWRvE66/iGNu5eby/Z4y
704p4oIZly0chKF9OC/EkiDN1YWCfzWAN+lujkW24jRyyqB9PCmMjtZq9MDU2pXg
5yEdAAAnh+e3OifWe6KwVytCQaZaW0o5jTTkkJKzNWT8+up8J6OQWwyqwkWVs9ze
TEHgxnpzFV6O9pHtR14GGBsQMCARhUUSqtTvm9WzHvmklaK0ZHvxvKLYVQkdd+DK
7G/VRpwqgdyj88Fd5hJ52KBAd0k8KAxa3umJLfCKMrZL98l/C0B2O8CqVAFKb+V0
mPfZCZ39hK15dJH5+WGwHcTn/rPVcvSei/XE+GGTfJqKAPnR7aLX+ld+dGjOIqhx
C7hQnaMjs/5XilOt+m1lPjNqsFnfu02jRLd3micZp/RQ5weWfT8rLdOriB8a/gcT
UwQCjbnwYM6O4MDQcv9o85SgOqDKcQjRLcLF67eCjtCcfXQ54/bnuQR77JsH1DgJ
uwsGrE6j0UeYI4TeCetb+WPqzS4z3U27Ipi3cxIuwaRDbrP2gkBGz+aXgzqdTfNH
F7jenPTcR51BrJ1OuMPaXMDLbnxloZfcZw0DFjZOvfHLn+86v654TYbX2lMSXowC
dO9psMWCBX0CSS9+bkZ2STQzQ7JZg71i457oouVUCNrGgqmJ6nNfvOkuAHv1z9Bn
UnH7yhec4lJRODhtJmxLEbDR3b1S0qZUHECw0lAFqQzNH1Uun6CFDiqyGCB9hiPM
+j+3VCwMWRUQaV16ZIwMDFjQmj+ylVBwpYhB7fLpmtev5M5MiJ4uecMkrGNzGMG/
CLRdRcOZJIAuZLh8z5g7sJH48+P2aWAwMAC8Pe06hgY21JHdDg2MrPCT/f4RkTqh
YhjEsC7JpKZjHwDQ7Ei8GV5ztyt8Xvc005S5/oZI7QW8WZwsP0xUGXwefYCeBCK3
bPJ8UdeD++HCPP8ev04hwhO/EdUD4HtHVgzQBwato6ZcmpES01OdmQolPU7zKpu+
9J763RYO6mh4qo6WV21dSvLNmINAU3DImLZNeId4jYnTp4fw+CBwOnfavNV1Qz8S
Q/+7E1QVPyXuhbTud0JjmqJRv1qbAgD2cB/gb6PeXgKQeicRRPrZQoSe8vLNhMDh
8RLVpRgVmut4WGTknPRnEqDHHw3ZdlaHM221AFiYuhsmOgum7APagdtVnZZHKaLu
nE+HO3D6KBEF0MVbYVRJiSKQWYpuLyUV+petomHAg7PHapw7Nsn7qDFvQrh8ZDpS
MXLWBjTfTSQi4yMWCZd3w9owkbVbeVS5BUw5IjGlcVwVShAGeUEg2mqt1jCaJNoq
Yrjt+EWMrYLpnZ1gdsgzRafBQXg/BG7p4rsSWFBHWBnMkLJsO5+wpVFkUoYDF68x
591eSD2qLcGGPP7HVZfNvBlFvHXNi9Riq3LJ7dafbTTV1tVzAobnxcEsrSWz/rOZ
xdgrRj9OP2eZc47y0T8p0VmJTcOsDMzkRy/s5G0h/VnaffDl0VSUgyen+1YHwgNl
NDgIcbDSsVD7Q7dvTKYquKr2yuicN5go/vk+qy4K1vFfCHL4Mfr/XUxlr0dj/q1a
7zhP/NtSAhmsAuCQSS86Vqvk0NWTkRLnr/PXso9y8gI5CIyeIlSoEE+GXx8LPWr5
C1ZaeMItfLtrgIOKMRpyJE2UQGNQdZ6XaPUr8BFJitp102GC8syQmbABqyoiDxoA
MVaWesYvAzVYfPh6iBoV+M/siikY4I0RaAYf90rvirCa/qw+bpeXhIf5BINKAEVm
xxl/efX0TN+66jxoJqws6hCAr3Dif1s6VqGrUmMePFFA6jBcfxOPeu2+A6HmYCWt
1/if6EB6I4eGsn+J5aR5jzg7DiIpwTyxWKPfcDDhjXeQT0N5QCgla1MsMIBwpNrx
NzoZWc6czg7Hn/wjYX3YRlK2TBHnNcNNhrOg2JUrsnkNrk8B42WluvNwzI8YHF1o
mf6ZbRQ7OhCXgLGXkw3uTDGttHYtAPZ7mRy+/2MFmN0QKn+5eish1x+42hnIWmLd
U2jBIhuhJIYjd2KnycBpBJWjLmHFNeAD+BjDWaP1D70yEur3C41owI+zKD8Ma9CD
+4MKbtVUM3Zelet+0GsSp5Fxos0AbqMNa+ZQS6gGD02PJt2AwDa/NQGm40gb7bc1
9yUZWLnbZZipbjus4yxxtd0C+Qiudq09iOoRuCPhB4yur38uhE+WwLsN3YFJ3hh5
tbiYJdaO2E3DeAERkYGzIE/IreT13JA/bB09FYi29NrlcQlhim5XFW4WBrWvH649
DiA/YxhzTxT2HDtlH1sna51Zy4wzGh1emIfUyaDP/ilv1djCMePuWAPJvso6n7Pf
9X3aB0zJDM9PaalOW99QaJ4VXHKqnIP/meKiaR2dHjCjmuAvx5wV4y5nc6scTpSZ
Uu8sWk30rRTsTa6EfCxsSAeCNKjOTWrYa69m+TVKZZhXl6JC0OK5Jq+LBKvcqhJQ
++2F02b548ujLT6dvwQ0ls00/qyHmdrTemWTjHFAv+5CHuz+6UFx3JP/PT8qRLZ7
fTDia7RLtKl7lnoWlIPR9kihG8RZObdzLzYPyTSO7MYbR0nDMq9zT48/45B9lN6n
EZ/T8a7bFWyD+pj0IDIczu9GQFcUbyTvWbjRzgVxBMTh3yIBhOUR4bjjTuhR/nG2
BoqMO8+53yPg0qdrrPGnpYLqALLpwF+0xY5b9wGw35ExXqRmc9UREtrim/XKIugG
Irl5QegKIKZJZ/Un4oZr6ZXwkXsO/QeNbYpluGYubfENFU+f9g73jpP3e7VCKFPS
hmxqRmWkZRDdZuDrwlBSMXF84JmYRcpPrcM8Sua7lWmDvuxkK2R5aRRFBxgYrV1Q
0KxO1jGAldUPsw9dj/VG7B9LB0QXQBs9om5oON++XzsVZeAza36Bc5g/2y7Lu+9A
k8X/PPU+bo8R+dfyMMXmRdXrfx8FuxMGv96dSU4Lah06JZuQE/nUeAWZ+fugo/xN
CowbYIqo20zowStlJLwBbZo1cYM9tY3Ksv02J5OdoBi249ppkGnF2rvgaNee7H5b
kaxqJ36ZR+X/I4kVdgLmOTAJ4lklk1syucueZ2ujyNJ2MFugMUY2La1hG+kUM3Lt
C0NjElNjcNbmAHI4yhJvTDDS0Zor0v4qyrx3gsHxTZ9N4b+VvgcDttewCXbdk6Zl
N283nASqL+Z4iEo0wdW/nJopAS5qbTRuQsA/hRafwsmJLqkP/hZZEY+BfX3mYy3j
0ULUgUW2ykDGnhs87JdcnoqtAakbsNRbPO1N2eb7x9ym1GdjCdM3SU8+FK/U8oOC
zJ0XX38nmQUCoBw9qibNHe96FXGmutVJ2N/3vqA9N4fowMBtQnjp3Yd9YnttegoR
WM2/6FnkUEu8EiDi2hVt4twvDPlbc8bzaBt8Y4I80kMMnm3ZMZR1lomyXadvpKd0
wKyjr4F+LK8jEe6CcFTdpgtfEIVH/6Binz8JByv0B3HQMjTolL5fhxZ/9Qqg100F
xGDsCuTrVFmeDkq2CGLOp2DX+gfN0RmA0Vgxw7N5WGKpqgfRacNyIQPHbzwGhjuv
5AE9d88A6puUzo9Vfslx4Pq0dtlqJ16NzpNH4Yh+CZseOIWCEalUr9ZrK9ljqzRL
GFMOupkL8QNW2r0GgeiIjC90NQ1hPL/uy3lrGLCF+geCyHI8vJse6F5L10IzdBcK
rnRUZQWjJQq/kSBjAjwKxjPFXsot6UfolwFgtMFYZwj1sq0xAeiiiTL0pmsaHsw0
7b9O7ExHzS4qbIcT08dZJI1tZcmmRGPvaOgfZnQo4qNw6oH1McaRqtxtUpnUsXBC
DAHmdr7mj913szhB8y1JJ4aYVyUwqu3KEMxYfeNDWABuBEOxEH7EQEDK7AWUQZ2j
CZa0nHoO/Ka7Jce462CvnSmnYBQTOlZEekngNEgVzhHz6YM9lzP7eNkJx3AfVBRr
dbXKE+xQeNMwdgsadY/wL/jdIjALgqy7nRK6lLd/KOgbCN/aJGGzOcpSWiJq9YKS
d/yMtTKM+EuCPDRJ8dUhjL9knBKv0Uk06Vg9MbkTdT2n5PYP7G8JAZbL1ZT8+qCR
AnA312WoztYpN4/3uEq4KHEEB/viV3Nc0bHmNaDU2Zva3/mkEwt7d0uk77qHQfbU
hRYKr6HtFtfpm1MTi5iGyKSUHP8eiCxkMg1WIcjFWFCXnN/WwwM6lQctVlbYTPbo
380APCLg+7GCUqVNU3RvdoMU7wYygim2V3ejTLfly7A1mmJMUMYBsWqhTDpDN1s2
NXYmnSWfGrRizLIAlppSu5uRgFbp/eKsKCOYEeRlefMYYeTLjpnHhjEg4d+HHdKE
8ugj3fQJzODUfgoTrG0+T/etxNPmc7bpRmryChsMiPMm5BLrcBGfGvBBMw7dq5mg
/PxSknv1PMPRvPKW6K7aPAXym25kfXJkIh7PyZRhVNA/iwbPoHxASo3pa3dkQay7
FaVCNR7BK9o5U66CBDY4VRkjlBb/v+evd45aiy/Cfk8r9MLawExEIKZ+c7YsN4ry
EpyyEdbQ5BSVO5MzSIwcZ/0jH6n23HP03EJnWGudwHKayog7M6VxiZJesnvzSpN9
0hgZVMn86/LlUVmSXGZVmNMYMaC7X07jAdQ8xCZUh5Dno8OInHNn/W5AATNg1gV2
pAPmKnYWaVJQG5FJ1cdp2dZ27aa+BX5qaCOXnym9Ttzxr87rQ21ZobDYbYRSoBP8
zP7pBHd+2x2M9Lbk3opUyDkpWlSz3MZga4WU6WA23Evakmc0w17JpkV2qDDXIptB
oTfgHTuSy4/kre90YwixBLThufwVmid2Wz2R2PYWBYx5pM2ezSUDo7vUMMp74ZJe
12BgZvKG0xXPXzWo9NOxV076c8YS6v+dhb5WcJk26adJGFzmpP9W4W4DyQ95/gYN
cR2OlBS3pm9E2uUDXFKJrwjnXGG/EVMD80vAbYIR57NbpoCZ6XadXlL0sVBUHglT
kuIf2KqeqbRKfy40b9v1VQdbzNUolUvkcNCwDVHx4wfXdknpDmLyHEbzZXRGRN0w
I1i1lEG1enXCd7fKhk5p4sCamXoCSC2yyPmDmFb9dRHbb+Zf6aNsNwGfgAxE2g0B
df0U/l/kKn+tkyFV1lxwHQ8E/CPJ+eAGIsWxctSyYaxJZw8h1kZVZeS5MMjgMrJT
kOCUerHAtvN92yT/bJ5V/pwGfg0C5PRbTE+vNkNBNvW+2V/+V55ALnaYhHfJiu7v
74vtdC1Io41jg/D+pT5Rzk9OYyn3JE6Me5Osozy3uSlZUssV/KW/n1BOqLqfNOQQ
6HAtwet9yjyUO4v0axRtYLHqnVNED0JXJDgIQrGeLK+6kQ+M6LnAzaQS2fDaCpKt
al2OfFMdXwF/Iwd5Wwn4qWoHz4iF0QHV2Hima9m2uPHTbKo5lom8+3dPZqqXqcsc
yI2zfFOFnw5N4cXFWXkrfQh3d8q4QeutgjX+8BuBPuRS28tTWP5FXgXZbn+PYbMq
71DvxcWkPXLBP/9yWI15jWUiPfPCvXtV74fyS+llz/YrIOIIY/HZyCq8FMraj3PQ
EHuKWcKX2++z/sHrMNIeo092Dyh74dIKan0EHmLiL8PxgK9FifrmVv2Cgs2rRgNq
vfCRbu0HxKuay0yURxPVnyTLp4Df8CC84NqDFxVaf3D+pr7uOb5tt1H5WXBPiFgo
xtEeEuUTYTlcHEcDIEWqWlpWa9bK3Vi6xBi3P//3QOQpMbty0YHTg4Srkc1DAsI2
A0B9ILRDSsMBU+covMBPJ++ptiyXNoVZ8UzLpBK14tQzb+CUnM0eUfsqmbegVfNd
ZCx1TMUvBYk5m55HiNp4vB3WvQEFF58ROOsLs0yg5+VKmPQV2zZJBUmYzT4YkGUD
SYY3cKRbsA4FuyZ8EP7aRP8tKjRKWoJ3QZTOkMC15ihtEvKYibJP098r3r9bi8gU
1mKDcGuwvtK/cLS6XNYeTUWXpD6ZhjghcKs38s+xjEP5JfAXlQspf+7SF+sD19h3
IE90kZ+V3/RPjooj7JWT05EjhpO/s7hx/d4wUFvPMuz4rKTBl7DdSh1kXyFHB5hT
5ZuCKXvixbbKw45UF8IY17gMLcQz8X6btEtlXfu6YyR7k013/aAq8vjZUffijn9U
xebIRoDBN7UaG3pcBNoAH3kOTZjb/EDFGVys3nhjbPaDoHMosKTKFKhuEv7nOEfK
tYlWZAEVg4wENiC71sVDp85QNOdiR8eA3xer/KbKksFkX/Sk8FBm60s2e52iTSv6
m6Apg3xr8w1d9cwCDxKITsnzCjZxtw6BV7EnI0Fk0cJjWDiq0BNDyncBvTEARXmo
mhfkgpc7epj8FT4Hmj1+bhsedUtofMPfP8Rfj+sobiSPmgWUWERqURr95aOULwrs
lwJIBcN7Lzhlw6fbLH3fyAxp1hfKWKKacn7j0i1Ba0z8WBXt/LlQz43DcZT3Axk2
oBdDtLYOTQ3LXPj8vjLUT3lbVte7NrXeGGLZJaGSJPdPMzwaqvpXSkzuQljlDSM3
0jwot9v3h8swSekntpDV2vLnea7bhmsfLaUzhjmSKsbpcXJoNH3gPHvpCgQ5YN0T
keZ2Fj0YuzkKW/s/o01DXKxZ0+HU+f96229IluV7b0227epyXoMkPm86MqSpzTHg
luFBmesPu0pC/iev9rmJeZOpvKC0TMRKkR59Y4l5eXSTpFReI4kMq4yEnD7ZMtbd
ij86Y4LBRpqd1FHGcnG9Mw1lGJ4QB109k1Zm4UwwTffWnonGaJiIxYldA16gDLhW
swY573VgDoHUD7/VNRY+P2unpqj8HWP0NVQfwrGeC9H8PamS98/y/jgYLHCH9/jf
4YmN1bRRHrETimuZwH4yGH10wPLSVzyT4hLopF53OLlVh8rw80kMflpK0lirudEw
UMfnSDg8GZHL6+E0TUOUIsTbhT2T04r6u+2wJ07vmH80dY6Gs24/Ad4Zao3nOaGn
yOpCUgd9lVctmCQMN4i6RJ8HwJxxX1XiGvaAjo5tA/8HERLgLApREHDOWoyxdMYz
neOmIC2bBukA9/fC3Kdj8KoEFJ+GKOF9CErZrwteCKvu3lH2DFoa4lxDhhhoDgVf
jAyYp/pHilAX/cR3vl6ZVdOTnXcuJRbazRS3nOtUZ9ga6hCoMkxITUdKfco0KoJ1
2zaOadHiIIlghZIgd72RY4AdU2dxIUQcSO95tuL0Xbtn89L2G4ng1T1suCSkZ5Ip
j5hOQe/mQlsRTREGpT8lN/tC50b4RMbsYT+W6ykqbmPGF+0DTc4RFUFHfT8vSbYu
1XGsA+y2iWkWQBRvyH+lvLxc53Do9wRhxZ0IyLUoo1bvYB0hl9MUpyDkT0mJrmlr
SyRm9H8EKHVE2iMj+vpwqysMChOGSzDXHnDrhQAQ6H9gCnK+e+mpphc1LRtNLxnI
KDMqroZONwv+Awp/fcotOoab6ptk2LrJDWlVL61VY/Su9sYAtmeh/JISRb6H03Fq
ZIkDEfY2VU7j3mQYGcKEZ/yBitVu1BxbyimCkeRkM3lfrv7xA4wBgCF7UvTDmDgH
W3gypYR4FWcLhK92ogdAcP0d7UV9Y6kmODQsbT/arChampnQ0foIZItnnQS1GX9/
1PTaQeYcuv1IFeI1xIfiBx+zJukkR813kip0yMSyJJphles45IvUFFg/XhO4Vt50
1n0RTFnb5Zf/RD1vFN/0TAQOXuaho7erM5yeUH8J5s/7qZ0EPlj10802h3e8PeHM
dfmWjuOICWtxTduNXGToX5a9+WJN8dNym2rxkWKGriRu0K07BGUlAdNmOdztOpLM
4BK7YMNJ1DCIESgBQkyxsSLbYL9R515JuwgrHXdFkorkcpB/kMmx2Jsrm66ebZop
Kuxm6c4OBc9cfgb2y6L5f9WRF/A3Z67hfAwrXMg1c8qL9UeJeDIZ5EFCIUH0K7VV
KdANAjTVAeSCMHIy08b67aZzex0COQTB+vr5ch1CSF/YEtt3+zr/TtGR9bqRsA7S
YWmoo3CgzrKFpkYGXFSy+8Hh+QepT+RjxgdC2kAvkd0ZMSXgAvKG+vDZRDaOlzGQ
U+We0Sy381fF1D7PIBSX7c+eAPTejSvtZO1fTc55vl8E7gFhSkhf+F4URCFSkvyK
z2nbHV8wrj6NLKmlbuWHGGN2A3QXxtkUgIGpi6D1LfP1HhVthSjhMvz7s9wgnrLf
R5M8mWAj4Zm71SYVMtWOg6GsBaIjkXjWfiRxF84ghOE8oVkM3ZaaZWH/UwrjbJl9
iOaHAGiKw1HTUIs2FCMb/P7nxXSue6LlW2kP1Hlptz6YE1EH1MNPq1vAyk03IKP5
Wpnj0XItnVCyM33GJKKrEPy4O/zlxAmxY7aWMVvHd85TVk2g3h0JUGlnQJYAH1yz
jNrlGqZF18aYaegjD5biqrOULa9gJFjQUiDsUELwFveUwwHCFPtUpxmJF1kd5FvP
quFXR61IHdpiiK8Fl45kdMWBZmJy2rL7Gnlh+Xzynfz7He0BnCdMpCDmumzNa9SM
KWfQ3ycCwPIo5OT0mBlQr58bv+nsKhIZK4vfwbnJ5W+e9XK3//Vz0fVyQLXl7CDP
vC7o5lLR4c0r4NglZI8nkoI+emF9s7mtQfXE+P487wgV5q/5Yxt3DMHFpXo8C6eM
/WUfKb08k44XN9aVT0UYgrGzXYovK9uYn5zqdkqaEMdHgO0mrLO2yK1gcGiT2hyL
7yLK7GF0rGC4SnLkp/CFoNdCEr0BUwpc78ol0HX32enaB3rfUpLWE+XjTAVHaWDo
1GPY9UFBQz726oIUy9wbBDdH1fF91lqU3tG890T5yKZQBt6i1QsNXUM8RvHXdXJW
8jUjdzWlh6jZzBVJP3ZeoorUbxPWhg1J4WmmWxIAC4hJY4QPfBHcuLV0pH+Qzc0n
JsNQybNFre6Prnz8zsHYDrj1uAKgOmczwvv247sYlafL3rWVu94Ns3n00f7nXoi0
3EcTd7VQc7uvH+GiUjdLccntt830NCCtY+oFfRAxNjoW9WKMq1X7cknnAcEk98/m
aNMyiH9U+tEEyRHwqCOgJw34X9BxqEG7vR6PPAiA731qiOrsKOjyC+LBoTRgTWmy
VJ68QXffSurEtyxDD2hMV1lLkTU94afBfSjZLi8UJOcAUHuyOdNp/akR8GTdtCxA
FAvut55Q3kx0vd+s0M37Xfa6oEe+2twq3zVssFXoHlXsZIfvrmz2qitIQ1kBoYsk
AbjpehSeJ1FixBvQ//PTyST4gIpdC5GAFsBo+QJYNzHCHaL4+/SG+vf98q/25tq3
8iAydqM1mhwWoDJJNdF9251Vo0EMUaebU4uEts8Ie3aplP3btVZAHOxSaxguDCDt
ZW4mJiivVjbMezJawASRFpprO0oBQbJia087jvYyIhFskxXKFIUNpuGZO8kHu0WD
B7Fcc0gh4wP+Mz9QNY5fztgcIvseTlPJKxiH0/DMbs8U+foh0WmZri8BHGEZdeS9
HzefRdTuSTuQ8OC+LvYIflM1hhcakYuFpyu7XQP/74tpPt9jHaTbLhVdbv29ZljH
/BBx6ogKDxfmdj8+GUZxGt7Q5SsPGKrRgqwk/XMsqg+5azqDPD9CpJnXQr8VShFD
181uJkwfrxtD4KWE8oK1aloHHhEJIw+oqaL9eJZgikvfZdxeaGkVTGEVI0ElL/hQ
egxjsXZwIn8CQysN1uERM0DJXlEbGogF4onnUdNAjbBTq7Y78N8Ty9CeXT467k7d
Ew8OCgU4RCyK7VGbw2qFG9GCAE3IlmEwysyjUAWRKpg5ji3FjUqPPUIWx3fKgIGf
t49mVqB901cWblW2eTzU3i6XN21+KxE+nGapqAjxT9r6QnvEcfPVv0L4+dBSeU2F
eEatW9GdKGs+ODYm7BmnKDstqMR+ST6h2NxpH3FTaBTT4Z68XUrFH8FWZBzTVLsP
W/f9vBZrYb3vnb1E1dPgXTaZONjxN5+ldI4OnSMMRmkKcQdt4iSjslA/J1aCNELK
OOduHsVAw3XVeqbTGTcHPpkUs4yJc+vaDlgL62ZlWOHvmwTdvaEtA/6XoohwbcA6
y4tcy9KomFlwGQmjoRdWq/yu6yoDO6XbAIDSS3+llMIauPWtU71tact6G3cyA6Z5
mQuqu74P52Nwy0Q0ExNdzX9lqJsnPetxESTiDf/Yqdtbb3uKNDlazyYqq+X5Vlzv
DxHHeExNQ74t66XycKUI5UgvS4nOauMdrkdnAulA0JNBP88yMNGblAcx8/Nmrd8n
SyJXHxP5WzagS3kV4nJ/+NPLnY36xt1NxsezBAKfvmZ13awRW6Oi++u+YtEWsiQq
9kxAJ2AOS1pUGyS+YEwolTXCAkNOfRTDC0o5E+q+bbvYrdLkeesuPg+OsTX+gR7a
5miS+DRgzZ7MOowP8Q3518OH0nU5sfqqwyCSXyreVMdLRB/Snbp/mF2BVUoVHsIF
xreagRbIZgOxA/9kP50DKZzRhzKJGPNLt5kNT9zyFQTJfJNNFMu+PW2angLkUTHG
qLZXzHmfhUaxDk9VAXi7N5PFxzWYe4pEaED3xgtszJoVJxaGqWb2nO3VxS9IFNUv
uRodIqFrR44YXVFii7RbzlqSpxT0zwcJCNILAtx9KjJQ8K1Bh+/2voR5TISAeaXy
JAqL/xjXP4IyZ1KmcERwFt2NV44gumcTabytVy4jYeo6IC6H87x2JjnMK9ZyOcMB
`protect END_PROTECTED