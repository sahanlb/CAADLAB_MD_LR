-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
hYJ3vTEi9CrK3DaPtba9iuqxCcJ4BFS8NWboP3HnAEhQ56llZZrPxeLSnMS2TfyU
Nbgo8QJfR0+xl2Sl4t+Q8SbEwdHG9Nm3KVPzMrjosYT+KM805ywsQj1GfCxSP2Uh
4cHYTNXVzvy5vL9GpPfXpsXiP+eX+58JYH7TcaK2kKg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24915)

`protect DATA_BLOCK
7l9aFTsxm/pWtHdKeAT++1Lc3v/oXECkEmmu9X02Xz8UPEUE0qeIjsTSqrM3pH4f
wSwub8no1b9O2qGsZHNVz/kdq11xfJg0rX2zYt5BQr4lNKV80lEWiFiZaBE6P8Wg
LhwUDi4hvvA7OHSfA/MYoRGc1ploR5Vht5AlrMwwFeJVjs/TP8mxZEdx/vyeR61B
GrVgiInpadeBfO9w9dzgwYYVSBxMJTn9u6MsmRhRxMa0xs+nrOfyeuqWt6B4qXKK
+Wm2YXobGA54Jn4vVSzdC56+qlf4rVOz59xXdJYY5bcT5TDTiyQfTmrGKRNK+mG5
2OsD8b9UePt6UbgsRYcS7CJQwrGHIzhuXYuhyx2anCnVR7orjZgb2cdzJdBvLtTL
EPOEzURUmxzNYuOd9nz+lI8oDntRjFPFi8qe/7sXNH2IOW6JnWdqxTHloz12x6Al
JEPo38GscC9NowuOy7actqLRQPq5iM+iXMvMOM7swLlu54PVrNRiv8F8Ws+BglCV
9Sg9PiP0rG+xTYq+e5OlPVsVrrY8w1xyvKbzUa6EVlnDf4Kcz6BzrGGH/dHS6hsu
4GHHGUTbugnXxiql0s1GUV3hsLxa0EIDU4YexEclV9PjPZZvCPvWq/87JoOCfwW6
NXHCNkLoAgYpBqsQdWgeDdNllpPu8S+3ZI4XT+Vl7or8W3i5gVxTjlFEEYBDiidM
VqQM5PEMMb7MlQoN14rXZed42aZ3mN6dHF+PAKoVbnlqoOW1nOls5zTYZoUqJGiI
UcxkPyOa99ErDt75aiFbIOIn7ghN3GtSPXG37hPJZX8mpuPutNK6fAUa6qPp27gK
hel7gQ/LE91JLmF/odHECYGAvrGbQCepjDeyLEhvuZLUHiYQ47VZkERucNZG38Bd
2PyrahFfWmgv3NVz4rVFnaBe5IYhP6LwEB+rKt33khepedCoWyU0bCWOktDC9W7g
CqVgDyVxc262K8nsN2dV1i+/chdLhLNPzSaF9uU4qQQmh3ikAEaKkgRgUvoE/Amq
Sq4idOiXkM94WxoiFYhir7PngZNNq+F94BIhCpKxtZPhQP8R+39hmJF8osaVf/pT
zVOJeH0hLNd0uBEXJU6AZo45CcWhwEOFkbJPkk2t4qDCZhdfF2NAH6qDiyvuGInf
fCEQkn3Y21cg0s5YAlR8PGgV9Rrpkqpg4viLgMMC8/CpFRLeH9K4xa+J0/+D++B/
mLnqhTZ81OSPgYvxiy9AeNiRdsfJVy/yi0i6jnyfJ/WeRqwsdB8uq6nVbnzBHJsh
KPMxgiRpcWCWvmsD4wnkZ8SkxGxRmw+a7ya1VGVaerd9jaZFhQR/uz0sI2sLWcxC
5yDbabJdwEL2PcrxuXLwV3JVuSWjLNy4rw8COBasiI4Bv+4NigplyCXEFaD4E+4h
vAHD2OMkEdQkHh3Y6JsEsYDmyCTh9haAs77q4pvMprTiYT4j3LLBRVxP9pI6hjCT
g+Wuxi1kkv3SEe8QspUp88k/UqysFDitPDyjClprwXyoNGRVo3wz7FqTgfUfDrUo
RbcVrQ8faQn3nfn5HuHjsmXBIKW5Wbl/w9FGS08oHUAzOef8bGjjoq7oYhnrIM9J
2CB02l6aR91XBrVjyt7zXcdrShQy6CFmLq4S1VY+ONa8z4ZaFJ9WB2jaSvfCYhxm
JQp6xSuQ4KsK7s67i4e7rJa6nqm3I0amnNSDjZStQe6Yb6t66Som4oEzChhI2cIz
CC6xm14ip/yGLIuRV6eDYwNDTnUkBa0ga5Jhkd270Dqgx3M6Iud2g2JGGfcjMths
hzlA1Yz+CrrKDz2e82n7950CzyVsmvnqfJqKSsZeNYWhMRQVrZHhEmNDFuvjjiq+
P7kkr60u9iICJerVQ9i90KsnjoOdX3eCPvxjfpFq/Ms4uXWwjKQYR3lv6Ml2mnsT
YrsHRQBeu8c1ceE/3I0867HeMnP0+B72wWOmZt5nreZOkCN4ppzBG3l2Y4qwPPwQ
RXO1SCB1/3SEY8wHMpn/14PWRC+na9MI7lzuAeTyw42p993vFlhvz/dQkvxJYnmV
9vWMUSP8eFZdEBjAENvNdFmk7E2j3fPr2yeNYaRrCa4WEh2Pz5KS/r2Gmi9Sxi5P
Bzp8xqABwKQ2ZOExKzbRUwf/dHNogzvpYkL845duIIOwrO4kSx3TvyADXzbahWgf
rsGF+C15MuRkDj7rDvAPxLp0nNMIgpTUxOG2gwcWZGqHGW8pMwrHpW2TLQAf9iQQ
6zKtxzMGjRP+2pQDW33T26kTpYC8y0sRofg9MVMWvYy73ZEyROwhWgrbrQv0I1Eo
QwTLPeUiupCnEgwBhl4L08ajP37q/3x3dTrckGQF/qo3I028AOxi2818qhEhCvq8
PiVmkRGLjDW0NTqNbM01/2D7MwqfM/3g5ehS8OPSAOWuBWM4RgJydG3SX1b8gAGK
PPVe21yNQZ4l7PF1oKoKG6PxxH7lkrq5P77u6KztsosrQmifKBrtJBF1Pkd6RLjX
gtEjOvcmRSrKT9fHd2wEYp31btXKmtbsrefCbaGOGnP6FOq71yKz2Q55e+D6FuR7
Dnka9NowJZDXjnQYZ9rL3/+ysrfN41yVL4+z7Lyc1hqBzseQKvKVOR3juep98Ph+
IGzvwK8POzxXBC5ZjcZuQEDAv+Z26nirdo/PPbsm3IAIG2JJ5XBxdgORehipbygz
w53QQpRmIAW9a1C4pJVyO+DkiHUa5SVIcsW+ZYHU26KJtJl9nfgIrrzcD4CsTeqE
t8hQ5JfDZOorMin2dq1edO6zppO92KNFEO+ep6mTqUO3ls2jYg1CzIirfNA/eRti
C7UOmqOpFE5JS2giu+jslaUY3kRsa2gf9Mbbh26uDQn4TGNy+L2RHFavZlXFIRHu
ouUeQUelqaeloYk7BjaoA/RPp2RU1JoAMI8c6bW4uA2PImBzowzwH/iJPy0YFFhy
xZSj3X4pjz9PD6dHGkE4gzmuWaiadgjPxJj0RlgsX4mko/2LkGAqduEADXiL/HC2
eypCURcEHIPOMX/2ziCtkVCoRTYpHm88LyRH7LGCib509iW9csAh0virWZq2/t64
MKqj6y1yDAbsf7lVxzbDlh+uhXPHccaQVu+DI3G83Bn6N78TY8utMzWBefb7Kmk2
RYFyCO2zLTcpPWdxJ3OtX/ZXIvNerwaGwyF67FXExnwCcXidopWEdy8fN9Q5ce7V
NuLEOnRUkx3m/l2ueRmCpsCc66lL8N42oWjVOfmU0/yN0uGZ2DXoyBS0DwesmsBj
42L9K671u+DeWPbES9sk8hqXnn89rybddj/WVxqtT6kAmyaILxf6AMv3loLAALVt
qRDpPU6hLHy6nHQ+tZuGUj5xE0RH2LLUq1GmhkXArMJ51PFU70PWppz+cOb9Dm4K
8uTieY9dVdYOWIiYMEHD6AYDuyAm0XVAkoLCVfzfT+pVQkF/NUwO9V86yiVqMfzt
KKMUvGDD1XkaHUDjB7tq/xpvZ/y3k6dbRZlbeZyoUW0kM6Wl4GwKe1PmtdAIA0px
5eCCqDsMwHnL9QMriBAF0ZkTr5j3HV6zdl8aWmnyEdK+M0sN9u1fPeFzQu0mh9Ei
mNx5v04hY2O5uWwnamhorlU6aEwR2p1JsLq9AkH2mARZ9gTE6Bqa2NOwmeVeoyB5
28mc7XFA3DgiNsI5bEMKooGmY6vCts8krzCCOxQA5Ym/4RoDVOda6BEJ6b+FzuC/
BmvxKX9y9yCG3wo7ID3XVq/7XSe+tOrBq07ycFSG4mmo251pIjTHpemZtup2JKBq
PAlQfcJ0BrZ3O2brUmwclEEgRLUxNHRl/XmXH2hVc8JLxl8GWM0zAGUiwYY3GqBd
VLvvMNvYdnvC/TMGci/8DB2dJJwPNKAnnKY3yhtm+PpF6SEa8qOFCMHp0oZCEuTl
1Iri1Dt0Kr3RlsDz0aaVgrcoakTpWGo2HufQZ5D0gOa6OeCP9y/I/pdcHNDT7Gi3
+BsOwoOLyQJLgSMxMSTzNC3QjyFswlZJ/dAtr1Mi4GtvafxTp/NBBmzJfWaBYVHx
DEksvPERcopKcHF+rp7er4aH6pAr+fwMri8fuSmNW8xDU1EUxjZRYErZFkubgWYr
cZNwE2Lg3FsWoZSnUTAGgG3y5guTYOvhk+kqOvZ0dSh/nZWTgTNI5ZjR1n+JOgPx
JU/Gf2BH+YTRZ21Mrw0nsgzEECbRik4imoqK4krrmyJGJKLq9+mK9OIumRFbusvD
IWkE5ZUCSLyd4TKswilwjEGqC1vlciVJY7125AE2NzMwgqFuvnC9HE3s+1bu518N
EiU0QHpUqmSrHp2QbHTiDgQkWa67aEMorHb9U2nhmyePoiwo7NNi1K4OSR6dHp4v
etcLn4nCZozbRRKbVgIoRJw6Ynww9bv1ph8pivTt8Vlz1jD2rsDWIPCOVLC73SN5
/pHy6PoqTn9B3cRWuHfbkGV8z3VkmCtudgQPBhRIvPjXaOtyMe2wFAVFvRoOPcxy
d0znoK6IzDnVQjKT1PNrKbvAlvdO2J2BRxMJFBuWqt0KoGJxwCxsuI5YFhh9fYuF
f60C2sNQI3Wn9JB8S5CkOtXe2xENJBzyTUO9eh8RfND4WZs5ZDvdS3fUAbw95OKE
ofUIui5u3W+K1y9ChX1YqJwd2CY5SWrX/eszqSoEd8YQNO9MC6oCgw5MBHz+SEsa
Qqvt2joI1AIEpptWWK0zJiAaLcmJMi4A9UIT6a0PHX4E5uafOeL8xQSdldU1sYmS
A9NDQ0Jn1l1VcJooebeX2RKAidi0dQ424NxNRntnuN1/cAgET4LRKyi0HffeVdW8
vTGREhXqFqJXZiQ5AUNcIZnrstNTncE7/XWC+ENzHV4F40SokggBxDfFLMZMQ/cb
qB9c5YCLIZRLoaz+e5AGFsh6IgKKsO8jdkhiVxV5Fodfe0TEc99tG1l6yNIF0fw2
BgPewKBy4mH5rr2BTqQKoYhprZPWyiCoWTdzTTpcJutFh8X9LoOWGKHrZo5Hqd+P
M3EAhG5hIrri3uwG9xTpAtqvXYlXGFGXNfmqLIp+hdqr6/IHEBTvj+683AX7ix7b
mvkDhJp88WTkchuHxVpO8qIV32P0klbL6qyzFo7vKhf8g+uGfAm/PqjoRQLOlr9C
YXwWGrdsxdxXAtG+8U9nHchlK8nR9gKqhBQ0AXuonZ7f9HC1tBaGpCHFXPHjLuCR
zgGc7MZrD+ZvfNK6m1ykYFxxCdtmvrkc+5i32Al7ZqeCnRndngA+6myPJ0O2ovc4
BgTDiG/f5XBaer7hG01/rDxMab/+6DJXLpLQdL+823l80RfdWvFAYttn2Ti0XW1V
UVulDJ2GtZJWMXf96GImUxHEQBNeLvOU7RREj2tGl37oGpdcFvqdhtbQxvJLqr50
dp6MOmx/y9piwa2tnLUckqimxxZ8sPms3hPU4/Cv3UIvbCi0+VQ0Nz1JIGjEAzId
EvCjazocGUi9w3XvFqES2gVnpAH99mnPAHsqaTDKkyEejrGIO0bZR/QEqgIW0v5Q
swRcRjxowmSmix6Lm1VhTx11/CUXTlyeBFHxXfOgt0uaMa+wunE0YrIPnLwR8u7Y
S5HErNOeAjIh0xaBwVQoEgUJC4zqrPgy07Z/6sXq8S2RHyjYyOtHlHc0BUP7Mp03
Uz0Zo8Gc6Eq+jrxiOhFFI9MlCsQihkOvbkaz7xGP7VfqSaDjDog1fssoYV0SNyA2
GGhWCs70g2syZQ6MyaKCH64xa98vaKRrN/ptlZkQL+1tVRQA8WsuSfBKCBnuz/mq
h3icSgrXbFDX32CrgZTQ2DmYnfX1pNL43q/HZO2vvNOB624HotU3y2cmoOR+lmSI
n8BwWPUOlR6e8/YoqSEm/DkqCMLHblkZPSe+RZoxv5SF5aHe310gRuPUOaPkCRle
heneJZGafaYt+zRSMLouuBE3CRabFAihsTEuOAdJNS49zaPr7zm7FVpawJVl6cm3
KemX+JTheUYbYQFiYJDVfqbiTm2fC5akGK7srLC5ECglCD5MEapeHImeFmApVSE3
R4MNOIOSHFtBbVVBZrOGDzbYYuNC4wjB8OnBusSuZHFtdvoXlH3DlRIGV6AGfltS
enTViilbmB38vtyGz9g3+Rs9hwrbd7hcaSxlIY8MSgPtMQVHg5s4CsbfMk9J7TdX
Gcm2IS+H35ByFJG2rDYzVW6yBmxMzgbMQTbDrcVgHzKlMgTAQzw7pl5tksWenjtg
X4ES1dP+utZEWEv4MZMI7LtUs3mJwKEZ/B/WIR3NJSz10YNC57cZVzShTqRKeeh4
jmlf4rFFkVBjWCnwvt2ZESncZ1PQubrenGoql12qxvLjalopRGlnO3nqWpG4iO3t
dJzvCpJZ4zeHl/qQoSXdihaV9mpRR+2+YdsswFQyt/9xAs078G+OYZ5K69J8QCjt
FpFeYmRZY67KSdTQuWwk8ix+5kNZf8+5+jx3pvjsFrGAde4+3MozQcvGSyZOoV0x
r9VEg6IlQ15sj3cOyXu50lAoHiy5Auoslc+VnIFBK6kBO9T6Z6rUWC3MLLpg930v
+qC79VZQ9oCqAFjx/qKBrAWdlSerQhxAIf59OyUYGiY/OLkhS/TiySDrtoJHH/VA
FR/SwOP+2/haJHdda4a4I6ljmtrUSnsFRXAwq634a9TA17uZYNQZvWS7wq0XwhJE
MdprO/fgX2S2Rs7qWeJI5pXwZ6oXIIz4Edbopoy5L4ON4pA6BZlfD4Ak+UsAH7B4
LBEtNSA2+qEKcG+Zkpakv/6D2blGyUxqij3ZqfLaycQMwLtFaKe2qk8UmLI21CIw
Y8Z0VlwCJsGLTyn4H8IGwGHYc025WqAew6J0Dr7w4XKuR1OyEuWq/8eh8s2pJ0YR
t0My1RHrKZ4cAzzUZoLxKaJAm8QrIKtj/OF4LQF9SQ3LMUPzHKjhropOJzhe4OaN
8uDhxYZKyDoeZqX82+VAngdi+QJphmAu4hF06UMhFs5rtN8mus2Io7Uhd/LYEWVm
6BvRSFX6HD/cP2tTy5WRppWvUrvQSs/Dfk87YFhSEkwYr0fp4IsjNKMhHJ3OMg5M
sjE2M7QonRJnBHCXqBUsLz4k2SjvQj9bsaFPJuiOhOaQEhJtTSFBKjgstKveJREZ
3Yf55IfQNxpXCmk87tNuri0ImMBUm/4aEaUkJTYkNVnaV45npnwVDMxqBM7w/S70
Ijp0Y3JHoIQHlEPUyU5ftXCdBsD3utuLtYWTB8AdubJj2w7ylngXsLhIbCRLkmfC
UblTY1Nsn68Oosqiv290sVBXMm179h5iSzCOPB2PYeGwMHUruck19bdyYZjVYoev
TVh6yvbuqV0V5iUIjZJIWtJkwMBJ0fIQ0Jm7oxYUQb5hkVYX1Udk+yQSIbqatGiM
plARhoXM6X29gl0jLex+XijfZ5D0xcDRF9z2AKmULMRP+6urhf0jp3jw8N67B2Nl
QFgfEgEjWZu+8zy8cVFoKQ4J00AprcFqUenzWpyK4CjF2mXw8K51TQ5rBaY9GB28
AYEvbDK+6Etvg5OpeMMk1npzcblqiw6VIAWgCGTCakAY5sBoSYX4KF4mWz6I4R64
9BCa3wtzBKsxFZT0rg85uGQYQdX3F6xGmFdPkAoCc7nSFWKbuZWv5ftidrxWYBB2
FXnldg9BFjUblWgBH3PtVkhpaxvtaEORBlkppTpP0dm3Qh0bU3yOfEgxDHugxNSl
QwR8H9zXR4gkgwlaW+4cUALmumW/KnYHA88w94h+N2M7XxaXsCCPuRvmsOx0CR/1
sxSuJrvFX8v6docaS5MV4nCIxRfkxyjpSdCekOjLSopwzhzN2PMQBc/Qav1U05QB
9VnSQ4qkJNUg9xx8feHzf0wanKR5LzWhJB0hFAfb6hLpSca7flafGD54fnQVxQw3
G6PgUOBxfXp6j86HjygtKnNhMxuXI2j7MIw9z4eKRZ2TbMdkL5+lMYt1ZfqcLraB
8sbG+Uhkzx4cWFn56rJIHMR5HtLmitB1URMF7yI7k93bttuj0PgEde4Upw2TQ4hU
kQ/kbO3oA4r40WTWS8yYqI+jnNX71RkP59C3QGnw7pEXAmhcpQgVx8b0oU0GODrI
i7Aykv/G86TuaZznYfZCrEwdMur14UYLEvpuCrWAnOqIK+rGjEhxODFY26PU4caL
ebx7h5bZV/dHRkzmP4Shue0NS3uWdgwzT9S460zoGrdKrBq93/QDZsay628oWa10
m4JekeKTFGHP+n8uW20Ji2gI0aUwHMprhqeaL8xJiPuqzE11E0Jk/jWohZ1/9cfw
W06AWcS5Jk/ucZELi4epoW40IOpbN8fNj6bK0F4Rq9wM6DGEBMADDbwsRHz69I7z
JXByIvbMM8YvH7pCgcU0oFTCkkKt8xm77rOdj2sz8Y3liK6IgHCjXHyrDJNWxPs6
QrWcAm3sOBe6m/fjYsCm0CvYSwX2kN1yIhiay/SguTb4H6iMdtmU/dG5dTAkD/B+
NLjEgjpWnc3M0X9lQCtNxFrhhU+lufUb2WJA44W+1u8FHpt6cvx9jqE9mfLPTUUY
DS7Q3mpmufcyZ4G9GnhVyDqvXFo4OJaHLeBtQ1JhUEpkS+IeI5gcxLBAcnqe5Fvy
L/IQFwORAAgoUcZ0x+kO15ncl0LNZrFwz6C95OvNL+t4Yr/Ge0xXJHQzPR4Ev5o8
1FPOO9xGLnm5tTbrkQQifOjRxI3bnUY3N32o/xuPFIc+4+scH1n3MipfBoqWFrkK
SA3sKo9Y/o4YysrvbgAeFPxBLMr6ymAGNXOErs83NQsxKBn6AQXpFnTFqgUYqlX/
BCmWJnLC4+riqUOG/3mJM6I0pib4a0LYMXAtDmLIuqDeSS4OKUwjY8JcGbG0K7iH
eB0XXymcutKirsOKWugUOCvZ1it7Z/brA2jbfkFJYL8snFWvcDQLGWPQuDYCwL8g
iQ27nsqaJF/2fUoL4DAbBc8MkM9axM8oELG3+xKDJTmfVheb1cX0JkU0XewOn5oU
5TVWpUcM9IfIRGyt7HduXXuImepqdpN/d1Byh2fIiQ6/3pYW6sE7Bnxv/2cJb0F7
20X/DlTpKD4oz7B0XYejqL3g14RA6Sn1ebcJBQXP1tTOM6BKHN1CKv6Xdh+051ZF
kaUfcEy9YBB+mDtIQpddzb2Ok3V2GiwsPyjQG/DXPsFmAXXyHdpYjMY5YKivP00F
XW3YeiZMPQhEI6wDZa5B6Dgjvt6G1m/8qwQ2YESOLJ4mGhUeLiyh0lVa9NETEmEg
W+XYCdO9WgXsj5r/VaBmMz24SMgLAnzgGQhD1gzAIzk83HBbs7sBbtUHWNBLKVcb
sQ/QbmOb5NhPCS2eFiSlcyPik79DBSUHIIwq0RmGvPWmrDTE3H+V11m2E32jcCoM
Rbm6vKQoyoS0GSKQlfMjtGN9RPmGeKuhFY/Nh+DKEh9TX9CcV63zBhrzFjJU0fSA
HAc/GOKTVc+/hlBbVT1gR/+sOgfsDbT65nVWPsGJv9pixk84lSx05ng3IcS6ZVFt
2dIxgOqWC7RN9PmFgswbfq2uJ+PuGrDSHuiMIvVOI76XZkiXTWTk68MkFiczKtQy
NrgcTgNIilsMhVDeEDliDOnf9dOEE6Bi0cz0v3APov8RWSoXgkl2grhn2HXu1+W4
oEyjNlWmwMWTZOUJu/uXRxo3r0Ow/YNV48VHpvxGPrOrtr2Z2dSPpFVA8O1p8Y6S
HlfNy7tqKQLdk2nsP8wR3s1P8MYfkhdSfnlkBBuaJWfh5Ab4llxXakpTaogTvSkH
z4iYh0JCZBqJA00rDXjatiTqiieqVwdCbjm3k1UwTtufVgYzDROul3HeNu+Ecuec
SM1Rwmfk9pJktsf3u8jsoCOxVfwdYJ5jGsg6LeAhKGb/57zb1p7aU85HtJcGhTH9
gj/gzCLWCPZkDugcU0cGSsufA+1bZTAhB40r31SiP6ssPPRK4bjSZvCion5B60Mf
NdsFny2U4XU0GkrQxS2yM4ZSBo2t5NY2X7Wveb0H3hoIvjFmXHHqvr7BBSVCt4gB
8xCS1Y4VMXlB0AzZicIGHDI/3NIhLtJYOhMgs4XVJNIdNQufyyUE3luXAJ+odsnl
IDssKjpGUyu7ESRjI5uRr9QS3vKJ9ZPeDCP+FG3CtG9TbVuWZezf+wDAceimTXRf
xH66PbYWkUAas6m3p/7ZfKGU6B2peRT0F5VkZ3XBWZrwoOueDicu5WXE5O723DOW
R1377bu6pOUV5uKnE8wiVTtAx77Z5SzXyT/ja99P8ct7xk8v5P9s+yuDxsIOJWD3
PiZKtg55Olaws08MMl3xOW7Zn2SEfh9X7oop6+sQWVwfO6vBnDu6pCV+jbOxgPaM
5RAqPnQk3hqbqztcKAPRfI9JZ9zRLdE6FvAH9DsWuj+THyEyZVnCVQEOrN1hP/Es
h2fXgs6ZA99qVu+aadEDRyaCAgs2BEFQJBsBzMfFsbkr9F9IlH4iV/X2FozlwZ8g
n1qB9TvZnDB7XaDvVkvz2qQ52YBSSO/I/2cMEk/vFw8aDqrXrE88qg6JMjQ63VIT
eanqrsTzQDRqE03UI76pJcavv1QrFr6Ig8bjPmWKMCjQbhjFQQMSoq5uKARcVcj4
BpSiU0ToqpVb8CDIbeCRh/TsKxoMsz5NHy9VtcF3vpMQePHoj4V3ZcvQUgKRhlmZ
owznO3wh/JLiKPXTZ94hmGxPdwUt1ByiYrjRtPSzmBGRwUgCByox5T1OXM94uwMf
6p+sPB6cC3JnaqX5/+fDIXBZjgxDaO+F8t1YAwCpRqi6Z+5imI0txRP6czIAJRgn
n6r8yNEl7xgJ9pdhVA6euNQPjawJgxrE6uRqMjdaJiZPqvCvRB9RTTwKiReIYnc5
gE6LoeYyoYXCDtfyF+Koac17VRi3MMawCTzuzRZZbyAP0PusKlmdzYf0poX1nUHH
OfprLyNpj89QMULwKFn5Ay95hxH7e9qSqGAcLPLoMYKjBZMIBlaNqWWhQL2CgobU
B7kFsz9EUyclLsCRz8f0NYEbT54EZqKHwW2icDhH91k5om9j0I/hF3qgcOg7tlby
vNT13ioF97gmvoc2mikDHL33dvUwca0ICLNz0ElqUC29feQQR9JjjO6NXNSQ9WXM
eOxz7bpfOuGxDwkefPTfaRhnDeafjoP6TtQWrEzfN7v+CRvyVtv+JZB3dt7QCeM+
Xm0q1pDTcmpEVthyDlCio+GKbJO9vjBbdHJgT8w+VSy9VFP0sGTXuaa8gpKpoRBC
eEFwS4isuBQayv7l5a2izEb8ZgYTRShqykT6+juVG6a2NWEP5Oyq8a1qmtkv25gI
f7oEe+pmcsYn3jScW8uAEl8pQep9kE+gd/R1baJUvCKYV3Y8to7VwxnnhvsysQGF
jZECGXwWg2nkv+60+mXHGEzoI2t5I2IoAQl07ImjoDvuYgrlhOp9JCa2FJLHPGG+
/pIN7i9ksV0gmIjROjmVwhVewm4lwObnIJD6FPyfEpRCXiq3ZQuyvW6mBtiLgeS7
gd9xgnPoiMT9Df7MDUGrJrthfvQaK8pcBRIl3Ll43EqfvezpzIcQl7z5xkXpXTEi
ZMQoxnBnVbJABTRMfLzCt9yTEQa1qDkxrHxGTkEYZRru6uKg11Qd0kWYm+ElcKrq
6delW4ACj47x7/tmxwpNsj/yRIvh/V6RUe0jcRfNaAtJTggMaY0v9xDyRKMiDCPv
SZnzy+SvdEC6QhQPIwBRO5jERqT0t0NRWgRF5LM8Ybj/LZhrJZEtMRDXyjs14hod
v34TX2FynfGlQhU6+ZvfDNBa7ZjrL4UHrMu/wcAXFDHheUqQeW2Slln7TKkk1Uu/
CSM76uWmikvWFewNpc5bfUjLHM7Ci2kUsg4KbGWIbNQ6BsWk+/i0aRbe74cEWvk7
ze2po3avbCzrOuC6oLeVDjs8hD3wYq9bGL/yjs9MPI+BZhP/KRk8bRCFELqavVIR
b08yYJ0J8ExPyJ5GBKvmi5QvQ3+3TrB5y3qBoPpPLI+knUVyNojC5LUdegZnFphU
P3J2jZkCUAbFOWhR8kOooI+4DwKQ8io374dwYn8vIDT8DPIp2qxojWdZazAzFHBu
Fcu4kx9IXkLCbi2+wIZGCicrNHSBwVIEO1mYaw5yYcm6nQjSarAws6835pCmhqJA
ZiMaR4fowT/75WTOwxpp8hUqGzj00v4LCviaFElTCW2RuC8OBgoSOCbGjBwh+8gN
hfr1+RXBza+dtV68HieC2vu+/DVyIPUIuXZOSQZbLfoBBlj0tevWsXdSiJhUD1HH
lOJXKoXbRssjGq5OJqib/XAznoshvjayfW+hfBOoOZI/Xnn9NVbNz6QaMjcTZNhU
e0nitCYQrnbmVM9bacrZUXMuppVULGw9Bk5NpTiNopH5VRjFvxsilgxSY50A9y7G
DYMAjdb4lenfcI9pM+SO4XN16QCIfnU0jXsuijTdcsTAmN8/Ke3vDWxbNsYBvNWB
FDtNm1uwgZz9bAz4ATi16K8FwT+fpe8T5GZMZ1XMuX26im3AIBoBQ6+FVsZ43uyc
DHnGds+TSz8z2JXXsheh+g//nQknLHmA6uv/etfsXSbEiAP1V7mTi4xqWD10L97h
yUPaquomq5n7ub4ecF3qsnIKSTmRZwS+vm0JoGWv0H7wdPkHuY/I6paYaZOvTbuW
E8YV9MDHJoYMeyctBWTtv0awwIBrTIlE9p6vcTuYo4UBYWc7cVgTqeU8kDIF0y8P
g2XoqeDBm2O+V0sn71CmAXS+hovyKQ8pn5ZkGH600jk9e/V+NsBxtaPzPS+YSZWk
FwHaDVOQXQuUWyk25hNoh0KPv+uwq80Y0gakPnBens1xodn3NiD6fLgOofFGe8yt
OTFflVxzoT2O7vZ8nyO+LuLljWeoSAjf9RNNMiRTdL/4nzfVODh8ByHGhJszpwgp
1TXSpguyfvGf5g6AR+p0yy8sJvqs0i8qGS1jPPgV53YjV2tUNOdxe8qTY8j2WT/d
mDBjPP9RcczhYOUHc925uDBSMPF7KXCGdEvjoh82Pc7Hzv5PZ1yaPGPyjE0j8GhK
O38kbc6FlMjRZL46YMMlExzxWHVQEVVx7jtTpNfRKjwI9h6frRv3+oSs9Qh1s3Wg
NdvtM6yHVvfo9Tc4LHuHoNNn8AYIwrxRJh7c2fqB+Cb8SRUti2ZNHIrrtM23fBDH
tx4y1uZ2P1szsQ1oE52fQuF6q4w3vbvj7V/6mFNvf1hwGN7kTMoEy9gUtgbsgGot
PL7ZCy8lxfh62znSEIiPAxUUmbk7DuAmiYK8VEc1bx9B2V1QUc0wLzkX8stYh2wZ
mRleBqPg/wMclnz3+4BOsLg61JBEbrzmU+5sJJamz7/JEeClV7viw6QtxEuSKmuN
qeVm8kQ3dre3UpnsUFgzQne+tneX2bBYfNKaeEYeM9jLFWkNhpqRIed12/5SfvJm
G+qngNyTyattJRYBFssf6Twaj/sKza9a0FcKs2bQZvxIEciCyPCSqhbZwmwELAsr
wKtwWvvD3HLJlXuMYb9oXiwDux/9OpSRmOTgvQmSaq3xenWDfrIPi0lTv0ExdO2E
A2vUwJYUwKyWEt96VpWMGRvnsSRxEih/c2bB7qdI2vf1o5Q3gEcpqEbPPL6E6WE+
/aNpLNIsquG1ZnSKVCV0AC8r5GG+RCtPlfkZGZyed3slW9en4Sv/WlqiSpjna6g0
uK2Ry3Bc5o8HL+lfvrTmHhCqZ2A/jadRrqxs1+knpRRABhELm6LKoF4VG6s0tJLS
J8fseKFT4fQvQH2YgsAoM7Drkqaq9rSJWzupNCQmztJILdovQHo9ZEtqFnlnlp5L
WaXG0YyJaC1s1icBswJz+J0MF26Cb09zp32IgfQ4qNhKQuM/CFsRcQxWZ2neFHVd
aND5BpAZdPUMUOyS9quEYXyxQGekXj48omElGxq7L6RHt49DW03bfxtwuIM9PrFq
AGPfqD3v05GRdZDVx5hEORoOHORx5QnYpI1zH5+lsfeAC3ngrDV5czmqrdDE54Lx
nTozEWOTxlyGXarG3AyGukM3n8+UWEjjiQXGolWP3ZL3VV89iRUjq/AOqfhOcVoO
tk53rgBR8z7iuiBeeMaTd1vxF5n6tNJMHSFjd4Uk4+jIDN11sOQiPTJxHv6In8UR
BPOswTYWv2v94w6/1GksogZM4bfwsW1+pXl45yofAE7yko5gFr2O9lX2p6ZVrPtm
UrbQoFpmY2EnHngxlJ0QujMLXfXXZdyb2DeVNetNAUxKLl46T4A2TpExkpv/1PP0
4SeqGCH6w5EU59vzraq6GoIQx2BT/N5jAtEMDHjc9ceAI6fw1vpt/1GxBrd5RI1N
F2Y/BWS3THEZJoJzCqz+if+IkYuiFVMmWgIS6hdvjnT+0plBUQOgt55vZkXh6AT3
pwjIljSYp3D6kuo3UNf+MoRqGMV3kvVCn7ads1n8UJSynaL4PQYIP9WhEzDLmMLt
TmXMOwC6SKX7U5y4SjfPZhCPkoedKimwAAKoc88agJr7nnR6FLu5jOE/20YD4vye
JF/gkmvx/jWbE2ZNf6jpvtpnxIy1XWVcZwNmTq8I8djL+WywsnbOoNcAR9eFCUgi
WMUcMUi2LAaD1VQCoKMvP/G5IAlMh3r95wD/0ZRsdF03T3Q/FEpLaRLi+WWQ6j2U
QoGkO0ISk/CvHVIlhrRjZWbj9mF8ukTKtfMXbDO6FehrmEFfOAIbELUE9+GzOJKH
Z9WiYfMVN8MKHGjvsIloNM/jxjH/yfk4UtDu8Lui2EaQbPrUnDHbB8y7s4oqNZ9y
RzvEnFqBMqaMEWyaQhixK2FDbEf9taKllfK8QGwPAH5iHekTjaBZE/IOrwkljw0r
hX1r3bMN9mndI4QrwN+klm6x7chlg6BQPTAGBlYwCuph0Vu8oXwTQ7bisR5o2D5z
bnn6j48i94XoZ9r6hWHpsghO4XjuLSAd2qoOFPDf4YFGN1RZkRbSl0r5M3mc4ySl
jyXG4a7a+9vAT3a4cBz8bRcQg9zaysXexy5s3vFE4Tj1oGMtvS4PCMbzAmbCJ4HS
00iBbRCINPMBgyps1G6SF/Rhi2yTOvO6iAwZ4opxOeliqDQLN+Ct5zIwzIt/Ppoa
TqyhDNwjP3zXSf4NPBB9k2q6uzRsJtYxAYiewjAWWFgxG07fPaTpXxhzWyW7vFjh
N9zOHeS+SOH71tPDmYgowQFp0O7qnkq8p9adLOV90d84m9kftJu8eGydKl/FxK/5
bWeRuOZ8if9pL87rXll3bRGRVE+sUPUnUJvLrQYlX4KRDgXkC5n2U0QYtm+Beqyi
VH122UcxiK4EmsNsKGIGuXgkB2TkBmym//ighhQJltvl9qzAN1Alhmv2hyTjE7Nx
+aHn5n5g7avaBiA8D9BHApPSHUY4SRqdwGuNp0hEhQWfCGeBcOz92HfqGD8coSz7
1Uq4H/wg/WJviEoN2FsauDTTCBkZNBinmPgkLeVoh7ayBhEH8o0Gs8K7/vVcaTpr
zVN6sSK0OXTryyduYSU2b6AmX7US9gl9hRgvCFDfZYgXolrC2dDIq8mH1EuXdmiy
2QaiRApEqi5Z/Ik5h5kVnQyLbQAzDUa+HK/Sku4FrgRVpZVXFddnp1JD+g/Dg2e5
cXqgLnZ55ziqF36bJMpwI6jdq1it7rl+4xQMSq3qVTl9/rIn7RX+T9oKCvX183dn
nx1Slm6ZdRLu5b/lObvsLyNAvcU72aKAWFC6C1ywPLfqvu5VKExn7oe382vjPHp5
jF4sdcKhNyqKoOXVGuURdGMMKQgMTmvSQ5h5zqJHIRR646ox3t5cYz3TAZIFk4d/
RXLI+JQU5p8y+0fS5dGN3zVUQsWQKMkHPGJFfcx/Xn+B3WkQiIEPkJ/IYSCQNe1W
UCN+Fibh5aHj3T9vMMyD1CD7BC8GvUshHsHZSUd24sq7cY8VM3h93faI34ibFgUw
Rj5644/xAA/XjedW7OU7x9mI6jEy9yFjy5vGvGZ+5feBJpVKW2EAbkw/GR0RB0Ub
9DVX3nJDKSV+CGQahQm8WJek6EfnWEbHlPbTqBPFxywhOVpg9TNOnNLkj8lDorpB
j6jNfzpaGahdRZKbPTvIKN3YOww9M2eGdkFvlXydFmapdvQJUPxvVxry7W40ffZR
LnqZMv7qJFD7sO2KDrM1Jj2caJfGqZVW03JhXeZ72sIbfdayz6KXaGbfdIXfLsc6
y5ySmsqZuGH1InfEjirpHgwAtTC8vbhj5bgxCZ8Nmps5nfIRFpvrn1DkF2zuN25J
2gxZCYXcwHqilkPrV0C2LHd0x3pwn3stbpveX+FNJw5UNRgAhbxbQMq3YIpVUWqI
8MsogS2QdXeSWd7MkRhHJi8X6pR2e3Lh0jqdHPbtUdOLxaofVlrTHqInAz0yK2o6
YoZwHTQvFkdWe36f3XH29Mh3F/ZhOJHn2bjHjnxDxYk/e3i+J9HCIIwvm1YRokOS
Pf11LatX4uxuwhYq+dvG6VTVdA1Gs9ZEOBpO9fFQsw1JBSmdl6QgVe1tlSpRvjQ6
OkvcY6CBNn4juNsWkQagfdAf+Af+CuewphLEmloA7nZl8lzHnaNoNtn5/yG72C8I
/9nYE8pTAl0NKfxzr7b87d1WLEIwHux4sAPy6BlDZbaNRRHH+TuZ3NQQQBoNdubV
Y6n0+1+QEzF+ngtxcYmhG4RqzMurJXACjEhNjRQaGl9FE91Y3bRDTF/BX3OI2TXu
QiMYYqqPyX6vYiKmI5mbW438vPOA4XL+sS8BU9PEVzl7Jrx3eYe3JbB1F/5Gc4sJ
nwpfKwtITV7daD+SqNeFbgG4bUNYCvpXwopPx9u/3ZWZpuZDpobAOSDs7li758r6
YORIwHXbzjKQTqkxU1HJ0yaIHx6nnXyGJnM/eQrZYbRtg5/r5M+HapcAk+R7clXf
oR45BJGSyrXkpF4PX7WfZP623SPp9kAVNpPx5uzLbeH4tMK22GfrgiDq4PU0gZ61
wDEN/NlolyJBm7QTdukYjrO3WO+zRJPglZZZ78Uwn31gjMIAjG5musuw+XXaxvRc
qW3OySqflgJOUbbLOGXWV+tk7uBh7B6ROc/vsID795XiSYmBLsIy58oqdLQkNxRl
TrGpp4qmxvHsGz0Iix5jIwWVcfk4xlI0UYYV+VqrAUQPPmAJI5ntPUXMVUAnMihY
fYZ9r6BwxRCLJv7xo4bQoQlIB4Cq+JiATmmCriHZRyeHwD69eQB2KZzo/uiF3rsm
an+duUuUhps4RiNUN5+YeeZiaKB9TAl3S6/PL4w0DTr3aJBV9zhatiAXqq+tSrju
L36PqxNAcqo+vJ3JNPyj4BaH4q7ciImll86q87iA8/qoys5hLsbgGa5bsxLDSRyr
cuIQId9YPojMuv0edMXkA75GpHrACjyFysoO0zKajHOMcshWYM/2+B2PazRhMvMi
+hW5a5gN8LdBUNf5LFkmRhXjpnWSHqL63hzLBsrv802/wle8pewUG5heA2Csw2zy
fePMXaqJxrtZrN7pWYOKj1aiWHLY/C8zKRVRYqVtJ13GmGY8YiUfmD4UmWCfxhD9
bVQnvN4u3ks3YBj+8QiXb+Jl+2zRjLsH8uUu9ORvZkfgcM7s6w7OU1qYPJk7BliK
8Esf1x3hrlShbvWuwDEw2YG0X1GO5rsC76wx8ZiCxUBXHLhn9osfLOXvcXfODnON
Ejy8Ls/orHNGn89m4mHVpRw0FtcAgQwTwr98MYw+AjBor2HUX9q+KHY4Lov5PAwU
/5u1zKd+ueWrPevVFZ/NeK59s0lAtw1JsPDpjnkEJEDtbQZAjWN28pZSnQFiwBNK
yyRxJgRBjrp8TJLol2wfR0x1zd2wTn0f2iU3guLimcZnNLFWIBsYJMYML0wL+Zjw
a9tMj1glX3HegABRvabjxqyrX/I8Cv9mGU3oVHHhCmpzblISqkOWui/M1g8c9AUK
TpCo6ZPF4OuzV9BZ6sQ4s8nsPcUuFACua+CrlgmxCO2Jdf7YiD1VQhejwOa6jOiO
AuYdDsB/EpjP44kM98aXHO5mVCjGyarhy0MKf56CfjYUWdanlHqCpJ2gL1wElcoC
5tl3WO44Ndz8VJ+WjA4Eg8WWnrZAdo+I4KAeTu4qUCW3hbq317lbNWnJ8c/yyFSO
I7zFiN4RLEMY77Ao065PmX06Prs0crJQlD7APrtiZgeYzJtIQzVHw5tp7tC1jN6C
5tNH/6S5aYL+x+lRfhTXW9cNy2aXSqjW6FyRW4jWYWq0S98pSYeX+ko1P8xPgRYJ
Pq2LMs5dmcTmfPcXgTXaKTr3J3TcYMX3cIy63e87ftjz763qxB0OcPtNZzeaw0oF
6NqR8XIdl4YQDzuHYhTrNvvcfawTxklF78Lntw4dptuAUl+nQDzzFb1IGeTQYT6q
viQrPvitP3F+MskwT0IfbDazCvsyLbXGkzDNn3NPR3DjgtzrnnTh/FHC4+y/Q6y+
KH0g9V5viKRHo3nEEZcQinX+oh7tcnekNX76sVu7WvEmIoojct7JEAkVcO3k2guT
hmo6cH2Olf5bwKozzf8MeZ3SesTc0AYRMroW+9uZXV51aMaw/vWEOKhHxzjHeWMF
sZcNW8j5r0blMmiy3vfeqDeGsJ5e8emD5w918Nst/lQx113LDj6QmMReBfU669FS
rXGRc0z5WdWqt6kaQ9mlqjIz5ux+kyH/LIlb8Jf5KdJPbDfoMldurzU3SUw8AZwg
57XC6ifWB13+zJzBIE8HIlYZdw2ZlrHJ5tm62qLkaWX4QDJPHptN3gfKcn4EX3/K
5y7fW9hVjLByrp8GNaG/Xe5qNgYZEqMHY7Q6gKFdydZumbuIsbnLg4sl2aSF+yS0
SJYwxq+0gkGwMCUx1lM1PWAGIJ+6qUrtgNVyRaKwe5GS/bqQufiE2Do6bdZYMa7U
MsquxpWOUoeQsCEkM3vig622+EYLM2YWVSRrmImO/4rCvhiEMjXC2pGQPOZS/TC4
Wt81GD+p34lUHa6rxgIKhW2R0JzI12NJoX+Nm3A3/a3hQxhssRdbcKg5tXMj6ksq
AnPA9cyug7rFfRn4B9A9E4N6jtY/eeHADWyzpDJEGZSJ0TnVKhLjCfOVtKb822oS
ddQE/TKqcCnZNI2Z99D7DeXNx60eTummcUeh9GOqqlZdStaBFybtGP8b4kfacaCI
16LYPMOZeaV/tq9jFMiyXClkRk1U5uGVS8djMKSoaJ3WwajJw5h+oaNqgGkef0FZ
BO/TwNXuAh78w0BqalNRFIWczLpfI9VUTWUAzNIfKd/lJu6q16O1JbnMIxjMN76S
Eqkj4BOs6l18eVlCu/up/Ojp4pjSwVfLJeV5g6Qtkj1EmsLTz0X8k7feOOCatlxL
72Ph79iH5spByKZmhCdaLSNGCghG65H7vOhgbIDRKaPtb42J6Kna9orF6uPZfgFi
Snoh5sDTGwupdYZIO/grx3bwOxj5ZMsaRK8J9QSw6L1FQambv41RVhun+C/ouOP9
O7mBw8rMK9kBg9271jbaAt9BLxAX3WvkVrdR7kN30BN8b6VrPfoNDYnmxORpNdQG
Uw1xdHMfTWpU7S3RuesKtwaNPQfngQBnpYDyI8vWorJVAOrryHZxAUa6a1no8n+1
JDaGopdT0hkmOuolyudC1Xe5GYMB/t30LF4I1Vjlo/CekMqGxOjshMapL5mRygl8
D4vq2dwalPUwLB5q3+MPdhudA5QLXvpaoq3UM1FGhshAdT85Q0i3zQL7YyohJK9y
ReoqdYKHS3p8tyfMlK0X3G6ogGw9vObrQBitDgjPoPf05EM8ainFPbkIGYdtDzrB
/zc8ynnhK8S+STSix/kH9+WbBcAsUsEu/kdhMmczhXlf47IlWNrDdtSHorTovTq6
R1NPTrCZhMsnSABovXrA1siAhLGefxUx9y2G4xZaq2/hgStqEFPFtcMYHthi5NBT
jIzGU/vECD4jn9E5c7Wfuo7Xo9zkSeXkSDfxGBp4Kg93glQVyG98ArRufiKHEped
3l9YINaSGoXgGakJXBQ0adPk5BveHR7DApdgGQbb1thQwCEsbl/2U7vz6OEhM5ol
PEb3AKWxofcSD2BJVwjkwURwGVyHTtXCnjgnNJiw+jlhF9U5eO+zbIY8lq2jV1mL
k+MLc/6hTfkiT/GuwQiNCzIwgjnt4RukzWoym16o5sGBXaC9XwEfDiDQjj94+h9U
vlEd2LzqThJq9kxR3tLNv3UDwsI3hjFXltKdAmZr5hK5CoAsSz7qPZsSfRI4b4DH
T6P/YDayL5HV4tmdTlISGrtNEq2zKpJn6UGfrD/s5XskDBm1YRiwa2EITI4TZr0u
yx1VNvvRJD5teLiNoJNWFpl7m695559AD6yWgeyqxjBAsqnDrSnPdj6p6gmXGDE6
9JVI9VQaQm4/EpaAzyUdx5gEOy7Mx7Pjd9N09NYXkE+FF9SfRiNI3fedUgvk/U2A
1NVXoMua5AdJt664lxuLB3/WJDsiOOqs9Fl2F94Qp2/QGTITIyEqFGxKUjvJjNpj
L+sujDAoaZl6OEacBPb1oMHX324CzCOvOva+QgpRz0dcXR5tGnVMYXzpMeHgDd7l
VwMLYSyT0CSXzUA1NyG6YjUsQMR7vNzTKZ5kSN3/E8L8gV8JJ/Iw/Agj5EecUZxe
h8l+PJmraLb/sgoLVtUe1iFVKydFv+whEgL1mvugBRle92Z17rz8ymii8NPO42Mr
SR/G7XHAlDJyvI80T7BRry8wgJJJQswlUIUz7d4mIq+WI3Cb5MwxIqjwcMaTeumF
wCBv8+N/qDdBlCKsvo/w/fgxUCWlw305f90GyOCPg3ZsodL1nvXBGhjZWPDBFdDg
VkzRECCoy0UCuBmqENfhF86tgFCrVi4KQgh4XfrAdgKKnc9gN3AJhsAfdoPPwq4t
hWkwqDw0636Psw9dvGVVvLN4dwKai4zmGADuV2mj1z/R0hE0VlOUl5ceEzBDHsWg
3qjszfRU+rol6E8Q3XmGYAXBsCUm7TzVSaI8y0z/36iS8slxtBaHJJBDTWS/hHXv
mZq4+h3+Mt2eIT6+Fj3LDjt0ySv6XaVOVI6xrcHGWklBdcwkNl9naSOAX7Z8fO+u
krLwxUbQhG3SC0x23A+hbWCRQ8P9cv3Hr536f+44nUAGyhvwe/6ZshsjQOBpFGnS
jr7NMcccOlWNANci0oP1AL788LSEZ0QYopZxa3s1p6hFSZW3tyQ0xz1nqL12djaG
joTGGp2HiZz2IKr6AEkFdH9suZNzyr3dcg3tmVHUaR+MsPPSdsBGeTjIOblKJ6QD
p6HeNYcFm5UqE+MVBtYc6sUEp2pTfzqOI4NYZhOdcU+lXz9jE6YdLQ//L4oRxvHO
FtE8AbLH4VajYA9wUrixoA7RZFUYAHxAtPz1bhtgI26AH9y03mj18CDUGk1posDQ
UeY25HyW64c0LfDHS8NN/jaqMVHTHNWCvnoCgYgNB8euOGJAqBE1QIvjSRNIrBDY
Bfymf2YzA2qQ+w5QKaKkxAV4p4MtbqqwD8kW1soxMIKLYbXLlo9DUlXMJD54Ng/H
TTXYj8Mi2Rf5gYhb+kh/0TaetOStEuP61xnKUtx2HFFTSnsoBhWNQbC7+jqFZkQg
EwrQABLfmwGO5ijtM4rvOPNbumj84BG+QW2NfhAR2Vncjd+1FcGytBI2ojQ30AO9
ZcYf+Nl2oF49/o8KNATl7tz2zbgwXL622vEyG3Hsw9iwI/qSBHs5jxSW3Q77+b0A
y0Cn3Mc0kwWE7khnSKelAe52i4ZjIoBRtLLEIihTrxs+LUcRISDGdWpAxXksjRnW
HfYQYvk/gpPVEAE0Xg/n+wyCA8MjmH6gPm19rCi3XcGDbDkNU09xb9N4qre2Vgyg
dUcYOL9EYAv14cb6lCevgXOUpD/yndpbmB2Jq7QnPMjzzZ+KVi2b+pgOzY/Ng4ql
qWyBPZ8LXwb81LZxCztIwZYJOj9MEsLrggLIj7TonBav8XsNHW6fU+rWZ54AD4Ly
PBkEwe3P+c+gS1VQxb2nM8kqJWE5VZeB4y/chrpZaQbs+ef+Ie3mxfKSakw+CM3r
+ZxPU8V68x/cHI9lqZIC/bvtkbzQ/ld3AoUxcbISR6QVkm8ge+FvaOCwASXbiyQg
hZMapblxsWa90cxHyCrmFVM5qbAxNragW2aBEebEIGPk3b3JNUnS9Qfd43NVfX4j
e80cVocct7v+ZhIjchEuD00I8InnwDDIL7VvC+gUvL0A0GRi6Ku0nP9zrLqCsNDG
LsmQULm6nW+FSIWK2D16Q2i6tzCZXtthe3Jyi2efMxTeU8XYtjPCxGhe2I97sawr
rjdAe+BYL2ffArp8FD4L3YMs9rfcEKYj1UrpPEE5gycrVwu1ASclnkC3UmHSlG/R
g/4K2noErwEyBm5RLlkxnb+IYz2clKro2k4zVVVChNtbbeLjQuEXjYu12Xe5xfhg
51bAxnuRezrD2xy9YI4m3axDQFizXpcsr07yzuxyPczvrQTNRz85MVmjTU6JjY0v
OQJPkyNCKskuNeOFNcJrgMsfZC8YKgR/qR9QaCaFkABXXDHR1mZ9CAn5Fly6RcUb
bB/x4gEvFazv9WttNIdtaQKPSRkyim38Awktv9w236Mm3aTk/pXVe3iUKa1eVBcC
ZWQTl5Kg53qUnTtGP8vhr2Z/ChHFDTxZiq4dUclLxTIHwluCsipYDXfFX9/lYO5v
K5LIHLNzm1kovjXfh/ak2EX5ssifwH1FN+K18H8j9SpFuACFbe5CCVGe3D83R1Tm
Zf1P0h1rxA6JM3CHiaiLLko4hPu36s57JpqWz+yhkRGS0dGzylx/7enGyiANxXxZ
sQkAp9CdsFV5c+Od7ESyS1D2yi6LkNVxtd8YyuXwsRoPf0dP54XrgV3AYzCOgYe1
l0V58BKVDIlwcpecLtFvA9fystUevo5enHrMEAITYpfKdEt9/EdopgNjnUe3pkK6
FgtycXjjd+aRD+86Zx470kminEvoB0zXxjIb9p2rwzS+2yV8bNhlXCnKy7zKy723
9AYfN9oCEEwph096JuD+gTNpVAtDQ5sEpaJNv+c9qiHqidJjcSGIwUllIvjw51tn
+lef5ZEf3C2c4lM8pduBs8tpYaAGReYun/xrzm6+TCI9OthGdZGIcnF13yc9Wya0
29xanCSFxULOogIvGlpIWFzrz4Mxchc92Xm366hsfXhFZ+TCc5PxdpAEIuxtJ6wN
CDH/Wkev+x4WFyGuOixYLI+rxoWoZ7KXaqLAD5jw7kKL5L9fPS8tH3N1b5LMenTu
I8BYBXj4ZtFw3TPoNxJ3IMwGqxMlB7zCFdIPpl9lclcPggqSCw0POol43ZOmHkE0
oRu+7b+5d9EdMJtaWzZEdNPvkvOgeDHw+VTNbee4OnKobktnaOcsAga23sAjfPcA
wF10V1vpWO6Vg2ccSi3C4mgJRbrhDXpDht3PFg/qnbfTuIe8kLuFAeu4KS4zDMKP
WNSTrXLv9zFn5rlVyam+VjCfmKHb7YKnbR75lzNp8vYIWi8tn+KERffERBkBlkDW
aDBwJDSvzyL4+UqlAotkXxhNXiFiz5EkZVRuQ6yGcumAFMZjk+E8/m5DmCU+Vgb2
HbOzPbKzSbqSHXChROAev7sr4v9ZVYTW101xxU4W7twnvkfTmBI1JZiqKaz8TdX2
jWJHZy6LbZs0L4xendXPy9p0AANv56l4AZLyAJfPVyy6srLGVKhHlL9WdttMDZLi
IxRa+pA2noiAMO2l/4La3N1CriRi6/lEaar+dVcaM5NLOi7pHn8Bnt1eQHc/KUoN
4ViVQJ+eyKVwaAy7qDyu3cupwTQRfztYpLtP996ceXSptp1rNlGVYR6PwozhFWEZ
+O03ikZggrmw6r8mFNNiGkwTnPTwo1qGKk3jaMnN55zOC8TlPyJzE/kBOSeG5rCd
8kRvS3qCojmd5ad+Hs6i8U/1StUoVcf0MARr0c3tHnuNF4HBbFJ9ESPuqSqZ19do
12QHoOAVfgz0cd6YrhvC2nkEdNEN/d1I5fl4YO/BayA/+uqdz2b3IknDyqRnwiCD
2LQ8AkVkK1Hmb75RoFeID8FS7P3jNk8/Vrqf/p2g0rQDkfRJZZC1MhmfPbVMtqQj
atz9Da6Xt08g/+JDV0hY//eq7eLzD0E3gAwxDK0eCmexnn0PI6PNUzMkbp48juWl
ckKhnuC1S6/4xvnYSO/Sm+9z4a7fO04aZRieoFtAtAv8ZbdEJWE+/kvWm74LDg+c
J4wmlzxDkvYS13jFvUVLxornpBHVgI1hM9/xEJxhMyCD2PB82rfHGW+a3uC7723y
qnz4eDPfdR58IuGDaLpjpknCThUsdhJKnFJEyNO1kvK/NDhirm9ZZYAxq8EE6Taa
Fb6CPVR8yWf58Pwl4x3mJ3+E5OO0qdR7xR74Nwo8EaiijBUZ+j/WDYh6tH8xJHdw
HZTlfTS6LS0kTDEhH7GZZ8y5xwVZzmAaEPlgCloAFbW8LV12TdbwV4dMnnkk/yIv
GYkz01ZQxpJgNKJYnvs8iuXH1qPD4DZVrTaNeyurS17SxgsYX7u5BOy/7TOg/870
fxC1Mp8ABOho3b+LB16Vs8qtrcqv5VaZugu0vt5dtwkRnEqRU1PPZCsJYLPT4+zf
7ePXQNotb61sk/jmvNOpLD+mg1IO44E+eMY/ricw0L9HXEhwJcoc5n6AmW1J1rFs
ilvrGZqXHi+ijtJfEIup9Q7UEAW3pQ7HuPvH0Y5HzWQ9NUUCr6FZyI8/f2CWomuA
7Nfs060HSpVV1qHXX1z2xGvz5nQoH72JS/wzcz/GjHwR4PWxo30RCVSRRLnI397m
En8Uk9kv/bx3mKXbWeosjAmVUaVxn8FLR2o1vjbFR/ViOXAmFOMFlOA8sxnj26sK
0tO3vGj0315VUKEkPJ6dvn04a2AkuBZrO/fPKDF0lBFse9YV5GL9ombkrF1cr8ej
S35yhINVfAt/OVJyBu84AkS5EwhL/6SvM6xo3EaCNKEXW1qnTCk31P+UR9TBeyx1
h5hr4qehSySAPFA3MVay+JGkCvWH5GZy58eeq6kBnhAfBodKMRZUF05wSZygv3Fa
Sve7P/vo4kiFrPKgZ2dJAfPpwk8ByEJ7r0PZzifI/3tJjNY5TH2Fprxs1N7kfxZK
nRY/toiMTFFQTFSH81NUovApBo4JJ3MTf86mFVoTNN7L0H4ItVMxOk24PX90p6pK
8N/jThAHaJ0rVT+Dpzmsckjkpaj3NFkWa5GXXYnHscQKOmGRddoMmq2oCgUBKst1
FpAJOkjwSGh4WWsi4P1NgP05cl9CFDnRcNYTBdGuLrXh+wl5f7l4dxncB+aFWBJj
Z8la3/q0hiqTrMGobwVEtlLme4dr4/NUoe9f95flO1K+AhLiQoXE6sk4CloveT9E
uz4FfWBTstbTIEOKY4EiWo8K6YYwMYzyxN4IaDpIuHkDqxrBvBzvB2bAmccagl3s
DdemPACpJTZGuSfjfxpRoIMup50rniud+PuuO+P5iRFkFZBweUwWxG52DTDGh9p9
Ee4M2BwIx9GormtkuSgwvXqSAPdhmvMGVwyh2bLxSdxbRSchSbKHvdEpBPiI0GZA
YnGFl0rjRCishbB+sKiPzlM8mQ7ZDZ7VnCSZ3vQo9nf1WryKC6nW1ljIqKdHi4R2
cAoqgo/+XeCmyAfNPuf9syRseDrIIzzrJxDPKQ9AIOzE9jjVuGg2Or9DLUqAFnek
kjO5M+Un9JhnF1GmJ+j6yvnJpRU115uEqj4rmp4ZEomZo3lWkb060KKeriu+rgl0
Nkii9cGi4wnxRli1EEGbiZ/g+/2sXM/ZFq9uSN8ODRIroz1hvkdHyNbATfceucBy
TaqBm1nVEvqZu5AZ1tEFswdcyK7O46yWhHq3YPciqT7BpZ6RnRChHvZl4H1CqrPn
GiSXB0ebchgmrjQpwUWNt79v1aMt6GTKqRc4vdNMDvOcgG1eoFebRqi0vsQ4rNGt
blETEpwQBp5s8bEAL1/4cnXuI6+t/RKqibZgHS+1v3ckqXOJRlhIfLLrBZQ+qPIR
pswxmD3Fc1I7eDQHHM+IhyRa1NaXQLNtjKTdNvQBJOY8HVkFyC0TUjzmrdPjRQSM
sRYc3rgKpOqrGSPMqB7vEDs3hdqLKaQ/JASAi2u2Igmj6SCvki5E1Dt8Vq2NGs4z
paJGi+lQKsYKSeiMkKR5xrIe3yJrPXNxeLOoUrhoRsxiK5hIAXCmyVl7i78+qxw8
B2p/Kyw4Jtd0tb3ErMfQDkqv+Yqp7+PZRlo7jRmjlFnTpQhpNvGVErWfKREPUVhx
yY7dIwNb5cIgvCrTsdi7UhMc4ByLW33ia/XQN08mjTd17v86gIWgGNyzef24QDRT
lXWojw2+9L9Ryhqoil5BCIg6wbEK0tT/DgzLZZ/w/0LGbTTOq5t9K56lzGS5xj5M
f26jGJ/Ww5oxIB4nP36Xh06M1s3m7edYlJUSpp/XIG50KZ2b68eGI4kRjCxcC+Xr
TP4LqGlwlCUw09qlG8HxJwNcUhUi7DdiMR2PAnZ4yW8teHrcczxIjoIqNz/jl8wv
Z8PNiqpIJy3qeGhZAWywidMgC/ZvNUE0FfoLCPnc+vbb8Dz2pspnavF2nDGIpGSy
NbjGtmL0ky4/F7H9QVM8oGDxzLIn10dowCpZ8MzUxVzVDb23PPf0QdlynoQsU7sZ
6dOUnH7uGHybQ84qt/dY94+iL6OcsEpZ7uKOtzjeVo6DSt4bIY7G7JWmEArZpz6R
xUFqg+MHOqazZLbanpUc6Q/X0RCt91b/g6Lt5vwe+jWIitmZsSZjaki6uOSL4hee
mhU6cOVo4MSy1I7blxNRxnzjiRAGwEpn+iP9hvuoAqdvgHd5OKN8WrJ6SbORn9tN
UM23vyZPzH1UdNO4+ElZR7fF8OS7YW5VcYqhPd5TAPFA/bJprtCgtt5JcP2TeMHP
FPq/BTGkNt9N3beA0r97vEYfAMp3cbkUdS0vE7yVBk94Ipr64wQFJXtKDutR+0lV
ZE89/SkB0P0179ZL5V4Ee7zhCBfXtEv1QVXzbQr3oL8Efd8ecDMyM/QhHrkjzOdE
Uv8YQMOzT2rhlBhVSD54tJIudGkwgNcPRbltH8P8sjb/NwofKAl6sGeGZF7K9U4x
vzjKVxIa5d7ajscxHfgirCa5PteaZbTbQT5ZEY0nfFZHQDXiYvn8i7Xl2I7/Dmtk
nZxfays4hXclTGUjNDJV8+isT4JKlzyhV4Cv7tLaNmlUwi0ggdtcPh5zVcJa6XE9
77UfpngqXHiHW3sOG/M6Vry/DojXsMhrHTtwKRn7VbOd9MABSdx067zktzn+3YDq
lcCV7BX9IENEnEYaV+ARhBbns3i3N2t2DJSO0I213X70aCgAVbqcrshDrVW0bQfy
LkFYbyKp8DcVJh4buzT3wf3sHagTGC4MkSsJUYq/sfmRBdDSvxlQL6bdZCcy46cT
Gr3TuVbLu/8tRGMKmIHiVxPndeLiFb/FMFuF7ffTSN6dD/1wUl7aeR5eJC+HRJb4
GOXQDkjdriev35UH6FOwRqetxx6sOTbxn2QrrbzZbOHZUDw+H4kuNOxuK7YucZ5u
37P3NXTtOaZBEYIG4PHalwgL/+t4OrQIyDW8XGNmZ3ni2XPpyZMT0IVOuxD7khkJ
F/aorCMX92qmqO8i6/jxGPzw7/B2Ma939Jx93zb7zwCq86c4t0es5WIuYXpvUAll
6McSFmGbUrd19FvG4KWTTgOqCcPHFV7u3Dcx7CpSVqVueGuHfGZnLF2WywnW7W9V
uNvJMYMHqL+VX7hOQRTJAFPii/oQxq602SKTXuC2oAlScLJ5rtrTM+wMIFvFt104
jINLy+MCr2H9U7XAGIhLfCmrSEVj7bSUS0KT1f/5/KY85fwjqiuhNHR+Cx/AJPBo
/7ZoHJVdyeVHhmRE43DhDHHXfoOQ3Siua+8eMzkIMS3hbtnnEyiGnoEE5d5dCLA7
k4IX0b5lN8SFTon8swJH14HRft5VWHYM4q66wezPzSVUNwGvT2JhvLzWer3dMUhE
8owMjrJSp4OtVr1OhVYNHxuQvXaO/fGw4MDMIBMlcr8oKuo3QDwFrvVxbdqJab8I
yIgCL12hINrhvBFpY+hIAfxKfbUB7e8cWZ+Sk3AFfn26Bd3EJSo00LnoPJxKLOBS
tQdNcqC9T+YqeDdrx26Uv1A7Fe/pWTr6zXOd6XoR2KS2VBLewARFTznMuT8w82yl
idqNv87Qc93w5ZtJ7Rx6LZ7/3JugL7JWEyKTo0x3AmzLK/OVvagUsGkpQC6hMv5Y
lajJYaIUj6JKvMB3+YdOxpgeEiXjAdbHqx2FfQEG2guu6Rlm8SpXxwiPsenPwi1j
qOPIY2lYKOOLFZIUjFNFY6cPTxwa4WEpHOWJ6+3o+7/8oJ53iJ8DCHackNuOuFi2
7qxDCqBLzxPbcm8QwuMntQcFeODv9Kg9AlHh7e/xwQ7XwD8WrkMWZV22SxEqMmfe
8I74LeE2DDVsbzvvBIlCov/c3OwPPwh0qVdHVwz+EWv4R1F2ONlYKCMEf3mQhKhk
0xtFQwrFfLR3BsnKDPmzwXSYdXj+sTPv6Tq082TvYUzYqoICwizGOPpW+YcaeCv5
6FNT6FBOM6yqpOc/8/tYVlJ/Xr0EyvLySNFLa0icsFM45cnrLp3f4QDcljan3Nu1
rN9xNhoBVfMtuayQKXGXGOu85GIwQmc6+V/4DV05hxf4IDWmGlGRvfX25/XMiqAu
5P9Fj7le9VnLEIjPzWn9mSVb+eJdi3gaWIS/PjL2ilUDmNyeLRrsi5UFC+ygaCeh
jj4+TPqwJODQQoN1M65GwWxJKlAOKEbGDkzAvXf7xg0qVv62mEiYqLsv5NOIPfa0
cEA45KeTxFKPBMBNZgQwzITZ3S/kMCaMnAWig1dlpynE2jixqVvLSMWwMxdTBVbU
m6et7yXFK6AA0XjDfbQiFs/C/Ubnik2BZqpqS54NNTO5cpEzchNSz7DMnkL/2MII
/lEJGku9QZb4wKrzuvaggaEpTxv5aSzl5WIau+qiGbWzV1RgnukPgwBXUX0N3SjD
0ilGD+orYgXaK5+3itctqgJkvIBcwG3O+TM1XsEf8NsC4NO+4B5rG0EtIG6Fl4re
q9QTg5GjlY9B0g1gAQtSJYoXns+7hwyC2m/gkmGIvihVBaZ+T2/LnUl3Y3vJbQNk
3kDaJc8dprdJcsGtn+XTcVqHNMCV2AvwEcfKjuEtCjSaO4AWAoVuhI6RG2BW9+fl
vJp0JyzaRkzM+egaB49wcN8x4OVQwgcwfJR4cQE7txN9k0ZFH9/9KAtKe5TvYV8R
GyRxp0wsfm2mi7fXznQ/3Yn+2mMy51yYZQ2lcpzOP/hkmMzclDqWIkrg30zeMt8v
tBlrFkrm/VFneHYzRBnpbTIWCnc7yrASW8LXP/MM7azOscrNiN3Z9hYSDmR3WL2F
Fgc9yNu2ImGOxvbV22+z6mAQ8wdERiMgvk+9KIiI4dIJj/UZxVi26JI2DAjn29kZ
9/HyGC2ju/TrnQW5/FDZoljGpTjHp4EW/vuslPY5+mC0iT67xfxGwMuiZChvHRVl
y7qtwxJ/lDrkqQtnkR2BYNVbAvdS78tYZptTwdZq+/hgBRxDZxRLoADN8V6wpJvk
Gw91ut8rvdjfoVGPts0vngRn0p1LmlxPOw2VCIBDnDseBXaCzpEBAcJTJy0cKK36
oV2/KhDDfO5MCvsXWLwVdg8n2m4C7TPdrEm/+0xloJOEHRh+lvP4XU0QQN4mKAB3
nISX1uj+bu+goPuFE+Pmj4OrOjesQ0Px/ra27jTpOYisHVl26M6FiLZ4h/TusErd
X2bXsUEoCnC4ekFMSrM7HJp3v7PVkX7j1dm4YH0Ic0TMUdh96IdGmtL6hxjjR7+3
fje5z/eWQhX3zvAKufsyN5ar6yDciGHAS7Tb97q8bzD5TvAZIQAdeDWJeMI11HCx
RxVxDSuSt/cFCl/4ortnDxIzmWCzTr0w9OkOt3TzCtpJvknySrZgtLV5Y0hryTm6
pWUuLdhMkbjVBqyiACNThHYv0BkLuj7LtZrSgjNpWnj39Cr6fXRbtpxisGurWrXv
uzSZnQ/U9s4vZId974mbsUClEE6NS55WF9gGGYiXzq2G/gDiJHEUsAV+wTZIQmdn
2xqg8wEozXe4VFE5bZbM4L9QwP5xSHb/hkFC1cU4+T54FW4TeAfBRY4QAy/WIgxr
+0Vb7W0I3gYcRboQQpLrFXDdfOIvlx6cIF0q/dmCNu5W05VWTuLSx9eTbbHzbnt3
8geNyonSrzFF/eai/KioA0d+Lu4VPxrX9D/8f5EhN+AIkox0+padiYZNlHyUj0KF
eAT3ojjtgwa4Os6tO90Hb2RW/P60qOYGbFiRC+Qk33XDjGGAoaCcbbgA5vTS7phF
DtMJ4ihQVR39/oXY59VJ3Big7VMB/eXvrUCeNiKrAj3DZ1Twul+hZwAFWORzvtxP
N2AetuO/c6Yvwgg+4wMReFW3dSHltlZ30OeO0nmNl9gn0R5ZRkdos2Fp92uE1yYK
c0hBvxYV1HP9NFwv/j0Oi6lVWd18ZvnMAwul8JLJtkBWhyIsLlM6nGcxVHfU5URB
N6tKeAl2xGGEXMdix23LlNwIzFTydjAbkpK2RAN2nZZeAv6ZLgoQQrrnKmM+cAnm
JxPY9X4CmIBsURn1FT8sVi19cLI2cnKOwOCNE/R8Dn1VZn5PJazYfwUn/qeEvbT7
kXwU/QBZidannuZ7tSA5HFeV84HDqUI3sS56svk5Vh7VDnnT7HROOPbRNmh8+SL1
mBKyobgpObIi8iDK+z1A9sbWNOVF58t7XnZzw0kRq1P95uNpSbEPRGV9HFNULfrC
BS4xAoQujoKyvpZT0wcPwvZycJ72LXILDYwXG6d8RGJL933PwTeapfRwoBMjyRN1
0FXmdJkXzzhuja2HAPqfFyN2/fqFxSyE2qe5HJfMN3fpERitxg5ZDQYlqaaCegI2
w8sbglf8nNcuVPfCcq9/WgE2S7OsU9QBqfk5uakDGR8CGL6IuVlQc4Sab9hCSOEO
L5G9iT0YZjlw1Chfu8iPlYRESPxYd15qvf9JYt5h7vPWq9BFd1OxoQCujs6sQ5mA
gFE4GiHXjE5MZUuAVFGiqLsSV6h5phyNz3Yy+ntuz1FTFe0rpCp0IZ3Jp8QwFFH8
/+sjJeRsPrVn9s6uy9BSeuea+cCVcf25QCz9t9HwF8AkVbIuRAx3BmSYkX9n5lEn
Wa3NgAK2ffw6BuLKREU8FzRzgzNXM7yWKWA5SpUmHeaBvhJzzLVnCSZOcgNa1gzl
PDxnOjIUEWsDJwwt3ZC2qqDiBH3b1CPLvFABYDZF8YXJ//SAK3xXaUO0xZCBthux
e2QWp1eC2TBLJqwr4XfEP5FzaslKSgCfnkHYzh13fUzT1vx8IGfSwjrFj08ysJ16
lVNdJ4L0H3w0oXDOSuXL4P1qflUu8PMGxCUzwYCG5b24zH39ul6csImLDGazBC0w
sMXJhHBf67gb24hqwCp3vw0T5V+ohf13vTmBV+9e7kvFfgCfLTf/IUPnMtmgzYQx
vmuVvy5nSG3raK+izK30kgNv7ow39tE0cFDQTBV7tYu1iIRw63duT2qkj/YDJULe
eyuiEaAK44+IhZL+KUoVUHRSvnkF9sCyMU9tNgL0bu6vJg35pal/XYJc0cJkWbgu
0k/4HESu4MfrjXMZkEGFdQnDDKZulQT/n71sdfTw0ZpraNhBxdrFWCyJ/OwKjyTA
09qnWSS8aLdOuQB7fC4UiFDCnJCWQ2b8GIzwMCD63WiB+hTWYrfT8MW8VXoxN7+I
f9ckmNsKqz1TYn6cJUgue1ycLoNYig50CxcCi68wOUbDym1psm1ZsmLj4tWZo26K
rmCRT40nveT4kPZmoNNlahbxhYnQGGVvO5sfSVT1uHma/5lIkbuW8rkgBfQxMslh
8MRMm+waskCFhsMji2PwswRqQARiCg+8aK45tZk6tSkZjPdF5zUczag3V47Rq7VU
XTFvbI5hC/jZGpeDe5ul21aOl7NSXUmfk3zjZHomL15ysvsLhDZSpikaOO0Y/k3Z
x1LVIFor+dbyzQqPHFyRfIk41aK0taZQzYv7lclL8RFto0xqxx6lLY+U4f7YptFd
zcZcdDl8fNkXZTpoL88+BimA97DOo5+TCdQAgyTAzhxsVqtv54IWDrtcBEtl/Uuo
4qpDqh/rsNWApuYa0f3PIT0ZzCQueUOpg9oD66/VBIF6w6E7SamYhwzCEpeDXV4C
RPFObbEE9Cr2VnttWlGxB0Sunk9GOGRncNbJUs4adNKXgsp95+hAjPpXWMJ9pfgC
72bEljWcBvmcScxGqQk1TH0u6gu0xG0Ggt3pUTCCur3eXBZTdw9RkxmtPCJ5njd3
pmqGVQIDTmRwiXrx6mIhPClOFk7sOYa36jcL0te+qESXPRzcX0zP8zjfx3ECnpUN
nwLAGbtmm+BzHNuJoC1PbvnP49/vSUW8f91ay4sW03jn9WzfNojaco/dAWJgaWed
mMh8dwa/MVD06K3TIIE+KQS0JaTxxqvXP/lKjXJJNu7Ladhx55MUTBCBoZghyAln
yoxVdyNDqNMe5I2tInc0/oeH/pT0Txl8i/mxigz/BmqL5XYO6v5eU6evYeWHmu0F
S531n+6Opd9ZFH5iT7MTAWD7az2wPyEcPYOVO5FypoIK/3K8RCYKy3t94yWpx8Jy
2X7uc7C0F9DwZiAaEdq0cGtToD7CPEEGKBQByOa54AnSjbxNVqi/0gEUMNKJHHjC
384QC3Vc75qNBnqv27/N4Zcrifn9Io6X/iwJZgGPG4qakdR2Ht+r/7k0ZjIZfAK8
G89pxopi74Q6oSs4LkYvEn0HDkBXzyfeeCwaZPwQqx0zFDxZL6N5877DC0EPgYCF
LY8Olgxt+2gFf56glUQ+cHySf3kVQbWt+yH7IxhGnBn0zLwHEIRvozP+nGv9xmdb
q6nh8cVhmfcqQb8+zKfzeMDdBfTFMDjsINWgLmETIpOghDOZwgMF0JPgbAvb83E+
Ylavj9KBKTGQfqVYGTqr44GNYHSpN/nVovbiTh0upzKtQTqqM0s7O1ZzEZPvEpr9
kc0diD/nV93B7LGhul9d0rlhX3JpsSomQ3+TM8J3Ap9RzE14rL3zNzZT1YIEafdS
00kk+sYh5merl1FisQtMVC15z0o4QVwNXlIaMH1/RVBq7O0ffKHBiK3TR2rVTxx0
Ly461G99jdCt3Wn8QonMjqIddUWwhTiV2G3KsVsbQ1XvHCSzlI8gzY7A9NfzfAQA
nnOmKsshkeo1wo++Jvx+E81hFhetGhSj5QPUv1fxZQEGhp843lx5Ak/uIW2Usxqt
p3+YtdJBARSmWAM304LL20syeHRGWOKB4hsODpNvleg=
`protect END_PROTECTED