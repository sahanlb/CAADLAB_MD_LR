-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sP+xl9X79Sqq1WXSHfpzNesb5A+5JXe8h6YvYO0ak9Wg2XXb7HfQkaSmlRumUWUI
YVyub84JT80/nvm+zDRxEIc5pnLkCG0WQTIC/Zgze2wghYjuU+tjTFsmIu6z7w2b
erqF537G/Yysm7Sr/YjWCu+4vhgL3RNLRqIEBSdxOCc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9280)
`protect data_block
p+dT1izJIcETboxFOp34UstOseVz152+Zq1txjh00VAJysYUM9AOHMJURTBI56oL
hiQkO2z240gBi1Qsw/+TUA4pVFr5HGGcTWYEXUfaCfE7hAQV3ftyTmvmw7O4rDwa
vNCgg69lAK0qzuGuMC4MT/aLwUVluSmJtOyGC1pCI28x8FwuTSLvN2A/RMHd9/wf
RESnIq2xJw97Anc+A/Q4rsrzYKkUPEBMBAMiUMh6k2HQH1GmbeqxZv+lrD5EwmFb
FXQI1wpz9YgJx3VHrrGMUbqpgMqtuI/njnvO9+qFRhaVEUE6mWWTEcnyXB4cjROg
XdcBQuJYoUR9EFc0V7ygpGghb9O3e84yt5BrjHfBjD8Eyc5aGYPYiKylTOzCe5fF
uSahhu58NIaCnftKyDvsxMeGKD41jBIXV5GtJXvcubU9/Q/rmNiJPNDdNxSL/mPM
DsY+NwFn3YD9S/D24fkzuDwT0L3GOyoaW+rLbt+RE2Ke8/z2I8ZSWRgrkSCW5gk6
4KfrL0/e0RxRFPWoxcL4SKi/6FlOpgBAEfh7zkZ6Nq8iu+FpFpNY4jQ1FSQNmbPW
uak01LGZ2y77/wEzm8FdCCN8GBJ79P0/3jsPtb8ISpZ8kJEoh49x1H4QLMg3Kx/Z
ZBXzgBa7/hbDH29AHtr/2Qt7q0PRlg3PZaXkzhYAxy6RpxlUPWdUQ8Wlr9+wAzO0
s38Hv+V7APhUA6j/z+oq7LZxJo1Rs8DfYnR5t7w6x0k1jfBej9mepZahsD8ZUIyQ
b/Lc3N42ieNr6NBNqJfyLkOHIpJndxfq22ut3w11bdikR/FDKAvQu8gSGL9rST+J
9hVuXVdGazasFPXXfzDvsoNPOvvUeKD0c8la56rmXOVqHslOQ7G5aAHmCtDQKwOL
JN/ISheZ0EC+OqR6p7J/a6fUoM16Z8hqbLEqfKeFJ06v4prVVocEYAVNAJitlGa/
MDCas0jzNcuonflhKQlfeHIe8cx9YvwcRfL1De5tNvVGa2d/rI0nWhuYKHm01gum
Fw04W9VB6bpJSw+OSrt6Hc3EC133dzZX9sPXiCZ8Z/VHLOwhPAD8XtTVcdCVwlZ7
Him7xBa9yqqlHl9hTMHqy8sT2jEwZUPyxo3FbxzEXFjxsbVTnGd2ai4nM/iK/piJ
B8XQo0Rfp9Vpw5gKUsnD1PQXoHpg5bSXg7Q/UAwq7AK237id321paZBMLvCUQxwG
ImjB7GCayXYeNLMu21L5HzJEE4Ab2P1trEmkbgRv1eRp+wZbzoVGtK7MUJBVoBC9
ilsndMnvH9D+j6N/NV3yIth+3KoDyxT7EfGCMTXg1Ta5Xw6h1u4jbD4x11uyo/Sh
PXwRNIquXPm8xHC4wDWqQxf1DkEyHBLeItXj6DOMdu1K7f41bNKy1uE18sl9D+Mz
/RqHJ1lGazvuQ/riWU95BXRDABf2qy7i5y2s+OspZUBtR3dpvkKE9r+W0M1Mwiqy
Vp4ul9vWks71i0Cu0OXfDGv+8d5UstXYmF3CjcUXysdPeVMFq9mt+ctUbUl0IygW
EqWXd4aDWlSj0VUhfGUtXTzg6Nv84nkqSSD2NY2BoDjqeggBmhJTEQtrb9jRLFTr
xrc8JlnKlt5VM2tBZNFI674ZYuj+mWeR/CPq7P6hrAT71VqYgzzpwf9S2FvcjPBY
ckEPNTAUgWlwHjoZGW3B244wrfL7cBIwa1/frGYGz704TJuuczWXcAPB7i9yLxFV
fcskVzDsAHVmX9jEcDp23c9qnneYU5DL1C+fCeyj5qeSqIUVG/N4/uHY8f7Xt6qK
g/6Fco8DH70+Qgir7fA2Fk0eQma/ulaODbB9F+NGDv80WhtA3Y09T/lGUWjH/mL3
Wk5PBT46pvAP6B5hUYlwXaSSLIC8fXicUhOo/HlrG76Q8kDarTq5Lq+zQ7hLK7Mf
aNrH61JY/ud5IJBsPgszT0gRikRR5TTsgnI61HxVMDpdgJbaAx6TPJ9n9ulbORS5
iRViTvBTgcO+TcL+M5QQnsFxt6MzqnPeAKZ0jzRlJmD72bXigucDkOtYknPkXHl0
kBt9OSpIhnpG2//Oed6QK0ftFtu35vclG7v4KUTM5DtKUVlM7DT4W5zaLWfx/hac
pL0oVl+QxFLHI0asVPZlzoFxNEwBIJUK3OFMzdby4quWG9eIEpfloNbD0pm5H1OB
Ld135L+gicX60th3FfdRoX462XaRMDYTVuXvoi9AXmb7/1gQocbupQ8XPwTKneh3
d5r8uB5eQErRvAFXpCFweNa4yzO+G8L5+VS4CUO7BZicmviV/Jz/UC3PUIFhv/Xu
NmHkpknCVFqgG0ANAZ9VxXPVKJkAhE2MiuO5PnlGZXt/Hz3uLwpxPfJMGjF0sc/g
lAPwTyXSEQC5VRTR0R8E89atlQjw58L1FDucxFJPLdvY61QSfCgQwhmIWgpAr6eF
hSiF1cXTU6zblU+mjySTvUURZKyVQBmsRKygsWOPwPG7E3yBqUSovaFS+HTAqq+W
+Yq56A9Q2YBYYZ3Sky38LqIzBzmBZ6ptjZWdY5qShNy0ZyjiX/lZoiAskokFyWIX
WsG6DJomXgBJuPRguFyjwgQSQFGjnVG3T+T07NpsFd1Mxo3K0IgEmluCUubJzqiR
FWfwNteogReLLi625ZrdFEbDU6ZvimwXM1+zcIDWE1C4N94RADDc0TFAF/7jEdAY
/SX468gci9zZyg8WK6RrBTSwGgnVBNY+qVrq2Z8DrvyyuJ9sFKqI3b1oP56dburQ
m8UYoHKII000md0ALNByCMXFmcTW7IwnFwqYrQmnUSKv/3jTtQqBKJURFJqcCws5
chB11y2nXs4Kbv1ygm7WWcQakOVfKVch0ZZy4yVKasgrCXIk7Hv8rWVq900ibdBs
kCpJ/TEePKZYKARJeOHj8LbwReirJEFqvD2UkvSdoPrPjeqNSRNvGVugyzLR0vF4
mhw8elkgrpdt/gGidDhkZZAXhmYm8hg69U5Q8qpLWlMJ8tf5D0Wv4Yc1c2kzVuQJ
y9kNr+oLeqxLIoIdW84+xumhg3os8qQz5XYOjVjjSH9d1bNJXTW552aBweYdGSDn
bpxhyE5ZzDwTUwTLTyPO3CxKtzaQmCNOtpEvz99irMHkUOS12loMGxCilXj4rjRi
uNjDZZNmyho7YOFSwJOWMV5Wiq9Uy9FDhwxlRR+5r78pHXyQNU8fXXgaXwAR6l5N
B3Gr+j5iRAf7la8HRkSjMNdDpO0Vaio1QGja29vynGngPkshPNxW95TdnxWEWOXE
yQSKlgR5F1QWudpgeB56Rx0dpMoQZcEzW0Jor91mBW/aS9iGUl1DBUQHohv/lpnp
hhknViOGlxBQtH/qH6dPDJOzTyG5g5S9c2/hgxyi8RuL0oehQdtA7hxCMDDHn66O
FbTwsz0Md2K7u6fjqUn28SmhiL9WPTB9iADujCrG75mb/bvb4FjalGIfrMCtqzE6
Qhrm2AfiEv+JTDhabtnQXrxyKIYjKHq1uAW9kZe4LLS1yazygP9tB0ZhTAnng9Qu
HPh7D7fvP3TXnQdDtzbc83hkd7Dy/cRHtmRtalAfzM+Unj/gqQojbUzmJS+UAV+G
qndeiRFdF7uAAG2MPkD5nThuzBJIh1iMjOB8FaTFetQZSnLGr8St1CcEquOIMUI0
IjfDoMJpBbos+NLZN1HSU+I4/OdNjpxAnRBB1ec9Lut0lXkX2dK8sIh4mjgqhwzD
GEB9NUkkhqcbXAn2XBF3B+YV+dck9dOk1EvdR7MGwHWoRYp0H2X3UcIptv8WtAzW
FpFO/9spJTj69Fe1Joc3j5s2uX0WlEKHk9Y/vJD2H3nOTj862GZrCsN6l2f6yEvk
cI1lgDdhQFYhr4K5oDpQUqirDcYASKfcz2bluIOKxZ2uEfHZsHde+SbG8dillrEY
jsn59M4/44n6RKxL3S22XEvi3M6thve+Cl9ECxpXbkmIkhrokNDvs1e39WQeCBm9
eUNdcnVCqzD4JXEd59Pa1oyUu4dWFyLj8IkC7qXa8wpNkCszZqQWW0Kdx+rEOQ/y
oeoiSXdMJUXgVTfeyckJPD2vgHONDkzRR/06gUMp7UdlXEPK706brVWIKD19isbA
7mZbvuARrB9hj+U6eSgNH37CHQi+YtTYg0aTpd1JJ+Q6NuOqbgdaC5ArE5wmjsXE
ULXetGX0U+kCg04PvrWxd/dA77J56y+Jy0qAaamRuc5ewWPNbSs4jsU5XLQ1JmAc
B83mq0rQRXj/rmfSiuKG/VYOQ/W1iXuH+o95s4oVtP2lQiu1BaDstKiQLcxNhfE+
oGdjfEVYAswJDp7rcRd8fwj4gY1esUhpG4k66eJknueS2k2SR6N1Amac6Rbu22So
8RC20es0iwmASLJr0KCh8A3Vw9nVTfu6U6sQVv6I3Cu6kiUZAxKE3eleBhk9kL1j
QjiFSm8Z/vfveojN1CWwcCYlvFbbs7pHibo4noVOnl60DVDzErfNER5+6u7OmWB8
AsEsJ832HqHrd5hO6APaPSAjLTiTqI8ADkas8Driyr5KsW85Hhq2oEM0GIJ5MVhO
x4vcRLkLO3sodfVs16kyrvIO30jaIPM3X0QgRZBuhsSZJYqJ4RITLizaY8aGKmyd
pkPY9xW5P5wRyqXLsvHw+GQGQm+3Ow58bMPIXq8on6OwKJgDAXcf+EP54B8SYxPG
ianKou2B4ngPBhL+vM4waGpnPZQ2sxqsM5E/N/+KHep7UMZ38dKCMsjSwkLhpjct
FJoP1MyuWBdLXFvUFb/YKvRzlunyt63XfPX78Oo6jRGQY0SOo8Mrzpv9mpvR+FGV
YRMAtWf3Fzd78kbeqTtNlP0jDkQtBBhw8d5LhqwV15jTQuiZdmAtPMOohZlM+Qo3
VKcDesDyYfgCvt9rFj+/360YDYysmgfnx3BQDRVyWSx8GycmL+ZpRx2fWo0889QC
ZMOKQgYpsmw+GUA+Wow/2ir1+RYqURYcvM7Xn1zjwfPIQlJXh59NiyoZSdA0zraj
sfiMDnnMsd65L/0RO9oRRpHGOjcA/pWt6PbzD4nI1NkDcZEYp00wFPoh8KLnup7m
+KdQ6wTb1Q8mMOW9YIy+PR21vLxAl2IFU/FHj6qv1xI8djYJDe+jzpJTMpvv94Os
NtNAnlxymIH3j4YnwKBrSA7/i49oUcZaXw+gytL1uXBzFx1bAYROSlpI5effat23
POhdOMpHYw0VNdOuyx6ovWQIYwN3WXpCBVTwlfLGZrBpU/t7EE+RyDfTz/++pfHI
1FFJlvoLpM7+2ic+wHuVDIRcMYEI7pRfnE1szwHOVDjsTKoKmWf7RU8pcJ/jebxA
8+k5uWaODLvjRYHAGwIEmk2F6SJg3lwDzFcQ+vbj9TpOx9v15dTTE1Jb2sSsMbcK
4Xb5UKjefVkav/kS43qDS8eXC95Q0ahjFmnuxIXFYSFK/UnC/vXAHImOFxkV4x+b
THMMRv7BFZb54YU3J7YgMRLHlJotSEbAaJ4F1YENa/0e6VpMmpAbs7FDHvPuYTuK
fGIpNm2wuCCDLtXPYStln9VUJCNsrbc/f7Lfo+orp94TrFoSmnm5w7dCx2V+A+rV
7lzG/2AyajrEIIuL5Ib6j+JEmK6qXgoLl/ndxBsMrO2KzuHIS2Q971Cg4gGU7MEJ
mYo0Aj+W/RQwD7mq55/26ThyMkVhF3vMaLdVjpZ4GoXAt7mcDfFcG0eU/k6yUSR6
VwlzpBtaupLj9XvYAWH+BRYeGPsdZDzRXKC2Er+GvU6b798ytwaeGvAQS2K26xCq
zrszwpMVC1DLZFCCwOTC2d9FUQKNMnjLuNlpHaf+XE+bqAR9ju5ydnDCZ+ti/0bb
QNcq1E2neLKkW2rJh/W+id8KnLSya4iXjWbiem3tPl+vC8DPOBzW/poe8y3EAq0o
YrVkJNsR2anqpm0HfiC9TBHVJ5hyBB6LFMC0mNkck5cpqebbQ4tpXMSMfxN2y0ge
0PksMBh5trB54WHVJ4fjamHfFgOLpF//vIf9ibBTsE93dcmj9NdpD6fDVBpAm52P
MPtsJ6HwC9EyuFMu8lnGQ+wBM62nCB/O8GsV9Mgy3/0uwAkhjVhe2aP0S6j6h2Oz
iM6lteRHePhYiQMT32+NawsrdF2V7pFslCDtkacTMwr47YlwfXkIoD4dSp0WgFq9
TPqS/ivMmIDWi+SKeKVqFdC51h+U91mgkhO93/9y3S3dk7kcmsUWElxgZeJr12cJ
hLITCRGLd6x2eZDSe8lNxLbOALNdU4CjMq/0cc/KG0ceGVxMWqVECABSsCi97alY
22Feca4oW3UmrUYxMusy7RsNz5Z4eUgFJW3x5IRvkG+1CoM2HOAxEPu/01W3IwmH
hzB2WAM2+uGVqlqClMMmQ0phGSWxMpRs6HD4htEr6OxaHd7WObyNziUouOI7A/em
GrEuCQ34UFeAwduZKqwBgnaj6BVgvyZCzXcyb0OtPP4mykOcCQrRGyhF1oMl+cHP
gD7j54I2PGu1TQf9pQ12u3RakafWiJ36FXt9VjK6X0gA0Ki4immpzJOXwfLI05HL
hyZgOQWwzfNP1TQZT6il0z87HAoIE2OO6jUgQqwwCyYo1Gif9QJ/iIjkEDTLWW/Q
To3lMRuyXBsiBDzafQhtGyOPWeP2e7QYMQTUSNE3hrMVZNFamI+RpL+ME9wlRe7l
H5/smew7K0ncTEVm6/ic5SHxc8dnDlVRW5DIVTvrf7mHgSjfY/aV4jUwlZwXE+rv
W1KPwVHCROjFzWv0ZdgxgmgPt2ttz/wBft+92kMXijDR3jkV769u6pmFJ+2eh7Qe
zh+D+owezNnDG8tRFyrjDeG5b8FyYPXVulMSIC6X9mYmhAmDu68rf7CgwMRT7eR0
tr86R+3/rrIR8OkbRSe5/30dVt3PKT7hQJi5eP7F5iPIP7TxmqSnngKxPmIDf1fy
IVq+Nviv1Lt8pqwoNK0blVc+x+58YYB2RpsEUw+k0tcmAnH5y1gQWJQzmlnxMu/V
zf3MiBR3yt/lB4IEMgjy/ciUG3xpHunxSmm7aHgxeNbC5QjQhQadcy4VeEy2B7eU
O0eYSbRb/10+RCZEVXmcSSKq58TlLR/fAWOy+XX9DkeEHygeuZgxZ03ekSxz1iDL
DJQCRQPkwpX2uKb/xcFsym20h9uYVzwRiOuDRYC8ldWIw4HUIuiQNamEdCKMKkor
zkv6grzLfubjTyIKqoIFVZBhgaT/L9lfJzYCiAQ1y742FOkkF3we3U4D6R9UHGvK
5Ykpv8jbxJh2+P3eVrPJoEKGQGZ+7pB0IlF4EvF240jJCZwhGkYbgRDWno4fiX+Z
o5uKuXLqZ+kvKTBnqcf3jLJMUCTRA3/+geySdpm/IH8UOdsT4Z/MhMpvwxWRbmAc
XnOXbVx3ZAnrUe7+iuERCEYomSGkBNn632gvhG1AsXiwBx7if5ffTayEDalxFz7h
0Rj7Lsn8bSoXihnRj0jjQrzU4/o0SLk8R3/MOBdgiJsXRkreJrVJis8nqyX4tfMs
w9gnV4+EProvmIaHX1mDaKo5UUzERHDI3y2fWUVAabZDAbwmV6259U8dHun+KgTh
JnjbATptux8niDKbNOMlccbFZRrJenzqHOLby5b7ER91DQ6+M35HDDYFPL5ini1X
hRrhfDXtJDK3n4D40Kfu/ToNsydcZugHF3Vv6XlOWcs1OhY74wun0lhpLmJz85BN
9iD3tbTYbQfc8k2xY6uvSmdWq0oTjZkxuK444OoEWyXlj0c1dePGcqPclFWS47K6
90LGnn5APAjzSaAUjeT3zbUumMmpaoSb25crRA2fafosJVgwJ4rHwiMvAX/mhY++
ynwDN4nzGIfSnHtnsWIw2N35tET9RiQXhspWp94IZMNTGtyPqd9m1zwKsI0O6D8a
H7SSZ+p7dbyQ2tyHYm1eO49R1FR71N8hwfRfNEXxVLtko9KwnuZhNOx0oTbngIzc
Tm7Tj0WK4XWDpI4BmwGvj5WOVqiEdHa4JHlyApZbHT1RvEBtMxzM1iZMiAM/G1GX
990+Th/OaIzkTyCzD881cgztiQSTWtxTVm0laO/WLJIwkz8x2y524SyROEntPhw+
L/Md/58L9RX9Dn154Fyvij1O0ZmCUcvdR9sazqwkyHBdqVdCxUjodrb9MrLv1eBa
gfYFGUA9ggkVyslNJV+NvRc7up/cBlk6IWgBxlEyRFKLKuUZL4YC47iKrE36l8vk
KJ8LqVx6BFt1sjZHftcLvdHjqrCJvVGhXWB24fPN1jpeyL9Ac6BOaignDRCQ+LTQ
XEo+gt3R6bCpKgAWbk/KxTIcoC9Vf6BKK9kAfXle1m8/KTMDtKkxUtfbH7SxlPMv
NSNq87LqPCHgqHSZGovrps9LN6neGG2vkqx/Fj9LVq0CsU5S9AJM2b1FfXDF1rLC
6KnZgWvkCAe5Sh7fu4vNm1s8m2cxHxF/3MPfIa97oMYc3N580/k+TXy7kwAEg79u
rEbv08bKeU8gI0XeDQyIM0mhnYPTGqdRQ4MvSyCEV6EbpV2+mCfHG3CticXR337m
75bjdBHSwSZHpRxbzlcfi29mI95BhVzYkfOUYbdOn4x/3J31ufKeOiB8Ctesm0hr
arHtiu+YqpCrXQ1x5Oc/qGdrSAWaU0vQJheO2C3CwGMqzeuW87cgZTQxY2lAs2Qg
Yofs2uee0s51NQ5Iz3jWU9HcL431MC2L7io6ZJa94IWYRv2zfrZs1VXFZYzQA3DK
mricK+ZMKDFagfzxR7x+h5hzxe+7L9warEH3PpTrd5yQwCdT90g2QrapPr6RTOpS
h8rVNzzoMhw++S+g3waQXF1e/VrSDqvIyKGIibo43A4jIdWFKLoO3aEyNRfxAEex
UOtHyjoZ1+Lp++cPssxO2Eltg8eWulgm1JsnJ0x4jEOoBAwa2d8qX0FOetAXsCfw
t4yl4VRkCDnLMMto+dXzHKFH6/SsgQPiXlmXykuPywbZOc/zDX/ddSxKZVsd8T3e
jCs8Es8XdPwJKEafH6SZkau+rCDwWutUnFn9Uc1sp9sAOJ2Voeh3VLdH1O0rQioo
ccaJDyYbIqwmz5Hc20RJVruJ7bfr8tCJb1CGTJ8k4SB6NR+USObHP5J/JhF4khbc
/hhzlkzZ4p6QN4Gltn+ojxcbXzIPvIaC1Sh0/pwIrBfc90g1az0DQyc4TtHtEe70
wLSHPAvR0bc4ml+6v0DQ/Elvjlnty00M5/WNuz2Cdfw76pFsNpbI8sdr1FpNbOBc
nXLlMpCss08gx/PsAnUuwd12J67Mz7i4N/JJo/DTbZUFq2rhN1OwTZH3yoo6Qc6L
GOi5gGBmXR20iR9gQw3dzaldUQjjaud1d2ai2g8rI7XkDaClYhX9qFyagG9wlgK5
dHSnq2j/tQQkc6D476flr5B7PzZcZIZiAut2BiHUTlDaj7GpYHGx2+wYEpTzWehq
FsyGK3nXQ5Yt1ztuvL7k+ZGlshzLUBTFQnHISapXXEpygjH0BoPi2+JfjMsA3kwo
kybeLkcg2zLIGfh3dDZer+NLeeMQJ+dvGkzttzDQjqxEwgoWoAYNh0GDPWaWsUUs
qAp2F9NUrsXe7eSZXL9QXjWCOaISkYbawl7rDjdO3yDLNWEZgg0Argecyc8hIqQw
HsuYG2QBLYMNRWBPpwOs/+VemQBNcwpKvA1W23qTlskyfCEMxTuDY7gw/o5cFo/s
J5RTEgDhXLNZtb2hsTGeRMky7ojY09UYm2U6xzPAuigjRQEALx2IxijWB0C1vhb6
H/429gzkhSa7psI8j83872b9KujTNrtyQLv+ZakC9EDZFp/A2iHpqxNIKmaeQ7P5
FDWw/2ZNCgEZhHj0gLRSIgGNE43Kdy5gVI87J/m2uD6kCNANzSEKO+AcjVb5NcTu
fJ7rd2ANilb4f+eh9xUfYoeHagols0meJOM650OGYobh9HWEmkxwnbbM1VsMWeck
sDkvv5TSM5TiBMkTVx4qYkUBNqOnFYRl/J1OSCRKk8/iJNTAWP0iZgExtjclGA0c
H1/G/foLJnZwv42DGyWj3Fo941Se7B7UQveIuWck/HuQ0COOnGz4LhqtljfYPk3g
o3+O/yv4eAIhRn9N+XfmGaGvsw1dUpwR8mxsYKzUuaMVlZXlEjtGBq9PrYJChtw0
eU12ymsEbY+3oOoFgKZsrsEdvUfcLA86s5Ql5XcMFbpTzMsZmLciarRtDwX0F5mw
0qQKcFr0JZpziod4GzDletPFZeHliuNloIyxi2DewAxG1XMHGPEYaBaS46qrgdr8
JxfCJPYKdecbStfTpsYxWvwpqlozQN+9SL2OKzqOSTXskX7EjrTNi0HGrMzoLLei
wdN2sd+MZEaChMCzPS01rDRu4qV5rHNriKOtHnELlsQoP96S6U5cdj6PmAyUc9Z+
cA805rIFKWEDFkqwRLo5gaMI7IJMH2jw8d7rXxpabUuNdauwBFCNcRe6L4Zj8YnZ
5I+4pJ6/q9oKvng/FRPo+Y6MfBWJoPTHU0fbWche5jKooBG46JkcOf4MUVyH6vuJ
B55O+c6EcDUs8MV7ZswkLD4jT52Q+4KBq258KiiMPvXn9OrPlMNTR8nkgNamUqU4
wApcO0bOJNWjQ0VrS3JeDpZpfOFrv9wOUtLSOXuBjmGzP+9/3nsElKeVLrFKbeAE
hpW2/Fdgtud3n6xUjN/LiBPh0X7TDE6U+i6FiCysO2i1YHkOOdWZvn9NQMlYgt0h
ida1V9yrRQHqzNtcKqqIzdoa8+EgQllxusr1rC+H/yho73LeIXc1PJQwLFiKN+NK
Tlys8A5hdWkcf9MGejqQ9ptO+8106U47qrfI3+5AexySvQ+EmPKLraDPUDwhVHYK
u4IgmP+BR1HV3bi7U+rBPcot7VwXthYJeJxZOxcfDVutRWkZS0ARz5C1jVvXqiwp
RCJg5TqkfBqlfE3ydBts3O4MIFYhMqt7AGpXyXQ0XVcKH3kkWPXVmRAQigjwDhXo
MRAP6QnyaKhjefPCDraoGDtyS8HlUD9WQXMVzVM5JnAslKAFA3zZX7hiJua+9Iel
sYE4++BF5JoMkG+RsHHypb1i83mk+GCwRU3b4ncIZuQmjOKPRYkKlWQROrjkMNv1
5hV7Tvonm0Ok1Io6AP/WZI9oT2McH44R/f8wfCG7z0WlFzBezgoM2mHnE+wi91Ta
tsoikAwG31fOiQlyYq3q+XLk9syjaBX5VxTVeFWqfyghY6ZO9LpfEbU4D728r8Kn
ZckaURgIEalo0T8un1KSOJih7dZ2hps8RwGPfHP73NTq3tVXmdC85nqOB9asK7un
pm20g9Y7PXmzBe0AL6/YrswkUEarzu8Eaemq+vqZx67FOfSLGVmjLIV6n28y2RCK
3DGLmv4Xxdr6SJoSrGfrEs8rjk/fKlYhdARMqf5ooLs7hjFQs8f2OTcjV/AUYaIr
CzWtjRK/BKtxUoMoiGvg4lsshCNgQqye4n7HgCMQvd5hBdkzj13DXsiRyzRHfxxq
Vwl70TQVdsaRIrIVSUBxWoL3sbCW/bWdMtpIAmNiwQsXg8Aq0Ghvr8WjS8MmluIZ
mJ6WyLW4m4oTg78zX0DOE+GW/HWfxUB/kS30IUALpiFQHjhvhNI0V+2L5bIF1L4h
jDKh1IwvPXIJ8CnnCKcpZHUnUd6ucmK1hGXYKnmPM0uzlbaZvNKSpkehaXpTzwWz
HeQwiFUTRh/GOjPZSQWl32sCIeN8Okf//PXwQvkoT9NfB/Gtmbwbv5uIL2TSe8I9
S1BiftwAW95vIuiWRzmvAhOzenLwbDwOhLD0edxyC6odP7D0FnAJBm2t++h1VK/v
BRE3sbytbrXvV9OOWWKSsvpdg3BaVjsabPTVnT7j6VZjlM68/KIpTBgmeHIwW1Xb
vmNLxlkWXYkSdpkSi/RPnIpOj9fTbWsrfE16TedEuguPgO9ZXaVuXD1Cg8GnxnOS
jXTPgmS/TU5pkxGq2CVAPDjw4kEBAJfxBQbLEZFfvrJeYcHrV06OpIzxY3CjQEXc
ecBa2IEdLUzqYDwsVydsd6Dp6CzDjzCe9lnSe9++sttOwdY9Owj2sp+WwxyQlwxs
vo8OB+xRQS+TuR6YNpFk5V+gUPIxzNmNwEpdfECyHd5XyVb3xyqCZDgz2AMAUNYj
k9nDiR+wscNDWR4BNurfTBIeDzJVJ3PJZN5c/Y3PaDCkunCRDe6+jLs3wwxPcVGQ
QZu0Hfm5k9A6ZZ0qQEXRrgwQLEKUU+nPkUCqpiN3gfEP+8B4CAoxFIAYR80yy+G4
TNmQPGCAkvSvsEzVz/27s5jwa3lner+kcv+GjAIXhiW7SZ86P/oIlo1n75I4SKdC
wBbM9oDk3qIgOuYTNZdzapeomi6tToZRMNH1kZt0b8+sdZXYlg4ST31xO/1I8xAK
vFYrRqPbOOISvb06eTrgWQ==
`protect end_protected
