-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
bxYFhHdRc97lUP+9wIiPj1ATeCWppGY7y98nRZKDcs68AEj2aJOcAZaONfcNnjde
pPOZsVsziAdGG8CSCYgna+1iihtylODH/TtO3RFCiryFEujQ99kfIlLKPZHcWt02
1A8eIZpoX46NwnVl2QRPL98W4ehOBP6kJEAAKYfcu5k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6812)

`protect DATA_BLOCK
1VNfQCllzDgSvyMcW4gwX5EYG39sHNElGHJK4jdHTF2DpsI2k06BbCoRUq2xjn/D
QcaHJM5UfQNCXKkumorqlsDdDtgU2FTsWo1n0xbbsCI7WBNzwePo3I8qRifKpilH
1/vgwiwob9R3SnG1yFbjZoip7YdcHlSRcJ+6PJpVnM5JJ6PTtT1i7Qm/tPjXN20m
S4AJFJi3xuv5mcSzrUaT/7kIIie876oE5ShUStVXB2gWpvekpwHhsYuF8gkYabAp
H41GuHHGI6EdHcOTyMZtwkRsQ21xUfUtUTK3c4ClRWMWyEqB2X6H8K3B9ZTTIS7y
dgR+MY19iCKqhzA6NnWsgPR2uqrg8vhdKsCFy1oCsnMazFsEdZKBzRryuaTgNpeL
UHROJFra6JCuVyLw/vvqNHpA8RbPB6SZekcoG4r5uzyrnxX/zYOLx//aygWlO5qf
36cYcRj7S+1aU61aKT7zmKWV1SbD+YMj53izTVMU8LXINZO7TWSGgPD0B8ueLCXk
fVElq0/t/XC8E/6VBxAvel2qv1O27t1/IF+kkBzuXQa+fO7gBKbXcwNrbj90ZvCB
dQl0JuoRQPDVTPWHwLZgq86oiyYMWwVhnMqgswdv1RDvdp1ysxLLEgLZ1qHg2Sty
cyTCAy+mt6fAGVJP8PuMXaF8w6RB4E2yrGzJxhQf+9h54/5n6YNZVhq5Y7zIgHk1
qLfU8OwtF0HpASTkbI3H7Sgb3ORUrfoSWSggaBEmtKADVMwNi2YowBey3Db9T3X5
4ah2zGNXyXprPZlsovSmIXt1wMkrnEbzC7gcxdscmjma8/TNV9+80uEh16Hdd7jR
puwwomQZuDo/wTldS+ztJpmrAhpl8khyu7QD7cQHJdIAIWRlv81WTUBP+jXXp17Z
cNmKPwARxHrtJQ9lvN5J/T7Rk58plhYAZLKAR0td2YeHCNLlMN1NtGVkfTM5Eb0A
RsID93cpRtRjCAJ7ONvQ+3zsrdIcrlAp3mgxnSjmz+sTCu7j149wPpKs+8KlC2Df
8m11qUYGH2NSYSUAd+se48H0F5jj/maZzZNxySsTdvxUakQQi7WflVbLNQnIFv7f
toRfALSo6j6j7to6rb8JdYCKYPY4Vuz7oue/LTWB3idVQlClw4bB2a4kZLeahg18
AkWcYBlFRY0SPGJOos8d77H/78ezs3Ud2G0Dh9f+kDWL7YtwZNfm0kAUnBJgdIOK
T9KK77EOcfzVn0kdRMV8/2jaswMR1qbzmbnfnQ8dZtK+dpFILPhJxDel1zpyrTIW
KNGwmP0yVwLMO730iZSSxuyctstS40KKlLLQDhrtyqMJ3U6DC6U6AeVJhCsEIKBZ
nfDaHY/VHlR40lPXk8yi3T/no4IUDRuILNTLsb3H05DX+X+SITCsNHMwrW+QcwNn
ZsLPf/jkRm+jEpaefz/SN0we1piAu3xPObVbqdhfIg3VsS8W5X4RMz3nwQVIPDlr
Rt1OYaaVJamNWk77l03/hxo0TcDeo4TqN3jTQNVqN054DNLF0DBuIO/RHC5XYyUY
QKBkTbr0kYqH+6U4EyhU9TlJJi0dOgayrezlWfGr5SbDN79joSkRl+MRVKrrxWDW
pqT908P0IZpVyUIwsg3RO9S5LDZ9UH4ZLugbPhUTDEMmzL8Tm49HFjdd7Jj+1QGb
AmJ/FCOTSwsPXKJ0XVgu2OYUVgokcdz97KS82/JfnTE9zN1/6UEBmoIwXozeAFRr
ssQc09tf07kYGh49UDedJ3s5y/9JlBfi3nNUxt32r9atghNuOW34ppThXetQN+0U
3Cyki4O2r7cfGNvwT8glWsbDv/pG341ZeFP5Dq/GgP9jP/VzOETg1gmpMdLSxUD3
6aBmcJ6XhNCWL3t/wRocsl339H+ut/diEBSS17jYd5WUIlJ3Dv3NPc3ttx6iUew1
+ajR4wEHtiDALcTr5WPa3q+ma91c17zEbnqdXk2pcSq/hvTYtwGhW4PnOD/+Eb33
iHtyw/u+YJN70t4UwI+Cqva++hBe7dJ2ekF3UcvTimTSNx+ceBmw2B2uSgu9pkin
WjX52DRXh9q82C1XXrP1yjUvjDfsxyudNDnyE7bEYNM1O49CeCQn638ejWnzVKkW
stcMR+dgc2fM9MXT6CXNGv60tb2kAfKADFF7jeWO53TOVqMmgcO3ZnX6asHQDm+H
Fc/V29MfZ0GSTAmxtvfFiOzeJ04tuKt2VNNPXEgYkYGcMMZcwC3SxPW+mFZFJ9JH
PO0YNQj7hrn7haSPb78s6YDOwucIc0kqzoGbwCOd5xFDRPqYBFrrp5/QBlqRAI+H
zE8bsZEkds+fx0HlBzvdr8x4tdpLOydMgwxQa/AgdJnlSxWVSXfn0g5A2N5xA97V
NcykJr/ovE9F3uTPLLOc1GigBUZRhL+ZBYLaiYNAJRYLsdu0RJriw7s0aCY37x5w
0kUuXRhAqF5/CE3ICZ53TPBfBjf8oZngkCBurdHKlfKbS2OwEgBiQgvKkGLU1Kuh
m1xyzhKzBU1T4afn2Vbg1cxlmWeQjG6qXz/8CMZ/WEneLSm7YdaZqc7D+MgYpJkU
HIgT7Kv+IbbhxW5Bumkfzkf6KMhLhE9lX9mWP4oVlOsEJUP3pJRtWV3SW1HTn1tA
nZw5Wt/9f3DD6rbiRcfhwLDq/CXmYxdDni40GzHQTxl0U6LevkFPsr2KG/cUOIQA
d70V02PQhiiGp/hhU98c0cVL9N9AXeBgKimlsAY0ZBoMxSBc8swembJQ7c8MZ3wX
IHkewfjhXcCysgOXOjnQf0oJpUAvWAuWzgi/sQ5egoDYK11wB1Ny6QuGbMPS3/Lc
Vx6xAuUFmuEdnObtvTVveJwu6VQR/ncGTzMxhwfydPj304QqKS9jscbsEo97EQLc
Ixprbr9n7jgMCbWGp8lVHlLUYbC1NRs+FGl7YvIWW60H98UjB1PymCPU+pwCH1c4
ZVChS9RnyvxlC0yHnCVPkcoEP2bKbpiN0JqonoSwvje0ZTJ8ByNZYDDFvH3c4khI
8d4cYq96VddXxaXAYhFbCfUwfTMMOd4+I8i2j/9Mw5MA9XrFpRyAJKzBB2TyKhXg
KbLm6QYwXcX8O50uqNRrJifAXUgW69ZXFZvrZO8HIWliD6pxqFABI57QHMZTUcms
4XI9oi8LCPQ+mjoanQz8G+k0t5IFUr4q6WdD+ROnkCXBegyQBYGsAR5MpusaNQIr
8bOdCWQnFB/KiIZEKt6+meEm+YUC1AyvsTCP/HhOKxDkDNIuReKhpfdC8iXGub2f
1lbdNXp7LR5pcVQgA/oaQZ2nLPepEmhqYaKz0n+DIcdjIELeUOBOTmplu+jvhZtX
Ljyd4VyA6jelzGT+fWkNx8O9OD1l0sSj6AsYR0Tu8oQjsxD533W5Eegoov0hT5dl
f4iJuSXtrfKoLhMeFS05luAYBBGigCcl0lgkzFls7yVYAI53c7QdGbMNV3hcxb+W
yZuBPxgpTg+o4Rf9kMmvE8I+UkLRZAtUkKANVj0rXij7MZwSdLC7qnyxfD1iqS79
ftCfYXJ0OFgeBWPMWB0mo6adbJhQm4yX71DI7ApLMuhKtgglSquKxYwl6SQZoV4k
Tm1PaJEypFX0bbp0rkCYZJJp77y0BHqOCAyIaNRMeQaILKeNTC3Huz1aZEdTwbzf
7rg1VkihFrWX/ZNcHAjjWRE3SKbYoJSZhUN+gHtZjSA9nzzHMNULTCCaTL6/l9tG
RCCrP0BOxtt4zZkcSPhzO/Ez90y+7/vGkxIbgFUeYIbPFhwxBGQKUGmXKdwc6z7E
JcX+aKUURHE/TTCT60gznAmrZccHoJojQX7CC0E3rmjrYRRLM2O5f9CSR3PD+UF6
9eRRdp3Ws9ZAuDOry8muPN3/ecc0z0VwSx6buKUF6wBb4vcg6VuIhfvfj+73gQ1w
TE4tfSR9uw4WFl99Pt0oasNE9D6/muINEjwBiZaE6aif7mn403fbL61US0wXlJAj
Hs+7bhgXrtnqOTBaWYewuC7tPTxp8u8LX5XHi/z9NFYTvWPX3e1WPHaW0namxnJq
DCLUcrxYIhNKjj0FVmq8xbwO6BVsvugXMRleM+w1K8n3wZHiMkECL/beRYFgCn+F
1+T79dm+PC4MBPKKps9trbmcYHx5YU60JP0THCyAcnl5pvTnr15AMcJexlu+OpJz
zG71Rwa+gCLSGrIFTd3EzZ/YIsSdNFKxDR4YnLQN2IRJz44ZQRg1Az+sg3e7s0NC
NBxX8oZqjAov5cbcKQus7g6gkIAG7JYANaQtIMeDRfvOtH1G4gWsGiPdU2Z6po/2
RqlKJjRhYCpID/aKpwGCPZC58U+pt7DuIzMmhIrSnkzIuS+SjCWaavQ95NgsXQVL
i8pQTNjKdduDr1EJ5lxMY1jhEqoNGWNRw7572zAdGpw8/w7rSqH2NLxRtrhlHwke
EIcQsBi66UzAbVkiI/DoWizjUPjng5wabV/Hh2CASOlpyjTh/2DucmfVz+icgh89
Rj5VhV9JRPdfBpkKj4QOrC4ef96M5iukhE7p1FVh+qVNYHbS2Ocuhok6+RiKI9Au
CcpQ2NOOLq5FOzbF3tkiQr6kSS23qrXSY2gJ+EZiGGaA+kMIrgwr8XTkfUhob2V/
nnuoWJEhpZcONLX/a7uhIx0/H4iooZYPILo6npaMAyRxa/4rmT5wlgqbOGe9uGBE
wEJAKzlBcUdwZCGm4wqsBNlyKCsTT0EPNQIlNOU5MnteseIvAx7mCP6Whup4NwH7
Mevw2DyE+Meh6lmh96wqjDwcgX1qVhpqb9iXOmxjIt7d/dz1MN/YVv/NWi6tgUZy
jNB3yIFAAUApJd6bWMBq6LHApJVkp0o13P30PYvEDch41prZ9yMjM9J8/ImuSSSk
yxZEbCkvyoY6ogVrHIN7LWNoRrqtHG4F6dAbWSawzs4ups+IEpzpz1rJ445sKaVO
K25Ei0s8m2/qc4KRfyURt7SfEx529nX2ghnKTpGpkf28P/6zs7KgpExD4SVktZKv
Hy+pIL/8SRLYHKPGaCPV1ZWgv6LY+lVonFg/LXFHDpBqLanc8rvdMnUzty3idPT7
IjcFtFY4BP4P6b4MqPqn8dPiGqK2s5NEHg/iTi1O2vkzl8Rg3lFQrqIG8SUIgqD5
CtmbYyWvXJD6JSyGgR6ZRHhf2PWXHClb5bdBBSyfpN2zKtynej2BEca15OXe29af
xVIVKYbcpMEoo767Lj6a4tQ83Z4zX6+hBYzE8mSd/p8Gbtt532V1jF4Fz5CIQBjr
hXGvqFZNuA2z+r2+IM9SwEIBXKKOkrnIZ3fp1dntGLheV8/Ppo7uCkWpBBNHtq1V
ZEmnIS74uXMetykULqvdWXmMsB6FICq4ERqZ4la/+bdC1zHibFM9ImJqUb7H5+c5
Q8xWuQN4w+p75lqZRgj2Z+j5uw9aT53gbFZ7EeKIOyIDgRCnUfG2KpmhSeGdfguz
Hvx3KIEq5Z4Gh3NNCBPPz5u8Z+9BgYCU4qv2gyE6jjWdOlEk0wPXxVXXg4cyBVpD
27gwkb4RhkmRz+rJwMZrBlYTrRe0CvKROgk6X6FEBDSJp7RZgSt3cXjMweT+qC/u
7gJgAp8YvkZ+418fA+XcyRnaoASZ9qmgvwBdZVF0+Hc4f7fxxx+Qpx+bBeUn0B0v
IAkoguwLnM3/hXYV+EPdAcFMEmXKFLZ/Rrv4LqHdd+bE+ZWNouhwBxxampTfAgPb
SLTsRXUoogRi+GEXRxywxl2nFw4VxU9m7qZfWH8rTH0qI3vwi+u3y+EQYJiKTSsx
n146nD+tB025onF9rvhiGF5nOBh/iqldotktXXYd3OBK1+RWafgJsd9RqXECGAsG
AbxV267yhFG2Q0Ecw6FUKvqgqj0+1R5hLdLAhsZYIfEonkLnLvL4dDuO8TKp4oha
Sn1Ba3xSDSYGkGtFmtjQxtneLp+7mOXKNgTuwgf83Ml38D+TfMEmIL1fCFP6Gm27
3xuGpQGaoqkJ1J5h7qbTaFPMqx7nEgP7Fh+WwP0yldyV4GL6BdnmKVDkk8m7PMVp
MksKXz9PPKXWCo6BJNTLgeEif5XwlEw9CkK1F+70vFqJWqNWXJmd9ru6jOsxaCsV
3BsfqBj6a0QcN3W+5S+dD/Nv2Bk9btSh0U9f+hYY3JQ0PBL3/wUJK3Vb8b8oL169
vWeSz1UQ+n9YtXGfBXfMDbZ+yl1gmk2EyGl3spvu83xggs3xwjYy914YSdz/s8AM
FZXMbIzzE8zDhp8O+2Bb+h+MpunEK75TwKA2ZgZ62IoBtltwGaIgkHksWiUKFEcH
q/rBdBjeP87NsbDJvXBCu3aNC9swYaEZtBASNg6ahHN7u0IeLXBFoFgSh9I3L1RA
ng39+7CBQ20oTai94NagpuM2Kcg3OG95zdNqcv4qcAhJRJi/KTYqBnDccxpa71z5
R+oXQ6MIgAb60LCjBlsSGiLWIkzeZtr+B88Rv2PC5nWpuzmRxpvKqgPmk+WhgHhP
Y1s62q7LyE38Fcy4oKLbBsdWlr5M/j1HAtTCzRrKLML3MYi9RX03FLKxpTaKOGHs
m4FIZJ/ynSbExoFGbJy43pxECFuGIyLt3jOdS4K1DQuuuyfbbP5XoXUyKPFmxHRv
u9JBBkO+KwKXjSzq23vZtc3LQe/jB1++RqXM+/TLDAu+LJrqwhUYt8IM9WSUSEzg
3QTFpVTShHIuUFS1pRfR2U/elmCJxQ/SZ0LxbrmvBaUGJTlC9k4JkeLv1Rj2pBS0
eFoKg63Gos8BeQHyGtQqEXCwaxVhGuqnTrTWOPDQ1U7f6RLalANHGRGBfjz3e9KR
yflgxfde9ZnrThsh0XqkO3eamkgPF2/xG1KpXHUa9wp3mDyCwhAucwfWcfa98YxG
d29DdJw8GH7fpKp1He5BunnRT8J82BCUkjURt9LHsXSrYWo5btUppA7IFy3P9QEC
GtqdFRR+3dNFx6VM2RSDEzNTN+z2ogPoU1UjxD1MVnO0coo4atTdEsRZ3tsUx55c
FNper3jZ6Cs24VrfmGcEWHwBMDwdYlO7srrybU4q+uU1pNQc64AAcZ5qbCbTaxm7
+am+GTdeoZeAdPvmTZqbuspeTXWl+0THrVqf1bSvmqcA/K5jfwGBSxSXHoVOjKny
mSLkFiKkCdTyQ2A+NeLzjRQfZTEltFmDg20v3BHFOlblb/SnGJFC8FoRq6VJV307
oycl6+ZoQIXEBCK1MQiNSwdc/aa7XAi4kpEVD74exuN3m5jWr8v4X3PCtYfKgDoL
foU1LTkI+ye/eEM6VDblDyyoVA8m1sZ4rxEVMJ/OWsfNYoOqLy3Z9JSp/wA5+ewx
PxCo3Y4zsnQbrLEiu8zKLOKOSvZMYmkgRS6zmaoLLLyeGXPQHUiIA8TZo8X7ThyV
wdg8JaWPEOjpoH3yEJR7K7H2LfZlL/k8utSRC3XNXrrvUYPNBs8qMyJKWy6OYdVz
308g7WNAQYk5qkGzUuGf/Enk2oee0rj5kZcLBdSXhWcAs1eFMfy/tLE9L4vhNYKF
qulGKXTOP7g1UWzBuzr4b0/kPOZMPG50Js8TKv+sxpF86e2DtIIBYEdwmQ7kLHTL
rCkLmCMjQ4GUKB/bnuohUmCXOclYeWRUePcLrKSkIlZb3RIEfChcK7BitcBMInjL
drNXyRco3pbKSIu6UuKTpU2ihTrPOB2fnmNTwpUvsqdt7opt/sj892fZMI1QUhXt
KXh5JugsSGWIbACHliKWOCNKfQyMthhRD+E9bmZvH4+yf+Q8FFwpzgc/aGX4xHFS
dOcB3M7b0zvXSfuw5pUQ1qmUYi0KO58RF7/e2OIJPHj2FPHn56GMU4E3WrToGWCi
7OLKS43U6GqyZ4xm9sSasvMyK97AgeHwhC30M3IYG6olgUm1ZUslp+YE0qJ82dSC
mzQAy2lNsDnL0CaYZXGZq6jGqsiVtKkgAAjWP/B6uqKaIPoAbDEZiN1X0cgirajo
qI9XLJ4suzGIHKpg47qvBnrqUNXDfW8pc+FXMayBkFoy62JJq50QPKLKm2/1FE5Q
xjvVF5jJtkqoO61+kPG6GhWDJ5UnWvJFHEUEdswXSx0YORaBWD/0a0HGv5L34g8p
K7aRNVtiKM2QutaNgzCUaeuo/H2nxDL5gxCAptqZ1xO35yl3q06bdugJRod6TfSq
7Ib9Zv/p+BZWnEiKc1LZV38PDg9fZXaTb+s2MlTh33EIpf7mQ2j7+VG0giyu8lV+
zCNc3L5f6tJAnAURTrCSSj3LSkH1PhoLyfw8gwxYMHqgBKM/xTF8lVtzEKyvBVuO
2v1QZVWY/TrnkNEu0sLCknfG/YTuDGi+suJ8eIuyfvMOK7Cr2iY32QNn2IOtpHM+
qFZciLln93yC1MzW/Ag6ezNTmHThZu/VJyHXiKCEeestjC3V4EGkDfPSuYMpaCaR
gvGAxJLJwpySRoOyU0DdZ88+SZGbRrLGAoQ1lox7shV03PZVqfrCq1fPP/xBxF4T
Q0Mmx6O9DoatV/kcPxmnFn/sT6ya85N19Ce4Sc7iRx8KP9AlNYCNCG90FxrzQTqI
/x/NzebeMQZdJBXbtTUfNxfWto3UaLgRc3Y7UNVgaXSB/eixXsQT27PYcGcWoikA
kcBshd2KyVuYdADTy7HF4+DGKhZgCz6tk2OInizBUqhOEtgm+Y60d4Enwcr0PLrL
EzfbdX4gYh0EijFfxqNn8NH0o42wFzPsHqHrvwMZoyPaIleTyDlKFmkkjFO5uz1k
qRGX1OW6o79RAfppnEnVH9qHte0o8VR/1UFuOiR8o8U4yxctZN+gzHY4Sm87UDAx
od00DPUWTVGntuwAnrXPjUizA4tw6dOwZFCdKtLJUsNC9jnOmK2EY7sXP3xZDNER
JeGHnGDcCOCk6lt1LAB/P4MkB457h6PDOVpWI/5riE1eFMpfbycJlX47bgREJh5z
iSDW07lM6e6I7gh75jg1+Mbha2W+Ip8lauptW7BX5RU7OpWCZtCiYbihMhrZxNg9
Uiy8mTQF/WjHg/72naYAZ//0X6lf7FyWawIpo4KGcpscJ/Us6QIav2Sqe5Ibml+r
8d6suC4oXOyKtiIVwMqVdIzzHPrH0v9aHNazYwDDaBR719tEaN1/6PNE56QtrgmS
Nh1gE+fHQI71HLyg0kOnUQ==
`protect END_PROTECTED