-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
RkrBRB+2jVPxqLizLjKT8pSMqA5etswuu4wnnAIjedL1ttETo2L4aCBHNi+iXvjq
A49lNHy0CgXFDJAkDPnhDnqBGFuLhU23TOgiL+cG5Jbdzs1skTa9saE3YlFEe1xB
L9+aUp8LQuaRF9f+xIChlyp5pESZ4LJLqLjgDBwQgjo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 30000)
`protect data_block
ai1gaPGqbPEqfa9OujHK4UmCylMpgGNWEDEygxinz0xyDJ2dgUjbUR0iDG+yE/qY
BfnyQ8Dgn9xNehdJb/PnxK1CyV6KBNAYmV/mVeIBqPify4a9yWBwroNNXuR5L6KH
CCq6TwWzD5Kt5UCZzrl0RZWUyvyOXJZp2OzLGlglBeLqNyUn9N2BC927hjr+aCY9
LObBLbkpY9axAkA8x89lBjyDhc2ErpYSQ8j/g4afhrPvDNYRJ/p9+X1Tr1Q9r2DG
o2h7mNZ1J1ajODkL6siQKjBU/DRcrY/P3ry3d7J6CqXtfDuc+orSe6mduPOndjva
tKixso5s+++qFfZOCGB0rJk2rFd6CGtoN2u9WqNBAqwSURT1NpKBYJ0M5nL4F9TY
CNyHC9C4pI4cokoVN4i4K9zrFccaJARSXeQ/e9wVtUTauOnuxNeuaANt8KYu77xf
gojpzgIRcE2GT3hpgxvAHHGJJl89+GGOASpFHF2gKfYE7wLo5k/52HYZ7yycIKka
l/XEYmvfmQC8uWQj/3PBC5+lHYdBey2nZqOmFnEMNqeS4BoCdtJMU/tfpz0DtkNj
1nJt/HNzWYx5IKxNUT1ntFTFit17GEKeMgTT/J8+X1OEZkMn4c523xP3moqlDbP7
fw/XlGD8HwwRSDVP0qPBym1i1A8MrUXq6BFuUyqg9z2VGhrAt2Uij98y4VaRw2tr
8OH7XfHJQhZLnOJVz3aZKxEcxWtjMqcdvsgkjCuWBayyRNZt/d7OzKN+fqBF5cTH
vtSFNZgBGe0DixLBlPsdPn970Z7F7xjsKS0E60/hoy4ieMRLz7x7TdecfnxBqgeF
clYbPhPYF7cz1ez06r7UNggDF3eT9bmoHjYtiQe8IfnoCIMjgZvwgfY5YalGNUhw
zRzkfFJvlF/Nu5zMYVDIHdJlmMxNi7GgNzif/klqESXT2MelX5ZA9tXQEeE1lyLL
saOeCvLZeLEeObYg2g508XM0wEXonVjaTKkx6zHplNruRrNoFz3iv82EODbHOwxh
MaYh5nIZh5dSD7tY6GKbC9lLA/pJxS3IfubUGzQsAPK7P9GglwrXTdtiQB/fOk1R
Ksr8GcSwQvwPo8Ol9RDofrGDG+4yvVgnoNlaFMxg7fbPcaAdFzpUnpTCyzCfxsFT
/kV/vxeCWlw3QVlrceL60mmgUdXK7XuD5z4SOSnPjLGxMZn5T5HB2OnYRaTjqKQs
Oxm6wZODtLUAefhlr2PhNGwWlhRxcMigzG6PuGT5ipDP8HsmwoaPzusynQoAM0pW
Sn9amV1Pua/Pzlmjv0x/Zb0fxdeFhPUBj/J+ADzH+yA4tSvDf0q9RLWB+xg8MExE
ZJ7h3FeQKVF4geZNdHZNu4/47OSEOKAkjKnRY6/X7kkPHBgM4cQKBjyFPQbNasKW
lvO5cgTzsWOL9WJcoHkun8quWqjnrZa7ZBviIn9IU/kiqVU9IngEoJg4KqH8mFyH
akyizUG1NFzGX3IhqznZrzygsTNAwMngVaXYVnhiAvz9SLeYhJkpmxtuZxZgzEq9
CRCOAjcs+ct67MbCNws7VLp1mdXtR6F4b/s2T63fcqyBwfwqarCMcoTpu/JAyOPC
2lU+obXgJ8dVBEH27NpFetG0CUhpATKOlOmzGyy0NKGqLKmLq22Rfaw6IqZ6QZtE
r/rergXoJ7YiRi2W6kT61rf+hej8uQa5+Ws3M2EfzPBxWncA+ro3dDx9TDFfim95
MEV/Fo6/8NzCjLShF93TXkopPe7LQz1xWPD/BdYGwjSkDWgck9cVGIeWzPqF+tDs
hexPdR63m/SrTwYR0aPqzJTCvwaCTfCpC8umMSp3tzSismnObwSaIeALj3ej4mMp
ppo7hM3CM6qfp228Ncu+SSbK8zIpUDr/ZuFfaBCljnzdxsOMXDz6aR/nq+Y4O4+D
8v5t6OcPFGhIZLuZLb32BmtNXnz90VKhSMIYtTCrutHY7kO3RZ7RK0eaPSSp20/M
g/JcJwnX8DZIp+LdCyyYel13J/dd/AvzCX3hn5r0ohW+JOkN2mDpXxrLM7gOiWoX
Z1R0gLaF6hM14yggUBozGKMM7uQMm8sF52/GQnBO/zgTmw9rYjb6t9WC4M1brJJa
FUdMkixLvJTBqOpiz+DNbqr4fZRXz6FCO2GHHbA/mES9Q6jowRTtr/Dg7mze4xPw
iqKKYiAbsNYeowYzKqtfVjx8oRhXHgoe6Z7TQQs+5UX98HVFG2hUCLoZ581JWOJm
zlPdx76+pJiU3BfF7FxWRzq0l9JiLSq72AGvbzAV7KvWkiDUL6cO/ei+oh5ZLTNV
X7k1MoJGzBY0X45NDFgujPzHSa1tACt3PBGk5khG2MP1AW7osbC5Un+Xm9KJJzi5
dtsZ0YX8L89Kv6m2tLRq61GNAZ8kx2ERMxk2fYg9p+7fW5gRN3g7Jrb1P596ZnKc
KDjn07Rm+5GWgLJUgP5hAql4lQU7h5qUmqq1I/LVAwoHa7DPw3BN7nd+ROe4aPYt
qVo/17ZX+pe+lR3TWKLUBGzF+HhwpwlRZi+VbQHurgzWN/XxiPTKyCC6T5nbLiWa
84j5Tg1/5kVLgrxlYny0TqfoECPvp9mBDEB8y79NhD+g6E1qc8OcjaHHMTtcK3JV
ZJn5W05KqgFZGKRHHd77L21zbk2J0a5pxTKAyfmRD6BOt9URzBxlXCm09aG8s0yA
JxfPh4T+01yWYSbmJW/iJZLkHlhggrD/9Ki6xlio1ion5YP8KwZJu0lV7kvmMYF1
fB25LJWAN2/NqfDN7fC+BpDVKbX5KI0jfO2+bdpWNvOjlQV5FMrhdSiZCedSL+cP
iXrqnIdJw7+oJSK8v9IpkACXpsXtUIUDyJAs/6s+81oVidn0mUeXXZXk+8yKGCpx
niOlx6kXljjR8dimudb6pz2sjvxqEJOobUW2jb+RDoLtGSD0l44Yr+kcwb9Suj/l
P9VsL13SXk4J8+VsO0E4Seh9aEcTRdQjRdBQvszXLHkzGgn4QkgkkQUbApZiUPR9
KS4h3d5piRb7tqQdzdKMTokR7ldNyLFJg5Zep9KpGFYkI+zpM+xhKTX0gtlyI/VA
UqkpY6qJXPUWzSTCnBZ7iHt3IgKi3iLzN2ty4AhdBNLA65YSzJvS7XI0c253M95q
UGKiX/jd5LuUQSnzLBJpNMu2Esa4HbkJ2GbyR9oEeAMZ8TR+EybZ4pAJcITbIKM1
3rDqUyMoIykjNIsr01uqU0JApdKSNFKPq/3YjJUCYsXKwBq9Y1KarFzVCDe+hx5M
LIiQ9Knyy3atHT3KzxP8JZPdciU+OCKFQLJgJCrofnybDhN0DFymdFDNhSFJw5Od
PG1Rdursprb5+9/iVl0Vezcyv54oiTCmWfjMv5aJPYvEjxQqabEqI4xTyEIAfW31
hOUkR/dAKKMcAb7bNz2bYFOt65Jx0MewqdC7LEbgADfTNLjBz0sRjEdaweLPRWx0
ISFR9QzJAIi6StqfUOQ5yI+flAlL+6jx7+Uv+jMGywxQd6SbBW7mnIZxPn/Nb8wr
h6l+O+l0IOagvLwAQh6WsksoB15eiMqARLpana80noxlvWfU0QsEsagM/LH75B4a
P8R2i+Nb1RKML7DhRWCoMPRcG6chOhs4hz9UK1ruLSFC0bLUnJMTp5t7K3yE1M+S
Abi2a4pi1EFVhTFr59kqQBAWSconVrgLLAahKLYZd0MYfDENhMFIliT+AV8nx7tb
TVDTfctZ8o+Mh0rbHKFDlacFhl+4dcKP6sJ13/L6ONiEYp06Tuxt6SonCizbWjgY
mGpGitq8BCBF2N9NaW7awFlcacxcQ8ifSyJ0z0JgbCdASGh0NwhlVxwHiRyZ/KlG
YE1pCGONqd6cJUOd6C2DNavhljIjXpyc5TLSddA3lH38fKosN5lAOS0educvHh+E
/jIKSrnrwxT5EJ81PmBD8S4Kuks0sYGRiShhYkKW4+44s2N0CF4yHaswx40X4fSi
jmxxBkyzczplLhWwV2T1ZiPILZqiWBc4rHdIoBEojp1ptOUfIyhO/4qgEN/IIKZZ
VRrm+GEL2WiQxy6cN3gPuQxS8FsMCEvfob4qSmFMTYQH1tXVBnYr6T4Lz44MnfI7
jnUTdrNroCkKnO37C5ZYfVswQUHjRMgWAQTsZMyZfI+FccXH4XNNd9o/WvBwqC0F
+XaXbMsJAYtJZddCon1P+82B65juvCBIzzTVTteMMFpQ3NCwCl36Ns84j+5kuLUW
cKqnAV6KrRd+xP7D6HRFSZfotAZaXgDbfE8ks0GBs03+3NKyFizY6SPF+2Ys2vmI
783rV/lelsNcezgAxW9+BOdFfQs59rtxdUWYM9AhjqG+/4hl+ta3BGSYlZmmq3Xt
Rm7UQvUlEXfeLqtVBSLLCJ8sAMhAlR+5xciy7YWJqmdTkRzUIVVUZrq0ff17Wgxr
QoVOb6LdYBUFgCrCU1MbDucHabDPiH2nvMxXSmWbCFhZuuNhSuG1JMm3aC47CcOC
KxzD/OpaFtDH3rWAss5qBTeZ0oaYMjboXS5uiA5GIsTC8k4gEGYyTZPzXW53arLy
N7xwWhvp8/r+4iJB8MhFDgCPcS2Yp1Ndaw2nHnZRczqThjD3W+bD24fvWGjHRtir
pwx/OhcRneV7KsndmyueCNkX0YNfklMWgaFSyyd/bg8Ipw5ukFULEMKh021JfZKY
xrF24aBsLRZNmcHMaDisk2FoTNBTTveIO2NadcgAyayzJaUSQn9mql0Npi/Vidgb
KPX6R1+TRq2Q9Nb99veIkAKt1xOwP+6jXn6rCKO+byn84j4qrVEtAfb2KqufaCN2
HXJ9d9itGZ3y3Gj6j3YiT5jSrxStdvH8EY0lLYY+6i1HeGYUfUbSPjcpGAuxU5p8
qV/3mev/e49UO4ooSU6uYPrQp+cgvpENR2omlhddGzcdMHKR8T9Av0KZg+L/x411
t7wdYNPEhb1ZaL3RFaPIlzppGE52kI3a2DxMjBUZz1wg2qjO4AOhCrIDzZTgEaCR
2nGHtcf1z1OSgnwfE1PNkt2e9jst16KAZt1tdWgxg63XbklxHm+NYphCiRBdQz0a
z8Vnm4lTm0oE+IoXngcgoYrXiVsgtgR1eHuduqQJmLwvRWZhRA6Ty/q5hRd3/EgJ
OunpxtdJi9psqnPc0WGhjzc5UBohvfic9O5yQbDD5sasjE8KzxlkFTTBGKl/cx0F
r0Ga60xWvYNO8dp8nhFSrX/2FhbV72gd9H9mchsOZwAAU9kZpOTCXozmAEYGhfKu
G1WRgNMwupkbpo2PkRNbpVYfEz7HtwmvxHEVy1nm9FCVmiZsShGIXNmc8R5JNdQZ
eb/JxT9XA4DXy6doBt4RVp+MZaqlPRoPrL9fnKOrBk4hrZDSYaA9ba5POPN0Gg+B
HBftvlxk7CXMtuAWCeNzJfCkudzL57Kci9AMuZz5SY6HTTl+lR0OO9z4nho3zoVj
ZAOYm21WEtzdRTWZdqxdNATPEJ45i9c1cjWM05TGkZPSGM78mBQdRW3RSVQc7Mf8
vp7xNgx9aJZV2WnYBQsDxa9Y+/UPM+A1/W9DXo7bvKass+rUDAak9GSDVG66tLsh
6O4JwLzD4wucIyJqIRTb5vNCw0PLPuslp4ht1DwGCrzDj2PTrDRd8rjRV9onGnHI
GP38XQJUsX4fDXAeLk6Xo0aHX8yDw8KQ+UAmedQKA8e5oQv+asBr9pfd7kUeYEaS
EY+YcF8GtJnB7KHBI5MTe7okw+gowEXaM/IvBqWaqQZFtEfXBq6UwosluAeW8uml
5gG2yTYeYY57gSptuNhJ4mTyEvwGGSSdLsptnqDuSpuOqDI20T/j0Haqo71M8lYp
Bq9u6M3naEYhOeu19IbXUtd02uQqu6mI3rh3ekZmT/WeUt3t584brxDbwZjqRJAi
vp530kWV3CLBYN2ogAwTDCPvRwWyX50w1uCND76Z43dN8q4+k+dwu7L+v0XXkV4V
215LsQL3ILUb7A7CTgdEeghQCfcow4kziqWm7KMsDzHW+2dyNvqCLtNUhExRb4lJ
tcMwPwPtW4PjxcrWMkdd7gyOeez6v8lcjvGHT8FZ7KWE5hrOd5wq1L4F/ENGXxv3
ZcFWDwzm/ZXv2IIO9rjJbSH1TgREmYkzuV1svDpJ3WtOIfixV5/or2UXW+ld8Qng
3QKxFH+KY128pBZFN0UJjO2dawizpHpl67+k572Iy1sTfA3cFZ7VGJfViHjZDV7f
3A50iujNltoOKbEUaJY3PMQb8/cedP6SUkfid7JuJH1u0OB/LMD0hd6RvkM2woc6
rKEQZCR99jCtEZW+6QfvU3ebqj8WGR6XoUm4gDlS8hP3ojWo2mz7dvs+0VUTISFQ
kAbqmimpRdV0+L5ugbUSlQatryiIRNLsMUf1fb469/4V7aLXoeGMUnNwuwCOimtQ
RPOzSyYETem3/xB9v8Ty48LUK4PHT7tvwR74nasudeJ2NLSkuCYno+++95KBugrP
rRfJxKUQSx1ie3JJig317TxJdhUWm0RDLWIn6RsPl62UkCnUedaiqT+BswKrkVah
lHxm6+MnWvn8mtmIFZKXEU3Mu7Yx4oiIMMlfb4BxqFnB2uFzFeomvkcRivGWdaX7
zjIzXx/eG7fni/N4nnrlcV/REILaYiRlPZiw9A1gMeH/lZ01M71wEqoXu3faS/eR
k3XWPzNRQoio0WPN0LWjNDnauVWPMHc8jNI54nvdR5SGWFyd5YShF3Xa9f1w0ti0
8ItTNw9559Gs6liLhocWIYBVnbzlqhNaI5LlBrC3MBxHAFRjzm0j4ueGWTg464HI
RPBSALbjI82rdPRlhSmUHZm5MSrxrGsaptCqPWrf2IsxeJHN3GDxLci5n03GMaff
YNd88MH0znBKf+EzPZVlGZcgEN8Y1RYjaOoUtj2IA16ZUOtJhKfAMngxM8vJ1nzK
cdjFkGur55fU5HKAOLWDWWHmPyicnsqC4bUZe2O29mdAe83Wcig+KGwk23ShFp9X
dWHjSizf2fRAuHVFr8BCEzBkj5c6okTobOjE0ugQFSOuSaNEbAI1TLnaexU0IYFI
153NCOVsZTrwGvACpK/HiGTC+0j07EpiFoXdjszTqIwMvZkDv4gKbA4JXotfpHEA
Zt2jHIbb4aJDKEN+NtIL1RhY+7ykU3aXijGyZfofgk5fT2bG5CZVKreeCzarxnQn
t/9C97VXGz7jj5DzkPHs2R/0aKXvL0ZlhxJSs2ayz95sIWAl7EPkrH/H/kACCHli
+pZx1jczKpS2C9ZaDTa2drpAUOwiID4Tul+M5T8mxcLxWp/QCXISl19YukNRJpDT
0s0L6y3EBiVb51rvD2LBEaWmxh9+XVnt3mcRtGO58KysuTfGPMx3zUzg7fAMX498
7vRkDiheowujPjAZ6AOOOJOPCKivqeHAmvKKVZnc7b7rAiiiT1pMoll4H2IevEJI
VHEdHBKjGGgc6mDqyEgOLd84aBwYl0BCGZ3cXbLMn277BTjHR0rpuErqUaBBDMKo
9DqcRnZdQetm3tmtF5xxUSMTU4AHHcOsHO3uefGDcxyLsRgqgAat6mGPMurMWqY8
F1OnXwYMqsCeCadyK8f9hcs/rs5+IWYE159GU/iZtcbUf/Q9dm2EJ+HESp2hqnf7
TTZTU3Fupz0SygGyPwwWUiCNuJZLUopNdrH4Tsd8qOcLJ+9SyQZZ8osbSFqe2hAV
xUK5jhy7tUsef17vhDr67WfVKxDIvDjoJNRZqmCkqb/lG/isUoAim2gMigIspWCZ
0I8jqDgkoqz/cy7bjp3SjexLhRzTRgGKdXfyG8qeF21W3Lr3RonKSx+ikPAPI0TM
m+1zDIPC2nZRpNV42XWx9jrqr0aO2+35v1EsOfcNX+HzOa9BoWHlx/MCaD0/hL4p
5qx62vf/pe+nF1fXnLem0hdIbDL+nKlZt8UYmMLDjWOn1QzAK4Sr0fxeHNAN2bdY
U2V/EQK5uecXSWx5G8XEbb+5JjW5HphpCqlhaqUYY0mcQK6uGwR3k6iP5dA4HWTX
MgL8+k7k1nvpIGxFbFhQ5DTyGNUV9GzqeKm+MRt2v9OuAi+w/ptLb8GSTDV4O+ie
4lc4O9KEemShLdOSCLLL9JzpTlaSChm8E+IgucOsSq5KUKbpyKJGSsty2Bp/2zyp
fL6vS7ur3RKbFReLNnmdN/ua2t09S5GRflcr6YD6Ady9BTGXVsHC2IS1TiFrsoPd
Xwx9RikNGFxNRDGiOz91izhYY//bicG+/TAsTKeNg4yRGjOL6k06vIUXFpDIz/bm
bqOlzf2rV/FrtdRQSlDOKm+Lg091fl5w8Eqch8LOU3ox2HXnhX0ZIMNIJIfxbRPn
6UgZ3shn0nNU81ZBj43Pu8QB/EI+PUnKDGq6b+XYT2oFWElnCxFXe4p0vD0BbMO0
EHjnTrsg8ysS9jDcnTZZyC1jqmzjvJwQKfWDQC87909oE3lXzBE/ttFhieVgkHc3
Ozdogevo6a5rxWLdczQRnwVy12jk/J53JcBjZkptL5/Cyd97h54jDcm4q0GgTRT2
mQMHHeLrIrkrbaRQlISHJCCY5pl87zMz1Eq+1BMUq205s84gZpHpwRfB6Nx3e9BE
dB1Mjc60/r4KUFfjEiHP7w8ocTznBf/TZIWNyj8RUgAOWcPiuUZl7WeB8x8LH+4B
vDg4e0aDlO9AVwJOc36BB5Af7q80vOuAw1dt+z9zkDLc4BMk6ijEow3rbGKaigWk
bJE58/XE87PcfEjNSRrksRLiz0KIw5k7r0azC2eumI0HVXbCJ3EMf5Ht27JYvSDv
ZNT5PLXRa+mAtzb8AlK2t2SRXKfj6PgnQdWmK8dryJ8gxgrJoEoqlSvSVnBhHRsT
bhyX9Fjy9lbBhbUOoZJuXGl3H+wvaW2CDZba00KRJ3XBbSFJ8UYyUPHfAeMudWPV
CpC+n2ZoQXNVgNS4164U6EPR1eZ3d7KJ9BGz/JxPGvfGffULmRZFwHrvjKlaO7WP
KRA9wOIP+cANtregNcBNRoC77X2xDfEB6RfCI6y3oTKLDf6nGBsknFJSAEE5O+8V
cYHei7x6ivSKCmUuqxSgSnmgld7HLp599DMZQ6bH0N2G/gKrWwxzSuY0PcXOKSfI
Q2RcYWiaEXbZQPGiSb2XruyLeNKjAvw+Zm0G25gfGZDAKF2UcoxUN6LRxpxUq0k0
+HId6UYCxi9XCByuM2lLIVyJVWZLqQVPd0nOdW52TTfWM8mRpDtPGUUaejc2QFcl
RozU2C1IpTYAeUr3uA4MjMKw/2bSbWl1AgcdGjqp0Hs8dPX8yQInWshZEVkKdw81
kaL0AN0sRgKjRHeSeXypuKpI7qHJm/h2AADmaz2PkK3ApWZL7v6Q3WCA0w+WIJ0O
UETqXHJRZuhSDpTywYPLHWFoYTd49aJXyMyo9aob1kjk4wU/3yQqVnoOpvW8sjYV
PQrx049C0Y0LRrG31Wf9IlUluF7G0BZcZkz3AxrxKr9jGCp7s/ORmeMsfiKTx5j4
PlqBkUN8H0TSxto4szGr1Xm4Nt2WU7tpbr4VeM3M2GVdXqHP5xZ0K04OTpO8XncX
+mAMJsWIMMnXZKKqW48JwX3i0NrYGaDZYBwDc/ca7MGlOPN+WIrMPG2SEV5ENbHW
5T6m9wWN3OoGBeugVPT38TtaDb/0QmQDjum+JioPvEL8O13vGNqwuZ40PvLB5Mai
BPjl/rfr0Us7L9ZHNSD9meK5bOLNNqL93ayi/T+EUcHVnsyDpDk1I6VG6PASVdSg
vJxY8pJG+mI4ZfJUlEc9skP7GMAJdpBzxfk7ycRTOz+nWcDGATnd9YfVr/3QEtye
W1zVy11HOCfu7btqk5xzr4aHzZ5gBJ+xkxhkS7q0XVFW4QQwVD2pcwztpCpks2lI
RaMOoSbYftLzsGR6uMtFkp4wd3qUurBlP8pFf3Ub/eKJYoB1udB2wd6JecTOXnYm
djqUJLgPz57p/L0IrgdOH5VLcwBr0aoBrB2mZywea6dFfKpHIjeLehz+x8RKgmMh
5MFxviSrzkU70t+o+2CnmdNvczy1PiYZ1IsbRGSUCgEF7aRzqwHaIyqyTBgyq66d
Osb96ugpBbStghsEWAcPw6E3Wbf/XL64H4DcLrm45zfx+HxLgqnqEWDkglfOY+C4
etNuX3zCD7tB4k8YNxHlkIiCquLXwjkYIH31zkDPJR8ST9bMnOaAme//t7zQ/FDD
3Kvbshgb32cqUm5PILYaU/TG6Ux4gUe9rFNLiB7aKxxcU+FpRhLsnXtIG/Tbu94x
Fq5x/PuL1AE7aKESc+iwy4ZtphfwVaXk4KfYWwZV930b7d0MUGnC9z3UzocmFH8e
EjbASS9e5Wlkuv95QWg3XO0rwehppbId1SPDJeqQ9e42PBt2NJXgw+OCnQMV5hII
iTvPRC+cLxQwtZIXwKl2idy6soIsJV4jvmi3efc+O1mkH42Gw5TSlqfVTmJuIOVK
HzXpRBVBzw9jB4kngd4w5dcQjWEyJU7FSuSKH5zFMbknyBuEssYgx2ALwF41h9tG
hr+tYCF7YcVdzobr6kxT6jF5VkqOauWutpONJK5vomu2zur/GIczMMgaTETVgAim
XsuzkG4JrfX0lsvlrdFqn0bMFmzMlG6ZEL9YDu0iJSIFX+I4E/JzQhm1rz0G//LX
oqC70I2tRIQ49Gbz7WxLRsuHmNaspnlLjpIyKarxywnnioFe4D7Kc4u34bJNV1rK
7yvbFWtOg7Cq00H/QQxzNs2nuSdVOgVIopZvG0MCjKVORzv1doG75w8LdGx6S3t2
1XnqATwY9FKKgiP9cTIFjhkcZ4yA3M3M1U0NLPLl+7SK/jsTICnOZtHcJw7PaYfJ
ZwJvSw2L6g1YbEfbkeUw5LpG7FeNAucJat7eRw5Urc4EzGE4o5TAaa2WAa79aLfx
3re+QZ9wfoNjbgNvdJUle5jH4aSok7LQ5zMGPZAoDV0I+FwU9hsi9piG2ZnuqPEN
r6D/gQmx53VkG1rkVffgThhnXcARwOlmxNqi3sXVs30k9iqy39vqQZU3Tz3ktn4g
t2Khs9e4/K/Gr2SdfpF7aFJjjiq+TZQCYCx9I1/c7RfwWyhqvBG7V9+lQcb1UVtb
gt2XmWD14U1hQb/MnlT2JBfnq3LSMivWraD36l+9e9g4/JECILWIDN9tVdpjlq7Y
+4pSfEJzB6JiAJckm97xRWSjBHL2h6s76qC17g9TG9+ExU065j7N5+0Y36AmUJ6D
0VeSAdr1dTQz03R1bGXr4+2vpTNQK0y137fsHx4TQo3TqDNYjsPb5bXE/bKHRPLc
1knX11ypANAatVWNN0WVtC2Kml1nIoQVdwCJKcDNFBGJ9PAsMBdwr981zlbNOfT5
o/vnAQLhqk8iLRRBPdfj3hwqytyNKbWNKGEVHFGzSx27TDh/gDxX6GXyuywS7qpK
hnwJddGhS8E+nsFzZJHK5CGkv9yJV0qqK7E4CPGNUg5pe12tLpl4/hby42M6Iq+0
m03d/YU1n3MxAHshhNh0Av194xvnDutUECQsDU5KHv1OUdL25e7krbGQ9tT2t0oj
hl49TMFG1F2daC/yQaKaKXKXV01C4KPyVw9JcWjfkxJkP0Y5Hnog+dqBjjC0XnM4
8q1y70hC5bj4CYZO90AveuUdLPhOhd+YppM6Si0xFRY1bD5oLYfv78JIYKXGIwy2
6SnPUel+QfI+5CpCSxO5BtGE1Q/D84Ak/Z+uGuiOnE4wruhj9fJGWbvSxz5kLj+3
P/L+ebKNsIWO47RHwSwwtnBExLCJjW04aINPnpAm7WZv4K+O96QARU9OvEVDgLyt
o/Y88RA/5nPLehTbfXT9VJJETBkR+spaWp5hQFhG0V/CrSzpBycBWlSSm/YD1yWf
x3IOe68Vby0+WGWSb33eUjQa7Oo2u370Sg8SBhCgBrSs5hZK5ndcf5F3RiGv8+//
L0D5+8Db0eMavuc6Y75xXOU2VaQeMcoxaf+Kvdu7kCXqSyHwus6I3psWeyxJAlEL
UnCXY3b6yzbEIx8HPTeThYWScNfku3A7IjnyULEPVTUwEW0dkgstxlaXUAcqAIrK
Z0KKgt/n4EuFbww62dBvLSuWB+Jy6tZBLwMXfcPIOzEJMqzLaeczEJnclm/NnXZc
wHCks59Mw6i+BNMmhDVk597kXP134vYl1yl9IMqPyLJBfYtEwDGcoHOEJNVhP+8b
jcFJok1e9mxC6GcIGjfOq7iI2v9Z23qKXz2pH7b0GXJhJz+Qlvq/zK6LXz3tKBdC
r5Xw4VEI/FJRoGMTyP3PBJwjN8gwnNxB6X2/pqqgPMCiumKv/CbGNmNi67GOMKB3
JFwaCeRWTaoVMo411L7FDlcGoVLXf9y0Vz+0VvaokTiq1aSzZeyGgamd2VmyLhOr
KPCLToig9wmO6DUzy5iA7QHJ/c+Eb4PxFcIthR94bSE54Lr5shIaDBN+pHSDY6By
jTQpTSDKd+rw+lJ9CQsDcfqcvgb677SX72Ro417DqfDK2qOuzoyaSLAiv43yUMxN
fhBV0PFd4T08F6Oy1+ohiEX0gxRNRxt5vQMNwBlzSyA8iRN/M6i1s1UBKWxD1icz
CIh92sHsB+dn50yP1we/NyVwN4VfWo890qhyO875zDFgdK1WBJYF08HsONVUteOm
3ML+BJIMwN6mZWAsgj/zVn8BtA9Pr0fvO3llT6SrqD+HmV+rEV1WH2YksxA25Zzh
o2SgPCe4YI1mzWhDZ38HGdXBXJDXP3XriArQsGzO7Kw1asjYZIEyoXWttjIQBGmS
yx83QEfCxuoYlms8EMp3EeOfdRnujkJdsUeKYLUxcnFkJJhQ48O/kNuWVnxKf10h
Elc/MkmhqTrbr7SUpsOCK+MYaziPYCPCaVhVK7eE7utO0nElYkyvCSaxz7i11g+r
CfqRrwchfexg9iNoO6i/mmYG2kzcUU9G3+MJy3T5KC3ARUktRwwInCrdRXRjUm8S
m2u7QEqQUeD6qf+xGGpr7vJOsT3Ok+f87HNvQfPlqIBdoyzspn/udi+uOqCxSI1o
xenH2Drk7vtob51sThlJ8vrofmVMkhQ1H65btA9jNtVgFySd+gansyfCzj3Tu8q4
CSO8mSzcJOEXiohSBRYqTGNzrAyhLvlW5SIPLpAKJhRoSXB/lLotZh8T2+joYX6c
WM56TpIc/tXp/Ndzh9FLiymBy5q8HYhFb65EFBIMLlsd4n24+h8Wty+eFHoqFAnD
WuZ6ZSDg+1GwYNvgoaOpTfyp4f1FwVY2qBqqjBHSvSBSy5C9wkDpxZ5ZBmhxW7Yj
u5zOlgesnSC6qU8XpwXwJj5RwYEgZH1LVNg8CXc8Db9vyoTiJTIpP5/bFnIf4fvX
QFTh7Yl1qEyZQsWBe0ZVOJGtdpCTmhqaad76rxRnLdlVLB5uFFEZbIN2OnYVKlsP
wMXPEcaniOfaFfpV7LasLk1TGcsnqoUt8hl1pjSmlm9OL+7t5VO+lh3xSoQAhafb
M9VHxaeDh8iYTOza7EwGTZViTt/Xxma/hyaV+42MNyzTDr2emrGxBo4U8a/4cjT1
qe7OXyUlT2vovOypmNneqlxOh2DvT/F4FJNTA7YFFlL4tFjVaCAMLx3QBVcBZlPJ
y5qHGksMx48fJ16lhkfqqPPbIGzwZoRxvWy5puPMBo11VJqma28t7EMPZLkY6LxB
zEf1Wv+sRKvD+1oQRavcvUKimbMGA/waSqk3MuojXco2iagCF+QRshd3l16aGYGF
WbYIoOpiVdhHWtmfdRQL6EsML6Ey5QAUFYjQLOxFeUxhVLA/D5onKL0WuVqjoDdb
NgSIFIV8S85E0gWWnlg8ZKC8Y/jL3iGN8/MttvkGkkMSvZEpRmpLyksAYg3MWggi
InFu3vJ6XWGuGzY4JM1GMiZpFRmfrH9SynSn2dz8SsS6IjL0KfjudmDgfrWhXFRB
SGiECn21J9tNYTan6lB7p4IO2aMB1srao/3h67dTzlXGbBc6s82hLXCny2jSEsLs
y1ffPLhGJUWhrk9Y19mRznIUr5GjjAaufPyGXOH7sSRW9D+uFV+PjIy6GBvPiHb3
QK9mu3XEnFdgADBu1H82ZM87HAEA5BXagfpccITgvtcwAP+7sG6ra3fchRbWJmZN
PZdGU4/lRqOgXkGKXBCN5JfHkAqSbzakyAhtVHntTl3ZgRdoucqZ6f964FG0gTjU
qe6SJQfFjaW2EH1CwBSu3PWfkSmKKmAISD5LuwLS35yA7tDv5FuauO+WCuBsL6Xw
uHhrqotyUcHtASy4D8vG/uzeGNhDuRAbeiOonKmpMkwhu97fROR/v9m2fCNI0xqQ
AHqCPyYYoJWJJHyDP/UmiARKKLXHctwbe0MBolRCRbRuD3m4NHoGTeEOQE6Ht9ZG
o1HYfJj9MSGjxT3FIHI4WVnknMNNkcbLkod7+k06d51Nw9UJv/+GZm8YRnP5D7WV
I76VhsWK+0u+RLwvqUiEHj51fCFm2MRv+KXrK2T2i6K17X7dCbcrp+1KBcZb2zQE
Uht7bCH8d7+gEOV87dNbUz6Si4Fm3vkD2tZc8zAgjaGmp2izZ4rr4jyvvLB9Bte+
UEkRg259Fjp/Me10h5W55es7m05qE4QrwdukscRNpDkHiNPBPooF2VDLjahEEalB
vM3Jkd4V86LDK/Ube9THQkzuoxVD5BijfXsT23QalZrES9qQIttqYjAs6gMPx1y+
qCUAFGfb1DWLtKL8I93Ff11HgQRhZGP7ZDJTBds+vDqVrX8MM+69q2dl7m+9YIDN
Mi5y8FfiWqKyYhxU8hC7nd6aDDPiBiktBTkuh70TuDU9BzAc0PpqOlKFc38Gyboz
vAwGriRSudKz3vKCuEq8uJNpuqMLTeucl9ToTZaPj7kyLgCotEcTQ6OFPfVnv5XQ
XWr203LC3dvRs+N7saYcU24cBvPLDs8ix0jC/Rjueuv8xjRsVF1ZdZcDUWinbbgc
nqL1/8Io6K5Qowj/kTOxLOuVT1sEQFU6uPwh+RjmcS4UR0XYcI5EncJijfNSlEbM
KV7FMaw7Q5GnZhyzJFz4VCgnpwNXuiyVBG7hvXKxavMvvnWdoxk2YM9beuY1P+RE
OTy/RIqhGb9AiF2tG/pbscR7q3SzVAA7aZkWsZpSrxrgtM+IvAwIYEpkdrdU/90n
JmxRHMM/moLld8vFImtsMeMleYkAwiDX+jcyM7lWE4Gqcp3paC+A5zJDAZ0s/0VR
KfPZt2gkrhzS7syKq9xKfTBkfMBzrPS3TM2cgl5PAYBBIwZhgAwYCntGWhEShPdg
ycH/H4Z1tVbld3QCsTs9KX7H+tO+C3Ge6WMpsSGZhefMIJmZkidaY1XvBcqgqfEM
UNKVtkwXCNj/7ziD0k9Zo21aACQxx/745yaelKl9kq5mLugLddgliRZmpQtscWRX
sqxKKFbw+6UJAgX77+ysTTTcWPFSoGQm+vtzlHyVgARAEepoXYYiT2axIe1u8GoR
igU5ZPXZr+DAVNvdIYkQnw0Qlm2qZNi99w+yfs+H4SRahAxBH77BFJ33F2YsRscW
Yb4Ea0X43nXQaSTvT2jaPLekvdoXUHrHBb4ux5RvSguAi3zp5MqAIJYMdZZjJR65
Ix5L354dM6eTbE1liWKXIM1YUKmaMymd7R3bTqlCKtFnXtBDydge92jGoEUy2h/q
jpIlAHik1y4rbRm1OHgHnjmlwriG/uMA7bTjGXcXBOIEWhXzWgl9rIC+ZtGwe7vm
dEXRZyojF6INUdRHRt5PCe3GtnKsFH5M5/d2RrqGpTcbHcxVtGpbG6OhVsPWwEOk
NDysUs3GBUubsmNndBoaKM271b8eRvP723B0LxmHFg8nHYAEhVQoePRsb6/2c6Ku
7yzJFXdE20WD9bilXzJCdkm1t3vFUI3y3HWUz9WKQr7LJLSa/yDj8753F0L/4GK4
QnFwT08p+8EGZkoklMIU4GUCHRDjwr9baykAFF//eSvaVDHN5GTOUr8hihZGFnhN
9GrrUe4RoyY1lMUYhwcQKax2NYOak+vUmCxC5horXNobHsiK6C3DQsO3t3e3gSlH
wRL4iAD3aXpueOSbaJ0EVqR34QO7l1+okYjzRjsldPedVoNnOy+shQWB2uKAO6Am
nfCE7e3k2CMgjF52oanpep0tTfGXgZLq7wOg+BJBwXc8aQA7oFw0l3/MwnSN2/oi
/NO2K/KAIz9eoSjTTlL+aMoRau3e0szwZ2M+g7kfEYqnC505navNhTePGEMyjhpp
Mh4Cl8KlOKu1l+2EJrijWbf8wQH5Wx7P/uPU1/MOuEE+0PaqapYWj9c3PMQ9aIOn
xtc2MIJm2S3gaU5c+YHpsWqZeenwa5Yp+uapPiqrU6AigmKt5wBExP9TIxwYbMcf
0xBZ5zbhy4+0RoTrsfvtFilkBQlEjGKCHE3Tc2INOWjrf1k9eskXTbnTfuBg/+c4
jm9YkyIz0AOFv0zwpSS94HYKsd/QDQ3Up9pcciYwRzMIhBQiMuTAPPpwjwXoqSS1
owuNnRPN41nGepnKpdzhG+DGWQ/EaeNZmNr5ESjx/TfIpynLtZBYV6uNyBhG1sT+
cyk9mT+H3IJskgMZcm7TLbLYiRv9vWwJEzZCu5bDeY605TszYcHt8mxEqaa3mjcl
mU6Yq1GJiefk+/aosUoztSMoufBqRztPPx4YdnqdDKgYe6DHaA0uOIIb3Kx4S9dD
RNRxWwZxQrTVu0ocp1Q3LtJO4w9Bnw+wF9CH8dy17p15XArLJDQv0nShIhd0WIgl
NXz7qthGdnvlxf54IoYBIocTsR9xlXr/E03eRvkk+weaUEUbmSWaAVVXNjEJcsLk
15FN0rV6h80icdxbcado/mgW/XS/EU9MIdAoP3jhaRy7BSJR2GdL2DKqPz+F83fu
NItgc23aslTy2N29v6Poc3rwPq0OKtfH9wPOIahi6lkcYjLPi52FAnG5xo34BIqe
F1DpxKcxFzuO6fwgswKWM53OG9kwiDpPLgAQfY85Y7eLQhN04Jzr7TTnokVxT3NZ
tX2NsGZCc1RGRX2y/8wcqPNG6NcLLhcJ63hw9lmAWQV44umbF/qfWqZy58KtjcLR
ekBnaXCsCEIm5JZLmJNvYfvXm9+zg8BsB2TZsCEGZmleD3tMxC+XdYc3+hR5MTXy
9EMryd17qXzofq+nGNk+qQLhmppVVevuZLVLHf7QTGSGBuhB0HucCuYff+k/giVM
A726xqxfDF43I3yBMRzn/QjdJw/vrEfwz1thPYjcusjZRYUxFosiqHhrW1RBFB1v
4hv7O94YN5L8TO6YafIYeZvPPtdgY84AX/RFuvmpzhfUwNuLpTJ0s9v3K3BhIF62
WCIZKO0t9u4NMxlMBRnobVuRBc1lnY910fLZO2IkMuujuMAmN/yY3qs6dIGJoiAZ
uMZD1ayrNtXCDhXfC2YAmZL2dX1sP5tskjFsV+AsyElDXz8mJuS2xke1YONeuK3x
rSVvllvaKT43j7QQXFwapfWR4OBrCewlyZbLmSCvjz6rfeMZVSCxggHCcW830K9d
UK59KCDOz4dsZnc1aCF7rjXdOp2Hs8ZnFdLPWrj+h9eYZONoboztqsjYKRaJNS2p
p48ShLUgZNX/r10zpPnefUUJSOwi5srQxOITIh2gIOw8Snaed0uU131n7wtcaIjI
xM+qouH0n/oUzTIVdD0fK1PlWyCDrlAeAy4h5TLhQT1XW47y20pqt1hrc8u33SWQ
xJKlPtF+rM1ABHBNU59bL4sOBoUsdUVCB2GXilNMXL3CsdyOXY3kaWEb9h7cvNHv
UWbWKy8GOzi7DAH3QBkwuIXAsICllr+4puh6z89AuLHv+5HTnE5AQEfZnsdZrQ/S
3xTuPoI4Z8dGkAuvQNnUoPOOSeLEH6FiV7Ep5emb36ITAkwLQv5tW8mJUbVdrMrc
Wvb2r8PzicgGlBG3YR/cfEnEM/mDoWn2IAwRRHCc8lqYF4D/97eCaCcBDU0vRucy
G+/6FiVhKvfYwmET9oc0N+mpZErRNQ/chV8is9BIwP/0sVnyKlVxdYybSQOW+W1X
B8QoDAOqrEKa6F6yjTNycIqPxzwEZ8koz/L7VgZzkqE9P8vKHYd1Lzi/PtmLjqxD
YHovUfDjExUDjKsWI5nPWjtAlveaG6wnyACPXSQ1AuWWS8u8fSATD9aB32LClpSD
xC5F02BQtcilyKCFNyh6IWFiiK5YnHjs6e4IVCE5/TKMWNeoAft/zLAbRI2tNyJ7
MgVXADP1hyPk/JuFQZB/JggKSejavIBylkI+8i79crzj2tmljQq0bLWiQcfYmh94
a7ugtmw8SX+YYdWqHGQ/vpPNIHSOVEyB2w9w7aHdOoNEDfyGeLoSTnF6g9o4Z95G
ERDrQsbljRuYnubNIDzsCTKnT2hGWjDFyhuK2piHKM0AD+dD4fvcz2aKytwaQPu4
EvY7+qCYG1mr2MsKDbcd9T/cKEu/ySjCBDv8SUGXZa5SYjv4DPWJzzzP9zJu3O4e
DhTFeyYAFe7p7ebf84npWc6Bg4VyUkcNVkCEivllgVly76eunSAIKNEXrGsOnqP5
M5UQ33I1JFf9nPwzVXvRxfOhvWSxDVBHBXynRlWgPmifa2+a1D/r/JoKNtLUernU
kytj8Pp6wgM2EqJUzhDs/ptB9Kf7GMvTpIb/f0CikpJWCIcI+MPIehrfWB5xDFHz
4hrWVDPBiehXA2jea0/iLwru6zxxTS8ye6KhPcwm6GUfASd2PmK+C/6xreJTbqBj
cEWXyxLixj1oaJjC0QUDCJi/H65z548JuTLIr58OAG+UGn2lb3XtVAUo1ZJlsr2s
/JtY3fMwdyjKlODhFTWlL36OZVwycI5hd9b4UrpXA+zusDCPxOv+SKd+KOSrmh9S
NncM/ZZVo5HTKZJJPH9mfeC429bDoDJwf+8CdUyJ/PWX8+JHCi9JEVR+fvuUYNMW
vWD5aG/kRqMDkL9k/oB20MVK4EZlXexEl8RrG/JteLnHsffqy6RESk8C0TyXbRwT
xrGIYj1jsqQp5ertqHT/blSpYqdaihq7ewovQnvcOZ/b7LS8p35yIEogAHZC2tVz
oJntxScvFDk5Lz7yjvexMgZJKIEEVKhYZcjxtVrBMpH4I30jYWWKJgJCuKLHKXcR
mXjhUBjWwT2xLct7e68l1HSsBH4MSuHHfkPWAiv64PGG7iiCvQjX1GnQmZKyaaOk
+IV3OTcV+7l8R5Iglktdn2bV3/vHw5HU/W6E41x1FJ2XlDzk2uLyMzd+RE5l4nxo
zjudsIvnCGF78Nj3TldBfS/WpdcnH7+Me3dhAvmnV4gSuOtDj8q/ExbDdFoxFeTr
Wr5Vspfdr6Q+ysVtUZhzCz1niYL+Xh70AXNNJtFa831050/rInC5T/wcBgzu6c0F
2wKeVqAIvrQkOnS6zJpdCxsiCy1xJDUbPzWhbpC8sHf55gYxh80NvZpKS9WkWFCO
bqfIpQrlgp7NsOAKZpcbOn0DWGY6pjwWIs1Zd1TUWK9pqLPTTa+pql/+baFrfx6n
YniW7c53IYp66nfMlpBS376wgiQ7QQve3DNGPZ1RM82a4ZHODwz9Z0oeBYS2youi
vAuZ8bEsYnuBPodH5DrdkmZKbb20PKm9K7ZjM2XwlskTnQS8B+mdZxKc3pLoyBNN
cfaPK9UaXIz4qQFjGkIubYd719TScHf5h4/MxjepxjGaEMsG8ey10YUapbmtXu2C
XLsCR1WtI0NBvv/Oe6Pls/O/+os7ny/8SNarZR35wFcoEn4DBi7DWKFOS5HrvMNH
u70IVZCXrKTiLhktZH5qk2KBPmzb8gLnLu7qKFKfR7dk9aYcHlJu+rBQeIkMxtTK
97IkVUhkz6vPYpMzvF34Z7XPH0peNA7NLwJWHO/iMSqljrkhNa++MguAnQgX5j2S
coYQ0egbQ/3UbKSBo4gBH5oaM//ZrAKSUZOVGVYK6At+oPuF8QQTgmG/LEcoRNHF
hF9hC6+/MrcbbRailluMe4jcEN2as6HxGqJ3O0CqP61s/JVQufxCVeryFdxswCe3
XcOO+8AC1lxOClDRKxO5KYYHEui02VM/MvL8vtMolO9L+agZf+oje0TZTeKfPuZX
hZZld57+q0nqfmRXKoyCrTyav/j4OeO/Z1mgxB5mM15Ksqp9WAtLdyDKlhN9MxUh
5jTNqpGHkhWhDiV+t49bgWyLRhAahhXtOoexgM3T83+JD+wr0qMx66A8DhiqP/Tl
9TzF0/Zu3gzFp0ij4pCVuRsR23yGTeQpoX8IBid4FPpIwLkJk3L7F5NGzyPh9wRn
SEy1FAn7/h8hEcyiSxGI99lsarprYjnBB5MC6O9sl8LCGftJaiI9+lylWieRkJW8
2I1wGh7x8/XGfLMBRhAgTTRER4udFNv/y0WnEZxJqwYwdgc2D9n7XBfm72t2olrd
bXHE9oLSrc0Iyf+of62LkxpLmYT3/rhCzkKD8zVDSXOr/AXoduli9vDc69hpfFqd
P1g/U0w7tzJTk8wD4X6Fp+0IAX+vPZHzaUJGb7Nv6SgKFxJgTwgYe3qdmo54C8VN
g9UtZaigwRJW2+x9qwqkLDXsUsp760jXxze/8THFSNcjhbu1vWM6Hsco2siNZiX9
ePgpnpbYPtIqZHKtsiBYXMILL61PI0ZX+7DTL4UefA5lOogjvLGAEDsHrJHiWctH
cuPpFcy70Fu9aPmqSaHj2gxaP7d84/ZQmjMe20Y0PcDnDAaM5+Ste4+ZMBs7kmdR
hVNPAMjhGaxZvfWxZ9X0MCvfae8PiQH0EZRDLB3Hl7ahXT+J9nBXsD+lLHVZAovZ
Tda6+6dUTZLTdEEY+wcrC6syixYH00pu2b8xfetBhUFQWStArccoboFtbp8veWEX
w1lkiOC8+IZPuD5VOgzNtOsQ9K3qS9sBXAJslsd2BcLoHNs17HK/ni/lSMS+nLZ9
WpKKK3OKSKCGpYhL2YMKUjn9gS+UMoU+ED9fZpZZU4RlNzStoTXpz48dv2u8WGPH
MQU5b3CAtf4hk13I+Q3PbubMfkip9zf+5o1itaa7Q5/DJZUPwAY3CGxCduDp8SAl
Xx5vRBXzwQHUHmHgytNY28jnRwfoWDIC7pluNniUKCPFtwgqsOOoVLt26Tag3VvB
YM20AkbX+fO9sz9rKvbAt0jZ9z3Z1nX2pp3GJ99SFwEXKbsnbnXbZetn9HBLctiw
qP0D6yegu9eYE0DZ9w/z9yaDxtuKUnl1UGbcYy3brsr/s0jZzi7H6XbRdzAQjIoH
A4v958wvTsOZDJXPluqPA20ev2Av9LzzliYJE0tRgexWQX1NcRC/vQqtw/3z1yX3
/jfDq9KqNq4UHGbgtDBbPpc5T6MaIkLLHX7u7+VFkaDVOLFAvKbBaXYIAo0XKbJL
OOF4ywhWRJ0f6T7cRZD7YTP5IQ9wvm3ucnQ1f2vJkzRX3Fy2sv6oZqjB1+v0drup
kk3U1OADMlLjoiH1ivdKDBMTmcLIkJsDMlt6yJkX0wLwX67gfGf/teSjxoMH5yCJ
Xio+LktACIMdELST2EvFTTEZL/Uv00P7DWt3euX51DVqVpVxc2Erh1teA98BbQPK
E3+PGPkSTntqHY+KNqUTT8BPicydEULCpl8lf1S3lxUcOrkyYPy4bU77VOtW5fD6
QPxw0RNeseokNSN9OpQ9aAJO6C2Ol7yCd+1QhJR9UmxfzywE9hZ4Rp4iB8RKU4Vs
/WkpRMRC9y06LNUZHdV8S8rlf7keP9Ea6kcdd1Tv1F02LMvnMY6hiLD6yd1AszXu
l1ViKVrpumSVBhxL1GrtO6oYDPFlzp/HRJz0n+Ck2qJ5Ebc+l9sIinyZQ/2SCxFE
RoKlrmGs7xm7NDPPm8RN8vpZi8IlRQEQjJl8iS5NvTuNRxfXBBni6nvhcDPMCmD7
mIFEnVdO8jB2DUmDffMh+2AW+DGu5FfjhFxYVergSbE8G24IvCg5vsW5x+/vg7OY
zcirWgz5+zpHSZTnyrH/kY6yyIfkZxF1TQCnIqUBjVOVvzSTfGZtsfz7gcjFaImo
BFhJsUqDRAomyYm/sRYEYFFhWcuFduS9bbEtUKYZFe1xIiKIYBb6UkjN5QYZHv5E
Kkj5ut5u+6HV43yLbbdBCx524O4eBAv0IKCGkmrp9WA/MRx47dg7EMuoYYBP4r5+
tL6QKrqIt90nmjyso+upNOJEP+oOzPaJ4b+NfjSeLSBwAslVyj9KCQE+lFU/kEip
M3djE9wt9zOknsDxQSwA+0xKHaodDFk9VV0cgGwmDdpmuPwotwdV6tLv3eaLNidz
0JwhZBSCkyk7WoeAoBaD3yeU7lIF8LNPCVWoI+XpnbihK6JvZjDNVGtQC2jirvSb
aaoWjaQZn52ckSBlEwWwnVzKtehgYsVKWgh8yC9oeHKXLuP98zVYR830PzIZP6ym
FivCYsykLSHnt4ZJ/M90h1w/z/dQXiZvSQ0YvBLDApYTtSqy7HEq4h4HkfRYOgne
XAfOsXHg7Cin4CzJL+jRx4QHHs2nOY+OAxh5ZMEmv6Fysb1ad8hAOLbhT5+31C7o
L1X9LK0VTTYrerigj05FxA8AiezpwAJmyKoZH5lAkk07g8hjogBXcifiPgFQob+6
4tk+YtTlGvW9iZNfK07JDaVR5UhNNZHPojHO0VaXmZNixBituUh9bRQpamVM7CQy
EmCGZk8fDytPw1e5VxFtFJ7kVmxjEyKxVoSKgnmHiiTmZLVPd1vEIrAmDvWOeO4T
NT8Gx+htbr6INrf/t55/MfMI39eaVg5KTwxAKl22YFGdDcsnGV/Y1k2oDLQVQ4DR
s1BMeG95gosQFbz+sFyI49Vu0BYqv3Y3YuuS/iOW5kBEcn0/deYVf9NjFb4cme5m
iA6zDEhgJ2ELvtgZkA0YlYlEitRCiAWLxZbWO3b2LZ8EmsA/iHE3vV/bT9wn713S
cCjioYzVOJX4RP+aZHqi3yrEnASqbzfzLeYMQ4ltH7l3RHHX8cxcL1UXxcE0cMGP
a4pho4xzj1Ga+7de4MgT1MO4Ng5DukmzTtoEi0L+rRv+PqKkxI53aEP0ZEDprd4R
la36ii1yfXeoO6tP7fEj5JJr2Bt8zPOVa6/BHVxy8vy0De497XaRYZouINDksobI
QrZ8rbROU9ZdUo2EYRH+HRowcqbVclG7IIENjlEoIH9zU29wdE9T5qGegKEeApUx
1jZJzJkEH8wn5G+GHC1zd2q8ghJ5k3nnytyJ+HlkEID2gpLZPaDloMpIpUbM9YCq
FCjVEc7JBQpxIfqdW7IyUydksKHoo28T/PUYrXGYBRwgO/A9EjRTvEwdrgLK0Ro8
/hhL6o3ik48nN4gCEaHK8OUParfa5Y7se674EWtjxTYdUYeQAUdUGuC/uxBTWvro
fUq9/Ok7G5Xkog3vh+yoBY6owRN5iX9HcWV5hmNLyCiKE5mhTiaqH7MTlHLGzOZU
6ksh+86v5l8akZ3D05/CdTbHhyEropsw43a0SOYVQpwdJtJx+4xy8uVttleIwQnj
VK2HfHKldPqvb8gf3160ns4fiO0k+v3gdtntYfpg04R6siPBTACewDmMrQRihjwI
VDjfh//3ooXJwjfkO1pwhJ2dmdYGXStpoyphItosORe7MNJvCiVadHCVPPm7oeFE
DO+B1rc+bnK/rnKKF67m49llQ1TYXe7p4x2UPlv04w96nLXbQ0WhaIBH9bO35jYX
wk0x1WeXrZzTJmvaTDxRipZ32gqL4OWlasUcpI7ak97Q0aLaM2nHArn9kbqwx7ni
x2GaKKVnQECI5Z3WPtHpvS5daFuHPLSy/JKfeVV4EWITui+FqRvEtj4hTJbiD+E3
SGL0z503fM/jBg7eicr3PV6BMT4IEDrJSfHcfAfN8zpFHVijOW1cNenS2nKeJLEF
foUtBIPRRFrwW1lRWkBqZsVtn1rH44kJhkEIgr0M9QocYNB4K+Tbtc27JvboGxLb
DTQQGWF0A7hPoml/q66PJtgk+/1smQSDrrc85LKLfF6v1TSRfQ9pUUJkGN008reX
ZPtt7BM4GEnV6oAasyNA+owHTifVWfjTpwxzVKP4v11tSqIimMNXKEStjRGFNns0
Bs+BW56277w4wkHViwcMFl5CFXGaQ74WHkzLIkeEh99Uc49hTDQCBeNq8zWeVmow
U5XY+KbcF4ws9C0oLdQfRHrM/cczm8czNZjGTgkXXP9JFA3TfWvV2X/gByd3+B81
wz/WiQ+OdfQyLA9n6DavOvkHNtgsVdqLJy8KfS8D/O9IC9DOKiyx+LBCUj27IIPk
uQQEMETBlOfjWUKwD7WfSNH/9AJ9xZr2+Wobz+Sx6LdIU1T2kYDFOfcr0zSMh+88
JynkjiX8q8a/0hoHl1qG25KqzcMaC1FBKSZ0cOcgXud157fh6OF4PQrsrsrUl3bI
JC/+6K8xbA/kpKa5HZ3NSM1vYqykkM0HzJq7r8bNnmALvhTmAwe6b7zZX28og1wm
U+E5d9tpUZunnEV8MMsaBycH/NCLzhL7BCm05YjJg6MZEl1lb/ZC095dWda2Ozg9
B1GSiLrhXA2em1u9OCb85QRri9pVmEm7Wp3j//Np5xSBaao9J1APKb80ekDT1Nfz
aomKrQfsxTyBc8/xBOc06gKS0tyjshmVWOW0ZW6uIauAzh9NI7RU9nowESLgq8Gu
EMgA1YqnKQPaVgrK3ZRlN2VLp6NvNZ1OfXzIenrSSnJ5+/LXbyZO6bA7g+d8TcsX
nLax+hZwcaulZfqfGJv+3HqwCmsKByj9EfM/RtucaDsAtMLMV7c1CMOB3DElPDIW
7o7bcGZa/aAUb7rAnbGuRPEpTOVpkOEN+Oo9PvSKpN3AJdwTSLzZsIiVfHURl+iZ
mAHddKc1qRsD1FuLqokownKdYqBYBQpnV+Aon3n6xTgIQrN6zTcqj2YULunEqik4
WZy6pzUE/emL7MSRECcfYlwR9S9TB21OcE4AavfSwRffH5xIoisQsV2KjcaFz5AD
LkhhCVWmy90yLIOV2+xZWifekP367yws0Th32acp31QVDuxGcSR5ROZKxXadpAzM
waMNONxUY7E4+SwcT8ZpCWBr4XaGJ8Zvr/lQVeILluzt7VX6ohbTKvNCbawwIam9
1cWYZxHFxE3dlfoH5CiuipdHw26C2EJ/0bZHsNLVsjIq/jQ5qG1z6CWK6MqKBHb/
v3ALjI/u9tHNj/gch77bGNgzQ7pCZK29D/xTdySBsBJNgvriIJjvJRsUSSwbLSdQ
CJDfbiO1bAfWlwJGTBMOOwqckq+JwM2SPiILIwtbYTxLeZAUsoEgWpLVgI7Cu2gM
txTXUAUqEfHB7BnvzovJZ4xYmgIAjtRVTs8FRvUIO1cC2jf81JWT1myUg1ROK+yq
gYfQIFPb3a6NAfm67DLX3/K1bVrutfMNQCpq76sma63hqeHuj6Y6UuImQ0ESygMV
FWs7hMbNqtPCOVbjQRiFZuKiGwABo4AQKja1T9l8J0DYhOTFZOtpgnK5y5x0QH4/
/uzo8ZI66hxCacRXBt4cOU6Pp2bO1fR1edor8/ye6RJCZw1WLjxd14JPqsoQToTt
Typ8B2yO2lKIsdRN17pQzeasYupjzjBj7TDxHxoTenFWWAmdi5B0T6JNB/ZQjYuK
TvglpH4tpajUEainkdyB3PtXTM8u4L62CyrpxqyxExp4hSYe323TdXqdIuHw6az+
UvA03goR3ieAxYMbNr0lGTB9JPEVKP2bbQUKQJ4uMezMBbIQTCWVLWqhgZH6XL5u
IbkU72hTW1eDXgzlw+mjVmP6ZIcv2tKjIW2j31IUdtwSL/xQ6GcQlN40RqFGMXzz
qduE3PIAhIATY+jPnQRhacA5TBDofxOkAU5+J1G6goYVA6VDlttvMY8bfcGhJNDe
OHwgJ/Ovxf8psgbPyImM9/rUTyB7wRJZ8+/HISnFRenIWB/PXR/BgBfNlN+HhLpq
FZbzxgF9dLldL2lpGBfuzAexoZEi9A0hETEMC+cC7P6/oxLrAU+EZ7m0quEXs+DH
4fNW4PxlvVw6Brn24+I6cX5oA7G/PBAw94BK0vu6+dSqSLpL6MajvPK7JWhzeQJR
+DlWQa15d5nv3O07+tWqG+Jmvy3nwHQjR1N/+ZEBn7V5nIxMSciQx6CeRCLdD/dq
MDG1hptVKCUjux4l1n9olEkmd8U1UqNJswcNmUQY63eO+uJnLN5ZhTvGrs5q3JYZ
wpqIjPiaEkr2J2FgkV6S2ZjMOu9yAXyMIDRfs9eDYYJoqeE1/ZatmZvfwMDdwl7S
eHNQxqny9CG1W65uC512QOBDwHH8dCj151C/WdPahTFivekemSUbq8+McJnKnBGw
bwDbbgzmREToBdIj841XfnNSzXDHwfk5WHEL20m3MGBfrQZSlR6SqAK5NGje3IvP
3jKN2BSvor5W4VdF+z2+jvXgVwwREA4PqLp4+A/0jIOdeCXy0xkmn6M/UFgwUcrU
9tj168cWsAYBJJGMm5zx5m+zXW7LTy/5p100tTg7a3BFCJrbJ4yuTadYIYmJjIF8
BDgniLoO+QdHnbkuwXniZp2NnGfKdfpNkvoWnyY3ooR3iSaSq8yUk8UqvdK6tChZ
I3YndlLEX53n2Od97JIfLJAjnrt+DOeFreHSH0f1hQivzgiZTcapNV3oWdm8UFFZ
d1zyuqo3WLoBHBIPH1gd4J+yROBCUjzI2se5cfuMqq6Hkaszdc1f0o9g9wzHxuN0
Vd6wDWjAxWAJTuX7x/Ea31q/LdEP+ITTHySk4uWlPElCytt3lasR42kZxt9vAOXd
ezPx0B/qSbTXhLQyxzEcQTCmCZeuSUZ3TUMrluQuZb74tL/HXlyNpsuihF61wsDv
SULakhnhQTWlo9/x7vtr+9LWxLEU7DEqr0K9lfWk4AF2lkR7iYq6U5Nio5CWQ/Et
txbk59w9Fj8A4idu1uy+6O4PP49X8hd242hoyr4LJORrC/cgZINj4JnlkVuayKlU
pNBxuwG7rj5/+n4OXteZk9H6juEI0zadAmR/8q/ASaebXWgqVpkJnmgjMH1Z2VeO
TJaKGzCD5wShtzts18OSPK7N8LZTL/aDt96urPg2Nx9g8YOa8yl+WNO+IxW9hXdE
lZg/hcw7b4TU81aaw0sqfo3iiLMRuK8u41Zs03C+g95grVw8chcw/OZJHoLQBF/A
Ud8yPxPTsSLmoKkYQB8tdHEm5+5J+cRyW/vd6AXwJiGpQWl5bEoqJiFXlixh80t8
2MFAM+Tnrn7VN4IjGlXicZv+SmwXOXIqvjfMtxENpPxmHW1EAuPnu96bkGUoJgiN
fNLQ6CDCqsnIjGbCWBkJRyIrvDKLtqRzIYGw9rPe/Zj3r29xx8rdU0aQAmlskdTV
l8n49T3tOubC54Qy8ae3f92HMHB9wB1UuMQziArZjDfoealAROpLIYeMhkJDieDO
0sUpPcAcuBkKqlSw/45Pfg4Qhq3/ij00Yg9W/Vgu9/hz6MVnoFpMu3YNHBp2vptM
Q3U5j0OQrDP9VymQNrdCvV8AKr2ETSI/BEGFtz7+EaDyHktzIoQVdnZ+sBCbn0Ps
WtQaZtRj50qc3RKt8dzvFL3IbYxEzWnfpYVeDyQejD2/1T3wfuKan4/vNQeaBzPR
6KNcvbyV3YTAK7yQ17gr/NWLPu1epd3dade70VjkCiNA2utWz9faDiwuHurewfgr
kcGA/YyIZWqnEvXgBk17VGXmurw4kZ0QQ0Cf2XJXc8lZE6oaBZ8xpWOtMVOooTJy
LEONA2uZiklpDPxF439MesJm5CwUalUKTswqwuZI0EygvQvxFO+RfAhcQxSp8ghO
i2qaWZHwbkijz0gEOAQ6fHkpfoV0/QX97mdhnCfiWxhmaMRtYiN/TQEPZUj2W3FX
7sd7mXYakk/0MEfoivGHEHCe9pHRWL+KFmEVJn+gwpqi8e4cPabDaM4Xy71fiJdT
R5ILeu9vbUc3p93/6eVRDo+b07rUpDSYpQI5LvFWjwiCSDDdK8fXD5xwyRni6IpE
7bCVv3iURgOyVakDvNQwEEdjl5w5xZYW0tKlLwfjX25enJwZfXlhIKQYyH5tsOdK
+cvHdkV8sPvxNSHKKaELJKyjY5tRmZqslqDkLh9apAUReKJj8DTWgWIVbfE4js90
WAFLvdlKOQiRFx/DLX4nZ8TYIO2edOHKsgbLqwE5FJxoKcVZdgjkvUOmLTg8Jf8B
dXwNHTmfpytwnXBvcvvm1FmPiq4DuUArxpJiRCaZUJWEIRxynpwPHqDBNlMMdgiN
M0zxXFRNSeZ88J+FjNXD3VMIY0+lsoAU7usfPoHml446Cf2BhIjBFs6+qwPFMTEo
sdiJepgjUfeunme6cyx8Q2m0X5tOEJjLgGCFlvEjWR68/OC8yjAKQ6VhSzVyJjBm
VDGps+DvuZe9DVKWB9UwDAkDmFz2UTT8yOts0oY+EXqVMSXNG5ZdpQ3+2LbJG5qe
/ugHFFLu7r2bK7ZbzjaKaw+cnhfvWmXopmafmTVjgNsC0Mhirj8RKHfB5v6N3lvq
Y6beI3OjQrzeOnE+VOhjQYXHTOxS2b6yy6O5VsoXIWOaKj6ipfxBZpp3X7yJWh5F
hficpGN18aoV1ODnz6lc4aCCXTP8IExt8+7bGZu+ILFcZ4GfCeCa79mIUuonrmJM
5PrBFj0xkd6fMVYZaRLZtRZgtlhfhBfCNuouDqS4UE0VcxAMMDdCYVQ0vfJrfhyB
YtGJhmOGiYTsIDYahu4IHvjGaQFXv7QCN6dUYcKZ6BVhjQGuFUZDuYGC46u0wgtB
OivghM4zbo6z0U7J7DuVyKs0+zFgAJjkI5sCwVweA006AIntiQoLa7lHNSkUORNv
c+6GYCj1LK/c42Xnli2UJNG9B8GrsHXQIU7bSmhVGtAPAl8BCOO+X6uXXOaYCqj2
ByAr7qhG/IzVZM61OGxiqn0SO7HVO7PqPnjAkqfpkPoa2tEDRQv7DYrGqTH6i/72
gsq3QnOMe0/Rs3crvhzS2yzGnydQe5JwfWdXsmYpXbS4gpEm/72IEpngcgNLxY9A
U3bvo4wgY8Uh6njbtLU0Wfm4AgsJKioAWJh3bXkOzBbnCoY/9SPBcsoCnHyrBGvs
vsMJVmCi/zLAIdVDNZhTJVI9I2a0LOY1typm7SGWeEsvaFqL1LfnURfvmhSP+rjZ
iXZC86Xy5/c+X1TPS1eoJVXiawF4CMCDLR0x9NG6VaLNEDZwHmZu40/63dw2VnfW
XxMKANCizay1Q5KWaivGHO1huANMEUD19xdb6+3WGMyAyfUP93Fd7UDS0CPqMoBP
lBuNCObKUzomEzeHH26NJHgRUJcd14V05xbEhNTH1dCQVTT4Qps6pLzPIlcKw0hz
/KoXIhsuePYl6+eXTswQXBoWVIjRLhIZ7qTGMKIBAz+LD+NjtVdY8jVhlFJdkNZk
GeB+/mj2krCkj2dZbmdPdnKJhRMcSggq4wmKB8aydgYposEJJ1kJjJEQpwa3djIU
QUf+G1mUeoDtB+moTIZ1Iw6J7B6QxRBaVJ2o0r5eWD4WODpuPtDgG51QEyNvmGnT
RI/5DshchbjYD0zYh89xifEl/vS7hjruafbUhgq41EW6/8k3Sd5xQZQ7KX/qOivq
oSU0kWlI0FmftAA1aFaku55MKmcogD/mPtZLYB7wy08aW/RVeNO4XyuRl2GkiL/g
lefhmmNWD9iJd+tL8QZ88eQBf7bWzx+YkZqhc688+BP5NH6tCGbF1/mMlltXsbkv
vebiyEuj+63212GBVS5XDFuyFBNhjoq5Uj0okksfRiNvM4+fUoWxdjqkjmkLGAFb
99Dcl8+IV0SPQlowNWF79ULedut+VB3dOTkBxtibz0mH9UihiiLtLtAArZzHaEXr
Kzqk6aTmjObaYyrHGjUuOYoQwAsvMEX0Nz27J0mMf31c1EWltLdbv2HV0X5ZJmT1
5V8R+oRdECwqlxTPEM+6siCPvVETVxP+7dDJBeLOoJoLUdrP1eR3NskvPb4Ijgtl
cSOccm7hzPlR3DqtNCgMOel9sYj/z9fXmCLhNH8rlwA1gTXMyiFb0bkUeGfEYhlj
yPI4eZKOZZbZIUo66sPD4xZcnyIWKJq4xRDdqUm4GuMig7ZQPG13L85zX6bKpjTC
bLVyJf9+Z6cSi7z3daZhAz/KJNIrge6perbbS1i8T9qOgr7VwdwYfD8jC7fXwH96
bg3HrfXtYj3kV7F5dEtF5ZpwWEDPu9urcJ/c9q2vzTqCEGH4yJrhPjrPAzeKQ6EA
m7wImBHAgyW+vnuJ9seusRiwBGIR9p4PMLtHm2dNfT4UbOyNJCuN0H/0sXeL6x4G
G2pm1ydFPu0PVYtw7Uv67UC0PREaT/dbkahHuJ+Hc6+jlB2p/urVIRGS5AXRsW1D
ZVEygCZalVCE2QOoFnQVBUqtlBsR2pv/Moldl2v7ACKI5TOQaJgUa2QqSJXkNzyU
Flyaw88S0Y0zAsIPa/gWxFrgk4ijIePR3AZh2fcuxhzK1BdxabCWD98ArI8wGhY6
z4q5KPDcu2NzOPgbCPAMOuN46FD5yu0l+qMrFFUMBCFjELogz4ZcM0KLAZ+QbNVb
u4HTRbwvDFlWiiWrtakjExCHv5b0HNAKmHgRv58j/5fO6gunYi+DKzCR6hbceJU5
xH6+xz4zzUuhg/gth24dvQhI7r+kDnSIvCuMoL15Gz8+XbVCnBHJytvK3yIrgPMu
baDrTrm722td5xG/++vCKEzlp7Q2tL325786syW7ZfdmI134xL8I5NJmlASfoHAt
d2y81ROUs2gjottCp9ZoM4s7HPFEC6X0eZreWAMvX89se3pv6niyrGh8D+LCUu+w
0ROd3iI+Sz3Yxrhqi5wKhtwfD95YsAqdQeYOeOUT+BSRpKuVec+qy170CgQrbQwj
CmG3S5xwa/b4JbuIahT4SvI4QiTR0Umb2HUeleg6IcQ5aBHkI70DO/JluhUtX9m+
FyxMT5K3DBfQmrHm31NqrXPWLfGGRgjg1kAwgvJESuav0kMOXO+YcFLbguTqR4J8
AIInjjTlii2CB39ZGMyYoESXtJWGlW/OF5acRp82288+fiWi3oLZ+oYr7zCLdzwi
RzyGZreIItBpW4bchWgQuahlfbTFhtMje3AypirD/XXfgoQz1ynf2BPBmJ00E8F3
E9cPJrLMHUdU3uXq/umPGEmmNlaV5tvDaoYevW8Lh0uvDMRLkDYlt5VaIvdOWtFg
8lQTnUVl/DRJ+7YYTYEF7tYM+3RTJytvMK1BKgmaABvBrZXcMOL0EVNXoxKeUDz5
jTEsjKgXHJK5viIrDtH/WgPS2NbGWbzLJrwB4/YI4muKEzcPMrXePPicr0KLjdb+
0bwKg+/I1YOf39PusVV/xteJTefs1muadrqn9LuwIqLUv1xSyzXzppjj0K1cp+9i
VcyROkkzTs8dreaZWlO92K5H++Gpmw2EX2XsD9odzyXI6MLBrkPtsIv9HEgxehZN
aMSbsEJKZnreN8w3peNasFZuu8SZvBDTzJCCTAJkmPeAZVtMP5u2Bjyp4L0M7dtY
KKJiW4Ae/UYeqzsVjav6Q+ONEnL2g4QyQF69TuIQbFrL7O5yHmDReZjmhhXeHDCm
/OGZ7eHqGLOwFI5uasD3SWrkOQ4UKtZHQPbYvbf+N5FFXsDPEz+xkIh0L/kBmpM7
D5XXN/epajsaqtKx7ZhJ+3oAGi6q8/JShlok6XHWFru3CgCrVJM8Q8xv8h9RFOtG
0Vekp1N34/tvuq1GYCIX3gYCRIgwodNXTIeocxSlUxnoo7GfguBlI/6bK8mYnDxr
2SgWOHMN6ZuQFuntl5AIAwGZ7jCVYW+VWXtSPfx1PB9t/ovAmXAWwckmoV5E5IPv
Evi7WKm4X56cEl6Ym6J5CUdj1FGhj7i075sH/71LF8PcsWZKoZ1AoXuvV9ltdhXa
OASTarELZme4o0rH0OU0W1aszDFQ6OylJ0ZQ6c637DMPocMrHx9JY77q9anVK988
G28m1Oa4d3E37LJzwRVYNTgCSKwIADeSPM1WgFboR0/Hzf90/065kXMecoQyV9uV
dG3XTYTYK8vXtjWGAVoyLELv4RnYHAHooBW448Vh7Ik+cnPVsq9ARheGqD6EgoQW
x0RLBr47uVx9r6/3oQQ6mHsipRvnOe2fxJT0fmck3fZCzBnjhFLI5wc3IZXPAHsr
cBGXy7VuPy3Oc/KQgcc8uNEQavNSVrQulyIIKTDZUWeM2GIH+zPgr676ztiZJlLb
4x0KHWbO2+rVvkeNoeIcP/K1PNLMhIQdxhLRWVmPrnMXAs65Tpb6Hdk7/Kwdwgpm
/j+4i+hMuGNm5mWjjxzNjiInAwrOcZFMMdxWNRhrN7wEgb/UDDCuh4haxBzqHHbv
CFL7b2aiEq3pbgUjgAjyvT4BjddQx/b84+mkLzcs1dbYCc+z2xDj/uje3P/U8e7c
TlD60PefULy9i/fhuoW5bj4rMBCBC5uPBA+pGFTCE/itRAZ9JltgTNKStbGxZLAV
ZdK2Xl+WEHZXznUwVVRmTnpoZNAtoFvpLiVMbwfXETnrjNKtWOBOFfJ/zGkgjJnk
JuKlxOz9GgTujUc+y9QPQjJSkoXQLslwZRNqoOKWniKJfUvZNcCBqKrhsqxq7fB7
u31/ed/2jNXCpaRGvb2p9j2pbKb3VgEBZj56msj7GgvSmu3ZggM3pvZPIAssUeEH
Y42lwzNBC/oIsI9AA9o1qhJ9gSu8uPX0z2H28Di3qJ3+iEnn3mqdCvIF+wLPArK3
GRS3oGd9YN18h7YZwRnKU1bK+fNP0JQ4Q9VnggzZb57AVuwokBYJkjzq0ONkGV86
dmKehoc0VzRK20LVsKyNmwBdqFN1cNDq/EgUL4WzZnZk0G2vHqO++ACMs6UOK5Sb
9zZy4vYjFlg+EVzFdRPWag5/tAKhu5dVQBqST+X9aL2SVLYcpYlylqgllMEuC7lZ
WCvQ/sHeypOrBcoyipcjNqocspWfMIjSKzna/rNa1PFUdeTHEkxtl/rsyGx3IxHi
xSLdQ9wUD7xA6bESERrdHvGExVYG8ym5POfcbczV7lH0ixU0dqneGHHNNjqCbexn
8Nyzv/B4iNeWkVwwSSiQw1/Udmtp+7Z/vT6TSGRLny7Ci3AP3jnA4n1Er9zALZfM
oQyt4SPdg54eNPY2+w3VvuN9HEA6Cm91DJHrCj4/9RZMdJ3PS+EkxKSzuOZ5cBjC
YkPpyMFGjT6MhGlxH3zBPubsU/MVePpeyqNmOemmUnNm0kMPmh1c/bagdXnLZ1zC
VX/XlIbSR9TtTXgpaxhQB0Iky1IwKXROd28vouiPpmwmYYwFbLdM6DWDDUXjVWRx
pM8D+FjTL/71kyj1PQz4HUYlKlofteSN99C2STsjTZFA+n8Z2GmyEFgk7c0cy8+c
azf7mTIed783gKZD/07tV95WV+W0sGa+RLSCTJdD+sbSjaCbUg33UKdW0BLDLnft
DuAacapo2+2ImI271UqHcVUkI7hcE+WR9DJmgDDViuPDte9TWexQgnfQiFahvjmb
2lpxk+XIsI/DyvP2c2qv4GbCKNJ28z2wHMtHxIKmbxPBRbi6mACY0NPk4rqvj7wc
sGHeWON4mV+1m7xy/iQ2uq3QRgkfehiL3CerAkj1sTnJrTAuouZPjRo2BI4DxsfW
124wfzZxAeRJpUk+/PWEL6BKmdTksZgbI0HH45qWsy/fW+q3Ywau+FN3wFdl0/ef
VcAd9lRuLN2wGskUgM1ZSaxrT6JIA2MT2IC0URBEDIe6YRmfwZwsoWk+/sDP1d/o
+BjazFkXLsymkGtVWmIGuspezIT5UgLi1tLcqVUOQqC094PXpNcMfGtpGaq+daPc
k6yzfZhdcGQS2FWpmJQ47miC3glNutsbW7v2ny6eQD0OFHmeILMhiE6PSFoUkJct
UopAf3lvzAKB0XhVpgkHYgci0ZdKG+D+WcfpCf1gGA7JZg26CdDKsMKYpTgKWEid
C0uxsoHMCZRkgOua8bzqtSitEIk1On3sc4i/eI6n4D1Z3824t5JPpBO3BLXGd68G
wHIri8RgvlTIkzTcHsMi5eFXHzGzalY3+QX9gwdEnFS9aVJLd5qckMw5J+Y+PZ21
abTd3atRzc0ZDpytyL4aEsIYig0mzK/+qJyT4KkHqFBJbx+jJz1aga3+Ais/Npwh
L0rb3IHgYRpEbD3/9f1jgnvBfbRfLveGbryOyxxBRJGLdQEwPD5WA8uwh6zut4S1
uLJAzWQkQwM1NNxGGuPtMfUitcc4d1B7KP/pJAxfzYzI7BWyeOvnSYeGZpVeBt40
b1dYrpkZCGhsYIFeQiawAaRP7LDOhdcnjbKzONT0YomYPjx10l579CZSgtSfmAC2
BsQg/VSGqdJfURBAf8jBU1sA1dUxcXwZldJw3MCO2zBCN8IBXPTJd1mOFSPGH8ZC
Ugda4EjpfL/wMOnAbJ3/2S73QAg+jMWxC5cmA3E5lRf+YNkoxeIMDJthPvBs3L+f
5KNTJoTfB4LNgHjEgpbPdqqmdV+5shAdX4aMALX5E/EpbjrknjRcPzJuSJsExPaf
EzMyDoYt4aGyGx8vWVFu/UnbOzpJIY8/XNKPmSpvZwV2grGp81X0a0dRO022Fqyy
pF/iBxoDrTLMdffpB9S5nTqX+QMR+UEoNDWeLvMqQJrzTt14lXHGlRp6RG2b6yQ9
OWKexuID7VsBto1Q625bE7BHAsrqOyigjKYXs9Ab1bB1zReg97rF2O9vMHzc64Yo
YMwjdxuJJWBHZY0+yQYoJPpqrkOTdulmvU7EKRpuiRZJfpI/Bg4rQGCQgX8KRZEq
koq3fI7pnm/mE75eR7MZE3U1CUdrYkX/Mga/c3es8NUPcccNwfJjPOrnThKo7Igh
cHLpTQenqsJdL8R36bnxCTqyzTUdq0Y3ar3O78T64Y2YJrFXn6AMY2L2ZzV6kOZ1
HTQmKwgkJMJTEkDBnLdOZ9op2STl2TrJndqFm3/EnDvboHQWi5Trd+CLc+cj4Q9F
rmQOK3mWq36f4irCJIpSzDJlbtg7aLY717afiZDnrvT+v+nI7SjHiEAlDEszXehr
LQu1NvIU0Y0hny1FcsRrO9Uh0cX0VXc4dNeEcJUbDByvlyAe4YgBSrFs6QA5NTgO
/3hzRWBqC8SylM/sn4paWqwoJR0Bl7Cq7cWSHeF0WSkFxLLVBBneDSv9XwJnXyS6
j8SUqE2VGCvoRy3qDy0I130IU9duRxSX4TEjAXkI+SL4oqUXuxeHIl+KncP522cP
/9LLlFXxFVwH6ntjMEBK67sXArPVERNH2tPuWO9WAKU46x1W+i8KZEIxhlCEmp9o
Dv9p7lVjIPKmuhjJs3KnOmokrurS1QLLBAwu733LqkZiuRHwVI169msxTaQJwiQF
CmYvAivuVmfsVZXwt45r9kauJLvTaCkHHRTq64LhtCPJL57/KQ0F5hn2K9oT3Nwb
HQbB1rnzdgudFm7aOQrxFxrLAAlyIYfY6mSvI4qMN9OIE0bq3PWoRSbbyfdf5r6g
GbbJZyHHQjiv0bguCCIxdmNEqM5B+mRyh+yf1GZaYXAEt9inA3/CPxlCLkVjt/Oj
TEeceS7PclgWhUQk8VQJ7ZLOwCm1vnoscQcXooq0nEHcSAmTz2LURM5Z5g/v+qPz
DUwyfg4vddk1d/JP2D5RULbvdjUCDhu+P456AfSG1ubHZnYFnLXReqX9920UQX+x
8Rg6D/jeazxeaXKpOWzUBvewL6kQZtiTFXMW/l0fhdidrgpUB/jNU3lpYM1pRYNF
YhGmu816LYxvCpXvqJr3+46Gj6dY4jdCpeh/h7SrX/nNk3WdxKs8OaGgjNKvT2dD
Zu2DLOx5IDsWHpS9zf2gW/DE5KrfPb6Xm6bxGP4zJmTXIxeBqvecqeurkVIJxtvu
7E1+0kGJFKAiOrQ09eySXAMbQHKWACsdvA/NruSf7fnt6h3F4jK+grVtw5C4zyX3
qtPaqjFou2JuQWm+f1yqIUE/Qq7vVJ218oe6UsTxnb60svQ1IoG1uj4S4/6VIfPH
pspTHGjQbsK6k/QPSEPQQV23CHpixGuySIRbE46ghlUOGdwArCcBvGi2kp4c/0Ky
jHtN6sws3sGUFnEuGSZnxK+ph2ZkrjNuiex7XWNRanaYPko5ZR47/uBgZTrT8fvM
ekRsmwtQ+KI3YVvDhnHQSSEiVV28IGZkU23Z6qLcth/tgaNZ0oLT++fkQgNMb9s/
mgTmFuLsu/vLfvwecEH4/rXiCKZ1ZuHVWXPe3Y5qR/XcTP/UsB7Y1Jm5w8N4ymcU
VRTcr8iiADyBNKC1mMU/F0vULMqz0BPZmHaDEMMIWj6vLVXHVQ7SnY+DB03hi6B5
PN2NXIeOhtbry8vkBbi2zZQzDtYaBfetgjcn29/My4uz9Wj1vk8ekLMxg7G7r72s
3iaYhMZzPLTNa4rP8sv/Kw7bo/OBA/M3MbagjXS+DfZ7UyxcgSsYLK0bPgau10mD
jWIV9+Mpq+vfRI96omhNwFlhUoIns1d7iorou3f1jIZoe/b2fRCSy/CAb5GYZ4I9
BZQ3QcWIDfAQsYp7oPp7Plo5Hb50Ee9X0ghOAx9ojLATo36NQHYL53sDqVQ7nSy1
NcesjNGTAwouh0t/TdvTygxsIF4hHHw7lLk2IOhdQo1kHpLU/MYzR9fo9JyypYgc
1x8XkqHIBljqpyW2snMZLMTmx5fETCRfOoJuYel0R/b5fvErFiU3JI5UNYXBc8Pb
X658S9VbYbtXKgVAOzmtlz7ewFqkM5rtqMpzeALNoAbO7XBBnd4FkkyRNnqhPd32
WrGZO315/ghmxSORLABQCqh5ez7pBF63j+Hvr60cgazv9RuQ1ZFsc+/PhrVZ/8DT
J3CADrmJU7wOoK0rFwhBYPOyaltrTcVISrimOM6JBArQ2lWQBbnndifJ2TvItLvk
RsMB86fvAdo8V6aM2WFviFCzrm8lEFHiJyiQmqagHeu0DO2W9+JSU+3MLSNEFRmi
1vyOPxzhhLKMCxJ8ES9DahnBiKB1LS+RwOajZktGNgHV2F4gtZqsYCn/L9t2bOT7
Zn9ZQCXXDwMah+7tnw8tA0m9iczo9mQjAJ9FkVNdeqYrQttoUchWAXvHBQbpOq2X
zkhmjPsCXrXqT0SDwr0tiCDlzBhZlt4oMAwybdpxbyzZZa45Epb86/aVWJQg8TSi
kGAdzztN2J2VNqraCXJ5SmIeHusKKFWX8DonLk/e41VAse7jXiQMA06UQIz04As3
dutPaIMqU6qS7OQtPVvFyqukigsTfqDWW4yZrfmWSPby7uMSder6p3QZjssttaEe
OgUZrX90G1kk6a8JQb6U8dp0s/cIm1a/Rev449DKPxL8aPXdhzST3NirASn90K7v
g2KnyopsGqAXD+PFbKDq5Y3XUwidHt/qh9Mym+il2y2LDAR0IrhIvz5l8ULh9WL8
yIiM4MDc27pmmbkWdZXZPI8LE9YiUrXWGWZqfdjN94GeD9GLfQ1qGKErG9MMlHoW
AgpvJ2gI5DbNzuvqA0WsM55mgbXgPWawcL96d3fIcepJ0bipj/sJYQhUYFjlOOkn
doarDdFbLOf9js2p+/z3Kr7Zje+W+mYZQaiKwIBAdz+sCVoIrfTnMbfqWBqUir+A
t6TYsIQMAZ7Zgen42pKN/443bKe0RmuYIpgdNbfZrOO7aEqVb2mVoelmaRhABkW+
7Kg6tLeN5W4QptI5WegMLL5hut2OnJyw5wi4lo9ob/MoNLk2qpxnAD6ne7KhsWit
JOjSJlz5ls69+APLO6WpyCM1Po2aeyoa9lAzMcZkX5uYl24SsRnokSnWpkl3JMYc
DZpIxa5SZf2EPO9bULb96IMPQS+cQPspA/xIELDCEPbp/iaAhirOEXWt+aut6zxQ
u3uiGB+AKfvkYeOc2XOguiTR+p4L20v4dE2/k5l9q0RSUw7u2sjMjlvPe+epXejk
Y5Q5D9Li1/4YQ9Eht7mmzS8qsUw6YHneakzuwQrSxnqLHkXDbFhu2wn8NwZQm2Wt
9w5yaDsVYpSNlsaonW8Z0BGnfB0NBHcL4h5vph86KCSKzgfvK/j1fNieDC51Ixt4
yc539oIX3Ay8WzEi/reajp88C8kiPJpyfH2ctI31ZJcchdn+NnHpFMoJpmv1OXSf
DnuTyYs/O93feAI+M6NePP0agUAN44QsnVK8oc7YgahRMIFhIZUw6YSLRzZvZgFG
tY/dkag0Z0zhYiG2sbC2eqADWGgTxi0mkEw6xPScWBPKob7LMG3ldC3PpLuSm6es
PP+v2wQSm/Ju8nrn9MfH3grIeRGSX6bu820vVHPfJvebkSYAyWcd/xzRI5L8byX4
kASUVt1Tf1H+vS8Bx71/JeSt95zj8Ma4EEcDZCdnSH+YP0HqIjbRcXucnpjuSQM+
PY3/7rPxfGDV8saY+y176lldaYxh/dMEj2xvm/iDnSUOJx2ga2JILvXtYaYy3s9m
Z0Z5rrzHZHhov4iKU7TI8JNohwCRp/PXPabMIW85TI5cy3zbona8O6xv+q4fOm3Z
LbPked5tJkZ8L690kwVomS74puBef2VqslNI2IL+QHX3wohI7EWfi4VTeQqoPBnR
65JQjcCLGZ7WoBnlZMrSaX1zg16rtSup/Pc36c4vedCXqD+RIqGPYTV4nJlOgNjR
A3hIDhxkAUH2ictVJ9Mj3/uMoMzW8S4FFHw3O/ya0PyB4ZS8QPPKR8oGKhm8MdWf
9vKF76GnfETV9nZ7FyGlh6djDe6Pvk8zamBwMrbSJA9Rejwv9lzE5Sp/7yan3HPT
bTM4egoWtgLP5RIhsrRgwN0E0S2NyJSm3V4KhMARNps/oaqUmfZTT3qKXH+DSjUP
VtoWOcUBBw9iUgqa3HsiBazi9JqfjdoCjyEYBAKFqqHHlTYing/4Fb+eIO8f7/32
rRAWkDYC0n0/e7xJuIg6zlXUvcA9AkfHMp0vyqvXuGUyRTknaltyAIbvoix1ok2t
k9mIWGa+5neXFUCdw70zx88PfzOMmn0H/yr3kL2N89Cd1Vqk4ttxioED19Ndsd/p
bZiyS2AJQEnf0+/YVM6dLJQx28TmHadiY3azYVoLBMVvNmJLbfAoT09acSoWzYgP
aH4A4dYVzwH+fHrcskBygqLyBJ3rslbqW1QR6B9tDOZjL3PDmeoqdUIxeYROaM23
07OERel1NlnmUEj9ebGHd9RIzK4rlGLut1Rg7P6sXkUxSWViTxhkvlIrIrz92iLt
7jjVPrdXGM2bvfk8/ayRor4tqAGpE5mVsf8jSfECHX/6kzjeGWEYmYym79wNLzAW
oJD35wzG6cGU7grPpAY8krGZNFpyFN0iEUZRFAc8OnAe87LIPSrn5k81PscVZVe7
cyZH2BcmQCt7lwgUZDHWXtp75r60p6h+tvDpULY9/YkeapEEF3lnFOyFJxYEsiHr
SfHBDW1mdtDFGhlAt1Ays07oR6hhW/h/TZEdm9uefY4X/wPk7tev/BT9Eo7zIUf3
+iOOllSk51svHrfy2Pm9vlLXD6BRhnuxAkhKWWf7D5xgtvMr7SuRETq+5cAHB+9Q
KItq6m8jFXrKVQF9jcn5kH3uAPgS1Jj3rwFxJsjOngeUloecIRTek87EuvCc+qaG
aTMlHM9Oc41pT1KkuEcoRDeBeTPMrO1cFp9u/HnRbI2MNL6fVpwE51SSu66Xb/Yq
FPsLMf+ctHiWpp9rtJlJVxQen9QzEpPm1aP2OoOx0NSj49VF1oWjZHRGCqh1dhvu
kfMglEVKbwnzyEUlN9OceWbU5ms9xMSpMioedNk8hdcbxCbI1xrz5Y0ktsjY32uB
gtAqS7owCvJGUmkx+TZpi3baVi159Uk4KriPPgzsk47RVIUj48X1zjWEl6bmrWOr
f0omHQ0u3nRgtkCVfZGMHiZQk0KNYTp8+waPQzBXOoqV1kJklhEtAbC+SqQQR7wd
vc3kN2K60fQK9Pup3I/7FO5SZQtBncPaWde9/kFsoTTv5J8B3ndbWJGZVtqHwRLC
/IcqGs+pkJKyc6pLmAcAU49uJGZSWHVoBO60yntq3ZBVWWmNRMwN3vkcfcQbRwim
SaALmliMuf5HQHT+VoK1TviiP9fKtVIbBePlAbV504x19o8ArN0nFygd/52arGjG
`protect end_protected
