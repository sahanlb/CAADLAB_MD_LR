-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
me6ysFjKLk4vhmYDnXznYhAvJWpVOFiDNAiifwwd2oo4wbrX7AE0AVpmajOpJ5Jg
fb6prjGqRtj+GXxndaCSkqjdDkh7p6YNcvxpsHbnIEtL0GKfwdcj6JcJ6ZfkzkP7
d4ZxbqNmW4IB0DM65PbcUHOkCgHM85VKR+cxdW2kgqGUBwmQup1BHQ==
--pragma protect end_key_block
--pragma protect digest_block
AhNEgk9WojdyRpYrDAypKQ6jtlU=
--pragma protect end_digest_block
--pragma protect data_block
KwCED9U6jBZALNmdI03qXyfFeqDYsLD2w37tJY4dXspI44y4W1FVBMxvCNXsmykl
sIEs0ktsLCyJd8DRezIEviv/jfORtrTx1SeYG2m2v9BgSLJI6CD8/MJPMkscf88Y
w2peyfXxYcXvW/yPOR09lSlW0yy+nCuwVgHQCPe148HhVEivWqqcaQaTtzhFzjWR
7gjY8GKoGM3T0kyHj/DwOMZJ8jtY5wVOY0qJN4T2vkji/KXAShKfy7PwilVT2il2
hhlWKfHWH0ibnuStVzvyialEDGCbjy537hDFPaJG11ZRSLvpl7VSf+2fL6nhD6Op
xTGNjrmBIv2DBEU5OYivN6aDgq8MaBUzC3dwRI08flzb5S2wFbnrIxoDZEeKaZ/m
NzburmjZ1ToKMAgg+Yqp+A0PHbP8xnybP9AzJ77zFbkTXafSWc/3NDYlRdm9NUxO
eColh4W3UxOrtZcMw6G7ttV3hm9SvxYjRhhAMgKnQEq47wbQPY575bMyXev84kSJ
Ubpxz5X4wm9PBTOAW3NFtJ8Zxw8WMso3dtHlSkJkzJJ7tc2v8MzIkkFnN654Pk8G
nA/3gXiansGTXvfSZdvfGrp0JB/9hcWa6dHoj2RLx2QKqLI4AmYPtlqUfnk/oBlZ
wb1xvJvcUKURp1rkElu6oBK2VN6D05OKr2nqNvwvTlVFJHP2hZ1Q5D9GKe4czxyx
L36RUxiTe+D9XWpm556lLMXJq89gnCzoLtn6hBDGxBGs5l/wGvq+IhE5BzJ6PvPv
073E4CYP5lucEuGja6O9UWuu6nkvXN7FAwWB/l4BlTeQQUOgL9vZjdFO4HDRAAsn
XFhkRUayvPJ5l57uBF2DuL1ax24zb1yhxi70ITunfPjMZqWJEkXhlsHN00Ht1Uhy
E/kxELnzxIj0/SZ6a3g5/++BFFa3IGrSpR84EhzmL/1ow80vr0Ce1oVDGKIu1krk
FZq/5QWjaCSVLcTu58aW4HBScaAKBG1uVFSlJCwifrNSBiVhSNYGxE26g+9/MWlC
hZDeUFN9SmkFrWxUuPGLjAbDCVAen8rY57E02orkyFFfyRknbmq+t6EQUiXejkL4
vt1HFozKHOIC7OB0TMrLBDtUgi+eIkl2uEV3zd2f4+dFC4qrKiWWPlnovNRj0F6X
9jdlSoJQNkUbTweoGnpGxmfj2ZKSL899/HdA65OZ6SbaOIhNjWkK0gSOlzJ0/AZi
oESZI3aYxI6S7l301Z+S1GeLWpwr4RcW7vdb1FMfHAfqsx5vWqdtS8+f6dh1hGLr
0Ya6qy0Fa2GUKqgfWohFzeke3jEsJwcGyc5MeOyCyDQvqKp4Hxk6rsKQs9t16Nl7
a6gGpclYk9A6itJr+4F0J56xsvm+4Mm89lDEdh7ipBCpD+tGoTt4pv2yFr3c+tDW
HDc1N7MrBnO0wXfPq7+Tmw9c0Az9Ph3GUDfD7HlhLi+lOtz8efctouKoGTE4FATC
c6DPL+PvQLoXC37Nb6HJNVJgZr7YWx9ubAhJQP4SyT5WPVFDiCIj1aHdOUl0upM9
kxSh2qYSzdGxqz4zBZzhxyZ9As1wy07sC/mEEiA42tdYzsxPOY8YdiIznULGsMz2
V9Sr+iBdqu2e+oU8wP8D7hAocbF4jK/YmMSiJmfaP+CWaf09nzNuVjiQZU7Lhi1n
8DnKfKW/1WLc9ou48y2mDgPVrt0YdBSxXRzjSrRaNF1+FQ1SolmN3U7M2CDSYcZc
1pFsDn6yVurZZ4EZUahOdR9vEcP5h9L+O4dWrqrw8DWog9T2k2E75ZPYQsL9wPbT
cL7Yu+Y3swKHzeSOFddY24z4DjbN1p7fkyHL2Y88lbWSyvd2wBxCKY1fZftlJFL2
oZCLhd2kOTo7PKUA40VdeOvG3af2qKJirVJiQKsRgLV9hxCfoRBH8UZcCyBU2awD
3NyLiBVWlsrr51ydzfrqYe25FkSUyV/jJ16nu3R8mgwCW+Uf0pT47kHa249q91u+
/HBVLpiIefcwES7ohw18oEQU98kaa7LO18kXhaXzpezTzai+C1nz11UADJdxVh/E
q0oR/9o497mlOQ5Dsvnctj9i2jsEBROb99Mg6rQpaRgZeKYYHOjSVQQ45c3nJPpV
PfBlYCybCLyVyk1wfu9QrkjSqNMNbZbZe9spJ4Xy3FHrsyF2WAGKKX2c2WsmP18h
T+6vLUSjE0/cuW1DglMqAaMai3n/h60d8nWWoLEFm/KX/Mk7XXsVetfE3+6duW8W
JE1nU1yrPPsgSJlpmO4e4ytF9i6mhViNCp+ZS2wuUHuXRwwctD8k3mNng5TN/680
LfKPPinMAclT8Wb+pA8IRzf5X3dlTRq9Q/H7sN/KQEyPtAFOHc99r3T60uxANoe7
bd0iT9yMA/JCrFTjZXp+38JfVlYDApYDW+x1c34zc1aXmf3A7KHMoQdkO2rFpPYR
KbvX2GqFnbXnxHVARGi3fmnnQwf89OJS2MK7oXuWDC5zI27/AkydKFrQShNU9hAI
YX2vY6ERDOTsedSLe+2wVDNcgiYL620PcGTa+qR0YiLOFR1FyQDmj/RYmdtNYabN
5qggyuAblTzpNpZIfUcpboRTakYF0MnqkL1SlY7QbBSqtF+QqYy4QhEf/i0Q2282
MYDGTTLjB+RnJbfKnWbdc9gvREU8E8iYumptVFtb83ZqTs1Fc48VYEMbHH9vxg2b
ooyaroCT0/grCZ5LcsvhrJpH5b1nOp3zJRTwOQTEfmFZw+97PVIUcCWrXpO5/nGD
tZLWsNT+SCc734MsF8VkryPrts/GRIYnffxdJfTKoDmlrtGpm29lYiNpF6m1FDDb
8rmjPMCQcSCzul119bSjxAqC2R9Zp4YNYk26NMJZbMiAZHxVGrArRYGKEMNPeGnU
Cgb4sC4mARJ8UFV8wDrtzTE3PZPxyQRMQLDe92JvO23/sJxW9Cshnx2Ez5+KVHbN
yrL4XmY4sMxe3+bUsJMXsfU7J+4J4s34xjIPokPXpZap+PvWpGWLnzXBeR/Te9wj
bc2uPHKTdDkces2sblZhGSNQVeS9xNWqOXNETkFNezWhEzQDd3/cb1hvbhbkX4P0
umOQCmLaNMPSmhq+iJHYk017cEiN4LUUnp2wUgjeHf7E+Q2P60IDYItAyKTu3jr5
6tG8b4iva82vgHIf525MnNUWhWDRw7Bq9suH5ber31XeuNnhCdRhlTw04LNHoPhQ
HeN6/LUACBTUYURMjezZTPRt/GJFOtRBi+Z7DzyFtErQU6JpR6udHaUT3BGCmd7m
gmOPjJpLtHGkykUSdLC/HL6Rfkq/gWKtRe6prU21kefgbJBZMdTO7iaA0OEk7BfN
56RAMA61MfJBV16vJw4rbXBasWd4K4ctzoBTT91yvZYpgawOeK53xMChjOkFFRtR
kKKnz0AryeEU7fYN1QOgHIyhgMTgsA3mtkHLI/eR5TITs1uz78cHqzNHMS74vO1J
V01CcqT9X8BqSa+LTChkfpN5DESDi0bbzJReFPI0VeQNBCGJlS0yn+NkQAQL/ePj
ZjqqnxpIjC/bLM6tOp7O3WVqmmCXRdsK6FnCME+q7p0qqNs01DXKZ/SNVpkELrkC
OT20Lo47sxFvfU8jkDT9fBQaXxe2iclAcW2Olg91e0+kCzj8Ov7dTu+S6sFJrOf/
LXh8xdx9I7bN2PUj23YFANG/j9q8hcHRA09/ybO/L+ZEC2B/zIV8cCr1ZzmUM38P
Ti9mHih6OYRFJAEqVvY/LVxGW+WgXDCQWBZqkeYeC7x8qlefu+Hb6+7inKRbOqCI
Hwtp0Vl5YHUQxtecPPbqDl9HrefznphIIy+D4yRTUbs+Oji0uDyDT7R+KqWe95X9
Gni5rUy30nNeYgM+tTb+reewM8YcI8RGq+pFMs79bVhPZ+J+bfA5HkH76STdjXzv
kvbXDouMNw1EGA5w08OE5MhncfNV4LYnr6Bx3tNS6bxXNR69jG4G4ndQh3lYHllS
5ahHXD6l8tXkKqDDZaHJCwsFNqrotk+Hp7en6fTOAYforgUVIm3canBLzNNoHkhD
kJI/cG4uyCNYuACfjZU67pOemOFLHKPXSigOo4wfWPdfskvK7v6hOAm2r9H4wh62
cBn4fz1vWs3ZaEqWCis0dL7Q++xDWP0CuTzILWwcMGCKcUGe/Ga46ySy/QOOoNPp
H1+owpmKCp0eCfqM/YEPQLoabinkq3jHPvWsyqDqhSuXLCFRsId3nztRAW/UOUAw
TiZeL6UNaqEeBzCg4qwsAf8dkqjuv4brbjUP1Qapk4frM68DL2zXFgt5CKN99d8f
hhofsOAvwAPxSdTZDyeYki8XdjMNd5mlYFw54ZohhjRJeou2AQqa78HhWH+UcYgh
B2JxTXIChG6xiVWh4PHIRLKlmRsEVvrcwaEhlcSbIygnRG1iYvZ3EFqL9m04ytZC
3Ge0zAcjWbCqAN5y/o3YlbRKQ3AD5Ul7jyjfk149gazSESJ5GZQUWJxdkpYbi1OL
xeUVj0rL9PM3XDycGPWhtek7sckicBhXNFW25woADteQOUi+pKy5TpfRh3PI+96c
rupa1Q5aC3QHtCKzLRh0T0KT+nv/AOM8yzZ/IY6tJlbeejT1VsA4J5xOi5+FHivR
+ixddujHrgL5T7qk7r52X1ebOfdtj46iH54zJaxoF/o9AGHSdAoYM6xDarzLrTKp
zplBPjFIJvFHaLBLH6rZD8zcUuOguUTHjpZMlf6VyjnUpG/QIbzwF41kq+5StEtM
LhgOrmX6KMk0VDSoufqbRouX2Y22w3YkXnY9cm0uDnnbrADDa/6eosHpGBh51a5s
7Q5q7ZNGflQ5rZkNEzbID/TdPjojTdPOi6yf+V3/J/87cIJyGlC1Vu90L2dja74a
lht1FL+tLNeNKGDLqkR/yR7dbk7aOpWgxkU3zv5PWGmtPUHo9svtdHrlmS7zcwp+
GOTfesIAQ8EAFNKsX9VmrjD1gGgRgfpnwcTzLuDDN2Sdopmrs8Fgw53BPzPtnYcN
a9r87sWPfRzj6WLTByEOYsdRItwm/4VHF4bgTwp+DminQJYVgdgXB2jxwG6e0al7
RdEN2emTDEw0ieV4VMReXC0+PINV2Wvdncz/Qb6s92kHV2YfRlA5pINoNdYuvjev
CyhrZmAegsFwFfeJaq6FuHTbl+McsgHT46IKefCbyNmqJLMvi1wl00ybPV7mKnz9
Z49kzgOkPppsP2C0bJ1jzpK6pjHIUFi7EZvwaUHpVvwqA4zz/ckXVEcVIcPLyU0B
LKXf9F/X0DZS3FlOopWPDXkHxJHfA1Gl5fz7uJdPrN1PsMWb/pa4sF9NVLzaxNAX
jrh9UlDmDG3pRsWjo8IeOQaqtohlOeSLuFd6tcmOGiimiMIne+2NcpITKH+IMsEC
W8VvemAcwqdutBG5zj3j1KC58kLK06XTq43kTh6cIxxL9B4bYYfSYGp6VfKfuINV
aVeG0+opbtWotYWMboTAp5c0cE6ntvTo9xXZRYJKEw8BiuDR7C1L/Soi7/vZ4ov6
bslxhJ/HnmcNISz4eUf+8f5IlgD0ZRp44By3E+rk3IdVKY3B9B+RKjltlfsORZ+W
mqD5qTakkzSBThn6Vy2hLSIj32S55G79Wra/jzUrusi5zqUdcaSaMMNF2MzR3XN8
CNNMIHToZu81UfPCmGyjnd/G6Jad1cfx9zPtR/caxr+FQSZliD2rH9DVEpPGK+9H
xw3Br/N0Jcl0RewWSYpgHRB56awhUmJFPL3BB5ELhE5zrl25YXQpNC12d1Ru0DdL
Wha4ji1gCibKuMssKOofAg5CMUzHW5e5X3C+IcbaJkWcU3Jj6IRlcjByhAtPaQGu
jfcflT1KPuCPPVZjMVRlpYbW5r584YQxC+Bo91jY5Xvxo5Kay+L2OgTZ55JtPqFA
mmW0Sty+WJPZjE3FSqTw/A/LMdr1TUBBOvY3PcQixRk/ia+4wXTNGbyzxE2opZcx
quSSIvlyRIHuf8ij8fmMEEE/ICyQagKZWUeqsvmPk2Ec/CXpaG3/YBNQ+8bUOV3r
LCFwz1syK/wZxLFrCfEo8RVBOqU1o55b92OrBdYeT02Xtfq3WYJnuqE2vAfciu+f
G89lSC0svV7xoUC5yFMsd2U9SzkLb5cecSfeF1kmSjMQLGEmYBCxxHQmymidLg6F
PGvZVkn3YqbUtdjA0H9XFW/SAWgEjmO7fVbeRJ3Gq6Y1tBrJ9ZjADM/wBAsYdugq
Ab5/J8npIrk0HD163nauagJ7QH0qxv8LEeTlfrIeIv+HSW3pyaIU++Sx1hsLymrE
6FbO44ZApMcnhcxaI6gntgjAALFWm1yJwqBu8F9IZ/M+WM7BR3blrFMjIV16hl24
L9aOw5fjnwTGIYjSC3yNeqasy24F2CptoN+Q3CIwRfUWxpVdS/EZsSJQ6/CYEAiN
jHrctcUUR19rpJ64nyk63eWEYJYRwPzGmZY+eRQ+CRSqodAbuFqAFBD+h/Z7JjPw
rahkFVP5BSJGxjIh3Jmdt+gArpgyolQ82vhdPHYt0ol3BhC35NKR1lIekOLrrb68
lx89KqqZ0H2cPHnPj5PgtoJE73JX0IB+PmrpKTW8i6+RbhYK7qmEM8CZUriiSRNl
Q6E6X8OsYHurGb5yN4qZURBMTht54yK4Z7wV3IwbMVdQtdy759hq1u3jMAqrqz0K
INSX46KlNy5VV+eS/eHdPsIHuVNUDghea9Rr3YXFXl/GweAyv0KYYCp/1dZmvS83
y1ekLmT8E670D1PrVZBBuPhbXCZWy8oMI12Zd+P/BuKKhWF2tR7aTUf4afNkqy9n
s0dj5HFqh+VvKiKqG6AtYKiqrUkFiXg6NBklAGpPYrJ4rjmtvElVZ2vaOewwCz9X
v9SyPedWZZxcfPxHAnCMVj0L4U3r5C3cAVDqEnl1Y0ZQ1UAt001DqFCrtV+Y0l1j
wWHPC0dpMfIxY12WtI2Ghga8CBl5fh27aF8XI/3hDRXe9/8yUrFGQD5pv2lQNaaQ
osueQDT19XmVzVLBonPYO3+jPbw1WmUmYOGuSlLhTvOGFcG6dxEsn7tzU5sVRAf2
t41nFFjY6kiewsGsTwejDd9Fur1lit7ty4W3yChYadJzc+R4f8g/7SfrA5Htil/9
RDlBeuIEmMlMo62VjlXDHoM73Vcv1TVsbhRE0zf/OQAGPjbPUrCWbttPRzcbPNqf
Dw3c1b0yi86NZunlsEy+NQnY2bCx3cmoxTPKroNruM1XepZw1DmXmBMYDHqyZMHT
N6NGSrFu+qZIsmBUcB85C4axUPOY1LcUKmQz9auy3VcAK86o+irm5fNJ0sM18Vg7
fh4SZKwRo0JOOBpuQ2vsIBjruuZslab5l202WpVJdxsRe011rvsNNj5P+g6947QG
4bdTdPmX+1ur4omGIqNTlrK3iHExYHyX2FCwydaEZ99YBbC7crjONNCX0BATt122
rvwswPDr1CL9L0Z8Gt/8G97anIcp7qASqCvROBMIfgWKwtDPZ1v++qxynJk6HLh3
1zDX8XClD94ddbYTJ3CTWG8XBbFYHIViPKTE/GgjoWW1kIXMDIFAGLaa6xIWZMCH
7181SxYk6VnqdkKKDTp/eLy/0O/lBBBQ1LzxHAG0+UKHya30C59XfTZaBKF+dnHL
8dfdnGmhApPiqVLgnRYwGuxfTOy0VDCsrKAFW5B7tzpCmQS2tKX7Zc2SW+jQvYI3
OM4oYklseq+LMsbYggVfbK47PFFcq/GpPnjhZiNhZBF0XKpIuRqIM6PtKGfYZ7yP
2QUa8aDdfjy7lfbSZmj2wz3QpZavG+hHv6INpqxKITfg+RvTWQhD86TTSl8tAZ8k
MyEaPKYVVrybDRMCFs2oKir2pvr6NQoeamtxV+CFJ8TZndHvsZJamMxgsz3XPdaS
dAAojlwMRSmXU2Ohyn8Nxcrse9myRzR+PpVuGqWNr/iOixX3jJKe9QRxQRALL6sY
nBUZNdFyMppAAfmks+XIIeFAYu8Xr94S9ztRAug/dsDIpDDUdW4XZX185V18z4eg
RJ4BFkNyVKTn83j04mISoXW3dot/q93sl0NB3u+pFEhAAzyG3fj19sKYfRxSNpav
yU5OBgIeuTqaqKPvQS/wE27c8eS2yz4BTokSCsp/ozRbLpD3wo1nH7/nciQxdVk1
lRDb0+U5NPbThjA57lt6u0bauNde3jACm305hjes57Koq8p/di1U+lzKt8Y1FKz8
biAMrv0KljuXlDQITCuyTGDsTzRohZ3w5GsSzMURID49A0tYa6ZovpSCaQYgx55p
2L7i+zg8ZmGXUBTbvXUMBxIIUZQ9NeDcSBf8NrHdAvF1X1Gg5BbgUkzyj3xr9dRR
lj9UWJ0ZMDXdg6uRzGgt/42FFifUQtgaWTgpvlGi1fN0ET3cTiYt+Z5qA1D4B8gO
c2lLXsdbbhpyql/juQ04Fp7/zumBoDu7xIIn4VO9SOQhn44ay7+JuldNJ4l+HHfH
uCMhSKDi/0uk9QxqJ2ktKLKL4Y/x7AgggaTGVy6ULuhj1kzsadfpnMxAEkYgitVJ
LbAXPqG7nniUU23bts3nHMSQlU49OGJeSGnX+fxitavqYDZlik/bSh3/PV6NS2Z1
rgMaQD+madhIty7NAH1pIHIH1UShsOh++j+SSY2IwHF9z8N266EEwmtzNiByiecR
X6k9rmCLJR8npPJOR1UiVXviCGR04EoSK0cL6q5gikKhfpOL1KoYjqIJ7BEOqB2Y
nbYQ5m44ffh2kZPO0c5mmv0damNMskVTSlOs8GTBEO/8B0i8qQM91V3anZ7AG6xX
IK7+Jv6TTNTJV91F4BmNcqdFWa0ShHzUJpXjl/dQAyHQhxKetKUpXV4NKeEv5+pC
q1zhemFONvpu4jVbzIzQv7nLe+q6pw2Hrf4Ul0FCslyGBtldMx7atX5vLTemycyJ
9RsbK3T032anMV1v7AXJ+0T2SxmGE5ZpUEl1muxzpdczqmIgQLDN4xauMPT79Fp1
VZbFljYdxZB+DlaTD3Kzd1JD8U5gEctfSLQP5BVedOZjcvk+gef8QbM11GCXphtu
HwzRmsEwBJVAMO6MT1aeriSRaJtbuW53M99hcLbDF4+Yfre98FIW6b4eT1awuiNP
kry7K1TKEBeIKPyF1Le28yA1u+uwkSsE+r1O8qQ6j0ydX7RN9aRTFldb4ALMmdUj
isz2u+0BqBobx8yDqFBnwjX1J7tpmYuli39YrzgiV5/FtkB6Ue6MkpC+GpioPG4O
0/oEyoLa4rKaEV2wAdRPF3+tRIFMkHbeEdvXpyzqHMBZoLxRsacs+E4Wp4oHUUPw
5vPb1EPjPQHEZCHFY7ihMhMZw2tmSh6RfT928OuY22sR4aPa3wF/AOz83dq4Irzz
rHttPnej3HXEt6NFI/JQjZDB3rs2AT1vTdUyQmibO7EWQ21a0SLOnKnspb/cURWn
wRjqKH6xqw3yrbx42w8S46tLNeLNDdCAFTuYTS9QcQx83aFwoWQEkw8V/HQU9YNB
kzVoV2FdzoBYu/P2qPVF6DPDNn8FqAzS1gq1t9LSzvGVBbSCT/EzisOVQC8yaxJj
uoGPh6IgJSMcQf3c7P/U2pTDuCc4e4cTujgkxmRvEtvcFkJT7d4JvqMWTtq1qedn
ejRL5VV4wtmcBfumlMJe/9PMiOKt49HinGVYZNt5CBHFbuYEjkn4ImkCiGj0QamO
etloYQuOO+rwe2N+n1Tm04F9F7nZl+YnyJeHaY97owUuvROFMnLN166EjEE0tMl2
DPXpuocp9cHWmC4lp5CJ5bSt1wYDBkgMt6nH+e0GuMxGQMBYfvvP4Gri0pPs5nAC
PCEAU8a1QkGZPP5tp1feMk0SMeAX+9a+sI9NnGppwW9X1iYBrjNMDHsz+RlR+EIU
tuF6fc5yYGAnp+Z2uTX3mJVrzKeKgjw1seIEb58XUwoScecl9gQCRChwvzPaCmbo
Q5+4mEUq4J4qhLQPl/tnpOCp+V8/6RtZlNVE+31YAEEY78FbcZR+MX3VlkO5eJIe
uB0V0MGBCXNq7DOpSDe6O0bAV34dVdXf4Gh8jMLIowC6PqD0ri0hASczhqMcDQYH
B0MEu38lK5onKt3+pRVdhsT+IBMkXVsTXHQujpcMQrdGju+VTWq3lgjYrf788L94
vXlWe17WCKsFAj31FZUjyEubn37UNJGIA4SiVXC7niVoeCXr13JjdS5ePTR6XE0O
C8Y5MxRGDyYA2RHQfLtJnpXE8682VRcbitxFUbSDXa5TRGYktwPQ409/nHSKy/pL
bjSHs4AyXsHETxHSOdzXAJLPz9iQ9sR5Gshs0ztHhsyKb9W5GzkUwAyyo40Wtbqd
s2xeihueEVF/Xkp1SwDOtC+wpW6svAkCoDh65vLNmyk8yZDanRFRFgdcCb4kj1wO
Mjp7qkBsyzEJjq/Kt0NizRq7MIkz1OryZ9T27TOf8vVygI2SFqCJ9JmmjENvBNtB
iArqzhnbwHDiL6c5Pq8Y64FHY7y1z4JfAzPtNipXD9BwWQuaUa3uqMc3Hh3dIKaK
gEyAKQvoHZ5yRPBg4h6vlJ9JssT9QfMYa/Wh71rNS8dzd9hf39Mxwf20qCZ3pU9q
i2ES2KGA3MzhZtajKf2dhA==
--pragma protect end_data_block
--pragma protect digest_block
5OTfqjji02U2iwG4xjSBLoqdMiE=
--pragma protect end_digest_block
--pragma protect end_protected
