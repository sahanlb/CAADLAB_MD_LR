-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
umnACYN4To1cw1fhoWFXFP5T3h08ZFw0tUBqb4EGwcxZzezSdvAWMP7yP94m4L80
bsLyGnOWaRAdYMZ+3zfzyLOEkDXCBYLYdp52DhScLsv6wM0xh/sIr1PGPMrai5qb
6EalkfZGyXK/FnDJeAKs8mOR2+q4R2Ln9U3COIFCb4AoDo2M7JATpQ==
--pragma protect end_key_block
--pragma protect digest_block
Ir8rcbFgS5C9Dsx5CyPo/qLR1jc=
--pragma protect end_digest_block
--pragma protect data_block
ATxD+o3TMP9KVxvDlP6MdSBum3nZmJtt5FnRU6d7QZAT7UVywhMT/kiQEONhJ14/
RqT9w0bogHjiQstOJIpnVvv0WiySxwCewRdS8p9TjG7Lt6boPoCR9uQjkliQjc0G
H9AQKJ6IiF2lW4Dqa37BJrQnLyYwB/7g7ljT6/zxYIg6TIgZoC4DkXomrX8fMqq7
3vXd7NVUbDdfJxe5laPZCbPhjMCAZe5Z3aOJkB+am5wFeaBHypENx49SRaHF4hVU
URdYvXkicz/eRuILh0RBsMTIpWlWSCMKWGZxOKO5j0gHxrZbiwXL9UbCnYLf0Yva
PTjkkJsNXng6OskTMnIaLAph17yHF9CA5Fambvdz7IHKg3UypTdYXJWUxqzGeUw6
o5FkGhVoYMtSost6/m0nJwY7Vbz+7OW2yAM1lnzPs8LO5RIoMtk1M9boKMAzvwXy
rE907CzOnU9R5lRoQmYtP8Z39g6m34gqgBjrdE/NhYT8NmU+Y3SGB69bplALvpsd
UyqZQhIKAeoEZS87xMv3aowYAk+5g7yaZtjF6jKk2T1SX0xC5Lzyqm33h0Pn59tt
VEdcnkVNtbQpH8WKAjUTeZrzAHSvz3pX6Eh2gKWr2cJobMpN2rLNyqrR6r1XIpg8
/e6r2rTsrHuUzs2CjQbmEX+r3ItuhzdhiLGGGGAiZC8Mk0wr486WjQQqiuaAWlcU
/26+DFB9yXNQTScaIWKObmEjaKyj4MssERbGN69KFMwO8ociDxhdJjKWiU/sQq6u
VkqauZ9XiZXvRd96CsbCAyMSSrFusQLyfFW4p7yaYR9nV+MPzfeU1OR0PPaG2vYS
/rBEB4eAC7+eJehJAWbkR9pP+kbfzAHgs8ToUGn3Kp/7p6ATUfWhQV6MPMty0zbW
zCTuHLu1x10k4PyJTF+gtVrPe/437DWar5fxavJU+57ccap1I7zE3aQ3kYD9fwEb
kZ+AzHhxKJkoQM+HThRxNMuQgk3rgoqczJB/h4BSzYPdQ5Lo0RA5RvgYaSPQL8rr
cVZ0J5g1w24ybFfjCB8hyY5n94d1otFUV498fZy+wR2tIUx0fQ+Gh13b+L04qVwb
Fz88Xlw+xh6fqCd+F6oOEfqlnBOgRkwBZaC2ydSqkSJOy1FMITzP2kh5wnMFjUWf
gprcNYlXV3rql+NlKlG4UC8VBjcLz1svuHHq04YojZ7UPk4sfr3nendWnrMDW4/y
hF2nlRdkXFUczQCJvInEA/yMdBgX73xZEbelYEFgMpdVfCSvkUd8L0MRhwCNBRqp
Ibmj/CYR4VOD4jbxJjd1HOlg6u60zCzNjdgWZT70HKzYO49gakKtYcU3OZ2yYJXA
RVnZvccA0GStkNz1ofGHN7C8DvTOIh8WxNWpnqnlK+BrI5ZpnpV5is3vI7zI49JB
VRVxIsUxk0/bpsTjBgnd/xUSCALcOQkBkiMD5yCaCMnbw82Br9EyXNOk9hweA1Na
PrLy2rJHRxVOgX3CkMuHL3yZLsdmyPC12XygNjq/IhNVgvT6m2WypYhtjdY5xi10
lsESi32Nt1nsCJuzwbiUKB7lOn89CNIqhm/eV/XgWQq25U51RcADfPLSKBj5LevM
EjgzDB2B8oSDaKo/Tn+oPFWFKA+DADXU/qIVgznTE64U7oqvA0yxIveJbkiBGKyq
d9G8k9w6zb1CU0Ykct5g5wjkBpW0v7VEXATg/k6OlKvrLznskzsuuvKOJTDLuRAW
YMbpNEzASWrx3Tsqj+zU5lb49JUCn9H/T2u9A56T/S0vms8X/10fffNvH3/zfpil
bUOPxuBgkRC5/DXxG3P4RNSpioa+9PTvw1MGh3SxmRSWnut5zijpFnE7nlQCNW4n
IoiCAyUDdvSNWT+QamXBLLwOQV6DEpP6ZWR4g4KHvwOxMdjcZiHQJW0QqG23CssX
GUFFkMggPmv4jPc3Fwl0HJwjgLQDfS3t5WVRsBgDD/UrQ3JZ5odF3nry4XwON3f3
so3sgCfVm17T3PMg/PSQUgOARJ/AD0f/FjzmeEgMRrsYDYzLNIelRxsd/ds32gs6
nhJQGqgOgFALkod2kxTdyPPg2dfRfy9XVKPrB+VeN54mivg1WUPYgkiyQ8Whubs4
XdAXnNCbSfXPktqb1A17i1/CM4UMSGLJY8Mbls5oMqkClYI1SZAUK5H5oPZiKUSo
K67iC2sy46W1tl7GMvpo+wkCOIlHgA8X0RqwqcrgpsU4D1oycvlvoMuRXQvRf0rQ
d7m6WfBLZ5nYtWk/Z1n9SiMHxOPKAnORvGITiRJtEANETDCYgWSF4mhg4G+ot7Mr
RuXZoSzkr7QtTa7MmebGbf6BTOM5ONlj+Z0mCqoi0ALK+iiYwXKxcXL2TuhudiXH
BGAH4+OnJLlnAuYDL0OYUoNCC/RdVIVr/2wURbPKmHxz9ANWy9sUgcYiJ5TVyV9H
YnO++Ek/XV3ixNWPPvNP4qS5DotruX9RPxBCUn2vhLT2oWNXQXMqShaQzgYY06KB
shyvIdTLt2XtH0A2l09r8CYyzwtAe1FpUPdfOTap2LL/OWnQr2oI5IDhvyc8b0an
GDLElCp5sXgPANUJJLf3YJwXSFSe39OtGnU8L/d/K8ACP2dcVZ3/RPnUQgWgypSU
8XsBThP4K4KakGIPsjaZZd1mxgm4+xRs6825dbQMBDreoIyUjLD45CmLhEVn4Ke9
JPtkqJiZUGhl6rzw2D2TFe699SNeiXQ0j5FQDGZZNBxHz9j/gSurDHcN2ZQGHA3Y
qOflufvJn2wiMvhvD+6wTAagFat/zjMWKh7ulJ3ixXn7Do5V5oNRPDX/TQd0l2Jk
5ctk2wR4TzcBQHvngIoGmHUI/Y0FbaHBVPGUW9llZVP54wKJ8F6aHkEHbrkeyWAo
TMZ1xtCImmtenh+K4VVhpL1DTS2FKNB/rWBbl4e88K4W3axECQWP44v6ayvC0mxU
9T82TLnvu22PnwM96Tld62lyspGwDecAaAhnzmW6W9SCrRP0ofszVJOn3rlLoE7c
i24Ud2c0BVh6+VmzoqKpeQZB+43XBjggcVaRdLEGkpyycGQ9qsoyQygEJeLuLldq
vP7jCUbLm7gQMPBwJR0J+hsprQXHeJWA9iFQGXckvfhtCbDk2C47GoKQ/zqTffLp
bnaNyebQzsp8lS21pCtJcIcnCemt1bzkpEFgn19R97gX3In3Fr6sn9ne9I9zanFo
Rr+wKf3EFtAbSFO2VlP6DuIRC2bktkErHCucdm2YvT76EY8Stv82ErNYuXR7vPJi
XpKX747yYQ6KrJvtM5ScLLdX6FO1OU5sOofZdIcE9LXwWW3SLxQu79KwDxMcMSfg
y+SLoA4AeiWP3XQMq47p6PlsxxJHXMrkrB7E/zEM2wlLhB6ssHvyKtpJkV5brisV
zW/TXnjSy+aX7Xh7mot6QmuW5FPuzQ1j2GT1e6ku35SN65KUIfjVbcRPBMqonxMN
779Nyqil/CWErsVxcgvklIBT65teMN1UQATSSMFwZT+Fh8r90XtPDrIgWsPuuMVi
QAui5bxRaAjQ1Gsn4u9/fnVjAfKt/9xERyhYlpkJ0EBp7wpjX+ZW6IAJw5q3bKcn
n2hAm0vN6rCAuRch3m8GjaxBhsa+I9/wSbs4wg1/P0iK7tn+sDj2seJQHjti8mxg
oHVUxUUpe2bQnXKr1sxe4tvWUjl85UK90J85L8zFSF9D3ofrsXvrgSHnyGrqAtix
4DkHAOgPhqoWkrh6O8kxV2NZoABf7GQmCYNNYNjAW0uW23YIeKlpXYkvVBC69kfq
WoGoH+iySrqE4PfSEvT3+BHhQ4oDweB3K2V8ARTNrVmBi5DZ3olNjQCcWsjBFk8y
hMU+gaz4JNEDtqVMEgqq09XwtCEUKbCe6PDG29vEXqn6ATGw3uaSAm4WXe+D0Aqb
sq4u+9x1ify3eJv+4Y1NEMNegVNMJ/u9sHi52OV3S9nnjvw+gAFndbA/NniAulvG
vMRMkKFB45gIk/WUAzntQjLKS3MlPO4QZ+dcnArnMEwOMThFdm1P1dvG0ROMtFSP
gJiXt/3en1Cp69k+o9iHomgj4XqyReSms/X3morqLrVIbyjZ7g+/Tyr7fcmy0lA1
UNq5ChkhtCrx3EtIrRuGiYBsKBWjaqogW+bJbCGjIwhm7nzJsFXDj3ZQCuUiaqgf
QWMgY2/wn5Iw9X/GpbsIyN1yBvnCS8gNeF85a/AMQKLIZ8ovyQchVTI2fzZ9fqpV
2ZsxN6VY3HPe+rgOurESlSY19+EYomTQM6ngPs9heb9rfMU6XZ1Ulk4CDxIW09pz
jFJiddi6AM/361Mx6VG/KT6E8a+kHfXgiO/Fu6L8nvZ3Foq5UjJ8nq8NcuQ3+Yag
1+R3KFqN1NMshuYwjDteBx1HIQAvBnEOcX/WNz4J0N5m/bK6MJGhJyLh47eQlz99
gkZRWvosVQJvT0rYkUL9Dsp9XVUPtp/URBVcGnIHXy0XowZGeoGwjrfPgoTl0XqP
4doQgdFdu45GgAaj7s0a++Ao0QyACsomwRj+MaW05B1KVEFKjRPCuLGxpFg9iRnb
Zjs5zSLxKCOSwj/JeurtHORX64qhStWvkan1ojcgKK9gRL4vD9/bxghc0lBOED8X
AYSGgmXmiS1j0HYAkQ00IJP7gI2viSG2eq1EHVcE21DN278q0OKz35Y0ESYtuQiw
/S4+BLoJh0wCPHkFvxDamaHF9dz4Afb3BCAquJSdF92tIMh9JwIBM8tSjmgsveeT
NQVqsGfVZK+22qDHouQhN//YHtP/RMBJO1egtVB8b9nIKUrupzRSWxW0Q9n6HIM9
V4vzFYGdvc2LIsiUFr0wgb79N5oiu6d/3wwfz2/FEAW8nWY9Kfd1wWAVsNacin5g
ibP5LwaiaE02fohzUbbF8GdK9iZIV5hXw8Qgj287R1IDLHjutsc1Ok7VoWvJ0Ml2
/zwEdSo7rOoBk5LgIc6S4OXYiDV9rWZBo3KtZziawUyFiIQ47LLGoACBFa8VPmdo
G76JU1AhiaZ4YIH2u4zX/trhSEou64TxXbdG6VWYnYuy68ajSfRCzGNgx/ch2xES
Qbi5a2ZPJruFtvf4YmWAIaFNmghZtjiPPteOh1zB3tVGT+TVaJpbQIOKFTaxPmfV
dP9Uyx1WtAmsorFDf+lN5mljKt9JPWID+TizCU9rzud5QqzPOMVPrXXzWRNtQYhJ
G4IxkMx0PyDDRlOCz2f9VQmN1Ey8XsbLhpqwxTcILdGSbL3M/96DxYMs3JrM0CrS
qLi/2YMALLqMY38hGlKo/q4iYN9IGN27xeEGTnJhlP1qAanzfB6vhiwEwpqW2Gge
taCUAX1HvEyjpBIprP9vQAPEkFuj3VEsfXZSgQocye64tS88Uu2GU6YyVQx9MLr2
MFsTZqP0Y/bkoa4GINNPNRraFgpkSF4ED12OHNCVxfdj0BX9943f7OAOHEjn7Ghx
4ScnlzWMbOiuDLjvRBCq162VMr0emfMIfJVxL6aOcqJcpp8+bCdL+jmgiW/tzhXu
5NxemiHcrIOxS5AfcdGhHlAwH2ooVzsLNPrGgoqnsmUF7RpKtd61Pk1W38RI8vFm
b3WYALE5AfvBze3TgeMkExwlxNdyw1ma3sos0WumCwew5MG6UInIWCkMsemYm4ZQ
MeR6fNIzZpA/xJdBgD+9V3DPwqc5MWBvV1eU/WKS0Rw+1feVMHDzVOwiCjQgTGzv
GaHk/8UqyI5Xl6vvrM5etCF5daBx5pl2Y9BDrmoOVuBFtpkE/L+hJbLz8ocXWmh/
dIEgH9ioCEpPYCuMlo+oIXc5TlJcQUBBlN3M+sYhj6juzjS9m0QlolBPxhV41XF+
my1wK6w3aWQuq3YJuwkXwLdEQqiAHrPl6RART8uulvYEbSSXOy8+/1q4aoqGzaeA
nEEIt+27tFxCwqxgUWeA0XyW0+QyPwRM5SO+TFRv0dpNQKiE+mybVVV20eaBAjyL
bYL1zVn5v6FvKAYvMARvvpgRNCA2l53v11Obk64ucaWCd2kQRGj9k9CRuwJs2X/X
xBK+32N0gykoeMFvLOWhfWuP9heRouxZ0laKZd6R7oTU6NnAgp4wPZMSjv2NkLgE
jF11gWnxGe/qc6YremNr4NlXKhxcm+X+twn1d8Smyzew+nI7eL9kZuTzBs59DxfW
dtskqXkplmgWcja4jwRBMZYmhAo9ZEnCRdFn49bMjyPoQtEZ3+yHrzf/pIxq3L6l
wpkh/pRJLqcLgEqyt1vZTMvQOE4fI6gmZ81mwvMgzB1cw8sspdZxn09tzp50ZR5D
vZpzyBjCDeqZ3ZkEEzUoWJNObjpRsfFU810n1cd8eIXVX72ABn0/0+25a8i5fcEw
2DCwJj/O1HKk1Ykq0Wajiti8wiATF0X38mbuqlOsMMLHPd3RENjTMWIsgOuCxiZY
D8F95wYNchCzkUr6WYQ8Y/u3rKvYaV+xV6ZHg8gTXnS7KQoQ2r4cSPihtGRA1Mp5
K0VY7VxUetO4EfLWkb4rXF9Zk6hXONBEk9pqKMPU8ydp4XIgXcXijp7P8a/DkXYQ
ydewnymz5xgMchfKDPB6gMBQaWwmcDBM2tZnS81DiBo9vC2gg2z1W3jHgVZCNSNd
zYrIy2AOr7h3TUuFEy1SLwI4/ecvL39nO5k7NGGWDrf0NoxnCPUjHBf+s24+SwSu
BEV29qvIbtqSwNUbwyWhZdF77BDb7tWWpWREza4yh+2b6/gstCdvS6oaaQ950V3M
2SRh22c0nZw4Q6i93xxCOjsJ+NgFw3bHtG6XV8ppIxE9GS25ZnRMSgJy0lBeq9ig
/xG6OPIj8X1xCHl7XmuM+Ha1QCUT2HhELLMaOufozo2OTcj/FABU+QG/YqTVBDfo
dNOxmIBee/Zta9Eqcl1f4/5h7/TJ34PhP2H9gs3WNfO/KPK2h7LApYX00J/qn/BI
2CW4hE30+p/ouqc6v7GRzcR0m+CGXrumE3SIvYrnb8MeJvcKS0jR1iewg4joKMEM
LVjXgYbGChurQg66HIpOT0G+Emo+1aDrRkYAhiuqI6bzjPiRRmqFN6lzg5MLkFd/
ckC6QAuFaU0BtLg0hI1eyAR+Hu4aCnld0XAT1DHnVJ3AdlVaCNDHxsvrVkeEwHOx
KfhhTA+KbzPtWK9KxR0BMQh154s+cmLji0WtRo1ArTUQ9iY2Dxho/HXHbzHcqc9/
f5CnLl+eLKL6ALu2kFnRkTMx1v851yJDJClWbQincsj6Hy87oI9kC943IFDcTblJ
dDAcGcMYGkTsK4jDw/csTG2iFRRvjGeaSKb4suqfjpAwVR6v+j2iLOGBhv/aQMtz
5kbYb+bTMJTrIDQN0Xt6ngtZZIKJyywBFrJeeY7JTuhwsbYx21JyyeK8qTOvgLL9
JgtWV0PRfCDWgpygw+1pc5prLrWPVtwlYFWzvO7XyH4YMkhpCMvXOKUr0CJlHlEs
BuV6ye5v2pgIDJYk+pQsAUsLTrCa5os7IDspA0Z2c0HsYEb/prHuvOL0bxD4C1E7
if5W7aKGnpQEwa0GfcUigAN/jhlvLIF4dN5ASgVUEiZLeplQzmy8QBzH9QaI6lWu
uiA+fszg9pc7p7A54DmU2sbxfznkUfW1NklY397AT/J6Ywmql5hPrQZGV8/xfiTC
ZKjaLba1TxKApHdQ4xpy8LovdguX0Nze0jANU0D8D3B0iGscgQxAUvuoLDkL9TkH
bgbJRX3zsDlEcapwt8nUyPegp2ynqHOQjPaaM7NoIjHCjxEWLQ5Nf6Dv0WPa/XHf
QnTBw1U3PdWomBt1TOf4DfyMkCsXF+FjgoqNRQluCXZX2d2Cjheac2H3iqvideAL
NAhtJvjgVf3mdGxywUDNeNce+XVm6Wk+AN0R3YACP9oxa8lWIwod37k2QTLEh5J3
mzufC1HWQbQMGQugSZOPPvCL9rw/Lq0Xfse+MK/d2krE7VznCw1H7hkGWh3pUkF3
0Tks/NJLxioMMFQgNaPfKF1HlVPt5x5mGn/UbMSPyvGzpaQdNiECqH2hUwUEsxci
IuqvxZIn0nunud8EEpnzrKqoydUXSAfKw277QOUclrb7J41b3uvO9w0ql0GJpVsV
lr/c2vNOAibAf/EzWnUoMwTgWCPQCcTa1JveKmf7FDkpr1TvPKacWTEIISDyys+c
SQWdXFnWXRzn5CBmNfhwMnYTJIGIsNrrOMqMJsC7BMLmIaDMvhDdfPK0ijQ8G6yd
FjJSD709xvVWA29c6+HjRkeFjkVAqGK3Bhkg7CXYZjIjh+oRZ8CX3qmrMlGSdfnh
gApJoNQH0ltPBXhuODXwuKmGAmNopW1X8HNt+SyCDI+0NWyrbotw3f5tnOrMj9v4
mRwOo8v1mGJDAzpAKiDLA8BZD7pfpECm+o9Fff4vjCtfhU7/bH1/LaNghf4NeEzW
NZ8oLnY9aabjiB/r+g74qjTgItAz8mZIYBfeCnXsnNHfCCi+9/y31NfYSZd9AO1x
3dvkFHolOjxKp2uzK0vmHE3PhXLfTLQ9KAO9yljdSlGPD2Ce59Mi9x3y4eVyEc6w
C2Ia7k+DXB1ocL6FFn0iH19+F61k8UANtW9RJMJP2trLlQhp/0OpOpVRRW0u9VU8
eWOqAgadoVfeXNj5Dtqb9oJyjD6NrN+HlfeIXFk2QKDKKNcJT6+kwQrZ/kIdkqNC
X1ci36obRNJh8ZtUpriM1Ne42w5GJFYLfUAk7lBIfn3VKkYYmaYWLhvzKdIHJq+e
B7PewT6NlqtQgnY/htg2+DzACaNHovFukFy2fhPGTI6JeMe+MaPEVL8Uk4fX1AEP
cYZlhHYWw7v4Tbrzv41BTzwkPI1yvMG8zf0I8ZmWgG8UpIh8N9wq15ur+Wa3o23s
JkripRx4zdRZ3XQ+Yz7zUB/RZ+sszSmywUigJSonhG63lwWyMlmzxBsPbKedmbr8
MCszCprhXOPISSy15nAUJsCQHYlZh84ukFrEjbfV4VCdB0SfjyTCil5MAG3B5jOt
XUhberefOaaI+saYrEWt2IqJo/w8Ftts/S0a7faDrCbivxCSl0d05AcSaCQinEd+
mMCSaEIaSTlFryXjSxUeWryv2l4v4v5tEy7h/MGw8oRdE+pALH8DEc7HlaoNr0F9
MQCds22vm0yV39gmYbtxiO/yXqkLuXc8yfWP2TGt4YEuTNXnOFLtvro7Yqja3pvK
x8q4DLSmrvY+2+3N7DiK9pgqdJfdKIh6BarxS9O0I7SD62gxXwhcq9OksJ1dqVQK
Fv/NEyPawWs91QawKqP3j41GupIb2zNKd8OKuea1yOgL2vZJyiTTxryHhWhI0Bkt
ql40B16ybJzpnV8BM0JVSpoE37YZS02JM9dQRW+739sOU802+rf965+UrMuDA43d
PsA9+bB0BNaBRdDMKgIxZglqa8QutWf5iuZJJ4oUEBFz0KjEkMlyLBvLynZ5orro
OVkAm1NMuRs+xAtXyN1qSiovrRbrGljCJOtqgpGlr82JjioB5WR3qdqiMqH46wa+
i3KFIg7Q9D9PCjtIfhVCBIONn3ajioiF42E+PqiSBGOEi9IicEoQB5MAHM/3nAb5
Sxlj8HUqXWO5yX/fO+i1lHT0J0nK9Wa/jFaSqf3Ywc8YAV456EuCB8QPxYzxunlu
yacecQd5rK8JNREDJh+m6IYeyVKoHfem4yzMz2s2Xozh+3iDQ17SsGJZ9gnrYPUF
LJ87jDgWPW4LdqSsaQw0e/wCt7QGA3cxUqL74CFLA1kQYukqMfIRFWNAscp1IZ/X
73281H9ysyHq22vyO4+ml11/5TYq5NZmJr1ZsZTBkg9+Pj/EZj/WmhCC2Bn5LVQO
ZoKcSnqqRgPe7X60TifDDKLnDdKsKSmUMWXBniegnSL28ixCfKglffbte7Y15oJr
dYaByAwc9n4tWjKAUGM/0I3VcFh7GpqLh1adbn65DqOq8UTmzoTu+u4U0u0ducxA
yy2XR9qMI6RRD5QEbXCINL8g05KvL1JOTOR58Ela2nJLX4CbfadLq9fsWh/bTwZr
WAQJqZVxno7QFS0Q3hV2QRrYHRbekBx4VFAtWO8hbpgNCpiioGqFtI7B4tdFccdV
zJfsyrjSW4rn/xB2GbZJVWVbYpjGK7ekUGZ4eJ5SLTNZJDhEza/0hJ7FyeO2kKdF
GATjglxAcoN1RZRq3RWl+L2cTtl6HRBfjKcncJ+pDl8/7J+1/7F+ViqKnj4wgHSc
pstv2r2WEru1y1F4XtKKAXTAtfPWL4iBUhGOi5HIrvNG0FdtwLD0bbfhmHKnCjPt
teVXGzSOcIGNhNa+ss0wrpMk9rr4dyldvF0/b1iZZBfJOn3DZh+mYcyGrEhwTDTE
kfPNbqi0YPWyzdAL4loG/ku/7vFYmdpGwhU47qqlZvvNti1yrQqgS/bL6abjfVmo
oL2aOY0sJr1WopP0UZHTVneWP1a2R+5VVkn8QJYPB616lBHVmjQtNZXyS5K+1p+F
eOHKe99PIYM7adrYA1psRcCE9pXI4lmb2+tEpY6nqS+05J8TY5+m9d4EpnVyooRt
asLYA4pRkYOMNtnWRMoJo7yBYi2gUlqqkwaqmmYiKjKVe9hGE3OEjICC7ZosE80d
Z8QQrkSVqauDlAkSpvyQXAjnQrp3hhzuRaO+l5KECd6j+okwYlmkTMbRQMFVyZLL
M+gjIaIWYUZFN4LeOrWf4VSLwwo2QxiWPe4uOLqEkgZ/cgbqu1ziEiX912kIrZ9M
qz8Ic2WNuYRzAKU2ZMl6Oew4Fh4wXSh3sqjaLqhgQJZpet7rf55ESpb0NJWH4HkH
j65uPkD0oIkyeJYK55GKFcgT3S4NUXqNYPB0S0jHKIuG0QgccoxHN08RC547rf7j
D/z5eJCVxrYweBqUTM8agi9GY9D8Rp50k+GmeaP49SN1gE2i4u9/ADfgQ2hHaImE
SLU2ubMkZQbSe5YbBt0WcQ==
--pragma protect end_data_block
--pragma protect digest_block
zWzSldPNCYedMKlMakM7UimtQys=
--pragma protect end_digest_block
--pragma protect end_protected
