-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
BXwriPsV3tC0XxsyOv0j35PYg5Zkm+iQd0/dUQtrHT9iwWfEx/aEi4rpZMqoSK63
Koae/8bUPxNQrAJ2zvCFwmNGS9u6ICzv0GZtqV4feYeejMY0e/MrdQtyDIxJEVxI
beFJeFFCMoFuUQx7qWIPAqGmz469PjPi4EhplyqUR2I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9468)

`protect DATA_BLOCK
ZMSoke2KSSI9QER0Ho010AOtYoTPN5mNA5H4O8fijA++GE+Ar/lvm5Mai98GJZmV
C48Zw+tHRH0ZcmSagzYn1sS9s9Dzu6Jyi1TPTLkubrphEnkzOCie5DjWXdcTBE8B
p3/fRTGuUYX+sgUSvSjzW5A5ApeFRYX3sS//JyQtSYef8tbbEZc+o86CkXiG/+Mn
Hfs0MKs6FWVdToJbZM6Zie4qXn+3rvkLD1DYargw6oR/lW35LmGGFURZlFG0h+SD
9CIBNYUrXvzxmMOFiRxwIygNBDYAxOJkz5wRMNL0h/t0zptN5omjEtSYk8BCDjzg
ry6bGO0bGvCZ5URqUChqlSl2oZfm3/320efpk/syG5DKVluKY3PxOTzHc9f1ZZtV
QDmhKoj0vKDuBPAWusJudIEVF9WsLcB69VJEE+RN9Oxjb9nuxZ20mzYdHu9M361I
Z6cOEnlcE59d+WIcM37/dIQgZzJYm4yoVCo5XiF8iy6PV9+P31QCsu4Lxc0gYEYU
sY7GH+oe67aGDl2aneU+aZfk16x9FGbLAMbH/b+6oJ6cp6xagnHN5hr9DExL+0qh
qJ/uTM0VJF+rzG1Gq4b8jKD6lgfjznBXVxltAvqn/WJqijjX3WM7Tw2W6E+0N39f
wCWLAmIy5GUZ+gQ1zy8EQrjbfhNBj/8lKBkc0ujQr7nTwI/3F1x7sKy5W9XOSoqu
XWwxCclXHhrh/aKRSmvcr0XXSue/sKFTJQZZwh4X8womneeGrZ632dn/ES9rO1GA
3tL11m7NiWczNQpwz7mEAFq7D6sfXw2beUpvdARypg3X86f9cPLlY+qC+K3DuTDy
A/DCKTk1hc4YzdSOXK89XLutQ23eiwlPdiNa4G17SB4+9Tqs/fM1yU8zfXlMRApd
oY3nV0CsjQNsWUBWhTrlEoC+xaL4V7+LESDjMTpexJ0a/QtKITAdn3Oh/KvcJtQr
UC5a/EiJILel45AHH9OEhr7XuQ5aNx81SR0g1bOKcbVefYsUZWIICbVnkFZs4NBb
LWt5E8P3LWQnQvM3DhtwcDcp+AzSL8szy8uM4+No2petU4BRq2vVc7EzFpQeTrVL
IwtfVe+1mD4cLWHEZNmyDWOgg0Q1terY+oL5BbeKzrs3tZhl7QRxalsghatXdbaS
3rMSlojPSEE712kEqku1BT2BfF9p06P7oxWyloHOHs6P3xpCbfeGkTtFzHxy57D/
AjJ4xC/7lWwmBc/kWHiy5P3fD8Ch2HnoA5vN+Kwf3rYMx1BlyY8FMZg+W5ZKxJX1
d0TfLSn5eTWrqL3OQS/3gY3zdRBuSx79fX2ERb+QyG8wEw56fB7FAxFG9rQetsh2
wPDLaFbyAhxdZq5BBff2h9QI/sKuONLhMo9+VAFppaDCfT2sChTpA4MwvTZwLUFw
VWWJUAId6+lIKNVkQy76lPHdhBevpUrsNXHZgOlWmUdRbMgI8B3clvu5FrVLIjbS
/kzV07CgN2N1yUowlyCNk28lXhgX071N6Hx60MPY8HlM/+3oHnvSKtGUT3OMpBF7
mqymQd9Fss8VlvYMs4slqf/piUoZ7wl3YEkb3n1EFaFQ/WjKZzO4SLsOjcYtGs3U
XdWhu4iCLZ7UuAwh01FEjV5lAOlCIFtN2JyVLWYJMgevsC5L9lEPtnY4+BBqwtI2
BSPOeaJIFWx0JNFw2/yJJeptAsYnm+daArjUw9oHZo1WjIFKHKC8+cvHL5OXMfI2
56AC+QxcwXsP1SbdEhbMo83P++iicqKV+LVSsoBBrbG5cdPmjMqdBpVyyovQ4U/q
Ju3/iSJOAQLiVVkmNnXNEsvysJAa3Tn2ylvuAiiG4MhZ40aJqSoL/8TGcTiNRUhf
HXCJ0d5SBUU6Er4VNRX41/VURpOyoTe3WwwSpYh8TD8GFCHBGZUEysZqKh0D2z13
IwCxyF8jMl5WVgkDb/MrKzzW6mpadRE2c4PvlMFl6OAXkLXZ8KZ4WaBi9IUef48a
9IG36ZU1MPJ4N4Slgo6+Im6wY9Z0fB9QRsddV6ERFt9+cg50JKb43q0jYRFhQaOS
nu5YJG2xcg4Xloi1pquRhVGTRe7Wmo/K9UeVXmftk3o2M5k7WSg1rtw1tVnYmeh3
+8NQ3Y/Kb/22ANUbRECBe0aPGiK/E6MMazwW56HCVp6YpuXaXvSKqRqiV8EHbkIh
UoVJoL6J37G3vvUIONsYt6I6YJ4ZAEhYBoHjNLZOJG1I5EWAqPnKDVzBSxllUqDw
joHPz/dFYURju5XgkO1Ky3WJIZi1CTlI8jWjDijGymhkhgTeh9v0zxRZIE2/BCCv
uQLD+YGkW/SePDrkspd7c/o/LyQ8iPr/ee/P5LwU1KysQ1cxkAmd0vw4q2kUyqX5
hboGZYEQMzkprz0c9n015fZs7RFJ/MdiNSRnsR4bJ/JrhLe1p5xkvGoICiwaDTGx
rCM4Vs4Zz31JRHWLlxe1GH4Qr3rLC7ewfET376cjtro9z+f9t9okOPY9WO/xdvuf
nmXrdYT0rWaCyVv5RPV0hboAb8iHD3LgoI/6+GynOaPBwUuCIFbrS5fZoxbI3mz+
AGs5lZ2C6at/eloXdO/lKLLKEAAhOu9/rTtp1RferXHDnzhkYKfuoKqM3C4aPg57
AOqyPljbG76+0JpvF2E/MUhBhM4Gcx6+UQ5ggnsqmlEfmssCtTqrqnZDDY2KzyZZ
+RbVQJ+EazlGSIN/GHk+ZF0xYqkx1kW+neEPVa2gqED2q1HYLfhI+pkXiwbH/5je
WYJWp8veU93Pc2f0re8r5ufYmHlBXALEkY3nDSOQ2tYZplS4S+AGsy/zHrRAz/L0
pnONAZW6pRwwYzJgO5jRRu1ys8uweBtM5UT1kqODxLRN43210ej53fprObfIKS9H
CYUGJFqVhVqGK4aOebx4XNOuALLkUkIPDXSHkAVT5T96Xh/C5tr0LILuYgbS7/aR
gTYdE70No+fDfH7QA8wD4nDR9NMmdOFvfQggeLzHQ3Uq0PX0KNpJTiuhTqcSHQcj
DJplIlndgMAZXBGVDuGa9Rq3WMhL4dkLDzH7Bro1nMExVoBDZpUYNI/X8WL386P1
FTrD/P8yvgAoNtH8mUfdOUqOY5f2z6WWMlYYiPjR8W2wE7kycA13zsbbn+hDTO0n
zgjNyC0Qx3ZMsdUonuOjt7Q3jA2Vrk991iQGPU3jRqIT0H22t+veGkzTKYs4o4D2
25sCe0I8kxBbijNBEXpCp2H4icwduEZnmldVU3xg7H3VHDbE4eEq6+gBUfBBcy+9
Dirz9SZCWqYwEaMACv12Cfkl0rTd3ivv9sloFNanf3UPv+6OMiegz8b0WB1+XKi9
H1OWI3CLl9AKIbNScp3ZyXS4HexjrKfyLlEt+6fHqPC15/OVUftdLHflwXMxk1tA
mvfZmuLDaT2rWu/zoDs9OCeGsqJ+Jyq5xPdPC+jwEQ7S+2+HzcvZqqAdIxq4fFye
D40/ucqyPesyJjjuPIQCpD9zedkKq9D/INjoRi7T/k8gNBLQFxJj1+AxGGwaT2bG
gWEbRvb5KK2lv6BHWFb2nu2pMUp9yntyPwFtUSLRSgYOC3ITfNuD3vu6AHQ5mBYP
2erLlcJHA2kiyX29wcOR2bYGnU7yVidfpU0IbBfsg33CXaOMpyPhLHmUUmqBLAgX
Oszq4eXgIU2DBYzb/+bAi+5Qxa1V60hsnxlEJ0vmuka6Wjc7pSItYQzEWdMssyJU
vibe9aPVTwJH4TTX0GgPws5dQBoJ0sE7Q4LgSlL53pMRqBKkgheArbe7rJB3zK4f
a9IGQmLOyQMMcFC5bUs4hfukvy6jnW4PEln9uzuDbZdoHgMW9/AB3P2oa30+QQKs
3N1aMP9jd2iD+CpR5WpPlH381S1coZaKHvw5/Yq7QH9trMtJgvtLwMCrQra9uiXi
Kw4acafqAFSfzcImryOzjeecIlasVOv7FzrvR2KP8DiLh2gRvyXZMpiAvpIW6lP0
spL83uRdE8IofiMdy2eyRLu1RTH42LJPBN6AV/6EdxHcHwtwJvaE4QIdC9VIFyDH
Vdqci7FccVV+Kl43NHosvpk7aq2VGKlez8PnzqAm0uQoeeEvctCCz1N/i3mSErOW
uVj3+XIRVEIV/pcHTNHv2cK8B7kOVVR8m3m1JoojAcH8nfWQPdHUUPcmi+JFgGyD
UPuae++Ts9D+awgdwLbYDttDOC+QyYd2NtFxp7fDNZ+cNM35noyEog5yczzBYBGA
K/VmUNxuVzkwzcNpddiTVhHP+N0MLcyjGSiT6FcgMPaez6VHptAT2+IZ6UMlKXy3
/Hv0t+b8RZoYJlz8zvHyG/C/e33mxCzsyzlaI8+YvtQBPohKWgG5TZvPbW033oYa
/wyKLZzDuo/KSUXaeoM9PF0W2kBeZjxJ/ckeikIvF7ssjmKWM7WbZkTsWqIUBtyL
csJN7tJ6wVXt5/qJEIrMM0Qsz0kvf8JuRCVCTYBo/pEx045gEPttZE36Zfd21sbO
4DZB9pD5qU2iOCZpYBh4qLFfqlDRj7rHZEu32/Jl8igtR4kh2SkNg94DnrNvnNr1
T+8qoli6VXREIPajruSQ18ES/euDIaX00VkIeuwCZh59BBcjNs+Od4zRczKDLDtM
bK9EiGRpICxmldlt6xe/7zQ0se14EejFqYULgStS1pcLgy7UQ2Zguyga+OFeU9nK
MP4ycp3KwN+grjZi0PWoshdJEsHHLIgyXe0KwFB5b6vfemXkc258smspcFy8/Yzy
C3RT8bbLxqOTBstTlo76cBwNey2U9fKV/o3iOVMA/zRs4HIY9yUKuT0kj9YJhKGf
7ZXQ25kx6ojXnZ82hDFbvFQdtEeN7xYFxPMOa1d6HHt4oTIq0rcz4X6jU4VGxVcy
/YuhOSkFDJJV8yFoJbPGWQ9ctP+BIKFElJ3kSIKAEjViCOgl9ioHAfSF/r8kAvBf
qgzdNvWLXdP5najghamj2EJdY7jSZ0t9rPv7+jKxFJ+Wnuv78YKJwgCsjxl4Hv0e
BCV/XPOZ3NvsImF/pEMwwl+DJ5fJSUj83l/QX8bVBYhbOlSqVawMH2yepvOIiIDh
kmqzJeHLFRML656weSsWfvwJ2s1/Rr+Y2CEUjXezlS3dh+VTnRwZwHw1lLyD07w+
vY5uXQ/nzDNirEjpYsShkWjacwwJSGeEC9dvWEE62XII+TnzRaSWyG8TiMuf2Khd
WthtKAQMaR+0N3eRN7MGLzRL4DyiaqNHDQJ/nqEbaNeKMUQaaaMLY9AdqHmY6NsM
4+p4IbDB0NFXm4qqIeSwR1Ke1/8Pyxj8pJCQbiSjFGZ7txgPMaU2KrOKmL90/Tk1
vzMD7sFV6hIZ8lbxY3ca2OHMENC4V5IMDW5D/QbHOlR1z5MVsJORXvgnARDwJFFY
LHbEn5XqPTH/kieWaCgpEOH6AFXOOeJl7VIFAlyLokJ8ghVFIyTj3lwFUJw+xgHo
ivA6Bmr9wamgLydGNF2HnLjLz/likmIwVZ50mwTjlSHVVSWBUiHsVmmu5hqkbiOo
goU2i/xhPVClH3UZVKcFsmxQoQoaxVwu1CwT81xKt50fZv1VULkrkTZuho0PhK1e
bEZZsUStUzVTjWGasiMV4Z4FrznHvg6dmV5XHW74AEqCvNaccR2IbMIFwS1rMsOe
sU7QoUnZhjfFYk2MadbZA8UC2nqEpA/1PsrZd4g97fBD7VtC0v9WaLehasF57weX
znC/MC0mnZr0aJpexwVEXC7K1Rgs70yzFMfeev2qKK62BgubUXosKdCcqjMpmhDR
F47MT3ZLSNYT1udUFsXOwHUwspvUBPQgbKgXVvVS0b3FYim2467aMA+xhrCXXE6+
qmyRYfDmxwE4v7DUaUy0rNI/qKxRCsW61SDCRstMhHEriE+bS7phfuUoAHGozFdl
m6RARJ5dkIgdiyzypsrmXxV03g2DQO5sXrHKUH39+WaNlPvRgs7TnhaDW4M8mPIK
u9XoxdGAeQjre2itge8+mTe1Tf4NFmlrNX+hEHrTziOtDH+mwXMUWbp4MWt+sIed
Hj+I5f/q8cRifgerG3ED8eDDETvxnX1TWKWKI4Pf7Mfgztvv+pchq33sxvG0Yw4Y
RcwCUkiyT2nZ1KdCnuTw1WAcNWmk64mheeTCErEC7pY6FZrPDY4Nt9yBygtDd8Wg
0Xa8MZuBbXL02NDrkpxpAlYNeXigx1uboVRqUaA6bbsFF6gRGRLaaQkSbcankAk3
85R0jDvERjxu1GLqBYabA8vALP4CqW3GDJInqPiS4QyH9fq5OwO9DUrwAnt4tenZ
ybk6PMkit7C9rczpNGQK+ky9m5NqwAbuQGlrhTXNr7he2/tQYIbS0bztKLo7CbGF
ZvsrghGEq5juclGEY6Ccbn0DJRHP+b01e6HqOhOBC/fe74CiEWinQo5Y5cgwdi6/
waVJf3yX0nQk4s10wnLvWJ0vj0z5Txh+bhFffriE5geZzlZeOMgIgWjU5yY4FLEu
Pv5A5BQWxKvFpU/d6LcV89IS3wOLsskUrwYO5MgaEyqOxSC+RlL0BkDaE1Chc+j3
BmzUEXYic17VwOJz+A91yzjh6OnJgehJjbuLQOAhUgXR+kjztUoiEZxTpdO7uuc2
NBJaI6YYFyz4faOdJpO8jEJX3rIC1LEpqlft/VkSaga0vksIsIgpz1tN/TkkXAfz
88yj5QPUV255GY8f7AMQGYAoTI9RIPEYkcG6RHIGD9ieKMO2ZHRmOrjdCxaffcbj
GaX/2kV3AYlvP8mlbiHsMkg7DlgyOZHIgaofTkonlEcTCC95HvmFLRXCWNDP02mi
QaBULnkJqduuLb8MbRxc6ViN0iaRl/AimxxUTl5EL2kzNyezKcxld5l29JJpTrut
QPp4NVKzCIOFpRAZIqCQ/m4MEdB0YWoazrsuFtGEqmbBUQvU29PpGT6DWPc9HXp3
AeWTjVxtOgAD6Q8mgr4PUwNEHABrbhm5rUi9nbZHqeaZRaKBySjVLWNfyXUk+bdW
+XIecfX+6y2AzHEUUcV5i5u3u2S+nNqGtDV/k5tZSM7BOmhOmedNrEMYYNUaT1rz
ZZE0zDOmOFTq6ZbsnxvpTmJy9IU53d0scDHSIgzVDTmBe145l1rz6+++1xShZWkS
q0i80tPIMzWNgW6f18WRQgTpDt1JO/qzlaWgAQ+JhAH5Viuv7LsGr7kqF1lbKCOu
rbe1bYCVgQJmH/r7MUNW1u9jFECbFi5Quc3MSfq9+BYRhZDbgdOdLYWswxVf1WZE
JMK8ATyjwcGeDsPV5zpVpAkEjndje+Iu4OOl8CH7ZkPKAq94U9cllR2ffWMWlZnD
z+wG/YWTdLO7s2i6JIivb8v4jqo1+yopuYUkKCtUiFBpG31OwH49XSlFKs6VWHCq
mkwmdxM6xJ6OORb7/kL5IishJebHumdTAlywnGM1Bhju0xLtcR9M1P0G/gz0dPhG
8B/sZzzHtTksNlnwp/8b8tpv4xhO4Ye86seANfXlXkZtdR93F537ZlPUaG/bonYx
6z6HWkXKrp6XiMTlKv7FsCT+2yIc7j12W0VIiT4L7Fj+6TQ8s6xcquQ5/EFW9Ns3
+sodsXwNHi9bO7ArvWo+PLFPn2vCbmY2MyIJYMtxJCqw36foBjjCgADViQs46nRH
eKYdh00ZuzDnm2r3JxSMRkvTGLHczJVmI42OWhO8NzGUzjcbTOm3QLGGH2aNNntv
MVudRUYmEAkzNC7g0dLz8EnVqiCrlSEpd6nCw/oHI8NbbSR1jpd+o0srpqWk4KX1
P1k1xX5E6j5YE7txZhzj4yovGQHhth4bu5GLlaJXnLOeUhrEzBmevxvQmHVPMRxf
tAs6QPRXUxUj+eIarlTHORdLQNHzqmZ5c52lqbvrRFTKPG0Zn6pDOm2kOaSICQCL
xIwxlno4fQW9RaeBpKYSfxKGjm7DsYUMx0ORmi8O3nBiqnxP6p/cJKloOwqjW0Ny
XhExQEdtQrCfCNwuBLy1kCCwgD4fTQBkna5YSTzHDG6xa6vIkid9RscfKtHAIy/G
Zh7NAvDAvIU1Ii0fs1zyxwUed5c/KHmrlYAF0RqX/yfbahLuGQHHOqy/BzaayntP
zGXr8oZNsKE2S2ClIUZyytmE+9+eydbNfBQk/z3/4bWR5dWHJVAMzZhPIo7g9JNb
dgSIvGz3nHLoDNOTCI8fzUUuAk+XpotrfDbi1DgTH7CZRBton9gyMwdrcgpAZ5ZC
FI/4Zf5gH7gfzsY/x2xHF+3MG70H7wRNoQ69uAVEPOtn6ZODsrtLYATZdTV6A6hK
gwdgyLSgKPIEh76CGle4TiVRps1jcyCthryzFUo0ZSkWZmPWzbYfwNjARCuMId3C
kEJcmEtfjO+hGu/WrClR+Qqi/snkQ9P68rmebfY0Cxqf4I+oicHlD8E5zVlE4KRd
mFomhGg5Ha12O62+04gPjBszxaUvMmofzawCrg8M00G5EM9OfIOkMc7roCShJUK+
BPaHLTui07XnyKdR4FTWTNj7YqpFT72axbazGtY5YgL16ydmur15kmPvIWm+4Am5
4eOS6IyWfdNi/Zteb+b/hLdexj2M/v+RoqGIcySdLStR+ww42xvKkVPSXYqJak9S
3wRrpjR5uNcPsUefPChu+8dJV+3pvSSS/1BIrV/Tew+3AqyjbMhlkrrJY7ATxSNe
gE/A5apijqKB/tjB3OpbGDOnDhnPh2ok4EfQw5zV7ElasGi4DoAekdnIuxObUBVe
fEQt13TbkwKcwJaifWHLmUS3eBwSQ18m+TKgCydGyJSWApjyeK5xAV7VI67Y95mt
/JAo5BcX7IaN4OkTXY6gjDmfdwxo7cOYdDt3cSmh9Vd4A0YCgShSouWg85uRNWGG
8fIb8VfxMF3V/G5VSn8T3DJHPeethNpUmfTxYTpBYNIM5neJZsunKNdfyDvmYmPB
Aqmx1V65ShKV73ZODWYgEbTklOffsqrxBRSK38mX5Z0guBEt9PoTutAGmnF0Trvf
Wyu5lZ6CCnzKWF+QPuHUbjIHqDhTIZam3zC2Ja1+cm36uHv/L/IvLU0IoBZVyi5+
93B+DS8PcCa5AdWhEfi00jvxRzUcEzX1n+44OsnnaC7s1zJOamW52HHqT5f43cD6
MZYQMfv3xa2hk9dJ2E7s7nd5WhjZz4UJ2nKH288TL/RVL4obVXtWBx2sUEGVYuGD
12OaJzryxxo9eR5BaNcE8frgadxfq9HQmQfQMD1ZM7NXpdaTi3r5yboxesTJ+QLb
y+h86+93m7PTIX4AV1BxH3oywZisDhuiiuV/73+JTecP0tE+2DnLXNuVr4pLooG2
RXsXTjBH3ym6jpsMxq/nlIAFdJDhwjdzBGBraANR6a4AMLXo62XGIA01rELMMgHu
Au2LhA2+M7DvE3GSvRcHg8fh5yH5OlWexcZmzOTA4GhAy0ZpdYZ8mvo4DMPYXQnh
WOg40bFTXBgxfBkGPZ6RxVcAdnAzPUYUkbGdIjWP9DsgN+Dn6wsomBs2SmVTuFpG
1Ebg8N+mZC9P6Fq26qd9vsD3cC1Uey+wAaOp2gMLsLNr+xtcFC0dZBqUXdB5mCkB
5jFxlu3T7fwSEwnZfun0HTt7Xo+KPPXj+nGRFI9EpSsbnX4KJQDQaBzFOTm/L6ED
VLa1fDU93SsXnsU6v6TiHHL591l75ACHVslKkBZaQKESWctQyZCjCznUrGOkHZNf
A6bIXkqmfmjOUwfBso5qibGtoWTOBsoMR8zXiDlxtEd55BgHws+HtSATOhZNJ4TJ
fQBCFgEzCvehInZ1EqcZo/unIUA/7FPtsgy120ERaK4PYMctaOJLwmTX8cr3yMmI
q2XP4E8Ozs3utBjQuC7yn9L7tX23zKSJVxLW390WKn+IFQpjMfWJOPJHJWjQ+1d8
QaKUuCx6yqvOHTYhMPcDjRJO0NRoMlDWwLrwPetKDkXRCPquMO3x91SQNlp68rKB
96410XncwxNjVT4pPwE9L73sHMc07ic5KvphvHUx2do74tdsM4rEudawQkgzZ7U3
2gDlKMipQTlUG5ZghX0sVaovn7Ur5PgSqunzJvJfq4uUM4XSkWFs1EbBQtPiMYgf
Ska4syKsF0aWohSY8j02u6RCWI9CMr2QwEYM8mmzlSZXk2ARWd3/QWUi8PFeolwN
lhaOvdQO4NBxGXMTzuSenVOSu1XsTx86SFhYo506vG8IklbbdT72jQmDjnDDwpW5
O/kKNLw+cnPOH5PoPORd7+CLg6/UjLUgJeS8Mj3jc8vmf62GJ0jVLKa47lJH64MR
HtuLxZJ5OAhIs0+UVRc8Ib6yk2us/92lifEQbY0YVy8jiompTWg5QJLEuoqLVJAm
ZbThpX18+LBudLGo4EqpSWeCpCUtOaB15zjfHl4ddhgsZYrPd0W6xwuHrXTU2Dal
XZf4f0sbayGqKmH5H54t4PU9deCitpq11+74Bp/+kvnC2VL4sOSnKNKnNccUfTEA
hCm7A8kSgBD8gtsOZrt0NhUkMGfStZRrqmfR1ytHaW0cN/BkdYqH4R/6dgCBcbhz
9Mor1yWFeTDydZwLRZWJxHXIoqKQtCzR0gdzY0W4mHIX5rXtF2lqjlM8ueAPYR9Y
53gZ+fT4aShJfXBippmRhmD5BjgJp/lllVo747j5bHZTAmjsCsgnvx3YRh3DaxBu
7N2UYREgqNwN/rb3WGennbxY9iZph2R9zZWnnHTMllfLT6fzLoCPFzKy+anE76Vc
llEMvk2HsxFYM9Owhlrquo9hi9lQ+smz7x4eitRA+lUQo+zQqqgKs5qtrbG04bed
q7a4jwCGP3S0fYS9YcI0kGdYH/u/TZcLU/o0uEJJTw2DmCi6ik8f2Cn00WsNpcD6
uDVFv8tFt4EnWKL4CtwouB5p95FI3Z/CUDOSmmlTioyKbA+qSgZFNSMXKLCSgHJg
jY2SOqE/l7Q2vwuQNWZVgOnO4Nk+np25ZuOr+VLDpCyD9NsE/Qrk2alwQ1GjBuZE
kMmLFA/kJIj1GvT77ZkhKyWhUumrTxHCxS79BWPuUZuELDrD1C9uqvXb2eVqTrrY
BgoqO7Ezc7Kq8tVaFON+l9Zew7/2mBmFqXbzF8M8KJMMqgYg7YMxuVKq/yj3/t8F
5Qqf549Y9pYIRcZz5LzPNIWyGD4ldiap3npRydBkpO2N4nwUIHRoDhOVnwEE0QUV
mT5GUSmjWC3DnJ9jny0LPHjwIJOCgf+6mg3EeFej3Gps4UbRkamAMWwlUlrqNwFR
6R2GL0t20D6UCb0SoJQIJWmKi1WI3X12C1Z4WMREMk0tTBFDUmRMzvgM5LYkJlI4
EvufZ+tmaSNtUI/rQeP/ih5SmsnckEtJcWvmpgu+qdjkOCwUjQhEKR/nRw6XVCX2
6J186aPSBB+ONPIXRn8le98gfQXlm6R/TQthPHbedCrA7RYFdOXGytnmFYRxPzZy
9E2OKO8GKlLhLT+KB2zEqu1NJvkMSjNEKfeFcuCqFI93rqwhY35jc1XZcBao+8dS
X/g8EwCCmdoTuWgZtXw9iGk+Lh7NHHCoEozfEh3TBXm7JZxKRRkW3BytO3gAVrLP
UYCQI0+GRLLtI3pjv5RZ6K+3lHwK5SFMEmJa0Bug5IPllI2iViE79Tc9yCwWVYXK
txVTAuFVYdK9F4e9X8yAGCTeFvl7DLYHgE7GQK04yeJkbEDC2LgSEWY+C/r6Uu8w
9JKX7Bz5rhVW7QGVK2np/fWHKK9O2rFnON3tVgCxPYbRWizHVKJLJgeJ09h0Gyq2
I8wmxh91QrGbOy9gUfRIz4JrO4y1C7UiXdP4Z/X47ZpAqLCLmANwsuqQpB5NNTyx
VKDykSdgp4NPVeVvpBKWuXzfcTkoTvOMt+kE5xT/YhHLvp2pd7HVJm4U4R7XWSnA
Ab8+Uudc7AxSlSXRfshR7N/fnInNQo3hYPaHy9q9dMNtvooaAVED4nw54aK+AYx/
rotZtN2W841F9JNYKf0gkxqslxqd4oVCZceYumhr/cJuzc1JmpqaNiD6Egv03xtS
+X9/MP9MN71XUtT/msJzhC9u4bjGmI/wmjPhv4607Lpv5EyOJuJUmRYqa3CI3NAF
QWeury0WYZtcpJ+mgO7lgWvgLnFtync0AmoUcQYwt4P/cz0b/LC63T6VsaijwtRe
Z8fB38GSL/uzNKiBBIwRKZ/PwtZg3DAgOOKfydkd08kCmvcIs/Rkwmc5dd5/ZKRR
zBSfW6F+u99EsOBWHSD5HFNtl4EtL08gn1BUMm80myBMfjQteDj7KvSOVWhGnoIg
PunZPIBki/BtKAhb5M2VF09aR8gLH5DV2tOHzq7jBeo18mMr4aEXKkkL3DtZ/GkF
iyd+TzDAPDCpWZz7M5WrqzQJBEELcDV70d/Jy6+LzkU0QcHeHfiQaV5f7IO5wSQO
Dz/t4+pD5IuqE1u637+f6T+9ly/d8gXdWY8G6A+22nmpM6B2ho4yuVHc2p/gl2m0
NIPlwtk1iCsdbpmHDQQN9CRSfZqSgl1EE6kBaZ6ddHhuuNsepVrYpPv2gQTBqiHv
dKyS7kmoga1GWR1c9PRoDad9v1Maokab8fZmV9Gi/T0N6Hlr6gjWLGUcme0ZKFIe
hIeBoyeofCS5O2b3nkZ+d0V0/ddgGEA7Stm9MflVmXueKtBkb6NGuVfitQbSd/Kz
dMvEfo8vdbY0pUStAjGc1cfPhC+Xxji0LqP2G7PsGFY=
`protect END_PROTECTED