-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
GB3O4rq6n+U7L6M7zVXmixRxr/GccSqeGD523w2srfeTgcUuwRchVXVh7WlaDwx1
mUoiJGCLX99HPkTQUJfcaVSArazlUX3UP855efP9vkw8qyAqiRnQ46v6sgtjiOEe
FUW3iG4sEeVLCK50p2Y3B7yDFGTsmwNgfEZqiL22Hcc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 49792)
`protect data_block
fCVDWFIFGSNwm32b2czbe0/VVxsiXI6Wjq0pbXvvJCGOXSGATx6KH6/zxrSEogt2
Lm0y++yZjcBEzyOPg0NFSj9v6Xta8xx9sJuTgvvtyKCOF818vUh8P9Q4Go2sa2MN
U8D5QYZ8gLYQbIQhXT7xuwmWt7gGkL1kHlTfsEWpmFzjINuwRnNKABUStOFu/9qr
OXWl9bq8RxIh0GA2e5K9aDvR/TKGgq4+J3JrNebsDRoueC92V2EMawZBbG69uNG1
1e+gDIPbYx45iW4LS30QyVCBMv3SBa/2iz/ZHrNzID+absspEk50ESYADDJT0j5O
NgHr2m9CjNy1EMJQ5lPTsZ4PPTe8NAnF51M2ixJ4Qxv31VqQ+97FGsBw8B5Rl7aD
nXyNG7VGVA7toiTt0XieUKkIq8oIMXO8+RI/psD9g4MwTgokLQ1+vyRNeMthnltJ
dS4LCf58Arhzbl0/vKpetOyF23Gsub/VVKoGev9tTGf5I8yQijiCpy9V29Vhm6Hg
Fjq+loHwQ+OxQwUezCyll+etwnm1A99UQmVSirJEYyNWEQuDDSU1LwKoNmeoDBLc
X9pgX6m2xCpGGGVqusiqW7nkDmR6j4v+33NKpt2UrAJtvWELXh/vMrrD1/PgG3Qd
SjKJLJh3oIKn67lmAXdsSShIzIKo/dRb5L8yzyK7f/2WYyaekMQBcEGDiSAW0BRd
MUwOxxXVQsUYTEqW+HwhNmNHrjBBEN5Q5Yxcytb6m74iYMU0gvTtHeF75lbgHdQ1
3DYq/MJml9U0hwKhrQe19jZeja9+TOD3WDCmWZ/F58qZcbvA6v9Bc5e3nhUM2n/O
Ifcha4RF4IYylP9yYcJACzGJKnJNEHiQhMlCI1/4ViTwUXzSL1Fz+o39WhYO/VOS
oACqoW6+GvzUCZ5bJ0CmEJa/r8jjzHLmp6m+xxcn4wGB89a9DThceTunpLUvvyP/
6YJf3MkLPX5iC1ZmoTU85AcCjixenWcyrnq2WKcSbTW+QnVWh7pUi8WRyhGtWTnv
94zN6XABAiZrR3dCstPJxIdXp/X6F8EfECIfVMV+eJj1cbmzp0SRLwSSnhsFq0cW
KsT2X2i0s27r7kH6EDy5qTbWbo/rnIri3M5kRMKKbwVk1/TvGfPNHIfcbkb5/tbK
ydnrtkN2aFux3fbHKH+oR6sbTnxH7FGlh06E5uwnxkdcBNMOYSwy4HixEgoFeyem
/2zn1fT5WYhE5I3Le+w41kHm+6cAbnaEkdFvqtdQQQnIU/b8Eyy0e38+Ky2+09VS
Ibr4lD0PWtAPF5EoffF1JSOd4Hvln6qvw/YkYFhMS/zJme62v8MV24GSYflULQ9D
tKuVkkZwmkpz8vrjCnljr7jK0kQm5CPXEnIFb3V6p4+NtFgpodJUyI4syfiLy840
EBhVWJaLc/hHyYYWBpnsuWfOR9SlWfNG1ZzrwESem4p0UAcELrXCS8VdO09kkwXl
e6IdWWpH8M0Zn90V1yKPCT7gIbWbQAJk8QMc7P5EGJT+yTX+7aULUT4Y6DgRTwYi
7Sbrxmj9ysixa6/tMa6LiaOwN45mZ/VNFC33/ZTrINBz3PNYbNQgb8z2NrVIIJqU
uWSKo88vzK0Yc+pgKbrY7QJ5nSDVCfwbVrCDIhRDNqjuahIBNlkpDt8njMDxyu73
p0mTHrBDliuAiNFWXk8meR+2JzO5D80Id36OpdJMSd0J3GoOekq3aDhuoJkbpKba
nQdw2FehDqY+1oD8TO22Y1sFM7I821zzGba7x5XiWTEUj7aR4L6H7vmtlCvbplkf
/e8qVG1nGcuArklJrn8z5ih+z7nqtfW5Qjdx7+1xgDU2JdxCtxuvmLMlOGSMr8AK
9L/suA0jpi5nnCXxH+SIWOLFdromelPBZbcg0YjzQATLoBpkdkRoERyeVCy2cKrw
K9MtFfgheCoM0hdcjl9fuw+9ASd/vRbC9ZbmmJh0v/lZLgW7c3kZSVbeEJoQaWN7
DyXPLosb4GL2FXpzBkmgj9zlBwGbNNdNwq3xM3Qp7UIoir24AVhqMeWkGDX7XXAF
CEQ/6+k5UdvQamzhpqxUwgGJwcfbktcma39X1vcrNZToH/xu5ilRTgS5PkAw69SK
hF9XR3pQQqIirWEKiOWy9f7Lp9BuYNOtNG2L3RcVrcL0ivVl8mpVdJL0P5uB0Mfk
UXdMZGxGocygHT0T59uDiF45JRFApRp/MDCoJiLPFun2p4tBz5wduiLu1R4wx2n8
zZC8AToX3BwHmc6SwQ/wXAfez2zykDqusF/vuwC2Sjt/T6KZvDVPahrUdHLquphK
6K2KYK0xdRMHXapapEGbVatxoAGzb4e83hNKU2jBxtiTE/BXbGXprwcLV32iwoLP
9RfX3LmnS27VjN9kM3tMKkR9o2KI2VGYuDs3jWPuzRUcFY9tYEm9hCgBjNSpaoG1
SpFwwSDU7MgyKRmyJ/KxddGRlWD5hrl3szmrMp47dPQsgl7smMBnkmnNJdoh4mGz
AphDVtUOyW430pWMnbUzXyS3IG6dFlwZROeSnSFoi5UwF6W3qDqXswRy6h7X5IJ3
hrzpujlDxvNEsXlqzJ7rUDMTkEzEvdc5L8Kdry6lkNu/Ul/vdKv3bN6baN1S3cgU
D8ZxjJibvzQbGqSBE340W90Rb6jujT9Zw6XDBLsYNV92z+/dHQq4MLqfyVbx1JgX
0pIqHqGdUVfVBsWrNocVick68DLr5qyZOuxXu7r3vY+tyaFp8rUtf9NJYGsxDBdD
kAsJO3PK5KphRsjSl7jHYLqSpBLbIoz/73TBTO3sInzK9e1WyINSpQA1mN0Yq4DQ
dhAAFMCo3M6nF/wMN8TDoUVqkiiZ7Yb6s83JPZPQhe0f/GTiLUv1zHJDo4pqDqqx
wXtyVzT37H1v2gzQgraqkqMigwCrfTbHKSpsSQdYaDiT8ehlUHaPi4dtfH83N2pt
2Wg+JtL7E4Y6cv7HX46PInAJorAvv0ydDRG6viE+hpOVTKXEaLFnQg+o8bvVvFy3
04RWVZJYrIP3E19NeeyVy4BbbIDAo82JFE28zDmIeR2vo6VA7FHrnwJmOIaelH89
nlqqHIstovNgGBtax8o/FZXbZPPm9N4tGRWVo1ZcVMjLFCKXCnkDwPmajUBcc9I3
/CATxx6II7zM36pYQsxdSBNxOzSGV3wqRqO5ZUzT3qAdV3ApZ3p53QpIww1i4A8P
IQfkdMtODvfZ1aaJqRFxRx7M/FGWej20gLYWuTujJN8dBNfKi9/pZbvQHnm4E1LD
ODPvG0bdVCa6xeko+39Gy7DgKP7cpKFJdaL3924bFM4beSuqN8XlPiU7aa1IU90s
IRiFBQr6o6zUaXwZgxczNy9GVSAZeQ1F0qgDThYHME++8LkYnxer58zVavXgBgnx
yQdzApE9Fv2Pk71TBfuUbnZaNIQDrtg8xRNAnThot6PRcAsPrePcbEO8/wIh+jsR
32XJOPC1WJI1s8V1edZ2lShwVTMCebWC/NPL6+IGgTa04ncJV2orntp1UrigJ9mF
kbWwtnD3cxdTjlY4b9dQmGZyBS1uV6HvIPtQ2WV1+9slrGG3x/cAy2ReVwnUB22B
LQ5RN1/7NUrWkQ0eWc7iY+zxu3ARME+xWyp7+TgfzlmnHTm3SiKGMU5GdfeSulU9
sFHeRdRmZ3/Tt4pxFJk/821teY2SOnfE6tLl+MyR4ehxc0CkK+osbG9AR7v8aVg3
CkW1oSFUWq4ta46PF0Rn0ZSVyTdceS0bsjEn0eojEsR6PNNtoPnByhYDhtTFmK+d
vn+3Qp95m3hdayfZzjfKydbupyIzrcFUkzcNMDAK11Qq8ITPG+btXP19jC5uw1QJ
Goy8LcqLr/kdmJ1IoyJ+S+RmywG/4MGJfgvaLJ7qwcQMQtSnlEqQ1l879/Y6YLRc
OqhHH7sSdLamYMDSFSZThmGhKXsyCyY/LVbww3o0HFTe8Vf/f3ZI4c3gKFcT4bN7
BGBOD5tmoZ+C4alpEoS6uJu2frjoHSzRw8Glfc2EgyQN9chLssv42ScrN4y5Q/cY
9UJ7b3qbAlNwb2OvEgkTZUtaB68pDJPhwA03aXEdxM9XmyxUi3MhzGe8XfH0ngQv
p4WdEzfCx3lHU/McG+ETxdp1cImqb3CWNWegPwBVVTcM/UucJD2uiHinw/w0q85u
n9H8PrfGFo9IKZvMfSHGC0rcGWJRgO2A/6tPczRzJ5wrv02qZUh4OObp66HoVOHq
PMw+PL5l5RPdkma8xj4DKC/MAayhqfxoHaplEPMAr391kgFDzH0uCvjnQ2QxK8TC
f92rSv1akqzLVaZWWd3M6x47FG5wchR/kteMBmwm0h421Q9mhsaGZoHA3VDyvHr+
bzfjg9yTGk6/f8g0WLHtVoOFgdglA+DhRbH9js9MCcPlNHgjTiaY5eEmfzbZXnnG
3xXyhIejGopWkulIFryG/xb42/lMerXOLk18+TF/p/7dQV3Nv+GW0PTDtNrMOgbX
ZVYt/gt0TY3W69PmswJOAbngBP6LRbltJiVT/JtZPjETZIbt2cghLW2mdFdlyO+J
CJ1vTgGRpEeHYvt9RLX5uhyCnyyMJOBqwxT0Zklw7hd5O0MCmLDWrgpnNi+snxHT
5Jz1SRl1eEWZ3EZLp/qCUt94c2Fqq6nN+pl+AouhxQen9p8qdiSx7o1Lmztzj8jN
mVxadNqISm4eqsB+lZxoYfDnotE7yGKCS2zyjf77YqRBDXXtW588+RZ7Ni+VGC3y
k0hueIASvk1iMEmJLKGVdegRatNmDhzj/Lr6YFITjhfKYcUI9cK5fq80f1epKp2/
AvxMaINrEmb8FfoxptyykTtLY12HgLlM8jhGBOdzHF7D45fjhSxpXjR3WdQBoqIh
mbyhq+UKK+BJ7gvORaiIJqN5A1cEWnDWla9f0yXWU+19paLSVed9SiphsBDyb7c0
s2N+8ZBpg6EGrkiAkmUFZ6Z1yWw7M3KcYOrt8lSniHIkZjYf+oZpezkHvfNybcA5
jlmPbY/yVit7aAM3uE1HJLEpvTMpkMnV84d6GcrrHfz4znw+3wzhWpgUNaplYBTf
mPlonYKZJ2HalfGn+rsulW5FLQ9tQqke1O4HkYK25L0lKsZt4DFB5ZYYGOgr8UJM
4cyJJytsLOdQa/Q8mX5uIm8RxMAv8TW5X06jW/lw6CwI8ezs0oeStQzKrj5C1xBC
o55bY4+0piUIX4zBHxMSMdiqH77C1iaUwSDtjrnJ/hl0k5oMEc6zELBASxNwUd/W
HSxEgU+SnNgO2/MvkoslHNBgofaKPjTFc3oBlVgLYlQHpHl0i12aaxTlg8auTQrJ
/zoh6AxvE89K8QooYEcKV0QmSkUqKyhLG++GXHNDNuW3LZm9El17ZiFJpBXmYiFj
lsMuwQVg157sSvPfhYoHQBQwEi4X17xQ4X2EjvS1rG5hVSC18/f42H0uNYWGIixS
5PcyDCGl9/wdfDapBPDubKls29m2oATRJUPesC53rMBxbN3O4aSQqdTHV+pqZVuc
5G3tzALyAyFvcwUm0E9KnmiSSDTIvQ8c7LdTl5qwWDZu6qdHDI3MJpa8XW6DL4qX
TnRmgXGcxcM5r953j3E8wqaIEpdesiF5bbyUPuspX8kzr2oTYFV2TXsRax8L8Sdn
ANhU17mTC0AO/f5P7n7tUP7+x69U5yQ/n21nH85fjnwNcMwff0PINKH2oxs6KeZ4
Sv2ev24QXDmPncSaFERyECAy5GEhu3HaQiX36RR6U45nlZ15IRCMYpticpiEsG3q
5Jx7ZpqbS4sSgRMx+A/y2SlI8qGwwYF3zC7SxcPrqlTnxxUgCuKzhRVYUPdCfCxp
E9cGWQveJGTL3adNbs5NFwA/Z84shbphmVtu0hdaYCtzeqVfMj+66BFcwK8vz5Ef
cw28bltlOd3vUEh/8ienKBCit4Mr+rbsAvPpkC/7Fp4zvRqm2y5yJcVjl7ba+vKy
/D0zTfFHCnVI3RjqlyhOv8NWv3t8t9SCa67S5hkolqIvc/T2qamNPHx7+SPZP8oD
E3dN12TOZtH76fwwJuTIGVdmWgQMAOg5Fz6s5ZEyylmnyluRctPWUxVnliAjHKZl
09KhnQ/ep+SSoHbTMnm3MtuhqWANFpfFvvIAXyyx2ZWAgUixVDJCMMwh5AVY4Rwp
9W9t57NOZnm6SLqCvg+dNh7o3jZe6GJm/TqGiNa13RZOThJ0c3nWLbGII6ZR/A1u
TGvQtAbzuqDhATDR8ogmsU2Fl5TQ+gOwFZGa0iy4V760A/jaUPXTEzqT/WtFCp8B
IHXFpGMBMaSAtvUohletsC/Atxut61e2sCam2fNuRbdtQSyDjJ2Zc/RGkNwa2hbU
6SdvdgF1S8oIYFRbm/5NEG+kNPVZs6lwkrWmGql1aGnR7TGl27Ka+XA8llAAf0D1
C/2z12KLHVgJA5BL5DcZMbffZEuCju4QZLCh/sdH+6QL4FZ4N75QrpgqRrdvxncf
d3nQKbGkHeizwO2OukYVZgKRAQdMLlXkgX1h3dv63Is2LtWf9Ckp6Ch/uULX6sHH
RaWRxTFrxVBYP6G5TjvNRs1GMfpkx+AZBnLbs/3TSs6j5g+TD2eABn3AEsnPPLhN
QdN1YmdIzXApMRvKs6O17xnXykgDK2YplKWDTrMo417HfVGSYSgg9GPdhTFjZV4B
OUupkOlCqPOsPYXhiNwVQhvEWMmcvCMxWCq0jIVnIJpJ56WfhUskCAY2PBrVdX5i
20SQM1UYZ75Zk6/Kh3OcEriGwoHMoZ8oCEocjNxhEGoa4YTLIGTfk29EYh21OF0K
VdlTLQwKNi5uPZzIEjcqnok/pIpQtfaNluaczykAs73IU+HSI5WXpnq6tOjSaIsu
dwtq0BFWNGOkmLonC0qqmlpUfppqdL0XYLXP5g6pOowabFR8l5zg+qRSB4G1W99o
YuCCqe3S8QLwnvFuCWn7YO16xb/v+Hl5qT6FCFTp4y5F/Nt9SnA0ffy9VQURnJrY
SyG+OA61qvRsntgH7wJ941ISk3YLFod9I77kLdpvdza2p9LhPgauviLs+ZZefj+M
/s6J12h/CTih22b2raR3+J4utrLzjrXFZbN1YkkR7obs7Sd3kgwMacWQ3jo0u6Tn
gPrUqhVd0f5m88FL8hKGm9jJpUQ3iWlqKcIWZNKZXEMvOGpS5Ey8xC1x7zwSLDob
6fBGlwQP5zstOgvpIgjPnfxBimKa1+Fw/8SYTtKrn+3F+n+XhDxnRNU/hYSorVFh
pGgAmOVMSZAVoidrr0IuL7K+/tCyC7MiX0MmlRkZnANpIsq1A6hX2+SrV/u8SIkQ
Hzc9GuAVd/VMe+AtRb2FI++IgYSUBS/aZhIf2ZNmFZ8Q3NgVquLvaAPe5bBzmbNN
2u+R9snMR3HT/30UhD9kQdG5onYahJ39WHidny81T+gQrR8DYgqiWpzuwjBSqqqB
8xCFd45u/mOUh6T+peuVbYpXX9hW4n6UIKKIZIs+fcQx8Qdsi8HKKr0j+E4Suxsw
DK+68mx5EnCi06ZF1YoTmiXoWrjS9ALTbTItoqDre8k1PLjj+HqOGuFFAugWdtuz
KnLNmc8I7nWZHbVL58Wm+yXoyK9W1ithXUbV+JK6C49NISdwme/7p5MMM4BnqUre
UX/utWdVL3cORFQhOiMXZb+KcPwtBZQ0Md+WCKSV7aZY36yqmkOjRYgUceXrxc7a
iGthPEPtvxZvBa1jkJHSxAvVleLMHQ9Ka/S5nEcBqT/o3lJ/fd1RjWeydRnweW7+
6rgO3b5qCk7dwS8bGhmfNiLbnxgCjmzZg/4qO7+C/ikULtU08EtHI5SsUpkP6Kv+
BMXg21FrTfsYXmBJ7A8ZSJ9vP+iHclohOvdFeOlFPB8bR/JoEnNhPVTvmSGVgK+I
BlGSQDwjp0KpBkHMiOK56w7b4m7f65T8QezRjiA3Hdr/o3C/2MIyTXALEgtEV5UB
TmjomUSFCx70YB4SiqykfiwYtriAWNqRv7ykdtV2kpgoB337GW/2X8nRh7L3FKiW
Cf8uLx90NlM2/0Xj+oIkueX/mSIvcDahdZrrOroy3X9viG976XyxynV19YsYpK3l
t9fvcoMLDLQwbhD+w2TF7qJXDw3+OkulZc6hIHtEQbCVdnPBR2t8/QvnFL82pgoO
Cim7xOaFSIXuoJkFR2gZ8PwH6sG03tOuaEqBJfrFO1SpaawXZLMJfSqIIIzscJOL
BdVW8+5Uco5wApgstw12Lq45BFFpMNe1gYNl1jL1Ckqdlh7A98hSxLLuM3inEJx/
5KjVYJjH5sIfe90Vi+FiKslI9yJd/QXaihzFCPaJsVkBjpw9ZlNuTjnpIiYkNYiD
z/EzXIqHDNxliOPmjLfeoRXwYQ1pGh8kV/Q4kJiZWT/y+DRCn29XuZpwUSSfgodD
OMeZG9HhGLkHuw5skkmain7qce/PNl4dbmU0IG6toYm/2qoYeP9EpvQzVO3OJRob
RRLp6QagargP+mcwILoVQjTbXDqPAypK5kZDefQ8RqNGDLw/09ESDYr2x3b6WWtg
WUFseXkeVnaqVcNYh0zWOFEaPwQlqjN4LtSZFtkdWQpx3MuUFQ5/DMg3AK5hd2b2
cXAcuqkuNvqbLpzaLayRjyMCo+Mn+mJ9HAmBhXMnc3CGHihkca2Z8O66rqG72xTn
pNgy5YEi6JdrtukTxYyOoSAVr9oqJgCwJRpH1fuC+hIVGAMdM3+88V66l0EINKQv
qLt0KM3CE85DYZd0dlKRMOXCBrjb248YEzE/MoW6mPo+cZKLlnYkMJTQh3O4IYM/
wJSRnR8EV4Ve270DOfZo6xv4HWDgrIrg8YkQxc8u5TBmdPAWMTk2GMgkMp104gQ3
/D+78SnSFYTl6fS376M1cdC6z9arM1Lw7LSl+hnbBN4fgeQnVmAHsDSa/0Sn+DnP
4lo4YBsIitW71I3Bh/241E6olm7omueW3t1oviMaw0enMZugmXz5CoUSn3o6wPet
NVfxfIjdcY3qfWzAmDWMYV6R91H8rNci7w3g6oPx/lu/1QvD2Cg/vBck7XjVkvg4
qVzJw0kYYqPruzvZDPO/5X80hBy0UR+j960JOhGJdBGyF1A9XpzO6GZZvzbo8/OC
UMAjUyakGGqfwhJ1KwSgr8H4iqx0gvjKCJYTMN8XUMzReLuJwvusorxQy9NxNUXz
0Oyej6NiY9oC3N7DUhImTTXiQ6Z0/YHvJs7Hh8bUNiofesZUupK7p64CQNYONi0O
03/DQpyAJEaLN4TV221wdpj9GkUgCMCNDWkRsXBrEUT+BgZfdipaN5HXkJIOfJ8V
eAFwFQyV766IuPBN8YQAMfULhzS0cfqWUVDJNPi7MoUgooXy7JvujHhNEcrDh+lD
bZlD+i4EzHbXi8og/kCJzFS3p/aWSl7CPtF1Zrz+C7zfiigqs1vy3DrSzc65TNbW
D1RqPW12y95tL8/uIPgGde3VWBYto0CZ9DPCvsK2aZePtZZn1UpT2Z0gdDnAUlBA
wB8NrIBcPZ/PBDupdl/qhghPXZlmq+0FArhblQtM480CNQ8/Gq9X1+wNkQ1Bcw+o
YlW7+06082JePyK9Ag93PYz3Ug+hCy8abiUON+sHMmIl9+0Ad4+Z8aRYKzJ0I51/
ktfH7trdz0+rx1BlVCOjAdf3GMwHWKjCNoqk2GfgKowpxjPCkn/uh0vxBDSvhaxK
b0JcGO3ceRlTvt8AHewjtq7lr8sFBQ9XXiLJpo+6BmVy2ENVCNYHPjNHUa0OlyTk
z/tXb6Qo1Xq2wZtdrQfDHTTxkM7M+hcJp9y7tgXFEWzBW6iA4uv8L97c0ZBgAsLM
bmvFqlDqOUNK4mGlvcpPI68w0NqJgTal9tq/kWiDQV+bTX48C/Z1iUPq2yxmu0j8
a7MbvgNEcCZvpwt1OYz7e1s1DI7iblHqW391huYpCgPJwwdjbb8EGRoBA74gSJev
3pGexknUQSDK0t6f+eEuVQNgh8yS2MgT5ARUMSkGyESPdmTRjzUu8rhD37U+osaV
e9aWWYrfDXNQhfrLeM6hXXrKEQtkTe71+OQGv7gIEJrnEk1JugX2VZsL+yyVq7XN
QiCYHvGenoMo84B01gFzV1fxEfyXbw9JlL/nWBS90t30xklSS3Jipucd/c4+lp2a
Mj7D2kJaCuo8qKVBdDKQFWnjtuq6iUPdRGy2qqHGlTWnKda+/eEWLQK9wPn+RFRR
mfozk80+fWIc8biLjcw0QMiNAMSgraV08GQE7AdtvDpwEdALpm9OfrfoyVhz2kKN
ujd86JWeN+Zcdv8QfQvdD3dpZdYN9bub061f6aUkxR/MJFDc6W+BvAobucr0uguq
U0Cc2G+521Nd/VOWSZLYvRIEpCPV9LjvqB6Xt7EAZkT4S3tE6+uzkeQcZZXASqFB
A4v+1b6/DeQNABI6utSiSU+7Fv26Kw5tOXlM4kQwdNBROJLmA49g1w1geGrKx8k+
HVt5hhuHkOKtgAjKCtp68v9BF+gcocthC1/CrI5W+AdpPecqsgDD78AYoice2PV2
EenLZp/CPR7NFzLFrhD6Pio5eJZ7KLOkS0daPPz3F/h3yZ43boKuBbZZm6IpSEux
BWZCCoLDCNe131ql8sohuyUd1c04yEH+j5lAHQLB18Qo/kkPaNdDnZ+ZuhjPn0z+
XTlPQN8hDBM/al6oe0ulsLkp7aOfD+5NVtEfFoU9bL4UgO1KtdSAhsMYus8eMgm9
D08LNCcyDIU1261WCwx9d3n2pSkujJikdlaIK/MNZPjPDYJp0EfCFH7NQ5Hkayrv
b7PiCpdBQR4NJQJQcGxh+qyIv+FddUG6nHEm3xugu/SE+QHhCPq7gAiAnx2yKDl3
oID12ar7TTvQ0g6sOlDYKyQDBYRRdmw5v8cQMUxDXPk8E+2McV5ILxz5jQ874TYD
tsZ/yyGPPdvK83GR+w6FSuGpHxTzKIeoXhDK6d4Xk+CdpsvJtwtXzcaLwGV3sagj
fZyaJFkqI7N7kjc6VcptQoQ2jrubp4V4kzq2vvP6dxZ3Usw8RObVBn2WiyrJSG32
VcfXP+0fW0oew7Nla1XbOuRZNxeXxcdQIaXJeyl+oqUKPQZOn+j7b6sq2G0sDLbP
jmlfGHzh6LJ3Bt2K3kmeCz9MbsHEKacArnKjoDbYEPNz/zstL0fuCAvyNuQHqknv
FjUXT2/LWAoftjAtVp4JpVzy+AlDHyU8ljg0BGDpfZzrs14aNMAYHZZp9Ra7uVQ6
4Q06fk4Xtmd+Lgv9G7cs3eDUAhmRV7xkWDPrCP4/mW8259eTf8FaLtci1AMaJiEm
+M/DRK5HpGbQ34tbiRUgbPwbwjhK4b/8rDSPsm1KX57msCuXlc7DmrfywsNRDI0X
tQ0HtFFRSh0jkz+PrUzxVgk/EHWlCvzVtuE2HfjHYY4OCvXBriMuIimhFf5RIQeN
RdqrYX9PvNL9mxmMwIii1Yi/EsutVWzH82kzU1uI5qP+8adJYJU/Z5QHCNsQoG5+
XVSgnCdH3WXJgRXFL7Yl1l4ZjSoGLDufC2hT1NZ9U3gFzg4SxhGgeG1GkwxL+pmm
fkuRbtnQn/XXwtsPM+GAlKQ4g/nATWlnM7q5GK8tm3Ywl6lck79+QFyoWXpoJdWf
+rcJTr72IahasAP8xUAvw/4GNCh5whAasmcZN4Fc8t24Pg3hENqFG552INTtqy9Y
ee7Wz2FCAfYi4b0vHXwBg76k/QbW2RVTqtE/pkC+DkmjW9vus5iuPA5xR6cig6Ow
M/nTLDrbqEa0Le7yuom7sJ6N5MZwgtjd7Yb+l9HkA0MGku6wPftx9M5AjXL1XY2T
a/t0xg9ZdLxAW2zOdPX/sKZXhucw8QziMZ95MlBhrH+nCdqeavP6/qeTISpSmFcl
NjVERwoC5epcOrOzzQbdZPsdlxod/lYGxZLtPVqAYLZfpZCbaHj82RX/xz5Pwqjc
tzTZC3Fs9nEB+D5SdFYJFcxmq39gxeD/6msUVOZz9d/IE/tyFgjiX93matFhgSS7
gqYK129SzZLENNdxkTz+0lM9BO9KrXiwhMjeOBSbRDeIQLo6rTDny9peUxGtL36N
yFCqByqb7+1YxczFvC8ljs8pW+EGkYkG6M523yl01wb111tubR0op8abV59taav5
zWjloAv0w3oHYzsCwhUMJLUH0guRw9VD+dS5PNbjZmMjPx8yTNQ1KEGH0IYonti/
NTDYv6yJH1nyhDh/1Wah2QEnHqUc7WF+OLlpsL3RULVUaijHXqifK8EOzVuAIjU4
10XfiVgZgfRPAc8MIB7UYiVXCAbYJiGEZd6y41vrJZVvcLmDktjhTBrC/yShygsb
tqoDLutYZOvbzxFH4gzzLUKk3YmVuQHWXgfNpxmQlJ1TRnR6vF7Zw5E4N4bYkMIH
I1Z79wUo5pDewKCL+AYJ1/WJr2XA+1z4/7tvV+P6aL+YyaJ98PptuKuLI2wZq+V6
kZ+WpJnEsPLJkmaLXGl1jkObRQFpQT7CiqPWeQU8I38oe1kytPZUHSFp760K4cYK
66O0nL4viWd3s4NHR9t2Pzc3l6WfP/h/L95FcoNIzC30WV3rTVwUrDb1KM73p8cm
VG8/uGlgXSpJATiiLI4B8rDmhSSXjq7wIh/j4oN+y3Wl0l4voQJagzcsmcx29TUd
yhDP8V5zo27MTrie4z6pNPOjZ01oDRvuiHSMkXDVzUUDL2wA+errQzdmWEeLwLT2
VQ3LOS0UMffSOWvwgfix5LrWenavFREmW/hfUW+MEyZ2mAcyoR3MvS2nfM+hGr+n
A2DPakf6vLN8+/STkLWfQfibrQuUJdphjUx48d6odyEhwGI8yo3PNDrMnYloyaUB
AYkD6eT3m1JBXX15qcHFN4zs3I+LyxH1V01qV1LOzjCtXI0WpzYAWUqJa54gvG3H
m8cQr1BUXBW13RYGYiMGKDp3O9xIqIFuKvnCgaRIlCzlHQnrNGbCNlMnAppFkiQW
E3DFLhHXxb5y0T0A41z1mRv1Zwd95lu3UmHKp86zqC0+B4NJ2ejd/UlXWPjcctx7
JTuqSnuzroOIjqpjqxzklO78arlViKKULx8v/rVzz+uFDwYDCKSQS/cyYw0HNwSZ
8tl9HqBA4rBhYhGM+qoiqYzUl+0kCbBHqN/7k/pVVIU7NeluldasoWhnn2tKYVHK
7upJxCeJi9JBnNgWlsEdhuhL7ZDtkOSzRpf6n/rHDSeOLF0bucUzOHQZbBFan9J5
pdzDxkICRXf9VACgFT81wRQ1EBJVXG/5wlwCshZKaMO0qsdd+/Xtxj+saKgb6hvL
B2UjerKuzZ3Bx7sXcXonLdnSnEvEeTJBq4hdvw++ace1zGTzesuW27Rj+yvgrbnv
qznIbtnyCAEtvvg+c9mzB5vVkd+ZUatOAD61QCg02xTagdP7w3N2aAVWYqg77I1V
6ods/QBU5u9M+FiCnqZHVcmGwdfhGrgYdFNeObcGb7GQb9UHV/V8a8rTmtyZ9Fe7
eoYNtKL8YyZnk2KJ7BczduaKt0kfdnfSa+iT9OrN285Eg+5oEmqkZ6bje2CmexMi
1Xn9PxodjK3scQ1guiWuyrDi4CQq5bpPR6VlKjEkJ1lL4EdhlMVLjVOyiGKEpHTg
b6Ulw01d1HHyX3VCT69JjuGryiH+/E5gxO/NpxMwDNtLGibjplXbB5kjnBwUDRtk
qvoMqDWBK/fFax8swDz5k4eLQ3GYlqDrly+mweR9W7HylCyrpjE3FwvoP9gOtfoQ
/3z8vyRHW04IozFNse2HC8FdD1U7wmbdkFKRpi71EAfyDxGYjr+9C5K8PbPxFmf4
g3STGkNxa0gqgO3S91LvPFobAj+4cGsdt57YClL53N3H4XTosX2/ussWRc5+Ij7X
QBmfCFj7afkjf28+IU7Dm01XLEEa/0nY7/L+UjliVHhxv8aSrNfwpFiTsC5CwynL
DIyviwv7XOgjfxYrg5cfpUE9y2glv7dkAlxdhu00NIRNgnze0xshCEP6OevT4Fh1
DrvayoIEwCFLi6gSvB0RmYfCmE7rDYTAlBU8hJqBo1EJ5ODeW1/MG9KlBPiE0Sa5
tVGFzhb/ZzHchRnq19frhdZ/u0knKo49TvBMG12l+t8CTnUVdbhHLmzR/I5qQOAU
iUCzQ5R3zQ/VRUAmxVq2hsKlNhj905c2TK9qQdNMAadtsGnoqWxb99mf5XQrJqrI
P0J+NsiL284VnF8DW2d/lmMHnJkumBZWshHQ9g0zsYjIB0XzjqGok+xrdojfh8TY
DfXr80xJ+Bbnkp4mejdsv+dHuBrhxGT5+/0Qt8DhAmlkIrHXNlMImBXrqzp/JrvR
Zmn9tKKSfQZu53rPPnNiwooHr25jwGmhHK94fQ72MbSn1RnWb+QzYBVzOuXOm3mU
5gYP4Pv/AkFSUnDCmAQ6cUIUG5qXa/0eNVgeo9pjeSVMDwb1UbewEGRaEXkOuNSy
3fwNG0+y4AOQOUCzpWS4fh8k/MLUzkMOxrLq2wIZnGHgXWX1Z88bW+xKzkDcD5MK
xzLoguDsKz6rLzeinXPePxznDmaLniVKuCsjguwpqwAQ4eQH8LkV9Kw+RVKdBxNL
clZq0l8LRqjrn+zG+1SQ3o/jIp2OC+E7gVOx4tsB0Z5aBRDhP6t9/YKGfkrIGk10
OlqJIbmpPBHvrUfCsG0loiNSxbb4DFmi+mYmERcymUmVa14kyqVLPPSQs8Re4F7q
ah6ZLpakN5jpBToDQ5ptXVJS6YaU9aEg5hhjiRCR1yLnGtBEb84XP9nXp6KJrDdl
tgsas1E9H4huhJlrr8oc9ToqmdTTD4qxlAOzS2av+PlmJVLallKrIOYT2b4k8e8f
Lxr4IvYIlN0nVLfq+DlSFMdKpcsM/QPbC3b82YhRDlTiO74j3NIbGk5P2w0Dq7Co
M4U+1qY6oM54/42HND/KLF/4UaUZnxzQ88GhY98Qf0DK9RGx/dEyLevnlxNa0bFH
Gjvo8vHa9lg5DR94rTojYiJcHnx+zzzUC4/Y6Mt5bU7yhOYDpxbg4guOESzgyodw
rNaUPbpGLFXqAdvpxPT3BmPbATM5WJ4Z6+viKqFPmdEjsKyhpQ9iybexBUvMbn6y
/I/0pQj6En0fBuAv/zJj57/6qqwBkw5m+q5Yb1taWUoJDcRB37gO9kg44Vj1/6Ca
1QWl/opkAtwTJUjCMpPz2aa1z0i1PJPYEVi2sFCXKIFva4Df3DjF6nvcR1i2+w6J
X/mpFXtRl+7oJTzGSoX7UkvyEf+natEJW8h1lcrf1zFphEo6EYPJiWihmOqr38eO
rbGHWkdijqF+hFk0Qq2/8nR7tNwk8bjp0PkICkhh+b6gI9YYGkxv0DfoFTyJClhJ
WcBc/A5eAA1fMxhMSJzOWWQKGda6wwgwl9TiEzJVgCwq6BCcVkLXW7Ywpd8kCbWm
TxU0b5pqmcB7XLTk1c2MKpBE2XMkBO6YjsRx1njKKvGbNRtBtjKGLKJI4TrQ5z02
hGTuRvA3egK9OUplVYhNLCUI/j1q9wtGK3rfQFvRDZsNPjq0a4QMpqV1SGZEapTJ
b3SiNjQg10v33aNt6bG+iLZQcdE0kluWZNqQ90irutFuHViWiWQmw6xhBC0yTmCZ
fvzuePM/VgMcMRhEzHHoZDD4rUfXVv8pF7y2DwQ5c8GMe3YJZni/6wNjb/J63Jaf
0nV9SO9wqAKMNBtu1gvJCBDQy7sMkCLJZ0BCABS9bkp/T67o32gu71jxWNa2Oq9f
QBLKSfH2d5Zfbesz1t/3APXKwhHGwZfFHzQXciXuEAzm4N/A6fJ212UUt0/Ydoqt
/MbPFAg9x5BpUQKiLbJwkCGmCpoXlauG/zp9H/rnSWmDYH7yTBOZQY8IC3AB1xCD
9cEdy1w6NiYK20krbXa6cuJEJmdDU2qYaeixEKQgFpUN6ET1hBEmseB5AucJ7fcw
Er48PBTI1MEUaDfsiazfZDTwgmlaCktUcJzTflWCnA19uK05erhO3xtS7LQdYzk4
kr8PFSVhnNmHaVp4hCiznWXzd8ZO2SrOSV91qVOFsSX/RQPgL8bJsTdUC0AIDvmH
tjEgpfVkU8vf/9+71FQPIHaiQS7aIKY8QE6xrL/GPKIXbpOHaCGOccqqE19rQTSy
e3biNG0vZxMBHuKjk/+0WEBKcBYMkXs+fRS3z1a3yNuQ+UUrcpW0wGCI0n2keL/B
QGVt0Nqb4Jyzu2XVJ3CDNusWwNffF3z/pRf28Xlbm0endXG7kSJ/alPigDMbxlkt
bZSpPZQnf17eBZ7UENNCbps/EZU7FPE11ZnfraP9rWUFB+VJvzHTA+ZSAIbNAlEG
1EomdwKRdOx7Y0LDJYmaNocu152c2gTni1zKGj13kicNA59Vn4oKRWrD+C3WWDLh
ugiE67g3hzdscb1hzPLYRuy3+OPn08PGoLOyJpa0qrwx1wz5dbCkJf7SEIw2wBZN
KqramW5wng22eahXOAsat1dmNpx9rJd9llcD1OWixxcI7V6U/js+dnaKH8cVfoLH
dsUil7kd/i1aB6ujesHVmtP9Kp5aY5BmacjYCcp9ODuLoHVqVNZbio5eR5QBwa4F
JWTP0RuKxzq0Pvvmko7WR4YrtsgIJm8M6/XWXqaLcjB57K3iMaBVL0olUq7UwSBL
uxH/ej1A+IDwp3i9o5kZzvTw4C/ywfA1nebnySruxzMyz570jpEk/zr2JM07P+JY
XDDXVRKng6Vv8aK1RgPxhiDJFikRlIG9cpY/iCFgtw12RuTuyzYDJ9THOIM37kSG
BTTi47m9v7JPeWyLwEr74JXE0Pgz53LBH8nRRglRQMpzw7FnMjz4kRwfDX5BodlP
X6BbAjK6LtJfYqkXRgIxy07ACH3FyVS9OKC5U22Cw+cKQcQk6tgxQuli+mQ47jVu
tmb8qAQtPqv5SwSPtAvrDMPH2zI3UB0jcDur9Fh6ws+MDgBwLHE7Py8NYV2CRPEX
AHJXI/d+iIkHxIXV7+Eo2sc/m0lmsqIOP+HUgAdLc4BIrJTJIl6vhVm6cjc4gt4h
zLPTEMusu31/6LgnHw0AvsMY0dsu55JZLiM0WonbWKib85xDIgepah/C55HfG4jQ
Sw/MLUrdZoVQsWaHg8hhhtcN/lj5ObdpapdHkJU8/JD+Kyf2xdxt8pLU1sUDukP0
iXjwhvELoox9ZGnPr86vDm8LbomFW/K5wt4PCTziKXTzSGi78orHNZqwS/HI9tQ3
ym/4Fgg0lCR4dc2Uuz9Sm+4xA3HDd/k0l1Vj2S+/5nuUP7nyybsXv774I6Z8PRWN
nk4VJ1nycw+w0YRxGFHZ0grCCSVZU4CePl8FvZEXqbcXyKv86TzJgpEiksmB31O3
K9TU07ra7cI+OW8oOFbbnMg3UhdMXCWFFnv/W9Ku2s3MyE3HAug45hQ4WtwmCndK
QZ8SnDcVmcsHa7eIp9Rz0GMBa+fuZP9BsLqvecCLxVPxIU/S2xNur62zAaeEgp6B
cz8dV7G9C78sQZzKCOMPvM31Tp5pllgdKqWmnhwWQk2HkBbGXP5lUx4PtXbyAiI9
yz4zYlcP3pet/5lePnbX1YHtRlykENFb8pa8vHRmAHlmWkrC+oZgldLQJimK+/mW
Zmb8xsW2SJrwZ9Bilo5EymOOaFxKS62q2LKFVMzAn6W7FKkvpqfF+KmlGOR2MgJj
4Hiy6GAzfrdIw/M45vY3DU+vP5uALK9aSWV7cbykcJMwFmqanIzR5Q/8JFsePfmk
FSrAZB0sGtyxP3TfWocvh+BGVSD6cO/qLsJvCxOLZsjjYWHYi+xVADcAcgTiK+fd
Wa868TqW8W+aWeNMegQ9IXwC3SBu+SoKuuHsdxpBtfXZ12u+yDimyaVm13xFyxXr
c3TE4UZngiEEUe1Z8GDceSUL11hNiwBKsjp5mZdB3bHHHaKywVB4Rau340RuC+sF
ph2fovzJZpDdv2CBHSPrtGAHL7ZGLTKBhDeyL1lGLjjmy9L3D7YRFPDFfErS0Yo9
At55cIfU06DbxiUAsks4aUv0qbk0MhrvTyqa2jUqXUnWQyQxh+ozUAHbXJnhuaob
flMs9DvsCAlbgUwRw1c9vip6CkpwRAZTD2mY1juZtJEwtqdJP470o2Si6Q1Zfyye
bqtC6Dhnv2HuKeCCHiHBeNXuO06351lMmKOKUA4jD5TXHsxeH/ucBIWBH3qhcbWx
/+KghlpaeeLvvLPBolnTPQCrbBwRHVRSMkoFhbMv4Umxtu1Ll6POA4L6TlC+tVUM
yxIFz4e2sHMnNwkGfKL3EAXJ2PI9a7DR9aiFu/abpcsd58r4+8lpNRnOsZp/CRa2
2AfHOTEJ8uWlFXZ11WK2aOrUzAk+4MbP4/mVyUvRif0DltFachv4pn34jYw/XRxM
yuD9LUY55oQ2B8RCrmD5iflP9OhpckiPY2raQRcoOPbi4B6fN7rLyL9toYj5vJlZ
Pqe4cUCOiIGL1VZ3rPoLnDGvQ8IcE25CUWDI74hzV4nP7rCr46iS7lzeLxpIhrzm
StsFJVG/j6MR5/57beUWeF1rL1etL0m9wsFHua5OYw/2P9vchDjrtlwBrAt8iQm3
nO5RmEiCI6zgida8h3XjQi8gj3d7uICDuYf6sHi8aHC2+rsAmINY+0E07XZO3zeL
9K25bXm1a7gg+rmRW3X9nkbAA93zf70mfevzREa+akLJSYXsbYwmRPfXfoXCsBzO
Q8ZazW4qMDvM8O6t0Uyy5MjnCuEUqNL6Qk/6scbCJopm4zGxf6WdPVGoC9URSYvP
qlQ8uFi9fmyXv5HQbBrxtWnIICQtdY79JPNkU8N47H+lDkoUUDGEWu18wjXeW4cs
+b06NuoVzPLIi0q7WyKS9YdxUAc6rHXOtO0Lc44dbiTPuzioe74AaClu4HJ/gk9A
xr5JjYuQTtTDLqCVjWVv9QiOg0XlKcTYh0V+A8yah9TM7W/55p0tqiOF2YsFM7hv
4lRDwKohyDRQW5AzckFPAOxLdOol1usYJkYX8MU81z7xYdKQHKpZBUek7RI2RpGq
675fvvu9l9CLA+acALhsrA/uPH/fuxPjVX62ErNdogjudM6GkA8O4Nn0Y/6hyz64
yCO6QYz5dhbiZJK9YeB4h2LLpHHuLzR+/Yr4Fm38uNFMYktVXP+KOdMorLL5Fnik
nsFMN8wpX69f6Z36h3mEBRotU+4hbn6VnpI1/ewxUKWcKqrpkt2YdvVxmCvmTQd6
GGZMDvZcC1cXxAyRMFWKnUh6cK2BZkt/4UVz8Yjg2o0Aaj5wuEnwc5zvwDlr2t6n
Hdsjvndvwf1EQmEd33y8VhwxIEFanoesuj1aAwpW+oBudnFThEejdyCujwEu1kx0
lrywgRjzKeTLy2RcgQnJeO8riPMYTFkl/Sd0UeZEWnmfnUnyeVdr9Fhvq6YlslxT
fGN2Me1YlHn/r4/1kSapBKL0x266jUb3AOMv1AbPgzcsRXqPMct8lv5nzYl1w09X
Z9QRMbBO7NntUD6aM0dFDd8SYuvTTnmQHmic4lIf//HBuGV2e08Q6UtUtOLK1XhM
d2Jjyhtu2ilXQnUUakKkNalJrymS8h4+y4RNMs0N93FfHjda3XjKsyeu8jWpDGk3
Fl8gb32UCcSsNOpzexBDS2BDTrauTWpxp1hSk0GR4xiITSwP+Lc6FOH/bwj8a9Ej
f5JxIFpAC1ISqmFrn0ZiHDfcFGy5eLr/+6y6mYC6cVM+Ui1Y191TnYUz/qx7lRgZ
ojVlIIDYXVmvzYrtBC2MABBoUiYgNQmwYVRCn0hLcn7iiek7XCYOAc4nqE+zDdB6
3EqozAsneD4CL0V6sVjNCNUhbvv1upsqixcs6B3Hpg3H5ENPIaTIB5d0qnEa2HCp
rk6TpBoWobYsFOLOeENBU5L/K4sjbPQcwAU87D6bF4Q/xUq6CbW6geLZcdn+ulTE
9c958xjeZtC2LcAEyFpHHojpJe8N9OsXyj+n5CXmpOYQlUuYNosAxizmi1ScxVYz
GABZzPpMykUpG6YDydDXRo9Ra1vtiuusAU5kbIfXSxI6Hx9SXyEVXOb60NEJqv4a
aOY+wHm9l78roF5WtUU2qeqA9VQ7CzYcoYeuN11VqVILDNCpLEJX1uPEKi1iOFSU
TCPh/emu+snkp8MBEx+0X9UcY8RYjcu9fuICrOPZFdvSrge/M3tnJR9pkHoCCj4e
F/bsdJerEunyjT8fO6BtDU/yqXOr2aTxs1E0AHSTd0gcLzfrPcUkYSXC84cZ+F4a
3XavZIBkqNl39UTqrJO2tCOVjMrYoUm8yU56MLe1I3p0r/stMy67zBT40hp+5vNR
Rvabg/Y95O1Twm9vjTmbHgIeAKjfzOwYswk4oKUKXOeEwID2NU/wvYXJSkg2P7Fe
HbfbISSHMYGVXpP0uuvBmyBX/KGAqo4QqAIoBBYVKSfZVcMYyjAksPccruI+kHYD
1IV12mqdQKlDSMjLcwY/wwCEJfgR8HdsbOrVHp//VcQqjWsItkjpE4TofojDydhG
1d2yAdv5LRzBFjvhUl2I5FZYh7n4sBxRMdbVOcOdTGRG+KDr6pItjteDQyddXey5
qStOYppQjlNf543/Nqbk1XcrL9KJTdp/FQ3ql++0vyoZOamssjjBauD+1cWlN578
/dW9ToGb5W6muyeFYzgELNSNbkyWPMehlFGOCRFHPrmvlx2eYqNSk6silo90mvYF
1f6lcCk5c9pmvRx92TRTMM6Y7NUNGtkZGCkk/ES1pGiy72m7s7KKGRJKzIsCDPM2
pg4c804s/nm7XEcASUn7/aEkfq3XoahoZ7+7LA893V847Ps3GmtP7AbUNQd/CStQ
r6FZyMEjV1M05+Hrt5u6rPAq4XPuO5AaN1KMcObJPfMh/24Ncw/0mj3PuGEj0YBd
6X2LcqpCfVWNb3dU7qOp7gSIM3sQIaO9KXYx4yEgbY5WH7y9ALX39ciViptiBqPL
OJ1TqMrvmw+XuxDJTNankVTmdAWWIZyVSt0MD7Pr1u9fewVMWKPHvIpSnv4IA/Xp
8otVJc/kg/4xdpj3M0E0ls2v0YsDDtIa1wX6jPvsCKXV8maNXEUSgDw9fCRC7YEz
Rb03nOD/jQElmHnihKLNd1QHHbgBq0FsHGvIK2NM4BdV6xnUk2Q2jH66iq9zEGzb
hGXB6YEniXeXTgBkrobuL0lVrxvJE/qNAWGfbUGai9XlB4C8KKONr46bgiyw9ukJ
v4bga08Sq9pcmQRY4LyTxDWF0UnlEShwql6sI2jXAgVdQDwN1UlTSkemgBqYB5AA
B3rdi/t/vgXWXmk7Zc3W9I6oSWQFeoJPLvoleszwm6hDc/uhYWYkE3DwKmOqM0z0
O/K+Ku+kF9phfpmYfntN+wP9ysVMvfNdn/kUXhRHvJ8Goq22UmosCBgMgxc2jsOM
egzc/ePMNQyJwMzaBy+6d7SOP+d0x9cfjk2oI5BavXzdSEGnRBGmT8jbA/H4TGon
oH+TZWFPDjMrsUdHVdkxG/8Cf7X4XEPMusMzu/lih/YFUUhLCuGDzJCCvpoyJ7gd
libBtREbk12tSw3ZAInAHTkByJ4daAbid0FB2NAa47LF1oirM2ZMk+satjgXwlFf
nlY/sVPDpPGVsyB6b3NvWvY8yL+IqDUWT1CMgAd7z1kuKzYDkl8isoaqS2pJMABD
562cVjLkqHmIY6YqMxHIXV/S4HIUbgUK0rIZlmRvs0Ke7GM7A/Qygp3HNC7/kRqc
kjkB8WBoHsATG3JwcC9W92ybHHBrFOgLXAZloLJ/v27pui9Wxib19rp4qyxw4Qss
NxUywn7ALNS5LpU68AqcXN1ge0rM4Tt0E+9b20UOaAiKuY1JZcih58EZn7yxhrLg
5wUAzTnD4u0GIHvHIfBpgZne6dfP8Tg1rHZmJNDLYKoTjfj+5jcPpZykN/ESFysT
ldy2WEtjJ8UjM5PxWbHTBlM56TrHtNIAd/lQKUbBlWVyJMjrME6L6TZ0jRJLY6XI
Au97EeaZV9IohlgZ6t3t7JO04dJdQgbcqPOlL/d8lOQKDpsmgwdOyD+jJipPM5v3
DK+Z1UuR0Dt0rdHx8jgFQVULnFGbiMyymSiHq0WBD1HzNr/441/nE3ZurRM8ZdF7
bdzQ6icy7meX66D7z+rLuTlIvtnl9S09MuhaKdYxWtK2CaUrMr4K98brTo236PO6
GiFPJTvXhNMby8F4TzZX/KdoF3lBrb4/DVx6PFTemZUATUgrXduWWrjy1p4WIdcS
gpdoAbDQkFILfrvvJNG9nwD366MIDOtsNugU/P11P1id/eAGcAci6/uLhIdbRxaf
jdmldBVizmu7lANyefJyOZh7hdwPInCzCr+eLauFe98bG8fGWy5j4SDjZ8K9Mm+q
ILo+CE7B9RWJ94unDDW2TdnLtVMu1G4xOMMNFXoXH41yTB1oSjFklMt8jVfgHdNT
HH0ofHlNkw0ix3dahBoqlG9LJ+prH+aO7iKaaaDhBFBc8H8UAmSNfj91cm3S7lVs
HQlyO71KE8ipB7rWChydx3yrQi9a9aKoCJZrVl8/A8T0XPejPocvzIX+xN/WNDFM
rt7rt0Bo/bvv+3NmCeb7rFSDlQShARVRofsqtuVyvzKQDSjWKDBG02VDeTG3dDNz
rba8twbq8cWIVDrWPAnLd3BB9FwJmkIFpokoxteXegmR66zNuxCu2NHGZLIvzk3a
LreVag6gccrDF59ToUBOOK+dl8O95fOxxSJ7iwFnz3Py5Il3hQmg+icChCPLNAmx
sOro2HGXM9mGcWnfiw6Rf0iYqCROFiTg9YcoR7BHO3+GnX3Prz8Zk3WQ5pC1mu+I
Lo+hWsMM6a1IfY+ECt+2TDUeweNREY53jTE26XBZ+7m2xWNQlNavuZNyBzZ7uGl3
/yW45coDtfuxfK9Y91/hjBjaHgT7aTBUr5uIPfKRbY2b/mKKkg+bK/Lqnq6osYgZ
bxPxgjihd7O8upw3ncQ3KEQHfNfVBYNnBpOQ+nPEb207yGNiNwZpZyhAMzw/L3Te
6K8R5TF7e1a34CjwjspqrCmFm1VqyJPjBTN5c5D4hwJrUhErRnXA8g952QL5tTzE
KJkbaN4vH6eA0mE9KEjcSzUB46Vr6CQDExkKxMEfGsiOEJSLlISi/OmGlGO2GhJG
jZED+OSJJHgdMpkMvletTgA1fjrMigVnvVZnulO/M2SYDZM6BQ0/1MqhIoUSjiMb
OYI0xs2eU4sfSbAvwuENRdqIMXoNtj4zgsgIf9cbDXdtYmrmXLZDdA02tKmw7GZL
30l56cPyEEM3Tf3dTo5YCIHbwBvfKo0jrDblXDRQFbe6SUSh4WG8vB8u6jGeA1Fa
W0WKooTezDcJ8Zn7m5qxaIYOfvf5E7Hb5/TgsNT3gxWTnX6Yv+qGJhI2ycJlFvFw
3aZL5UZ5O8Ez5wQRm05mdLiuuNGZazJJPvfumRACDujStioc4XBQHkWbyfVm+zAL
BA38vDEZLJgar4bVH/q/T2M/vWu87M+ebeMgT1Ybb1e8dBT9DFbDqC2fAV6tDyhy
JqSQB7xVVTrRqxKBSg4h9MOEVT4+2XDLGeLM7JmDf/E0vj3sGZPFzc1XjBJaue53
uvXpFNRFV86nlWu89BKaIoqKSbceAI6E0ahL7ltraChBf5Cw2oXVAphPX2K/fwi0
I+85PbPcuYK9T+qakCA98zQwQT421tf3/J49CMNJwpcZeYYzVlWC6oS9mvEHJYEo
ysDx9fIH1oPOXVLmCsrC9xkXKY3Er7bzpuIdeHlkJMKLOMp+/hlhEq3hpUpDReR0
8nwpf04dk8iS82Bj5F+s/9WgyVwNXOxbFQ6x6Z0T2DL7izKgzZCngecG2nCSUsQq
sMsJBHm2P53sf6TH5BOIT5cikn/mnTfy8grhFjFzfc8EUKk/bbGohmkBAH6VQZyj
yk4b+FbfUCW7Q1Half+kIEYV4nT4w8XeCd7VAPnXEo7YRbpJZDruz3tnoqmdoz2c
XglCBB7mPBPW3pSBzwLSn9rMiDeqOd5LPmhSHpzrqTdNco731U+jkVPwI9K0dXcD
VCHGGXSJydVggMyJq0xJ57RpXa62I1xyLAfCPjb+/goGGwKT9+/wvierTSgkZ+mr
IIwIFvenRSTScDh31BuAMiNQL9Xgr6EuPHE3+kw1h9PoXK8wUurSW5/XxlUKtghS
l3mKuZsJnHCs3mSTtL4nR1OZIsCeo/mDogg1FRthV/9Gm9n60qN8iBEZMcpR0uqM
kYyzToEkAGf42D3pw7ZqMixwWOl2F611oUrET9hMtygrvSsOxkjvjCNwOKiMQ5Iu
M5Igu+RhwCXZRvn6YlNqv6UzUMdwMEv352EpLq21vSWc1Avg43hz3JTu7dQzyUr5
6JzlDtsTG8HqNusLeO/XB5j5WZH5PZenUWRrgA2GGLf/hzRa8+UOrAFhiVex5K++
YOfnmnVQSrMpsiBYUzn+ZrXs4Ke1RxuKzKM2I9tmDA/RkHS9KL3iapOMRng/ZMBv
ImuIZV+3roWz3ARKr7yd5nO5GnlTzkNkVfR5tUcamCF299f7k8SOuI+2+KdIUW/E
48cYbWvwH190xaLNnX64n1y9puJTRcgzENADl9fx2cpht/ohkfAUBAZNSy98LyRx
Eccd1SIRc8A6Y6cHAVNEqRCOy16TD3F3R9huQZfOpPJzZfBlM92zHHFtv6cyZWW/
+s8TLqf9VALZ+m26xDCZRraBl1h6PIjeSIvIUZyP/Kmlz4IdusUxMs1nXMjJJHsA
WW+7SZ8VFn/bV4agYEhQe7lse4O9DfmqSTlV57/OMe1dwA0m0xSieIIiB6D0kAZq
HXEXoxhne9/QlScVwEWn20ibipjLMstwzUuMXPOXf2qXFZ3BUySTql8XptgIwJo8
ZTVbg4s4m8wldHcTz1WTT8ZWz936+FDLgPIge3hzxTLggEEGksphwQuO5fQqC/9Z
5BZ+Z+3ewt/HBr7yzpF1CVI6fZUDGdpaiOTVByrMrZk7g70mePiKaQQsWgQn5bMj
DuCYPnqFuB/O9wDjlEZdHAqobBUMlpjEiIXfUdcdVJ2FcUjXZO3sAGhoFMoX8If5
pjxkcwQA1tLbZRRZ7i6/Ul8G2jypIu0kihjdArKBXUxzj2fAwSp5wfVY1/jb4EGE
VuiFNXpQ5VOf3bQj9mTfQM1sz2rF0likoCiRH8bgsGx1YrqukzXKqqLW1V2MBlEW
5QHSnXVUGKkCkFvlXMC4jCgTSjsLvBc7LuUMjwBZDpOIHHjza9Vq82w3q4YmItxo
hTAaxTWc0XGZcN7P9VgAH+hSXB5sTzApAKtAJObhCzRRlrZXtai67QWuK+dcig6e
093EY6+dmxkJRcAEKbD5Ragt1A0Alcvw3f3WSGB/xw0OPsEQ4hJyJDZkAOtA0JEG
nJPCTXO92wLEFVruW2IVu8ly+ib/gMHZ43OB2kfkrOOv/dHiy2TUA0iwZqFzpt9k
byhT7m5iRlttu5BnxcG4qBEexkObzKrPEYjSVdV9cbG1m9tSVDivDU/fdySWL5Bt
5IYNkh40ncfWItQO9mGumfZoHa8sKMxuqMIKvrP4XirALexfhjD446V2E5nJ35ph
toPHAPsl9JB/yH+m8som8CBNt8F80On0WR+ptkdppj4d5BiNgXlZ7HGpUo3bOhTx
TmbyrUHZ1QHwvT6xo8RFcWu2N4M+P/RTEOMWsKEDzZfhgqLAf9GKsLxka05trqjX
wQRZHtdBIno7pulElb1My41qVPw8Z0s/0TEshKy8YK8+rvWXjSsH3RaRC0a5F/gC
UHAwBdscVWQm9S9wDiIhi2oOoMG5Otp3EDjm+A5tUtv6ytrB+0eSwcF13nJQs56s
1+tKj7xIe0SBQFyL3wM+6gXN0IkPSd17kUi2l/rCcFm46tJjKbo2vsb+QPGZHxBr
4qcaTLnTZ7aaKQH7bG1iYTDrrFA0RH9ob5fI0Jf35m+PWOtxG2L66GjKFfDhBPRN
OXpOyOmd+UCPBe2kpb0GND8F52MLdZkGuUxgmjyh0r34pChP4O8oTf5GzuBwLxWR
7GgjBz2Ax5t3W73s9evFZPnh1SCJd6z946XDpIPUodQAO2Xyv9LpBIvFaduxiy9q
jeBIIgjR/uMZG1ViCLO9s2Q+r7GyILh13WRcgv1ntFazqLrgEg+8c04Jym+IAQmv
2i3XHKCcveTlCeUbxkvYgELa1+DIw7sPs/e2F08/Yg18O8ixn1WOftzSacKO3LVC
dbqA/CbbhVJqlc2l48a/wSsEaXLk0t+cFS8j4ozO4xp7xDGJdTvv8nPEZ21PuQYK
4hsThOb/Pt4mtd5dpo30lXPSMsfLX8WxGM96tp/6ROVDfkW4aJPnDH11JovrLEsE
gYpLKJaeX54rJN2OeXWByftkHVK8jZx/hskDNeR7TSRxiFwstWm4QYuWyzOyb2hZ
31/92DhQGiQjEiGlQR6a0guHHYftpNYsgbw39vuC+zDjnrRaB+bn7lSvDqgO+VeR
4tBExKSPF3E/6KOS19j0dswjKE+Sa+fnvT8SOUaDFBgi/HKp1hXxDQdUMjGJL63m
hoDxuWZxj4V/pYaBeaMGov1n0vQTQRKmfln2udi0xlrqh1QCBMB/PpVz7mnb2VOr
VVH34ut2AGbw3yrmisUTdCfhnZDvmTwXhffDkCUYzGSDiXXUuBkHvDGvgnm/qpB6
4cfUOlHleBWOm8Dz/+C36IhSYoeEgMZUfuX9l5um02D0OlqItZ9E0Z93KW4OLKjw
l8layNhvoNJyv9/dtf3VUhKOX/32FiqOvz0CRO2WK4YmtgZCjrJWQMO0icmqmc9R
kLwbxlAuJAgye+I6lPRR/RFbdp7elGBz8X69YBGD9chOYCo2jzbu7Ru7/medn2DA
YYJr6NjRT2LXjmGAMG3ZvqSGEp2oTFx60GplImJoIRjWKx3IHkzB+zSnY2S/Uh10
OxGRkeldix88xBC/1vcKU+Wqlb9IuH8hThcnXuNJwYe1fe9Dix72+4P3OsyyzaRS
i7p/F97MNoCsTOqSj8ycZtmW+7FylWcLkVwEAbOToo2R2RQrmoDZxahxOJXIY0zM
QYXENnfHovicqT3SXx1Sl+ZwR3pbEvjMeyw3gmQjtivJMuATcz4ZpiGMZsn1LEDK
Zejpx3EMkinA+PFL4litV7JEt9PDnVio1q7lqLQrqqKf4c3Kp3IEzhWRKkQnkXb0
BalgeY8xTKX8vJjb8dt9saDXXMwkdWviX8fwxVybzSK7GoY+RRlD429zZiEh1BQo
t6dZPR6SoaxM/IXVt3BavMH8ordt1A77SH0PrUNMeFQKsdcOQ3Js2rfO96lOCbPJ
DXYHnIDOwTag771gkxT94JYLpKiSRmnJQJWLaHIogWCUupREsalFr3goMbgg5u4A
1lq40KhQw20L8ZJcEiCFYH/W6/2Rpof3XcVfx2zSPQemMu9DJWeVlN9kD3DuGltk
JyVfnNRNEgSKRnnZXp+bPYWznssa60nntGH6S8wRwykWnnRZRO+q/9r3czKHCdNF
PuHY1JM14yZngNI8WobuLG/YwmiliiK+wlbGi4bt+irv6paCoLHevwkkLvGqELQR
yEIMph3l3Zb5CvRM9rwv9NRrIxcL0EuteFmMzIrCikfCmdHW3jtRavvZoiPpdmEs
QRbO7UwCrA+VWqXctW3lYAhNic4mBgTWKU/AafJHVR6CAIcw2mZ855rPnAi/rRNm
6AVen1Cmue7NuMrFHvFTv9lUKnNo3NluDeE4zj9MYcIcV9MFNuvmYCHrRRmadKX6
CAr8WH+FnrJmMhx7bnQ2NCEkRp9ytos0DcFN5F+bDRx1F4UVYu4MTGbmKJfcmxxC
B2FBpZU6GQrlVMKLBnCU62JlqIDXeUipLEOzydhFlZDDYo3y0iIAlI8RsKHiCVgp
d+guRinakmjBaq2hmErRvHHjO1a3Zq/BKDCd+70r09Kfd3hH6ridSnskkA6Cnh/5
QfOggM0Up5M9xgUSWnyQuHUhOGv74alncSATzmrF9hgM6pqgEdv3DXnQjTxFJ2BQ
XjZ7WlM72HNr3xjEHESpzXRkdYJuTk0V3iofIFPFenxSpWQeFndvTkuWpLhp7GRY
bixJMVT3mLCnR9ZYus7NnXAnNOTN0M7RQhArukYTkzzUoJnwGWW8bMY4jHyTr4LX
ikQqNzuIV5qml0VrDZFBvqJR6rEjuOW9BhKk9el32qqKmoCvDkBAtASKSjR2yJdc
rgyVjzXaCs1XbCezTv3C081ZLkgXZ+0YCvY2lpIXZkHTGVBXzvOXHbBdGnc23d54
jWLm8qIiot8zebq4unuqv42HZb3ZLYbWg02Jpa9ocMywD/ENCsXtiPY4izgOxGIb
AMK8y4aFo+JmyL2oMFwUrE4mVbllx6PGHikGmAaSogod73uPwtaaR8k7zaRGByEv
ty+rOKuIDKZvCLRrIUGDSAJveO1ebkdF3bnzC9igkqBZ33RZfOiBX/fE5aHlPPCk
wAXE9vVJYn/V5AjK0KZ3uyWHAdEqUwhuoHYQqWkyuy+xLNanFCq8JiBHkTTuaehR
xWzfPFD1m8wdtUM4012d24rr0hnOPXZIQNmnz2bpj18FiC/lhiB5oAI+V7JL5h7j
yd1+E0BmWOdlzETb9AFnAn7fmYCPcN8wRNiKWxTCvzw+0+KUQDfDNKtm2yVwGq9W
yWWjjv9v4yJ0hQPoJehCawOvMn/CrJEH6bapausU02Bizj2DltK2JTpuINp8znA2
IB4PDVDpb45IPWIYV1SjNH/C9UNUWfJiKIQgovrQnkpz+HB7T7ey6v3jIz9Q2Wzr
9eDtE+zl7S7P2yW/e9g88ELjCletHbd1DZgEHGSZCeYmP6Oq+RseXUa8Mi0oJJtB
GI27TWhEpe1Qo47j44LMIA6vXLnLs02rJYUZbZFoh0rJvwPj2aMoacW7LBIXNiVV
c5TYkUK+uvD4/CuMv7oHIlIFmJ0ZEPksoPAwDe1oNEpxlikOGJ4erPOsF4tUZghH
5ASt87rQOUYwZSz/WzYyGk077EGQhTPbOkDGteK6s7oqmSi2KZTEnnw2IecE8FzG
Dg+DwhmnodCfrkXURuVnv/KtQlm6XqVOYz1N0ip9YFknIuo60e6DrabaqKhY9bWg
Yf6jlGAMgepifCDxBbHnayOMsWRnQ8Lr5Nrp7y86BTKgVdRMTKt5Lfw2Zsp63SLf
m/TpTevkpehDe5jgVEsQnlWI/+h44EFs+Azp/LSuUwEJ67xK/7TfIfVpgiIByWz3
X2Z//cGoR5MXXEMxwUBmHu9ZYQCCjtgiRv4XPnUEFPp6bmYGPoZo8opMjyMjlR/u
e7GIj+m17WD3b4f69rhtJhxaF2JYeWUtBKq+YaD4vpd7xAxjH4Qzwrfi7R3zlRAc
PIHDHHDuCoByTeoMPG63L9qR1ky2G83l5zPgYUObGEUw0zKWNRc0PEGjw0J+KPqO
BDlkTF+sHVzsdmWj/M7UphRiy5CwnUsZDt4RLsKu1dR27H9IrTEjovd7VUf7AY9M
EIDiutMDoLeVM7FUTV2d+ux6NISN8EyBKX9mXSB4VLRTf5ahq5awPmcXC962aYQY
aFzuwxYhfASdpqpQmmhOX+qxOLSBLrOrWd3S3PjqBu9nnrUsK/okYjx/5Cd0+uh7
1LIDNj4bGgON0siTmc9h1Uqv4PsqXeOSbIka9zTlXMuyQL8gaPVRgzfcPwSGoZVi
tWX/DWV3KbABOy5HLSkjjvWatm0zAzuU1WuGgHm0JaWX7hY7rWhXPgxnLcuGY4o/
cbcNOQyQMh2ZvUh98ae3nXfODzj2/YOkR+kL9b8yfKRJkeZhVL5znV9E6D7EwYhx
K54ErsPqCwqQEI5eZJ9OKMabUxNWZ9elTTkZxJb51t/8EP/MqE0b71y+UpseFl6u
+8RY3Po98hUoHHWfVfZZ3pELt76h6WqqUSlHyX/Sh9ruk6I+D7j1l2Pfi6fex5JI
yA+lhtk5Fe83JUe7RocJcXRvE8KPhFdQSSyJiqsVqHwVpn/4GwJvyRHxXQx7fKbk
QxL/ziI7l4KxXuIdiEFDarYiFhAdyvL5Z7ICbmU7lkwVJRwA1rwqbMquh1bxQTLR
NXg4iUjJYrI2XhSLeJDAtlKF+jj0aTX5KJVuFiPmgYQhL6/Mzqt/dOxX3wK0U8Oa
axe0F0Ni/HfvmlnWiesTtAZrX9ZJHPF8ijq94ygEr35LQ8/cs2/IfK8W6ZnPJccR
A7XIDBKEa23ukYQoWWC9nJKUbvbcJ4+YFkA6F+AmQLf7z997uBgxQIU+XKQehO7h
8wd3oxu8HAT/RFPgaWxa3x5MQMTDUo6vqC/eUm0hoyvhtCEaabX5/hLsb1u6Qx89
fm+Nc8i+Kn/Hyzw1fAbDYRrv9bVTWhtCGcOaCMNSxjsV2/UhYIgPZV+oitmGrZXv
4/Tj8mdGuavVw9Y06m0+G1iApI2NZX+VsAqm2zf82FYCNaOvyNUcR+JtM1WF0fWr
KxXArPAWeWCpww02jD7JOLtZryKxQgJ6qfKCqXgABFJujDazpizBnRjODoNnqCMx
XeTDOIN1g45yJnRHRu3Fxiuv/XfVsB37F1Cfm9oZk4Pq7Cfs/yBPkzYGFVgXk2Aw
IWqKQXPtsmiQxOH8ZK7Cuvw0V3gkKFcEf2ymhJUPFl4Lv2YQ/MoPNw04vfclXAuE
eBgnjVx/XqcR7N6IRIPeLTeCv6EGGtthJN4Owugg1pGAqU2BXPfIFmkz4mwhcilI
6MYhrCKw/LBJfaXxCbfIST9LBbbmLho5aBsGyoPt2GCDigAOP+cfhMlk6CpMUSvD
zvP1xRjM8R5Svq0lPEnP32wbxQXXa8OjSKYb24cpKkazYnrZ6l55df+AJN3M9zk2
sEMyDPO+1Gs3JGvqpiDYuuvf1pG9uF4cuM4Ty7Hg4/iDRaUPR5hyc8o9dCNwwy3E
8tyt/kbTC3wb9lo+3GZINFHHtHtRqNsz+J7JP8PnKN+5//u1lW6iqRYlNcV6LQ+v
TZznZYJJJzLq2YbDE3aK6wtOXEkPJbxecqZBH3xPEF7MHp9VIEQeUp7ukKkvrwAn
JvQ3nXldlUN3KtgLGk++hHIfAh2q81/smUUyfkVE1nQNkoft5ZhZKiyOt+YGyRBP
OsTscA0Q6ILwOxM8aShK7NJAlrqw6sqTCzMr3NspvmGSaasvIfcMo4A5Xdxy6BSo
szSdXhU97Lg3DR3ck6QbRigjcDkyZJqSa4/KEd+M80i4aRjYrtAU7Zp5cz16MPV7
FmJWSclB0aDFES7kS64gblxQq9oT7vKeNDlumivvwqmgc0va73ZfewBk6tPO5fmt
wX7TpXULMHCt6nKfB8bkw59UtT8ec2JrhwN8NmjgxEhhwCT7/uazDShVFrUvax1z
K77ui4DSFv3AHYeOIasCFFjJmc40gK9obYmwEuu1SH7ENm1pEIw6uvYmlVIDAQsS
6ihpiC4Suqhb1tNIdhwsndjOu4wM2jZuIPHr4Xh9S/ge7dyrojsDJwFST1joKaMB
xs06P4DE4VMwmYhooAnc2sJr9AHvL5aTGaI9Jwk0UVmIJuQzwyF5O+HE0yFu71s4
qrsKakCv4bbAyJ8u8Lyoof/kAjpVqomDTLnt7f8Ffr7D1zep1LMxgGtUaGWo1K+i
TzS0NorL2n3ipn4GM+xMnksgQ/gQQok4Da5B5RUdOPQyCWQcK2Oxh3z2OAbiHUce
Mv/QbfvcCk5DJEOLW8+NC7KDlGV6NRMAImMgwqr6FfHUaxRJ4bvlxhTfb5bY59Fv
DUD9X9cS76yet636zOv8yYiRGaCWB8eBzYy02QYnTrgcsfm1mJbJHlUTv69lBBZY
LfHRw8gQLsMv0SlcDQeObf6focZas8AP2h0BArQoy95TP9FjynaGaxwEbu814ouK
7SGXJaoi3sZHLLuVjNF+wwl2gwP15JP8mI2YnmSB2g23nX+ye5vFuEUUQd29UXRR
0wgpLSB6Kw+lu8EeiDbrljB5/ZOQwHplySwDoBjZFS16Sg/RIJHFAQX/44OmQNuR
iB04gg7y9Fqr8eoUofX/P02yen6fmyzEFkr4t1UYmo/SkIjPGlK7r95XvCQIqmtB
ljTYPSdNp1BNqIiD9Q+1j51/8/bZqpBKlX3yUfkhj9jLP/BtT0anCb288c9OWdyt
JOn1fjXji5xiqM2L6NjRUnk39IS8pC1d+iMRp+Q+dadDNZpxAMYQ0/5kqV6ksKfD
ebe4EPSrZ7IrR0BSmFuGAcBSgbFAmLsGO/u4QBoTHlgZ/+2irni+NmAOd66AnMN7
4g3Nlp8s7z+eO5UxLZr1dKakzj2fPPzWP/m0VnZAjE3DJJdQXiK5XwOVskGIxFWy
MTHRTE0pYiCwpuL4jONGV1c5RqVpsc48QZLddnj1jap6N9Pg5ePLudmf2idNIAkD
8jTpTWhnvILNrNAFUA1U8X2Q4uu0BxsrH2LQaJsciFaE5afMR86KBMYCnuCKIbZM
q/IdETMeNhyuBzzuSTlMGxxt6bN/eHlYQpafA+wDyq4XyW/3AXTgO3WszDD8hOxE
og74YIcTUVcmMsEPM3tr2+CICWxdDrhwzwxygBFFKEOoSEL6ObkXY1TvlkzetZv1
mCAsEqETI6zwCGbEvIkVyuvH7YIxgLZLOhmrJovh7bjHy8i9y0U3pEAf7LS78idg
g9IY4LuU6+Vgr1S4PIc2cmBRiv95GZ8sXmZhRY/o4SNORcwtGU3wpHOP55I1Mbnb
GPt3GvDq9N7KPcBNSuH2/y0aEV1HuzxguaDOedonCVK6idqqNcs1b8uncngnmxQO
VVFf0Ft1GoanKI1iTl+pEdyX9AVAms77vf70JgO8MXDLlKsUVPLHy4AEv3brqyJG
HgDX2tMd3E/VXyWlXeDq7/QrHuaCOYNYqS8Iab/KqKmWsChgNiq52ZqlHq+OJO/5
bv57I4dDPhgkThEvP0Q1UEtswMz332KuBWEuuqhmXe4sl2IzJqNpu+Yp6IY/w6VB
91AoAu17DfyT2Dj4NTf7lJ2BObCOPJGm1GNSM1kM6ZQEwjjoXKVXdAYft0/gXvdt
EvAur9lngROqI/RmQjjwGPyimpZuyVzePAZgUKkfXJOSU18+87P8Y7tzJAuj70u6
KBBF1cFkBz7aH4GI8KjK9d0Axhy6fkvSr6czdmXNgDShHpi77MctSwc/soojZYfp
GdofFGttnkGHqgefunxRj45Se0s5maTKb3q1H9lCK785UCtItJxSbeTAru/brTvl
G0QoaVYS1W4y7OjvMOOGl6NRLR49JHVC3gkMtCcvWvB/q/Q9ywBGRneng99AnFKw
eUD3CK/cCxhVaN2DiLmCmPwqp4wxhw/L5KJQk96RT1PmR2ZadiXGCblaxR6gC8PK
MTshSfRsUGT0eaAf/DqPoinJ/2vTQpLj9BHn0gfNXnAzDYZlvNVp3dn9h+XW/gcp
sV5vIWyMKf68ZbtN5u0J5Z8ue3hgxKTCZcfLxjaPSJ/FN7U/sfcrD95gEzIjwMvE
J0ZtU9nJS44G6dBAgklgBvB8+IO0klekInEvVszAFGWcYk58Q0hcqIUT/bv0gdOR
VWeU2ym1tkMkIlls5s1jEuhPGa6afxDg9xD8XbN3LHnpEhCCj3uiyklI4P+62G+Q
U5gh3sGE5FHOcUMtgdH4LNI9uBqf1OjJro4/bU1kMLXsT2y6fXePLZBm3U+vuRhZ
bU3B9FivqTGb5gX64EfkjkJ0UH+qVOPOxvUK0VsjXvBqPU36g+aZNiADZPvuOK9j
c9q5cXNh3WDNCsVaDBFGxfb2MsbpYCKIOqav3K93V7qaby5NbZX/y2/iFKqmYw9D
1KITM1VfdQhKnYk3uFDnbZmDT878aHbBlJl+DNIJ31gmRQj+vv2+csaxiANwc9rR
WZnmvFXqdxNc7qkQHxWZ4Y2stFPPNRX7oNo8J3Li9N0C2fzDrALDpZgoEmoOp4mZ
hdB2TOl85ul6gudpbXbGckFUQrwzcUEapnxQm2MR/rELcCQtirgJEDVdE7+FknoQ
gPZ6DvUi31jg4EcHHf5YQffSLSbxQ5734IiD+hg1OqkuaRHQ7J/hCvB8EXEQp1WP
KqugEI4+gC0m+J2ROZak5TM9yyhLhbVXgfv3+zxI5HhwSfgaA31btPce0JhdhBHl
I1KhAL3IGjEuqxoM+kdaPPuyGAlPvoXcTiHGdtQYn6vYTUlX6m1ZJYqzOVxzkNt1
AbydBqOa6tL+lXLaywagU0Ofoi5MVkU6kPauurIrCwvNQ4zvTDhoLQBOMK43zHV6
ct/4GtT9bHIrw5AwvS2nHrpoALP0Aoqtz/M8HQiC/WxuSIi2GGwtFbKVl402J3JI
sJBy9ybPOkZrtwsMmCKwwBOKdqQaYSYQjR/NyGwbELGgL3yi+fD+xbZ8zJRgXoT6
LwMmvxePVL3A93ahFxlVyGmI4aTw3oVnxv35ak9XzSJkhtAYrRAZR3M65L3wQT7a
71MyW96XvzuAdstSo0ntm+/L5k1p+QeziQRmwaGnxTKO9QLZVyxTpz4gkZKhK4gh
XTclAmE/ehjETxpwAQzoRWdh9nvnUnpAbhBd3Rhpc+grzHpqZpFhJpzFxMh9/X8a
w9wDmLcSM85UxTCN8lomgrQYqNggm9FFceifszI1zC70bWvrWjO1KG5c2pIMeHVV
+wqYcMMzSnUcaESHQXOEQlNWU4FrzTt5hLaiMdEsc/QnDtUZM/JSdTHoDpz+h4Uv
DIKXDtky64gK4fQuuBs7iBeH1gRniZkeh61q30Z0fG+xqQz4InBbvocUXLUosD4s
Aa2nGraWMb8cbOrliqGMy3cbmgWxYzWKzR1EYONRsM/48qTbAcbJQGnUkgdM/kBC
5GnQKxQjSAJ4sZJd+7WTEMGwqf/bEv1anNWyaoYC4eVueomMu4VKbDc0yg5OsFXa
dqIdyUPMyACrXxRjpm6pOzjCVdK8lL0ayNW+tFTZr4B3KdoXWiGTxPCBX6hRffwj
ZNDM9/gTaEiCMYElgkZelM82RV9NH0js1JI348ptb1SumBJGDTAD+YhVEdaV6joa
CLSkuGwFjzQG6+UCiFp/LCD/OskDhVHrhJB9NHKW1MIlk8h+0eZIu/3OQOsW2v0b
2zBMjzerh8WZ4HpW0YjhZ985LW6muANdXkYpNoBPN1YMrN3bvPpAronNJ/GXYZLd
1KHnUkbKO3EinQqCq3fFBZl6SXZjB5Kq4IOYfWF72z1mVpExyP3BRc2m4YtSzi8p
Umv9TCzZhDasXQjFFwBjeX6j29ivUiC0MuiU9kw0kEo9kQii0PVZl5Yrce+OLYs/
Egk48GbwbRjeO+UbOmwCb5YzeapIEcqOkAQdwtNkNlfleWEXtsy1AhdLLTxO/5Lh
arvkgPWyq1bqpbrw/TsQAfgPXXcH8v//vLU15Or4/q1NfmntlkKIPr+LqqkF1BE8
cxR/Ql5IAzirowd7rPFvNgOoygJjOq5jsXEVrT1APuy1OuGrRfGKQoHTBagfM1es
r682yf0gzk3k7Z9i7fT58DswVVde+NG2QfePBSY3B5bXW46xVY3aYZIpgRgdEY3+
hvvdFRTqFShJ154wsANwcCj1Tw1oDOQmAqzKRBDjxDa4ei6aH7Lt4qpd9ygGwnMr
2z5XDP816Z3SHp7FHaz7UrUntKcNHIEE93WDkzb1v4Dm5Nv8HaV+EdtY9ftJlX7w
d0PeA6dV9HJCofmT9mox7ZkAmxOYuWGI9VWbSDJod1jO3hzlifZ32hyn5NWOA43T
XkNPBCBNVT9WQVRFv1FlNBdzIdShV1qkWowzWVUPR2IPveCtRZ+S2gPIatDCCxzX
1zOZ040QGTswyobEhUBQBUY0rnEdPC3AiBSqNyuwRMRPrENwRm7jzo3BLHDynyjt
+b6GTFtU5lrHVNKHT4tHBw+xh8zQpXIDKTqkznPGni16NuqoeLqAd4dowyI4Gy2e
Y3MxXQNCRUUZcA51wb6WWm/oCGUld2C+9K9Jf/k/aeGFwNYI5j/u7+/EFrfA7SHP
AkJY+LiFlrXgFWEEUW2b270lFvEtBnQ6HaCR4DRY2eiGiKf+Ex0FNw+7l7+fLodG
MBMlZWxafsdWluGD/t0R0P9sM5KQRmBVh+M40P9zCooPAm6RwgvrojBR7Gqnw5Q2
iNqYdEMe+WgcuVUMwP0sdfnc9rWeoapkuMzsXcFZL3YGNqUxOCHM9FDk8ApBduQ7
9LLrRcuwZzwJPCadn4GP10rdxOXL20vv54Lu0wx0svNMSh3oFwFeMpQy1p7M34MJ
KVigh7eAW1tk4boPzdBh40Q0t2XXixYet4PTqNcb3z++OUYt+b0d4aGpifq4wehq
CYHsfrDwyxTrrdzgv2BNMnDBPXLdWgBcBrH32dWB0y1GZuGKhRl3JZMHe1ApIWKz
J5PXlGDfxPx4y6BHYhrzzMnpEtORqTi3LBAQVMF/LOWNyJUbY9/Lj4ENTUaUvRB0
f2qNI6Usw/2Wgv3DBZrjrHJr8JMuIL98tXr26Zo41Lu4AbAPWew6i96byUsdiGis
O8II8F2lMp94rKcAXGE7MV1lQJSbaUoBAFB2LQe1NOczJvEjQjNIUgtvh8ViYQ98
n667bV+pHtoepYDXY7EwUO1yLx5SMafVlaOhOFnwood/ly18RFwISDQx8CGiZN62
ltEAQpUWxzsLVNYvf85OtInMLn3ZAyJrEsMN8G0k+ctjIgtjNoPBq+FVvjRdb9V7
f8aBiXuVUwX1H3+P5XwpGSGSwxM2G22n+pIvYzKGayWPrdCBoNFKusk3alf/uMUP
qMDTHXsInuQqhat8ktGbEyHWOZzqDxJCPAYQfIQDET9SUVXfqJVHR2FUYv9AJwXq
4+bWatN18V/IbgT71wUgNM5aFYi/vQXCjpLRjAYSyhTmIl54q68g0hJYa3HrtAmX
Ge3YSxnzII2ZLQk0MqxZoklxUhgMx7/DXRRPOm14zAm5V5sIaakih8NS1dY5T8L7
8v0f+XtFnJTmlbhSEbjUXhTutOZ2EcFXomDUkihfmhMyVIhJf+rUXdXR2XF4+hLV
0zFFigLI7d802s7NYc3hJ2adtGK4SNXwpQyMbORNdf1erO4buAWrEyVlHau+Ktqr
YmsddVezO7Ei9W6JWy2AW4niW96yqTSfSRIWsf0ZoVuZDmjo/JL9WrL9Pii7rDsH
qg2EJfN3mQNsgpD3zZ3FY5D4axg+vvzD4pWgd+peoUO6AOQI25rrdOvE6A3U/gXL
D9CqG+qGPiNcn9Ea9+ELeoohbGVoHcp/BSrJCH9Hd/atL3xsbfmohzigzz2/WFOg
uU9M+OVSf6VzEB6Mqa8AhCq5bLFAgWvrdBpbZ7XuqHbWOFxgCry1/8aZ8Wbi7ZRG
Ya7yVEH7paQs9pGzbg3Q6Zaxwn5JTnZfu4GCF461qBSbJjQKLs7bNLW2BwTQoSRw
a3VdpgiVC+erQrZWg3G381Ka+oebinNpf8AfxIyb4fGBCA4jhNMk+dh9PK2mxfcF
kda6OnR3QnGjoPu3IW2st2ZWiw0Exb5v10VL+Eewx9WvmrAL2Ph7eHChCVgDeV/h
kzRafzXLrpZltvv6I+IblW3f1pTAZhyHAGx7caqeBGz1F8D5+v/6Utn+ANATJqET
IxcQSyU7V+OpIkxYS2fG5BvYQRjcC/AAqtDX8oCBhZDI5AQRsj0Psi/QrkAwhFf6
ClTGxSx5W6a1uFP7MHH2YwWCMttMCnZt+w/+wc2EXbmzB9A3ssofr0pgrZ5k1SBL
ARE7crv4SQTpvkqI4pz/8QV5jzylYwP+Ag/RsTUTT+6JW7FYoFgqhOBGvEXu5K27
XpIdb+AtqUJVEMVmsPDUvZdJVg9jJkSNSXjOuAzaTnKzqYnTkKWRPA7gNdlrZEEZ
3/nbtzZsB3mDw8K/I4LyJ2sLcwtaUqz2m1WbIdkLFMerogQTv/eHRfJiGbeKE7s3
vbk8gV2B0rWP7GAqQDzpZTH4CwQnkFnVXRK8YhVflJPXmS7dX4Kyuj2l3Iqu5NRk
9DheHTgnbL8Ty7lIqqHhmniZ/ZrG71Sqyd3S2oiuZceg1DReszROlw4Dw9W0Htyh
N/43JscsQPDX7FvDZQ98gHnZDujzGV7zIgmWJa+vXfxCwQL1MGlm5K8v9IVUTi/y
mjBUzcvfiF48WDFCPVSKVszz4lcTLu9k+fF8pYLGhVh16609svRzqmqbfOL5GSKK
QzUGwFoemy1t9GN5w9HpsatJSLlDGnz+8YkwKTaFXqkcq9FBHzBz9y5Xmt5yGfbU
r2ltS/bLGqjNfhATihwZabG+C6/xkWL8iayRiffdSMPTXwqmEQ+kgaBuLmDBqOzx
oGUtJmK1gefbCayOMKsQF9YbhWe6D6yKUXMAiaGJekxkVnhRqpL0rC3cq0agty46
SF3uAOww1AA3eJBe0rsPgkWVE1amDEQ7DsZvr7GkUHaiojncB9mJ3LK4D3+3WP9m
P3lD/ey8PwPc/vqa1y/2emYO+Vc6K9oTvcQmcPTO6TxdPT65D5C10OaWGlphBMrU
DYnB9XsD5Nha+0EwW4grtioetccQOtwO82EVgnKpHa/QBBENVNd26Bf2rxNDBjN2
5vEGyR7BitjV9KWuIzT11qkDSxjKnAVRtZjf+rTIk6m5lpFkDz89IFfjYR94/Ihz
K6fQKOBjDTg80twgrQ/gJxVWAi8r5eiJL+ahnJ+U/e5zzTjGhOj8DOQYrciN2fxz
GsagtoVOpHAiiKD6jogbaFd6FruhCPlCOafYjGW+cyqhXWee53kC9HC7uVArPT7U
fgHGW1qEetbm4ne88DEFl07RzlIGc6+AmN3vOo0C2/ZYtoo/8MUGS6aM1wTJ1lzT
QTFEMPmiT0zkHNHSCEJph8bN+b7qeULPRN52xHHtgWuPjG0QhXdMQAsFv2RrsvVx
WsYQdhAo54oCbnVQpXsrB65xwOTPutquqzOHtkn0YbeG7AEGoWcQmp8s0Ft08Kv6
GhibYi0zftOiJQtl2xhEjNWdUs4QMLaWy87kMJyLdbdj3eeEQjbTBK9pr4PtGcMe
tjCbGP3oK0CnhV6qMKLLIhx+e3Zw+gxXyu5jYcA2mAzLEXr7Q+NAu2UEjDurgZU1
i5q4aYuf2xB6IGjyMHdqJ5S522urOIdkpADt4XCsETCA9NTo72Id/q1VxZNjOkN2
uV3VQigcTgaU/8zqu3xF7HuIZrD1mqKgBRBNrCv9OyWMkwMdy3cy67SwEhANwHM5
6akXglVNl8U6CUVrtsgoihS0alc3b12FWn5E3WfCtSPFIcaFiSl49BnP6N7645co
d+OQtNhtLbAV5x4d5JGiJjqbX8lvPN1TTUhGNVYyuwlzOGmYxfJJTQRnJv8iX9wn
sczmjvrA4BNchN86/ye5izUEnXxc1yDTg91ulcFeDkBeWtXBViALhF9KYMOWj+6Q
0AkU2JopUlz5rBDjnUNX/GNxWlKUXCf7WuhaZ0cVr4IxU1izItTy8fy0ChFvf/LE
eKl9w8pctrKoI6F3coH+SHp5J/lsc+IZvzjW8dDbwfmWWxw0H98HkG/VVdH44LV2
dTgRVqh0ZGGvxstW7i7xIcvndhad2iCXbUq1SN9IqfMgUqXrJVsSoM/3RmMyhdSD
uI4lhtVuXvVufqVrM5glDtS4q4srG1B32jGmbYEZuzxJRDnoPUhbjk/G5SFhMMm5
UUJoI5jN8uQnYnAN2BkFdphKUqnNn6dW9J9R5h5FltDOO+YyNRktEhqYLAuxw282
8c6Qpg6sxbK2QozPLHNbrObtFnrc+vLp4u1zjxX/GENCbi1E3MLO6F2QrijoKfI1
IiPhK2XkkB83qId0zcR2Zc/078GOjGQ0/jx+In0XpGmEOlvFvB7eweeA36FsZfl+
wFYvpPINyVZZBIQf0OQ+6LZG8j/NriFE8/T4mboJdLiMYDzItKmpfiFXUKvfqsoE
LT8TvKZr5lZP2K8v+EKkKoULI+XDq2kjj3UhYeLDi5vWdeFXYF0a2CgR1eI/d9FV
9gg4+i/gCc3AUHORFqGRCEiZKVRNwUcHetw7lfwC9aU565MAufdkPCueAFzaDZ8z
B9n/GjCVtIKwYLqzzJ81oFVC2r7VY5ezlYcH6M5UeXVueXbcdfI904tQgYO6umI0
LLu2LtEhcRqG0J4Q/0pRSzsJIhR/y0tDRqtjDRvk10XkyXfiy/UiO89UWXupgOTN
sp8kIgyH46rnQHtKQLDh1ahw406cC8fzsK4P3eT9iLtbwss1K0cwEgTQyCCC9lHe
YZ6Lw2sTPAcntSjZeTLUQDUgBGGDyUsH3jx/QkzTUW4tj1Zchw5DYBh1R3XqcN+R
MlR3CydxduuKSyNphjddvptnlpt530qjrGTlEenvhCcTmeNYnl5G3w9K2gj/Q0mc
udEtppMYrP6BiOz3SSK5aTA9I6kKggUJNSbSR5i+y7VlUJTqKcPf3A0nUdLRe4PD
F4pi18fqBhJqrduZ2pnIFnsEQxnJwvU/g309poSywFyprFg4eFU6qpZ57azfhfuk
F6ASiL31SuR9h8Ba3rS9Nz00bxTgM3hUMSnLAWqqOpWe3LhpJdRN3sqhG1+hRq0H
jLW6gPNA4J73/NqaFa7bKmnSbLg960NC5U5tWpb4o7p67o431m965tqsKZuHm/D6
t7j4+mLyfogENURbAg6IaUJAjYAduz8csEFLVwA6cZARpjzCYqY5e0LSjRmgCpGN
aK3bjgX3/6GBhPTvOFLLJRluazvkLlIkPpLSHTZwhwQ+n8X/pockKcYAjc6roded
Ol8y93999kDURHZ107+68RQPd0ZgFG8WtWhteFTJVWXDu5VR78rfz1san9IO7pou
p33aV7W74SPFKWZbysqB2ixsMP/qLXk8vhPpLPWeHf6B+vJLVBm6MBIhYm8UjsdT
PJ6iitKfFPCLk43n9yuwuBzdlUGKAn+9GZG8CIpfu/useuv6Jd8UIQvDdANhZoxK
JxIzUKDlG+eXyCxGr7LkPGFxfkpgfMNJiKXa4JkEWriMf8aaMDPnU7mIqebKwoWu
VQqmQZ+Z9vFwdVAmdO90o6pP3uAFZuWGvPKmrytHLrx0j8reIY8lpv4vJv7AtdOo
reowjLWSUk4i4R87JO+1yGTaY38TdXqY/z39CcTRO96Hqu8wqdwyb4aEbPD6aEkz
e3yKZ7QV6eUQhiAA1IjWB/vTdEzWudo+WKYJKfiYQrBHxHyhSMv9Xn+AF6uKRKYt
4J36k2ziJsdVM03wS+ojpcabvwoCURpjKlXx04M4znSAlzjMFru7V/y7Q06KMZs3
F+8h2Y9F3Toy6C+7xfCImFxq1kE1bAr8H4S2lnhziSM10Qt0W1zavDHMCCG1I0Da
8h4QRFacN4xukLPlGRpTBROR5bOICsB358kwGQDwSf8z6QaEQn001DwciBH4xFmV
iizE6y0THogURYuDQ8iON1xk0wtgAW+8d0b3OA8AZhhLqa212i8k8avzCV47pEWX
ioeH8gH4L5tvbJEQtvA/JzJ2I0Ho6nfBgZRj2tptkHx7gIU2Bg1Dnd63S4l5JbJy
X76XPJfERDktmYFeA8tOfnV8nci1bSMC0LmLyHZl0RLpDM4oyuzoWxMhz2Z31OAc
y4XHXXq7Nd7MDewUBx+cBxTniXuwOVNh+oYIuElOmwIqI8S7AnXUrh9nM2/gO68a
2g6HBk+kKA/m8r5rfN9Cyu7mLevTWcb7A2k3MDTfdv2SzbH1HPYfxh4KQh1RPV0n
eijHgmmz9sPiMOM1AH4LtpO6wFoDLBAxH7g0C5KQUjf9wP28ajk7ot3Ic/v7TTWZ
vHwJZoRXvwfHqweA1uIAaKWyznXqNboquauPah3mP8zl03Hf4pKl/XiG+IyB5W+8
3NFCunBhdO0uBm5sYf5F7kJD7Anecx6EQ9B82bgbz+DupU+NyGPdiTGkYEb/6cN2
N2vBURwcQXA0bQ659mJH1AEOjZXFCe4KOBzpRHm3SAEha1bRsXbTHft09dne5NNq
7isby4q3f/T92BYiOAkVmRrUrayZuZVqaUjATs8BmnFdrFWdkW4YL8SKo5GeKUvo
j+dPWaBe9nlm9du4yOCWZ6afTloqHfewwYbpRy3O6zAemmBwE2jo9c58+FFn6hYO
EoYnEU6hUX/ZFWplnfLQcDRjcJfzxNu5PCuYSOnSvrxal2DZliR5j5L81GL6+FaE
rofk0REXTitY2Vp4yxNSVOctRWJbKA0tTe4qYYKaqvqG1DYkk0FG1iIond2HoZ4P
eUHourpEGD30SDOXkKKOkXkJ5EGN1mGU1D+VJoresQ3lyDUlwsJ98SURiEPt4kfG
HFNDBAh92pQdqBwAfGqHnm3nOLF1rY6w1aqgpHfbAnxFDLsPDLWa5Ee4T/auVvpy
GRfTSTXggguchEeO9YVNdGSZVt8at/7oX3koyzhYTSApSCxXwpifSMWwrYGrqQxg
U8eJjGfk/GCJQe2vMuKgKr8n+KrY4eADf0roKqa/xLNQezPr5FdIZMJcpqysdo8E
fWTgm08aVImbcBd61VW28ZkwgJYUZqYil0SvJEYRDdx8wAjdKhL6H1JuT6uvOml/
My061SlBU++PMNYJw7OOSabRqpAyq8BdgNg1SPHXwtMG4BpoDM0C/LXelaWgOHto
s9ri2EnGz6h56cTTSd5tOgzeHjdu6teEpDQTc//o2/utSo9YYUQrOSeuEH9V9dUr
Fx67aPeaK0oNftn+rrtPiBErCLmdotagiKqoKdI4EJzYetxgidHpSlTiv0wat5Yy
14jd6J76xxr6HQpk80ppJuHHAcc/HDhfADAX/IuQiW/AIb5TwJwxY4Xd0256WLOA
SEh5SWfyreIcjuPgLtfHNMD1cIJ0vuNtP59Y2oG9W3saJnlLs0ifO0sfjtoTdvvs
+Ej/3QvsKksyyCPk0XF1UKXEp8HT4thSwaplIlEHFqnFzsfCrYZ72McNbeExVv7M
FNsO2/K+3lPUReA0PlqEyvQY6Hdf3pIDynrZlM0/i4FkmDlQfCdCV/DKc2ybcVd8
dj+OXEqCOtkIW+X85I7yHV+6hsHgBUlanzgU2N0Kn5CzL0Dgc8WaXCAPEjesNR+H
ee2inbukUTE9tdDdY8MWM4XOnIP2No4JY0Trm66S1NAB3i9GnUYVpTUURclsQqai
2jK28jBsuKiQoiD9xLPyHvY0mFaG+NqxKsY+B2Kh8iWKyWMbhN847p5NOzaAkp8L
qrCnm1kLiI3tEJI3B6HtmWwY215g+EiyBBWemL5frVxwpR1q6Qhg83Px4tT0cGQl
/WO1txhGj/QUW1dnxrUZXaExQHm77scBPes/wNfFIl7+xaV/I/a6BZ4bgwH5QTCs
URjPe8JoyCtidSjBr2er9J3kUiTNjJVbH/IC1puMfeTaQMDayeLGYgZS6qZ9K303
AgcEH57RABqhsv3bIOZhuNCc1NhkECm8FKRkzT182hUFRrEk+WqTFb1TYnhX3M2r
q5WgdQLdwic6vEFmO41t4s83HPryJyvEWpgq5eX+Tn7vLXJb42/JtAzEs+bEOk6t
GjG/gcV/lT2JRuI5mATZ9x6qpmUnuW9UV21EUidQIs27AaaUcSQk+1eWn44cWOUq
gFU50VgRKWbcTdqEKQ+sa2WN8xm6VdqQKvtlGt3+rohq4Aib8B0eOBSB11MKu7yC
vF2ROULRxd/uQc1HLNFxK7DISW6TTjyPyDzk7Ct7l3anmYbBXgbhlHL1LlROK/JH
uR6gfRtLGgeJL2jTDDjXjUV3z6GyOhBgO2WaKWQypgVyKl7SADzdF/p3oqivBMcR
l2aPo9qYuiMfS4eA/lZ3kiYo66fvnMncS311+PoB9rAEbXAQB0hbSp6hoba2oFyP
Hb+wtEtyOyanuEQ/q6tmFlrtog/US/WHlxCSZEN1DCanJ5MN2VJDA62ZBISXJNva
y+pM0UBd8heKKJYzT52HN/TFcuQi8r1teGmC3rQE9DBt5JwdV2uQI2GneaJcsu82
WfLuemb2NVWRF65PEx1eXI7SbErgGHwnFAy3nmeww55ImjSRuhZZb4XYyWy/J98t
pYo/iExoIdPN8vOBSJisxzVVR9IZsQI/pPGkeHEUkBE6Iw8uyGdgbyso0RT/QqCj
LRkK64F6NYouOxG9UL9bHtyOFumLDNtpGF9YR2ulWwygFaoeVQ0URTAfqVQz71Ce
LDe0/W0zPnKEZ20tnyreLUBcFTETcoGk3uYpa2SK3f2ZTwIwPUmI8/oarzlRH8r3
xZevPUpuaWMeei5dQ2eRAE7BiWWqzeL4nOxrLyzoDzFCjQo/+c9WDqVfLnohWCdB
b/NzYN0IWJZmHmFhEJO5jmCifyZMO10f8MzhgY841/gK3Qd9MnWHf5uQ3dpzh5h5
/SSr6WFUimQQ28eFyxaPvmTq+lRv8JdN46DDEIDW/HWoWnos8ru4rV5FtiAOq9yB
40zbNyzQISbp2bY3v/u9ZoM9DFPFltl/NLdEaJvKnrQ2FVrD+29WlttQD4cApZqM
NCIPcKcQSLlCZXiQEZFg+1PmCn3zgAlYjTvq0Ajv5pyArLuFuRuGjzt1M8DraoJl
zAV+dMeADv49NKijP4HUmZVf3Mv9CafoIpnnjWjmDRy+dbPYIueH8zzm3SLgGcBt
eQZljhDZXRlpP4rmJDdeX/Q+PT5pIBN55Q3UwkTsHWmaRHvhDM+b52w2OG1PquJd
RKtHBrluFfywJvJ+3Yn40IEu/VdqOQUNhTtnF2jYW8s2CyhpNYeqHg8GW/8MSOCQ
qp2ZgrG9dYgmC5cBOZK60ay0W7RZVW5qZaGSLTACajskpf2t5Tw72/3fhqrU40tX
cL0tC99DuFAOyAqWNI7RFmZxW0BFUPGJaO+SemafERZ6hrqW5f3SkUzjtmfOFDXJ
lQyLid6ZHNByu8/zGhzU7nxT+UfwpW7V8o+PYLWLzG1cq9QrmTLX48ZPDr3/k2L2
Ro1YPwfp6fYnHBaB/Izbj7xq0mlhgWYqx4fCKxRWQSdY6XPcrly8GXFye4EOCJMt
f1g/g6IYwsVBleasstNB2mKxRukZY/Y5dtO8DRBvq55635WZ0rZej0Vz5biiPgWS
Nj1vdMpGuvd06tmntGYYtiLgOa+xorWoHnHiS6j1vLVRCjaWftB9gEtEkhxNjcyj
qIYnpqDHFJUWX7OjTPOETWnbFhT5WYqNDDleowuJYqyO0mILh5wq9dNcxvs7LCGM
InruPGKB8RiIorvOMwJEY73EMryGYpy1JaJIBwZHqUcfyETF5wxY7VMBxJ/spMkx
jo3zSEuIsLVFr0aXlHEWybGfltKI+hDAdb201wNcaepuHAVBvCZyn5JOiOl1cvAw
Y1qSZMkB5cDPg4MzGvjxkLoI4bmvyfKwWBMeUaObvPY8xGL0pG+TLR98iKa6WUUd
sHBWZhv7w9K+XqpKc9944o8W2k6Dm6XNW4mkmg2udATQ0YOZ/nrVSsFaFS7atXMv
vH1l/hq1dwIyLr10i8hCyB1nacVHtGMYKeBkf171nyPW1NZisgCcRNJLr09aM+lo
0bNS8P2nX41rig9wbDHIsRrOYNTxOd78ihORxUURRD2ApbVf/tv5M5MOoDZ7pXtf
4r9hMelItRm6au39dUxVbrb55FbOjaVNH8XFPe1Avny9vEOPGSYgsJkf6xz/1I2M
UhcuhDykfNLiasveqke7u9Two7jnWBn7XOtRwcNtCqHvnkPAyoCpaSw2+lKc5wx1
M/R3E3w2Ml2BsqPQ+Qq+W4U+T9beWNGOsGogbAE3KXlgRzv9FU7J1SLaRcmGezX2
VN8ZKjgRtNf1eu3tfXOlcvefmBbXlf0pEPoXKodKwKc5HbqEkqy0QdtuduR8cEsA
hk+FFjdHAucPtYAX2FtSvObKCoCnFFwutUR/Bqow2HfW/CniHsqhDZ1nbwJzGnoq
fy/cl1A5dxD5QrPdMYjpicMAHYjj23Jq2TKsdTtNMJd0w/4UAOct/Q2V7wneRxYH
rsCD9WiYqE0joqw5K6FzIa1JTRyUFPHE2tqeRqwmlISfqZKhzMWP+X3p375WNa1U
8Q5CXEnt8rKD6o6/hwcB1c2+OFaRHf1tvD/qif9Vmkr513gLETcPKmgBpjos/hIC
6utAoWPH7WsJ2nH0PSy4V2XwvDewwiu5sxqqcL5bzeqW+zCQMabCkWCEKBU1BXpm
4zxYsf9P55SNlLgIpx27HjLh8S5zL7J0pffLBL27jWAXsNZPJCwr26ON4XGl/E15
YB0BB/YBLkdiAa1jTPmH6bqcDClcHumvcrOto2TIn6RbTBNu3XhLTFT7f69uLzho
nrKCEUpFKdGp8neuidHVMSg8Bg85nES8MX8aMqSo9oCRoRAOtdEwqllIRZqPGcJi
mStG6tI1xiDTbdEMtVUJwmY1hVNyLQkKWVVE2G51Kl7zMPiuWL+hz4LG4SfeyC6d
H1+wcVmML1JDEow9HgkHGmJ/K5+P721GsTn1l6do/QAH4r94VM1lcGlHBXZLGf9m
12sMWqWHrYG7Ubhh0rWoAfYvOBeTkctAC4nCict/L2m2g9VENAfgpsFqNJ3kqCjw
auhNceCqlUPpGATvxCHwjTaoSOz7Lj9oADrAbkKoj7+dwl8U05stc7Q2g1D54OP9
5uzJnCenM648kPlDjRjs92iuRTqj7WenqrkaCMlTEZ9ttEiam/2e0cjAgy0l04c5
pU5rPkUvVmnkJtq0P00/eXNA49Ec/pghqV9W4h5WnRPl8rEMJn9Ug5wAtZEnoP1v
Z+OgYw5WY+wvzGi71/2S5+Vn7MenHUJbtUMg/XWjeb4lWIrnDA1rGWh9J9GKnYpy
HVO4aatDXZ/sYH92w2YyRQSqd6s5L6b0jq98zMvd+0fk2dV6kqvinQdHydOT1Z0p
ls3/z2EEkdxog/hCMNMglU0rgeZbBQ/WOK/fBEq8GaO+2oozqwVnf6YVnV9FOS0N
6XrVIslKnliWuRToDKrw/QBC89d4uSGPCWYfgHMCfF0IYsI30hkBQoQPcBHf1+Ba
26YsyJUSD5q48GLC/1Ck6mp/L5VHwPkL+Kdhd6/RB/asMIyazPUNHKkWqfkBs/jm
0PdxTzmT6qQBS4OAZsMxkTrINZRaFm/em2fYfA22WyP6qZ7oKdbYBa72Zgqvj4DY
i4hHeZnMDFJbC+OBAjPpHlNOIXsgU5rdwIfV59DTzKO/LPjQs+H4j8fFeAFYoXjy
XkcBvWiwmd1ivd6vsYrNXL+wvviv22iJ+NCKFOF8vo0bqLTslY7blAhE/RnSi4mC
5xo2Q31MA4ImsCrlPXDSl1/UqjVFOUzVlg6gRLQ6uCLk6iXOfl+Ly6A5dkYSxpF7
GgtN+qUn8dEjlpvNvIRcTSQraYwx7pIolbuAHqWaC/s8zrezoS2+UAUJRVqRbTto
0SgXcPHlYBHw/fS4VndjsUKwE6vrLOJ/Nkqx3vl/STv2xTBljbm6h76D8OKjNiyS
ayQmD9p5krzQAoD6Dk2q1x+cdOHR2HGu2H/5ZlxqLuijxYIbE0Fe0eAUFpsiCRqp
P2uSvddJQn/w5OZS0YUjXpPx8imx8usVgififu5EIc5H/fYNa7ku8/JWkJjLLOsg
tcDm3xz3AXRVLt9j4PSNVIqTZEJNZYZt2qPeo+ed9y+2sKrPjkccZHXS1TszyvHK
xXUp3NxbSTPX38SU9PwHn0oqr1dWVvxDACAA43iT4oJ6WWzkOzigP+f+TZPhB6G2
EYpqA0yaNGepbjzH4TkJKHlFv7oIV/AEp/F1dfv7rXO5VeFhnCtUWFfcCcMPRW8T
dhmPEDU7bFj2P8b4eRXCqi2UKvVwhKLKH1XY2fhCQ/HGqNdgMwexmmaNXooocS1i
8okkwySRi46akcpEn+VauYScXbpbcuBkoYDbZQEnbVjG2iTXU32vTM1J9Doc9A9T
BL+tjKjz3oYk4NA+PaqIU17kI6zu02E/CdpE14f6VJWuZQ+V3sCLONRTzav9BR3s
+Y9HL9SL+GLa21sSHh0etDVl86C0qIkuSfDT+uPRtfFMr5fB7CW6yq9dVZjLNxNZ
OZbK2twAwTaUHPgJs/K4zfmgcBf49SMgKN6gZ/n0cT/vLCZfQGrr1phGIJeUryAo
4fOmXfJh90bX4hMgh3uof1ADYvfmsg0NQSRBwcQEkibdyBd8Ipnf8AJioy/X8FYE
nHYhTv8OjaUI1aZZgstBHBMUWuHbbb75Bd72nOaaqKajzNZLPS2+xNKW0dmKH++L
8b1vQln9wzOX2W/8A7+x+rNVU4dQuPwnJ6x/Rko0uHvBtEN4fOquVnl/yCIasF8i
CaMmgStFjCab3alRdWvE/vquqqAabKM0xaY/afVCfDojsM5qmDwTW9Y7e53KBGWe
BtF4pUp+Y4zrQvRtvzwB5Gy32QmJO2YE1VB2e1kagIFDuHLwPVINiZhX3sNxUylC
Hx6VeydI5dCRC7OW4uO1kUISvX6gZCTVK29L5FGqrKevZ/Mjnu9iBoozK6tlYCAW
YgvpeaYh0IWdlIAlAGXXqOWQ65maOU+pXujV5rYVl1ZjPzClL6OqQWxnV5LzMiJm
/Lbtx+ZzwGJFgaczwxU9joPHP8RRTcRbS6VewrEh70b21CmIhzdDIubgJtqcNXck
arlczTapyBWET50JTxFFuxJMQOWZPdghw64DksL7wS/i0bes4ekBjS/s1vLExUiI
pZSHXIE9ch9YafMHNIf2tO96ciGkrJUmSbLl4zpZQoBZL0QiW1eQn63v+txmu5ti
qYV840E/fEJtGHmmK5Th99n9hjf0wCa8DcRjCLSw48knzDUTSmzw9A4T4SkKLG7K
O7ZowsdJyvezO2psuvqTXH7I6q5pjs04ZIYbgY06PtW5E6A69knwiRcET52XqOtM
dHo2NduuHG7sGJjuW1N4SrkQgGGk9hxDQ+b0Dzv5/oc2t9Go4CVw2YzCmiEt0wpw
cnvQliW/HcNcjr4hSQUdGiOKPBIF3j3F21Av7FR7ObPY/DnsIG5IAU1Qa50QlkCe
pUZl01IDNbOldzU5xaqPDtrqy7UlWd1AIg3DG8V2TWL7GbrbGzBZZgdsvvuLG81J
RYz/Kd1+flm+SN9Qam2DvkzabSC7NXdc5VDS+ULBH2B9k25pZFhgRV7V2Yb3mzyT
5uAx7jaL4vZC+aKEz6EHdddhQx55RCnnf/2ncnrO0MWTjCF2AXwHfJ/rm5WITltx
p7A3ncUdHwa56sfIvUr1auvTC9R/vo+S53vSIKU2IZk6xqVIt9DSF5DXtmmXxrTs
5/FZf3Xw3sXb+wrbnVa6KdZCSl3f8GPJnL3LSNDsvLfT/t1oNUff72f6gD1KYHR/
V7ONc3pyw35Xa9cjZhrFX96V3hqdBSn6YLPppbF9V0iI6bmlOEkVsaWiYFiLjKZb
ZT8lT2qIlhNzI8d9+2JSnskLWHKgnyOaNZX8buaJSfBnpsmPtfx5EA1FZndbX8K/
L3l2881b62X4SjCVKWo5DLJf/AAkTvPafqk/IK4hMi805exCVX35qxZzaKMLBIJi
GaEyTD+UzYcHlI1raLjoMxos5C0UzUuX9dD4fpVlwrTVq+jn7q8+ftvgn1Ij+LeX
qDxBouwMXQxyl2tRng8DACF1cahPqpUK3w0GTYMMagyXla8kisSlsLS9MHbyGRe7
vpTxOoHZuJvfIOOAvKhlNXEm4R6sAjYDMmpDAlkz2nbs2ybMAYygxaQsbMHZsIP5
iei5huzcsCNZz3007TVdbImFn+1GmXe50NlZ/lvD5XBqoJoV2qyKdADExao48oTt
97kvLYyvUM0sSLJRdSq1dF/UK84asNXzJE9lZmS9HYvAg8bfg2ylXpDG5YfzfY6Y
jh/Xg5r5X0SrsY1YrAaj5JqL7epzd6IR3I61tUVfS8GEsigVrqoVBozc82EFRGn0
d0CMBvlvMcrr1urVabBkM8bPoiiVJwsZ88nCpUalsaqiC6wNrE2Eyw2QSESIs8Nw
brmGf/QfikuD4o1KgFutrjf90Yku9xLYcQ/NYp6HXlXij5ylTf91dcRT/bnFENjs
W2TyiEVJveo4QIa4oYBnRjWqnMb8OOYHdnxAGfxRISWyMhdlOZq8otxA7EGnYcaS
rOmabHndkQtyM0ug987NEmgVEFyBvpIXM8OqtmtmR9A+gb7dD/9s7iUBdFVHkav1
Uoio5dleoFqqL5HNnNCwqVrrpJnF9tBuuxNqjd7djYyRcblOPTYXTc1IS3zxcmU3
l+qPNZHTuNN6iPnTLYEtGAQKUuUM5pewHa2pKUvC0bCAFpvxBqPV/IMtbOZtGvmg
/wBFxpRMRc5v2GnMb7o3SHalLN/gCQTnWjZBgLDUe3LcFht3KWXooP/MDVWlGfRr
rTnnO9LPENJjvHyskeKIkPqNuyzBshlc0/DonysUWjWgwDY6++0f30nR+ZQMmJfr
KIPMJJCu5F4hArF0HEjTLWHPSEDSCjlkZ7L8pef6KGyKL9TVGz78UA6digc3QtBn
K7zV9mR3cohKFyt4gcqWEZvzZL/g14w6PhhJqOR1Mx1wNAKP//nZTUhwwiy+5Syq
97fmLIXGG4Kjvdr8p+PDM/iVDqO3BzmOOGri6ZbbTLB699yA6PE5L3IS7Enkpl1+
Zvw7GiaV6n+s+PIMJDoZP2l98zdzPxwmUyTVJmMrVRyFk1FFVXd5jn8Uo9cW4+3F
XNdzVMTByN3jGC4Oq4VVqKh4pacTts0dy7mT6ILl1m3Jsrsv6uB+n1qAHJ8dRlrv
DLc0K7or/YKN30k095ILPXSPxRkwyQ+oVPw5VErqGiqLt7+iuCn5fcyLx8iAK5tL
oBc+sJGdRYzNs/RcxjPGDOAuBY5fU9YqqA0GviX7UyrlAPjzc5OEk98J2EWq0Lag
VxOD8a09uiBialTFQXR73Srg9WPVL9qTGGPOt72Ntr9dGJ4C+sxmse2zIbNFREpz
BBvSeZ8uttZ9D3/OcDH4viOinWK+G7rHyZkETxL78qo+JGBJIDid8L583aa0dxXG
+jP5R3J2RG3el5oqEA4PF5glxZn0dwNVYg5AlfOfwIknkI5OgP5lanDpQfm4I3vg
fxAWwIv1/AP9796LESQZeHCgw33iYt4+OQ3MsUqugFAuxZxmTBxgzvK7T9VrnDPX
eflvven9kubjNkH2UXKgzpnSFLXG9IKcx0kNzchs+p4StZ7DeLwmjlGZQko5KmeI
dqGS/WzvAIW9oHaVfsbDfonLR9ewdKzphzmgnGTqDSBQNgsK0aKKNRE8Tn9jbwzc
1M2tZpKjv/JSyLLVoWAcQH7exlOyY1AxRytyPuKjfDGzPYVCcwu2JQuu3+wM3/oD
qqzMvABZPNSj5aQIEzXmyonTxIUGNNeFRuj4ZQAmty4h42HXS1j0KKkq83AC5yZu
US31wGwHDASGc9AIf6oCucu6H8YXJpavZAakaQN7XGAQcvDWgjXLZOrOhpYfErB+
YDmYEjFkE0ZkOyzkjoO0Cr5ZG4skAOWaMOwm++IQzPFM5D8m+Q7Ov1XV+el0A7m1
aEl7i4pQhirLoERvxQ8sTQZOfUGYczY/T9t43/y8Fawj1QISakwgRAxvVCitXSLP
lDOAuCcLxp5HasdH11KyHgstRJEcjb8DKJuoNH83aIlwxbrZ09b7odcAn1DMrC76
FK6YRF2Wr80jmfOEuJ0IvlsRuY+OQ1hOmFV2CthoDGqBqmRg636zXyC6xpj4ZdEK
6KvuahYppNNAG5kHVTtknDpaSYYj9Vj7nNPF9Zkxmvcl5gc7pQtIsT2DozQ3Z8Yl
/uE5/CQ0v9KfQwIJxIUm0kLDL3xF5gf3CYaw8tHoPBPvGtHTEf5zxICrh539mTVi
lULbghq9PNBmDUY2snwwvFuhrN7NeYDxUO+7VtgwrodThbDjMTHrmE13XzQBMfRH
j2NpXpng8Wab1u19Va5EM/Jbdk7583Z6Wl3C7LmLFBqPms/096D7/G1Nas27svhL
sPUUG7advNBU6wrTnCr4iToJebX+FZS71en/0vu0zz55Sp2sxWHH3S9euUGcy+PE
xK/IoefY2US7oSCU+UVi+6xqcP8oQbMF9XavR13PfQ6dJ9rztcQrt4T0Jwq3JT1P
iJ8QohalkoeY95qIstVf7wHrZ+8EXT9KLNs0y0QDzspR1fq9ODI6RbfKh4+Gcknc
r2I4dRRUByDEQeyRPO2pRb1V0cXO55g28LhjlQ/YN3ZWNoVbYrHokqjRbxVtuVW9
ah8LCIA4xfU8k9p2PqdRWUvbMYr/gES7FN3VcsSHuMMyTxnc9cfm1pqzfjARK0M0
vMXHszXGtJ3pL5XcL+NZTg6EjupQhnde4K3ygxoEnAG/irSXfZ1VwY0iOFrE+BOb
TTt912v3AZEzj451yUF66eZDTd5Vp+fea4z7u9+eKq7w0hD7iarZeWuo/5o2qXe3
BTCVYBEb9u8qEpR1ni69b+t+ipGOvzplji8DRgf15ZwuTLVy+0otngN1w+9AfNFB
nKGEdRYyPMi7OEWM/0GtN/BcS+ELIkd7HvKU1MTPBzVt04hwtajh4+Py5zUWrJ2/
uqbIVzk71TiPXJvYIzCpA9SO0j+HM/vohJAQ/4HM2sJDnwq7mATbz9Jgyvj850Gd
KTotlgbsF8xmDovXgYcvlUnh5RDzfjeWL/3JH3NtPpYPoS2v4JEKoEzpyyUeYWoT
tDGvUExGNS372bdRSRIFCDr2rRLRmbO2pHM/azqNQWUqIMuYJDREBssayVIjuCCU
19cwt9GnTJh4J/UfYEItzz7gCrDatRTXCs8HIXla8voM2gfmU4VQ3MEHmbkjwP8+
OhpV8ed7JOJ6jxfbWSAQrpJ44hUcTHiSotQIK0Ot+7YB8kx1FNKe6woyH6eqvOoW
wM1qvRiUzCj64QXhkUB4MkTvxRSRhvxCbfVYEaEx8mfcul8mg1C/rDcUrVsfZEGh
cywu8LUHShAGUMtB4SHCHKrsskh0APboRho9TG/CjO/1Rlo/RBKYyEV0T5JiLJDB
qO5ljwZ275fggPG732umTHRjRb+UKUrwuC6rno9vhLW1IuqD129AdJSVf5g7AWgH
ER1uQQ2VxEki/Gy4gtQ4oPMuj65UKjztblPe7PX77PE8Pl8zjjbijn6V3hG4x4hO
N9vv9YYP5l5bQadE/higTSCM2Is3DeuTkJhevjX4VoSFD7g9nv61HyTtP+PFKiuu
ekhmyTqK568kYlL629vHJsgqP8wGTsXMogAyzIp+Fsqiq51WT5krynMv5zdMHfD8
wdAcpuT6xHggpUdLC7Rm5gf1LgaFvwMvwg+D71IlNe1kqMMZuANOFhoHTFl4FRp8
HnzejQ6A1j6yWTlKukatH6WV2VtwE5Qc3abDp+63voPz72iySgwLpUXqL2m/6XlA
WTMIx3v+FlFxyBs2+JZL9BEBt1EJ2fwo4FUq6cC27MuOwZSBX212TW8ZT7/OPfxm
mUhu6XOfrY+88WXYsjamQZ3SlPFah/BzHezGwtUS9t+rrkgzOqA3RHnj2AnGEmrQ
iAfQoKDwJDZXOrefFa84gyjyqIN1EYh120Puw/3ESg3z432lv/PVF8v+OiKZNcrS
S8Jau0WkntTJ7nWxnA2+liy/3ObdQ8iIs27ml7Rg4xVxBkR6gsz5zcvxz0n+tAIa
916a0Ja+VTstKo0RhOYzKUvue7skqaB3qKFQcSCsiKu4XofdAPCMoxhmP8ovalwY
WuPZ4CZlJZfwKOlyfqieSMToGbQL95qmmB+iXe3Kh5wx4xNicAw7soqeZ6aohEaU
ZAaOgPzDDoGv0eYzY15JvvwgdtaGoazFXIf1OQgx1QKveAttQVkX7/TqzHEUSbTk
IGQNhRo4UmdSSQo5aFngHCLoInWhjGFvW4nY+Fewix3TiEIOz2NFY7u0bKBIsS9m
DWDMowSFPfwyiG2WZwpjzCGPuyWlQfuwfxbAA+gbGBZwqszuDN2qaGlWvuwQGZRA
g4tQ/OkNmuxcpbUmALexBflABbMW3r/D5DCxrxkpbjqMyI4I/CNGavQESYIJBIK2
HJdX+o+nfWEBgORhsZbzGtV6DuLlxYnDeroQkJZNN0fuGVbhqNFwc8inglz8OO0E
stt4W4y+0QnWBYMFHHYlluOwf0gpFbaS9iHu48Co3+oCJvSoco2rA3zSN+YjTtn8
dijje5L1W5MOTe1lNUoDwvE0mxZ0pAInn85epvR4ENKhHrWlnowdiJ0WkW8bs9mI
Xpsty264Jg+98oZOfOnKqtbg/i7sxdLdbKpqkfZSFuaJUnlUzyezapzKH1e1k6aM
MdTkZfYvIFN4fVn1QeO42RU9MM/0z4F1urNAVedvoqS7WolOoLhwTjmISFVeNkOA
nfPJdqb9CSPwMpF+CRd4CksUUGaNtpqUSA9fcMMwADMWlCAqkKLtVO49Ag8eclCX
85VD23kz037gaDs3L4JRdhlH0Ds9AsOetvAMkNlspW+v3oPOd1jV6jJn7n8WSEt2
swKWUPK9TUlQ4Hu4f3TqRYkY12qaCxFX3/pEEXIdaw2wIXThS+E/dGlxDGb/LcQt
QXo1CqoxZkfdywN7vxzcbzzfOAev4S4YEK3UZx6gItvVkD/cdi2LvZxpnxhO5uxF
SFLT3GlFFFrS1m2kA8hyNGGA1zmNyOx2ZGXn1Kb5gNZZf1HtBQHmVXXO67I7ED7z
LrM0aXm2C7VAfnFUeY+F61a8xhP3YT5fRkMTLcKhUgexTFD9DzOH47iUS3OScVNd
oh5cwEv1xTncQEXNFM8aXyVOY7QliUBawCTQ1S9fQAu523itxzdcicMp4fCYqEUE
m6JJ9MqA9b8XPXinwhXj6mO4gr60vaaHmh1dQsr8Jp5FL5wr1eGaCAxTxS4u9KhE
5SbEC7ihCKqT5zmbY06bh2mizSAXgMJXu8YXB1k+A9qhrgGyiTgjTWZK9Xve4hik
m1iSqCmQwhqI6GzXbgJYqJJFl9vlRa39xpCHsNlFJdc15cIZEOQRed+Ezn46kNX6
L64LTS1Re+yRIDAQrcstv5tCSuWOP4jLCeVOueXxxQpOuWk3xlQnX32WLl9gWQQM
rxj03yaafGsQ6JiVJVj2AIJc837sVfeZ5htLupLVhjYEj8a7Lw/NHxGOU42BbyyE
2JrQBLDa7dVvpWCT8dr358ae6qsW9s4/qv3bL11mtXl+5PtUHllCG/YREGt2pgOV
U9hrGZ5oDEWxPRUFEgqTTeLY5ZqxjOVS0THe37z4ClxdktacXzuxUPZqjoOzjSQz
e62s4LOR3AsLBD6t/4p0Co/Lei3keS9OBwVh5KqOibiNOPhwKaDU9Vw9OH6Bx7t3
XvqqP5V+W7JxbFEQ1CI+xQBHsVc4A+98S9DW+cTmWK7skSFDxjRUe2dCj2apWQNF
bpSNG71EFYIwj+rC27+2+SWFtZ2ajbu71iJ36b4q/fha9M6eH9ugYuvw7yGyplR+
MmtncRrEZvqyonoV+FW3+nlmVs/7QyuORqP7CsMNETrE9Ohu6n6arZ4QtPFxB0Pk
kBIeTinLXTEdjuzKdweKpkYDY5evA0eY2U5XgHAtqSI5R6u3Hk+LcPeyQqxpx+Fk
gNybuutMDiyQFQOLPbx4Ojltf4EBtESB+uxHS7otZoW0K+d2zz4U7anGm2ZfBHO0
fvkAvoRDbMJupgYFiOkDiyL3VBdYZWggCgQ/A9N0M268vKbkV9wgQObFgr2eOBhp
66KTsfTSPXvg6fSOM0NmfYVhKPooV01dwdOlAEtsaWgYxVLZfr+EYHd+ciWOvuYW
iYXanrg2BLZYiwGPnB23xtiVnYyZcAgzIavL7Xh2wUZ62VuTv5B2OLWicIAD+C1f
ew0eOZOLsYjTcOBfxAFDqj3AdkZ089wVeYkimxra8vRDo1xTRFMbSwP1/mhOCpg9
Ql9KkuE/aK0l5MRRVsb1/TFywlO8tkNIs3ZlHHMJe9b1K7cAcDMmp24v0pxQXD3G
/lkda/qPCsFpdeb1SXVuhiXrJnt53E3f//kdyh6vo10/VgSmhx+JYEst4yz1NtSY
PnZQN+OTJlHNuJSyC3oY7gpu47Tw+ifM8G1F35l7UyXTYldqvFhYjLFQTpuo+K1e
8zyr8m3bGkAUee4IgEhPV4saWwFTYWDdHQ1DTaLaGltFHOvb/P0OfJNRBKSvPNZW
cUEKGflMW3L5FzFWWt1g6g9ocXvXajpuaKKVjG/V8dhuS88ja/R3xGeaW2vVbLCq
aZCk57GLecrzCJQhQRvgv0he0FDW9HoS1XC6BD3dBAtx5WaSQa8dSrRu2WAOKVFl
t1Hk9cu+SC/tXyI8rPs2IVRZh5WFPjfbG3sxGuajU+Wqq8XUTHJr3ptkYjOZUnLp
vpNn099tkIzgNHsgAfnIDVlVTyDkCS1g6hlKPX/VvGHbOeqUiw3FHtqltpZK7SAG
GxM3fI3kZkrcF+gVzg6Txwf0KmELzylLXwn+5Zry1NWxgo0sXXihysoozS3JynVX
sAjYGRJZeuhYcW1wmwQjt/YcqKVamHCLjHLFl3DcFfWHG4d3jIyUvAwbomopTODc
z3O1rXWiLkQaQXKTXfX2i1bulrYt5BMQHR7/GRYmXe2hK2CJTgbdwQLoowfHC4bz
OmUPRdV+15/PuJ6g3PJJj2RBulM7F35zZWs81U170uGdvrlpLijL5Kd3uCmL/70w
gcVb08aKRVr/J94wpMb+GVyIi7wE/kdasgPZrYZAP7PAUTLVD/IV9rF2zSoq8ovu
ws1LLpL89ayCev/rUMNAxnk+sMH58+Afi3hqHmhhCazk6n3eQqT4pEeFgX8bM8hk
ucWwaOq591u1yS3ABUddcgapBpK1LkUZMFYXVwTJ1WMXGRKbf7Wd2rc9IfuGD5qA
xbriUNmCb9AA551QQNqxIMGPrSiBsvhXYXNFzqBt6VYzTu8IfsGIMlPNrh+JRz7N
2dbtsS7P0yn6UyiXiypV2+/DqSzyARZERYr7vxJUStspNNBWOc0V2F39t5sNnYm5
00UKXObOqECRE3ll2vIXhJLXniCHw8Bv+rkGjRPwUqnN1Md1Sou7OXBchTIOPMvf
rKcP32FM8I1xuvSnb2Qcd+KAMHvdNkEVTGkI1Gb/ZqtwausNxn/e1318W51ZUBTE
qEw47UPPyDJeAOX4jsOxsLyYWD7NnEof2cgCgWOY4rKxEDxwMXMPrHis/q350B+V
Tm19yyRp3EIDf4yXYbe6JLFbjt4kn3ChVQMhXTtcCnL2piGOa52q+sNATigXwI9E
rar049GJKznRPnu36SBqdUmuMCJWOPwsYZo4CiwMa4b7tqEDSvor/Yp+HUZzfeMD
JTBIZrjwwtZUnxWsZg4zus+RAoareu3x35pfqjGZMH7omMCjJV50k+BICyZBO7Gg
Bc5I/LtqAVavgixKI3+zFRHBAA1XyCy2m8vgjqOgWdIjbFcsiTWSblXPCDE08EE4
xTJwPhTqky8uHtGCQvt8x45BvbwwSNJwLLkYLKeUtJrJc5AtWcF1LbZlRn9wVag2
CAvVunhAMwRcjSKRey9extcJva95JFI+TTqrTcD8HuNPN0n0yDfrQhXYZIiN06Wz
CPSg35O/2OHC+NjUTtqTeaQNwTk1gWU1lGhqEDbUiKLiyfqZA3OuiPGfC5MPSG0J
qF/fGsnldMSI+PaDlfICA+ksN+OL0N1fKSdLmzuEzvxWFAen6BTLYb3lCNhXmU34
siCpOJ4v0pGiyPCHVXE0t4hwbIPiAudNfv7d6+W4+RmTfE53QEt8hvjcUQaU2KIv
++isxfuqIV6GK1L5n4H9xxPep5nuqByQqfpLplMA1iqa5f5bb0Ee6GQ3BkvbDKXJ
Z//o617naZCQUBseDOC8PwNbgZ/5NLnOv3gAYnPqxRU9B86oUJxbbb++97yxvPsp
Jaq//GpT3KxfbdDRAY0HwpudqBNYBTqMr11JKkaFaj8+NqdHRJRx8QfiZJiO2KPN
Yn5kr5yEYYxnVeS6RHBLQ3sEl4T4n9Gnra0tQcPxvSIXTv7cGbVGnQfR3yuesl98
hTVj2Vu1CU87jU55zmmNcjpt3NZQ8gM+jX0kRZqVrhs1/Buj+RvgdNdGOT68Kzsx
iXuU3ZguEf7agb0KK1/0wpYcE02h5erL4gf6dZ8y9l/EgdSZ01qOozGuAmogaUMn
bJmjc8cWbHfBl+up0F0++hsznnboMOehsTQZltuMc09V8zUFQswmEkYI+kyLu9ei
WF0nK+pnT8Uc4/lfix+vZeRGtSGH8ry+MbQDXvmiF5foc5YYZ7dN1OSjgOz1Ixrg
1feuHfYsIrvjkjeenZtQOmZAtomE3HieGCva1Fcr2DBnwove5p0LuK1GJTprneMM
aiiJ+RncrRXR/kX9ThX2AtDglCQo7Hl8Ow0XSEp4yuuHJV23cb/HKrcQ/KKdiYVF
okG85SSDbpRipRVDy7TKkzG5buNnWZ+OCKbV771WvNNy/XGPuKyti4XKBAU7pCvT
NuKDBNKKcyiIIkcyaBbiwCn73E/W79zhzVsUzYv9E07Bnhp7GTC9btrVRYJ4+dLX
sIJriy6k5w5HXowALK9XZqoz2FJSXAKYUck7w1RQf9nq4lB7iSZ9S1PP3mA4OIxe
vZ7x5qZwwegWQLtHdlboRvJErVrmL89zkxSR3dwO0x64leKin0iC3LlqMxu3SSUK
y/lcUjt6/kBw2QIiORnSyuUmdxeO8BTLVQZPh6aQ6XqW2cSjWbXU5md880ReigDA
FKakWObJdHEUkzzkVquT+pbbCtEBI7iV4Vg79EC4mW1VCyFnVGqSw+JMv5DjX/t0
ZCeSrKpw+182Xj95JoDPZOAnXYMcdkvPt59wE08ep1bpFdWjq+DlZ+XqbvpGcbGI
hlBZhkBBLtH7sHU8+MQ/ZGGQOpGSo2j2b4R1APMS1gatulGj2Q5pOGZDsKXEkw8D
MUz7maWkAEDoaANLJAJStCoFK7LEeDEusE18rtZWUnIeBEmYff8tGweYDdxPyXkm
v3gXDAiF1NIL/Prsh6NJGiQ+BDARssgIm9b+p4yddMdNALP8epV2HRWGE8WktN+s
eHUMAZiTyVqC4RdxeezpW/O7PS02cf+7NXhDC2nxRZWokiPV614SGcx5X6eKjrbk
4sbeqR/39UWRPH5sB3XKFBV6pCblIsA8Sc2qBskYJP8frHcsfFJY/m+vLMQmeQqx
yO8R1PXvKhCq7XvI63K9/WOU1vPRWwfdXans2i42oYfBrBbtrYnmyVwDiwk2nVLi
NRuNUDzCX9J0xZ86KqphdEHaWW5OUoF4ynnOSfZnyY0Wsh3++ruCwqUAziWOlFON
HdcW05k6zxFF4fzf0U/8Hlsl121CngscmtKJAgCvf28fupw8+C03HeDdgNSCZ2+d
AsQkIUH/AnNW4BMKShuiRg5qMVDDr5tbISCfLCM6SbbWZeshTnZ7TQEzRl2OtYDu
rr5A2pKmH2CsCoPM9m606bTMnJVVgmheqrjtPU071/43T3EZS4D/oIMhvP2GLHob
WD82xYjf0wsDQpzIXDX14+FXUtYo5Vj9KlC6UCxTRWpVfRwA6mn73waa7O0wrMal
6elL5OuIsh4lQJAtr/ams7nRbffEmVLL/oP3WKYQqfcqqgsfviNKsdh2CRCDxc2i
kCB5Pch6Y8G7XwEFVY57E+N2YgKeEqF/55Ot5h78KB9G1EPU5IZAUn7EnMyXApzs
HVPX1/V2zMF4lFpDIxWkEm2KZ5+Qjde/vxH22vN/mpBAyiSfVELMSD11PXIiauPV
68hG2x/cDqnrobrie7u/Wb++Il1lUv+yUkGwdX6o2yl2jJEh6kKH5pZrO3rrB9Vw
BMQCDkE5MeQD78ORtGcblNiJTjYTfPJmlOP2/EGKgoD0eXrhvmiYYfq/8Qs7MTV2
ZffEb0colpSp1tPEOiC7tKiUwAANSA8rOUI7lKFMlUpAIg49L25uiiwliBylvu2r
3ZvEtKiOqW0m4IJDu8o6NWGLLQ5qcrcrxxEBZoBUI8vv/SVnxpmdVtdlgRAAZDkr
HELjsaWUSMDAczTdjzorMaPPyzOA1aePMuxOFvXrGc2VelYIKKL3AY4iQSI5NkEI
Y2jCSvTaxEKsIAJXr4BJZ/myHZfGUZEIVITzFSkiLLX31trBqliekT0qhgUcPykc
poLrI/Unz4Y3RUXZSJ26KYQtNC8mGGnwwkj8uRgTzJTKZ9i9xEKLqemCFrg6wijV
BMnATGUOF4DE7XEEh5iM0yTzSV37L0BOk9mnQzlEaN6PmZg0sWq1ZMg0Z6XJor8z
MJJfbdpnz5B/4cJlbbzVMcJwEJRyXeCwL2QTwZGvC4RLaWNXCNDKkwx+sjJWvhV+
lQdVS0hu4lMaDa6s01j9Daso5bRuGLzP8OIUpdWCWn3jmCN7cpU9R346o/zPLyw/
IPYPvbMig4/eHoymbmpZzBhaLeE3gQIhxVjl0PyjkALGWdy44n/l0URSXFclL9t6
SZi1GO4ffB44hS9bzH9otoqovbgWPf6k3WJkzN0tAKaIPJ5hxtGizxB4rFhYXEVP
7ntMRL7u1aMVfwZpkelHNUu/hC6LFqHN5UA0tlqlfWZ1Sn6elDScsTzYrnsMF1hk
hRRs3h/JHbeBLoSfcayhdbb+VWqX4lpJ2Q70QYXYCDHyX7Q2bxoIi+hEVhoVH9pC
uSeCD9Z3/8Kr3LiAVyCc7vsPOL75p+xYja0kk2vApSPO5KzVfbpAXbkGXz9YO9rF
3EsZwo9hoztjGyyB0q2btuVySv/nUvT4fEaUCcp3Ig7hfOg2VoWIS7Y+WB52ILhm
XX7LuFzptsrZ8I+L27H6Wl19P0KGdcVD1GQmgeEUCxU0iM0Gqd40gQh9Hv3rfh0j
L4/tXtvFhf78NGUNk9RBruQgBaWqlvDdc2szg2xsI16HBwgEIFmRh0+vwdItNiMW
behmjpv9Qae5K/lbECuPe0qmq221agxWCPh9aVHOj1R5vLayYctRUqFl6in0JWHs
mWYh17WCNRnWe8LxixT9Yt1816srrWtfJN/EwG3tbnK5orvCr3xqw0lia1tXGyM+
HoRKVXwFjXtYhe3Q28tYbFJ1f90h6Q0A/+iCRhblDomVlh9k3Qc8BVKz3bHYoNuv
/1QQ6nCgge9saf4i6qVgGd64EBjHZsPVnMmsMSlhryl748UdFOLZvxSY6PKGPBpE
siA7uLjpvEI2f3s4MxetWk3YsYeSnk/3YgQRkzYLRJQwgms/fXV3hwlhxjdI1oo1
Ljhr+mcIICT+5+XXPDRkSOuBreTCZApIr95eFnJ28Gi6nuF3WeCeSJKWrHLXbHXY
uVpDZeIcphPXGLCo5/DQShCVSeJOGcsXxV7q6fWXOikLZI83+VoCa4C22iMJoZPB
Vvj47YPc/aDU9y6AvNrFsS70NN7Z8tDwRV1uPolUrtqWw6L5jXJV5YFymTPOW1oG
CXOb3zmSkQXQY3AVtdLhUR2BAkGES7ZNZ9ZuZb2TH1OTrSNM0lcrmO6AD5sNpxAp
NEnAB3TcKU+yN4776XbWccksjuWFB9dptQ8mOw0EealPe2+R/uH1vkowmm/fjHuB
aGnuqf1Ko/qGb570ISu0r+euX3KXTt1oRqqtEIXSeAIIZi9wNvoEdhqUZRd+truo
7WrQ/W0Jsra6B4ROg/W5l2KOyDZ54Rx6HlyxwwTL8AULmJn0cKfAd0Sx+xDGzZfG
XzOCjo1CuWI5h4Z09CjlmZEHfzUs5Kfj6qbEKfi/IbYXQiFNLR4FjSgSAWBulAe1
XYeySQC/vjpbhqp5ZYbkYJN2udCelxY0TLHpjAKT8tjWhwfJB39ycZe6P+FgF2eh
hhWlmPwuc8BivQuiRsK80nCtRRYY+sYHWL897Y5/DB4kqdt4UqrQ/XMZj2K7zHfW
A03SaXr4JRWPQsAPhXaV61kEdZ3jMc6j4aOSc7FId7IrzHU54Q/VbO1LGGY/BMVz
yb7AA3RD3dCGD4ho13L0DC9NsNfKBR/WFhESVsS8482h5dB3Pnx6VpmpW/MzDZH4
hhMedszX0juidYsGYOqjRKPbKTjPU9hQkdR/57g4KpxHzvCTCLhUzK+nOteMACj0
N0AZqNw7G4EUfJNhpucPpSHAIzq5vKpIwmXPyiZzttnuIUxieF7pCHc/dzbKbgHf
mMmfVs8R7CcvrT8CefMZ8xUYfdzw73put9Go+umwBLfozDUh+HtCrQvNGGmFNuxv
HB45LHakZSgdDkSKbDZQ6bM/68S768/KbqBeNXIyN14wCyS0omW3SBrCAcrX2v6K
UEXUma5KXRf04FFSNCCIpKsGz25lDzrilTsQLg0DutemEA3VL5me5GzYUgBCzOq2
q3fd7KmIZcrfXUJtQnF7TK4DRQNwNR7fUkhgofw16p+6p/eQfQYCRAZOovLpFsrx
bakY/qSLbhGft9mpGb/BjNzdQ2jNJPAkZcAh1/IjXt6AQH+azZdguW19h/pCH3v5
zYMV4Q6ieTjrTXx3Pnm8tWtpnGXZR7sN+TwxxEvDS9FkohF4PACCd5CF3PAzzRpm
VIoZ0Vwm4FWXf6wFIe8p/joYdKi/NPwuwYgkU+6Wl0S/Napr43I4UIBJpQeQU8fa
1bR6k9kx31ZuoYB8G1r+AZqH3p5djLNn57FEq+X2zinT/NE3CsqKuUMf9qJudSmp
tk3xcCTX4+xzdnE9pm6uNjftxKgm3AuBNXVFwjWzWWUoD5F2cHOfsaws1NHGW4S1
Ff8YWUo6k3Iaqnxnwxfe0uf4i620WtVd8nJkwdvQHBIzv98Ocv92ec9n4saxT/8m
YLHNsBrIGgn+RxKcAH87IAEoT6qY+w5fdl3zrzK6+aZU8dDYaTVKINM5YzFpOS9A
JK/GfS17/33ACNaPH6hC71cQISIK0bHZnY6yXW2rUgwgxxn9B+lKmQbYnRge8tt3
3EnT95avKtw+Rvlefu6jjCPMLnXmn60XHNgVWx8JWdmX/ljmECQ/fSHe6wta2MpY
TdR5SHnomko1NZcI4zpnW2yGdsBLWvkg7cF2gzfJlT0xBmBDAQRjveOeTwDuOGxD
FX4dcjJEbQLi1Z5ALDNZkIujfi1G5lRACuvtT/cNQivhwZUjFP6NA220fuIbVZML
dQ4BW35AfPbSx9Q0DvffJ+KXHUDZuU031vmgkJcdhaOuHN5VZY6mPPUIRudCYfTV
2bbBCleADITEy3x8avUDbHDm1ZWRPZ70q9Nkwrn3KSCMF3tN1RAf/Ww6vpqgKn9J
WdGjHfuRWl35gejUXJWAwW4xPIBOSvWgvM19XV6BtyBneLzZBqSrcm7T4/+tx1OM
c8GUTEQFuH+yqeWzTqvbZlMtRM1NnzZtGmbKUhipwA5LbPvmOO4rO0tTCqQbsfhR
wpNv35wO2MN8yKVrvGskXCA0x4NQV/q8vcrQWI3Fufi4YjM0bWD8+esN2S3HPFo3
pQ30yS86EfpHAHVWN7IfIGfX9G9VdTc8EU5Dzuj85CBvWVDHbGIbAPcOfu+iwHn+
w7N+XM6sCeRHNGoYcneszcbwMn9wUntyVDlUgHveWW5zCK7goX8Cl3WPR7Vz10z0
V03Dcr3FbYiDajcP1lC10Qimz0CgDxfivmELtURQEzLTST4ExDVigUODQynr9to9
/59Nm7KoiKbrsSJCqlOYmpd8bHn9L9oWiqXVx0pMzwqY09yWHEgGzL28MORFXxzx
i2XhWROcOlfpcXpR7pENOg7mDAzx7UdQ76HZC4754R5bLBaIW1jKqIPinO8o5Pr/
lVyaEbiKeePhf3M6RGsNVr67iwz36jj1bvMB23aU2JfaQkw1Ek5UiDKod7+Czf5L
C5G9w2tgs2/8FSnuS1hLLHCZBhd2vlcRflA+UIVJo4yzHiNQC+hGNmCjajtmcdS6
Rn7sGESPeqEZrUtHIM2rJF1y8L4gdUTcilh8i1BC/FRlvDyFToPVUZD2wAbhhAh0
3UkMSV+7cqUEUqc5G86bOqHk+bl0MZuLqXmT0DosT46xzcazYdeOE6kdOmqqkumY
wseBW6svNe/ChvV4nrJzbLdorhuGOrkZyBal7OAIfUHniVtWBf52z8FNFjEnUPG4
llMRe4HxZTeWAu9C7A/YNDV6r8edLgTYz29DypkiEFOvIMbHCS7NrS2FSuVmjjHZ
pv5mqS8uJDwUVGUlCbnuf/p7ZcCtWICcOnRuSnt3H8YDrT7CN2+tZVkZj9854AHE
mtxc1NCDs7J+Hiot29UlCOqMpcxIhRQSvhhE37/exxbJ7iNgJAlsbWU1vcoaSxKv
8sLn6rE/9bngKm5vVehTlHw5Um9gstrLVtZwzf+QqB/xI6LwujeD9I88opVXBOaf
1naRSFFOdSDUvP1HgaW0ZKKVcBDmrrTGuQp7YJOcIpfT0njiWRgFQ4JAxbEmGDEO
YyncwY4diJ47VWYw3b94H5dYXLImyB2X+HiN8vjJrzyL+KXbmyKA3A9HpAeizgJZ
px6NiihC5MI5Uoy7jy8KhOO9hGSNDQ1MIYXYbvWUyQ/Sd7JNezyVHjpONC8DxNbr
cCoYj0LT2k0W+J0Ul2wP25ReMS80FYaQnwPXgnb0Y0goDrglaEmk1kWz/6Ymlbrv
lB+9qK1wNOp0etXrvIQdGvrtN21EUX2iID2J6DwUTMNpUlGMX3UCYT9gyrS1ihuD
0Kl+PRCY7ZgCmDviqvDLXBprwChdZTiRkUCnxQi+jW7VLpFXRuAn+uwl2GDAybrB
wXfZ95E/3tK1hL3EvPwIzwRWMJ5QmZhsTHfr0utja5ICQX+v4Cn4IDwC9XChulY8
8CVO+zbgFv33bFz4l5Viy8d7wmU9gd7RPG3PubX6Ydmt2uQoj3TQZSsKnF0BQAyJ
yD2kM5hlbZcC0nJzWIj7KD7zexaIeqn+CvUGgje0UQZR4X2oytaezatStqpQMOkO
NHB1ZdapzshVqXgcqPnXOURqQbI2wI4PVqLh/Z2GFKTqiN8xPkMnEzqCLmtyK/PL
Rk8yorF37/JczNBFJ29QXUZjMTlEvF9XSj3fVu8XQHGNPNzph5E3Yudwt3YbO8Al
xLUWucO/yqziyHm8IgRffRL3rwiqH9OYUoKKxytc4u9wdDigHz+wOC+XYTJ/2JvR
LKsvv+vt8Jz4dGxwDUPk3NLwDxR6scUDtXUQLBPpRGBAU2wBkC6FzR+ZWQdSZnIR
oAmKysT0W3kh8p14HbR2HzOuKzCf5Ru+nl39jkbcD5OIPDvaOYgxrRyWNobmWayj
8DJ5y6C0QzXTbNYTgePoETBbxs9W29d7hjHLb3eSNxpM5tnHpbBTw00ODVDPARvT
m3dqElmEkZ2VQ3v/DdSRdCmdyKgqbw6Rf256erPrnJu53KUNPfVCU/C9VoLK3V2g
1926KxfAhzZKd1kkSBR4dRm3+kK+3W47PEcfGEwZCCYY0Kn7y/KHQW86rWLwv155
cwyb1pBm8YUPbXSY95olRkmPhwdkUfnexlKapYiq0HUh2iHp1V/GuxKU2JNp/M+T
zTuw8ljWf4cVQ8vfay+ubT3mONCsldyHfV3Ncy39qybn7baSurbvKiIavcNhE7c7
KjTZGWcIH3geC9zbkjUI0c1QI5ZWvGm+n2FCMClRQDHH8E2vbbpsQT3hLtdKe+CS
b4S+iA3wW9XWhSbjZvNNXxBLDX6Saw1mxECBfXrj/3TpTJdG6BCn4FAL6EIrVemd
deKZEIgRLjbDd3CUGu+Mnb2IUMM/i5+khdHqoWvdgQh4TzAsYpfE56Iq1/oD6nRt
WGvlyoMGIHwP1Ye2KHs3F2D+ubeCWLxllyu+F4hFckqxEiI7wROABf6xuLqJd9ep
ov05A2nHIdV5YrLx2GQeW136nN0p/r7L0gK7hHYaOc5k06BaOwVKhY0gIn7ClWdU
ojAxAmuKWdB/KHp4VVr1ct3PY/kENwjdFl9Rk9KYtfpSsT5AQ2wH+Q6KWzBd7w3s
1Vx7lIB3Pp0/CFnCUvDiv+rd/pfFUVC4Uo05l8shwG3ZylYrPxfXWYG+DUv2MbP0
nm6VBzgqXE9cCDs5i7W2ZmW7C6Dn+SOoWSIEUpWCI5vhPl8AamzgO+2XDqL3fcqr
jwLZj80RcNXGiARRenKCUCorJ0CzE+tUoptBl2QHc7+jJ2BAlfSiDjlJTPtFkdpk
vlrsnspulf5IKedhOGA5XJkM8KMHezV+Y5WL5zNm9Oyw7dO5TPdGg7ZY3TAuTqjQ
BRgwTLguNng9VEx6hKyPSKWNKQUq+7iqs2KH5dY5RbrKyJVvGqDRJr9vcig2FZZT
lr3a9ee7Mb0htC9SJQj66tIHVreB9BdGp2djNQKe1AFNyxKVxW4VrT+CHS/7w8z6
1IEIxNRbW2m17mVO8ZKu1r4bPjHLzr7RA68V+NGxhBbzcberjJXBAHFBAm2XVQpd
RCjkKDZdIjhfil92PdPVKDcB8E4UC5xHtPQb6V1HF0/mQh1fl1mrxVE3QVWJbit/
oLWzHFra+ELJZIhYC1i/tf2/oRiGNUPayQFRzJ0I/+s+wp98U+gWJgzMUqrmz2hd
3tq0Som9zOOWnTamws5UBwIZGU8ln4o8nLr+J+PRNXFHuh8Ni4mNVrjJQOi8bJPx
ZPWLCzbRbzgN4D2IJfEtwaaiuMCuwj5tHlhoO7H/8fgXtfQDjJZy0jzJXRK0OcWN
Y5Ym1mO0CTFN27Bag0bviDrHmPKVx/hEajWnlgkkAFLn3XHlz7Og5ALNfBXYl5kW
weFtf2bngbxycezchyGmRg==
`protect end_protected
