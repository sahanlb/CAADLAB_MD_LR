localparam [NNN1D-1:0][NNN1D-1:0][NNN1D-1:0][BMEMD-1:0][31:0] ROMVAL = {
  32'h3f5a3fd8 /* (15, 15, 15) */,
  32'h3e93e191 /* (11, 15, 15) */,
  32'h3ea4f994 /* (7, 15, 15) */,
  32'h3eaf2a10 /* (3, 15, 15) */,
  32'h3e93e191 /* (15, 11, 15) */,
  32'h3eeeb6df /* (11, 11, 15) */,
  32'h3f2b075a /* (7, 11, 15) */,
  32'h3ea7dbb1 /* (3, 11, 15) */,
  32'h3ea4f994 /* (15, 7, 15) */,
  32'h3f2b075a /* (11, 7, 15) */,
  32'h3f88838c /* (7, 7, 15) */,
  32'h3ed1d4cb /* (3, 7, 15) */,
  32'h3eaf2a10 /* (15, 3, 15) */,
  32'h3ea7dbb1 /* (11, 3, 15) */,
  32'h3ed1d4cb /* (7, 3, 15) */,
  32'h3e953797 /* (3, 3, 15) */,
  32'h3e93e191 /* (15, 15, 11) */,
  32'h3eeeb6df /* (11, 15, 11) */,
  32'h3f2b075a /* (7, 15, 11) */,
  32'h3ea7dbb1 /* (3, 15, 11) */,
  32'h3eeeb6df /* (15, 11, 11) */,
  32'h3f77795a /* (11, 11, 11) */,
  32'h3fc5882d /* (7, 11, 11) */,
  32'h3f17cf64 /* (3, 11, 11) */,
  32'h3f2b075a /* (15, 7, 11) */,
  32'h3fc5882d /* (11, 7, 11) */,
  32'h40278361 /* (7, 7, 11) */,
  32'h3f6365d6 /* (3, 7, 11) */,
  32'h3ea7dbb1 /* (15, 3, 11) */,
  32'h3f17cf64 /* (11, 3, 11) */,
  32'h3f6365d6 /* (7, 3, 11) */,
  32'h3ec9097c /* (3, 3, 11) */,
  32'h3ea4f994 /* (15, 15, 7) */,
  32'h3f2b075a /* (11, 15, 7) */,
  32'h3f88838c /* (7, 15, 7) */,
  32'h3ed1d4cb /* (3, 15, 7) */,
  32'h3f2b075a /* (15, 11, 7) */,
  32'h3fc5882d /* (11, 11, 7) */,
  32'h40278361 /* (7, 11, 7) */,
  32'h3f6365d6 /* (3, 11, 7) */,
  32'h3f88838c /* (15, 7, 7) */,
  32'h40278361 /* (11, 7, 7) */,
  32'h4093adcc /* (7, 7, 7) */,
  32'h3fb9d98f /* (3, 7, 7) */,
  32'h3ed1d4cb /* (15, 3, 7) */,
  32'h3f6365d6 /* (11, 3, 7) */,
  32'h3fb9d98f /* (7, 3, 7) */,
  32'h3f07f0f8 /* (3, 3, 7) */,
  32'h3eaf2a10 /* (15, 15, 3) */,
  32'h3ea7dbb1 /* (11, 15, 3) */,
  32'h3ed1d4cb /* (7, 15, 3) */,
  32'h3e953797 /* (3, 15, 3) */,
  32'h3ea7dbb1 /* (15, 11, 3) */,
  32'h3f17cf64 /* (11, 11, 3) */,
  32'h3f6365d6 /* (7, 11, 3) */,
  32'h3ec9097c /* (3, 11, 3) */,
  32'h3ed1d4cb /* (15, 7, 3) */,
  32'h3f6365d6 /* (11, 7, 3) */,
  32'h3fb9d98f /* (7, 7, 3) */,
  32'h3f07f0f8 /* (3, 7, 3) */,
  32'h3e953797 /* (15, 3, 3) */,
  32'h3ec9097c /* (11, 3, 3) */,
  32'h3f07f0f8 /* (7, 3, 3) */,
  32'h3e9a814a /* (3, 3, 3) */,
  32'h3efc66bd /* (14, 15, 15) */,
  32'h3e9f454b /* (10, 15, 15) */,
  32'h3e9f454b /* (6, 15, 15) */,
  32'h3efc66bd /* (2, 15, 15) */,
  32'h3e99eb68 /* (14, 11, 15) */,
  32'h3f14d2ae /* (10, 11, 15) */,
  32'h3f14d2ae /* (6, 11, 15) */,
  32'h3e99eb68 /* (2, 11, 15) */,
  32'h3eb430e1 /* (14, 7, 15) */,
  32'h3f62162b /* (10, 7, 15) */,
  32'h3f62162b /* (6, 7, 15) */,
  32'h3eb430e1 /* (2, 7, 15) */,
  32'h3e9f2a5d /* (14, 3, 15) */,
  32'h3ec1987e /* (10, 3, 15) */,
  32'h3ec1987e /* (6, 3, 15) */,
  32'h3e9f2a5d /* (2, 3, 15) */,
  32'h3e99eb68 /* (14, 15, 11) */,
  32'h3f14d2ae /* (10, 15, 11) */,
  32'h3f14d2ae /* (6, 15, 11) */,
  32'h3e99eb68 /* (2, 15, 11) */,
  32'h3f025da2 /* (14, 11, 11) */,
  32'h3fa39217 /* (10, 11, 11) */,
  32'h3fa39217 /* (6, 11, 11) */,
  32'h3f025da2 /* (2, 11, 11) */,
  32'h3f3e2f24 /* (14, 7, 11) */,
  32'h4006bd24 /* (10, 7, 11) */,
  32'h4006bd24 /* (6, 7, 11) */,
  32'h3f3e2f24 /* (2, 7, 11) */,
  32'h3eb2cc97 /* (14, 3, 11) */,
  32'h3f41f419 /* (10, 3, 11) */,
  32'h3f41f419 /* (6, 3, 11) */,
  32'h3eb2cc97 /* (2, 3, 11) */,
  32'h3eb430e1 /* (14, 15, 7) */,
  32'h3f62162b /* (10, 15, 7) */,
  32'h3f62162b /* (6, 15, 7) */,
  32'h3eb430e1 /* (2, 15, 7) */,
  32'h3f3e2f24 /* (14, 11, 7) */,
  32'h4006bd24 /* (10, 11, 7) */,
  32'h4006bd24 /* (6, 11, 7) */,
  32'h3f3e2f24 /* (2, 11, 7) */,
  32'h3f993b79 /* (14, 7, 7) */,
  32'h406912bc /* (10, 7, 7) */,
  32'h406912bc /* (6, 7, 7) */,
  32'h3f993b79 /* (2, 7, 7) */,
  32'h3ee6ec8a /* (14, 3, 7) */,
  32'h3f982d5a /* (10, 3, 7) */,
  32'h3f982d5a /* (6, 3, 7) */,
  32'h3ee6ec8a /* (2, 3, 7) */,
  32'h3e9f2a5d /* (14, 15, 3) */,
  32'h3ec1987e /* (10, 15, 3) */,
  32'h3ec1987e /* (6, 15, 3) */,
  32'h3e9f2a5d /* (2, 15, 3) */,
  32'h3eb2cc97 /* (14, 11, 3) */,
  32'h3f41f419 /* (10, 11, 3) */,
  32'h3f41f419 /* (6, 11, 3) */,
  32'h3eb2cc97 /* (2, 11, 3) */,
  32'h3ee6ec8a /* (14, 7, 3) */,
  32'h3f982d5a /* (10, 7, 3) */,
  32'h3f982d5a /* (6, 7, 3) */,
  32'h3ee6ec8a /* (2, 7, 3) */,
  32'h3e9508f6 /* (14, 3, 3) */,
  32'h3ef2a853 /* (10, 3, 3) */,
  32'h3ef2a853 /* (6, 3, 3) */,
  32'h3e9508f6 /* (2, 3, 3) */,
  32'h3eaf2a10 /* (13, 15, 15) */,
  32'h3ea4f994 /* (9, 15, 15) */,
  32'h3e93e191 /* (5, 15, 15) */,
  32'h3f5a3fd8 /* (1, 15, 15) */,
  32'h3ea7dbb1 /* (13, 11, 15) */,
  32'h3f2b075a /* (9, 11, 15) */,
  32'h3eeeb6df /* (5, 11, 15) */,
  32'h3e93e191 /* (1, 11, 15) */,
  32'h3ed1d4cb /* (13, 7, 15) */,
  32'h3f88838c /* (9, 7, 15) */,
  32'h3f2b075a /* (5, 7, 15) */,
  32'h3ea4f994 /* (1, 7, 15) */,
  32'h3e953797 /* (13, 3, 15) */,
  32'h3ed1d4cb /* (9, 3, 15) */,
  32'h3ea7dbb1 /* (5, 3, 15) */,
  32'h3eaf2a10 /* (1, 3, 15) */,
  32'h3ea7dbb1 /* (13, 15, 11) */,
  32'h3f2b075a /* (9, 15, 11) */,
  32'h3eeeb6df /* (5, 15, 11) */,
  32'h3e93e191 /* (1, 15, 11) */,
  32'h3f17cf64 /* (13, 11, 11) */,
  32'h3fc5882d /* (9, 11, 11) */,
  32'h3f77795a /* (5, 11, 11) */,
  32'h3eeeb6df /* (1, 11, 11) */,
  32'h3f6365d6 /* (13, 7, 11) */,
  32'h40278361 /* (9, 7, 11) */,
  32'h3fc5882d /* (5, 7, 11) */,
  32'h3f2b075a /* (1, 7, 11) */,
  32'h3ec9097c /* (13, 3, 11) */,
  32'h3f6365d6 /* (9, 3, 11) */,
  32'h3f17cf64 /* (5, 3, 11) */,
  32'h3ea7dbb1 /* (1, 3, 11) */,
  32'h3ed1d4cb /* (13, 15, 7) */,
  32'h3f88838c /* (9, 15, 7) */,
  32'h3f2b075a /* (5, 15, 7) */,
  32'h3ea4f994 /* (1, 15, 7) */,
  32'h3f6365d6 /* (13, 11, 7) */,
  32'h40278361 /* (9, 11, 7) */,
  32'h3fc5882d /* (5, 11, 7) */,
  32'h3f2b075a /* (1, 11, 7) */,
  32'h3fb9d98f /* (13, 7, 7) */,
  32'h4093adcc /* (9, 7, 7) */,
  32'h40278361 /* (5, 7, 7) */,
  32'h3f88838c /* (1, 7, 7) */,
  32'h3f07f0f8 /* (13, 3, 7) */,
  32'h3fb9d98f /* (9, 3, 7) */,
  32'h3f6365d6 /* (5, 3, 7) */,
  32'h3ed1d4cb /* (1, 3, 7) */,
  32'h3e953797 /* (13, 15, 3) */,
  32'h3ed1d4cb /* (9, 15, 3) */,
  32'h3ea7dbb1 /* (5, 15, 3) */,
  32'h3eaf2a10 /* (1, 15, 3) */,
  32'h3ec9097c /* (13, 11, 3) */,
  32'h3f6365d6 /* (9, 11, 3) */,
  32'h3f17cf64 /* (5, 11, 3) */,
  32'h3ea7dbb1 /* (1, 11, 3) */,
  32'h3f07f0f8 /* (13, 7, 3) */,
  32'h3fb9d98f /* (9, 7, 3) */,
  32'h3f6365d6 /* (5, 7, 3) */,
  32'h3ed1d4cb /* (1, 7, 3) */,
  32'h3e9a814a /* (13, 3, 3) */,
  32'h3f07f0f8 /* (9, 3, 3) */,
  32'h3ec9097c /* (5, 3, 3) */,
  32'h3e953797 /* (1, 3, 3) */,
  32'h3e94e1d9 /* (12, 15, 15) */,
  32'h3e8d5b73 /* (8, 15, 15) */,
  32'h3e94e1d9 /* (4, 15, 15) */,
  32'h3f9befb2 /* (0, 15, 15) */,
  32'h3ec28d9a /* (12, 11, 15) */,
  32'h3f1e09be /* (8, 11, 15) */,
  32'h3ec28d9a /* (4, 11, 15) */,
  32'h3e924c17 /* (0, 11, 15) */,
  32'h3f0271c0 /* (12, 7, 15) */,
  32'h3f8374c7 /* (8, 7, 15) */,
  32'h3f0271c0 /* (4, 7, 15) */,
  32'h3ea04e75 /* (0, 7, 15) */,
  32'h3e97a967 /* (12, 3, 15) */,
  32'h3eb9823a /* (8, 3, 15) */,
  32'h3e97a967 /* (4, 3, 15) */,
  32'h3eb78ea1 /* (0, 3, 15) */,
  32'h3ec28d9a /* (12, 15, 11) */,
  32'h3f1e09be /* (8, 15, 11) */,
  32'h3ec28d9a /* (4, 15, 11) */,
  32'h3e924c17 /* (0, 15, 11) */,
  32'h3f3cbfdf /* (12, 11, 11) */,
  32'h3fbe36ae /* (8, 11, 11) */,
  32'h3f3cbfdf /* (4, 11, 11) */,
  32'h3ee7f590 /* (0, 11, 11) */,
  32'h3f91d65e /* (12, 7, 11) */,
  32'h40258eba /* (8, 7, 11) */,
  32'h3f91d65e /* (4, 7, 11) */,
  32'h3f2521d3 /* (0, 7, 11) */,
  32'h3ef076ff /* (12, 3, 11) */,
  32'h3f558e61 /* (8, 3, 11) */,
  32'h3ef076ff /* (4, 3, 11) */,
  32'h3ea49cf9 /* (0, 3, 11) */,
  32'h3f0271c0 /* (12, 15, 7) */,
  32'h3f8374c7 /* (8, 15, 7) */,
  32'h3f0271c0 /* (4, 15, 7) */,
  32'h3ea04e75 /* (0, 15, 7) */,
  32'h3f91d65e /* (12, 11, 7) */,
  32'h40258eba /* (8, 11, 7) */,
  32'h3f91d65e /* (4, 11, 7) */,
  32'h3f2521d3 /* (0, 11, 7) */,
  32'h3ff29d82 /* (12, 7, 7) */,
  32'h4094977b /* (8, 7, 7) */,
  32'h3ff29d82 /* (4, 7, 7) */,
  32'h3f836079 /* (0, 7, 7) */,
  32'h3f2b2ff1 /* (12, 3, 7) */,
  32'h3fb4be0d /* (8, 3, 7) */,
  32'h3f2b2ff1 /* (4, 3, 7) */,
  32'h3ecb578e /* (0, 3, 7) */,
  32'h3e97a967 /* (12, 15, 3) */,
  32'h3eb9823a /* (8, 15, 3) */,
  32'h3e97a967 /* (4, 15, 3) */,
  32'h3eb78ea1 /* (0, 15, 3) */,
  32'h3ef076ff /* (12, 11, 3) */,
  32'h3f558e61 /* (8, 11, 3) */,
  32'h3ef076ff /* (4, 11, 3) */,
  32'h3ea49cf9 /* (0, 11, 3) */,
  32'h3f2b2ff1 /* (12, 7, 3) */,
  32'h3fb4be0d /* (8, 7, 3) */,
  32'h3f2b2ff1 /* (4, 7, 3) */,
  32'h3ecb578e /* (0, 7, 3) */,
  32'h3eaaa637 /* (12, 3, 3) */,
  32'h3ef65451 /* (8, 3, 3) */,
  32'h3eaaa637 /* (4, 3, 3) */,
  32'h3e960c85 /* (0, 3, 3) */,
  32'h3efc66bd /* (15, 14, 15) */,
  32'h3e99eb68 /* (11, 14, 15) */,
  32'h3eb430e1 /* (7, 14, 15) */,
  32'h3e9f2a5d /* (3, 14, 15) */,
  32'h3e9f454b /* (15, 10, 15) */,
  32'h3f14d2ae /* (11, 10, 15) */,
  32'h3f62162b /* (7, 10, 15) */,
  32'h3ec1987e /* (3, 10, 15) */,
  32'h3e9f454b /* (15, 6, 15) */,
  32'h3f14d2ae /* (11, 6, 15) */,
  32'h3f62162b /* (7, 6, 15) */,
  32'h3ec1987e /* (3, 6, 15) */,
  32'h3efc66bd /* (15, 2, 15) */,
  32'h3e99eb68 /* (11, 2, 15) */,
  32'h3eb430e1 /* (7, 2, 15) */,
  32'h3e9f2a5d /* (3, 2, 15) */,
  32'h3e99eb68 /* (15, 14, 11) */,
  32'h3f025da2 /* (11, 14, 11) */,
  32'h3f3e2f24 /* (7, 14, 11) */,
  32'h3eb2cc97 /* (3, 14, 11) */,
  32'h3f14d2ae /* (15, 10, 11) */,
  32'h3fa39217 /* (11, 10, 11) */,
  32'h4006bd24 /* (7, 10, 11) */,
  32'h3f41f419 /* (3, 10, 11) */,
  32'h3f14d2ae /* (15, 6, 11) */,
  32'h3fa39217 /* (11, 6, 11) */,
  32'h4006bd24 /* (7, 6, 11) */,
  32'h3f41f419 /* (3, 6, 11) */,
  32'h3e99eb68 /* (15, 2, 11) */,
  32'h3f025da2 /* (11, 2, 11) */,
  32'h3f3e2f24 /* (7, 2, 11) */,
  32'h3eb2cc97 /* (3, 2, 11) */,
  32'h3eb430e1 /* (15, 14, 7) */,
  32'h3f3e2f24 /* (11, 14, 7) */,
  32'h3f993b79 /* (7, 14, 7) */,
  32'h3ee6ec8a /* (3, 14, 7) */,
  32'h3f62162b /* (15, 10, 7) */,
  32'h4006bd24 /* (11, 10, 7) */,
  32'h406912bc /* (7, 10, 7) */,
  32'h3f982d5a /* (3, 10, 7) */,
  32'h3f62162b /* (15, 6, 7) */,
  32'h4006bd24 /* (11, 6, 7) */,
  32'h406912bc /* (7, 6, 7) */,
  32'h3f982d5a /* (3, 6, 7) */,
  32'h3eb430e1 /* (15, 2, 7) */,
  32'h3f3e2f24 /* (11, 2, 7) */,
  32'h3f993b79 /* (7, 2, 7) */,
  32'h3ee6ec8a /* (3, 2, 7) */,
  32'h3e9f2a5d /* (15, 14, 3) */,
  32'h3eb2cc97 /* (11, 14, 3) */,
  32'h3ee6ec8a /* (7, 14, 3) */,
  32'h3e9508f6 /* (3, 14, 3) */,
  32'h3ec1987e /* (15, 10, 3) */,
  32'h3f41f419 /* (11, 10, 3) */,
  32'h3f982d5a /* (7, 10, 3) */,
  32'h3ef2a853 /* (3, 10, 3) */,
  32'h3ec1987e /* (15, 6, 3) */,
  32'h3f41f419 /* (11, 6, 3) */,
  32'h3f982d5a /* (7, 6, 3) */,
  32'h3ef2a853 /* (3, 6, 3) */,
  32'h3e9f2a5d /* (15, 2, 3) */,
  32'h3eb2cc97 /* (11, 2, 3) */,
  32'h3ee6ec8a /* (7, 2, 3) */,
  32'h3e9508f6 /* (3, 2, 3) */,
  32'h3ec29928 /* (14, 14, 15) */,
  32'h3eaab74a /* (10, 14, 15) */,
  32'h3eaab74a /* (6, 14, 15) */,
  32'h3ec29928 /* (2, 14, 15) */,
  32'h3eaab74a /* (14, 10, 15) */,
  32'h3f3f980b /* (10, 10, 15) */,
  32'h3f3f980b /* (6, 10, 15) */,
  32'h3eaab74a /* (2, 10, 15) */,
  32'h3eaab74a /* (14, 6, 15) */,
  32'h3f3f980b /* (10, 6, 15) */,
  32'h3f3f980b /* (6, 6, 15) */,
  32'h3eaab74a /* (2, 6, 15) */,
  32'h3ec29928 /* (14, 2, 15) */,
  32'h3eaab74a /* (10, 2, 15) */,
  32'h3eaab74a /* (6, 2, 15) */,
  32'h3ec29928 /* (2, 2, 15) */,
  32'h3ea1d2a3 /* (14, 14, 11) */,
  32'h3f242ada /* (10, 14, 11) */,
  32'h3f242ada /* (6, 14, 11) */,
  32'h3ea1d2a3 /* (2, 14, 11) */,
  32'h3f242ada /* (14, 10, 11) */,
  32'h3fdbd2f0 /* (10, 10, 11) */,
  32'h3fdbd2f0 /* (6, 10, 11) */,
  32'h3f242ada /* (2, 10, 11) */,
  32'h3f242ada /* (14, 6, 11) */,
  32'h3fdbd2f0 /* (10, 6, 11) */,
  32'h3fdbd2f0 /* (6, 6, 11) */,
  32'h3f242ada /* (2, 6, 11) */,
  32'h3ea1d2a3 /* (14, 2, 11) */,
  32'h3f242ada /* (10, 2, 11) */,
  32'h3f242ada /* (6, 2, 11) */,
  32'h3ea1d2a3 /* (2, 2, 11) */,
  32'h3ec56b70 /* (14, 14, 7) */,
  32'h3f7ca6c7 /* (10, 14, 7) */,
  32'h3f7ca6c7 /* (6, 14, 7) */,
  32'h3ec56b70 /* (2, 14, 7) */,
  32'h3f7ca6c7 /* (14, 10, 7) */,
  32'h4039abaa /* (10, 10, 7) */,
  32'h4039abaa /* (6, 10, 7) */,
  32'h3f7ca6c7 /* (2, 10, 7) */,
  32'h3f7ca6c7 /* (14, 6, 7) */,
  32'h4039abaa /* (10, 6, 7) */,
  32'h4039abaa /* (6, 6, 7) */,
  32'h3f7ca6c7 /* (2, 6, 7) */,
  32'h3ec56b70 /* (14, 2, 7) */,
  32'h3f7ca6c7 /* (10, 2, 7) */,
  32'h3f7ca6c7 /* (6, 2, 7) */,
  32'h3ec56b70 /* (2, 2, 7) */,
  32'h3e9796af /* (14, 14, 3) */,
  32'h3ed22ea6 /* (10, 14, 3) */,
  32'h3ed22ea6 /* (6, 14, 3) */,
  32'h3e9796af /* (2, 14, 3) */,
  32'h3ed22ea6 /* (14, 10, 3) */,
  32'h3f7e11f4 /* (10, 10, 3) */,
  32'h3f7e11f4 /* (6, 10, 3) */,
  32'h3ed22ea6 /* (2, 10, 3) */,
  32'h3ed22ea6 /* (14, 6, 3) */,
  32'h3f7e11f4 /* (10, 6, 3) */,
  32'h3f7e11f4 /* (6, 6, 3) */,
  32'h3ed22ea6 /* (2, 6, 3) */,
  32'h3e9796af /* (14, 2, 3) */,
  32'h3ed22ea6 /* (10, 2, 3) */,
  32'h3ed22ea6 /* (6, 2, 3) */,
  32'h3e9796af /* (2, 2, 3) */,
  32'h3e9f2a5d /* (13, 14, 15) */,
  32'h3eb430e1 /* (9, 14, 15) */,
  32'h3e99eb68 /* (5, 14, 15) */,
  32'h3efc66bd /* (1, 14, 15) */,
  32'h3ec1987e /* (13, 10, 15) */,
  32'h3f62162b /* (9, 10, 15) */,
  32'h3f14d2ae /* (5, 10, 15) */,
  32'h3e9f454b /* (1, 10, 15) */,
  32'h3ec1987e /* (13, 6, 15) */,
  32'h3f62162b /* (9, 6, 15) */,
  32'h3f14d2ae /* (5, 6, 15) */,
  32'h3e9f454b /* (1, 6, 15) */,
  32'h3e9f2a5d /* (13, 2, 15) */,
  32'h3eb430e1 /* (9, 2, 15) */,
  32'h3e99eb68 /* (5, 2, 15) */,
  32'h3efc66bd /* (1, 2, 15) */,
  32'h3eb2cc97 /* (13, 14, 11) */,
  32'h3f3e2f24 /* (9, 14, 11) */,
  32'h3f025da2 /* (5, 14, 11) */,
  32'h3e99eb68 /* (1, 14, 11) */,
  32'h3f41f419 /* (13, 10, 11) */,
  32'h4006bd24 /* (9, 10, 11) */,
  32'h3fa39217 /* (5, 10, 11) */,
  32'h3f14d2ae /* (1, 10, 11) */,
  32'h3f41f419 /* (13, 6, 11) */,
  32'h4006bd24 /* (9, 6, 11) */,
  32'h3fa39217 /* (5, 6, 11) */,
  32'h3f14d2ae /* (1, 6, 11) */,
  32'h3eb2cc97 /* (13, 2, 11) */,
  32'h3f3e2f24 /* (9, 2, 11) */,
  32'h3f025da2 /* (5, 2, 11) */,
  32'h3e99eb68 /* (1, 2, 11) */,
  32'h3ee6ec8a /* (13, 14, 7) */,
  32'h3f993b79 /* (9, 14, 7) */,
  32'h3f3e2f24 /* (5, 14, 7) */,
  32'h3eb430e1 /* (1, 14, 7) */,
  32'h3f982d5a /* (13, 10, 7) */,
  32'h406912bc /* (9, 10, 7) */,
  32'h4006bd24 /* (5, 10, 7) */,
  32'h3f62162b /* (1, 10, 7) */,
  32'h3f982d5a /* (13, 6, 7) */,
  32'h406912bc /* (9, 6, 7) */,
  32'h4006bd24 /* (5, 6, 7) */,
  32'h3f62162b /* (1, 6, 7) */,
  32'h3ee6ec8a /* (13, 2, 7) */,
  32'h3f993b79 /* (9, 2, 7) */,
  32'h3f3e2f24 /* (5, 2, 7) */,
  32'h3eb430e1 /* (1, 2, 7) */,
  32'h3e9508f6 /* (13, 14, 3) */,
  32'h3ee6ec8a /* (9, 14, 3) */,
  32'h3eb2cc97 /* (5, 14, 3) */,
  32'h3e9f2a5d /* (1, 14, 3) */,
  32'h3ef2a853 /* (13, 10, 3) */,
  32'h3f982d5a /* (9, 10, 3) */,
  32'h3f41f419 /* (5, 10, 3) */,
  32'h3ec1987e /* (1, 10, 3) */,
  32'h3ef2a853 /* (13, 6, 3) */,
  32'h3f982d5a /* (9, 6, 3) */,
  32'h3f41f419 /* (5, 6, 3) */,
  32'h3ec1987e /* (1, 6, 3) */,
  32'h3e9508f6 /* (13, 2, 3) */,
  32'h3ee6ec8a /* (9, 2, 3) */,
  32'h3eb2cc97 /* (5, 2, 3) */,
  32'h3e9f2a5d /* (1, 2, 3) */,
  32'h3e939519 /* (12, 14, 15) */,
  32'h3e9c5e8a /* (8, 14, 15) */,
  32'h3e939519 /* (4, 14, 15) */,
  32'h3f10451b /* (0, 14, 15) */,
  32'h3ee9b2a2 /* (12, 10, 15) */,
  32'h3f5576ec /* (8, 10, 15) */,
  32'h3ee9b2a2 /* (4, 10, 15) */,
  32'h3e9bd472 /* (0, 10, 15) */,
  32'h3ee9b2a2 /* (12, 6, 15) */,
  32'h3f5576ec /* (8, 6, 15) */,
  32'h3ee9b2a2 /* (4, 6, 15) */,
  32'h3e9bd472 /* (0, 6, 15) */,
  32'h3e939519 /* (12, 2, 15) */,
  32'h3e9c5e8a /* (8, 2, 15) */,
  32'h3e939519 /* (4, 2, 15) */,
  32'h3f10451b /* (0, 2, 15) */,
  32'h3ed1ff4c /* (12, 14, 11) */,
  32'h3f30df4f /* (8, 14, 11) */,
  32'h3ed1ff4c /* (4, 14, 11) */,
  32'h3e97b006 /* (0, 14, 11) */,
  32'h3f753c17 /* (12, 10, 11) */,
  32'h40037a14 /* (8, 10, 11) */,
  32'h3f753c17 /* (4, 10, 11) */,
  32'h3f1019ab /* (0, 10, 11) */,
  32'h3f753c17 /* (12, 6, 11) */,
  32'h40037a14 /* (8, 6, 11) */,
  32'h3f753c17 /* (4, 6, 11) */,
  32'h3f1019ab /* (0, 6, 11) */,
  32'h3ed1ff4c /* (12, 2, 11) */,
  32'h3f30df4f /* (8, 2, 11) */,
  32'h3ed1ff4c /* (4, 2, 11) */,
  32'h3e97b006 /* (0, 2, 11) */,
  32'h3f104c25 /* (12, 14, 7) */,
  32'h3f9420e3 /* (8, 14, 7) */,
  32'h3f104c25 /* (4, 14, 7) */,
  32'h3eaee5c8 /* (0, 14, 7) */,
  32'h3fc4fc22 /* (12, 10, 7) */,
  32'h40686d0d /* (8, 10, 7) */,
  32'h3fc4fc22 /* (4, 10, 7) */,
  32'h3f59ea43 /* (0, 10, 7) */,
  32'h3fc4fc22 /* (12, 6, 7) */,
  32'h40686d0d /* (8, 6, 7) */,
  32'h3fc4fc22 /* (4, 6, 7) */,
  32'h3f59ea43 /* (0, 6, 7) */,
  32'h3f104c25 /* (12, 2, 7) */,
  32'h3f9420e3 /* (8, 2, 7) */,
  32'h3f104c25 /* (4, 2, 7) */,
  32'h3eaee5c8 /* (0, 2, 7) */,
  32'h3e9d3fef /* (12, 14, 3) */,
  32'h3ece2dc1 /* (8, 14, 3) */,
  32'h3e9d3fef /* (4, 14, 3) */,
  32'h3ea34ae8 /* (0, 14, 3) */,
  32'h3f15625b /* (12, 10, 3) */,
  32'h3f91854a /* (8, 10, 3) */,
  32'h3f15625b /* (4, 10, 3) */,
  32'h3ebc86f4 /* (0, 10, 3) */,
  32'h3f15625b /* (12, 6, 3) */,
  32'h3f91854a /* (8, 6, 3) */,
  32'h3f15625b /* (4, 6, 3) */,
  32'h3ebc86f4 /* (0, 6, 3) */,
  32'h3e9d3fef /* (12, 2, 3) */,
  32'h3ece2dc1 /* (8, 2, 3) */,
  32'h3e9d3fef /* (4, 2, 3) */,
  32'h3ea34ae8 /* (0, 2, 3) */,
  32'h3eaf2a10 /* (15, 13, 15) */,
  32'h3ea7dbb1 /* (11, 13, 15) */,
  32'h3ed1d4cb /* (7, 13, 15) */,
  32'h3e953797 /* (3, 13, 15) */,
  32'h3ea4f994 /* (15, 9, 15) */,
  32'h3f2b075a /* (11, 9, 15) */,
  32'h3f88838c /* (7, 9, 15) */,
  32'h3ed1d4cb /* (3, 9, 15) */,
  32'h3e93e191 /* (15, 5, 15) */,
  32'h3eeeb6df /* (11, 5, 15) */,
  32'h3f2b075a /* (7, 5, 15) */,
  32'h3ea7dbb1 /* (3, 5, 15) */,
  32'h3f5a3fd8 /* (15, 1, 15) */,
  32'h3e93e191 /* (11, 1, 15) */,
  32'h3ea4f994 /* (7, 1, 15) */,
  32'h3eaf2a10 /* (3, 1, 15) */,
  32'h3ea7dbb1 /* (15, 13, 11) */,
  32'h3f17cf64 /* (11, 13, 11) */,
  32'h3f6365d6 /* (7, 13, 11) */,
  32'h3ec9097c /* (3, 13, 11) */,
  32'h3f2b075a /* (15, 9, 11) */,
  32'h3fc5882d /* (11, 9, 11) */,
  32'h40278361 /* (7, 9, 11) */,
  32'h3f6365d6 /* (3, 9, 11) */,
  32'h3eeeb6df /* (15, 5, 11) */,
  32'h3f77795a /* (11, 5, 11) */,
  32'h3fc5882d /* (7, 5, 11) */,
  32'h3f17cf64 /* (3, 5, 11) */,
  32'h3e93e191 /* (15, 1, 11) */,
  32'h3eeeb6df /* (11, 1, 11) */,
  32'h3f2b075a /* (7, 1, 11) */,
  32'h3ea7dbb1 /* (3, 1, 11) */,
  32'h3ed1d4cb /* (15, 13, 7) */,
  32'h3f6365d6 /* (11, 13, 7) */,
  32'h3fb9d98f /* (7, 13, 7) */,
  32'h3f07f0f8 /* (3, 13, 7) */,
  32'h3f88838c /* (15, 9, 7) */,
  32'h40278361 /* (11, 9, 7) */,
  32'h4093adcc /* (7, 9, 7) */,
  32'h3fb9d98f /* (3, 9, 7) */,
  32'h3f2b075a /* (15, 5, 7) */,
  32'h3fc5882d /* (11, 5, 7) */,
  32'h40278361 /* (7, 5, 7) */,
  32'h3f6365d6 /* (3, 5, 7) */,
  32'h3ea4f994 /* (15, 1, 7) */,
  32'h3f2b075a /* (11, 1, 7) */,
  32'h3f88838c /* (7, 1, 7) */,
  32'h3ed1d4cb /* (3, 1, 7) */,
  32'h3e953797 /* (15, 13, 3) */,
  32'h3ec9097c /* (11, 13, 3) */,
  32'h3f07f0f8 /* (7, 13, 3) */,
  32'h3e9a814a /* (3, 13, 3) */,
  32'h3ed1d4cb /* (15, 9, 3) */,
  32'h3f6365d6 /* (11, 9, 3) */,
  32'h3fb9d98f /* (7, 9, 3) */,
  32'h3f07f0f8 /* (3, 9, 3) */,
  32'h3ea7dbb1 /* (15, 5, 3) */,
  32'h3f17cf64 /* (11, 5, 3) */,
  32'h3f6365d6 /* (7, 5, 3) */,
  32'h3ec9097c /* (3, 5, 3) */,
  32'h3eaf2a10 /* (15, 1, 3) */,
  32'h3ea7dbb1 /* (11, 1, 3) */,
  32'h3ed1d4cb /* (7, 1, 3) */,
  32'h3e953797 /* (3, 1, 3) */,
  32'h3e9f2a5d /* (14, 13, 15) */,
  32'h3ec1987e /* (10, 13, 15) */,
  32'h3ec1987e /* (6, 13, 15) */,
  32'h3e9f2a5d /* (2, 13, 15) */,
  32'h3eb430e1 /* (14, 9, 15) */,
  32'h3f62162b /* (10, 9, 15) */,
  32'h3f62162b /* (6, 9, 15) */,
  32'h3eb430e1 /* (2, 9, 15) */,
  32'h3e99eb68 /* (14, 5, 15) */,
  32'h3f14d2ae /* (10, 5, 15) */,
  32'h3f14d2ae /* (6, 5, 15) */,
  32'h3e99eb68 /* (2, 5, 15) */,
  32'h3efc66bd /* (14, 1, 15) */,
  32'h3e9f454b /* (10, 1, 15) */,
  32'h3e9f454b /* (6, 1, 15) */,
  32'h3efc66bd /* (2, 1, 15) */,
  32'h3eb2cc97 /* (14, 13, 11) */,
  32'h3f41f419 /* (10, 13, 11) */,
  32'h3f41f419 /* (6, 13, 11) */,
  32'h3eb2cc97 /* (2, 13, 11) */,
  32'h3f3e2f24 /* (14, 9, 11) */,
  32'h4006bd24 /* (10, 9, 11) */,
  32'h4006bd24 /* (6, 9, 11) */,
  32'h3f3e2f24 /* (2, 9, 11) */,
  32'h3f025da2 /* (14, 5, 11) */,
  32'h3fa39217 /* (10, 5, 11) */,
  32'h3fa39217 /* (6, 5, 11) */,
  32'h3f025da2 /* (2, 5, 11) */,
  32'h3e99eb68 /* (14, 1, 11) */,
  32'h3f14d2ae /* (10, 1, 11) */,
  32'h3f14d2ae /* (6, 1, 11) */,
  32'h3e99eb68 /* (2, 1, 11) */,
  32'h3ee6ec8a /* (14, 13, 7) */,
  32'h3f982d5a /* (10, 13, 7) */,
  32'h3f982d5a /* (6, 13, 7) */,
  32'h3ee6ec8a /* (2, 13, 7) */,
  32'h3f993b79 /* (14, 9, 7) */,
  32'h406912bc /* (10, 9, 7) */,
  32'h406912bc /* (6, 9, 7) */,
  32'h3f993b79 /* (2, 9, 7) */,
  32'h3f3e2f24 /* (14, 5, 7) */,
  32'h4006bd24 /* (10, 5, 7) */,
  32'h4006bd24 /* (6, 5, 7) */,
  32'h3f3e2f24 /* (2, 5, 7) */,
  32'h3eb430e1 /* (14, 1, 7) */,
  32'h3f62162b /* (10, 1, 7) */,
  32'h3f62162b /* (6, 1, 7) */,
  32'h3eb430e1 /* (2, 1, 7) */,
  32'h3e9508f6 /* (14, 13, 3) */,
  32'h3ef2a853 /* (10, 13, 3) */,
  32'h3ef2a853 /* (6, 13, 3) */,
  32'h3e9508f6 /* (2, 13, 3) */,
  32'h3ee6ec8a /* (14, 9, 3) */,
  32'h3f982d5a /* (10, 9, 3) */,
  32'h3f982d5a /* (6, 9, 3) */,
  32'h3ee6ec8a /* (2, 9, 3) */,
  32'h3eb2cc97 /* (14, 5, 3) */,
  32'h3f41f419 /* (10, 5, 3) */,
  32'h3f41f419 /* (6, 5, 3) */,
  32'h3eb2cc97 /* (2, 5, 3) */,
  32'h3e9f2a5d /* (14, 1, 3) */,
  32'h3ec1987e /* (10, 1, 3) */,
  32'h3ec1987e /* (6, 1, 3) */,
  32'h3e9f2a5d /* (2, 1, 3) */,
  32'h3e953797 /* (13, 13, 15) */,
  32'h3ed1d4cb /* (9, 13, 15) */,
  32'h3ea7dbb1 /* (5, 13, 15) */,
  32'h3eaf2a10 /* (1, 13, 15) */,
  32'h3ed1d4cb /* (13, 9, 15) */,
  32'h3f88838c /* (9, 9, 15) */,
  32'h3f2b075a /* (5, 9, 15) */,
  32'h3ea4f994 /* (1, 9, 15) */,
  32'h3ea7dbb1 /* (13, 5, 15) */,
  32'h3f2b075a /* (9, 5, 15) */,
  32'h3eeeb6df /* (5, 5, 15) */,
  32'h3e93e191 /* (1, 5, 15) */,
  32'h3eaf2a10 /* (13, 1, 15) */,
  32'h3ea4f994 /* (9, 1, 15) */,
  32'h3e93e191 /* (5, 1, 15) */,
  32'h3f5a3fd8 /* (1, 1, 15) */,
  32'h3ec9097c /* (13, 13, 11) */,
  32'h3f6365d6 /* (9, 13, 11) */,
  32'h3f17cf64 /* (5, 13, 11) */,
  32'h3ea7dbb1 /* (1, 13, 11) */,
  32'h3f6365d6 /* (13, 9, 11) */,
  32'h40278361 /* (9, 9, 11) */,
  32'h3fc5882d /* (5, 9, 11) */,
  32'h3f2b075a /* (1, 9, 11) */,
  32'h3f17cf64 /* (13, 5, 11) */,
  32'h3fc5882d /* (9, 5, 11) */,
  32'h3f77795a /* (5, 5, 11) */,
  32'h3eeeb6df /* (1, 5, 11) */,
  32'h3ea7dbb1 /* (13, 1, 11) */,
  32'h3f2b075a /* (9, 1, 11) */,
  32'h3eeeb6df /* (5, 1, 11) */,
  32'h3e93e191 /* (1, 1, 11) */,
  32'h3f07f0f8 /* (13, 13, 7) */,
  32'h3fb9d98f /* (9, 13, 7) */,
  32'h3f6365d6 /* (5, 13, 7) */,
  32'h3ed1d4cb /* (1, 13, 7) */,
  32'h3fb9d98f /* (13, 9, 7) */,
  32'h4093adcc /* (9, 9, 7) */,
  32'h40278361 /* (5, 9, 7) */,
  32'h3f88838c /* (1, 9, 7) */,
  32'h3f6365d6 /* (13, 5, 7) */,
  32'h40278361 /* (9, 5, 7) */,
  32'h3fc5882d /* (5, 5, 7) */,
  32'h3f2b075a /* (1, 5, 7) */,
  32'h3ed1d4cb /* (13, 1, 7) */,
  32'h3f88838c /* (9, 1, 7) */,
  32'h3f2b075a /* (5, 1, 7) */,
  32'h3ea4f994 /* (1, 1, 7) */,
  32'h3e9a814a /* (13, 13, 3) */,
  32'h3f07f0f8 /* (9, 13, 3) */,
  32'h3ec9097c /* (5, 13, 3) */,
  32'h3e953797 /* (1, 13, 3) */,
  32'h3f07f0f8 /* (13, 9, 3) */,
  32'h3fb9d98f /* (9, 9, 3) */,
  32'h3f6365d6 /* (5, 9, 3) */,
  32'h3ed1d4cb /* (1, 9, 3) */,
  32'h3ec9097c /* (13, 5, 3) */,
  32'h3f6365d6 /* (9, 5, 3) */,
  32'h3f17cf64 /* (5, 5, 3) */,
  32'h3ea7dbb1 /* (1, 5, 3) */,
  32'h3e953797 /* (13, 1, 3) */,
  32'h3ed1d4cb /* (9, 1, 3) */,
  32'h3ea7dbb1 /* (5, 1, 3) */,
  32'h3eaf2a10 /* (1, 1, 3) */,
  32'h3e97a967 /* (12, 13, 15) */,
  32'h3eb9823a /* (8, 13, 15) */,
  32'h3e97a967 /* (4, 13, 15) */,
  32'h3eb78ea1 /* (0, 13, 15) */,
  32'h3f0271c0 /* (12, 9, 15) */,
  32'h3f8374c7 /* (8, 9, 15) */,
  32'h3f0271c0 /* (4, 9, 15) */,
  32'h3ea04e75 /* (0, 9, 15) */,
  32'h3ec28d9a /* (12, 5, 15) */,
  32'h3f1e09be /* (8, 5, 15) */,
  32'h3ec28d9a /* (4, 5, 15) */,
  32'h3e924c17 /* (0, 5, 15) */,
  32'h3e94e1d9 /* (12, 1, 15) */,
  32'h3e8d5b73 /* (8, 1, 15) */,
  32'h3e94e1d9 /* (4, 1, 15) */,
  32'h3f9befb2 /* (0, 1, 15) */,
  32'h3ef076ff /* (12, 13, 11) */,
  32'h3f558e61 /* (8, 13, 11) */,
  32'h3ef076ff /* (4, 13, 11) */,
  32'h3ea49cf9 /* (0, 13, 11) */,
  32'h3f91d65e /* (12, 9, 11) */,
  32'h40258eba /* (8, 9, 11) */,
  32'h3f91d65e /* (4, 9, 11) */,
  32'h3f2521d3 /* (0, 9, 11) */,
  32'h3f3cbfdf /* (12, 5, 11) */,
  32'h3fbe36ae /* (8, 5, 11) */,
  32'h3f3cbfdf /* (4, 5, 11) */,
  32'h3ee7f590 /* (0, 5, 11) */,
  32'h3ec28d9a /* (12, 1, 11) */,
  32'h3f1e09be /* (8, 1, 11) */,
  32'h3ec28d9a /* (4, 1, 11) */,
  32'h3e924c17 /* (0, 1, 11) */,
  32'h3f2b2ff1 /* (12, 13, 7) */,
  32'h3fb4be0d /* (8, 13, 7) */,
  32'h3f2b2ff1 /* (4, 13, 7) */,
  32'h3ecb578e /* (0, 13, 7) */,
  32'h3ff29d82 /* (12, 9, 7) */,
  32'h4094977b /* (8, 9, 7) */,
  32'h3ff29d82 /* (4, 9, 7) */,
  32'h3f836079 /* (0, 9, 7) */,
  32'h3f91d65e /* (12, 5, 7) */,
  32'h40258eba /* (8, 5, 7) */,
  32'h3f91d65e /* (4, 5, 7) */,
  32'h3f2521d3 /* (0, 5, 7) */,
  32'h3f0271c0 /* (12, 1, 7) */,
  32'h3f8374c7 /* (8, 1, 7) */,
  32'h3f0271c0 /* (4, 1, 7) */,
  32'h3ea04e75 /* (0, 1, 7) */,
  32'h3eaaa637 /* (12, 13, 3) */,
  32'h3ef65451 /* (8, 13, 3) */,
  32'h3eaaa637 /* (4, 13, 3) */,
  32'h3e960c85 /* (0, 13, 3) */,
  32'h3f2b2ff1 /* (12, 9, 3) */,
  32'h3fb4be0d /* (8, 9, 3) */,
  32'h3f2b2ff1 /* (4, 9, 3) */,
  32'h3ecb578e /* (0, 9, 3) */,
  32'h3ef076ff /* (12, 5, 3) */,
  32'h3f558e61 /* (8, 5, 3) */,
  32'h3ef076ff /* (4, 5, 3) */,
  32'h3ea49cf9 /* (0, 5, 3) */,
  32'h3e97a967 /* (12, 1, 3) */,
  32'h3eb9823a /* (8, 1, 3) */,
  32'h3e97a967 /* (4, 1, 3) */,
  32'h3eb78ea1 /* (0, 1, 3) */,
  32'h3e94e1d9 /* (15, 12, 15) */,
  32'h3ec28d9a /* (11, 12, 15) */,
  32'h3f0271c0 /* (7, 12, 15) */,
  32'h3e97a967 /* (3, 12, 15) */,
  32'h3e8d5b73 /* (15, 8, 15) */,
  32'h3f1e09be /* (11, 8, 15) */,
  32'h3f8374c7 /* (7, 8, 15) */,
  32'h3eb9823a /* (3, 8, 15) */,
  32'h3e94e1d9 /* (15, 4, 15) */,
  32'h3ec28d9a /* (11, 4, 15) */,
  32'h3f0271c0 /* (7, 4, 15) */,
  32'h3e97a967 /* (3, 4, 15) */,
  32'h3f9befb2 /* (15, 0, 15) */,
  32'h3e924c17 /* (11, 0, 15) */,
  32'h3ea04e75 /* (7, 0, 15) */,
  32'h3eb78ea1 /* (3, 0, 15) */,
  32'h3ec28d9a /* (15, 12, 11) */,
  32'h3f3cbfdf /* (11, 12, 11) */,
  32'h3f91d65e /* (7, 12, 11) */,
  32'h3ef076ff /* (3, 12, 11) */,
  32'h3f1e09be /* (15, 8, 11) */,
  32'h3fbe36ae /* (11, 8, 11) */,
  32'h40258eba /* (7, 8, 11) */,
  32'h3f558e61 /* (3, 8, 11) */,
  32'h3ec28d9a /* (15, 4, 11) */,
  32'h3f3cbfdf /* (11, 4, 11) */,
  32'h3f91d65e /* (7, 4, 11) */,
  32'h3ef076ff /* (3, 4, 11) */,
  32'h3e924c17 /* (15, 0, 11) */,
  32'h3ee7f590 /* (11, 0, 11) */,
  32'h3f2521d3 /* (7, 0, 11) */,
  32'h3ea49cf9 /* (3, 0, 11) */,
  32'h3f0271c0 /* (15, 12, 7) */,
  32'h3f91d65e /* (11, 12, 7) */,
  32'h3ff29d82 /* (7, 12, 7) */,
  32'h3f2b2ff1 /* (3, 12, 7) */,
  32'h3f8374c7 /* (15, 8, 7) */,
  32'h40258eba /* (11, 8, 7) */,
  32'h4094977b /* (7, 8, 7) */,
  32'h3fb4be0d /* (3, 8, 7) */,
  32'h3f0271c0 /* (15, 4, 7) */,
  32'h3f91d65e /* (11, 4, 7) */,
  32'h3ff29d82 /* (7, 4, 7) */,
  32'h3f2b2ff1 /* (3, 4, 7) */,
  32'h3ea04e75 /* (15, 0, 7) */,
  32'h3f2521d3 /* (11, 0, 7) */,
  32'h3f836079 /* (7, 0, 7) */,
  32'h3ecb578e /* (3, 0, 7) */,
  32'h3e97a967 /* (15, 12, 3) */,
  32'h3ef076ff /* (11, 12, 3) */,
  32'h3f2b2ff1 /* (7, 12, 3) */,
  32'h3eaaa637 /* (3, 12, 3) */,
  32'h3eb9823a /* (15, 8, 3) */,
  32'h3f558e61 /* (11, 8, 3) */,
  32'h3fb4be0d /* (7, 8, 3) */,
  32'h3ef65451 /* (3, 8, 3) */,
  32'h3e97a967 /* (15, 4, 3) */,
  32'h3ef076ff /* (11, 4, 3) */,
  32'h3f2b2ff1 /* (7, 4, 3) */,
  32'h3eaaa637 /* (3, 4, 3) */,
  32'h3eb78ea1 /* (15, 0, 3) */,
  32'h3ea49cf9 /* (11, 0, 3) */,
  32'h3ecb578e /* (7, 0, 3) */,
  32'h3e960c85 /* (3, 0, 3) */,
  32'h3e939519 /* (14, 12, 15) */,
  32'h3ee9b2a2 /* (10, 12, 15) */,
  32'h3ee9b2a2 /* (6, 12, 15) */,
  32'h3e939519 /* (2, 12, 15) */,
  32'h3e9c5e8a /* (14, 8, 15) */,
  32'h3f5576ec /* (10, 8, 15) */,
  32'h3f5576ec /* (6, 8, 15) */,
  32'h3e9c5e8a /* (2, 8, 15) */,
  32'h3e939519 /* (14, 4, 15) */,
  32'h3ee9b2a2 /* (10, 4, 15) */,
  32'h3ee9b2a2 /* (6, 4, 15) */,
  32'h3e939519 /* (2, 4, 15) */,
  32'h3f10451b /* (14, 0, 15) */,
  32'h3e9bd472 /* (10, 0, 15) */,
  32'h3e9bd472 /* (6, 0, 15) */,
  32'h3f10451b /* (2, 0, 15) */,
  32'h3ed1ff4c /* (14, 12, 11) */,
  32'h3f753c17 /* (10, 12, 11) */,
  32'h3f753c17 /* (6, 12, 11) */,
  32'h3ed1ff4c /* (2, 12, 11) */,
  32'h3f30df4f /* (14, 8, 11) */,
  32'h40037a14 /* (10, 8, 11) */,
  32'h40037a14 /* (6, 8, 11) */,
  32'h3f30df4f /* (2, 8, 11) */,
  32'h3ed1ff4c /* (14, 4, 11) */,
  32'h3f753c17 /* (10, 4, 11) */,
  32'h3f753c17 /* (6, 4, 11) */,
  32'h3ed1ff4c /* (2, 4, 11) */,
  32'h3e97b006 /* (14, 0, 11) */,
  32'h3f1019ab /* (10, 0, 11) */,
  32'h3f1019ab /* (6, 0, 11) */,
  32'h3e97b006 /* (2, 0, 11) */,
  32'h3f104c25 /* (14, 12, 7) */,
  32'h3fc4fc22 /* (10, 12, 7) */,
  32'h3fc4fc22 /* (6, 12, 7) */,
  32'h3f104c25 /* (2, 12, 7) */,
  32'h3f9420e3 /* (14, 8, 7) */,
  32'h40686d0d /* (10, 8, 7) */,
  32'h40686d0d /* (6, 8, 7) */,
  32'h3f9420e3 /* (2, 8, 7) */,
  32'h3f104c25 /* (14, 4, 7) */,
  32'h3fc4fc22 /* (10, 4, 7) */,
  32'h3fc4fc22 /* (6, 4, 7) */,
  32'h3f104c25 /* (2, 4, 7) */,
  32'h3eaee5c8 /* (14, 0, 7) */,
  32'h3f59ea43 /* (10, 0, 7) */,
  32'h3f59ea43 /* (6, 0, 7) */,
  32'h3eaee5c8 /* (2, 0, 7) */,
  32'h3e9d3fef /* (14, 12, 3) */,
  32'h3f15625b /* (10, 12, 3) */,
  32'h3f15625b /* (6, 12, 3) */,
  32'h3e9d3fef /* (2, 12, 3) */,
  32'h3ece2dc1 /* (14, 8, 3) */,
  32'h3f91854a /* (10, 8, 3) */,
  32'h3f91854a /* (6, 8, 3) */,
  32'h3ece2dc1 /* (2, 8, 3) */,
  32'h3e9d3fef /* (14, 4, 3) */,
  32'h3f15625b /* (10, 4, 3) */,
  32'h3f15625b /* (6, 4, 3) */,
  32'h3e9d3fef /* (2, 4, 3) */,
  32'h3ea34ae8 /* (14, 0, 3) */,
  32'h3ebc86f4 /* (10, 0, 3) */,
  32'h3ebc86f4 /* (6, 0, 3) */,
  32'h3ea34ae8 /* (2, 0, 3) */,
  32'h3e97a967 /* (13, 12, 15) */,
  32'h3f0271c0 /* (9, 12, 15) */,
  32'h3ec28d9a /* (5, 12, 15) */,
  32'h3e94e1d9 /* (1, 12, 15) */,
  32'h3eb9823a /* (13, 8, 15) */,
  32'h3f8374c7 /* (9, 8, 15) */,
  32'h3f1e09be /* (5, 8, 15) */,
  32'h3e8d5b73 /* (1, 8, 15) */,
  32'h3e97a967 /* (13, 4, 15) */,
  32'h3f0271c0 /* (9, 4, 15) */,
  32'h3ec28d9a /* (5, 4, 15) */,
  32'h3e94e1d9 /* (1, 4, 15) */,
  32'h3eb78ea1 /* (13, 0, 15) */,
  32'h3ea04e75 /* (9, 0, 15) */,
  32'h3e924c17 /* (5, 0, 15) */,
  32'h3f9befb2 /* (1, 0, 15) */,
  32'h3ef076ff /* (13, 12, 11) */,
  32'h3f91d65e /* (9, 12, 11) */,
  32'h3f3cbfdf /* (5, 12, 11) */,
  32'h3ec28d9a /* (1, 12, 11) */,
  32'h3f558e61 /* (13, 8, 11) */,
  32'h40258eba /* (9, 8, 11) */,
  32'h3fbe36ae /* (5, 8, 11) */,
  32'h3f1e09be /* (1, 8, 11) */,
  32'h3ef076ff /* (13, 4, 11) */,
  32'h3f91d65e /* (9, 4, 11) */,
  32'h3f3cbfdf /* (5, 4, 11) */,
  32'h3ec28d9a /* (1, 4, 11) */,
  32'h3ea49cf9 /* (13, 0, 11) */,
  32'h3f2521d3 /* (9, 0, 11) */,
  32'h3ee7f590 /* (5, 0, 11) */,
  32'h3e924c17 /* (1, 0, 11) */,
  32'h3f2b2ff1 /* (13, 12, 7) */,
  32'h3ff29d82 /* (9, 12, 7) */,
  32'h3f91d65e /* (5, 12, 7) */,
  32'h3f0271c0 /* (1, 12, 7) */,
  32'h3fb4be0d /* (13, 8, 7) */,
  32'h4094977b /* (9, 8, 7) */,
  32'h40258eba /* (5, 8, 7) */,
  32'h3f8374c7 /* (1, 8, 7) */,
  32'h3f2b2ff1 /* (13, 4, 7) */,
  32'h3ff29d82 /* (9, 4, 7) */,
  32'h3f91d65e /* (5, 4, 7) */,
  32'h3f0271c0 /* (1, 4, 7) */,
  32'h3ecb578e /* (13, 0, 7) */,
  32'h3f836079 /* (9, 0, 7) */,
  32'h3f2521d3 /* (5, 0, 7) */,
  32'h3ea04e75 /* (1, 0, 7) */,
  32'h3eaaa637 /* (13, 12, 3) */,
  32'h3f2b2ff1 /* (9, 12, 3) */,
  32'h3ef076ff /* (5, 12, 3) */,
  32'h3e97a967 /* (1, 12, 3) */,
  32'h3ef65451 /* (13, 8, 3) */,
  32'h3fb4be0d /* (9, 8, 3) */,
  32'h3f558e61 /* (5, 8, 3) */,
  32'h3eb9823a /* (1, 8, 3) */,
  32'h3eaaa637 /* (13, 4, 3) */,
  32'h3f2b2ff1 /* (9, 4, 3) */,
  32'h3ef076ff /* (5, 4, 3) */,
  32'h3e97a967 /* (1, 4, 3) */,
  32'h3e960c85 /* (13, 0, 3) */,
  32'h3ecb578e /* (9, 0, 3) */,
  32'h3ea49cf9 /* (5, 0, 3) */,
  32'h3eb78ea1 /* (1, 0, 3) */,
  32'h3ea63161 /* (12, 12, 15) */,
  32'h3eebb725 /* (8, 12, 15) */,
  32'h3ea63161 /* (4, 12, 15) */,
  32'h3e962cf4 /* (0, 12, 15) */,
  32'h3eebb725 /* (12, 8, 15) */,
  32'h3f80d0e8 /* (8, 8, 15) */,
  32'h3eebb725 /* (4, 8, 15) */,
  32'h3e88bc50 /* (0, 8, 15) */,
  32'h3ea63161 /* (12, 4, 15) */,
  32'h3eebb725 /* (8, 4, 15) */,
  32'h3ea63161 /* (4, 4, 15) */,
  32'h3e962cf4 /* (0, 4, 15) */,
  32'h3e962cf4 /* (12, 0, 15) */,
  32'h3e88bc50 /* (8, 0, 15) */,
  32'h3e962cf4 /* (4, 0, 15) */,
  32'h40148d77 /* (0, 0, 15) */,
  32'h3f12b00d /* (12, 12, 11) */,
  32'h3f8a9c45 /* (8, 12, 11) */,
  32'h3f12b00d /* (4, 12, 11) */,
  32'h3ebddc83 /* (0, 12, 11) */,
  32'h3f8a9c45 /* (12, 8, 11) */,
  32'h402594bb /* (8, 8, 11) */,
  32'h3f8a9c45 /* (4, 8, 11) */,
  32'h3f183f16 /* (0, 8, 11) */,
  32'h3f12b00d /* (12, 4, 11) */,
  32'h3f8a9c45 /* (8, 4, 11) */,
  32'h3f12b00d /* (4, 4, 11) */,
  32'h3ebddc83 /* (0, 4, 11) */,
  32'h3ebddc83 /* (12, 0, 11) */,
  32'h3f183f16 /* (8, 0, 11) */,
  32'h3ebddc83 /* (4, 0, 11) */,
  32'h3e90f1d9 /* (0, 0, 11) */,
  32'h3f59849a /* (12, 12, 7) */,
  32'h3fedbe1f /* (8, 12, 7) */,
  32'h3f59849a /* (4, 12, 7) */,
  32'h3efc5be6 /* (0, 12, 7) */,
  32'h3fedbe1f /* (12, 8, 7) */,
  32'h4096cd97 /* (8, 8, 7) */,
  32'h3fedbe1f /* (4, 8, 7) */,
  32'h3f7cadff /* (0, 8, 7) */,
  32'h3f59849a /* (12, 4, 7) */,
  32'h3fedbe1f /* (8, 4, 7) */,
  32'h3f59849a /* (4, 4, 7) */,
  32'h3efc5be6 /* (0, 4, 7) */,
  32'h3efc5be6 /* (12, 0, 7) */,
  32'h3f7cadff /* (8, 0, 7) */,
  32'h3efc5be6 /* (4, 0, 7) */,
  32'h3e9bd51d /* (0, 0, 7) */,
  32'h3ec4d2c5 /* (12, 12, 3) */,
  32'h3f1dd43f /* (8, 12, 3) */,
  32'h3ec4d2c5 /* (4, 12, 3) */,
  32'h3e964277 /* (0, 12, 3) */,
  32'h3f1dd43f /* (12, 8, 3) */,
  32'h3fb27927 /* (8, 8, 3) */,
  32'h3f1dd43f /* (4, 8, 3) */,
  32'h3eb32545 /* (0, 8, 3) */,
  32'h3ec4d2c5 /* (12, 4, 3) */,
  32'h3f1dd43f /* (8, 4, 3) */,
  32'h3ec4d2c5 /* (4, 4, 3) */,
  32'h3e964277 /* (0, 4, 3) */,
  32'h3e964277 /* (12, 0, 3) */,
  32'h3eb32545 /* (8, 0, 3) */,
  32'h3e964277 /* (4, 0, 3) */,
  32'h3ec24b89 /* (0, 0, 3) */,
  32'h3efc66bd /* (15, 15, 14) */,
  32'h3e99eb68 /* (11, 15, 14) */,
  32'h3eb430e1 /* (7, 15, 14) */,
  32'h3e9f2a5d /* (3, 15, 14) */,
  32'h3e99eb68 /* (15, 11, 14) */,
  32'h3f025da2 /* (11, 11, 14) */,
  32'h3f3e2f24 /* (7, 11, 14) */,
  32'h3eb2cc97 /* (3, 11, 14) */,
  32'h3eb430e1 /* (15, 7, 14) */,
  32'h3f3e2f24 /* (11, 7, 14) */,
  32'h3f993b79 /* (7, 7, 14) */,
  32'h3ee6ec8a /* (3, 7, 14) */,
  32'h3e9f2a5d /* (15, 3, 14) */,
  32'h3eb2cc97 /* (11, 3, 14) */,
  32'h3ee6ec8a /* (7, 3, 14) */,
  32'h3e9508f6 /* (3, 3, 14) */,
  32'h3e9f454b /* (15, 15, 10) */,
  32'h3f14d2ae /* (11, 15, 10) */,
  32'h3f62162b /* (7, 15, 10) */,
  32'h3ec1987e /* (3, 15, 10) */,
  32'h3f14d2ae /* (15, 11, 10) */,
  32'h3fa39217 /* (11, 11, 10) */,
  32'h4006bd24 /* (7, 11, 10) */,
  32'h3f41f419 /* (3, 11, 10) */,
  32'h3f62162b /* (15, 7, 10) */,
  32'h4006bd24 /* (11, 7, 10) */,
  32'h406912bc /* (7, 7, 10) */,
  32'h3f982d5a /* (3, 7, 10) */,
  32'h3ec1987e /* (15, 3, 10) */,
  32'h3f41f419 /* (11, 3, 10) */,
  32'h3f982d5a /* (7, 3, 10) */,
  32'h3ef2a853 /* (3, 3, 10) */,
  32'h3e9f454b /* (15, 15, 6) */,
  32'h3f14d2ae /* (11, 15, 6) */,
  32'h3f62162b /* (7, 15, 6) */,
  32'h3ec1987e /* (3, 15, 6) */,
  32'h3f14d2ae /* (15, 11, 6) */,
  32'h3fa39217 /* (11, 11, 6) */,
  32'h4006bd24 /* (7, 11, 6) */,
  32'h3f41f419 /* (3, 11, 6) */,
  32'h3f62162b /* (15, 7, 6) */,
  32'h4006bd24 /* (11, 7, 6) */,
  32'h406912bc /* (7, 7, 6) */,
  32'h3f982d5a /* (3, 7, 6) */,
  32'h3ec1987e /* (15, 3, 6) */,
  32'h3f41f419 /* (11, 3, 6) */,
  32'h3f982d5a /* (7, 3, 6) */,
  32'h3ef2a853 /* (3, 3, 6) */,
  32'h3efc66bd /* (15, 15, 2) */,
  32'h3e99eb68 /* (11, 15, 2) */,
  32'h3eb430e1 /* (7, 15, 2) */,
  32'h3e9f2a5d /* (3, 15, 2) */,
  32'h3e99eb68 /* (15, 11, 2) */,
  32'h3f025da2 /* (11, 11, 2) */,
  32'h3f3e2f24 /* (7, 11, 2) */,
  32'h3eb2cc97 /* (3, 11, 2) */,
  32'h3eb430e1 /* (15, 7, 2) */,
  32'h3f3e2f24 /* (11, 7, 2) */,
  32'h3f993b79 /* (7, 7, 2) */,
  32'h3ee6ec8a /* (3, 7, 2) */,
  32'h3e9f2a5d /* (15, 3, 2) */,
  32'h3eb2cc97 /* (11, 3, 2) */,
  32'h3ee6ec8a /* (7, 3, 2) */,
  32'h3e9508f6 /* (3, 3, 2) */,
  32'h3ec29928 /* (14, 15, 14) */,
  32'h3eaab74a /* (10, 15, 14) */,
  32'h3eaab74a /* (6, 15, 14) */,
  32'h3ec29928 /* (2, 15, 14) */,
  32'h3ea1d2a3 /* (14, 11, 14) */,
  32'h3f242ada /* (10, 11, 14) */,
  32'h3f242ada /* (6, 11, 14) */,
  32'h3ea1d2a3 /* (2, 11, 14) */,
  32'h3ec56b70 /* (14, 7, 14) */,
  32'h3f7ca6c7 /* (10, 7, 14) */,
  32'h3f7ca6c7 /* (6, 7, 14) */,
  32'h3ec56b70 /* (2, 7, 14) */,
  32'h3e9796af /* (14, 3, 14) */,
  32'h3ed22ea6 /* (10, 3, 14) */,
  32'h3ed22ea6 /* (6, 3, 14) */,
  32'h3e9796af /* (2, 3, 14) */,
  32'h3eaab74a /* (14, 15, 10) */,
  32'h3f3f980b /* (10, 15, 10) */,
  32'h3f3f980b /* (6, 15, 10) */,
  32'h3eaab74a /* (2, 15, 10) */,
  32'h3f242ada /* (14, 11, 10) */,
  32'h3fdbd2f0 /* (10, 11, 10) */,
  32'h3fdbd2f0 /* (6, 11, 10) */,
  32'h3f242ada /* (2, 11, 10) */,
  32'h3f7ca6c7 /* (14, 7, 10) */,
  32'h4039abaa /* (10, 7, 10) */,
  32'h4039abaa /* (6, 7, 10) */,
  32'h3f7ca6c7 /* (2, 7, 10) */,
  32'h3ed22ea6 /* (14, 3, 10) */,
  32'h3f7e11f4 /* (10, 3, 10) */,
  32'h3f7e11f4 /* (6, 3, 10) */,
  32'h3ed22ea6 /* (2, 3, 10) */,
  32'h3eaab74a /* (14, 15, 6) */,
  32'h3f3f980b /* (10, 15, 6) */,
  32'h3f3f980b /* (6, 15, 6) */,
  32'h3eaab74a /* (2, 15, 6) */,
  32'h3f242ada /* (14, 11, 6) */,
  32'h3fdbd2f0 /* (10, 11, 6) */,
  32'h3fdbd2f0 /* (6, 11, 6) */,
  32'h3f242ada /* (2, 11, 6) */,
  32'h3f7ca6c7 /* (14, 7, 6) */,
  32'h4039abaa /* (10, 7, 6) */,
  32'h4039abaa /* (6, 7, 6) */,
  32'h3f7ca6c7 /* (2, 7, 6) */,
  32'h3ed22ea6 /* (14, 3, 6) */,
  32'h3f7e11f4 /* (10, 3, 6) */,
  32'h3f7e11f4 /* (6, 3, 6) */,
  32'h3ed22ea6 /* (2, 3, 6) */,
  32'h3ec29928 /* (14, 15, 2) */,
  32'h3eaab74a /* (10, 15, 2) */,
  32'h3eaab74a /* (6, 15, 2) */,
  32'h3ec29928 /* (2, 15, 2) */,
  32'h3ea1d2a3 /* (14, 11, 2) */,
  32'h3f242ada /* (10, 11, 2) */,
  32'h3f242ada /* (6, 11, 2) */,
  32'h3ea1d2a3 /* (2, 11, 2) */,
  32'h3ec56b70 /* (14, 7, 2) */,
  32'h3f7ca6c7 /* (10, 7, 2) */,
  32'h3f7ca6c7 /* (6, 7, 2) */,
  32'h3ec56b70 /* (2, 7, 2) */,
  32'h3e9796af /* (14, 3, 2) */,
  32'h3ed22ea6 /* (10, 3, 2) */,
  32'h3ed22ea6 /* (6, 3, 2) */,
  32'h3e9796af /* (2, 3, 2) */,
  32'h3e9f2a5d /* (13, 15, 14) */,
  32'h3eb430e1 /* (9, 15, 14) */,
  32'h3e99eb68 /* (5, 15, 14) */,
  32'h3efc66bd /* (1, 15, 14) */,
  32'h3eb2cc97 /* (13, 11, 14) */,
  32'h3f3e2f24 /* (9, 11, 14) */,
  32'h3f025da2 /* (5, 11, 14) */,
  32'h3e99eb68 /* (1, 11, 14) */,
  32'h3ee6ec8a /* (13, 7, 14) */,
  32'h3f993b79 /* (9, 7, 14) */,
  32'h3f3e2f24 /* (5, 7, 14) */,
  32'h3eb430e1 /* (1, 7, 14) */,
  32'h3e9508f6 /* (13, 3, 14) */,
  32'h3ee6ec8a /* (9, 3, 14) */,
  32'h3eb2cc97 /* (5, 3, 14) */,
  32'h3e9f2a5d /* (1, 3, 14) */,
  32'h3ec1987e /* (13, 15, 10) */,
  32'h3f62162b /* (9, 15, 10) */,
  32'h3f14d2ae /* (5, 15, 10) */,
  32'h3e9f454b /* (1, 15, 10) */,
  32'h3f41f419 /* (13, 11, 10) */,
  32'h4006bd24 /* (9, 11, 10) */,
  32'h3fa39217 /* (5, 11, 10) */,
  32'h3f14d2ae /* (1, 11, 10) */,
  32'h3f982d5a /* (13, 7, 10) */,
  32'h406912bc /* (9, 7, 10) */,
  32'h4006bd24 /* (5, 7, 10) */,
  32'h3f62162b /* (1, 7, 10) */,
  32'h3ef2a853 /* (13, 3, 10) */,
  32'h3f982d5a /* (9, 3, 10) */,
  32'h3f41f419 /* (5, 3, 10) */,
  32'h3ec1987e /* (1, 3, 10) */,
  32'h3ec1987e /* (13, 15, 6) */,
  32'h3f62162b /* (9, 15, 6) */,
  32'h3f14d2ae /* (5, 15, 6) */,
  32'h3e9f454b /* (1, 15, 6) */,
  32'h3f41f419 /* (13, 11, 6) */,
  32'h4006bd24 /* (9, 11, 6) */,
  32'h3fa39217 /* (5, 11, 6) */,
  32'h3f14d2ae /* (1, 11, 6) */,
  32'h3f982d5a /* (13, 7, 6) */,
  32'h406912bc /* (9, 7, 6) */,
  32'h4006bd24 /* (5, 7, 6) */,
  32'h3f62162b /* (1, 7, 6) */,
  32'h3ef2a853 /* (13, 3, 6) */,
  32'h3f982d5a /* (9, 3, 6) */,
  32'h3f41f419 /* (5, 3, 6) */,
  32'h3ec1987e /* (1, 3, 6) */,
  32'h3e9f2a5d /* (13, 15, 2) */,
  32'h3eb430e1 /* (9, 15, 2) */,
  32'h3e99eb68 /* (5, 15, 2) */,
  32'h3efc66bd /* (1, 15, 2) */,
  32'h3eb2cc97 /* (13, 11, 2) */,
  32'h3f3e2f24 /* (9, 11, 2) */,
  32'h3f025da2 /* (5, 11, 2) */,
  32'h3e99eb68 /* (1, 11, 2) */,
  32'h3ee6ec8a /* (13, 7, 2) */,
  32'h3f993b79 /* (9, 7, 2) */,
  32'h3f3e2f24 /* (5, 7, 2) */,
  32'h3eb430e1 /* (1, 7, 2) */,
  32'h3e9508f6 /* (13, 3, 2) */,
  32'h3ee6ec8a /* (9, 3, 2) */,
  32'h3eb2cc97 /* (5, 3, 2) */,
  32'h3e9f2a5d /* (1, 3, 2) */,
  32'h3e939519 /* (12, 15, 14) */,
  32'h3e9c5e8a /* (8, 15, 14) */,
  32'h3e939519 /* (4, 15, 14) */,
  32'h3f10451b /* (0, 15, 14) */,
  32'h3ed1ff4c /* (12, 11, 14) */,
  32'h3f30df4f /* (8, 11, 14) */,
  32'h3ed1ff4c /* (4, 11, 14) */,
  32'h3e97b006 /* (0, 11, 14) */,
  32'h3f104c25 /* (12, 7, 14) */,
  32'h3f9420e3 /* (8, 7, 14) */,
  32'h3f104c25 /* (4, 7, 14) */,
  32'h3eaee5c8 /* (0, 7, 14) */,
  32'h3e9d3fef /* (12, 3, 14) */,
  32'h3ece2dc1 /* (8, 3, 14) */,
  32'h3e9d3fef /* (4, 3, 14) */,
  32'h3ea34ae8 /* (0, 3, 14) */,
  32'h3ee9b2a2 /* (12, 15, 10) */,
  32'h3f5576ec /* (8, 15, 10) */,
  32'h3ee9b2a2 /* (4, 15, 10) */,
  32'h3e9bd472 /* (0, 15, 10) */,
  32'h3f753c17 /* (12, 11, 10) */,
  32'h40037a14 /* (8, 11, 10) */,
  32'h3f753c17 /* (4, 11, 10) */,
  32'h3f1019ab /* (0, 11, 10) */,
  32'h3fc4fc22 /* (12, 7, 10) */,
  32'h40686d0d /* (8, 7, 10) */,
  32'h3fc4fc22 /* (4, 7, 10) */,
  32'h3f59ea43 /* (0, 7, 10) */,
  32'h3f15625b /* (12, 3, 10) */,
  32'h3f91854a /* (8, 3, 10) */,
  32'h3f15625b /* (4, 3, 10) */,
  32'h3ebc86f4 /* (0, 3, 10) */,
  32'h3ee9b2a2 /* (12, 15, 6) */,
  32'h3f5576ec /* (8, 15, 6) */,
  32'h3ee9b2a2 /* (4, 15, 6) */,
  32'h3e9bd472 /* (0, 15, 6) */,
  32'h3f753c17 /* (12, 11, 6) */,
  32'h40037a14 /* (8, 11, 6) */,
  32'h3f753c17 /* (4, 11, 6) */,
  32'h3f1019ab /* (0, 11, 6) */,
  32'h3fc4fc22 /* (12, 7, 6) */,
  32'h40686d0d /* (8, 7, 6) */,
  32'h3fc4fc22 /* (4, 7, 6) */,
  32'h3f59ea43 /* (0, 7, 6) */,
  32'h3f15625b /* (12, 3, 6) */,
  32'h3f91854a /* (8, 3, 6) */,
  32'h3f15625b /* (4, 3, 6) */,
  32'h3ebc86f4 /* (0, 3, 6) */,
  32'h3e939519 /* (12, 15, 2) */,
  32'h3e9c5e8a /* (8, 15, 2) */,
  32'h3e939519 /* (4, 15, 2) */,
  32'h3f10451b /* (0, 15, 2) */,
  32'h3ed1ff4c /* (12, 11, 2) */,
  32'h3f30df4f /* (8, 11, 2) */,
  32'h3ed1ff4c /* (4, 11, 2) */,
  32'h3e97b006 /* (0, 11, 2) */,
  32'h3f104c25 /* (12, 7, 2) */,
  32'h3f9420e3 /* (8, 7, 2) */,
  32'h3f104c25 /* (4, 7, 2) */,
  32'h3eaee5c8 /* (0, 7, 2) */,
  32'h3e9d3fef /* (12, 3, 2) */,
  32'h3ece2dc1 /* (8, 3, 2) */,
  32'h3e9d3fef /* (4, 3, 2) */,
  32'h3ea34ae8 /* (0, 3, 2) */,
  32'h3ec29928 /* (15, 14, 14) */,
  32'h3ea1d2a3 /* (11, 14, 14) */,
  32'h3ec56b70 /* (7, 14, 14) */,
  32'h3e9796af /* (3, 14, 14) */,
  32'h3eaab74a /* (15, 10, 14) */,
  32'h3f242ada /* (11, 10, 14) */,
  32'h3f7ca6c7 /* (7, 10, 14) */,
  32'h3ed22ea6 /* (3, 10, 14) */,
  32'h3eaab74a /* (15, 6, 14) */,
  32'h3f242ada /* (11, 6, 14) */,
  32'h3f7ca6c7 /* (7, 6, 14) */,
  32'h3ed22ea6 /* (3, 6, 14) */,
  32'h3ec29928 /* (15, 2, 14) */,
  32'h3ea1d2a3 /* (11, 2, 14) */,
  32'h3ec56b70 /* (7, 2, 14) */,
  32'h3e9796af /* (3, 2, 14) */,
  32'h3eaab74a /* (15, 14, 10) */,
  32'h3f242ada /* (11, 14, 10) */,
  32'h3f7ca6c7 /* (7, 14, 10) */,
  32'h3ed22ea6 /* (3, 14, 10) */,
  32'h3f3f980b /* (15, 10, 10) */,
  32'h3fdbd2f0 /* (11, 10, 10) */,
  32'h4039abaa /* (7, 10, 10) */,
  32'h3f7e11f4 /* (3, 10, 10) */,
  32'h3f3f980b /* (15, 6, 10) */,
  32'h3fdbd2f0 /* (11, 6, 10) */,
  32'h4039abaa /* (7, 6, 10) */,
  32'h3f7e11f4 /* (3, 6, 10) */,
  32'h3eaab74a /* (15, 2, 10) */,
  32'h3f242ada /* (11, 2, 10) */,
  32'h3f7ca6c7 /* (7, 2, 10) */,
  32'h3ed22ea6 /* (3, 2, 10) */,
  32'h3eaab74a /* (15, 14, 6) */,
  32'h3f242ada /* (11, 14, 6) */,
  32'h3f7ca6c7 /* (7, 14, 6) */,
  32'h3ed22ea6 /* (3, 14, 6) */,
  32'h3f3f980b /* (15, 10, 6) */,
  32'h3fdbd2f0 /* (11, 10, 6) */,
  32'h4039abaa /* (7, 10, 6) */,
  32'h3f7e11f4 /* (3, 10, 6) */,
  32'h3f3f980b /* (15, 6, 6) */,
  32'h3fdbd2f0 /* (11, 6, 6) */,
  32'h4039abaa /* (7, 6, 6) */,
  32'h3f7e11f4 /* (3, 6, 6) */,
  32'h3eaab74a /* (15, 2, 6) */,
  32'h3f242ada /* (11, 2, 6) */,
  32'h3f7ca6c7 /* (7, 2, 6) */,
  32'h3ed22ea6 /* (3, 2, 6) */,
  32'h3ec29928 /* (15, 14, 2) */,
  32'h3ea1d2a3 /* (11, 14, 2) */,
  32'h3ec56b70 /* (7, 14, 2) */,
  32'h3e9796af /* (3, 14, 2) */,
  32'h3eaab74a /* (15, 10, 2) */,
  32'h3f242ada /* (11, 10, 2) */,
  32'h3f7ca6c7 /* (7, 10, 2) */,
  32'h3ed22ea6 /* (3, 10, 2) */,
  32'h3eaab74a /* (15, 6, 2) */,
  32'h3f242ada /* (11, 6, 2) */,
  32'h3f7ca6c7 /* (7, 6, 2) */,
  32'h3ed22ea6 /* (3, 6, 2) */,
  32'h3ec29928 /* (15, 2, 2) */,
  32'h3ea1d2a3 /* (11, 2, 2) */,
  32'h3ec56b70 /* (7, 2, 2) */,
  32'h3e9796af /* (3, 2, 2) */,
  32'h3ea8c974 /* (14, 14, 14) */,
  32'h3eb7f7fd /* (10, 14, 14) */,
  32'h3eb7f7fd /* (6, 14, 14) */,
  32'h3ea8c974 /* (2, 14, 14) */,
  32'h3eb7f7fd /* (14, 10, 14) */,
  32'h3f54d412 /* (10, 10, 14) */,
  32'h3f54d412 /* (6, 10, 14) */,
  32'h3eb7f7fd /* (2, 10, 14) */,
  32'h3eb7f7fd /* (14, 6, 14) */,
  32'h3f54d412 /* (10, 6, 14) */,
  32'h3f54d412 /* (6, 6, 14) */,
  32'h3eb7f7fd /* (2, 6, 14) */,
  32'h3ea8c974 /* (14, 2, 14) */,
  32'h3eb7f7fd /* (10, 2, 14) */,
  32'h3eb7f7fd /* (6, 2, 14) */,
  32'h3ea8c974 /* (2, 2, 14) */,
  32'h3eb7f7fd /* (14, 14, 10) */,
  32'h3f54d412 /* (10, 14, 10) */,
  32'h3f54d412 /* (6, 14, 10) */,
  32'h3eb7f7fd /* (2, 14, 10) */,
  32'h3f54d412 /* (14, 10, 10) */,
  32'h4015a2cf /* (10, 10, 10) */,
  32'h4015a2cf /* (6, 10, 10) */,
  32'h3f54d412 /* (2, 10, 10) */,
  32'h3f54d412 /* (14, 6, 10) */,
  32'h4015a2cf /* (10, 6, 10) */,
  32'h4015a2cf /* (6, 6, 10) */,
  32'h3f54d412 /* (2, 6, 10) */,
  32'h3eb7f7fd /* (14, 2, 10) */,
  32'h3f54d412 /* (10, 2, 10) */,
  32'h3f54d412 /* (6, 2, 10) */,
  32'h3eb7f7fd /* (2, 2, 10) */,
  32'h3eb7f7fd /* (14, 14, 6) */,
  32'h3f54d412 /* (10, 14, 6) */,
  32'h3f54d412 /* (6, 14, 6) */,
  32'h3eb7f7fd /* (2, 14, 6) */,
  32'h3f54d412 /* (14, 10, 6) */,
  32'h4015a2cf /* (10, 10, 6) */,
  32'h4015a2cf /* (6, 10, 6) */,
  32'h3f54d412 /* (2, 10, 6) */,
  32'h3f54d412 /* (14, 6, 6) */,
  32'h4015a2cf /* (10, 6, 6) */,
  32'h4015a2cf /* (6, 6, 6) */,
  32'h3f54d412 /* (2, 6, 6) */,
  32'h3eb7f7fd /* (14, 2, 6) */,
  32'h3f54d412 /* (10, 2, 6) */,
  32'h3f54d412 /* (6, 2, 6) */,
  32'h3eb7f7fd /* (2, 2, 6) */,
  32'h3ea8c974 /* (14, 14, 2) */,
  32'h3eb7f7fd /* (10, 14, 2) */,
  32'h3eb7f7fd /* (6, 14, 2) */,
  32'h3ea8c974 /* (2, 14, 2) */,
  32'h3eb7f7fd /* (14, 10, 2) */,
  32'h3f54d412 /* (10, 10, 2) */,
  32'h3f54d412 /* (6, 10, 2) */,
  32'h3eb7f7fd /* (2, 10, 2) */,
  32'h3eb7f7fd /* (14, 6, 2) */,
  32'h3f54d412 /* (10, 6, 2) */,
  32'h3f54d412 /* (6, 6, 2) */,
  32'h3eb7f7fd /* (2, 6, 2) */,
  32'h3ea8c974 /* (14, 2, 2) */,
  32'h3eb7f7fd /* (10, 2, 2) */,
  32'h3eb7f7fd /* (6, 2, 2) */,
  32'h3ea8c974 /* (2, 2, 2) */,
  32'h3e9796af /* (13, 14, 14) */,
  32'h3ec56b70 /* (9, 14, 14) */,
  32'h3ea1d2a3 /* (5, 14, 14) */,
  32'h3ec29928 /* (1, 14, 14) */,
  32'h3ed22ea6 /* (13, 10, 14) */,
  32'h3f7ca6c7 /* (9, 10, 14) */,
  32'h3f242ada /* (5, 10, 14) */,
  32'h3eaab74a /* (1, 10, 14) */,
  32'h3ed22ea6 /* (13, 6, 14) */,
  32'h3f7ca6c7 /* (9, 6, 14) */,
  32'h3f242ada /* (5, 6, 14) */,
  32'h3eaab74a /* (1, 6, 14) */,
  32'h3e9796af /* (13, 2, 14) */,
  32'h3ec56b70 /* (9, 2, 14) */,
  32'h3ea1d2a3 /* (5, 2, 14) */,
  32'h3ec29928 /* (1, 2, 14) */,
  32'h3ed22ea6 /* (13, 14, 10) */,
  32'h3f7ca6c7 /* (9, 14, 10) */,
  32'h3f242ada /* (5, 14, 10) */,
  32'h3eaab74a /* (1, 14, 10) */,
  32'h3f7e11f4 /* (13, 10, 10) */,
  32'h4039abaa /* (9, 10, 10) */,
  32'h3fdbd2f0 /* (5, 10, 10) */,
  32'h3f3f980b /* (1, 10, 10) */,
  32'h3f7e11f4 /* (13, 6, 10) */,
  32'h4039abaa /* (9, 6, 10) */,
  32'h3fdbd2f0 /* (5, 6, 10) */,
  32'h3f3f980b /* (1, 6, 10) */,
  32'h3ed22ea6 /* (13, 2, 10) */,
  32'h3f7ca6c7 /* (9, 2, 10) */,
  32'h3f242ada /* (5, 2, 10) */,
  32'h3eaab74a /* (1, 2, 10) */,
  32'h3ed22ea6 /* (13, 14, 6) */,
  32'h3f7ca6c7 /* (9, 14, 6) */,
  32'h3f242ada /* (5, 14, 6) */,
  32'h3eaab74a /* (1, 14, 6) */,
  32'h3f7e11f4 /* (13, 10, 6) */,
  32'h4039abaa /* (9, 10, 6) */,
  32'h3fdbd2f0 /* (5, 10, 6) */,
  32'h3f3f980b /* (1, 10, 6) */,
  32'h3f7e11f4 /* (13, 6, 6) */,
  32'h4039abaa /* (9, 6, 6) */,
  32'h3fdbd2f0 /* (5, 6, 6) */,
  32'h3f3f980b /* (1, 6, 6) */,
  32'h3ed22ea6 /* (13, 2, 6) */,
  32'h3f7ca6c7 /* (9, 2, 6) */,
  32'h3f242ada /* (5, 2, 6) */,
  32'h3eaab74a /* (1, 2, 6) */,
  32'h3e9796af /* (13, 14, 2) */,
  32'h3ec56b70 /* (9, 14, 2) */,
  32'h3ea1d2a3 /* (5, 14, 2) */,
  32'h3ec29928 /* (1, 14, 2) */,
  32'h3ed22ea6 /* (13, 10, 2) */,
  32'h3f7ca6c7 /* (9, 10, 2) */,
  32'h3f242ada /* (5, 10, 2) */,
  32'h3eaab74a /* (1, 10, 2) */,
  32'h3ed22ea6 /* (13, 6, 2) */,
  32'h3f7ca6c7 /* (9, 6, 2) */,
  32'h3f242ada /* (5, 6, 2) */,
  32'h3eaab74a /* (1, 6, 2) */,
  32'h3e9796af /* (13, 2, 2) */,
  32'h3ec56b70 /* (9, 2, 2) */,
  32'h3ea1d2a3 /* (5, 2, 2) */,
  32'h3ec29928 /* (1, 2, 2) */,
  32'h3e95577d /* (12, 14, 14) */,
  32'h3ead4da0 /* (8, 14, 14) */,
  32'h3e95577d /* (4, 14, 14) */,
  32'h3ed08e8d /* (0, 14, 14) */,
  32'h3effc9dc /* (12, 10, 14) */,
  32'h3f6fbf1e /* (8, 10, 14) */,
  32'h3effc9dc /* (4, 10, 14) */,
  32'h3ea6b2c0 /* (0, 10, 14) */,
  32'h3effc9dc /* (12, 6, 14) */,
  32'h3f6fbf1e /* (8, 6, 14) */,
  32'h3effc9dc /* (4, 6, 14) */,
  32'h3ea6b2c0 /* (0, 6, 14) */,
  32'h3e95577d /* (12, 2, 14) */,
  32'h3ead4da0 /* (8, 2, 14) */,
  32'h3e95577d /* (4, 2, 14) */,
  32'h3ed08e8d /* (0, 2, 14) */,
  32'h3effc9dc /* (12, 14, 10) */,
  32'h3f6fbf1e /* (8, 14, 10) */,
  32'h3effc9dc /* (4, 14, 10) */,
  32'h3ea6b2c0 /* (0, 14, 10) */,
  32'h3fa2a180 /* (12, 10, 10) */,
  32'h40372c7f /* (8, 10, 10) */,
  32'h3fa2a180 /* (4, 10, 10) */,
  32'h3f390e8b /* (0, 10, 10) */,
  32'h3fa2a180 /* (12, 6, 10) */,
  32'h40372c7f /* (8, 6, 10) */,
  32'h3fa2a180 /* (4, 6, 10) */,
  32'h3f390e8b /* (0, 6, 10) */,
  32'h3effc9dc /* (12, 2, 10) */,
  32'h3f6fbf1e /* (8, 2, 10) */,
  32'h3effc9dc /* (4, 2, 10) */,
  32'h3ea6b2c0 /* (0, 2, 10) */,
  32'h3effc9dc /* (12, 14, 6) */,
  32'h3f6fbf1e /* (8, 14, 6) */,
  32'h3effc9dc /* (4, 14, 6) */,
  32'h3ea6b2c0 /* (0, 14, 6) */,
  32'h3fa2a180 /* (12, 10, 6) */,
  32'h40372c7f /* (8, 10, 6) */,
  32'h3fa2a180 /* (4, 10, 6) */,
  32'h3f390e8b /* (0, 10, 6) */,
  32'h3fa2a180 /* (12, 6, 6) */,
  32'h40372c7f /* (8, 6, 6) */,
  32'h3fa2a180 /* (4, 6, 6) */,
  32'h3f390e8b /* (0, 6, 6) */,
  32'h3effc9dc /* (12, 2, 6) */,
  32'h3f6fbf1e /* (8, 2, 6) */,
  32'h3effc9dc /* (4, 2, 6) */,
  32'h3ea6b2c0 /* (0, 2, 6) */,
  32'h3e95577d /* (12, 14, 2) */,
  32'h3ead4da0 /* (8, 14, 2) */,
  32'h3e95577d /* (4, 14, 2) */,
  32'h3ed08e8d /* (0, 14, 2) */,
  32'h3effc9dc /* (12, 10, 2) */,
  32'h3f6fbf1e /* (8, 10, 2) */,
  32'h3effc9dc /* (4, 10, 2) */,
  32'h3ea6b2c0 /* (0, 10, 2) */,
  32'h3effc9dc /* (12, 6, 2) */,
  32'h3f6fbf1e /* (8, 6, 2) */,
  32'h3effc9dc /* (4, 6, 2) */,
  32'h3ea6b2c0 /* (0, 6, 2) */,
  32'h3e95577d /* (12, 2, 2) */,
  32'h3ead4da0 /* (8, 2, 2) */,
  32'h3e95577d /* (4, 2, 2) */,
  32'h3ed08e8d /* (0, 2, 2) */,
  32'h3e9f2a5d /* (15, 13, 14) */,
  32'h3eb2cc97 /* (11, 13, 14) */,
  32'h3ee6ec8a /* (7, 13, 14) */,
  32'h3e9508f6 /* (3, 13, 14) */,
  32'h3eb430e1 /* (15, 9, 14) */,
  32'h3f3e2f24 /* (11, 9, 14) */,
  32'h3f993b79 /* (7, 9, 14) */,
  32'h3ee6ec8a /* (3, 9, 14) */,
  32'h3e99eb68 /* (15, 5, 14) */,
  32'h3f025da2 /* (11, 5, 14) */,
  32'h3f3e2f24 /* (7, 5, 14) */,
  32'h3eb2cc97 /* (3, 5, 14) */,
  32'h3efc66bd /* (15, 1, 14) */,
  32'h3e99eb68 /* (11, 1, 14) */,
  32'h3eb430e1 /* (7, 1, 14) */,
  32'h3e9f2a5d /* (3, 1, 14) */,
  32'h3ec1987e /* (15, 13, 10) */,
  32'h3f41f419 /* (11, 13, 10) */,
  32'h3f982d5a /* (7, 13, 10) */,
  32'h3ef2a853 /* (3, 13, 10) */,
  32'h3f62162b /* (15, 9, 10) */,
  32'h4006bd24 /* (11, 9, 10) */,
  32'h406912bc /* (7, 9, 10) */,
  32'h3f982d5a /* (3, 9, 10) */,
  32'h3f14d2ae /* (15, 5, 10) */,
  32'h3fa39217 /* (11, 5, 10) */,
  32'h4006bd24 /* (7, 5, 10) */,
  32'h3f41f419 /* (3, 5, 10) */,
  32'h3e9f454b /* (15, 1, 10) */,
  32'h3f14d2ae /* (11, 1, 10) */,
  32'h3f62162b /* (7, 1, 10) */,
  32'h3ec1987e /* (3, 1, 10) */,
  32'h3ec1987e /* (15, 13, 6) */,
  32'h3f41f419 /* (11, 13, 6) */,
  32'h3f982d5a /* (7, 13, 6) */,
  32'h3ef2a853 /* (3, 13, 6) */,
  32'h3f62162b /* (15, 9, 6) */,
  32'h4006bd24 /* (11, 9, 6) */,
  32'h406912bc /* (7, 9, 6) */,
  32'h3f982d5a /* (3, 9, 6) */,
  32'h3f14d2ae /* (15, 5, 6) */,
  32'h3fa39217 /* (11, 5, 6) */,
  32'h4006bd24 /* (7, 5, 6) */,
  32'h3f41f419 /* (3, 5, 6) */,
  32'h3e9f454b /* (15, 1, 6) */,
  32'h3f14d2ae /* (11, 1, 6) */,
  32'h3f62162b /* (7, 1, 6) */,
  32'h3ec1987e /* (3, 1, 6) */,
  32'h3e9f2a5d /* (15, 13, 2) */,
  32'h3eb2cc97 /* (11, 13, 2) */,
  32'h3ee6ec8a /* (7, 13, 2) */,
  32'h3e9508f6 /* (3, 13, 2) */,
  32'h3eb430e1 /* (15, 9, 2) */,
  32'h3f3e2f24 /* (11, 9, 2) */,
  32'h3f993b79 /* (7, 9, 2) */,
  32'h3ee6ec8a /* (3, 9, 2) */,
  32'h3e99eb68 /* (15, 5, 2) */,
  32'h3f025da2 /* (11, 5, 2) */,
  32'h3f3e2f24 /* (7, 5, 2) */,
  32'h3eb2cc97 /* (3, 5, 2) */,
  32'h3efc66bd /* (15, 1, 2) */,
  32'h3e99eb68 /* (11, 1, 2) */,
  32'h3eb430e1 /* (7, 1, 2) */,
  32'h3e9f2a5d /* (3, 1, 2) */,
  32'h3e9796af /* (14, 13, 14) */,
  32'h3ed22ea6 /* (10, 13, 14) */,
  32'h3ed22ea6 /* (6, 13, 14) */,
  32'h3e9796af /* (2, 13, 14) */,
  32'h3ec56b70 /* (14, 9, 14) */,
  32'h3f7ca6c7 /* (10, 9, 14) */,
  32'h3f7ca6c7 /* (6, 9, 14) */,
  32'h3ec56b70 /* (2, 9, 14) */,
  32'h3ea1d2a3 /* (14, 5, 14) */,
  32'h3f242ada /* (10, 5, 14) */,
  32'h3f242ada /* (6, 5, 14) */,
  32'h3ea1d2a3 /* (2, 5, 14) */,
  32'h3ec29928 /* (14, 1, 14) */,
  32'h3eaab74a /* (10, 1, 14) */,
  32'h3eaab74a /* (6, 1, 14) */,
  32'h3ec29928 /* (2, 1, 14) */,
  32'h3ed22ea6 /* (14, 13, 10) */,
  32'h3f7e11f4 /* (10, 13, 10) */,
  32'h3f7e11f4 /* (6, 13, 10) */,
  32'h3ed22ea6 /* (2, 13, 10) */,
  32'h3f7ca6c7 /* (14, 9, 10) */,
  32'h4039abaa /* (10, 9, 10) */,
  32'h4039abaa /* (6, 9, 10) */,
  32'h3f7ca6c7 /* (2, 9, 10) */,
  32'h3f242ada /* (14, 5, 10) */,
  32'h3fdbd2f0 /* (10, 5, 10) */,
  32'h3fdbd2f0 /* (6, 5, 10) */,
  32'h3f242ada /* (2, 5, 10) */,
  32'h3eaab74a /* (14, 1, 10) */,
  32'h3f3f980b /* (10, 1, 10) */,
  32'h3f3f980b /* (6, 1, 10) */,
  32'h3eaab74a /* (2, 1, 10) */,
  32'h3ed22ea6 /* (14, 13, 6) */,
  32'h3f7e11f4 /* (10, 13, 6) */,
  32'h3f7e11f4 /* (6, 13, 6) */,
  32'h3ed22ea6 /* (2, 13, 6) */,
  32'h3f7ca6c7 /* (14, 9, 6) */,
  32'h4039abaa /* (10, 9, 6) */,
  32'h4039abaa /* (6, 9, 6) */,
  32'h3f7ca6c7 /* (2, 9, 6) */,
  32'h3f242ada /* (14, 5, 6) */,
  32'h3fdbd2f0 /* (10, 5, 6) */,
  32'h3fdbd2f0 /* (6, 5, 6) */,
  32'h3f242ada /* (2, 5, 6) */,
  32'h3eaab74a /* (14, 1, 6) */,
  32'h3f3f980b /* (10, 1, 6) */,
  32'h3f3f980b /* (6, 1, 6) */,
  32'h3eaab74a /* (2, 1, 6) */,
  32'h3e9796af /* (14, 13, 2) */,
  32'h3ed22ea6 /* (10, 13, 2) */,
  32'h3ed22ea6 /* (6, 13, 2) */,
  32'h3e9796af /* (2, 13, 2) */,
  32'h3ec56b70 /* (14, 9, 2) */,
  32'h3f7ca6c7 /* (10, 9, 2) */,
  32'h3f7ca6c7 /* (6, 9, 2) */,
  32'h3ec56b70 /* (2, 9, 2) */,
  32'h3ea1d2a3 /* (14, 5, 2) */,
  32'h3f242ada /* (10, 5, 2) */,
  32'h3f242ada /* (6, 5, 2) */,
  32'h3ea1d2a3 /* (2, 5, 2) */,
  32'h3ec29928 /* (14, 1, 2) */,
  32'h3eaab74a /* (10, 1, 2) */,
  32'h3eaab74a /* (6, 1, 2) */,
  32'h3ec29928 /* (2, 1, 2) */,
  32'h3e9508f6 /* (13, 13, 14) */,
  32'h3ee6ec8a /* (9, 13, 14) */,
  32'h3eb2cc97 /* (5, 13, 14) */,
  32'h3e9f2a5d /* (1, 13, 14) */,
  32'h3ee6ec8a /* (13, 9, 14) */,
  32'h3f993b79 /* (9, 9, 14) */,
  32'h3f3e2f24 /* (5, 9, 14) */,
  32'h3eb430e1 /* (1, 9, 14) */,
  32'h3eb2cc97 /* (13, 5, 14) */,
  32'h3f3e2f24 /* (9, 5, 14) */,
  32'h3f025da2 /* (5, 5, 14) */,
  32'h3e99eb68 /* (1, 5, 14) */,
  32'h3e9f2a5d /* (13, 1, 14) */,
  32'h3eb430e1 /* (9, 1, 14) */,
  32'h3e99eb68 /* (5, 1, 14) */,
  32'h3efc66bd /* (1, 1, 14) */,
  32'h3ef2a853 /* (13, 13, 10) */,
  32'h3f982d5a /* (9, 13, 10) */,
  32'h3f41f419 /* (5, 13, 10) */,
  32'h3ec1987e /* (1, 13, 10) */,
  32'h3f982d5a /* (13, 9, 10) */,
  32'h406912bc /* (9, 9, 10) */,
  32'h4006bd24 /* (5, 9, 10) */,
  32'h3f62162b /* (1, 9, 10) */,
  32'h3f41f419 /* (13, 5, 10) */,
  32'h4006bd24 /* (9, 5, 10) */,
  32'h3fa39217 /* (5, 5, 10) */,
  32'h3f14d2ae /* (1, 5, 10) */,
  32'h3ec1987e /* (13, 1, 10) */,
  32'h3f62162b /* (9, 1, 10) */,
  32'h3f14d2ae /* (5, 1, 10) */,
  32'h3e9f454b /* (1, 1, 10) */,
  32'h3ef2a853 /* (13, 13, 6) */,
  32'h3f982d5a /* (9, 13, 6) */,
  32'h3f41f419 /* (5, 13, 6) */,
  32'h3ec1987e /* (1, 13, 6) */,
  32'h3f982d5a /* (13, 9, 6) */,
  32'h406912bc /* (9, 9, 6) */,
  32'h4006bd24 /* (5, 9, 6) */,
  32'h3f62162b /* (1, 9, 6) */,
  32'h3f41f419 /* (13, 5, 6) */,
  32'h4006bd24 /* (9, 5, 6) */,
  32'h3fa39217 /* (5, 5, 6) */,
  32'h3f14d2ae /* (1, 5, 6) */,
  32'h3ec1987e /* (13, 1, 6) */,
  32'h3f62162b /* (9, 1, 6) */,
  32'h3f14d2ae /* (5, 1, 6) */,
  32'h3e9f454b /* (1, 1, 6) */,
  32'h3e9508f6 /* (13, 13, 2) */,
  32'h3ee6ec8a /* (9, 13, 2) */,
  32'h3eb2cc97 /* (5, 13, 2) */,
  32'h3e9f2a5d /* (1, 13, 2) */,
  32'h3ee6ec8a /* (13, 9, 2) */,
  32'h3f993b79 /* (9, 9, 2) */,
  32'h3f3e2f24 /* (5, 9, 2) */,
  32'h3eb430e1 /* (1, 9, 2) */,
  32'h3eb2cc97 /* (13, 5, 2) */,
  32'h3f3e2f24 /* (9, 5, 2) */,
  32'h3f025da2 /* (5, 5, 2) */,
  32'h3e99eb68 /* (1, 5, 2) */,
  32'h3e9f2a5d /* (13, 1, 2) */,
  32'h3eb430e1 /* (9, 1, 2) */,
  32'h3e99eb68 /* (5, 1, 2) */,
  32'h3efc66bd /* (1, 1, 2) */,
  32'h3e9d3fef /* (12, 13, 14) */,
  32'h3ece2dc1 /* (8, 13, 14) */,
  32'h3e9d3fef /* (4, 13, 14) */,
  32'h3ea34ae8 /* (0, 13, 14) */,
  32'h3f104c25 /* (12, 9, 14) */,
  32'h3f9420e3 /* (8, 9, 14) */,
  32'h3f104c25 /* (4, 9, 14) */,
  32'h3eaee5c8 /* (0, 9, 14) */,
  32'h3ed1ff4c /* (12, 5, 14) */,
  32'h3f30df4f /* (8, 5, 14) */,
  32'h3ed1ff4c /* (4, 5, 14) */,
  32'h3e97b006 /* (0, 5, 14) */,
  32'h3e939519 /* (12, 1, 14) */,
  32'h3e9c5e8a /* (8, 1, 14) */,
  32'h3e939519 /* (4, 1, 14) */,
  32'h3f10451b /* (0, 1, 14) */,
  32'h3f15625b /* (12, 13, 10) */,
  32'h3f91854a /* (8, 13, 10) */,
  32'h3f15625b /* (4, 13, 10) */,
  32'h3ebc86f4 /* (0, 13, 10) */,
  32'h3fc4fc22 /* (12, 9, 10) */,
  32'h40686d0d /* (8, 9, 10) */,
  32'h3fc4fc22 /* (4, 9, 10) */,
  32'h3f59ea43 /* (0, 9, 10) */,
  32'h3f753c17 /* (12, 5, 10) */,
  32'h40037a14 /* (8, 5, 10) */,
  32'h3f753c17 /* (4, 5, 10) */,
  32'h3f1019ab /* (0, 5, 10) */,
  32'h3ee9b2a2 /* (12, 1, 10) */,
  32'h3f5576ec /* (8, 1, 10) */,
  32'h3ee9b2a2 /* (4, 1, 10) */,
  32'h3e9bd472 /* (0, 1, 10) */,
  32'h3f15625b /* (12, 13, 6) */,
  32'h3f91854a /* (8, 13, 6) */,
  32'h3f15625b /* (4, 13, 6) */,
  32'h3ebc86f4 /* (0, 13, 6) */,
  32'h3fc4fc22 /* (12, 9, 6) */,
  32'h40686d0d /* (8, 9, 6) */,
  32'h3fc4fc22 /* (4, 9, 6) */,
  32'h3f59ea43 /* (0, 9, 6) */,
  32'h3f753c17 /* (12, 5, 6) */,
  32'h40037a14 /* (8, 5, 6) */,
  32'h3f753c17 /* (4, 5, 6) */,
  32'h3f1019ab /* (0, 5, 6) */,
  32'h3ee9b2a2 /* (12, 1, 6) */,
  32'h3f5576ec /* (8, 1, 6) */,
  32'h3ee9b2a2 /* (4, 1, 6) */,
  32'h3e9bd472 /* (0, 1, 6) */,
  32'h3e9d3fef /* (12, 13, 2) */,
  32'h3ece2dc1 /* (8, 13, 2) */,
  32'h3e9d3fef /* (4, 13, 2) */,
  32'h3ea34ae8 /* (0, 13, 2) */,
  32'h3f104c25 /* (12, 9, 2) */,
  32'h3f9420e3 /* (8, 9, 2) */,
  32'h3f104c25 /* (4, 9, 2) */,
  32'h3eaee5c8 /* (0, 9, 2) */,
  32'h3ed1ff4c /* (12, 5, 2) */,
  32'h3f30df4f /* (8, 5, 2) */,
  32'h3ed1ff4c /* (4, 5, 2) */,
  32'h3e97b006 /* (0, 5, 2) */,
  32'h3e939519 /* (12, 1, 2) */,
  32'h3e9c5e8a /* (8, 1, 2) */,
  32'h3e939519 /* (4, 1, 2) */,
  32'h3f10451b /* (0, 1, 2) */,
  32'h3e939519 /* (15, 12, 14) */,
  32'h3ed1ff4c /* (11, 12, 14) */,
  32'h3f104c25 /* (7, 12, 14) */,
  32'h3e9d3fef /* (3, 12, 14) */,
  32'h3e9c5e8a /* (15, 8, 14) */,
  32'h3f30df4f /* (11, 8, 14) */,
  32'h3f9420e3 /* (7, 8, 14) */,
  32'h3ece2dc1 /* (3, 8, 14) */,
  32'h3e939519 /* (15, 4, 14) */,
  32'h3ed1ff4c /* (11, 4, 14) */,
  32'h3f104c25 /* (7, 4, 14) */,
  32'h3e9d3fef /* (3, 4, 14) */,
  32'h3f10451b /* (15, 0, 14) */,
  32'h3e97b006 /* (11, 0, 14) */,
  32'h3eaee5c8 /* (7, 0, 14) */,
  32'h3ea34ae8 /* (3, 0, 14) */,
  32'h3ee9b2a2 /* (15, 12, 10) */,
  32'h3f753c17 /* (11, 12, 10) */,
  32'h3fc4fc22 /* (7, 12, 10) */,
  32'h3f15625b /* (3, 12, 10) */,
  32'h3f5576ec /* (15, 8, 10) */,
  32'h40037a14 /* (11, 8, 10) */,
  32'h40686d0d /* (7, 8, 10) */,
  32'h3f91854a /* (3, 8, 10) */,
  32'h3ee9b2a2 /* (15, 4, 10) */,
  32'h3f753c17 /* (11, 4, 10) */,
  32'h3fc4fc22 /* (7, 4, 10) */,
  32'h3f15625b /* (3, 4, 10) */,
  32'h3e9bd472 /* (15, 0, 10) */,
  32'h3f1019ab /* (11, 0, 10) */,
  32'h3f59ea43 /* (7, 0, 10) */,
  32'h3ebc86f4 /* (3, 0, 10) */,
  32'h3ee9b2a2 /* (15, 12, 6) */,
  32'h3f753c17 /* (11, 12, 6) */,
  32'h3fc4fc22 /* (7, 12, 6) */,
  32'h3f15625b /* (3, 12, 6) */,
  32'h3f5576ec /* (15, 8, 6) */,
  32'h40037a14 /* (11, 8, 6) */,
  32'h40686d0d /* (7, 8, 6) */,
  32'h3f91854a /* (3, 8, 6) */,
  32'h3ee9b2a2 /* (15, 4, 6) */,
  32'h3f753c17 /* (11, 4, 6) */,
  32'h3fc4fc22 /* (7, 4, 6) */,
  32'h3f15625b /* (3, 4, 6) */,
  32'h3e9bd472 /* (15, 0, 6) */,
  32'h3f1019ab /* (11, 0, 6) */,
  32'h3f59ea43 /* (7, 0, 6) */,
  32'h3ebc86f4 /* (3, 0, 6) */,
  32'h3e939519 /* (15, 12, 2) */,
  32'h3ed1ff4c /* (11, 12, 2) */,
  32'h3f104c25 /* (7, 12, 2) */,
  32'h3e9d3fef /* (3, 12, 2) */,
  32'h3e9c5e8a /* (15, 8, 2) */,
  32'h3f30df4f /* (11, 8, 2) */,
  32'h3f9420e3 /* (7, 8, 2) */,
  32'h3ece2dc1 /* (3, 8, 2) */,
  32'h3e939519 /* (15, 4, 2) */,
  32'h3ed1ff4c /* (11, 4, 2) */,
  32'h3f104c25 /* (7, 4, 2) */,
  32'h3e9d3fef /* (3, 4, 2) */,
  32'h3f10451b /* (15, 0, 2) */,
  32'h3e97b006 /* (11, 0, 2) */,
  32'h3eaee5c8 /* (7, 0, 2) */,
  32'h3ea34ae8 /* (3, 0, 2) */,
  32'h3e95577d /* (14, 12, 14) */,
  32'h3effc9dc /* (10, 12, 14) */,
  32'h3effc9dc /* (6, 12, 14) */,
  32'h3e95577d /* (2, 12, 14) */,
  32'h3ead4da0 /* (14, 8, 14) */,
  32'h3f6fbf1e /* (10, 8, 14) */,
  32'h3f6fbf1e /* (6, 8, 14) */,
  32'h3ead4da0 /* (2, 8, 14) */,
  32'h3e95577d /* (14, 4, 14) */,
  32'h3effc9dc /* (10, 4, 14) */,
  32'h3effc9dc /* (6, 4, 14) */,
  32'h3e95577d /* (2, 4, 14) */,
  32'h3ed08e8d /* (14, 0, 14) */,
  32'h3ea6b2c0 /* (10, 0, 14) */,
  32'h3ea6b2c0 /* (6, 0, 14) */,
  32'h3ed08e8d /* (2, 0, 14) */,
  32'h3effc9dc /* (14, 12, 10) */,
  32'h3fa2a180 /* (10, 12, 10) */,
  32'h3fa2a180 /* (6, 12, 10) */,
  32'h3effc9dc /* (2, 12, 10) */,
  32'h3f6fbf1e /* (14, 8, 10) */,
  32'h40372c7f /* (10, 8, 10) */,
  32'h40372c7f /* (6, 8, 10) */,
  32'h3f6fbf1e /* (2, 8, 10) */,
  32'h3effc9dc /* (14, 4, 10) */,
  32'h3fa2a180 /* (10, 4, 10) */,
  32'h3fa2a180 /* (6, 4, 10) */,
  32'h3effc9dc /* (2, 4, 10) */,
  32'h3ea6b2c0 /* (14, 0, 10) */,
  32'h3f390e8b /* (10, 0, 10) */,
  32'h3f390e8b /* (6, 0, 10) */,
  32'h3ea6b2c0 /* (2, 0, 10) */,
  32'h3effc9dc /* (14, 12, 6) */,
  32'h3fa2a180 /* (10, 12, 6) */,
  32'h3fa2a180 /* (6, 12, 6) */,
  32'h3effc9dc /* (2, 12, 6) */,
  32'h3f6fbf1e /* (14, 8, 6) */,
  32'h40372c7f /* (10, 8, 6) */,
  32'h40372c7f /* (6, 8, 6) */,
  32'h3f6fbf1e /* (2, 8, 6) */,
  32'h3effc9dc /* (14, 4, 6) */,
  32'h3fa2a180 /* (10, 4, 6) */,
  32'h3fa2a180 /* (6, 4, 6) */,
  32'h3effc9dc /* (2, 4, 6) */,
  32'h3ea6b2c0 /* (14, 0, 6) */,
  32'h3f390e8b /* (10, 0, 6) */,
  32'h3f390e8b /* (6, 0, 6) */,
  32'h3ea6b2c0 /* (2, 0, 6) */,
  32'h3e95577d /* (14, 12, 2) */,
  32'h3effc9dc /* (10, 12, 2) */,
  32'h3effc9dc /* (6, 12, 2) */,
  32'h3e95577d /* (2, 12, 2) */,
  32'h3ead4da0 /* (14, 8, 2) */,
  32'h3f6fbf1e /* (10, 8, 2) */,
  32'h3f6fbf1e /* (6, 8, 2) */,
  32'h3ead4da0 /* (2, 8, 2) */,
  32'h3e95577d /* (14, 4, 2) */,
  32'h3effc9dc /* (10, 4, 2) */,
  32'h3effc9dc /* (6, 4, 2) */,
  32'h3e95577d /* (2, 4, 2) */,
  32'h3ed08e8d /* (14, 0, 2) */,
  32'h3ea6b2c0 /* (10, 0, 2) */,
  32'h3ea6b2c0 /* (6, 0, 2) */,
  32'h3ed08e8d /* (2, 0, 2) */,
  32'h3e9d3fef /* (13, 12, 14) */,
  32'h3f104c25 /* (9, 12, 14) */,
  32'h3ed1ff4c /* (5, 12, 14) */,
  32'h3e939519 /* (1, 12, 14) */,
  32'h3ece2dc1 /* (13, 8, 14) */,
  32'h3f9420e3 /* (9, 8, 14) */,
  32'h3f30df4f /* (5, 8, 14) */,
  32'h3e9c5e8a /* (1, 8, 14) */,
  32'h3e9d3fef /* (13, 4, 14) */,
  32'h3f104c25 /* (9, 4, 14) */,
  32'h3ed1ff4c /* (5, 4, 14) */,
  32'h3e939519 /* (1, 4, 14) */,
  32'h3ea34ae8 /* (13, 0, 14) */,
  32'h3eaee5c8 /* (9, 0, 14) */,
  32'h3e97b006 /* (5, 0, 14) */,
  32'h3f10451b /* (1, 0, 14) */,
  32'h3f15625b /* (13, 12, 10) */,
  32'h3fc4fc22 /* (9, 12, 10) */,
  32'h3f753c17 /* (5, 12, 10) */,
  32'h3ee9b2a2 /* (1, 12, 10) */,
  32'h3f91854a /* (13, 8, 10) */,
  32'h40686d0d /* (9, 8, 10) */,
  32'h40037a14 /* (5, 8, 10) */,
  32'h3f5576ec /* (1, 8, 10) */,
  32'h3f15625b /* (13, 4, 10) */,
  32'h3fc4fc22 /* (9, 4, 10) */,
  32'h3f753c17 /* (5, 4, 10) */,
  32'h3ee9b2a2 /* (1, 4, 10) */,
  32'h3ebc86f4 /* (13, 0, 10) */,
  32'h3f59ea43 /* (9, 0, 10) */,
  32'h3f1019ab /* (5, 0, 10) */,
  32'h3e9bd472 /* (1, 0, 10) */,
  32'h3f15625b /* (13, 12, 6) */,
  32'h3fc4fc22 /* (9, 12, 6) */,
  32'h3f753c17 /* (5, 12, 6) */,
  32'h3ee9b2a2 /* (1, 12, 6) */,
  32'h3f91854a /* (13, 8, 6) */,
  32'h40686d0d /* (9, 8, 6) */,
  32'h40037a14 /* (5, 8, 6) */,
  32'h3f5576ec /* (1, 8, 6) */,
  32'h3f15625b /* (13, 4, 6) */,
  32'h3fc4fc22 /* (9, 4, 6) */,
  32'h3f753c17 /* (5, 4, 6) */,
  32'h3ee9b2a2 /* (1, 4, 6) */,
  32'h3ebc86f4 /* (13, 0, 6) */,
  32'h3f59ea43 /* (9, 0, 6) */,
  32'h3f1019ab /* (5, 0, 6) */,
  32'h3e9bd472 /* (1, 0, 6) */,
  32'h3e9d3fef /* (13, 12, 2) */,
  32'h3f104c25 /* (9, 12, 2) */,
  32'h3ed1ff4c /* (5, 12, 2) */,
  32'h3e939519 /* (1, 12, 2) */,
  32'h3ece2dc1 /* (13, 8, 2) */,
  32'h3f9420e3 /* (9, 8, 2) */,
  32'h3f30df4f /* (5, 8, 2) */,
  32'h3e9c5e8a /* (1, 8, 2) */,
  32'h3e9d3fef /* (13, 4, 2) */,
  32'h3f104c25 /* (9, 4, 2) */,
  32'h3ed1ff4c /* (5, 4, 2) */,
  32'h3e939519 /* (1, 4, 2) */,
  32'h3ea34ae8 /* (13, 0, 2) */,
  32'h3eaee5c8 /* (9, 0, 2) */,
  32'h3e97b006 /* (5, 0, 2) */,
  32'h3f10451b /* (1, 0, 2) */,
  32'h3eb02eb0 /* (12, 12, 14) */,
  32'h3f036eaf /* (8, 12, 14) */,
  32'h3eb02eb0 /* (4, 12, 14) */,
  32'h3e939fbd /* (0, 12, 14) */,
  32'h3f036eaf /* (12, 8, 14) */,
  32'h3f91966b /* (8, 8, 14) */,
  32'h3f036eaf /* (4, 8, 14) */,
  32'h3e9727de /* (0, 8, 14) */,
  32'h3eb02eb0 /* (12, 4, 14) */,
  32'h3f036eaf /* (8, 4, 14) */,
  32'h3eb02eb0 /* (4, 4, 14) */,
  32'h3e939fbd /* (0, 4, 14) */,
  32'h3e939fbd /* (12, 0, 14) */,
  32'h3e9727de /* (8, 0, 14) */,
  32'h3e939fbd /* (4, 0, 14) */,
  32'h3f2bcc5c /* (0, 0, 14) */,
  32'h3f3a61a4 /* (12, 12, 10) */,
  32'h3fbe2ead /* (8, 12, 10) */,
  32'h3f3a61a4 /* (4, 12, 10) */,
  32'h3ee2e9d3 /* (0, 12, 10) */,
  32'h3fbe2ead /* (12, 8, 10) */,
  32'h406a2757 /* (8, 8, 10) */,
  32'h3fbe2ead /* (4, 8, 10) */,
  32'h3f4d63f0 /* (0, 8, 10) */,
  32'h3f3a61a4 /* (12, 4, 10) */,
  32'h3fbe2ead /* (8, 4, 10) */,
  32'h3f3a61a4 /* (4, 4, 10) */,
  32'h3ee2e9d3 /* (0, 4, 10) */,
  32'h3ee2e9d3 /* (12, 0, 10) */,
  32'h3f4d63f0 /* (8, 0, 10) */,
  32'h3ee2e9d3 /* (4, 0, 10) */,
  32'h3e989327 /* (0, 0, 10) */,
  32'h3f3a61a4 /* (12, 12, 6) */,
  32'h3fbe2ead /* (8, 12, 6) */,
  32'h3f3a61a4 /* (4, 12, 6) */,
  32'h3ee2e9d3 /* (0, 12, 6) */,
  32'h3fbe2ead /* (12, 8, 6) */,
  32'h406a2757 /* (8, 8, 6) */,
  32'h3fbe2ead /* (4, 8, 6) */,
  32'h3f4d63f0 /* (0, 8, 6) */,
  32'h3f3a61a4 /* (12, 4, 6) */,
  32'h3fbe2ead /* (8, 4, 6) */,
  32'h3f3a61a4 /* (4, 4, 6) */,
  32'h3ee2e9d3 /* (0, 4, 6) */,
  32'h3ee2e9d3 /* (12, 0, 6) */,
  32'h3f4d63f0 /* (8, 0, 6) */,
  32'h3ee2e9d3 /* (4, 0, 6) */,
  32'h3e989327 /* (0, 0, 6) */,
  32'h3eb02eb0 /* (12, 12, 2) */,
  32'h3f036eaf /* (8, 12, 2) */,
  32'h3eb02eb0 /* (4, 12, 2) */,
  32'h3e939fbd /* (0, 12, 2) */,
  32'h3f036eaf /* (12, 8, 2) */,
  32'h3f91966b /* (8, 8, 2) */,
  32'h3f036eaf /* (4, 8, 2) */,
  32'h3e9727de /* (0, 8, 2) */,
  32'h3eb02eb0 /* (12, 4, 2) */,
  32'h3f036eaf /* (8, 4, 2) */,
  32'h3eb02eb0 /* (4, 4, 2) */,
  32'h3e939fbd /* (0, 4, 2) */,
  32'h3e939fbd /* (12, 0, 2) */,
  32'h3e9727de /* (8, 0, 2) */,
  32'h3e939fbd /* (4, 0, 2) */,
  32'h3f2bcc5c /* (0, 0, 2) */,
  32'h3eaf2a10 /* (15, 15, 13) */,
  32'h3ea7dbb1 /* (11, 15, 13) */,
  32'h3ed1d4cb /* (7, 15, 13) */,
  32'h3e953797 /* (3, 15, 13) */,
  32'h3ea7dbb1 /* (15, 11, 13) */,
  32'h3f17cf64 /* (11, 11, 13) */,
  32'h3f6365d6 /* (7, 11, 13) */,
  32'h3ec9097c /* (3, 11, 13) */,
  32'h3ed1d4cb /* (15, 7, 13) */,
  32'h3f6365d6 /* (11, 7, 13) */,
  32'h3fb9d98f /* (7, 7, 13) */,
  32'h3f07f0f8 /* (3, 7, 13) */,
  32'h3e953797 /* (15, 3, 13) */,
  32'h3ec9097c /* (11, 3, 13) */,
  32'h3f07f0f8 /* (7, 3, 13) */,
  32'h3e9a814a /* (3, 3, 13) */,
  32'h3ea4f994 /* (15, 15, 9) */,
  32'h3f2b075a /* (11, 15, 9) */,
  32'h3f88838c /* (7, 15, 9) */,
  32'h3ed1d4cb /* (3, 15, 9) */,
  32'h3f2b075a /* (15, 11, 9) */,
  32'h3fc5882d /* (11, 11, 9) */,
  32'h40278361 /* (7, 11, 9) */,
  32'h3f6365d6 /* (3, 11, 9) */,
  32'h3f88838c /* (15, 7, 9) */,
  32'h40278361 /* (11, 7, 9) */,
  32'h4093adcc /* (7, 7, 9) */,
  32'h3fb9d98f /* (3, 7, 9) */,
  32'h3ed1d4cb /* (15, 3, 9) */,
  32'h3f6365d6 /* (11, 3, 9) */,
  32'h3fb9d98f /* (7, 3, 9) */,
  32'h3f07f0f8 /* (3, 3, 9) */,
  32'h3e93e191 /* (15, 15, 5) */,
  32'h3eeeb6df /* (11, 15, 5) */,
  32'h3f2b075a /* (7, 15, 5) */,
  32'h3ea7dbb1 /* (3, 15, 5) */,
  32'h3eeeb6df /* (15, 11, 5) */,
  32'h3f77795a /* (11, 11, 5) */,
  32'h3fc5882d /* (7, 11, 5) */,
  32'h3f17cf64 /* (3, 11, 5) */,
  32'h3f2b075a /* (15, 7, 5) */,
  32'h3fc5882d /* (11, 7, 5) */,
  32'h40278361 /* (7, 7, 5) */,
  32'h3f6365d6 /* (3, 7, 5) */,
  32'h3ea7dbb1 /* (15, 3, 5) */,
  32'h3f17cf64 /* (11, 3, 5) */,
  32'h3f6365d6 /* (7, 3, 5) */,
  32'h3ec9097c /* (3, 3, 5) */,
  32'h3f5a3fd8 /* (15, 15, 1) */,
  32'h3e93e191 /* (11, 15, 1) */,
  32'h3ea4f994 /* (7, 15, 1) */,
  32'h3eaf2a10 /* (3, 15, 1) */,
  32'h3e93e191 /* (15, 11, 1) */,
  32'h3eeeb6df /* (11, 11, 1) */,
  32'h3f2b075a /* (7, 11, 1) */,
  32'h3ea7dbb1 /* (3, 11, 1) */,
  32'h3ea4f994 /* (15, 7, 1) */,
  32'h3f2b075a /* (11, 7, 1) */,
  32'h3f88838c /* (7, 7, 1) */,
  32'h3ed1d4cb /* (3, 7, 1) */,
  32'h3eaf2a10 /* (15, 3, 1) */,
  32'h3ea7dbb1 /* (11, 3, 1) */,
  32'h3ed1d4cb /* (7, 3, 1) */,
  32'h3e953797 /* (3, 3, 1) */,
  32'h3e9f2a5d /* (14, 15, 13) */,
  32'h3ec1987e /* (10, 15, 13) */,
  32'h3ec1987e /* (6, 15, 13) */,
  32'h3e9f2a5d /* (2, 15, 13) */,
  32'h3eb2cc97 /* (14, 11, 13) */,
  32'h3f41f419 /* (10, 11, 13) */,
  32'h3f41f419 /* (6, 11, 13) */,
  32'h3eb2cc97 /* (2, 11, 13) */,
  32'h3ee6ec8a /* (14, 7, 13) */,
  32'h3f982d5a /* (10, 7, 13) */,
  32'h3f982d5a /* (6, 7, 13) */,
  32'h3ee6ec8a /* (2, 7, 13) */,
  32'h3e9508f6 /* (14, 3, 13) */,
  32'h3ef2a853 /* (10, 3, 13) */,
  32'h3ef2a853 /* (6, 3, 13) */,
  32'h3e9508f6 /* (2, 3, 13) */,
  32'h3eb430e1 /* (14, 15, 9) */,
  32'h3f62162b /* (10, 15, 9) */,
  32'h3f62162b /* (6, 15, 9) */,
  32'h3eb430e1 /* (2, 15, 9) */,
  32'h3f3e2f24 /* (14, 11, 9) */,
  32'h4006bd24 /* (10, 11, 9) */,
  32'h4006bd24 /* (6, 11, 9) */,
  32'h3f3e2f24 /* (2, 11, 9) */,
  32'h3f993b79 /* (14, 7, 9) */,
  32'h406912bc /* (10, 7, 9) */,
  32'h406912bc /* (6, 7, 9) */,
  32'h3f993b79 /* (2, 7, 9) */,
  32'h3ee6ec8a /* (14, 3, 9) */,
  32'h3f982d5a /* (10, 3, 9) */,
  32'h3f982d5a /* (6, 3, 9) */,
  32'h3ee6ec8a /* (2, 3, 9) */,
  32'h3e99eb68 /* (14, 15, 5) */,
  32'h3f14d2ae /* (10, 15, 5) */,
  32'h3f14d2ae /* (6, 15, 5) */,
  32'h3e99eb68 /* (2, 15, 5) */,
  32'h3f025da2 /* (14, 11, 5) */,
  32'h3fa39217 /* (10, 11, 5) */,
  32'h3fa39217 /* (6, 11, 5) */,
  32'h3f025da2 /* (2, 11, 5) */,
  32'h3f3e2f24 /* (14, 7, 5) */,
  32'h4006bd24 /* (10, 7, 5) */,
  32'h4006bd24 /* (6, 7, 5) */,
  32'h3f3e2f24 /* (2, 7, 5) */,
  32'h3eb2cc97 /* (14, 3, 5) */,
  32'h3f41f419 /* (10, 3, 5) */,
  32'h3f41f419 /* (6, 3, 5) */,
  32'h3eb2cc97 /* (2, 3, 5) */,
  32'h3efc66bd /* (14, 15, 1) */,
  32'h3e9f454b /* (10, 15, 1) */,
  32'h3e9f454b /* (6, 15, 1) */,
  32'h3efc66bd /* (2, 15, 1) */,
  32'h3e99eb68 /* (14, 11, 1) */,
  32'h3f14d2ae /* (10, 11, 1) */,
  32'h3f14d2ae /* (6, 11, 1) */,
  32'h3e99eb68 /* (2, 11, 1) */,
  32'h3eb430e1 /* (14, 7, 1) */,
  32'h3f62162b /* (10, 7, 1) */,
  32'h3f62162b /* (6, 7, 1) */,
  32'h3eb430e1 /* (2, 7, 1) */,
  32'h3e9f2a5d /* (14, 3, 1) */,
  32'h3ec1987e /* (10, 3, 1) */,
  32'h3ec1987e /* (6, 3, 1) */,
  32'h3e9f2a5d /* (2, 3, 1) */,
  32'h3e953797 /* (13, 15, 13) */,
  32'h3ed1d4cb /* (9, 15, 13) */,
  32'h3ea7dbb1 /* (5, 15, 13) */,
  32'h3eaf2a10 /* (1, 15, 13) */,
  32'h3ec9097c /* (13, 11, 13) */,
  32'h3f6365d6 /* (9, 11, 13) */,
  32'h3f17cf64 /* (5, 11, 13) */,
  32'h3ea7dbb1 /* (1, 11, 13) */,
  32'h3f07f0f8 /* (13, 7, 13) */,
  32'h3fb9d98f /* (9, 7, 13) */,
  32'h3f6365d6 /* (5, 7, 13) */,
  32'h3ed1d4cb /* (1, 7, 13) */,
  32'h3e9a814a /* (13, 3, 13) */,
  32'h3f07f0f8 /* (9, 3, 13) */,
  32'h3ec9097c /* (5, 3, 13) */,
  32'h3e953797 /* (1, 3, 13) */,
  32'h3ed1d4cb /* (13, 15, 9) */,
  32'h3f88838c /* (9, 15, 9) */,
  32'h3f2b075a /* (5, 15, 9) */,
  32'h3ea4f994 /* (1, 15, 9) */,
  32'h3f6365d6 /* (13, 11, 9) */,
  32'h40278361 /* (9, 11, 9) */,
  32'h3fc5882d /* (5, 11, 9) */,
  32'h3f2b075a /* (1, 11, 9) */,
  32'h3fb9d98f /* (13, 7, 9) */,
  32'h4093adcc /* (9, 7, 9) */,
  32'h40278361 /* (5, 7, 9) */,
  32'h3f88838c /* (1, 7, 9) */,
  32'h3f07f0f8 /* (13, 3, 9) */,
  32'h3fb9d98f /* (9, 3, 9) */,
  32'h3f6365d6 /* (5, 3, 9) */,
  32'h3ed1d4cb /* (1, 3, 9) */,
  32'h3ea7dbb1 /* (13, 15, 5) */,
  32'h3f2b075a /* (9, 15, 5) */,
  32'h3eeeb6df /* (5, 15, 5) */,
  32'h3e93e191 /* (1, 15, 5) */,
  32'h3f17cf64 /* (13, 11, 5) */,
  32'h3fc5882d /* (9, 11, 5) */,
  32'h3f77795a /* (5, 11, 5) */,
  32'h3eeeb6df /* (1, 11, 5) */,
  32'h3f6365d6 /* (13, 7, 5) */,
  32'h40278361 /* (9, 7, 5) */,
  32'h3fc5882d /* (5, 7, 5) */,
  32'h3f2b075a /* (1, 7, 5) */,
  32'h3ec9097c /* (13, 3, 5) */,
  32'h3f6365d6 /* (9, 3, 5) */,
  32'h3f17cf64 /* (5, 3, 5) */,
  32'h3ea7dbb1 /* (1, 3, 5) */,
  32'h3eaf2a10 /* (13, 15, 1) */,
  32'h3ea4f994 /* (9, 15, 1) */,
  32'h3e93e191 /* (5, 15, 1) */,
  32'h3f5a3fd8 /* (1, 15, 1) */,
  32'h3ea7dbb1 /* (13, 11, 1) */,
  32'h3f2b075a /* (9, 11, 1) */,
  32'h3eeeb6df /* (5, 11, 1) */,
  32'h3e93e191 /* (1, 11, 1) */,
  32'h3ed1d4cb /* (13, 7, 1) */,
  32'h3f88838c /* (9, 7, 1) */,
  32'h3f2b075a /* (5, 7, 1) */,
  32'h3ea4f994 /* (1, 7, 1) */,
  32'h3e953797 /* (13, 3, 1) */,
  32'h3ed1d4cb /* (9, 3, 1) */,
  32'h3ea7dbb1 /* (5, 3, 1) */,
  32'h3eaf2a10 /* (1, 3, 1) */,
  32'h3e97a967 /* (12, 15, 13) */,
  32'h3eb9823a /* (8, 15, 13) */,
  32'h3e97a967 /* (4, 15, 13) */,
  32'h3eb78ea1 /* (0, 15, 13) */,
  32'h3ef076ff /* (12, 11, 13) */,
  32'h3f558e61 /* (8, 11, 13) */,
  32'h3ef076ff /* (4, 11, 13) */,
  32'h3ea49cf9 /* (0, 11, 13) */,
  32'h3f2b2ff1 /* (12, 7, 13) */,
  32'h3fb4be0d /* (8, 7, 13) */,
  32'h3f2b2ff1 /* (4, 7, 13) */,
  32'h3ecb578e /* (0, 7, 13) */,
  32'h3eaaa637 /* (12, 3, 13) */,
  32'h3ef65451 /* (8, 3, 13) */,
  32'h3eaaa637 /* (4, 3, 13) */,
  32'h3e960c85 /* (0, 3, 13) */,
  32'h3f0271c0 /* (12, 15, 9) */,
  32'h3f8374c7 /* (8, 15, 9) */,
  32'h3f0271c0 /* (4, 15, 9) */,
  32'h3ea04e75 /* (0, 15, 9) */,
  32'h3f91d65e /* (12, 11, 9) */,
  32'h40258eba /* (8, 11, 9) */,
  32'h3f91d65e /* (4, 11, 9) */,
  32'h3f2521d3 /* (0, 11, 9) */,
  32'h3ff29d82 /* (12, 7, 9) */,
  32'h4094977b /* (8, 7, 9) */,
  32'h3ff29d82 /* (4, 7, 9) */,
  32'h3f836079 /* (0, 7, 9) */,
  32'h3f2b2ff1 /* (12, 3, 9) */,
  32'h3fb4be0d /* (8, 3, 9) */,
  32'h3f2b2ff1 /* (4, 3, 9) */,
  32'h3ecb578e /* (0, 3, 9) */,
  32'h3ec28d9a /* (12, 15, 5) */,
  32'h3f1e09be /* (8, 15, 5) */,
  32'h3ec28d9a /* (4, 15, 5) */,
  32'h3e924c17 /* (0, 15, 5) */,
  32'h3f3cbfdf /* (12, 11, 5) */,
  32'h3fbe36ae /* (8, 11, 5) */,
  32'h3f3cbfdf /* (4, 11, 5) */,
  32'h3ee7f590 /* (0, 11, 5) */,
  32'h3f91d65e /* (12, 7, 5) */,
  32'h40258eba /* (8, 7, 5) */,
  32'h3f91d65e /* (4, 7, 5) */,
  32'h3f2521d3 /* (0, 7, 5) */,
  32'h3ef076ff /* (12, 3, 5) */,
  32'h3f558e61 /* (8, 3, 5) */,
  32'h3ef076ff /* (4, 3, 5) */,
  32'h3ea49cf9 /* (0, 3, 5) */,
  32'h3e94e1d9 /* (12, 15, 1) */,
  32'h3e8d5b73 /* (8, 15, 1) */,
  32'h3e94e1d9 /* (4, 15, 1) */,
  32'h3f9befb2 /* (0, 15, 1) */,
  32'h3ec28d9a /* (12, 11, 1) */,
  32'h3f1e09be /* (8, 11, 1) */,
  32'h3ec28d9a /* (4, 11, 1) */,
  32'h3e924c17 /* (0, 11, 1) */,
  32'h3f0271c0 /* (12, 7, 1) */,
  32'h3f8374c7 /* (8, 7, 1) */,
  32'h3f0271c0 /* (4, 7, 1) */,
  32'h3ea04e75 /* (0, 7, 1) */,
  32'h3e97a967 /* (12, 3, 1) */,
  32'h3eb9823a /* (8, 3, 1) */,
  32'h3e97a967 /* (4, 3, 1) */,
  32'h3eb78ea1 /* (0, 3, 1) */,
  32'h3e9f2a5d /* (15, 14, 13) */,
  32'h3eb2cc97 /* (11, 14, 13) */,
  32'h3ee6ec8a /* (7, 14, 13) */,
  32'h3e9508f6 /* (3, 14, 13) */,
  32'h3ec1987e /* (15, 10, 13) */,
  32'h3f41f419 /* (11, 10, 13) */,
  32'h3f982d5a /* (7, 10, 13) */,
  32'h3ef2a853 /* (3, 10, 13) */,
  32'h3ec1987e /* (15, 6, 13) */,
  32'h3f41f419 /* (11, 6, 13) */,
  32'h3f982d5a /* (7, 6, 13) */,
  32'h3ef2a853 /* (3, 6, 13) */,
  32'h3e9f2a5d /* (15, 2, 13) */,
  32'h3eb2cc97 /* (11, 2, 13) */,
  32'h3ee6ec8a /* (7, 2, 13) */,
  32'h3e9508f6 /* (3, 2, 13) */,
  32'h3eb430e1 /* (15, 14, 9) */,
  32'h3f3e2f24 /* (11, 14, 9) */,
  32'h3f993b79 /* (7, 14, 9) */,
  32'h3ee6ec8a /* (3, 14, 9) */,
  32'h3f62162b /* (15, 10, 9) */,
  32'h4006bd24 /* (11, 10, 9) */,
  32'h406912bc /* (7, 10, 9) */,
  32'h3f982d5a /* (3, 10, 9) */,
  32'h3f62162b /* (15, 6, 9) */,
  32'h4006bd24 /* (11, 6, 9) */,
  32'h406912bc /* (7, 6, 9) */,
  32'h3f982d5a /* (3, 6, 9) */,
  32'h3eb430e1 /* (15, 2, 9) */,
  32'h3f3e2f24 /* (11, 2, 9) */,
  32'h3f993b79 /* (7, 2, 9) */,
  32'h3ee6ec8a /* (3, 2, 9) */,
  32'h3e99eb68 /* (15, 14, 5) */,
  32'h3f025da2 /* (11, 14, 5) */,
  32'h3f3e2f24 /* (7, 14, 5) */,
  32'h3eb2cc97 /* (3, 14, 5) */,
  32'h3f14d2ae /* (15, 10, 5) */,
  32'h3fa39217 /* (11, 10, 5) */,
  32'h4006bd24 /* (7, 10, 5) */,
  32'h3f41f419 /* (3, 10, 5) */,
  32'h3f14d2ae /* (15, 6, 5) */,
  32'h3fa39217 /* (11, 6, 5) */,
  32'h4006bd24 /* (7, 6, 5) */,
  32'h3f41f419 /* (3, 6, 5) */,
  32'h3e99eb68 /* (15, 2, 5) */,
  32'h3f025da2 /* (11, 2, 5) */,
  32'h3f3e2f24 /* (7, 2, 5) */,
  32'h3eb2cc97 /* (3, 2, 5) */,
  32'h3efc66bd /* (15, 14, 1) */,
  32'h3e99eb68 /* (11, 14, 1) */,
  32'h3eb430e1 /* (7, 14, 1) */,
  32'h3e9f2a5d /* (3, 14, 1) */,
  32'h3e9f454b /* (15, 10, 1) */,
  32'h3f14d2ae /* (11, 10, 1) */,
  32'h3f62162b /* (7, 10, 1) */,
  32'h3ec1987e /* (3, 10, 1) */,
  32'h3e9f454b /* (15, 6, 1) */,
  32'h3f14d2ae /* (11, 6, 1) */,
  32'h3f62162b /* (7, 6, 1) */,
  32'h3ec1987e /* (3, 6, 1) */,
  32'h3efc66bd /* (15, 2, 1) */,
  32'h3e99eb68 /* (11, 2, 1) */,
  32'h3eb430e1 /* (7, 2, 1) */,
  32'h3e9f2a5d /* (3, 2, 1) */,
  32'h3e9796af /* (14, 14, 13) */,
  32'h3ed22ea6 /* (10, 14, 13) */,
  32'h3ed22ea6 /* (6, 14, 13) */,
  32'h3e9796af /* (2, 14, 13) */,
  32'h3ed22ea6 /* (14, 10, 13) */,
  32'h3f7e11f4 /* (10, 10, 13) */,
  32'h3f7e11f4 /* (6, 10, 13) */,
  32'h3ed22ea6 /* (2, 10, 13) */,
  32'h3ed22ea6 /* (14, 6, 13) */,
  32'h3f7e11f4 /* (10, 6, 13) */,
  32'h3f7e11f4 /* (6, 6, 13) */,
  32'h3ed22ea6 /* (2, 6, 13) */,
  32'h3e9796af /* (14, 2, 13) */,
  32'h3ed22ea6 /* (10, 2, 13) */,
  32'h3ed22ea6 /* (6, 2, 13) */,
  32'h3e9796af /* (2, 2, 13) */,
  32'h3ec56b70 /* (14, 14, 9) */,
  32'h3f7ca6c7 /* (10, 14, 9) */,
  32'h3f7ca6c7 /* (6, 14, 9) */,
  32'h3ec56b70 /* (2, 14, 9) */,
  32'h3f7ca6c7 /* (14, 10, 9) */,
  32'h4039abaa /* (10, 10, 9) */,
  32'h4039abaa /* (6, 10, 9) */,
  32'h3f7ca6c7 /* (2, 10, 9) */,
  32'h3f7ca6c7 /* (14, 6, 9) */,
  32'h4039abaa /* (10, 6, 9) */,
  32'h4039abaa /* (6, 6, 9) */,
  32'h3f7ca6c7 /* (2, 6, 9) */,
  32'h3ec56b70 /* (14, 2, 9) */,
  32'h3f7ca6c7 /* (10, 2, 9) */,
  32'h3f7ca6c7 /* (6, 2, 9) */,
  32'h3ec56b70 /* (2, 2, 9) */,
  32'h3ea1d2a3 /* (14, 14, 5) */,
  32'h3f242ada /* (10, 14, 5) */,
  32'h3f242ada /* (6, 14, 5) */,
  32'h3ea1d2a3 /* (2, 14, 5) */,
  32'h3f242ada /* (14, 10, 5) */,
  32'h3fdbd2f0 /* (10, 10, 5) */,
  32'h3fdbd2f0 /* (6, 10, 5) */,
  32'h3f242ada /* (2, 10, 5) */,
  32'h3f242ada /* (14, 6, 5) */,
  32'h3fdbd2f0 /* (10, 6, 5) */,
  32'h3fdbd2f0 /* (6, 6, 5) */,
  32'h3f242ada /* (2, 6, 5) */,
  32'h3ea1d2a3 /* (14, 2, 5) */,
  32'h3f242ada /* (10, 2, 5) */,
  32'h3f242ada /* (6, 2, 5) */,
  32'h3ea1d2a3 /* (2, 2, 5) */,
  32'h3ec29928 /* (14, 14, 1) */,
  32'h3eaab74a /* (10, 14, 1) */,
  32'h3eaab74a /* (6, 14, 1) */,
  32'h3ec29928 /* (2, 14, 1) */,
  32'h3eaab74a /* (14, 10, 1) */,
  32'h3f3f980b /* (10, 10, 1) */,
  32'h3f3f980b /* (6, 10, 1) */,
  32'h3eaab74a /* (2, 10, 1) */,
  32'h3eaab74a /* (14, 6, 1) */,
  32'h3f3f980b /* (10, 6, 1) */,
  32'h3f3f980b /* (6, 6, 1) */,
  32'h3eaab74a /* (2, 6, 1) */,
  32'h3ec29928 /* (14, 2, 1) */,
  32'h3eaab74a /* (10, 2, 1) */,
  32'h3eaab74a /* (6, 2, 1) */,
  32'h3ec29928 /* (2, 2, 1) */,
  32'h3e9508f6 /* (13, 14, 13) */,
  32'h3ee6ec8a /* (9, 14, 13) */,
  32'h3eb2cc97 /* (5, 14, 13) */,
  32'h3e9f2a5d /* (1, 14, 13) */,
  32'h3ef2a853 /* (13, 10, 13) */,
  32'h3f982d5a /* (9, 10, 13) */,
  32'h3f41f419 /* (5, 10, 13) */,
  32'h3ec1987e /* (1, 10, 13) */,
  32'h3ef2a853 /* (13, 6, 13) */,
  32'h3f982d5a /* (9, 6, 13) */,
  32'h3f41f419 /* (5, 6, 13) */,
  32'h3ec1987e /* (1, 6, 13) */,
  32'h3e9508f6 /* (13, 2, 13) */,
  32'h3ee6ec8a /* (9, 2, 13) */,
  32'h3eb2cc97 /* (5, 2, 13) */,
  32'h3e9f2a5d /* (1, 2, 13) */,
  32'h3ee6ec8a /* (13, 14, 9) */,
  32'h3f993b79 /* (9, 14, 9) */,
  32'h3f3e2f24 /* (5, 14, 9) */,
  32'h3eb430e1 /* (1, 14, 9) */,
  32'h3f982d5a /* (13, 10, 9) */,
  32'h406912bc /* (9, 10, 9) */,
  32'h4006bd24 /* (5, 10, 9) */,
  32'h3f62162b /* (1, 10, 9) */,
  32'h3f982d5a /* (13, 6, 9) */,
  32'h406912bc /* (9, 6, 9) */,
  32'h4006bd24 /* (5, 6, 9) */,
  32'h3f62162b /* (1, 6, 9) */,
  32'h3ee6ec8a /* (13, 2, 9) */,
  32'h3f993b79 /* (9, 2, 9) */,
  32'h3f3e2f24 /* (5, 2, 9) */,
  32'h3eb430e1 /* (1, 2, 9) */,
  32'h3eb2cc97 /* (13, 14, 5) */,
  32'h3f3e2f24 /* (9, 14, 5) */,
  32'h3f025da2 /* (5, 14, 5) */,
  32'h3e99eb68 /* (1, 14, 5) */,
  32'h3f41f419 /* (13, 10, 5) */,
  32'h4006bd24 /* (9, 10, 5) */,
  32'h3fa39217 /* (5, 10, 5) */,
  32'h3f14d2ae /* (1, 10, 5) */,
  32'h3f41f419 /* (13, 6, 5) */,
  32'h4006bd24 /* (9, 6, 5) */,
  32'h3fa39217 /* (5, 6, 5) */,
  32'h3f14d2ae /* (1, 6, 5) */,
  32'h3eb2cc97 /* (13, 2, 5) */,
  32'h3f3e2f24 /* (9, 2, 5) */,
  32'h3f025da2 /* (5, 2, 5) */,
  32'h3e99eb68 /* (1, 2, 5) */,
  32'h3e9f2a5d /* (13, 14, 1) */,
  32'h3eb430e1 /* (9, 14, 1) */,
  32'h3e99eb68 /* (5, 14, 1) */,
  32'h3efc66bd /* (1, 14, 1) */,
  32'h3ec1987e /* (13, 10, 1) */,
  32'h3f62162b /* (9, 10, 1) */,
  32'h3f14d2ae /* (5, 10, 1) */,
  32'h3e9f454b /* (1, 10, 1) */,
  32'h3ec1987e /* (13, 6, 1) */,
  32'h3f62162b /* (9, 6, 1) */,
  32'h3f14d2ae /* (5, 6, 1) */,
  32'h3e9f454b /* (1, 6, 1) */,
  32'h3e9f2a5d /* (13, 2, 1) */,
  32'h3eb430e1 /* (9, 2, 1) */,
  32'h3e99eb68 /* (5, 2, 1) */,
  32'h3efc66bd /* (1, 2, 1) */,
  32'h3e9d3fef /* (12, 14, 13) */,
  32'h3ece2dc1 /* (8, 14, 13) */,
  32'h3e9d3fef /* (4, 14, 13) */,
  32'h3ea34ae8 /* (0, 14, 13) */,
  32'h3f15625b /* (12, 10, 13) */,
  32'h3f91854a /* (8, 10, 13) */,
  32'h3f15625b /* (4, 10, 13) */,
  32'h3ebc86f4 /* (0, 10, 13) */,
  32'h3f15625b /* (12, 6, 13) */,
  32'h3f91854a /* (8, 6, 13) */,
  32'h3f15625b /* (4, 6, 13) */,
  32'h3ebc86f4 /* (0, 6, 13) */,
  32'h3e9d3fef /* (12, 2, 13) */,
  32'h3ece2dc1 /* (8, 2, 13) */,
  32'h3e9d3fef /* (4, 2, 13) */,
  32'h3ea34ae8 /* (0, 2, 13) */,
  32'h3f104c25 /* (12, 14, 9) */,
  32'h3f9420e3 /* (8, 14, 9) */,
  32'h3f104c25 /* (4, 14, 9) */,
  32'h3eaee5c8 /* (0, 14, 9) */,
  32'h3fc4fc22 /* (12, 10, 9) */,
  32'h40686d0d /* (8, 10, 9) */,
  32'h3fc4fc22 /* (4, 10, 9) */,
  32'h3f59ea43 /* (0, 10, 9) */,
  32'h3fc4fc22 /* (12, 6, 9) */,
  32'h40686d0d /* (8, 6, 9) */,
  32'h3fc4fc22 /* (4, 6, 9) */,
  32'h3f59ea43 /* (0, 6, 9) */,
  32'h3f104c25 /* (12, 2, 9) */,
  32'h3f9420e3 /* (8, 2, 9) */,
  32'h3f104c25 /* (4, 2, 9) */,
  32'h3eaee5c8 /* (0, 2, 9) */,
  32'h3ed1ff4c /* (12, 14, 5) */,
  32'h3f30df4f /* (8, 14, 5) */,
  32'h3ed1ff4c /* (4, 14, 5) */,
  32'h3e97b006 /* (0, 14, 5) */,
  32'h3f753c17 /* (12, 10, 5) */,
  32'h40037a14 /* (8, 10, 5) */,
  32'h3f753c17 /* (4, 10, 5) */,
  32'h3f1019ab /* (0, 10, 5) */,
  32'h3f753c17 /* (12, 6, 5) */,
  32'h40037a14 /* (8, 6, 5) */,
  32'h3f753c17 /* (4, 6, 5) */,
  32'h3f1019ab /* (0, 6, 5) */,
  32'h3ed1ff4c /* (12, 2, 5) */,
  32'h3f30df4f /* (8, 2, 5) */,
  32'h3ed1ff4c /* (4, 2, 5) */,
  32'h3e97b006 /* (0, 2, 5) */,
  32'h3e939519 /* (12, 14, 1) */,
  32'h3e9c5e8a /* (8, 14, 1) */,
  32'h3e939519 /* (4, 14, 1) */,
  32'h3f10451b /* (0, 14, 1) */,
  32'h3ee9b2a2 /* (12, 10, 1) */,
  32'h3f5576ec /* (8, 10, 1) */,
  32'h3ee9b2a2 /* (4, 10, 1) */,
  32'h3e9bd472 /* (0, 10, 1) */,
  32'h3ee9b2a2 /* (12, 6, 1) */,
  32'h3f5576ec /* (8, 6, 1) */,
  32'h3ee9b2a2 /* (4, 6, 1) */,
  32'h3e9bd472 /* (0, 6, 1) */,
  32'h3e939519 /* (12, 2, 1) */,
  32'h3e9c5e8a /* (8, 2, 1) */,
  32'h3e939519 /* (4, 2, 1) */,
  32'h3f10451b /* (0, 2, 1) */,
  32'h3e953797 /* (15, 13, 13) */,
  32'h3ec9097c /* (11, 13, 13) */,
  32'h3f07f0f8 /* (7, 13, 13) */,
  32'h3e9a814a /* (3, 13, 13) */,
  32'h3ed1d4cb /* (15, 9, 13) */,
  32'h3f6365d6 /* (11, 9, 13) */,
  32'h3fb9d98f /* (7, 9, 13) */,
  32'h3f07f0f8 /* (3, 9, 13) */,
  32'h3ea7dbb1 /* (15, 5, 13) */,
  32'h3f17cf64 /* (11, 5, 13) */,
  32'h3f6365d6 /* (7, 5, 13) */,
  32'h3ec9097c /* (3, 5, 13) */,
  32'h3eaf2a10 /* (15, 1, 13) */,
  32'h3ea7dbb1 /* (11, 1, 13) */,
  32'h3ed1d4cb /* (7, 1, 13) */,
  32'h3e953797 /* (3, 1, 13) */,
  32'h3ed1d4cb /* (15, 13, 9) */,
  32'h3f6365d6 /* (11, 13, 9) */,
  32'h3fb9d98f /* (7, 13, 9) */,
  32'h3f07f0f8 /* (3, 13, 9) */,
  32'h3f88838c /* (15, 9, 9) */,
  32'h40278361 /* (11, 9, 9) */,
  32'h4093adcc /* (7, 9, 9) */,
  32'h3fb9d98f /* (3, 9, 9) */,
  32'h3f2b075a /* (15, 5, 9) */,
  32'h3fc5882d /* (11, 5, 9) */,
  32'h40278361 /* (7, 5, 9) */,
  32'h3f6365d6 /* (3, 5, 9) */,
  32'h3ea4f994 /* (15, 1, 9) */,
  32'h3f2b075a /* (11, 1, 9) */,
  32'h3f88838c /* (7, 1, 9) */,
  32'h3ed1d4cb /* (3, 1, 9) */,
  32'h3ea7dbb1 /* (15, 13, 5) */,
  32'h3f17cf64 /* (11, 13, 5) */,
  32'h3f6365d6 /* (7, 13, 5) */,
  32'h3ec9097c /* (3, 13, 5) */,
  32'h3f2b075a /* (15, 9, 5) */,
  32'h3fc5882d /* (11, 9, 5) */,
  32'h40278361 /* (7, 9, 5) */,
  32'h3f6365d6 /* (3, 9, 5) */,
  32'h3eeeb6df /* (15, 5, 5) */,
  32'h3f77795a /* (11, 5, 5) */,
  32'h3fc5882d /* (7, 5, 5) */,
  32'h3f17cf64 /* (3, 5, 5) */,
  32'h3e93e191 /* (15, 1, 5) */,
  32'h3eeeb6df /* (11, 1, 5) */,
  32'h3f2b075a /* (7, 1, 5) */,
  32'h3ea7dbb1 /* (3, 1, 5) */,
  32'h3eaf2a10 /* (15, 13, 1) */,
  32'h3ea7dbb1 /* (11, 13, 1) */,
  32'h3ed1d4cb /* (7, 13, 1) */,
  32'h3e953797 /* (3, 13, 1) */,
  32'h3ea4f994 /* (15, 9, 1) */,
  32'h3f2b075a /* (11, 9, 1) */,
  32'h3f88838c /* (7, 9, 1) */,
  32'h3ed1d4cb /* (3, 9, 1) */,
  32'h3e93e191 /* (15, 5, 1) */,
  32'h3eeeb6df /* (11, 5, 1) */,
  32'h3f2b075a /* (7, 5, 1) */,
  32'h3ea7dbb1 /* (3, 5, 1) */,
  32'h3f5a3fd8 /* (15, 1, 1) */,
  32'h3e93e191 /* (11, 1, 1) */,
  32'h3ea4f994 /* (7, 1, 1) */,
  32'h3eaf2a10 /* (3, 1, 1) */,
  32'h3e9508f6 /* (14, 13, 13) */,
  32'h3ef2a853 /* (10, 13, 13) */,
  32'h3ef2a853 /* (6, 13, 13) */,
  32'h3e9508f6 /* (2, 13, 13) */,
  32'h3ee6ec8a /* (14, 9, 13) */,
  32'h3f982d5a /* (10, 9, 13) */,
  32'h3f982d5a /* (6, 9, 13) */,
  32'h3ee6ec8a /* (2, 9, 13) */,
  32'h3eb2cc97 /* (14, 5, 13) */,
  32'h3f41f419 /* (10, 5, 13) */,
  32'h3f41f419 /* (6, 5, 13) */,
  32'h3eb2cc97 /* (2, 5, 13) */,
  32'h3e9f2a5d /* (14, 1, 13) */,
  32'h3ec1987e /* (10, 1, 13) */,
  32'h3ec1987e /* (6, 1, 13) */,
  32'h3e9f2a5d /* (2, 1, 13) */,
  32'h3ee6ec8a /* (14, 13, 9) */,
  32'h3f982d5a /* (10, 13, 9) */,
  32'h3f982d5a /* (6, 13, 9) */,
  32'h3ee6ec8a /* (2, 13, 9) */,
  32'h3f993b79 /* (14, 9, 9) */,
  32'h406912bc /* (10, 9, 9) */,
  32'h406912bc /* (6, 9, 9) */,
  32'h3f993b79 /* (2, 9, 9) */,
  32'h3f3e2f24 /* (14, 5, 9) */,
  32'h4006bd24 /* (10, 5, 9) */,
  32'h4006bd24 /* (6, 5, 9) */,
  32'h3f3e2f24 /* (2, 5, 9) */,
  32'h3eb430e1 /* (14, 1, 9) */,
  32'h3f62162b /* (10, 1, 9) */,
  32'h3f62162b /* (6, 1, 9) */,
  32'h3eb430e1 /* (2, 1, 9) */,
  32'h3eb2cc97 /* (14, 13, 5) */,
  32'h3f41f419 /* (10, 13, 5) */,
  32'h3f41f419 /* (6, 13, 5) */,
  32'h3eb2cc97 /* (2, 13, 5) */,
  32'h3f3e2f24 /* (14, 9, 5) */,
  32'h4006bd24 /* (10, 9, 5) */,
  32'h4006bd24 /* (6, 9, 5) */,
  32'h3f3e2f24 /* (2, 9, 5) */,
  32'h3f025da2 /* (14, 5, 5) */,
  32'h3fa39217 /* (10, 5, 5) */,
  32'h3fa39217 /* (6, 5, 5) */,
  32'h3f025da2 /* (2, 5, 5) */,
  32'h3e99eb68 /* (14, 1, 5) */,
  32'h3f14d2ae /* (10, 1, 5) */,
  32'h3f14d2ae /* (6, 1, 5) */,
  32'h3e99eb68 /* (2, 1, 5) */,
  32'h3e9f2a5d /* (14, 13, 1) */,
  32'h3ec1987e /* (10, 13, 1) */,
  32'h3ec1987e /* (6, 13, 1) */,
  32'h3e9f2a5d /* (2, 13, 1) */,
  32'h3eb430e1 /* (14, 9, 1) */,
  32'h3f62162b /* (10, 9, 1) */,
  32'h3f62162b /* (6, 9, 1) */,
  32'h3eb430e1 /* (2, 9, 1) */,
  32'h3e99eb68 /* (14, 5, 1) */,
  32'h3f14d2ae /* (10, 5, 1) */,
  32'h3f14d2ae /* (6, 5, 1) */,
  32'h3e99eb68 /* (2, 5, 1) */,
  32'h3efc66bd /* (14, 1, 1) */,
  32'h3e9f454b /* (10, 1, 1) */,
  32'h3e9f454b /* (6, 1, 1) */,
  32'h3efc66bd /* (2, 1, 1) */,
  32'h3e9a814a /* (13, 13, 13) */,
  32'h3f07f0f8 /* (9, 13, 13) */,
  32'h3ec9097c /* (5, 13, 13) */,
  32'h3e953797 /* (1, 13, 13) */,
  32'h3f07f0f8 /* (13, 9, 13) */,
  32'h3fb9d98f /* (9, 9, 13) */,
  32'h3f6365d6 /* (5, 9, 13) */,
  32'h3ed1d4cb /* (1, 9, 13) */,
  32'h3ec9097c /* (13, 5, 13) */,
  32'h3f6365d6 /* (9, 5, 13) */,
  32'h3f17cf64 /* (5, 5, 13) */,
  32'h3ea7dbb1 /* (1, 5, 13) */,
  32'h3e953797 /* (13, 1, 13) */,
  32'h3ed1d4cb /* (9, 1, 13) */,
  32'h3ea7dbb1 /* (5, 1, 13) */,
  32'h3eaf2a10 /* (1, 1, 13) */,
  32'h3f07f0f8 /* (13, 13, 9) */,
  32'h3fb9d98f /* (9, 13, 9) */,
  32'h3f6365d6 /* (5, 13, 9) */,
  32'h3ed1d4cb /* (1, 13, 9) */,
  32'h3fb9d98f /* (13, 9, 9) */,
  32'h4093adcc /* (9, 9, 9) */,
  32'h40278361 /* (5, 9, 9) */,
  32'h3f88838c /* (1, 9, 9) */,
  32'h3f6365d6 /* (13, 5, 9) */,
  32'h40278361 /* (9, 5, 9) */,
  32'h3fc5882d /* (5, 5, 9) */,
  32'h3f2b075a /* (1, 5, 9) */,
  32'h3ed1d4cb /* (13, 1, 9) */,
  32'h3f88838c /* (9, 1, 9) */,
  32'h3f2b075a /* (5, 1, 9) */,
  32'h3ea4f994 /* (1, 1, 9) */,
  32'h3ec9097c /* (13, 13, 5) */,
  32'h3f6365d6 /* (9, 13, 5) */,
  32'h3f17cf64 /* (5, 13, 5) */,
  32'h3ea7dbb1 /* (1, 13, 5) */,
  32'h3f6365d6 /* (13, 9, 5) */,
  32'h40278361 /* (9, 9, 5) */,
  32'h3fc5882d /* (5, 9, 5) */,
  32'h3f2b075a /* (1, 9, 5) */,
  32'h3f17cf64 /* (13, 5, 5) */,
  32'h3fc5882d /* (9, 5, 5) */,
  32'h3f77795a /* (5, 5, 5) */,
  32'h3eeeb6df /* (1, 5, 5) */,
  32'h3ea7dbb1 /* (13, 1, 5) */,
  32'h3f2b075a /* (9, 1, 5) */,
  32'h3eeeb6df /* (5, 1, 5) */,
  32'h3e93e191 /* (1, 1, 5) */,
  32'h3e953797 /* (13, 13, 1) */,
  32'h3ed1d4cb /* (9, 13, 1) */,
  32'h3ea7dbb1 /* (5, 13, 1) */,
  32'h3eaf2a10 /* (1, 13, 1) */,
  32'h3ed1d4cb /* (13, 9, 1) */,
  32'h3f88838c /* (9, 9, 1) */,
  32'h3f2b075a /* (5, 9, 1) */,
  32'h3ea4f994 /* (1, 9, 1) */,
  32'h3ea7dbb1 /* (13, 5, 1) */,
  32'h3f2b075a /* (9, 5, 1) */,
  32'h3eeeb6df /* (5, 5, 1) */,
  32'h3e93e191 /* (1, 5, 1) */,
  32'h3eaf2a10 /* (13, 1, 1) */,
  32'h3ea4f994 /* (9, 1, 1) */,
  32'h3e93e191 /* (5, 1, 1) */,
  32'h3f5a3fd8 /* (1, 1, 1) */,
  32'h3eaaa637 /* (12, 13, 13) */,
  32'h3ef65451 /* (8, 13, 13) */,
  32'h3eaaa637 /* (4, 13, 13) */,
  32'h3e960c85 /* (0, 13, 13) */,
  32'h3f2b2ff1 /* (12, 9, 13) */,
  32'h3fb4be0d /* (8, 9, 13) */,
  32'h3f2b2ff1 /* (4, 9, 13) */,
  32'h3ecb578e /* (0, 9, 13) */,
  32'h3ef076ff /* (12, 5, 13) */,
  32'h3f558e61 /* (8, 5, 13) */,
  32'h3ef076ff /* (4, 5, 13) */,
  32'h3ea49cf9 /* (0, 5, 13) */,
  32'h3e97a967 /* (12, 1, 13) */,
  32'h3eb9823a /* (8, 1, 13) */,
  32'h3e97a967 /* (4, 1, 13) */,
  32'h3eb78ea1 /* (0, 1, 13) */,
  32'h3f2b2ff1 /* (12, 13, 9) */,
  32'h3fb4be0d /* (8, 13, 9) */,
  32'h3f2b2ff1 /* (4, 13, 9) */,
  32'h3ecb578e /* (0, 13, 9) */,
  32'h3ff29d82 /* (12, 9, 9) */,
  32'h4094977b /* (8, 9, 9) */,
  32'h3ff29d82 /* (4, 9, 9) */,
  32'h3f836079 /* (0, 9, 9) */,
  32'h3f91d65e /* (12, 5, 9) */,
  32'h40258eba /* (8, 5, 9) */,
  32'h3f91d65e /* (4, 5, 9) */,
  32'h3f2521d3 /* (0, 5, 9) */,
  32'h3f0271c0 /* (12, 1, 9) */,
  32'h3f8374c7 /* (8, 1, 9) */,
  32'h3f0271c0 /* (4, 1, 9) */,
  32'h3ea04e75 /* (0, 1, 9) */,
  32'h3ef076ff /* (12, 13, 5) */,
  32'h3f558e61 /* (8, 13, 5) */,
  32'h3ef076ff /* (4, 13, 5) */,
  32'h3ea49cf9 /* (0, 13, 5) */,
  32'h3f91d65e /* (12, 9, 5) */,
  32'h40258eba /* (8, 9, 5) */,
  32'h3f91d65e /* (4, 9, 5) */,
  32'h3f2521d3 /* (0, 9, 5) */,
  32'h3f3cbfdf /* (12, 5, 5) */,
  32'h3fbe36ae /* (8, 5, 5) */,
  32'h3f3cbfdf /* (4, 5, 5) */,
  32'h3ee7f590 /* (0, 5, 5) */,
  32'h3ec28d9a /* (12, 1, 5) */,
  32'h3f1e09be /* (8, 1, 5) */,
  32'h3ec28d9a /* (4, 1, 5) */,
  32'h3e924c17 /* (0, 1, 5) */,
  32'h3e97a967 /* (12, 13, 1) */,
  32'h3eb9823a /* (8, 13, 1) */,
  32'h3e97a967 /* (4, 13, 1) */,
  32'h3eb78ea1 /* (0, 13, 1) */,
  32'h3f0271c0 /* (12, 9, 1) */,
  32'h3f8374c7 /* (8, 9, 1) */,
  32'h3f0271c0 /* (4, 9, 1) */,
  32'h3ea04e75 /* (0, 9, 1) */,
  32'h3ec28d9a /* (12, 5, 1) */,
  32'h3f1e09be /* (8, 5, 1) */,
  32'h3ec28d9a /* (4, 5, 1) */,
  32'h3e924c17 /* (0, 5, 1) */,
  32'h3e94e1d9 /* (12, 1, 1) */,
  32'h3e8d5b73 /* (8, 1, 1) */,
  32'h3e94e1d9 /* (4, 1, 1) */,
  32'h3f9befb2 /* (0, 1, 1) */,
  32'h3e97a967 /* (15, 12, 13) */,
  32'h3ef076ff /* (11, 12, 13) */,
  32'h3f2b2ff1 /* (7, 12, 13) */,
  32'h3eaaa637 /* (3, 12, 13) */,
  32'h3eb9823a /* (15, 8, 13) */,
  32'h3f558e61 /* (11, 8, 13) */,
  32'h3fb4be0d /* (7, 8, 13) */,
  32'h3ef65451 /* (3, 8, 13) */,
  32'h3e97a967 /* (15, 4, 13) */,
  32'h3ef076ff /* (11, 4, 13) */,
  32'h3f2b2ff1 /* (7, 4, 13) */,
  32'h3eaaa637 /* (3, 4, 13) */,
  32'h3eb78ea1 /* (15, 0, 13) */,
  32'h3ea49cf9 /* (11, 0, 13) */,
  32'h3ecb578e /* (7, 0, 13) */,
  32'h3e960c85 /* (3, 0, 13) */,
  32'h3f0271c0 /* (15, 12, 9) */,
  32'h3f91d65e /* (11, 12, 9) */,
  32'h3ff29d82 /* (7, 12, 9) */,
  32'h3f2b2ff1 /* (3, 12, 9) */,
  32'h3f8374c7 /* (15, 8, 9) */,
  32'h40258eba /* (11, 8, 9) */,
  32'h4094977b /* (7, 8, 9) */,
  32'h3fb4be0d /* (3, 8, 9) */,
  32'h3f0271c0 /* (15, 4, 9) */,
  32'h3f91d65e /* (11, 4, 9) */,
  32'h3ff29d82 /* (7, 4, 9) */,
  32'h3f2b2ff1 /* (3, 4, 9) */,
  32'h3ea04e75 /* (15, 0, 9) */,
  32'h3f2521d3 /* (11, 0, 9) */,
  32'h3f836079 /* (7, 0, 9) */,
  32'h3ecb578e /* (3, 0, 9) */,
  32'h3ec28d9a /* (15, 12, 5) */,
  32'h3f3cbfdf /* (11, 12, 5) */,
  32'h3f91d65e /* (7, 12, 5) */,
  32'h3ef076ff /* (3, 12, 5) */,
  32'h3f1e09be /* (15, 8, 5) */,
  32'h3fbe36ae /* (11, 8, 5) */,
  32'h40258eba /* (7, 8, 5) */,
  32'h3f558e61 /* (3, 8, 5) */,
  32'h3ec28d9a /* (15, 4, 5) */,
  32'h3f3cbfdf /* (11, 4, 5) */,
  32'h3f91d65e /* (7, 4, 5) */,
  32'h3ef076ff /* (3, 4, 5) */,
  32'h3e924c17 /* (15, 0, 5) */,
  32'h3ee7f590 /* (11, 0, 5) */,
  32'h3f2521d3 /* (7, 0, 5) */,
  32'h3ea49cf9 /* (3, 0, 5) */,
  32'h3e94e1d9 /* (15, 12, 1) */,
  32'h3ec28d9a /* (11, 12, 1) */,
  32'h3f0271c0 /* (7, 12, 1) */,
  32'h3e97a967 /* (3, 12, 1) */,
  32'h3e8d5b73 /* (15, 8, 1) */,
  32'h3f1e09be /* (11, 8, 1) */,
  32'h3f8374c7 /* (7, 8, 1) */,
  32'h3eb9823a /* (3, 8, 1) */,
  32'h3e94e1d9 /* (15, 4, 1) */,
  32'h3ec28d9a /* (11, 4, 1) */,
  32'h3f0271c0 /* (7, 4, 1) */,
  32'h3e97a967 /* (3, 4, 1) */,
  32'h3f9befb2 /* (15, 0, 1) */,
  32'h3e924c17 /* (11, 0, 1) */,
  32'h3ea04e75 /* (7, 0, 1) */,
  32'h3eb78ea1 /* (3, 0, 1) */,
  32'h3e9d3fef /* (14, 12, 13) */,
  32'h3f15625b /* (10, 12, 13) */,
  32'h3f15625b /* (6, 12, 13) */,
  32'h3e9d3fef /* (2, 12, 13) */,
  32'h3ece2dc1 /* (14, 8, 13) */,
  32'h3f91854a /* (10, 8, 13) */,
  32'h3f91854a /* (6, 8, 13) */,
  32'h3ece2dc1 /* (2, 8, 13) */,
  32'h3e9d3fef /* (14, 4, 13) */,
  32'h3f15625b /* (10, 4, 13) */,
  32'h3f15625b /* (6, 4, 13) */,
  32'h3e9d3fef /* (2, 4, 13) */,
  32'h3ea34ae8 /* (14, 0, 13) */,
  32'h3ebc86f4 /* (10, 0, 13) */,
  32'h3ebc86f4 /* (6, 0, 13) */,
  32'h3ea34ae8 /* (2, 0, 13) */,
  32'h3f104c25 /* (14, 12, 9) */,
  32'h3fc4fc22 /* (10, 12, 9) */,
  32'h3fc4fc22 /* (6, 12, 9) */,
  32'h3f104c25 /* (2, 12, 9) */,
  32'h3f9420e3 /* (14, 8, 9) */,
  32'h40686d0d /* (10, 8, 9) */,
  32'h40686d0d /* (6, 8, 9) */,
  32'h3f9420e3 /* (2, 8, 9) */,
  32'h3f104c25 /* (14, 4, 9) */,
  32'h3fc4fc22 /* (10, 4, 9) */,
  32'h3fc4fc22 /* (6, 4, 9) */,
  32'h3f104c25 /* (2, 4, 9) */,
  32'h3eaee5c8 /* (14, 0, 9) */,
  32'h3f59ea43 /* (10, 0, 9) */,
  32'h3f59ea43 /* (6, 0, 9) */,
  32'h3eaee5c8 /* (2, 0, 9) */,
  32'h3ed1ff4c /* (14, 12, 5) */,
  32'h3f753c17 /* (10, 12, 5) */,
  32'h3f753c17 /* (6, 12, 5) */,
  32'h3ed1ff4c /* (2, 12, 5) */,
  32'h3f30df4f /* (14, 8, 5) */,
  32'h40037a14 /* (10, 8, 5) */,
  32'h40037a14 /* (6, 8, 5) */,
  32'h3f30df4f /* (2, 8, 5) */,
  32'h3ed1ff4c /* (14, 4, 5) */,
  32'h3f753c17 /* (10, 4, 5) */,
  32'h3f753c17 /* (6, 4, 5) */,
  32'h3ed1ff4c /* (2, 4, 5) */,
  32'h3e97b006 /* (14, 0, 5) */,
  32'h3f1019ab /* (10, 0, 5) */,
  32'h3f1019ab /* (6, 0, 5) */,
  32'h3e97b006 /* (2, 0, 5) */,
  32'h3e939519 /* (14, 12, 1) */,
  32'h3ee9b2a2 /* (10, 12, 1) */,
  32'h3ee9b2a2 /* (6, 12, 1) */,
  32'h3e939519 /* (2, 12, 1) */,
  32'h3e9c5e8a /* (14, 8, 1) */,
  32'h3f5576ec /* (10, 8, 1) */,
  32'h3f5576ec /* (6, 8, 1) */,
  32'h3e9c5e8a /* (2, 8, 1) */,
  32'h3e939519 /* (14, 4, 1) */,
  32'h3ee9b2a2 /* (10, 4, 1) */,
  32'h3ee9b2a2 /* (6, 4, 1) */,
  32'h3e939519 /* (2, 4, 1) */,
  32'h3f10451b /* (14, 0, 1) */,
  32'h3e9bd472 /* (10, 0, 1) */,
  32'h3e9bd472 /* (6, 0, 1) */,
  32'h3f10451b /* (2, 0, 1) */,
  32'h3eaaa637 /* (13, 12, 13) */,
  32'h3f2b2ff1 /* (9, 12, 13) */,
  32'h3ef076ff /* (5, 12, 13) */,
  32'h3e97a967 /* (1, 12, 13) */,
  32'h3ef65451 /* (13, 8, 13) */,
  32'h3fb4be0d /* (9, 8, 13) */,
  32'h3f558e61 /* (5, 8, 13) */,
  32'h3eb9823a /* (1, 8, 13) */,
  32'h3eaaa637 /* (13, 4, 13) */,
  32'h3f2b2ff1 /* (9, 4, 13) */,
  32'h3ef076ff /* (5, 4, 13) */,
  32'h3e97a967 /* (1, 4, 13) */,
  32'h3e960c85 /* (13, 0, 13) */,
  32'h3ecb578e /* (9, 0, 13) */,
  32'h3ea49cf9 /* (5, 0, 13) */,
  32'h3eb78ea1 /* (1, 0, 13) */,
  32'h3f2b2ff1 /* (13, 12, 9) */,
  32'h3ff29d82 /* (9, 12, 9) */,
  32'h3f91d65e /* (5, 12, 9) */,
  32'h3f0271c0 /* (1, 12, 9) */,
  32'h3fb4be0d /* (13, 8, 9) */,
  32'h4094977b /* (9, 8, 9) */,
  32'h40258eba /* (5, 8, 9) */,
  32'h3f8374c7 /* (1, 8, 9) */,
  32'h3f2b2ff1 /* (13, 4, 9) */,
  32'h3ff29d82 /* (9, 4, 9) */,
  32'h3f91d65e /* (5, 4, 9) */,
  32'h3f0271c0 /* (1, 4, 9) */,
  32'h3ecb578e /* (13, 0, 9) */,
  32'h3f836079 /* (9, 0, 9) */,
  32'h3f2521d3 /* (5, 0, 9) */,
  32'h3ea04e75 /* (1, 0, 9) */,
  32'h3ef076ff /* (13, 12, 5) */,
  32'h3f91d65e /* (9, 12, 5) */,
  32'h3f3cbfdf /* (5, 12, 5) */,
  32'h3ec28d9a /* (1, 12, 5) */,
  32'h3f558e61 /* (13, 8, 5) */,
  32'h40258eba /* (9, 8, 5) */,
  32'h3fbe36ae /* (5, 8, 5) */,
  32'h3f1e09be /* (1, 8, 5) */,
  32'h3ef076ff /* (13, 4, 5) */,
  32'h3f91d65e /* (9, 4, 5) */,
  32'h3f3cbfdf /* (5, 4, 5) */,
  32'h3ec28d9a /* (1, 4, 5) */,
  32'h3ea49cf9 /* (13, 0, 5) */,
  32'h3f2521d3 /* (9, 0, 5) */,
  32'h3ee7f590 /* (5, 0, 5) */,
  32'h3e924c17 /* (1, 0, 5) */,
  32'h3e97a967 /* (13, 12, 1) */,
  32'h3f0271c0 /* (9, 12, 1) */,
  32'h3ec28d9a /* (5, 12, 1) */,
  32'h3e94e1d9 /* (1, 12, 1) */,
  32'h3eb9823a /* (13, 8, 1) */,
  32'h3f8374c7 /* (9, 8, 1) */,
  32'h3f1e09be /* (5, 8, 1) */,
  32'h3e8d5b73 /* (1, 8, 1) */,
  32'h3e97a967 /* (13, 4, 1) */,
  32'h3f0271c0 /* (9, 4, 1) */,
  32'h3ec28d9a /* (5, 4, 1) */,
  32'h3e94e1d9 /* (1, 4, 1) */,
  32'h3eb78ea1 /* (13, 0, 1) */,
  32'h3ea04e75 /* (9, 0, 1) */,
  32'h3e924c17 /* (5, 0, 1) */,
  32'h3f9befb2 /* (1, 0, 1) */,
  32'h3ec4d2c5 /* (12, 12, 13) */,
  32'h3f1dd43f /* (8, 12, 13) */,
  32'h3ec4d2c5 /* (4, 12, 13) */,
  32'h3e964277 /* (0, 12, 13) */,
  32'h3f1dd43f /* (12, 8, 13) */,
  32'h3fb27927 /* (8, 8, 13) */,
  32'h3f1dd43f /* (4, 8, 13) */,
  32'h3eb32545 /* (0, 8, 13) */,
  32'h3ec4d2c5 /* (12, 4, 13) */,
  32'h3f1dd43f /* (8, 4, 13) */,
  32'h3ec4d2c5 /* (4, 4, 13) */,
  32'h3e964277 /* (0, 4, 13) */,
  32'h3e964277 /* (12, 0, 13) */,
  32'h3eb32545 /* (8, 0, 13) */,
  32'h3e964277 /* (4, 0, 13) */,
  32'h3ec24b89 /* (0, 0, 13) */,
  32'h3f59849a /* (12, 12, 9) */,
  32'h3fedbe1f /* (8, 12, 9) */,
  32'h3f59849a /* (4, 12, 9) */,
  32'h3efc5be6 /* (0, 12, 9) */,
  32'h3fedbe1f /* (12, 8, 9) */,
  32'h4096cd97 /* (8, 8, 9) */,
  32'h3fedbe1f /* (4, 8, 9) */,
  32'h3f7cadff /* (0, 8, 9) */,
  32'h3f59849a /* (12, 4, 9) */,
  32'h3fedbe1f /* (8, 4, 9) */,
  32'h3f59849a /* (4, 4, 9) */,
  32'h3efc5be6 /* (0, 4, 9) */,
  32'h3efc5be6 /* (12, 0, 9) */,
  32'h3f7cadff /* (8, 0, 9) */,
  32'h3efc5be6 /* (4, 0, 9) */,
  32'h3e9bd51d /* (0, 0, 9) */,
  32'h3f12b00d /* (12, 12, 5) */,
  32'h3f8a9c45 /* (8, 12, 5) */,
  32'h3f12b00d /* (4, 12, 5) */,
  32'h3ebddc83 /* (0, 12, 5) */,
  32'h3f8a9c45 /* (12, 8, 5) */,
  32'h402594bb /* (8, 8, 5) */,
  32'h3f8a9c45 /* (4, 8, 5) */,
  32'h3f183f16 /* (0, 8, 5) */,
  32'h3f12b00d /* (12, 4, 5) */,
  32'h3f8a9c45 /* (8, 4, 5) */,
  32'h3f12b00d /* (4, 4, 5) */,
  32'h3ebddc83 /* (0, 4, 5) */,
  32'h3ebddc83 /* (12, 0, 5) */,
  32'h3f183f16 /* (8, 0, 5) */,
  32'h3ebddc83 /* (4, 0, 5) */,
  32'h3e90f1d9 /* (0, 0, 5) */,
  32'h3ea63161 /* (12, 12, 1) */,
  32'h3eebb725 /* (8, 12, 1) */,
  32'h3ea63161 /* (4, 12, 1) */,
  32'h3e962cf4 /* (0, 12, 1) */,
  32'h3eebb725 /* (12, 8, 1) */,
  32'h3f80d0e8 /* (8, 8, 1) */,
  32'h3eebb725 /* (4, 8, 1) */,
  32'h3e88bc50 /* (0, 8, 1) */,
  32'h3ea63161 /* (12, 4, 1) */,
  32'h3eebb725 /* (8, 4, 1) */,
  32'h3ea63161 /* (4, 4, 1) */,
  32'h3e962cf4 /* (0, 4, 1) */,
  32'h3e962cf4 /* (12, 0, 1) */,
  32'h3e88bc50 /* (8, 0, 1) */,
  32'h3e962cf4 /* (4, 0, 1) */,
  32'h40148d77 /* (0, 0, 1) */,
  32'h3e94e1d9 /* (15, 15, 12) */,
  32'h3ec28d9a /* (11, 15, 12) */,
  32'h3f0271c0 /* (7, 15, 12) */,
  32'h3e97a967 /* (3, 15, 12) */,
  32'h3ec28d9a /* (15, 11, 12) */,
  32'h3f3cbfdf /* (11, 11, 12) */,
  32'h3f91d65e /* (7, 11, 12) */,
  32'h3ef076ff /* (3, 11, 12) */,
  32'h3f0271c0 /* (15, 7, 12) */,
  32'h3f91d65e /* (11, 7, 12) */,
  32'h3ff29d82 /* (7, 7, 12) */,
  32'h3f2b2ff1 /* (3, 7, 12) */,
  32'h3e97a967 /* (15, 3, 12) */,
  32'h3ef076ff /* (11, 3, 12) */,
  32'h3f2b2ff1 /* (7, 3, 12) */,
  32'h3eaaa637 /* (3, 3, 12) */,
  32'h3e8d5b73 /* (15, 15, 8) */,
  32'h3f1e09be /* (11, 15, 8) */,
  32'h3f8374c7 /* (7, 15, 8) */,
  32'h3eb9823a /* (3, 15, 8) */,
  32'h3f1e09be /* (15, 11, 8) */,
  32'h3fbe36ae /* (11, 11, 8) */,
  32'h40258eba /* (7, 11, 8) */,
  32'h3f558e61 /* (3, 11, 8) */,
  32'h3f8374c7 /* (15, 7, 8) */,
  32'h40258eba /* (11, 7, 8) */,
  32'h4094977b /* (7, 7, 8) */,
  32'h3fb4be0d /* (3, 7, 8) */,
  32'h3eb9823a /* (15, 3, 8) */,
  32'h3f558e61 /* (11, 3, 8) */,
  32'h3fb4be0d /* (7, 3, 8) */,
  32'h3ef65451 /* (3, 3, 8) */,
  32'h3e94e1d9 /* (15, 15, 4) */,
  32'h3ec28d9a /* (11, 15, 4) */,
  32'h3f0271c0 /* (7, 15, 4) */,
  32'h3e97a967 /* (3, 15, 4) */,
  32'h3ec28d9a /* (15, 11, 4) */,
  32'h3f3cbfdf /* (11, 11, 4) */,
  32'h3f91d65e /* (7, 11, 4) */,
  32'h3ef076ff /* (3, 11, 4) */,
  32'h3f0271c0 /* (15, 7, 4) */,
  32'h3f91d65e /* (11, 7, 4) */,
  32'h3ff29d82 /* (7, 7, 4) */,
  32'h3f2b2ff1 /* (3, 7, 4) */,
  32'h3e97a967 /* (15, 3, 4) */,
  32'h3ef076ff /* (11, 3, 4) */,
  32'h3f2b2ff1 /* (7, 3, 4) */,
  32'h3eaaa637 /* (3, 3, 4) */,
  32'h3f9befb2 /* (15, 15, 0) */,
  32'h3e924c17 /* (11, 15, 0) */,
  32'h3ea04e75 /* (7, 15, 0) */,
  32'h3eb78ea1 /* (3, 15, 0) */,
  32'h3e924c17 /* (15, 11, 0) */,
  32'h3ee7f590 /* (11, 11, 0) */,
  32'h3f2521d3 /* (7, 11, 0) */,
  32'h3ea49cf9 /* (3, 11, 0) */,
  32'h3ea04e75 /* (15, 7, 0) */,
  32'h3f2521d3 /* (11, 7, 0) */,
  32'h3f836079 /* (7, 7, 0) */,
  32'h3ecb578e /* (3, 7, 0) */,
  32'h3eb78ea1 /* (15, 3, 0) */,
  32'h3ea49cf9 /* (11, 3, 0) */,
  32'h3ecb578e /* (7, 3, 0) */,
  32'h3e960c85 /* (3, 3, 0) */,
  32'h3e939519 /* (14, 15, 12) */,
  32'h3ee9b2a2 /* (10, 15, 12) */,
  32'h3ee9b2a2 /* (6, 15, 12) */,
  32'h3e939519 /* (2, 15, 12) */,
  32'h3ed1ff4c /* (14, 11, 12) */,
  32'h3f753c17 /* (10, 11, 12) */,
  32'h3f753c17 /* (6, 11, 12) */,
  32'h3ed1ff4c /* (2, 11, 12) */,
  32'h3f104c25 /* (14, 7, 12) */,
  32'h3fc4fc22 /* (10, 7, 12) */,
  32'h3fc4fc22 /* (6, 7, 12) */,
  32'h3f104c25 /* (2, 7, 12) */,
  32'h3e9d3fef /* (14, 3, 12) */,
  32'h3f15625b /* (10, 3, 12) */,
  32'h3f15625b /* (6, 3, 12) */,
  32'h3e9d3fef /* (2, 3, 12) */,
  32'h3e9c5e8a /* (14, 15, 8) */,
  32'h3f5576ec /* (10, 15, 8) */,
  32'h3f5576ec /* (6, 15, 8) */,
  32'h3e9c5e8a /* (2, 15, 8) */,
  32'h3f30df4f /* (14, 11, 8) */,
  32'h40037a14 /* (10, 11, 8) */,
  32'h40037a14 /* (6, 11, 8) */,
  32'h3f30df4f /* (2, 11, 8) */,
  32'h3f9420e3 /* (14, 7, 8) */,
  32'h40686d0d /* (10, 7, 8) */,
  32'h40686d0d /* (6, 7, 8) */,
  32'h3f9420e3 /* (2, 7, 8) */,
  32'h3ece2dc1 /* (14, 3, 8) */,
  32'h3f91854a /* (10, 3, 8) */,
  32'h3f91854a /* (6, 3, 8) */,
  32'h3ece2dc1 /* (2, 3, 8) */,
  32'h3e939519 /* (14, 15, 4) */,
  32'h3ee9b2a2 /* (10, 15, 4) */,
  32'h3ee9b2a2 /* (6, 15, 4) */,
  32'h3e939519 /* (2, 15, 4) */,
  32'h3ed1ff4c /* (14, 11, 4) */,
  32'h3f753c17 /* (10, 11, 4) */,
  32'h3f753c17 /* (6, 11, 4) */,
  32'h3ed1ff4c /* (2, 11, 4) */,
  32'h3f104c25 /* (14, 7, 4) */,
  32'h3fc4fc22 /* (10, 7, 4) */,
  32'h3fc4fc22 /* (6, 7, 4) */,
  32'h3f104c25 /* (2, 7, 4) */,
  32'h3e9d3fef /* (14, 3, 4) */,
  32'h3f15625b /* (10, 3, 4) */,
  32'h3f15625b /* (6, 3, 4) */,
  32'h3e9d3fef /* (2, 3, 4) */,
  32'h3f10451b /* (14, 15, 0) */,
  32'h3e9bd472 /* (10, 15, 0) */,
  32'h3e9bd472 /* (6, 15, 0) */,
  32'h3f10451b /* (2, 15, 0) */,
  32'h3e97b006 /* (14, 11, 0) */,
  32'h3f1019ab /* (10, 11, 0) */,
  32'h3f1019ab /* (6, 11, 0) */,
  32'h3e97b006 /* (2, 11, 0) */,
  32'h3eaee5c8 /* (14, 7, 0) */,
  32'h3f59ea43 /* (10, 7, 0) */,
  32'h3f59ea43 /* (6, 7, 0) */,
  32'h3eaee5c8 /* (2, 7, 0) */,
  32'h3ea34ae8 /* (14, 3, 0) */,
  32'h3ebc86f4 /* (10, 3, 0) */,
  32'h3ebc86f4 /* (6, 3, 0) */,
  32'h3ea34ae8 /* (2, 3, 0) */,
  32'h3e97a967 /* (13, 15, 12) */,
  32'h3f0271c0 /* (9, 15, 12) */,
  32'h3ec28d9a /* (5, 15, 12) */,
  32'h3e94e1d9 /* (1, 15, 12) */,
  32'h3ef076ff /* (13, 11, 12) */,
  32'h3f91d65e /* (9, 11, 12) */,
  32'h3f3cbfdf /* (5, 11, 12) */,
  32'h3ec28d9a /* (1, 11, 12) */,
  32'h3f2b2ff1 /* (13, 7, 12) */,
  32'h3ff29d82 /* (9, 7, 12) */,
  32'h3f91d65e /* (5, 7, 12) */,
  32'h3f0271c0 /* (1, 7, 12) */,
  32'h3eaaa637 /* (13, 3, 12) */,
  32'h3f2b2ff1 /* (9, 3, 12) */,
  32'h3ef076ff /* (5, 3, 12) */,
  32'h3e97a967 /* (1, 3, 12) */,
  32'h3eb9823a /* (13, 15, 8) */,
  32'h3f8374c7 /* (9, 15, 8) */,
  32'h3f1e09be /* (5, 15, 8) */,
  32'h3e8d5b73 /* (1, 15, 8) */,
  32'h3f558e61 /* (13, 11, 8) */,
  32'h40258eba /* (9, 11, 8) */,
  32'h3fbe36ae /* (5, 11, 8) */,
  32'h3f1e09be /* (1, 11, 8) */,
  32'h3fb4be0d /* (13, 7, 8) */,
  32'h4094977b /* (9, 7, 8) */,
  32'h40258eba /* (5, 7, 8) */,
  32'h3f8374c7 /* (1, 7, 8) */,
  32'h3ef65451 /* (13, 3, 8) */,
  32'h3fb4be0d /* (9, 3, 8) */,
  32'h3f558e61 /* (5, 3, 8) */,
  32'h3eb9823a /* (1, 3, 8) */,
  32'h3e97a967 /* (13, 15, 4) */,
  32'h3f0271c0 /* (9, 15, 4) */,
  32'h3ec28d9a /* (5, 15, 4) */,
  32'h3e94e1d9 /* (1, 15, 4) */,
  32'h3ef076ff /* (13, 11, 4) */,
  32'h3f91d65e /* (9, 11, 4) */,
  32'h3f3cbfdf /* (5, 11, 4) */,
  32'h3ec28d9a /* (1, 11, 4) */,
  32'h3f2b2ff1 /* (13, 7, 4) */,
  32'h3ff29d82 /* (9, 7, 4) */,
  32'h3f91d65e /* (5, 7, 4) */,
  32'h3f0271c0 /* (1, 7, 4) */,
  32'h3eaaa637 /* (13, 3, 4) */,
  32'h3f2b2ff1 /* (9, 3, 4) */,
  32'h3ef076ff /* (5, 3, 4) */,
  32'h3e97a967 /* (1, 3, 4) */,
  32'h3eb78ea1 /* (13, 15, 0) */,
  32'h3ea04e75 /* (9, 15, 0) */,
  32'h3e924c17 /* (5, 15, 0) */,
  32'h3f9befb2 /* (1, 15, 0) */,
  32'h3ea49cf9 /* (13, 11, 0) */,
  32'h3f2521d3 /* (9, 11, 0) */,
  32'h3ee7f590 /* (5, 11, 0) */,
  32'h3e924c17 /* (1, 11, 0) */,
  32'h3ecb578e /* (13, 7, 0) */,
  32'h3f836079 /* (9, 7, 0) */,
  32'h3f2521d3 /* (5, 7, 0) */,
  32'h3ea04e75 /* (1, 7, 0) */,
  32'h3e960c85 /* (13, 3, 0) */,
  32'h3ecb578e /* (9, 3, 0) */,
  32'h3ea49cf9 /* (5, 3, 0) */,
  32'h3eb78ea1 /* (1, 3, 0) */,
  32'h3ea63161 /* (12, 15, 12) */,
  32'h3eebb725 /* (8, 15, 12) */,
  32'h3ea63161 /* (4, 15, 12) */,
  32'h3e962cf4 /* (0, 15, 12) */,
  32'h3f12b00d /* (12, 11, 12) */,
  32'h3f8a9c45 /* (8, 11, 12) */,
  32'h3f12b00d /* (4, 11, 12) */,
  32'h3ebddc83 /* (0, 11, 12) */,
  32'h3f59849a /* (12, 7, 12) */,
  32'h3fedbe1f /* (8, 7, 12) */,
  32'h3f59849a /* (4, 7, 12) */,
  32'h3efc5be6 /* (0, 7, 12) */,
  32'h3ec4d2c5 /* (12, 3, 12) */,
  32'h3f1dd43f /* (8, 3, 12) */,
  32'h3ec4d2c5 /* (4, 3, 12) */,
  32'h3e964277 /* (0, 3, 12) */,
  32'h3eebb725 /* (12, 15, 8) */,
  32'h3f80d0e8 /* (8, 15, 8) */,
  32'h3eebb725 /* (4, 15, 8) */,
  32'h3e88bc50 /* (0, 15, 8) */,
  32'h3f8a9c45 /* (12, 11, 8) */,
  32'h402594bb /* (8, 11, 8) */,
  32'h3f8a9c45 /* (4, 11, 8) */,
  32'h3f183f16 /* (0, 11, 8) */,
  32'h3fedbe1f /* (12, 7, 8) */,
  32'h4096cd97 /* (8, 7, 8) */,
  32'h3fedbe1f /* (4, 7, 8) */,
  32'h3f7cadff /* (0, 7, 8) */,
  32'h3f1dd43f /* (12, 3, 8) */,
  32'h3fb27927 /* (8, 3, 8) */,
  32'h3f1dd43f /* (4, 3, 8) */,
  32'h3eb32545 /* (0, 3, 8) */,
  32'h3ea63161 /* (12, 15, 4) */,
  32'h3eebb725 /* (8, 15, 4) */,
  32'h3ea63161 /* (4, 15, 4) */,
  32'h3e962cf4 /* (0, 15, 4) */,
  32'h3f12b00d /* (12, 11, 4) */,
  32'h3f8a9c45 /* (8, 11, 4) */,
  32'h3f12b00d /* (4, 11, 4) */,
  32'h3ebddc83 /* (0, 11, 4) */,
  32'h3f59849a /* (12, 7, 4) */,
  32'h3fedbe1f /* (8, 7, 4) */,
  32'h3f59849a /* (4, 7, 4) */,
  32'h3efc5be6 /* (0, 7, 4) */,
  32'h3ec4d2c5 /* (12, 3, 4) */,
  32'h3f1dd43f /* (8, 3, 4) */,
  32'h3ec4d2c5 /* (4, 3, 4) */,
  32'h3e964277 /* (0, 3, 4) */,
  32'h3e962cf4 /* (12, 15, 0) */,
  32'h3e88bc50 /* (8, 15, 0) */,
  32'h3e962cf4 /* (4, 15, 0) */,
  32'h40148d77 /* (0, 15, 0) */,
  32'h3ebddc83 /* (12, 11, 0) */,
  32'h3f183f16 /* (8, 11, 0) */,
  32'h3ebddc83 /* (4, 11, 0) */,
  32'h3e90f1d9 /* (0, 11, 0) */,
  32'h3efc5be6 /* (12, 7, 0) */,
  32'h3f7cadff /* (8, 7, 0) */,
  32'h3efc5be6 /* (4, 7, 0) */,
  32'h3e9bd51d /* (0, 7, 0) */,
  32'h3e964277 /* (12, 3, 0) */,
  32'h3eb32545 /* (8, 3, 0) */,
  32'h3e964277 /* (4, 3, 0) */,
  32'h3ec24b89 /* (0, 3, 0) */,
  32'h3e939519 /* (15, 14, 12) */,
  32'h3ed1ff4c /* (11, 14, 12) */,
  32'h3f104c25 /* (7, 14, 12) */,
  32'h3e9d3fef /* (3, 14, 12) */,
  32'h3ee9b2a2 /* (15, 10, 12) */,
  32'h3f753c17 /* (11, 10, 12) */,
  32'h3fc4fc22 /* (7, 10, 12) */,
  32'h3f15625b /* (3, 10, 12) */,
  32'h3ee9b2a2 /* (15, 6, 12) */,
  32'h3f753c17 /* (11, 6, 12) */,
  32'h3fc4fc22 /* (7, 6, 12) */,
  32'h3f15625b /* (3, 6, 12) */,
  32'h3e939519 /* (15, 2, 12) */,
  32'h3ed1ff4c /* (11, 2, 12) */,
  32'h3f104c25 /* (7, 2, 12) */,
  32'h3e9d3fef /* (3, 2, 12) */,
  32'h3e9c5e8a /* (15, 14, 8) */,
  32'h3f30df4f /* (11, 14, 8) */,
  32'h3f9420e3 /* (7, 14, 8) */,
  32'h3ece2dc1 /* (3, 14, 8) */,
  32'h3f5576ec /* (15, 10, 8) */,
  32'h40037a14 /* (11, 10, 8) */,
  32'h40686d0d /* (7, 10, 8) */,
  32'h3f91854a /* (3, 10, 8) */,
  32'h3f5576ec /* (15, 6, 8) */,
  32'h40037a14 /* (11, 6, 8) */,
  32'h40686d0d /* (7, 6, 8) */,
  32'h3f91854a /* (3, 6, 8) */,
  32'h3e9c5e8a /* (15, 2, 8) */,
  32'h3f30df4f /* (11, 2, 8) */,
  32'h3f9420e3 /* (7, 2, 8) */,
  32'h3ece2dc1 /* (3, 2, 8) */,
  32'h3e939519 /* (15, 14, 4) */,
  32'h3ed1ff4c /* (11, 14, 4) */,
  32'h3f104c25 /* (7, 14, 4) */,
  32'h3e9d3fef /* (3, 14, 4) */,
  32'h3ee9b2a2 /* (15, 10, 4) */,
  32'h3f753c17 /* (11, 10, 4) */,
  32'h3fc4fc22 /* (7, 10, 4) */,
  32'h3f15625b /* (3, 10, 4) */,
  32'h3ee9b2a2 /* (15, 6, 4) */,
  32'h3f753c17 /* (11, 6, 4) */,
  32'h3fc4fc22 /* (7, 6, 4) */,
  32'h3f15625b /* (3, 6, 4) */,
  32'h3e939519 /* (15, 2, 4) */,
  32'h3ed1ff4c /* (11, 2, 4) */,
  32'h3f104c25 /* (7, 2, 4) */,
  32'h3e9d3fef /* (3, 2, 4) */,
  32'h3f10451b /* (15, 14, 0) */,
  32'h3e97b006 /* (11, 14, 0) */,
  32'h3eaee5c8 /* (7, 14, 0) */,
  32'h3ea34ae8 /* (3, 14, 0) */,
  32'h3e9bd472 /* (15, 10, 0) */,
  32'h3f1019ab /* (11, 10, 0) */,
  32'h3f59ea43 /* (7, 10, 0) */,
  32'h3ebc86f4 /* (3, 10, 0) */,
  32'h3e9bd472 /* (15, 6, 0) */,
  32'h3f1019ab /* (11, 6, 0) */,
  32'h3f59ea43 /* (7, 6, 0) */,
  32'h3ebc86f4 /* (3, 6, 0) */,
  32'h3f10451b /* (15, 2, 0) */,
  32'h3e97b006 /* (11, 2, 0) */,
  32'h3eaee5c8 /* (7, 2, 0) */,
  32'h3ea34ae8 /* (3, 2, 0) */,
  32'h3e95577d /* (14, 14, 12) */,
  32'h3effc9dc /* (10, 14, 12) */,
  32'h3effc9dc /* (6, 14, 12) */,
  32'h3e95577d /* (2, 14, 12) */,
  32'h3effc9dc /* (14, 10, 12) */,
  32'h3fa2a180 /* (10, 10, 12) */,
  32'h3fa2a180 /* (6, 10, 12) */,
  32'h3effc9dc /* (2, 10, 12) */,
  32'h3effc9dc /* (14, 6, 12) */,
  32'h3fa2a180 /* (10, 6, 12) */,
  32'h3fa2a180 /* (6, 6, 12) */,
  32'h3effc9dc /* (2, 6, 12) */,
  32'h3e95577d /* (14, 2, 12) */,
  32'h3effc9dc /* (10, 2, 12) */,
  32'h3effc9dc /* (6, 2, 12) */,
  32'h3e95577d /* (2, 2, 12) */,
  32'h3ead4da0 /* (14, 14, 8) */,
  32'h3f6fbf1e /* (10, 14, 8) */,
  32'h3f6fbf1e /* (6, 14, 8) */,
  32'h3ead4da0 /* (2, 14, 8) */,
  32'h3f6fbf1e /* (14, 10, 8) */,
  32'h40372c7f /* (10, 10, 8) */,
  32'h40372c7f /* (6, 10, 8) */,
  32'h3f6fbf1e /* (2, 10, 8) */,
  32'h3f6fbf1e /* (14, 6, 8) */,
  32'h40372c7f /* (10, 6, 8) */,
  32'h40372c7f /* (6, 6, 8) */,
  32'h3f6fbf1e /* (2, 6, 8) */,
  32'h3ead4da0 /* (14, 2, 8) */,
  32'h3f6fbf1e /* (10, 2, 8) */,
  32'h3f6fbf1e /* (6, 2, 8) */,
  32'h3ead4da0 /* (2, 2, 8) */,
  32'h3e95577d /* (14, 14, 4) */,
  32'h3effc9dc /* (10, 14, 4) */,
  32'h3effc9dc /* (6, 14, 4) */,
  32'h3e95577d /* (2, 14, 4) */,
  32'h3effc9dc /* (14, 10, 4) */,
  32'h3fa2a180 /* (10, 10, 4) */,
  32'h3fa2a180 /* (6, 10, 4) */,
  32'h3effc9dc /* (2, 10, 4) */,
  32'h3effc9dc /* (14, 6, 4) */,
  32'h3fa2a180 /* (10, 6, 4) */,
  32'h3fa2a180 /* (6, 6, 4) */,
  32'h3effc9dc /* (2, 6, 4) */,
  32'h3e95577d /* (14, 2, 4) */,
  32'h3effc9dc /* (10, 2, 4) */,
  32'h3effc9dc /* (6, 2, 4) */,
  32'h3e95577d /* (2, 2, 4) */,
  32'h3ed08e8d /* (14, 14, 0) */,
  32'h3ea6b2c0 /* (10, 14, 0) */,
  32'h3ea6b2c0 /* (6, 14, 0) */,
  32'h3ed08e8d /* (2, 14, 0) */,
  32'h3ea6b2c0 /* (14, 10, 0) */,
  32'h3f390e8b /* (10, 10, 0) */,
  32'h3f390e8b /* (6, 10, 0) */,
  32'h3ea6b2c0 /* (2, 10, 0) */,
  32'h3ea6b2c0 /* (14, 6, 0) */,
  32'h3f390e8b /* (10, 6, 0) */,
  32'h3f390e8b /* (6, 6, 0) */,
  32'h3ea6b2c0 /* (2, 6, 0) */,
  32'h3ed08e8d /* (14, 2, 0) */,
  32'h3ea6b2c0 /* (10, 2, 0) */,
  32'h3ea6b2c0 /* (6, 2, 0) */,
  32'h3ed08e8d /* (2, 2, 0) */,
  32'h3e9d3fef /* (13, 14, 12) */,
  32'h3f104c25 /* (9, 14, 12) */,
  32'h3ed1ff4c /* (5, 14, 12) */,
  32'h3e939519 /* (1, 14, 12) */,
  32'h3f15625b /* (13, 10, 12) */,
  32'h3fc4fc22 /* (9, 10, 12) */,
  32'h3f753c17 /* (5, 10, 12) */,
  32'h3ee9b2a2 /* (1, 10, 12) */,
  32'h3f15625b /* (13, 6, 12) */,
  32'h3fc4fc22 /* (9, 6, 12) */,
  32'h3f753c17 /* (5, 6, 12) */,
  32'h3ee9b2a2 /* (1, 6, 12) */,
  32'h3e9d3fef /* (13, 2, 12) */,
  32'h3f104c25 /* (9, 2, 12) */,
  32'h3ed1ff4c /* (5, 2, 12) */,
  32'h3e939519 /* (1, 2, 12) */,
  32'h3ece2dc1 /* (13, 14, 8) */,
  32'h3f9420e3 /* (9, 14, 8) */,
  32'h3f30df4f /* (5, 14, 8) */,
  32'h3e9c5e8a /* (1, 14, 8) */,
  32'h3f91854a /* (13, 10, 8) */,
  32'h40686d0d /* (9, 10, 8) */,
  32'h40037a14 /* (5, 10, 8) */,
  32'h3f5576ec /* (1, 10, 8) */,
  32'h3f91854a /* (13, 6, 8) */,
  32'h40686d0d /* (9, 6, 8) */,
  32'h40037a14 /* (5, 6, 8) */,
  32'h3f5576ec /* (1, 6, 8) */,
  32'h3ece2dc1 /* (13, 2, 8) */,
  32'h3f9420e3 /* (9, 2, 8) */,
  32'h3f30df4f /* (5, 2, 8) */,
  32'h3e9c5e8a /* (1, 2, 8) */,
  32'h3e9d3fef /* (13, 14, 4) */,
  32'h3f104c25 /* (9, 14, 4) */,
  32'h3ed1ff4c /* (5, 14, 4) */,
  32'h3e939519 /* (1, 14, 4) */,
  32'h3f15625b /* (13, 10, 4) */,
  32'h3fc4fc22 /* (9, 10, 4) */,
  32'h3f753c17 /* (5, 10, 4) */,
  32'h3ee9b2a2 /* (1, 10, 4) */,
  32'h3f15625b /* (13, 6, 4) */,
  32'h3fc4fc22 /* (9, 6, 4) */,
  32'h3f753c17 /* (5, 6, 4) */,
  32'h3ee9b2a2 /* (1, 6, 4) */,
  32'h3e9d3fef /* (13, 2, 4) */,
  32'h3f104c25 /* (9, 2, 4) */,
  32'h3ed1ff4c /* (5, 2, 4) */,
  32'h3e939519 /* (1, 2, 4) */,
  32'h3ea34ae8 /* (13, 14, 0) */,
  32'h3eaee5c8 /* (9, 14, 0) */,
  32'h3e97b006 /* (5, 14, 0) */,
  32'h3f10451b /* (1, 14, 0) */,
  32'h3ebc86f4 /* (13, 10, 0) */,
  32'h3f59ea43 /* (9, 10, 0) */,
  32'h3f1019ab /* (5, 10, 0) */,
  32'h3e9bd472 /* (1, 10, 0) */,
  32'h3ebc86f4 /* (13, 6, 0) */,
  32'h3f59ea43 /* (9, 6, 0) */,
  32'h3f1019ab /* (5, 6, 0) */,
  32'h3e9bd472 /* (1, 6, 0) */,
  32'h3ea34ae8 /* (13, 2, 0) */,
  32'h3eaee5c8 /* (9, 2, 0) */,
  32'h3e97b006 /* (5, 2, 0) */,
  32'h3f10451b /* (1, 2, 0) */,
  32'h3eb02eb0 /* (12, 14, 12) */,
  32'h3f036eaf /* (8, 14, 12) */,
  32'h3eb02eb0 /* (4, 14, 12) */,
  32'h3e939fbd /* (0, 14, 12) */,
  32'h3f3a61a4 /* (12, 10, 12) */,
  32'h3fbe2ead /* (8, 10, 12) */,
  32'h3f3a61a4 /* (4, 10, 12) */,
  32'h3ee2e9d3 /* (0, 10, 12) */,
  32'h3f3a61a4 /* (12, 6, 12) */,
  32'h3fbe2ead /* (8, 6, 12) */,
  32'h3f3a61a4 /* (4, 6, 12) */,
  32'h3ee2e9d3 /* (0, 6, 12) */,
  32'h3eb02eb0 /* (12, 2, 12) */,
  32'h3f036eaf /* (8, 2, 12) */,
  32'h3eb02eb0 /* (4, 2, 12) */,
  32'h3e939fbd /* (0, 2, 12) */,
  32'h3f036eaf /* (12, 14, 8) */,
  32'h3f91966b /* (8, 14, 8) */,
  32'h3f036eaf /* (4, 14, 8) */,
  32'h3e9727de /* (0, 14, 8) */,
  32'h3fbe2ead /* (12, 10, 8) */,
  32'h406a2757 /* (8, 10, 8) */,
  32'h3fbe2ead /* (4, 10, 8) */,
  32'h3f4d63f0 /* (0, 10, 8) */,
  32'h3fbe2ead /* (12, 6, 8) */,
  32'h406a2757 /* (8, 6, 8) */,
  32'h3fbe2ead /* (4, 6, 8) */,
  32'h3f4d63f0 /* (0, 6, 8) */,
  32'h3f036eaf /* (12, 2, 8) */,
  32'h3f91966b /* (8, 2, 8) */,
  32'h3f036eaf /* (4, 2, 8) */,
  32'h3e9727de /* (0, 2, 8) */,
  32'h3eb02eb0 /* (12, 14, 4) */,
  32'h3f036eaf /* (8, 14, 4) */,
  32'h3eb02eb0 /* (4, 14, 4) */,
  32'h3e939fbd /* (0, 14, 4) */,
  32'h3f3a61a4 /* (12, 10, 4) */,
  32'h3fbe2ead /* (8, 10, 4) */,
  32'h3f3a61a4 /* (4, 10, 4) */,
  32'h3ee2e9d3 /* (0, 10, 4) */,
  32'h3f3a61a4 /* (12, 6, 4) */,
  32'h3fbe2ead /* (8, 6, 4) */,
  32'h3f3a61a4 /* (4, 6, 4) */,
  32'h3ee2e9d3 /* (0, 6, 4) */,
  32'h3eb02eb0 /* (12, 2, 4) */,
  32'h3f036eaf /* (8, 2, 4) */,
  32'h3eb02eb0 /* (4, 2, 4) */,
  32'h3e939fbd /* (0, 2, 4) */,
  32'h3e939fbd /* (12, 14, 0) */,
  32'h3e9727de /* (8, 14, 0) */,
  32'h3e939fbd /* (4, 14, 0) */,
  32'h3f2bcc5c /* (0, 14, 0) */,
  32'h3ee2e9d3 /* (12, 10, 0) */,
  32'h3f4d63f0 /* (8, 10, 0) */,
  32'h3ee2e9d3 /* (4, 10, 0) */,
  32'h3e989327 /* (0, 10, 0) */,
  32'h3ee2e9d3 /* (12, 6, 0) */,
  32'h3f4d63f0 /* (8, 6, 0) */,
  32'h3ee2e9d3 /* (4, 6, 0) */,
  32'h3e989327 /* (0, 6, 0) */,
  32'h3e939fbd /* (12, 2, 0) */,
  32'h3e9727de /* (8, 2, 0) */,
  32'h3e939fbd /* (4, 2, 0) */,
  32'h3f2bcc5c /* (0, 2, 0) */,
  32'h3e97a967 /* (15, 13, 12) */,
  32'h3ef076ff /* (11, 13, 12) */,
  32'h3f2b2ff1 /* (7, 13, 12) */,
  32'h3eaaa637 /* (3, 13, 12) */,
  32'h3f0271c0 /* (15, 9, 12) */,
  32'h3f91d65e /* (11, 9, 12) */,
  32'h3ff29d82 /* (7, 9, 12) */,
  32'h3f2b2ff1 /* (3, 9, 12) */,
  32'h3ec28d9a /* (15, 5, 12) */,
  32'h3f3cbfdf /* (11, 5, 12) */,
  32'h3f91d65e /* (7, 5, 12) */,
  32'h3ef076ff /* (3, 5, 12) */,
  32'h3e94e1d9 /* (15, 1, 12) */,
  32'h3ec28d9a /* (11, 1, 12) */,
  32'h3f0271c0 /* (7, 1, 12) */,
  32'h3e97a967 /* (3, 1, 12) */,
  32'h3eb9823a /* (15, 13, 8) */,
  32'h3f558e61 /* (11, 13, 8) */,
  32'h3fb4be0d /* (7, 13, 8) */,
  32'h3ef65451 /* (3, 13, 8) */,
  32'h3f8374c7 /* (15, 9, 8) */,
  32'h40258eba /* (11, 9, 8) */,
  32'h4094977b /* (7, 9, 8) */,
  32'h3fb4be0d /* (3, 9, 8) */,
  32'h3f1e09be /* (15, 5, 8) */,
  32'h3fbe36ae /* (11, 5, 8) */,
  32'h40258eba /* (7, 5, 8) */,
  32'h3f558e61 /* (3, 5, 8) */,
  32'h3e8d5b73 /* (15, 1, 8) */,
  32'h3f1e09be /* (11, 1, 8) */,
  32'h3f8374c7 /* (7, 1, 8) */,
  32'h3eb9823a /* (3, 1, 8) */,
  32'h3e97a967 /* (15, 13, 4) */,
  32'h3ef076ff /* (11, 13, 4) */,
  32'h3f2b2ff1 /* (7, 13, 4) */,
  32'h3eaaa637 /* (3, 13, 4) */,
  32'h3f0271c0 /* (15, 9, 4) */,
  32'h3f91d65e /* (11, 9, 4) */,
  32'h3ff29d82 /* (7, 9, 4) */,
  32'h3f2b2ff1 /* (3, 9, 4) */,
  32'h3ec28d9a /* (15, 5, 4) */,
  32'h3f3cbfdf /* (11, 5, 4) */,
  32'h3f91d65e /* (7, 5, 4) */,
  32'h3ef076ff /* (3, 5, 4) */,
  32'h3e94e1d9 /* (15, 1, 4) */,
  32'h3ec28d9a /* (11, 1, 4) */,
  32'h3f0271c0 /* (7, 1, 4) */,
  32'h3e97a967 /* (3, 1, 4) */,
  32'h3eb78ea1 /* (15, 13, 0) */,
  32'h3ea49cf9 /* (11, 13, 0) */,
  32'h3ecb578e /* (7, 13, 0) */,
  32'h3e960c85 /* (3, 13, 0) */,
  32'h3ea04e75 /* (15, 9, 0) */,
  32'h3f2521d3 /* (11, 9, 0) */,
  32'h3f836079 /* (7, 9, 0) */,
  32'h3ecb578e /* (3, 9, 0) */,
  32'h3e924c17 /* (15, 5, 0) */,
  32'h3ee7f590 /* (11, 5, 0) */,
  32'h3f2521d3 /* (7, 5, 0) */,
  32'h3ea49cf9 /* (3, 5, 0) */,
  32'h3f9befb2 /* (15, 1, 0) */,
  32'h3e924c17 /* (11, 1, 0) */,
  32'h3ea04e75 /* (7, 1, 0) */,
  32'h3eb78ea1 /* (3, 1, 0) */,
  32'h3e9d3fef /* (14, 13, 12) */,
  32'h3f15625b /* (10, 13, 12) */,
  32'h3f15625b /* (6, 13, 12) */,
  32'h3e9d3fef /* (2, 13, 12) */,
  32'h3f104c25 /* (14, 9, 12) */,
  32'h3fc4fc22 /* (10, 9, 12) */,
  32'h3fc4fc22 /* (6, 9, 12) */,
  32'h3f104c25 /* (2, 9, 12) */,
  32'h3ed1ff4c /* (14, 5, 12) */,
  32'h3f753c17 /* (10, 5, 12) */,
  32'h3f753c17 /* (6, 5, 12) */,
  32'h3ed1ff4c /* (2, 5, 12) */,
  32'h3e939519 /* (14, 1, 12) */,
  32'h3ee9b2a2 /* (10, 1, 12) */,
  32'h3ee9b2a2 /* (6, 1, 12) */,
  32'h3e939519 /* (2, 1, 12) */,
  32'h3ece2dc1 /* (14, 13, 8) */,
  32'h3f91854a /* (10, 13, 8) */,
  32'h3f91854a /* (6, 13, 8) */,
  32'h3ece2dc1 /* (2, 13, 8) */,
  32'h3f9420e3 /* (14, 9, 8) */,
  32'h40686d0d /* (10, 9, 8) */,
  32'h40686d0d /* (6, 9, 8) */,
  32'h3f9420e3 /* (2, 9, 8) */,
  32'h3f30df4f /* (14, 5, 8) */,
  32'h40037a14 /* (10, 5, 8) */,
  32'h40037a14 /* (6, 5, 8) */,
  32'h3f30df4f /* (2, 5, 8) */,
  32'h3e9c5e8a /* (14, 1, 8) */,
  32'h3f5576ec /* (10, 1, 8) */,
  32'h3f5576ec /* (6, 1, 8) */,
  32'h3e9c5e8a /* (2, 1, 8) */,
  32'h3e9d3fef /* (14, 13, 4) */,
  32'h3f15625b /* (10, 13, 4) */,
  32'h3f15625b /* (6, 13, 4) */,
  32'h3e9d3fef /* (2, 13, 4) */,
  32'h3f104c25 /* (14, 9, 4) */,
  32'h3fc4fc22 /* (10, 9, 4) */,
  32'h3fc4fc22 /* (6, 9, 4) */,
  32'h3f104c25 /* (2, 9, 4) */,
  32'h3ed1ff4c /* (14, 5, 4) */,
  32'h3f753c17 /* (10, 5, 4) */,
  32'h3f753c17 /* (6, 5, 4) */,
  32'h3ed1ff4c /* (2, 5, 4) */,
  32'h3e939519 /* (14, 1, 4) */,
  32'h3ee9b2a2 /* (10, 1, 4) */,
  32'h3ee9b2a2 /* (6, 1, 4) */,
  32'h3e939519 /* (2, 1, 4) */,
  32'h3ea34ae8 /* (14, 13, 0) */,
  32'h3ebc86f4 /* (10, 13, 0) */,
  32'h3ebc86f4 /* (6, 13, 0) */,
  32'h3ea34ae8 /* (2, 13, 0) */,
  32'h3eaee5c8 /* (14, 9, 0) */,
  32'h3f59ea43 /* (10, 9, 0) */,
  32'h3f59ea43 /* (6, 9, 0) */,
  32'h3eaee5c8 /* (2, 9, 0) */,
  32'h3e97b006 /* (14, 5, 0) */,
  32'h3f1019ab /* (10, 5, 0) */,
  32'h3f1019ab /* (6, 5, 0) */,
  32'h3e97b006 /* (2, 5, 0) */,
  32'h3f10451b /* (14, 1, 0) */,
  32'h3e9bd472 /* (10, 1, 0) */,
  32'h3e9bd472 /* (6, 1, 0) */,
  32'h3f10451b /* (2, 1, 0) */,
  32'h3eaaa637 /* (13, 13, 12) */,
  32'h3f2b2ff1 /* (9, 13, 12) */,
  32'h3ef076ff /* (5, 13, 12) */,
  32'h3e97a967 /* (1, 13, 12) */,
  32'h3f2b2ff1 /* (13, 9, 12) */,
  32'h3ff29d82 /* (9, 9, 12) */,
  32'h3f91d65e /* (5, 9, 12) */,
  32'h3f0271c0 /* (1, 9, 12) */,
  32'h3ef076ff /* (13, 5, 12) */,
  32'h3f91d65e /* (9, 5, 12) */,
  32'h3f3cbfdf /* (5, 5, 12) */,
  32'h3ec28d9a /* (1, 5, 12) */,
  32'h3e97a967 /* (13, 1, 12) */,
  32'h3f0271c0 /* (9, 1, 12) */,
  32'h3ec28d9a /* (5, 1, 12) */,
  32'h3e94e1d9 /* (1, 1, 12) */,
  32'h3ef65451 /* (13, 13, 8) */,
  32'h3fb4be0d /* (9, 13, 8) */,
  32'h3f558e61 /* (5, 13, 8) */,
  32'h3eb9823a /* (1, 13, 8) */,
  32'h3fb4be0d /* (13, 9, 8) */,
  32'h4094977b /* (9, 9, 8) */,
  32'h40258eba /* (5, 9, 8) */,
  32'h3f8374c7 /* (1, 9, 8) */,
  32'h3f558e61 /* (13, 5, 8) */,
  32'h40258eba /* (9, 5, 8) */,
  32'h3fbe36ae /* (5, 5, 8) */,
  32'h3f1e09be /* (1, 5, 8) */,
  32'h3eb9823a /* (13, 1, 8) */,
  32'h3f8374c7 /* (9, 1, 8) */,
  32'h3f1e09be /* (5, 1, 8) */,
  32'h3e8d5b73 /* (1, 1, 8) */,
  32'h3eaaa637 /* (13, 13, 4) */,
  32'h3f2b2ff1 /* (9, 13, 4) */,
  32'h3ef076ff /* (5, 13, 4) */,
  32'h3e97a967 /* (1, 13, 4) */,
  32'h3f2b2ff1 /* (13, 9, 4) */,
  32'h3ff29d82 /* (9, 9, 4) */,
  32'h3f91d65e /* (5, 9, 4) */,
  32'h3f0271c0 /* (1, 9, 4) */,
  32'h3ef076ff /* (13, 5, 4) */,
  32'h3f91d65e /* (9, 5, 4) */,
  32'h3f3cbfdf /* (5, 5, 4) */,
  32'h3ec28d9a /* (1, 5, 4) */,
  32'h3e97a967 /* (13, 1, 4) */,
  32'h3f0271c0 /* (9, 1, 4) */,
  32'h3ec28d9a /* (5, 1, 4) */,
  32'h3e94e1d9 /* (1, 1, 4) */,
  32'h3e960c85 /* (13, 13, 0) */,
  32'h3ecb578e /* (9, 13, 0) */,
  32'h3ea49cf9 /* (5, 13, 0) */,
  32'h3eb78ea1 /* (1, 13, 0) */,
  32'h3ecb578e /* (13, 9, 0) */,
  32'h3f836079 /* (9, 9, 0) */,
  32'h3f2521d3 /* (5, 9, 0) */,
  32'h3ea04e75 /* (1, 9, 0) */,
  32'h3ea49cf9 /* (13, 5, 0) */,
  32'h3f2521d3 /* (9, 5, 0) */,
  32'h3ee7f590 /* (5, 5, 0) */,
  32'h3e924c17 /* (1, 5, 0) */,
  32'h3eb78ea1 /* (13, 1, 0) */,
  32'h3ea04e75 /* (9, 1, 0) */,
  32'h3e924c17 /* (5, 1, 0) */,
  32'h3f9befb2 /* (1, 1, 0) */,
  32'h3ec4d2c5 /* (12, 13, 12) */,
  32'h3f1dd43f /* (8, 13, 12) */,
  32'h3ec4d2c5 /* (4, 13, 12) */,
  32'h3e964277 /* (0, 13, 12) */,
  32'h3f59849a /* (12, 9, 12) */,
  32'h3fedbe1f /* (8, 9, 12) */,
  32'h3f59849a /* (4, 9, 12) */,
  32'h3efc5be6 /* (0, 9, 12) */,
  32'h3f12b00d /* (12, 5, 12) */,
  32'h3f8a9c45 /* (8, 5, 12) */,
  32'h3f12b00d /* (4, 5, 12) */,
  32'h3ebddc83 /* (0, 5, 12) */,
  32'h3ea63161 /* (12, 1, 12) */,
  32'h3eebb725 /* (8, 1, 12) */,
  32'h3ea63161 /* (4, 1, 12) */,
  32'h3e962cf4 /* (0, 1, 12) */,
  32'h3f1dd43f /* (12, 13, 8) */,
  32'h3fb27927 /* (8, 13, 8) */,
  32'h3f1dd43f /* (4, 13, 8) */,
  32'h3eb32545 /* (0, 13, 8) */,
  32'h3fedbe1f /* (12, 9, 8) */,
  32'h4096cd97 /* (8, 9, 8) */,
  32'h3fedbe1f /* (4, 9, 8) */,
  32'h3f7cadff /* (0, 9, 8) */,
  32'h3f8a9c45 /* (12, 5, 8) */,
  32'h402594bb /* (8, 5, 8) */,
  32'h3f8a9c45 /* (4, 5, 8) */,
  32'h3f183f16 /* (0, 5, 8) */,
  32'h3eebb725 /* (12, 1, 8) */,
  32'h3f80d0e8 /* (8, 1, 8) */,
  32'h3eebb725 /* (4, 1, 8) */,
  32'h3e88bc50 /* (0, 1, 8) */,
  32'h3ec4d2c5 /* (12, 13, 4) */,
  32'h3f1dd43f /* (8, 13, 4) */,
  32'h3ec4d2c5 /* (4, 13, 4) */,
  32'h3e964277 /* (0, 13, 4) */,
  32'h3f59849a /* (12, 9, 4) */,
  32'h3fedbe1f /* (8, 9, 4) */,
  32'h3f59849a /* (4, 9, 4) */,
  32'h3efc5be6 /* (0, 9, 4) */,
  32'h3f12b00d /* (12, 5, 4) */,
  32'h3f8a9c45 /* (8, 5, 4) */,
  32'h3f12b00d /* (4, 5, 4) */,
  32'h3ebddc83 /* (0, 5, 4) */,
  32'h3ea63161 /* (12, 1, 4) */,
  32'h3eebb725 /* (8, 1, 4) */,
  32'h3ea63161 /* (4, 1, 4) */,
  32'h3e962cf4 /* (0, 1, 4) */,
  32'h3e964277 /* (12, 13, 0) */,
  32'h3eb32545 /* (8, 13, 0) */,
  32'h3e964277 /* (4, 13, 0) */,
  32'h3ec24b89 /* (0, 13, 0) */,
  32'h3efc5be6 /* (12, 9, 0) */,
  32'h3f7cadff /* (8, 9, 0) */,
  32'h3efc5be6 /* (4, 9, 0) */,
  32'h3e9bd51d /* (0, 9, 0) */,
  32'h3ebddc83 /* (12, 5, 0) */,
  32'h3f183f16 /* (8, 5, 0) */,
  32'h3ebddc83 /* (4, 5, 0) */,
  32'h3e90f1d9 /* (0, 5, 0) */,
  32'h3e962cf4 /* (12, 1, 0) */,
  32'h3e88bc50 /* (8, 1, 0) */,
  32'h3e962cf4 /* (4, 1, 0) */,
  32'h40148d77 /* (0, 1, 0) */,
  32'h3ea63161 /* (15, 12, 12) */,
  32'h3f12b00d /* (11, 12, 12) */,
  32'h3f59849a /* (7, 12, 12) */,
  32'h3ec4d2c5 /* (3, 12, 12) */,
  32'h3eebb725 /* (15, 8, 12) */,
  32'h3f8a9c45 /* (11, 8, 12) */,
  32'h3fedbe1f /* (7, 8, 12) */,
  32'h3f1dd43f /* (3, 8, 12) */,
  32'h3ea63161 /* (15, 4, 12) */,
  32'h3f12b00d /* (11, 4, 12) */,
  32'h3f59849a /* (7, 4, 12) */,
  32'h3ec4d2c5 /* (3, 4, 12) */,
  32'h3e962cf4 /* (15, 0, 12) */,
  32'h3ebddc83 /* (11, 0, 12) */,
  32'h3efc5be6 /* (7, 0, 12) */,
  32'h3e964277 /* (3, 0, 12) */,
  32'h3eebb725 /* (15, 12, 8) */,
  32'h3f8a9c45 /* (11, 12, 8) */,
  32'h3fedbe1f /* (7, 12, 8) */,
  32'h3f1dd43f /* (3, 12, 8) */,
  32'h3f80d0e8 /* (15, 8, 8) */,
  32'h402594bb /* (11, 8, 8) */,
  32'h4096cd97 /* (7, 8, 8) */,
  32'h3fb27927 /* (3, 8, 8) */,
  32'h3eebb725 /* (15, 4, 8) */,
  32'h3f8a9c45 /* (11, 4, 8) */,
  32'h3fedbe1f /* (7, 4, 8) */,
  32'h3f1dd43f /* (3, 4, 8) */,
  32'h3e88bc50 /* (15, 0, 8) */,
  32'h3f183f16 /* (11, 0, 8) */,
  32'h3f7cadff /* (7, 0, 8) */,
  32'h3eb32545 /* (3, 0, 8) */,
  32'h3ea63161 /* (15, 12, 4) */,
  32'h3f12b00d /* (11, 12, 4) */,
  32'h3f59849a /* (7, 12, 4) */,
  32'h3ec4d2c5 /* (3, 12, 4) */,
  32'h3eebb725 /* (15, 8, 4) */,
  32'h3f8a9c45 /* (11, 8, 4) */,
  32'h3fedbe1f /* (7, 8, 4) */,
  32'h3f1dd43f /* (3, 8, 4) */,
  32'h3ea63161 /* (15, 4, 4) */,
  32'h3f12b00d /* (11, 4, 4) */,
  32'h3f59849a /* (7, 4, 4) */,
  32'h3ec4d2c5 /* (3, 4, 4) */,
  32'h3e962cf4 /* (15, 0, 4) */,
  32'h3ebddc83 /* (11, 0, 4) */,
  32'h3efc5be6 /* (7, 0, 4) */,
  32'h3e964277 /* (3, 0, 4) */,
  32'h3e962cf4 /* (15, 12, 0) */,
  32'h3ebddc83 /* (11, 12, 0) */,
  32'h3efc5be6 /* (7, 12, 0) */,
  32'h3e964277 /* (3, 12, 0) */,
  32'h3e88bc50 /* (15, 8, 0) */,
  32'h3f183f16 /* (11, 8, 0) */,
  32'h3f7cadff /* (7, 8, 0) */,
  32'h3eb32545 /* (3, 8, 0) */,
  32'h3e962cf4 /* (15, 4, 0) */,
  32'h3ebddc83 /* (11, 4, 0) */,
  32'h3efc5be6 /* (7, 4, 0) */,
  32'h3e964277 /* (3, 4, 0) */,
  32'h40148d77 /* (15, 0, 0) */,
  32'h3e90f1d9 /* (11, 0, 0) */,
  32'h3e9bd51d /* (7, 0, 0) */,
  32'h3ec24b89 /* (3, 0, 0) */,
  32'h3eb02eb0 /* (14, 12, 12) */,
  32'h3f3a61a4 /* (10, 12, 12) */,
  32'h3f3a61a4 /* (6, 12, 12) */,
  32'h3eb02eb0 /* (2, 12, 12) */,
  32'h3f036eaf /* (14, 8, 12) */,
  32'h3fbe2ead /* (10, 8, 12) */,
  32'h3fbe2ead /* (6, 8, 12) */,
  32'h3f036eaf /* (2, 8, 12) */,
  32'h3eb02eb0 /* (14, 4, 12) */,
  32'h3f3a61a4 /* (10, 4, 12) */,
  32'h3f3a61a4 /* (6, 4, 12) */,
  32'h3eb02eb0 /* (2, 4, 12) */,
  32'h3e939fbd /* (14, 0, 12) */,
  32'h3ee2e9d3 /* (10, 0, 12) */,
  32'h3ee2e9d3 /* (6, 0, 12) */,
  32'h3e939fbd /* (2, 0, 12) */,
  32'h3f036eaf /* (14, 12, 8) */,
  32'h3fbe2ead /* (10, 12, 8) */,
  32'h3fbe2ead /* (6, 12, 8) */,
  32'h3f036eaf /* (2, 12, 8) */,
  32'h3f91966b /* (14, 8, 8) */,
  32'h406a2757 /* (10, 8, 8) */,
  32'h406a2757 /* (6, 8, 8) */,
  32'h3f91966b /* (2, 8, 8) */,
  32'h3f036eaf /* (14, 4, 8) */,
  32'h3fbe2ead /* (10, 4, 8) */,
  32'h3fbe2ead /* (6, 4, 8) */,
  32'h3f036eaf /* (2, 4, 8) */,
  32'h3e9727de /* (14, 0, 8) */,
  32'h3f4d63f0 /* (10, 0, 8) */,
  32'h3f4d63f0 /* (6, 0, 8) */,
  32'h3e9727de /* (2, 0, 8) */,
  32'h3eb02eb0 /* (14, 12, 4) */,
  32'h3f3a61a4 /* (10, 12, 4) */,
  32'h3f3a61a4 /* (6, 12, 4) */,
  32'h3eb02eb0 /* (2, 12, 4) */,
  32'h3f036eaf /* (14, 8, 4) */,
  32'h3fbe2ead /* (10, 8, 4) */,
  32'h3fbe2ead /* (6, 8, 4) */,
  32'h3f036eaf /* (2, 8, 4) */,
  32'h3eb02eb0 /* (14, 4, 4) */,
  32'h3f3a61a4 /* (10, 4, 4) */,
  32'h3f3a61a4 /* (6, 4, 4) */,
  32'h3eb02eb0 /* (2, 4, 4) */,
  32'h3e939fbd /* (14, 0, 4) */,
  32'h3ee2e9d3 /* (10, 0, 4) */,
  32'h3ee2e9d3 /* (6, 0, 4) */,
  32'h3e939fbd /* (2, 0, 4) */,
  32'h3e939fbd /* (14, 12, 0) */,
  32'h3ee2e9d3 /* (10, 12, 0) */,
  32'h3ee2e9d3 /* (6, 12, 0) */,
  32'h3e939fbd /* (2, 12, 0) */,
  32'h3e9727de /* (14, 8, 0) */,
  32'h3f4d63f0 /* (10, 8, 0) */,
  32'h3f4d63f0 /* (6, 8, 0) */,
  32'h3e9727de /* (2, 8, 0) */,
  32'h3e939fbd /* (14, 4, 0) */,
  32'h3ee2e9d3 /* (10, 4, 0) */,
  32'h3ee2e9d3 /* (6, 4, 0) */,
  32'h3e939fbd /* (2, 4, 0) */,
  32'h3f2bcc5c /* (14, 0, 0) */,
  32'h3e989327 /* (10, 0, 0) */,
  32'h3e989327 /* (6, 0, 0) */,
  32'h3f2bcc5c /* (2, 0, 0) */,
  32'h3ec4d2c5 /* (13, 12, 12) */,
  32'h3f59849a /* (9, 12, 12) */,
  32'h3f12b00d /* (5, 12, 12) */,
  32'h3ea63161 /* (1, 12, 12) */,
  32'h3f1dd43f /* (13, 8, 12) */,
  32'h3fedbe1f /* (9, 8, 12) */,
  32'h3f8a9c45 /* (5, 8, 12) */,
  32'h3eebb725 /* (1, 8, 12) */,
  32'h3ec4d2c5 /* (13, 4, 12) */,
  32'h3f59849a /* (9, 4, 12) */,
  32'h3f12b00d /* (5, 4, 12) */,
  32'h3ea63161 /* (1, 4, 12) */,
  32'h3e964277 /* (13, 0, 12) */,
  32'h3efc5be6 /* (9, 0, 12) */,
  32'h3ebddc83 /* (5, 0, 12) */,
  32'h3e962cf4 /* (1, 0, 12) */,
  32'h3f1dd43f /* (13, 12, 8) */,
  32'h3fedbe1f /* (9, 12, 8) */,
  32'h3f8a9c45 /* (5, 12, 8) */,
  32'h3eebb725 /* (1, 12, 8) */,
  32'h3fb27927 /* (13, 8, 8) */,
  32'h4096cd97 /* (9, 8, 8) */,
  32'h402594bb /* (5, 8, 8) */,
  32'h3f80d0e8 /* (1, 8, 8) */,
  32'h3f1dd43f /* (13, 4, 8) */,
  32'h3fedbe1f /* (9, 4, 8) */,
  32'h3f8a9c45 /* (5, 4, 8) */,
  32'h3eebb725 /* (1, 4, 8) */,
  32'h3eb32545 /* (13, 0, 8) */,
  32'h3f7cadff /* (9, 0, 8) */,
  32'h3f183f16 /* (5, 0, 8) */,
  32'h3e88bc50 /* (1, 0, 8) */,
  32'h3ec4d2c5 /* (13, 12, 4) */,
  32'h3f59849a /* (9, 12, 4) */,
  32'h3f12b00d /* (5, 12, 4) */,
  32'h3ea63161 /* (1, 12, 4) */,
  32'h3f1dd43f /* (13, 8, 4) */,
  32'h3fedbe1f /* (9, 8, 4) */,
  32'h3f8a9c45 /* (5, 8, 4) */,
  32'h3eebb725 /* (1, 8, 4) */,
  32'h3ec4d2c5 /* (13, 4, 4) */,
  32'h3f59849a /* (9, 4, 4) */,
  32'h3f12b00d /* (5, 4, 4) */,
  32'h3ea63161 /* (1, 4, 4) */,
  32'h3e964277 /* (13, 0, 4) */,
  32'h3efc5be6 /* (9, 0, 4) */,
  32'h3ebddc83 /* (5, 0, 4) */,
  32'h3e962cf4 /* (1, 0, 4) */,
  32'h3e964277 /* (13, 12, 0) */,
  32'h3efc5be6 /* (9, 12, 0) */,
  32'h3ebddc83 /* (5, 12, 0) */,
  32'h3e962cf4 /* (1, 12, 0) */,
  32'h3eb32545 /* (13, 8, 0) */,
  32'h3f7cadff /* (9, 8, 0) */,
  32'h3f183f16 /* (5, 8, 0) */,
  32'h3e88bc50 /* (1, 8, 0) */,
  32'h3e964277 /* (13, 4, 0) */,
  32'h3efc5be6 /* (9, 4, 0) */,
  32'h3ebddc83 /* (5, 4, 0) */,
  32'h3e962cf4 /* (1, 4, 0) */,
  32'h3ec24b89 /* (13, 0, 0) */,
  32'h3e9bd51d /* (9, 0, 0) */,
  32'h3e90f1d9 /* (5, 0, 0) */,
  32'h40148d77 /* (1, 0, 0) */,
  32'h3ee9d3eb /* (12, 12, 12) */,
  32'h3f4b8235 /* (8, 12, 12) */,
  32'h3ee9d3eb /* (4, 12, 12) */,
  32'h3ea34567 /* (0, 12, 12) */,
  32'h3f4b8235 /* (12, 8, 12) */,
  32'h3fec2938 /* (8, 8, 12) */,
  32'h3f4b8235 /* (4, 8, 12) */,
  32'h3ee35c6b /* (0, 8, 12) */,
  32'h3ee9d3eb /* (12, 4, 12) */,
  32'h3f4b8235 /* (8, 4, 12) */,
  32'h3ee9d3eb /* (4, 4, 12) */,
  32'h3ea34567 /* (0, 4, 12) */,
  32'h3ea34567 /* (12, 0, 12) */,
  32'h3ee35c6b /* (8, 0, 12) */,
  32'h3ea34567 /* (4, 0, 12) */,
  32'h3e980196 /* (0, 0, 12) */,
  32'h3f4b8235 /* (12, 12, 8) */,
  32'h3fec2938 /* (8, 12, 8) */,
  32'h3f4b8235 /* (4, 12, 8) */,
  32'h3ee35c6b /* (0, 12, 8) */,
  32'h3fec2938 /* (12, 8, 8) */,
  32'h409a278b /* (8, 8, 8) */,
  32'h3fec2938 /* (4, 8, 8) */,
  32'h3f7759b5 /* (0, 8, 8) */,
  32'h3f4b8235 /* (12, 4, 8) */,
  32'h3fec2938 /* (8, 4, 8) */,
  32'h3f4b8235 /* (4, 4, 8) */,
  32'h3ee35c6b /* (0, 4, 8) */,
  32'h3ee35c6b /* (12, 0, 8) */,
  32'h3f7759b5 /* (8, 0, 8) */,
  32'h3ee35c6b /* (4, 0, 8) */,
  32'h3e844bdf /* (0, 0, 8) */,
  32'h3ee9d3eb /* (12, 12, 4) */,
  32'h3f4b8235 /* (8, 12, 4) */,
  32'h3ee9d3eb /* (4, 12, 4) */,
  32'h3ea34567 /* (0, 12, 4) */,
  32'h3f4b8235 /* (12, 8, 4) */,
  32'h3fec2938 /* (8, 8, 4) */,
  32'h3f4b8235 /* (4, 8, 4) */,
  32'h3ee35c6b /* (0, 8, 4) */,
  32'h3ee9d3eb /* (12, 4, 4) */,
  32'h3f4b8235 /* (8, 4, 4) */,
  32'h3ee9d3eb /* (4, 4, 4) */,
  32'h3ea34567 /* (0, 4, 4) */,
  32'h3ea34567 /* (12, 0, 4) */,
  32'h3ee35c6b /* (8, 0, 4) */,
  32'h3ea34567 /* (4, 0, 4) */,
  32'h3e980196 /* (0, 0, 4) */,
  32'h3ea34567 /* (12, 12, 0) */,
  32'h3ee35c6b /* (8, 12, 0) */,
  32'h3ea34567 /* (4, 12, 0) */,
  32'h3e980196 /* (0, 12, 0) */,
  32'h3ee35c6b /* (12, 8, 0) */,
  32'h3f7759b5 /* (8, 8, 0) */,
  32'h3ee35c6b /* (4, 8, 0) */,
  32'h3e844bdf /* (0, 8, 0) */,
  32'h3ea34567 /* (12, 4, 0) */,
  32'h3ee35c6b /* (8, 4, 0) */,
  32'h3ea34567 /* (4, 4, 0) */,
  32'h3e980196 /* (0, 4, 0) */,
  32'h3e980196 /* (12, 0, 0) */,
  32'h3e844bdf /* (8, 0, 0) */,
  32'h3e980196 /* (4, 0, 0) */,
  32'h46c4597c /* (0, 0, 0) */};
